/**
 * Editor : 
 * File : fc_top.v
 */
module fc_top(

);


endmodule