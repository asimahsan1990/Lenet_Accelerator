
module fsm ( clk, srstn, conv_start, conv1_done, conv_done, mode, mem_sel );
  output [1:0] mode;
  input clk, srstn, conv_start, conv1_done, conv_done;
  output mem_sel;
  wire   n_mode_1_, n_mem_sel, n3, n5, n6, n9, n7, n8, n10;

  DFFSSRX1_HVT mode_reg_1_ ( .D(1'b0), .SETB(n6), .RSTB(n_mode_1_), .CLK(clk), 
        .Q(mode[1]), .QN(n8) );
  DFFSSRX1_HVT mem_sel_reg ( .D(n_mem_sel), .SETB(srstn), .RSTB(1'b1), .CLK(
        clk), .Q(mem_sel), .QN(n7) );
  DFFSSRX1_HVT mode_reg_0_ ( .D(n3), .SETB(n9), .RSTB(srstn), .CLK(clk), .Q(
        mode[0]), .QN(n5) );
  INVX0_HVT U3 ( .A(srstn), .Y(n6) );
  OA222X1_HVT U4 ( .A1(mode[1]), .A2(conv1_done), .A3(mode[1]), .A4(mode[0]), 
        .A5(n5), .A6(n8), .Y(n_mode_1_) );
  AND3X1_HVT U5 ( .A1(mode[1]), .A2(n5), .A3(conv_done), .Y(n3) );
  INVX1_HVT U6 ( .A(conv_start), .Y(n10) );
  AO22X1_HVT U7 ( .A1(conv_start), .A2(n7), .A3(n10), .A4(mem_sel), .Y(
        n_mem_sel) );
  AO221X1_HVT U8 ( .A1(n5), .A2(n10), .A3(mode[0]), .A4(conv1_done), .A5(
        mode[1]), .Y(n9) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_0 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n1;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n1), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n1) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_26 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_25 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_24 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_23 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_22 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_21 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_20 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_19 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_18 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_17 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_16 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_15 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_14 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_13 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_12 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_11 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_10 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_9 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_8 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_7 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_6 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_5 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_4 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_3 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_2 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_1 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19688, n2;

  AND2X1_HVT main_gate ( .A1(net19688), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19688) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module conv_control ( clk, srstn, mode, mem_sel, conv1_done, sram_raddr_weight, 
        box_sel, load_conv1_bias_enable, conv1_bias_set, sram_raddr_a0, 
        sram_raddr_a1, sram_raddr_a2, sram_raddr_a3, sram_raddr_a4, 
        sram_raddr_a5, sram_raddr_a6, sram_raddr_a7, sram_raddr_a8, 
        sram_write_enable_b0, sram_write_enable_b1, sram_write_enable_b2, 
        sram_write_enable_b3, sram_write_enable_b4, sram_write_enable_b5, 
        sram_write_enable_b6, sram_write_enable_b7, sram_write_enable_b8, 
        sram_bytemask_b, sram_waddr_b, conv_done, channel, set, 
        load_conv2_bias0_enable, load_conv2_bias1_enable, sram_raddr_b0, 
        sram_raddr_b1, sram_raddr_b2, sram_raddr_b3, sram_raddr_b4, 
        sram_raddr_b5, sram_raddr_b6, sram_raddr_b7, sram_raddr_b8, 
        sram_write_enable_c0, sram_write_enable_c1, sram_write_enable_c2, 
        sram_write_enable_c3, sram_write_enable_c4, sram_bytemask_c, 
        sram_waddr_c, sram_write_enable_d0, sram_write_enable_d1, 
        sram_write_enable_d2, sram_write_enable_d3, sram_write_enable_d4, 
        sram_bytemask_d, sram_waddr_d );
  input [1:0] mode;
  output [16:0] sram_raddr_weight;
  output [3:0] box_sel;
  output [16:0] conv1_bias_set;
  output [9:0] sram_raddr_a0;
  output [9:0] sram_raddr_a1;
  output [9:0] sram_raddr_a2;
  output [9:0] sram_raddr_a3;
  output [9:0] sram_raddr_a4;
  output [9:0] sram_raddr_a5;
  output [9:0] sram_raddr_a6;
  output [9:0] sram_raddr_a7;
  output [9:0] sram_raddr_a8;
  output [3:0] sram_bytemask_b;
  output [9:0] sram_waddr_b;
  output [4:0] channel;
  output [7:0] set;
  output [9:0] sram_raddr_b0;
  output [9:0] sram_raddr_b1;
  output [9:0] sram_raddr_b2;
  output [9:0] sram_raddr_b3;
  output [9:0] sram_raddr_b4;
  output [9:0] sram_raddr_b5;
  output [9:0] sram_raddr_b6;
  output [9:0] sram_raddr_b7;
  output [9:0] sram_raddr_b8;
  output [3:0] sram_bytemask_c;
  output [9:0] sram_waddr_c;
  output [3:0] sram_bytemask_d;
  output [9:0] sram_waddr_d;
  input clk, srstn, mem_sel;
  output conv1_done, load_conv1_bias_enable, sram_write_enable_b0,
         sram_write_enable_b1, sram_write_enable_b2, sram_write_enable_b3,
         sram_write_enable_b4, sram_write_enable_b5, sram_write_enable_b6,
         sram_write_enable_b7, sram_write_enable_b8, conv_done,
         load_conv2_bias0_enable, load_conv2_bias1_enable,
         sram_write_enable_c0, sram_write_enable_c1, sram_write_enable_c2,
         sram_write_enable_c3, sram_write_enable_c4, sram_write_enable_d0,
         sram_write_enable_d1, sram_write_enable_d2, sram_write_enable_d3,
         sram_write_enable_d4;
  wire   n_conv1_done, n_conv_done, conv1_weight_done, conv2_weight_done,
         delay2_write_enable, delay_load_conv1_bias_enable,
         delay_load_conv2_bias0_enable, delay_load_conv2_bias1_enable,
         load_data_enable, delay4_conv1_done, delay3_conv_done,
         delay2_addr_change_2_, n_conv1_weight_done, n_write_enable,
         write_enable, delay_write_enable, n_load_data_enable, n_box_sel_1_,
         n_addr_row_sel_cnt_0_, delay1_conv1_done, delay2_conv1_done,
         delay3_conv1_done, delay_conv_done, delay2_conv_done,
         delay_sram_write_enable_b0, delay_sram_write_enable_b1,
         delay_sram_write_enable_b2, delay_sram_write_enable_b3,
         delay_sram_write_enable_b4, delay_sram_write_enable_b5,
         delay_sram_write_enable_b6, delay_sram_write_enable_b7,
         delay_sram_write_enable_b8, delay2_sram_write_enable_b0,
         delay2_sram_write_enable_b1, delay2_sram_write_enable_b2,
         delay2_sram_write_enable_b3, delay2_sram_write_enable_b4,
         delay2_sram_write_enable_b5, delay2_sram_write_enable_b6,
         delay2_sram_write_enable_b7, delay2_sram_write_enable_b8,
         n_sram_write_enable_b0, n_sram_write_enable_b1,
         n_sram_write_enable_b2, n_sram_write_enable_b3,
         n_sram_write_enable_b4, n_sram_write_enable_b5,
         n_sram_write_enable_b6, n_sram_write_enable_b7,
         n_sram_write_enable_b8, delay_sram_write_enable_c0,
         delay_sram_write_enable_c1, delay_sram_write_enable_c2,
         delay_sram_write_enable_c3, delay_sram_write_enable_c4,
         delay_sram_write_enable_d0, delay_sram_write_enable_d1,
         delay_sram_write_enable_d2, delay_sram_write_enable_d3,
         delay_sram_write_enable_d4, n_sram_write_enable_c0,
         n_sram_write_enable_c1, n_sram_write_enable_c2,
         n_sram_write_enable_c3, n_sram_write_enable_c4,
         n_sram_write_enable_d0, n_sram_write_enable_d1,
         n_sram_write_enable_d2, n_sram_write_enable_d3,
         n_sram_write_enable_d4, N2888, net19513, net19699, net19704, net19709,
         net19714, net19715, net19718, net19723, net19752, net19759, net19766,
         net19773, net19780, net19787, net19794, net19808, net19815, net19818,
         net19836, net19843, net19850, net19857, net19871, net19878, net19885,
         net19899, net19913, net19916, net19921, net19924, net19927, net19930,
         net19933, net19936, net19939, net19942, net19945, net19948, net19951,
         net19954, net19959, net19961, net19962, net19963, net19964, net19965,
         net19966, net19967, net19968, net19969, net19970, net19973, net19977,
         net19978, net19979, net19980, net19981, net19982, net19983, net19984,
         net19985, net19986, net19989, net19993, net19994, net19995, net19996,
         net19997, net19998, net20001, net20004, net20006, net20007, net20008,
         net20009, net20010, net20013, net20494, net20939, net20953, net21376,
         net21821, net22266, net22280, net22703, net23149, net23595, net23610,
         net24033, net24567, net25082, net25597, net26112, net26627, net27142,
         net27657, net28172, net28264, net28687, n459, n460, n462, n487, n1108,
         n1109, n1135, n1136, n1137, n1143, n1145, n1146, n1152, n1153, n1723,
         n1730, n1735, n1737, n1738, n1739, n2, n3, n4, n6, n7, n9, n11, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n23, n24, n26, n27, n29, n30,
         n32, n35, n36, n37, n39, n42, n43, n44, n45, n46, n48, n49, n50, n54,
         n55, n56, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n70, n72,
         n73, n74, n76, n79, n80, n82, n83, n84, n88, n89, n90, n91, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n461, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1138, n1139, n1140, n1141, n1142, n1144, n1147, n1148, n1149, n1150,
         n1151, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1724, n1725, n1726, n1727, n1728, n1729, n1731, n1732, n1733, n1734,
         n1736, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979;
  wire   [7:0] weight_cnt;
  wire   [1:0] state;
  wire   [3:0] n_state;
  wire   [4:0] channel_cnt;
  wire   [1:0] data_sel_col;
  wire   [1:0] data_sel_row;
  wire   [9:0] delay3_sram_waddr_b;
  wire   [3:0] delay_sram_bytemask_b;
  wire   [3:0] delay2_sram_bytemask_b;
  wire   [3:0] delay_sram_bytemask_c;
  wire   [3:0] delay_sram_bytemask_d;
  wire   [3:0] n_row;
  wire   [7:0] n_weight_cnt;
  wire   [7:0] delay_set;
  wire   [1:0] n_addr_col_sel_cnt;
  wire   [1:0] addr_col_sel_cnt;
  wire   [1:0] addr_row_sel_cnt;
  wire   [9:0] delay1_sram_waddr_b;
  wire   [9:0] delay2_sram_waddr_b;
  wire   [3:0] n_sram_bytemask_b;
  wire   [3:0] row;
  wire   [3:0] col;
  wire   [3:0] row_delay;
  wire   [3:0] col_delay;
  wire   [9:0] delay1_sram_waddr_c;
  wire   [9:0] delay1_sram_waddr_d;
  wire   [9:0] delay2_sram_waddr_c;
  wire   [9:0] delay2_sram_waddr_d;
  wire   [9:0] delay3_sram_waddr_c;
  wire   [9:0] delay3_sram_waddr_d;
  wire   [9:0] delay4_sram_waddr_c;
  wire   [9:0] delay4_sram_waddr_d;
  wire   [3:0] n_sram_bytemask_c;
  wire   [3:0] n_sram_bytemask_d;
  wire   [4:0] addr_change;
  wire   [4:2] delay_addr_change;
  wire   [4:0] delay_channel;
  wire   [4:0] delay2_channel;
  wire   [1:0] write_col;
  wire   [2:0] write_row;
  wire   [9:0] n_sram_raddr_a0;
  wire   [9:0] n_sram_raddr_a1;
  wire   [9:0] n_sram_raddr_a2;
  wire   [9:0] n_sram_raddr_a3;
  wire   [9:0] n_sram_raddr_a4;
  wire   [9:0] n_sram_raddr_a5;
  wire   [9:0] n_sram_raddr_a6;
  wire   [9:0] n_sram_raddr_a7;
  wire   [9:0] n_sram_raddr_a8;
  wire   [9:0] n_sram_raddr_b0;
  wire   [9:0] n_sram_raddr_b1;
  wire   [9:0] n_sram_raddr_b2;
  wire   [9:0] n_sram_raddr_b3;
  wire   [9:0] n_sram_raddr_b4;
  wire   [9:0] n_sram_raddr_b5;
  wire   [9:0] n_sram_raddr_b6;
  wire   [9:0] n_sram_raddr_b7;
  wire   [9:0] n_sram_raddr_b8;

  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_0 clk_gate_col_reg ( .CLK(clk), 
        .EN(net19513), .ENCLK(net19718) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_26 clk_gate_weight_cnt_reg ( 
        .CLK(clk), .EN(net19513), .ENCLK(net19723) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_25 clk_gate_sram_raddr_weight_reg ( 
        .CLK(clk), .EN(net19836), .ENCLK(net19818) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_24 clk_gate_sram_raddr_weight_reg_0 ( 
        .CLK(clk), .EN(net19836), .ENCLK(net19916) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_23 clk_gate_delay1_sram_waddr_b_reg ( 
        .CLK(clk), .EN(net19921), .ENCLK(net19954) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_22 clk_gate_delay1_sram_waddr_c_reg ( 
        .CLK(clk), .EN(net19959), .ENCLK(net19973) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_21 clk_gate_delay1_sram_waddr_d_reg ( 
        .CLK(clk), .EN(net19959), .ENCLK(net19989) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_20 clk_gate_channel_cnt_reg ( 
        .CLK(clk), .EN(net19993), .ENCLK(net20001) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_19 clk_gate_addr_change_reg ( 
        .CLK(clk), .EN(net20004), .ENCLK(net20013) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_18 clk_gate_sram_raddr_a7_reg ( 
        .CLK(clk), .EN(net20953), .ENCLK(net20494) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_17 clk_gate_sram_raddr_a1_reg ( 
        .CLK(clk), .EN(net20953), .ENCLK(net20939) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_16 clk_gate_sram_raddr_a4_reg ( 
        .CLK(clk), .EN(net20953), .ENCLK(net21376) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_15 clk_gate_sram_raddr_a8_reg ( 
        .CLK(clk), .EN(net22280), .ENCLK(net21821) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_14 clk_gate_sram_raddr_a2_reg ( 
        .CLK(clk), .EN(net22280), .ENCLK(net22266) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_13 clk_gate_sram_raddr_a5_reg ( 
        .CLK(clk), .EN(net22280), .ENCLK(net22703) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_12 clk_gate_sram_raddr_a0_reg ( 
        .CLK(clk), .EN(net23610), .ENCLK(net23149) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_11 clk_gate_sram_raddr_a3_reg ( 
        .CLK(clk), .EN(net23610), .ENCLK(net23595) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_10 clk_gate_sram_raddr_a6_reg ( 
        .CLK(clk), .EN(net23610), .ENCLK(net24033) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_9 clk_gate_sram_raddr_b7_reg ( 
        .CLK(clk), .EN(net28264), .ENCLK(net24567) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_8 clk_gate_sram_raddr_b8_reg ( 
        .CLK(clk), .EN(net28264), .ENCLK(net25082) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_7 clk_gate_sram_raddr_b0_reg ( 
        .CLK(clk), .EN(net28264), .ENCLK(net25597) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_6 clk_gate_sram_raddr_b1_reg ( 
        .CLK(clk), .EN(net28264), .ENCLK(net26112) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_5 clk_gate_sram_raddr_b2_reg ( 
        .CLK(clk), .EN(net28264), .ENCLK(net26627) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_4 clk_gate_sram_raddr_b3_reg ( 
        .CLK(clk), .EN(net28264), .ENCLK(net27142) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_3 clk_gate_sram_raddr_b4_reg ( 
        .CLK(clk), .EN(net28264), .ENCLK(net27657) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_2 clk_gate_sram_raddr_b5_reg ( 
        .CLK(clk), .EN(net28264), .ENCLK(net28172) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_1 clk_gate_sram_raddr_b6_reg ( 
        .CLK(clk), .EN(net28264), .ENCLK(net28687) );
  DFFSSRX1_HVT channel_cnt_reg_0_ ( .D(1'b0), .SETB(n112), .RSTB(net19998), 
        .CLK(net20001), .Q(channel_cnt[0]) );
  DFFSSRX1_HVT state_reg_3_ ( .D(1'b0), .SETB(n111), .RSTB(n_state[3]), .CLK(
        clk), .Q(n232), .QN(n1108) );
  DFFSSRX1_HVT state_reg_0_ ( .D(1'b0), .SETB(n114), .RSTB(n_state[0]), .CLK(
        clk), .Q(state[0]), .QN(n166) );
  DFFSSRX1_HVT weight_cnt_reg_0_ ( .D(1'b0), .SETB(n113), .RSTB(
        n_weight_cnt[0]), .CLK(net19723), .Q(weight_cnt[0]), .QN(n227) );
  DFFSSRX1_HVT delay_set_reg_0_ ( .D(1'b0), .SETB(n113), .RSTB(weight_cnt[0]), 
        .CLK(clk), .Q(delay_set[0]) );
  DFFSSRX1_HVT set_reg_0_ ( .D(1'b0), .SETB(n112), .RSTB(delay_set[0]), .CLK(
        clk), .Q(set[0]) );
  DFFSSRX1_HVT delay_conv_done_reg ( .D(1'b0), .SETB(n135), .RSTB(n_conv_done), 
        .CLK(clk), .Q(delay_conv_done) );
  DFFSSRX1_HVT delay2_conv_done_reg ( .D(1'b0), .SETB(n147), .RSTB(
        delay_conv_done), .CLK(clk), .Q(delay2_conv_done) );
  DFFSSRX1_HVT delay3_conv_done_reg ( .D(1'b0), .SETB(n144), .RSTB(
        delay2_conv_done), .CLK(clk), .Q(delay3_conv_done) );
  DFFSSRX1_HVT conv_done_reg ( .D(1'b0), .SETB(n136), .RSTB(delay3_conv_done), 
        .CLK(clk), .Q(conv_done) );
  DFFSSRX1_HVT state_reg_2_ ( .D(1'b0), .SETB(n135), .RSTB(n_state[2]), .CLK(
        clk), .QN(n1109) );
  DFFSSRX1_HVT weight_cnt_reg_1_ ( .D(1'b0), .SETB(n114), .RSTB(
        n_weight_cnt[1]), .CLK(net19723), .Q(weight_cnt[1]), .QN(n354) );
  DFFSSRX1_HVT delay_set_reg_1_ ( .D(1'b0), .SETB(n147), .RSTB(weight_cnt[1]), 
        .CLK(clk), .Q(delay_set[1]) );
  DFFSSRX1_HVT set_reg_1_ ( .D(1'b0), .SETB(n144), .RSTB(delay_set[1]), .CLK(
        clk), .Q(set[1]) );
  DFFSSRX1_HVT delay1_conv1_done_reg ( .D(1'b0), .SETB(n139), .RSTB(
        n_conv1_done), .CLK(clk), .Q(delay1_conv1_done) );
  DFFSSRX1_HVT delay2_conv1_done_reg ( .D(1'b0), .SETB(n135), .RSTB(
        delay1_conv1_done), .CLK(clk), .Q(delay2_conv1_done) );
  DFFSSRX1_HVT delay3_conv1_done_reg ( .D(1'b0), .SETB(n146), .RSTB(
        delay2_conv1_done), .CLK(clk), .Q(delay3_conv1_done) );
  DFFSSRX1_HVT delay4_conv1_done_reg ( .D(1'b0), .SETB(n143), .RSTB(
        delay3_conv1_done), .CLK(clk), .Q(delay4_conv1_done) );
  DFFSSRX1_HVT conv1_done_reg ( .D(1'b0), .SETB(n139), .RSTB(delay4_conv1_done), .CLK(clk), .Q(conv1_done), .QN(n369) );
  DFFSSRX1_HVT state_reg_1_ ( .D(1'b0), .SETB(n101), .RSTB(n_state[1]), .CLK(
        clk), .Q(state[1]), .QN(n177) );
  DFFSSRX1_HVT weight_cnt_reg_7_ ( .D(1'b0), .SETB(n111), .RSTB(
        n_weight_cnt[7]), .CLK(net19723), .Q(weight_cnt[7]), .QN(n324) );
  DFFSSRX1_HVT delay_set_reg_7_ ( .D(1'b0), .SETB(n156), .RSTB(weight_cnt[7]), 
        .CLK(clk), .Q(delay_set[7]) );
  DFFSSRX1_HVT set_reg_7_ ( .D(1'b0), .SETB(n100), .RSTB(delay_set[7]), .CLK(
        clk), .Q(set[7]) );
  DFFSSRX1_HVT weight_cnt_reg_6_ ( .D(1'b0), .SETB(n138), .RSTB(
        n_weight_cnt[6]), .CLK(net19723), .Q(weight_cnt[6]), .QN(n213) );
  DFFSSRX1_HVT delay_set_reg_6_ ( .D(1'b0), .SETB(n142), .RSTB(weight_cnt[6]), 
        .CLK(clk), .Q(delay_set[6]) );
  DFFSSRX1_HVT set_reg_6_ ( .D(1'b0), .SETB(n134), .RSTB(delay_set[6]), .CLK(
        clk), .Q(set[6]) );
  DFFSSRX1_HVT weight_cnt_reg_5_ ( .D(1'b0), .SETB(n141), .RSTB(
        n_weight_cnt[5]), .CLK(net19723), .Q(weight_cnt[5]), .QN(n275) );
  DFFSSRX1_HVT delay_set_reg_5_ ( .D(1'b0), .SETB(n146), .RSTB(weight_cnt[5]), 
        .CLK(clk), .Q(delay_set[5]) );
  DFFSSRX1_HVT set_reg_5_ ( .D(1'b0), .SETB(n143), .RSTB(delay_set[5]), .CLK(
        clk), .Q(set[5]) );
  DFFSSRX1_HVT weight_cnt_reg_4_ ( .D(1'b0), .SETB(n145), .RSTB(
        n_weight_cnt[4]), .CLK(net19723), .Q(weight_cnt[4]) );
  DFFSSRX1_HVT delay_set_reg_4_ ( .D(1'b0), .SETB(n139), .RSTB(weight_cnt[4]), 
        .CLK(clk), .Q(delay_set[4]) );
  DFFSSRX1_HVT set_reg_4_ ( .D(1'b0), .SETB(n134), .RSTB(delay_set[4]), .CLK(
        clk), .Q(set[4]) );
  DFFSSRX1_HVT weight_cnt_reg_3_ ( .D(1'b0), .SETB(n132), .RSTB(
        n_weight_cnt[3]), .CLK(net19723), .Q(weight_cnt[3]), .QN(n176) );
  DFFSSRX1_HVT delay_set_reg_3_ ( .D(1'b0), .SETB(n146), .RSTB(weight_cnt[3]), 
        .CLK(clk), .Q(delay_set[3]) );
  DFFSSRX1_HVT set_reg_3_ ( .D(1'b0), .SETB(n143), .RSTB(delay_set[3]), .CLK(
        clk), .Q(set[3]) );
  DFFSSRX1_HVT weight_cnt_reg_2_ ( .D(1'b0), .SETB(n136), .RSTB(
        n_weight_cnt[2]), .CLK(net19723), .Q(weight_cnt[2]), .QN(n367) );
  DFFSSRX1_HVT delay_set_reg_2_ ( .D(1'b0), .SETB(n138), .RSTB(weight_cnt[2]), 
        .CLK(clk), .Q(delay_set[2]) );
  DFFSSRX1_HVT set_reg_2_ ( .D(1'b0), .SETB(n134), .RSTB(delay_set[2]), .CLK(
        clk), .Q(set[2]) );
  DFFSSRX1_HVT delay_load_conv2_bias0_enable_reg ( .D(1'b0), .SETB(n145), 
        .RSTB(n1738), .CLK(clk), .Q(delay_load_conv2_bias0_enable) );
  DFFSSRX1_HVT load_conv2_bias0_enable_reg ( .D(1'b0), .SETB(n141), .RSTB(
        delay_load_conv2_bias0_enable), .CLK(clk), .Q(load_conv2_bias0_enable)
         );
  DFFSSRX1_HVT col_reg_0_ ( .D(1'b0), .SETB(n141), .RSTB(net19714), .CLK(
        net19718), .Q(col[0]), .QN(n194) );
  DFFSSRX1_HVT col_delay_reg_0_ ( .D(1'b0), .SETB(n138), .RSTB(col[0]), .CLK(
        clk), .Q(col_delay[0]) );
  DFFSSRX1_HVT write_col_reg_0_ ( .D(1'b0), .SETB(n101), .RSTB(col_delay[0]), 
        .CLK(clk), .Q(write_col[0]), .QN(n352) );
  DFFSSRX1_HVT col_reg_1_ ( .D(1'b0), .SETB(n145), .RSTB(net19709), .CLK(
        net19718), .Q(col[1]), .QN(n268) );
  DFFSSRX1_HVT col_delay_reg_1_ ( .D(1'b0), .SETB(n101), .RSTB(col[1]), .CLK(
        clk), .Q(col_delay[1]) );
  DFFSSRX1_HVT write_col_reg_1_ ( .D(1'b0), .SETB(n100), .RSTB(col_delay[1]), 
        .CLK(clk), .Q(write_col[1]), .QN(n235) );
  DFFSSRX1_HVT col_reg_2_ ( .D(1'b0), .SETB(n132), .RSTB(net19704), .CLK(
        net19718), .Q(col[2]), .QN(n167) );
  DFFSSRX1_HVT col_delay_reg_2_ ( .D(1'b0), .SETB(n142), .RSTB(col[2]), .CLK(
        clk), .Q(col_delay[2]) );
  DFFSSRX1_HVT write_col_reg_2_ ( .D(1'b0), .SETB(n132), .RSTB(col_delay[2]), 
        .CLK(clk), .Q(n180), .QN(n1146) );
  DFFSSRX1_HVT col_reg_3_ ( .D(1'b0), .SETB(n137), .RSTB(net19699), .CLK(
        net19718), .Q(col[3]), .QN(n163) );
  DFFSSRX1_HVT col_delay_reg_3_ ( .D(1'b0), .SETB(n145), .RSTB(col[3]), .CLK(
        clk), .Q(col_delay[3]) );
  DFFSSRX1_HVT write_col_reg_3_ ( .D(1'b0), .SETB(n141), .RSTB(col_delay[3]), 
        .CLK(clk), .Q(n181), .QN(n1145) );
  DFFSSRX1_HVT addr_col_sel_cnt_reg_0_ ( .D(1'b0), .SETB(n138), .RSTB(
        n_addr_col_sel_cnt[0]), .CLK(clk), .Q(addr_col_sel_cnt[0]), .QN(n1136)
         );
  DFFSSRX1_HVT data_sel_col_reg_0_ ( .D(1'b0), .SETB(n132), .RSTB(
        addr_col_sel_cnt[0]), .CLK(clk), .Q(data_sel_col[0]) );
  DFFSSRX1_HVT addr_col_sel_cnt_reg_1_ ( .D(1'b0), .SETB(n145), .RSTB(
        n_addr_col_sel_cnt[1]), .CLK(clk), .Q(addr_col_sel_cnt[1]), .QN(n1135)
         );
  DFFSSRX1_HVT data_sel_col_reg_1_ ( .D(1'b0), .SETB(n141), .RSTB(
        addr_col_sel_cnt[1]), .CLK(clk), .Q(data_sel_col[1]) );
  DFFSSRX1_HVT addr_row_sel_cnt_reg_0_ ( .D(1'b0), .SETB(n136), .RSTB(
        n_addr_row_sel_cnt_0_), .CLK(clk), .Q(addr_row_sel_cnt[0]), .QN(n276)
         );
  DFFSSRX1_HVT data_sel_row_reg_0_ ( .D(1'b0), .SETB(n132), .RSTB(
        addr_row_sel_cnt[0]), .CLK(clk), .Q(data_sel_row[0]) );
  DFFSSRX1_HVT addr_row_sel_cnt_reg_1_ ( .D(n487), .SETB(n1735), .RSTB(n105), 
        .CLK(clk), .Q(addr_row_sel_cnt[1]), .QN(n1137) );
  DFFSSRX1_HVT data_sel_row_reg_1_ ( .D(1'b0), .SETB(n147), .RSTB(
        addr_row_sel_cnt[1]), .CLK(clk), .Q(data_sel_row[1]) );
  DFFSSRX1_HVT conv2_weight_done_reg ( .D(1'b0), .SETB(n142), .RSTB(net19715), 
        .CLK(net19718), .Q(conv2_weight_done) );
  DFFSSRX1_HVT row_reg_0_ ( .D(1'b0), .SETB(n142), .RSTB(n_row[0]), .CLK(
        net19718), .Q(row[0]), .QN(n183) );
  DFFSSRX1_HVT row_delay_reg_0_ ( .D(1'b0), .SETB(n144), .RSTB(row[0]), .CLK(
        clk), .Q(row_delay[0]) );
  DFFSSRX1_HVT write_row_reg_0_ ( .D(1'b0), .SETB(n136), .RSTB(row_delay[0]), 
        .CLK(clk), .Q(write_row[0]) );
  DFFSSRX1_HVT delay_sram_bytemask_d_reg_1_ ( .D(1'b0), .SETB(n111), .RSTB(
        n_sram_bytemask_d[1]), .CLK(clk), .Q(delay_sram_bytemask_d[1]) );
  DFFSSRX1_HVT sram_bytemask_d_reg_1_ ( .D(1'b0), .SETB(n114), .RSTB(
        delay_sram_bytemask_d[1]), .CLK(clk), .Q(sram_bytemask_d[1]) );
  DFFSSRX1_HVT delay_sram_bytemask_c_reg_1_ ( .D(1'b0), .SETB(n113), .RSTB(
        n_sram_bytemask_c[1]), .CLK(clk), .Q(delay_sram_bytemask_c[1]) );
  DFFSSRX1_HVT sram_bytemask_c_reg_1_ ( .D(1'b0), .SETB(n112), .RSTB(
        delay_sram_bytemask_c[1]), .CLK(clk), .Q(sram_bytemask_c[1]) );
  DFFSSRX1_HVT delay_sram_bytemask_d_reg_0_ ( .D(1'b0), .SETB(n135), .RSTB(
        n_sram_bytemask_d[0]), .CLK(clk), .Q(delay_sram_bytemask_d[0]) );
  DFFSSRX1_HVT sram_bytemask_d_reg_0_ ( .D(1'b0), .SETB(n147), .RSTB(
        delay_sram_bytemask_d[0]), .CLK(clk), .Q(sram_bytemask_d[0]) );
  DFFSSRX1_HVT delay_sram_bytemask_c_reg_0_ ( .D(1'b0), .SETB(n144), .RSTB(
        n_sram_bytemask_c[0]), .CLK(clk), .Q(delay_sram_bytemask_c[0]) );
  DFFSSRX1_HVT sram_bytemask_c_reg_0_ ( .D(1'b0), .SETB(n136), .RSTB(
        delay_sram_bytemask_c[0]), .CLK(clk), .Q(sram_bytemask_c[0]) );
  DFFSSRX1_HVT delay_sram_bytemask_c_reg_2_ ( .D(1'b0), .SETB(n135), .RSTB(
        n_sram_bytemask_c[2]), .CLK(clk), .Q(delay_sram_bytemask_c[2]) );
  DFFSSRX1_HVT sram_bytemask_c_reg_2_ ( .D(1'b0), .SETB(n147), .RSTB(
        delay_sram_bytemask_c[2]), .CLK(clk), .Q(sram_bytemask_c[2]) );
  DFFSSRX1_HVT delay_sram_bytemask_c_reg_3_ ( .D(1'b0), .SETB(n144), .RSTB(
        n_sram_bytemask_c[3]), .CLK(clk), .Q(delay_sram_bytemask_c[3]) );
  DFFSSRX1_HVT sram_bytemask_c_reg_3_ ( .D(1'b0), .SETB(n139), .RSTB(
        delay_sram_bytemask_c[3]), .CLK(clk), .Q(sram_bytemask_c[3]) );
  DFFSSRX1_HVT delay_sram_bytemask_d_reg_2_ ( .D(1'b0), .SETB(n135), .RSTB(
        n_sram_bytemask_d[2]), .CLK(clk), .Q(delay_sram_bytemask_d[2]) );
  DFFSSRX1_HVT sram_bytemask_d_reg_2_ ( .D(1'b0), .SETB(n146), .RSTB(
        delay_sram_bytemask_d[2]), .CLK(clk), .Q(sram_bytemask_d[2]) );
  DFFSSRX1_HVT delay_sram_bytemask_d_reg_3_ ( .D(1'b0), .SETB(n143), .RSTB(
        n_sram_bytemask_d[3]), .CLK(clk), .Q(delay_sram_bytemask_d[3]) );
  DFFSSRX1_HVT sram_bytemask_d_reg_3_ ( .D(1'b0), .SETB(n139), .RSTB(
        delay_sram_bytemask_d[3]), .CLK(clk), .Q(sram_bytemask_d[3]) );
  DFFSSRX1_HVT row_reg_1_ ( .D(1'b0), .SETB(n133), .RSTB(n_row[1]), .CLK(
        net19718), .Q(row[1]), .QN(n237) );
  DFFSSRX1_HVT row_delay_reg_1_ ( .D(1'b0), .SETB(n101), .RSTB(row[1]), .CLK(
        clk), .Q(row_delay[1]) );
  DFFSSRX1_HVT write_row_reg_1_ ( .D(1'b0), .SETB(n156), .RSTB(row_delay[1]), 
        .CLK(clk), .QN(n1143) );
  DFFSSRX1_HVT box_sel_reg_2_ ( .D(n462), .SETB(n1723), .RSTB(n107), .CLK(clk), 
        .Q(box_sel[2]) );
  DFFSSRX1_HVT box_sel_reg_1_ ( .D(1'b0), .SETB(n100), .RSTB(n_box_sel_1_), 
        .CLK(clk), .Q(box_sel[1]) );
  DFFSSRX1_HVT box_sel_reg_0_ ( .D(n460), .SETB(n1730), .RSTB(n106), .CLK(clk), 
        .Q(box_sel[0]) );
  DFFSSRX1_HVT box_sel_reg_3_ ( .D(n459), .SETB(n1723), .RSTB(n105), .CLK(clk), 
        .Q(box_sel[3]) );
  DFFSSRX1_HVT row_reg_2_ ( .D(1'b0), .SETB(n114), .RSTB(n_row[2]), .CLK(
        net19718), .Q(row[2]), .QN(n179) );
  DFFSSRX1_HVT row_delay_reg_2_ ( .D(1'b0), .SETB(n137), .RSTB(row[2]), .CLK(
        clk), .Q(row_delay[2]) );
  DFFSSRX1_HVT write_row_reg_2_ ( .D(1'b0), .SETB(n134), .RSTB(row_delay[2]), 
        .CLK(clk), .Q(write_row[2]), .QN(n382) );
  DFFSSRX1_HVT row_reg_3_ ( .D(1'b0), .SETB(n100), .RSTB(n_row[3]), .CLK(
        net19718), .Q(row[3]), .QN(n234) );
  DFFSSRX1_HVT row_delay_reg_3_ ( .D(1'b0), .SETB(n146), .RSTB(row[3]), .CLK(
        clk), .Q(row_delay[3]) );
  DFFSSRX1_HVT write_row_reg_3_ ( .D(1'b0), .SETB(n143), .RSTB(row_delay[3]), 
        .CLK(clk), .QN(n302) );
  DFFSSRX1_HVT channel_cnt_reg_4_ ( .D(1'b0), .SETB(n156), .RSTB(net19994), 
        .CLK(net20001), .Q(channel_cnt[4]), .QN(n233) );
  DFFSSRX1_HVT channel_cnt_reg_3_ ( .D(1'b0), .SETB(n101), .RSTB(net19995), 
        .CLK(net20001), .Q(channel_cnt[3]) );
  DFFSSRX1_HVT channel_cnt_reg_2_ ( .D(1'b0), .SETB(n139), .RSTB(net19996), 
        .CLK(net20001), .Q(channel_cnt[2]), .QN(n363) );
  DFFSSRX1_HVT channel_cnt_reg_1_ ( .D(1'b0), .SETB(n144), .RSTB(net19997), 
        .CLK(net20001), .Q(channel_cnt[1]) );
  DFFSSRX1_HVT delay_load_conv1_bias_enable_reg ( .D(1'b0), .SETB(n139), 
        .RSTB(n1739), .CLK(clk), .Q(delay_load_conv1_bias_enable) );
  DFFSSRX1_HVT load_conv1_bias_enable_reg ( .D(1'b0), .SETB(n134), .RSTB(
        delay_load_conv1_bias_enable), .CLK(clk), .Q(load_conv1_bias_enable)
         );
  DFFSSRX1_HVT sram_raddr_weight_reg_7_ ( .D(1'b0), .SETB(n147), .RSTB(
        net19843), .CLK(net19916), .Q(sram_raddr_weight[7]), .QN(n318) );
  DFFSSRX1_HVT conv1_bias_set_reg_7_ ( .D(1'b0), .SETB(n146), .RSTB(
        sram_raddr_weight[7]), .CLK(clk), .Q(conv1_bias_set[7]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_6_ ( .D(1'b0), .SETB(n134), .RSTB(
        net19850), .CLK(net19916), .Q(sram_raddr_weight[6]), .QN(n315) );
  DFFSSRX1_HVT conv1_bias_set_reg_6_ ( .D(1'b0), .SETB(n143), .RSTB(
        sram_raddr_weight[6]), .CLK(clk), .Q(conv1_bias_set[6]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_5_ ( .D(1'b0), .SETB(n138), .RSTB(
        net19857), .CLK(net19916), .Q(sram_raddr_weight[5]), .QN(n372) );
  DFFSSRX1_HVT conv1_bias_set_reg_5_ ( .D(1'b0), .SETB(n138), .RSTB(
        sram_raddr_weight[5]), .CLK(clk), .Q(conv1_bias_set[5]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_3_ ( .D(1'b0), .SETB(n143), .RSTB(
        net19878), .CLK(net19916), .Q(sram_raddr_weight[3]), .QN(n321) );
  DFFSSRX1_HVT conv1_bias_set_reg_3_ ( .D(1'b0), .SETB(n134), .RSTB(
        sram_raddr_weight[3]), .CLK(clk), .Q(conv1_bias_set[3]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_16_ ( .D(1'b0), .SETB(n146), .RSTB(
        net19752), .CLK(net19818), .Q(sram_raddr_weight[16]), .QN(n381) );
  DFFSSRX1_HVT conv1_bias_set_reg_16_ ( .D(1'b0), .SETB(n145), .RSTB(
        sram_raddr_weight[16]), .CLK(clk), .Q(conv1_bias_set[16]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_15_ ( .D(1'b0), .SETB(n134), .RSTB(
        net19759), .CLK(net19818), .Q(sram_raddr_weight[15]), .QN(n355) );
  DFFSSRX1_HVT conv1_bias_set_reg_15_ ( .D(1'b0), .SETB(n141), .RSTB(
        sram_raddr_weight[15]), .CLK(clk), .Q(conv1_bias_set[15]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_14_ ( .D(1'b0), .SETB(n137), .RSTB(
        net19766), .CLK(net19818), .Q(sram_raddr_weight[14]) );
  DFFSSRX1_HVT conv1_bias_set_reg_14_ ( .D(1'b0), .SETB(n138), .RSTB(
        sram_raddr_weight[14]), .CLK(clk), .Q(conv1_bias_set[14]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_13_ ( .D(1'b0), .SETB(n142), .RSTB(
        net19773), .CLK(net19818), .Q(sram_raddr_weight[13]), .QN(n320) );
  DFFSSRX1_HVT conv1_bias_set_reg_13_ ( .D(1'b0), .SETB(n101), .RSTB(
        sram_raddr_weight[13]), .CLK(clk), .Q(conv1_bias_set[13]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_12_ ( .D(1'b0), .SETB(n133), .RSTB(
        net19780), .CLK(net19818), .Q(sram_raddr_weight[12]), .QN(n319) );
  DFFSSRX1_HVT conv1_bias_set_reg_12_ ( .D(1'b0), .SETB(n100), .RSTB(
        sram_raddr_weight[12]), .CLK(clk), .Q(conv1_bias_set[12]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_11_ ( .D(1'b0), .SETB(n133), .RSTB(
        net19787), .CLK(net19818), .Q(sram_raddr_weight[11]) );
  DFFSSRX1_HVT conv1_bias_set_reg_11_ ( .D(1'b0), .SETB(n100), .RSTB(
        sram_raddr_weight[11]), .CLK(clk), .Q(conv1_bias_set[11]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_10_ ( .D(1'b0), .SETB(n114), .RSTB(
        net19794), .CLK(net19818), .Q(sram_raddr_weight[10]), .QN(n356) );
  DFFSSRX1_HVT conv1_bias_set_reg_10_ ( .D(1'b0), .SETB(n100), .RSTB(
        sram_raddr_weight[10]), .CLK(clk), .Q(conv1_bias_set[10]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_9_ ( .D(1'b0), .SETB(n100), .RSTB(
        net19808), .CLK(net19818), .Q(sram_raddr_weight[9]), .QN(n296) );
  DFFSSRX1_HVT conv1_bias_set_reg_9_ ( .D(1'b0), .SETB(n132), .RSTB(
        sram_raddr_weight[9]), .CLK(clk), .Q(conv1_bias_set[9]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_8_ ( .D(1'b0), .SETB(n142), .RSTB(
        net19815), .CLK(net19818), .Q(sram_raddr_weight[8]) );
  DFFSSRX1_HVT conv1_bias_set_reg_8_ ( .D(1'b0), .SETB(n145), .RSTB(
        sram_raddr_weight[8]), .CLK(clk), .Q(conv1_bias_set[8]) );
  DFFSSRX1_HVT conv1_weight_done_reg ( .D(1'b0), .SETB(n141), .RSTB(
        n_conv1_weight_done), .CLK(clk), .Q(conv1_weight_done), .QN(n178) );
  DFFSSRX1_HVT load_data_enable_reg ( .D(1'b0), .SETB(n138), .RSTB(
        n_load_data_enable), .CLK(clk), .Q(load_data_enable) );
  DFFSSRX1_HVT write_enable_reg ( .D(1'b0), .SETB(n132), .RSTB(n_write_enable), 
        .CLK(clk), .Q(write_enable) );
  DFFSSRX1_HVT delay_write_enable_reg ( .D(1'b0), .SETB(n145), .RSTB(
        write_enable), .CLK(clk), .Q(delay_write_enable) );
  DFFSSRX1_HVT delay2_write_enable_reg ( .D(1'b0), .SETB(n141), .RSTB(
        delay_write_enable), .CLK(clk), .Q(delay2_write_enable) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_9_ ( .D(1'b0), .SETB(N2888), .RSTB(
        net19924), .CLK(net19954), .Q(delay1_sram_waddr_b[9]) );
  DFFSSRX1_HVT delay2_sram_waddr_b_reg_9_ ( .D(1'b0), .SETB(n136), .RSTB(
        delay1_sram_waddr_b[9]), .CLK(clk), .Q(delay2_sram_waddr_b[9]) );
  DFFSSRX1_HVT delay3_sram_waddr_b_reg_9_ ( .D(1'b0), .SETB(n132), .RSTB(
        delay2_sram_waddr_b[9]), .CLK(clk), .Q(delay3_sram_waddr_b[9]) );
  DFFSSRX1_HVT sram_waddr_b_reg_9_ ( .D(1'b0), .SETB(n147), .RSTB(
        delay3_sram_waddr_b[9]), .CLK(clk), .Q(sram_waddr_b[9]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_8_ ( .D(1'b0), .SETB(N2888), .RSTB(
        net19927), .CLK(net19954), .Q(delay1_sram_waddr_b[8]), .QN(n328) );
  DFFSSRX1_HVT delay2_sram_waddr_b_reg_8_ ( .D(1'b0), .SETB(n144), .RSTB(
        delay1_sram_waddr_b[8]), .CLK(clk), .Q(delay2_sram_waddr_b[8]) );
  DFFSSRX1_HVT delay3_sram_waddr_b_reg_8_ ( .D(1'b0), .SETB(n136), .RSTB(
        delay2_sram_waddr_b[8]), .CLK(clk), .Q(delay3_sram_waddr_b[8]) );
  DFFSSRX1_HVT sram_waddr_b_reg_8_ ( .D(1'b0), .SETB(n111), .RSTB(
        delay3_sram_waddr_b[8]), .CLK(clk), .Q(sram_waddr_b[8]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_7_ ( .D(1'b0), .SETB(N2888), .RSTB(
        net19930), .CLK(net19954), .Q(delay1_sram_waddr_b[7]) );
  DFFSSRX1_HVT delay2_sram_waddr_b_reg_7_ ( .D(1'b0), .SETB(n114), .RSTB(
        delay1_sram_waddr_b[7]), .CLK(clk), .Q(delay2_sram_waddr_b[7]) );
  DFFSSRX1_HVT delay3_sram_waddr_b_reg_7_ ( .D(1'b0), .SETB(n113), .RSTB(
        delay2_sram_waddr_b[7]), .CLK(clk), .Q(delay3_sram_waddr_b[7]) );
  DFFSSRX1_HVT sram_waddr_b_reg_7_ ( .D(1'b0), .SETB(n112), .RSTB(
        delay3_sram_waddr_b[7]), .CLK(clk), .Q(sram_waddr_b[7]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_6_ ( .D(1'b0), .SETB(N2888), .RSTB(
        net19933), .CLK(net19954), .Q(delay1_sram_waddr_b[6]) );
  DFFSSRX1_HVT delay2_sram_waddr_b_reg_6_ ( .D(1'b0), .SETB(n135), .RSTB(
        delay1_sram_waddr_b[6]), .CLK(clk), .Q(delay2_sram_waddr_b[6]) );
  DFFSSRX1_HVT delay3_sram_waddr_b_reg_6_ ( .D(1'b0), .SETB(n147), .RSTB(
        delay2_sram_waddr_b[6]), .CLK(clk), .Q(delay3_sram_waddr_b[6]) );
  DFFSSRX1_HVT sram_waddr_b_reg_6_ ( .D(1'b0), .SETB(n144), .RSTB(
        delay3_sram_waddr_b[6]), .CLK(clk), .Q(sram_waddr_b[6]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_5_ ( .D(1'b0), .SETB(N2888), .RSTB(
        net19936), .CLK(net19954), .Q(delay1_sram_waddr_b[5]), .QN(n365) );
  DFFSSRX1_HVT delay2_sram_waddr_b_reg_5_ ( .D(1'b0), .SETB(n136), .RSTB(
        delay1_sram_waddr_b[5]), .CLK(clk), .Q(delay2_sram_waddr_b[5]) );
  DFFSSRX1_HVT delay3_sram_waddr_b_reg_5_ ( .D(1'b0), .SETB(n135), .RSTB(
        delay2_sram_waddr_b[5]), .CLK(clk), .Q(delay3_sram_waddr_b[5]) );
  DFFSSRX1_HVT sram_waddr_b_reg_5_ ( .D(1'b0), .SETB(n147), .RSTB(
        delay3_sram_waddr_b[5]), .CLK(clk), .Q(sram_waddr_b[5]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_4_ ( .D(1'b0), .SETB(N2888), .RSTB(
        net19939), .CLK(net19954), .Q(delay1_sram_waddr_b[4]) );
  DFFSSRX1_HVT delay2_sram_waddr_b_reg_4_ ( .D(1'b0), .SETB(n144), .RSTB(
        delay1_sram_waddr_b[4]), .CLK(clk), .Q(delay2_sram_waddr_b[4]) );
  DFFSSRX1_HVT delay3_sram_waddr_b_reg_4_ ( .D(1'b0), .SETB(n139), .RSTB(
        delay2_sram_waddr_b[4]), .CLK(clk), .Q(delay3_sram_waddr_b[4]) );
  DFFSSRX1_HVT sram_waddr_b_reg_4_ ( .D(1'b0), .SETB(n135), .RSTB(
        delay3_sram_waddr_b[4]), .CLK(clk), .Q(sram_waddr_b[4]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_3_ ( .D(1'b0), .SETB(N2888), .RSTB(
        net19942), .CLK(net19954), .Q(delay1_sram_waddr_b[3]), .QN(n366) );
  DFFSSRX1_HVT delay2_sram_waddr_b_reg_3_ ( .D(1'b0), .SETB(n146), .RSTB(
        delay1_sram_waddr_b[3]), .CLK(clk), .Q(delay2_sram_waddr_b[3]) );
  DFFSSRX1_HVT delay3_sram_waddr_b_reg_3_ ( .D(1'b0), .SETB(n143), .RSTB(
        delay2_sram_waddr_b[3]), .CLK(clk), .Q(delay3_sram_waddr_b[3]) );
  DFFSSRX1_HVT sram_waddr_b_reg_3_ ( .D(1'b0), .SETB(n139), .RSTB(
        delay3_sram_waddr_b[3]), .CLK(clk), .Q(sram_waddr_b[3]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_2_ ( .D(1'b0), .SETB(N2888), .RSTB(
        net19945), .CLK(net19954), .Q(delay1_sram_waddr_b[2]) );
  DFFSSRX1_HVT delay2_sram_waddr_b_reg_2_ ( .D(1'b0), .SETB(n101), .RSTB(
        delay1_sram_waddr_b[2]), .CLK(clk), .Q(delay2_sram_waddr_b[2]) );
  DFFSSRX1_HVT delay3_sram_waddr_b_reg_2_ ( .D(1'b0), .SETB(n156), .RSTB(
        delay2_sram_waddr_b[2]), .CLK(clk), .Q(delay3_sram_waddr_b[2]) );
  DFFSSRX1_HVT sram_waddr_b_reg_2_ ( .D(1'b0), .SETB(n100), .RSTB(
        delay3_sram_waddr_b[2]), .CLK(clk), .Q(sram_waddr_b[2]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_1_ ( .D(1'b0), .SETB(N2888), .RSTB(
        net19948), .CLK(net19954), .Q(delay1_sram_waddr_b[1]) );
  DFFSSRX1_HVT delay2_sram_waddr_b_reg_1_ ( .D(1'b0), .SETB(n113), .RSTB(
        delay1_sram_waddr_b[1]), .CLK(clk), .Q(delay2_sram_waddr_b[1]) );
  DFFSSRX1_HVT delay3_sram_waddr_b_reg_1_ ( .D(1'b0), .SETB(n134), .RSTB(
        delay2_sram_waddr_b[1]), .CLK(clk), .Q(delay3_sram_waddr_b[1]) );
  DFFSSRX1_HVT sram_waddr_b_reg_1_ ( .D(1'b0), .SETB(n146), .RSTB(
        delay3_sram_waddr_b[1]), .CLK(clk), .Q(sram_waddr_b[1]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_0_ ( .D(1'b0), .SETB(N2888), .RSTB(
        net19951), .CLK(net19954), .Q(delay1_sram_waddr_b[0]) );
  DFFSSRX1_HVT delay2_sram_waddr_b_reg_0_ ( .D(1'b0), .SETB(n143), .RSTB(
        delay1_sram_waddr_b[0]), .CLK(clk), .Q(delay2_sram_waddr_b[0]) );
  DFFSSRX1_HVT delay3_sram_waddr_b_reg_0_ ( .D(1'b0), .SETB(n139), .RSTB(
        delay2_sram_waddr_b[0]), .CLK(clk), .Q(delay3_sram_waddr_b[0]) );
  DFFSSRX1_HVT sram_waddr_b_reg_0_ ( .D(1'b0), .SETB(n134), .RSTB(
        delay3_sram_waddr_b[0]), .CLK(clk), .Q(sram_waddr_b[0]) );
  DFFSSRX1_HVT delay_sram_bytemask_b_reg_3_ ( .D(1'b0), .SETB(n146), .RSTB(
        n_sram_bytemask_b[3]), .CLK(clk), .Q(delay_sram_bytemask_b[3]) );
  DFFSSRX1_HVT delay2_sram_bytemask_b_reg_3_ ( .D(1'b0), .SETB(n143), .RSTB(
        delay_sram_bytemask_b[3]), .CLK(clk), .Q(delay2_sram_bytemask_b[3]) );
  DFFSSRX1_HVT sram_bytemask_b_reg_3_ ( .D(1'b0), .SETB(n138), .RSTB(
        delay2_sram_bytemask_b[3]), .CLK(clk), .Q(sram_bytemask_b[3]) );
  DFFSSRX1_HVT delay_sram_bytemask_b_reg_2_ ( .D(1'b0), .SETB(n134), .RSTB(
        n_sram_bytemask_b[2]), .CLK(clk), .Q(delay_sram_bytemask_b[2]) );
  DFFSSRX1_HVT delay2_sram_bytemask_b_reg_2_ ( .D(1'b0), .SETB(n145), .RSTB(
        delay_sram_bytemask_b[2]), .CLK(clk), .Q(delay2_sram_bytemask_b[2]) );
  DFFSSRX1_HVT sram_bytemask_b_reg_2_ ( .D(1'b0), .SETB(n141), .RSTB(
        delay2_sram_bytemask_b[2]), .CLK(clk), .Q(sram_bytemask_b[2]) );
  DFFSSRX1_HVT delay_sram_bytemask_b_reg_1_ ( .D(1'b0), .SETB(n138), .RSTB(
        n_sram_bytemask_b[1]), .CLK(clk), .Q(delay_sram_bytemask_b[1]) );
  DFFSSRX1_HVT delay2_sram_bytemask_b_reg_1_ ( .D(1'b0), .SETB(n101), .RSTB(
        delay_sram_bytemask_b[1]), .CLK(clk), .Q(delay2_sram_bytemask_b[1]) );
  DFFSSRX1_HVT sram_bytemask_b_reg_1_ ( .D(1'b0), .SETB(n113), .RSTB(
        delay2_sram_bytemask_b[1]), .CLK(clk), .Q(sram_bytemask_b[1]) );
  DFFSSRX1_HVT delay_sram_bytemask_b_reg_0_ ( .D(1'b0), .SETB(n100), .RSTB(
        n_sram_bytemask_b[0]), .CLK(clk), .Q(delay_sram_bytemask_b[0]) );
  DFFSSRX1_HVT delay2_sram_bytemask_b_reg_0_ ( .D(1'b0), .SETB(n114), .RSTB(
        delay_sram_bytemask_b[0]), .CLK(clk), .Q(delay2_sram_bytemask_b[0]) );
  DFFSSRX1_HVT sram_bytemask_b_reg_0_ ( .D(1'b0), .SETB(n132), .RSTB(
        delay2_sram_bytemask_b[0]), .CLK(clk), .Q(sram_bytemask_b[0]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_1_ ( .D(1'b0), .SETB(n101), .RSTB(
        net19899), .CLK(net19916), .Q(sram_raddr_weight[1]), .QN(n364) );
  DFFSSRX1_HVT conv1_bias_set_reg_1_ ( .D(1'b0), .SETB(n145), .RSTB(
        sram_raddr_weight[1]), .CLK(clk), .Q(conv1_bias_set[1]) );
  DFFSSRX1_HVT delay_load_conv2_bias1_enable_reg ( .D(1'b0), .SETB(n141), 
        .RSTB(n1737), .CLK(clk), .Q(delay_load_conv2_bias1_enable) );
  DFFSSRX1_HVT load_conv2_bias1_enable_reg ( .D(1'b0), .SETB(n138), .RSTB(
        delay_load_conv2_bias1_enable), .CLK(clk), .Q(load_conv2_bias1_enable)
         );
  DFFSSRX1_HVT sram_raddr_weight_reg_0_ ( .D(1'b0), .SETB(n136), .RSTB(
        net19913), .CLK(net19916), .Q(sram_raddr_weight[0]), .QN(n231) );
  DFFSSRX1_HVT conv1_bias_set_reg_0_ ( .D(1'b0), .SETB(n132), .RSTB(
        sram_raddr_weight[0]), .CLK(clk), .Q(conv1_bias_set[0]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_2_ ( .D(1'b0), .SETB(n143), .RSTB(
        net19885), .CLK(net19916), .Q(sram_raddr_weight[2]), .QN(n209) );
  DFFSSRX1_HVT conv1_bias_set_reg_2_ ( .D(1'b0), .SETB(n145), .RSTB(
        sram_raddr_weight[2]), .CLK(clk), .Q(conv1_bias_set[2]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_4_ ( .D(1'b0), .SETB(n146), .RSTB(
        net19871), .CLK(net19916), .Q(sram_raddr_weight[4]), .QN(n374) );
  DFFSSRX1_HVT conv1_bias_set_reg_4_ ( .D(1'b0), .SETB(n141), .RSTB(
        sram_raddr_weight[4]), .CLK(clk), .Q(conv1_bias_set[4]) );
  DFFSSRX1_HVT addr_change_reg_0_ ( .D(1'b0), .SETB(n135), .RSTB(net20010), 
        .CLK(net20013), .Q(addr_change[0]) );
  DFFSSRX1_HVT addr_change_reg_1_ ( .D(1'b0), .SETB(n139), .RSTB(net20009), 
        .CLK(net20013), .Q(addr_change[1]) );
  DFFSSRX1_HVT addr_change_reg_2_ ( .D(1'b0), .SETB(n144), .RSTB(net20008), 
        .CLK(net20013), .Q(addr_change[2]), .QN(n182) );
  DFFSSRX1_HVT addr_change_reg_3_ ( .D(1'b0), .SETB(n147), .RSTB(net20007), 
        .CLK(net20013), .Q(addr_change[3]), .QN(n236) );
  DFFSSRX1_HVT addr_change_reg_4_ ( .D(1'b0), .SETB(n135), .RSTB(net20006), 
        .CLK(net20013), .Q(addr_change[4]), .QN(n380) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_9_ ( .D(1'b0), .SETB(n139), .RSTB(
        net19977), .CLK(net19989), .Q(delay1_sram_waddr_d[9]), .QN(n385) );
  DFFSSRX1_HVT delay2_sram_waddr_d_reg_9_ ( .D(1'b0), .SETB(n136), .RSTB(
        delay1_sram_waddr_d[9]), .CLK(clk), .Q(delay2_sram_waddr_d[9]) );
  DFFSSRX1_HVT delay3_sram_waddr_d_reg_9_ ( .D(1'b0), .SETB(n132), .RSTB(
        delay2_sram_waddr_d[9]), .CLK(clk), .Q(delay3_sram_waddr_d[9]) );
  DFFSSRX1_HVT delay4_sram_waddr_d_reg_9_ ( .D(1'b0), .SETB(n147), .RSTB(
        delay3_sram_waddr_d[9]), .CLK(clk), .Q(delay4_sram_waddr_d[9]) );
  DFFSSRX1_HVT sram_waddr_d_reg_9_ ( .D(1'b0), .SETB(n144), .RSTB(
        delay4_sram_waddr_d[9]), .CLK(clk), .Q(sram_waddr_d[9]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_8_ ( .D(1'b0), .SETB(n142), .RSTB(
        net19978), .CLK(net19989), .Q(delay1_sram_waddr_d[8]) );
  DFFSSRX1_HVT delay2_sram_waddr_d_reg_8_ ( .D(1'b0), .SETB(n136), .RSTB(
        delay1_sram_waddr_d[8]), .CLK(clk), .Q(delay2_sram_waddr_d[8]) );
  DFFSSRX1_HVT delay3_sram_waddr_d_reg_8_ ( .D(1'b0), .SETB(n111), .RSTB(
        delay2_sram_waddr_d[8]), .CLK(clk), .Q(delay3_sram_waddr_d[8]) );
  DFFSSRX1_HVT delay4_sram_waddr_d_reg_8_ ( .D(1'b0), .SETB(n114), .RSTB(
        delay3_sram_waddr_d[8]), .CLK(clk), .Q(delay4_sram_waddr_d[8]) );
  DFFSSRX1_HVT sram_waddr_d_reg_8_ ( .D(1'b0), .SETB(n113), .RSTB(
        delay4_sram_waddr_d[8]), .CLK(clk), .Q(sram_waddr_d[8]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_7_ ( .D(1'b0), .SETB(n100), .RSTB(
        net19979), .CLK(net19989), .Q(delay1_sram_waddr_d[7]) );
  DFFSSRX1_HVT delay2_sram_waddr_d_reg_7_ ( .D(1'b0), .SETB(n112), .RSTB(
        delay1_sram_waddr_d[7]), .CLK(clk), .Q(delay2_sram_waddr_d[7]) );
  DFFSSRX1_HVT delay3_sram_waddr_d_reg_7_ ( .D(1'b0), .SETB(n135), .RSTB(
        delay2_sram_waddr_d[7]), .CLK(clk), .Q(delay3_sram_waddr_d[7]) );
  DFFSSRX1_HVT delay4_sram_waddr_d_reg_7_ ( .D(1'b0), .SETB(n147), .RSTB(
        delay3_sram_waddr_d[7]), .CLK(clk), .Q(delay4_sram_waddr_d[7]) );
  DFFSSRX1_HVT sram_waddr_d_reg_7_ ( .D(1'b0), .SETB(n144), .RSTB(
        delay4_sram_waddr_d[7]), .CLK(clk), .Q(sram_waddr_d[7]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_6_ ( .D(1'b0), .SETB(n133), .RSTB(
        net19980), .CLK(net19989), .Q(delay1_sram_waddr_d[6]) );
  DFFSSRX1_HVT delay2_sram_waddr_d_reg_6_ ( .D(1'b0), .SETB(n136), .RSTB(
        delay1_sram_waddr_d[6]), .CLK(clk), .Q(delay2_sram_waddr_d[6]) );
  DFFSSRX1_HVT delay3_sram_waddr_d_reg_6_ ( .D(1'b0), .SETB(n135), .RSTB(
        delay2_sram_waddr_d[6]), .CLK(clk), .Q(delay3_sram_waddr_d[6]) );
  DFFSSRX1_HVT delay4_sram_waddr_d_reg_6_ ( .D(1'b0), .SETB(n147), .RSTB(
        delay3_sram_waddr_d[6]), .CLK(clk), .Q(delay4_sram_waddr_d[6]) );
  DFFSSRX1_HVT sram_waddr_d_reg_6_ ( .D(1'b0), .SETB(n144), .RSTB(
        delay4_sram_waddr_d[6]), .CLK(clk), .Q(sram_waddr_d[6]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_5_ ( .D(1'b0), .SETB(n112), .RSTB(
        net19981), .CLK(net19989), .Q(delay1_sram_waddr_d[5]) );
  DFFSSRX1_HVT delay2_sram_waddr_d_reg_5_ ( .D(1'b0), .SETB(n139), .RSTB(
        delay1_sram_waddr_d[5]), .CLK(clk), .Q(delay2_sram_waddr_d[5]) );
  DFFSSRX1_HVT delay3_sram_waddr_d_reg_5_ ( .D(1'b0), .SETB(n135), .RSTB(
        delay2_sram_waddr_d[5]), .CLK(clk), .Q(delay3_sram_waddr_d[5]) );
  DFFSSRX1_HVT delay4_sram_waddr_d_reg_5_ ( .D(1'b0), .SETB(n146), .RSTB(
        delay3_sram_waddr_d[5]), .CLK(clk), .Q(delay4_sram_waddr_d[5]) );
  DFFSSRX1_HVT sram_waddr_d_reg_5_ ( .D(1'b0), .SETB(n143), .RSTB(
        delay4_sram_waddr_d[5]), .CLK(clk), .Q(sram_waddr_d[5]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_4_ ( .D(1'b0), .SETB(n113), .RSTB(
        net19982), .CLK(net19989), .Q(delay1_sram_waddr_d[4]) );
  DFFSSRX1_HVT delay2_sram_waddr_d_reg_4_ ( .D(1'b0), .SETB(n139), .RSTB(
        delay1_sram_waddr_d[4]), .CLK(clk), .Q(delay2_sram_waddr_d[4]) );
  DFFSSRX1_HVT delay3_sram_waddr_d_reg_4_ ( .D(1'b0), .SETB(n101), .RSTB(
        delay2_sram_waddr_d[4]), .CLK(clk), .Q(delay3_sram_waddr_d[4]) );
  DFFSSRX1_HVT delay4_sram_waddr_d_reg_4_ ( .D(1'b0), .SETB(n156), .RSTB(
        delay3_sram_waddr_d[4]), .CLK(clk), .Q(delay4_sram_waddr_d[4]) );
  DFFSSRX1_HVT sram_waddr_d_reg_4_ ( .D(1'b0), .SETB(n100), .RSTB(
        delay4_sram_waddr_d[4]), .CLK(clk), .Q(sram_waddr_d[4]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_3_ ( .D(1'b0), .SETB(n114), .RSTB(
        net19983), .CLK(net19989), .Q(delay1_sram_waddr_d[3]) );
  DFFSSRX1_HVT delay2_sram_waddr_d_reg_3_ ( .D(1'b0), .SETB(n137), .RSTB(
        delay1_sram_waddr_d[3]), .CLK(clk), .Q(delay2_sram_waddr_d[3]) );
  DFFSSRX1_HVT delay3_sram_waddr_d_reg_3_ ( .D(1'b0), .SETB(n134), .RSTB(
        delay2_sram_waddr_d[3]), .CLK(clk), .Q(delay3_sram_waddr_d[3]) );
  DFFSSRX1_HVT delay4_sram_waddr_d_reg_3_ ( .D(1'b0), .SETB(n146), .RSTB(
        delay3_sram_waddr_d[3]), .CLK(clk), .Q(delay4_sram_waddr_d[3]) );
  DFFSSRX1_HVT sram_waddr_d_reg_3_ ( .D(1'b0), .SETB(n143), .RSTB(
        delay4_sram_waddr_d[3]), .CLK(clk), .Q(sram_waddr_d[3]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_2_ ( .D(1'b0), .SETB(n111), .RSTB(
        net19984), .CLK(net19989), .Q(delay1_sram_waddr_d[2]) );
  DFFSSRX1_HVT delay2_sram_waddr_d_reg_2_ ( .D(1'b0), .SETB(n139), .RSTB(
        delay1_sram_waddr_d[2]), .CLK(clk), .Q(delay2_sram_waddr_d[2]) );
  DFFSSRX1_HVT delay3_sram_waddr_d_reg_2_ ( .D(1'b0), .SETB(n134), .RSTB(
        delay2_sram_waddr_d[2]), .CLK(clk), .Q(delay3_sram_waddr_d[2]) );
  DFFSSRX1_HVT delay4_sram_waddr_d_reg_2_ ( .D(1'b0), .SETB(n146), .RSTB(
        delay3_sram_waddr_d[2]), .CLK(clk), .Q(delay4_sram_waddr_d[2]) );
  DFFSSRX1_HVT sram_waddr_d_reg_2_ ( .D(1'b0), .SETB(n143), .RSTB(
        delay4_sram_waddr_d[2]), .CLK(clk), .Q(sram_waddr_d[2]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_1_ ( .D(1'b0), .SETB(n138), .RSTB(
        net19985), .CLK(net19989), .Q(delay1_sram_waddr_d[1]) );
  DFFSSRX1_HVT delay2_sram_waddr_d_reg_1_ ( .D(1'b0), .SETB(n138), .RSTB(
        delay1_sram_waddr_d[1]), .CLK(clk), .Q(delay2_sram_waddr_d[1]) );
  DFFSSRX1_HVT delay3_sram_waddr_d_reg_1_ ( .D(1'b0), .SETB(n134), .RSTB(
        delay2_sram_waddr_d[1]), .CLK(clk), .Q(delay3_sram_waddr_d[1]) );
  DFFSSRX1_HVT delay4_sram_waddr_d_reg_1_ ( .D(1'b0), .SETB(n145), .RSTB(
        delay3_sram_waddr_d[1]), .CLK(clk), .Q(delay4_sram_waddr_d[1]) );
  DFFSSRX1_HVT sram_waddr_d_reg_1_ ( .D(1'b0), .SETB(n141), .RSTB(
        delay4_sram_waddr_d[1]), .CLK(clk), .Q(sram_waddr_d[1]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_0_ ( .D(1'b0), .SETB(n144), .RSTB(
        net19986), .CLK(net19989), .Q(delay1_sram_waddr_d[0]), .QN(n371) );
  DFFSSRX1_HVT delay2_sram_waddr_d_reg_0_ ( .D(1'b0), .SETB(n138), .RSTB(
        delay1_sram_waddr_d[0]), .CLK(clk), .Q(delay2_sram_waddr_d[0]) );
  DFFSSRX1_HVT delay3_sram_waddr_d_reg_0_ ( .D(1'b0), .SETB(n101), .RSTB(
        delay2_sram_waddr_d[0]), .CLK(clk), .Q(delay3_sram_waddr_d[0]) );
  DFFSSRX1_HVT delay4_sram_waddr_d_reg_0_ ( .D(1'b0), .SETB(n101), .RSTB(
        delay3_sram_waddr_d[0]), .CLK(clk), .Q(delay4_sram_waddr_d[0]) );
  DFFSSRX1_HVT sram_waddr_d_reg_0_ ( .D(1'b0), .SETB(n100), .RSTB(
        delay4_sram_waddr_d[0]), .CLK(clk), .Q(sram_waddr_d[0]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_9_ ( .D(1'b0), .SETB(n147), .RSTB(
        net19961), .CLK(net19973), .Q(delay1_sram_waddr_c[9]), .QN(n384) );
  DFFSSRX1_HVT delay2_sram_waddr_c_reg_9_ ( .D(1'b0), .SETB(n112), .RSTB(
        delay1_sram_waddr_c[9]), .CLK(clk), .Q(delay2_sram_waddr_c[9]) );
  DFFSSRX1_HVT delay3_sram_waddr_c_reg_9_ ( .D(1'b0), .SETB(n132), .RSTB(
        delay2_sram_waddr_c[9]), .CLK(clk), .Q(delay3_sram_waddr_c[9]) );
  DFFSSRX1_HVT delay4_sram_waddr_c_reg_9_ ( .D(1'b0), .SETB(n145), .RSTB(
        delay3_sram_waddr_c[9]), .CLK(clk), .Q(delay4_sram_waddr_c[9]) );
  DFFSSRX1_HVT sram_waddr_c_reg_9_ ( .D(1'b0), .SETB(n141), .RSTB(
        delay4_sram_waddr_c[9]), .CLK(clk), .Q(sram_waddr_c[9]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_8_ ( .D(1'b0), .SETB(n132), .RSTB(
        net19962), .CLK(net19973), .Q(delay1_sram_waddr_c[8]) );
  DFFSSRX1_HVT delay2_sram_waddr_c_reg_8_ ( .D(1'b0), .SETB(n138), .RSTB(
        delay1_sram_waddr_c[8]), .CLK(clk), .Q(delay2_sram_waddr_c[8]) );
  DFFSSRX1_HVT delay3_sram_waddr_c_reg_8_ ( .D(1'b0), .SETB(n132), .RSTB(
        delay2_sram_waddr_c[8]), .CLK(clk), .Q(delay3_sram_waddr_c[8]) );
  DFFSSRX1_HVT delay4_sram_waddr_c_reg_8_ ( .D(1'b0), .SETB(n145), .RSTB(
        delay3_sram_waddr_c[8]), .CLK(clk), .Q(delay4_sram_waddr_c[8]) );
  DFFSSRX1_HVT sram_waddr_c_reg_8_ ( .D(1'b0), .SETB(n141), .RSTB(
        delay4_sram_waddr_c[8]), .CLK(clk), .Q(sram_waddr_c[8]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_7_ ( .D(1'b0), .SETB(n136), .RSTB(
        net19963), .CLK(net19973), .Q(delay1_sram_waddr_c[7]) );
  DFFSSRX1_HVT delay2_sram_waddr_c_reg_7_ ( .D(1'b0), .SETB(n136), .RSTB(
        delay1_sram_waddr_c[7]), .CLK(clk), .Q(delay2_sram_waddr_c[7]) );
  DFFSSRX1_HVT delay3_sram_waddr_c_reg_7_ ( .D(1'b0), .SETB(n132), .RSTB(
        delay2_sram_waddr_c[7]), .CLK(clk), .Q(delay3_sram_waddr_c[7]) );
  DFFSSRX1_HVT delay4_sram_waddr_c_reg_7_ ( .D(1'b0), .SETB(n147), .RSTB(
        delay3_sram_waddr_c[7]), .CLK(clk), .Q(delay4_sram_waddr_c[7]) );
  DFFSSRX1_HVT sram_waddr_c_reg_7_ ( .D(1'b0), .SETB(n144), .RSTB(
        delay4_sram_waddr_c[7]), .CLK(clk), .Q(sram_waddr_c[7]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_6_ ( .D(1'b0), .SETB(n141), .RSTB(
        net19964), .CLK(net19973), .Q(delay1_sram_waddr_c[6]) );
  DFFSSRX1_HVT delay2_sram_waddr_c_reg_6_ ( .D(1'b0), .SETB(n136), .RSTB(
        delay1_sram_waddr_c[6]), .CLK(clk), .Q(delay2_sram_waddr_c[6]) );
  DFFSSRX1_HVT delay3_sram_waddr_c_reg_6_ ( .D(1'b0), .SETB(n111), .RSTB(
        delay2_sram_waddr_c[6]), .CLK(clk), .Q(delay3_sram_waddr_c[6]) );
  DFFSSRX1_HVT delay4_sram_waddr_c_reg_6_ ( .D(1'b0), .SETB(n114), .RSTB(
        delay3_sram_waddr_c[6]), .CLK(clk), .Q(delay4_sram_waddr_c[6]) );
  DFFSSRX1_HVT sram_waddr_c_reg_6_ ( .D(1'b0), .SETB(n113), .RSTB(
        delay4_sram_waddr_c[6]), .CLK(clk), .Q(sram_waddr_c[6]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_5_ ( .D(1'b0), .SETB(n145), .RSTB(
        net19965), .CLK(net19973), .Q(delay1_sram_waddr_c[5]) );
  DFFSSRX1_HVT delay2_sram_waddr_c_reg_5_ ( .D(1'b0), .SETB(n112), .RSTB(
        delay1_sram_waddr_c[5]), .CLK(clk), .Q(delay2_sram_waddr_c[5]) );
  DFFSSRX1_HVT delay3_sram_waddr_c_reg_5_ ( .D(1'b0), .SETB(n135), .RSTB(
        delay2_sram_waddr_c[5]), .CLK(clk), .Q(delay3_sram_waddr_c[5]) );
  DFFSSRX1_HVT delay4_sram_waddr_c_reg_5_ ( .D(1'b0), .SETB(n147), .RSTB(
        delay3_sram_waddr_c[5]), .CLK(clk), .Q(delay4_sram_waddr_c[5]) );
  DFFSSRX1_HVT sram_waddr_c_reg_5_ ( .D(1'b0), .SETB(n144), .RSTB(
        delay4_sram_waddr_c[5]), .CLK(clk), .Q(sram_waddr_c[5]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_4_ ( .D(1'b0), .SETB(n132), .RSTB(
        net19966), .CLK(net19973), .Q(delay1_sram_waddr_c[4]) );
  DFFSSRX1_HVT delay2_sram_waddr_c_reg_4_ ( .D(1'b0), .SETB(n136), .RSTB(
        delay1_sram_waddr_c[4]), .CLK(clk), .Q(delay2_sram_waddr_c[4]) );
  DFFSSRX1_HVT delay3_sram_waddr_c_reg_4_ ( .D(1'b0), .SETB(n135), .RSTB(
        delay2_sram_waddr_c[4]), .CLK(clk), .Q(delay3_sram_waddr_c[4]) );
  DFFSSRX1_HVT delay4_sram_waddr_c_reg_4_ ( .D(1'b0), .SETB(n147), .RSTB(
        delay3_sram_waddr_c[4]), .CLK(clk), .Q(delay4_sram_waddr_c[4]) );
  DFFSSRX1_HVT sram_waddr_c_reg_4_ ( .D(1'b0), .SETB(n144), .RSTB(
        delay4_sram_waddr_c[4]), .CLK(clk), .Q(sram_waddr_c[4]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_3_ ( .D(1'b0), .SETB(n136), .RSTB(
        net19967), .CLK(net19973), .Q(delay1_sram_waddr_c[3]) );
  DFFSSRX1_HVT delay2_sram_waddr_c_reg_3_ ( .D(1'b0), .SETB(n139), .RSTB(
        delay1_sram_waddr_c[3]), .CLK(clk), .Q(delay2_sram_waddr_c[3]) );
  DFFSSRX1_HVT delay3_sram_waddr_c_reg_3_ ( .D(1'b0), .SETB(n135), .RSTB(
        delay2_sram_waddr_c[3]), .CLK(clk), .Q(delay3_sram_waddr_c[3]) );
  DFFSSRX1_HVT delay4_sram_waddr_c_reg_3_ ( .D(1'b0), .SETB(n146), .RSTB(
        delay3_sram_waddr_c[3]), .CLK(clk), .Q(delay4_sram_waddr_c[3]) );
  DFFSSRX1_HVT sram_waddr_c_reg_3_ ( .D(1'b0), .SETB(n143), .RSTB(
        delay4_sram_waddr_c[3]), .CLK(clk), .Q(sram_waddr_c[3]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_2_ ( .D(1'b0), .SETB(n142), .RSTB(
        net19968), .CLK(net19973), .Q(delay1_sram_waddr_c[2]) );
  DFFSSRX1_HVT delay2_sram_waddr_c_reg_2_ ( .D(1'b0), .SETB(n139), .RSTB(
        delay1_sram_waddr_c[2]), .CLK(clk), .Q(delay2_sram_waddr_c[2]) );
  DFFSSRX1_HVT delay3_sram_waddr_c_reg_2_ ( .D(1'b0), .SETB(n101), .RSTB(
        delay2_sram_waddr_c[2]), .CLK(clk), .Q(delay3_sram_waddr_c[2]) );
  DFFSSRX1_HVT delay4_sram_waddr_c_reg_2_ ( .D(1'b0), .SETB(n133), .RSTB(
        delay3_sram_waddr_c[2]), .CLK(clk), .Q(delay4_sram_waddr_c[2]) );
  DFFSSRX1_HVT sram_waddr_c_reg_2_ ( .D(1'b0), .SETB(n100), .RSTB(
        delay4_sram_waddr_c[2]), .CLK(clk), .Q(sram_waddr_c[2]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_1_ ( .D(1'b0), .SETB(n101), .RSTB(
        net19969), .CLK(net19973), .Q(delay1_sram_waddr_c[1]) );
  DFFSSRX1_HVT delay2_sram_waddr_c_reg_1_ ( .D(1'b0), .SETB(n114), .RSTB(
        delay1_sram_waddr_c[1]), .CLK(clk), .Q(delay2_sram_waddr_c[1]) );
  DFFSSRX1_HVT delay3_sram_waddr_c_reg_1_ ( .D(1'b0), .SETB(n134), .RSTB(
        delay2_sram_waddr_c[1]), .CLK(clk), .Q(delay3_sram_waddr_c[1]) );
  DFFSSRX1_HVT delay4_sram_waddr_c_reg_1_ ( .D(1'b0), .SETB(n146), .RSTB(
        delay3_sram_waddr_c[1]), .CLK(clk), .Q(delay4_sram_waddr_c[1]) );
  DFFSSRX1_HVT sram_waddr_c_reg_1_ ( .D(1'b0), .SETB(n143), .RSTB(
        delay4_sram_waddr_c[1]), .CLK(clk), .Q(sram_waddr_c[1]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_0_ ( .D(1'b0), .SETB(n133), .RSTB(
        net19970), .CLK(net19973), .Q(delay1_sram_waddr_c[0]), .QN(n370) );
  DFFSSRX1_HVT delay2_sram_waddr_c_reg_0_ ( .D(1'b0), .SETB(n139), .RSTB(
        delay1_sram_waddr_c[0]), .CLK(clk), .Q(delay2_sram_waddr_c[0]) );
  DFFSSRX1_HVT delay3_sram_waddr_c_reg_0_ ( .D(1'b0), .SETB(n134), .RSTB(
        delay2_sram_waddr_c[0]), .CLK(clk), .Q(delay3_sram_waddr_c[0]) );
  DFFSSRX1_HVT delay4_sram_waddr_c_reg_0_ ( .D(1'b0), .SETB(n146), .RSTB(
        delay3_sram_waddr_c[0]), .CLK(clk), .Q(delay4_sram_waddr_c[0]) );
  DFFSSRX1_HVT sram_waddr_c_reg_0_ ( .D(1'b0), .SETB(n143), .RSTB(
        delay4_sram_waddr_c[0]), .CLK(clk), .Q(sram_waddr_c[0]) );
  DFFSSRX1_HVT delay_addr_change_reg_4_ ( .D(1'b0), .SETB(n138), .RSTB(
        addr_change[4]), .CLK(clk), .Q(delay_addr_change[4]) );
  DFFSSRX1_HVT delay_addr_change_reg_3_ ( .D(1'b0), .SETB(n134), .RSTB(
        addr_change[3]), .CLK(clk), .Q(delay_addr_change[3]) );
  DFFSSRX1_HVT delay_addr_change_reg_2_ ( .D(1'b0), .SETB(n145), .RSTB(
        addr_change[2]), .CLK(clk), .Q(delay_addr_change[2]) );
  DFFSSRX1_HVT delay2_addr_change_reg_4_ ( .D(1'b0), .SETB(n141), .RSTB(
        delay_addr_change[4]), .CLK(clk), .QN(n1152) );
  DFFSSRX1_HVT delay2_addr_change_reg_3_ ( .D(1'b0), .SETB(n138), .RSTB(
        delay_addr_change[3]), .CLK(clk), .Q(n357), .QN(n1153) );
  DFFSSRX1_HVT delay2_addr_change_reg_2_ ( .D(1'b0), .SETB(n101), .RSTB(
        delay_addr_change[2]), .CLK(clk), .Q(delay2_addr_change_2_), .QN(n353)
         );
  DFFSSRX1_HVT delay_channel_reg_4_ ( .D(1'b0), .SETB(n156), .RSTB(
        channel_cnt[4]), .CLK(clk), .Q(delay_channel[4]) );
  DFFSSRX1_HVT delay2_channel_reg_4_ ( .D(1'b0), .SETB(n100), .RSTB(
        delay_channel[4]), .CLK(clk), .Q(delay2_channel[4]) );
  DFFSSRX1_HVT channel_reg_4_ ( .D(1'b0), .SETB(n137), .RSTB(delay2_channel[4]), .CLK(clk), .Q(channel[4]) );
  DFFSSRX1_HVT delay_channel_reg_3_ ( .D(1'b0), .SETB(n132), .RSTB(
        channel_cnt[3]), .CLK(clk), .Q(delay_channel[3]) );
  DFFSSRX1_HVT delay2_channel_reg_3_ ( .D(1'b0), .SETB(n145), .RSTB(
        delay_channel[3]), .CLK(clk), .Q(delay2_channel[3]) );
  DFFSSRX1_HVT channel_reg_3_ ( .D(1'b0), .SETB(n141), .RSTB(delay2_channel[3]), .CLK(clk), .Q(channel[3]) );
  DFFSSRX1_HVT delay_channel_reg_2_ ( .D(1'b0), .SETB(n138), .RSTB(
        channel_cnt[2]), .CLK(clk), .Q(delay_channel[2]) );
  DFFSSRX1_HVT delay2_channel_reg_2_ ( .D(1'b0), .SETB(n132), .RSTB(
        delay_channel[2]), .CLK(clk), .Q(delay2_channel[2]) );
  DFFSSRX1_HVT channel_reg_2_ ( .D(1'b0), .SETB(n145), .RSTB(delay2_channel[2]), .CLK(clk), .Q(channel[2]) );
  DFFSSRX1_HVT delay_channel_reg_1_ ( .D(1'b0), .SETB(n141), .RSTB(
        channel_cnt[1]), .CLK(clk), .Q(delay_channel[1]) );
  DFFSSRX1_HVT delay2_channel_reg_1_ ( .D(1'b0), .SETB(n136), .RSTB(
        delay_channel[1]), .CLK(clk), .Q(delay2_channel[1]) );
  DFFSSRX1_HVT channel_reg_1_ ( .D(1'b0), .SETB(n132), .RSTB(delay2_channel[1]), .CLK(clk), .Q(channel[1]) );
  DFFSSRX1_HVT delay_channel_reg_0_ ( .D(1'b0), .SETB(n147), .RSTB(
        channel_cnt[0]), .CLK(clk), .Q(delay_channel[0]) );
  DFFSSRX1_HVT delay2_channel_reg_0_ ( .D(1'b0), .SETB(n144), .RSTB(
        delay_channel[0]), .CLK(clk), .Q(delay2_channel[0]) );
  DFFSSRX1_HVT channel_reg_0_ ( .D(1'b0), .SETB(n136), .RSTB(delay2_channel[0]), .CLK(clk), .Q(channel[0]) );
  DFFSSRX1_HVT sram_raddr_a7_reg_9_ ( .D(1'b0), .SETB(n137), .RSTB(
        n_sram_raddr_a7[9]), .CLK(net20494), .Q(sram_raddr_a7[9]) );
  DFFSSRX1_HVT sram_raddr_a7_reg_8_ ( .D(1'b0), .SETB(n100), .RSTB(
        n_sram_raddr_a7[8]), .CLK(net20494), .Q(sram_raddr_a7[8]) );
  DFFSSRX1_HVT sram_raddr_a7_reg_7_ ( .D(1'b0), .SETB(n156), .RSTB(
        n_sram_raddr_a7[7]), .CLK(net20494), .Q(sram_raddr_a7[7]) );
  DFFSSRX1_HVT sram_raddr_a7_reg_6_ ( .D(1'b0), .SETB(n101), .RSTB(
        n_sram_raddr_a7[6]), .CLK(net20494), .Q(sram_raddr_a7[6]) );
  DFFSSRX1_HVT sram_raddr_a7_reg_5_ ( .D(1'b0), .SETB(n138), .RSTB(
        n_sram_raddr_a7[5]), .CLK(net20494), .Q(sram_raddr_a7[5]), .QN(n313)
         );
  DFFSSRX1_HVT sram_raddr_a7_reg_4_ ( .D(1'b0), .SETB(n141), .RSTB(
        n_sram_raddr_a7[4]), .CLK(net20494), .Q(sram_raddr_a7[4]) );
  DFFSSRX1_HVT sram_raddr_a7_reg_3_ ( .D(1'b0), .SETB(n145), .RSTB(
        n_sram_raddr_a7[3]), .CLK(net20494), .Q(sram_raddr_a7[3]), .QN(n339)
         );
  DFFSSRX1_HVT sram_raddr_a7_reg_2_ ( .D(1'b0), .SETB(n134), .RSTB(
        n_sram_raddr_a7[2]), .CLK(net20494), .Q(sram_raddr_a7[2]) );
  DFFSSRX1_HVT sram_raddr_a7_reg_1_ ( .D(1'b0), .SETB(n138), .RSTB(
        n_sram_raddr_a7[1]), .CLK(net20494), .Q(sram_raddr_a7[1]), .QN(n214)
         );
  DFFSSRX1_HVT sram_raddr_a7_reg_0_ ( .D(1'b0), .SETB(n143), .RSTB(
        n_sram_raddr_a7[0]), .CLK(net20494), .Q(sram_raddr_a7[0]), .QN(n278)
         );
  DFFSSRX1_HVT sram_raddr_a8_reg_9_ ( .D(1'b0), .SETB(n146), .RSTB(
        n_sram_raddr_a8[9]), .CLK(net21821), .Q(sram_raddr_a8[9]) );
  DFFSSRX1_HVT sram_raddr_a8_reg_8_ ( .D(1'b0), .SETB(n134), .RSTB(
        n_sram_raddr_a8[8]), .CLK(net21821), .Q(sram_raddr_a8[8]) );
  DFFSSRX1_HVT sram_raddr_a8_reg_7_ ( .D(1'b0), .SETB(n137), .RSTB(
        n_sram_raddr_a8[7]), .CLK(net21821), .Q(sram_raddr_a8[7]) );
  DFFSSRX1_HVT sram_raddr_a8_reg_6_ ( .D(1'b0), .SETB(n142), .RSTB(
        n_sram_raddr_a8[6]), .CLK(net21821), .Q(sram_raddr_a8[6]), .QN(n338)
         );
  DFFSSRX1_HVT sram_raddr_a8_reg_5_ ( .D(1'b0), .SETB(n113), .RSTB(
        n_sram_raddr_a8[5]), .CLK(net21821), .Q(sram_raddr_a8[5]) );
  DFFSSRX1_HVT sram_raddr_a8_reg_4_ ( .D(1'b0), .SETB(n133), .RSTB(
        n_sram_raddr_a8[4]), .CLK(net21821), .Q(sram_raddr_a8[4]) );
  DFFSSRX1_HVT sram_raddr_a8_reg_3_ ( .D(1'b0), .SETB(n137), .RSTB(
        n_sram_raddr_a8[3]), .CLK(net21821), .Q(sram_raddr_a8[3]) );
  DFFSSRX1_HVT sram_raddr_a8_reg_2_ ( .D(1'b0), .SETB(n100), .RSTB(
        n_sram_raddr_a8[2]), .CLK(net21821), .Q(sram_raddr_a8[2]), .QN(n336)
         );
  DFFSSRX1_HVT sram_raddr_a8_reg_1_ ( .D(1'b0), .SETB(n113), .RSTB(
        n_sram_raddr_a8[1]), .CLK(net21821), .Q(sram_raddr_a8[1]) );
  DFFSSRX1_HVT sram_raddr_a8_reg_0_ ( .D(1'b0), .SETB(n101), .RSTB(
        n_sram_raddr_a8[0]), .CLK(net21821), .Q(sram_raddr_a8[0]), .QN(n229)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_9_ ( .D(1'b0), .SETB(n139), .RSTB(
        n_sram_raddr_a0[9]), .CLK(net23149), .Q(sram_raddr_a0[9]), .QN(n377)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_8_ ( .D(1'b0), .SETB(n143), .RSTB(
        n_sram_raddr_a0[8]), .CLK(net23149), .Q(sram_raddr_a0[8]), .QN(n375)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_7_ ( .D(1'b0), .SETB(n146), .RSTB(
        n_sram_raddr_a0[7]), .CLK(net23149), .Q(sram_raddr_a0[7]), .QN(n274)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_6_ ( .D(1'b0), .SETB(n135), .RSTB(
        n_sram_raddr_a0[6]), .CLK(net23149), .Q(sram_raddr_a0[6]), .QN(n329)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_5_ ( .D(1'b0), .SETB(n139), .RSTB(
        n_sram_raddr_a0[5]), .CLK(net23149), .Q(sram_raddr_a0[5]), .QN(n299)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_4_ ( .D(1'b0), .SETB(n144), .RSTB(
        n_sram_raddr_a0[4]), .CLK(net23149), .Q(sram_raddr_a0[4]), .QN(n290)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_3_ ( .D(1'b0), .SETB(n147), .RSTB(
        n_sram_raddr_a0[3]), .CLK(net23149), .Q(sram_raddr_a0[3]), .QN(n172)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_2_ ( .D(1'b0), .SETB(n135), .RSTB(
        n_sram_raddr_a0[2]), .CLK(net23149), .Q(sram_raddr_a0[2]), .QN(n204)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_1_ ( .D(1'b0), .SETB(n137), .RSTB(
        n_sram_raddr_a0[1]), .CLK(net23149), .Q(sram_raddr_a0[1]), .QN(n368)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_0_ ( .D(1'b0), .SETB(n142), .RSTB(
        n_sram_raddr_a0[0]), .CLK(net23149), .Q(sram_raddr_a0[0]), .QN(n359)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_9_ ( .D(1'b0), .SETB(n142), .RSTB(
        n_sram_raddr_a1[9]), .CLK(net20939), .Q(sram_raddr_a1[9]), .QN(n378)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_8_ ( .D(1'b0), .SETB(n133), .RSTB(
        n_sram_raddr_a1[8]), .CLK(net20939), .Q(sram_raddr_a1[8]), .QN(n376)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_7_ ( .D(1'b0), .SETB(n112), .RSTB(
        n_sram_raddr_a1[7]), .CLK(net20939), .Q(sram_raddr_a1[7]), .QN(n273)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_6_ ( .D(1'b0), .SETB(n113), .RSTB(
        n_sram_raddr_a1[6]), .CLK(net20939), .Q(sram_raddr_a1[6]), .QN(n294)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_5_ ( .D(1'b0), .SETB(n114), .RSTB(
        n_sram_raddr_a1[5]), .CLK(net20939), .Q(sram_raddr_a1[5]), .QN(n277)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_4_ ( .D(1'b0), .SETB(n111), .RSTB(
        n_sram_raddr_a1[4]), .CLK(net20939), .Q(sram_raddr_a1[4]), .QN(n200)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_3_ ( .D(1'b0), .SETB(n136), .RSTB(
        n_sram_raddr_a1[3]), .CLK(net20939), .Q(sram_raddr_a1[3]), .QN(n173)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_2_ ( .D(1'b0), .SETB(n144), .RSTB(
        n_sram_raddr_a1[2]), .CLK(net20939), .Q(sram_raddr_a1[2]), .QN(n165)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_1_ ( .D(1'b0), .SETB(n147), .RSTB(
        n_sram_raddr_a1[1]), .CLK(net20939), .Q(sram_raddr_a1[1]), .QN(n230)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_0_ ( .D(1'b0), .SETB(n132), .RSTB(
        n_sram_raddr_a1[0]), .CLK(net20939), .Q(sram_raddr_a1[0]), .QN(n362)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_9_ ( .D(1'b0), .SETB(n136), .RSTB(
        n_sram_raddr_a2[9]), .CLK(net22266), .Q(sram_raddr_a2[9]), .QN(n379)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_8_ ( .D(1'b0), .SETB(n141), .RSTB(
        n_sram_raddr_a2[8]), .CLK(net22266), .Q(sram_raddr_a2[8]), .QN(n326)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_7_ ( .D(1'b0), .SETB(n145), .RSTB(
        n_sram_raddr_a2[7]), .CLK(net22266), .Q(sram_raddr_a2[7]), .QN(n312)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_6_ ( .D(1'b0), .SETB(n132), .RSTB(
        n_sram_raddr_a2[6]), .CLK(net22266), .Q(sram_raddr_a2[6]), .QN(n323)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_5_ ( .D(1'b0), .SETB(n137), .RSTB(
        n_sram_raddr_a2[5]), .CLK(net22266), .Q(sram_raddr_a2[5]), .QN(n300)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_4_ ( .D(1'b0), .SETB(n142), .RSTB(
        n_sram_raddr_a2[4]), .CLK(net22266), .Q(sram_raddr_a2[4]), .QN(n283)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_3_ ( .D(1'b0), .SETB(n111), .RSTB(
        n_sram_raddr_a2[3]), .CLK(net22266), .Q(sram_raddr_a2[3]), .QN(n285)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_2_ ( .D(1'b0), .SETB(n133), .RSTB(
        n_sram_raddr_a2[2]), .CLK(net22266), .Q(sram_raddr_a2[2]), .QN(n334)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_1_ ( .D(1'b0), .SETB(n111), .RSTB(
        n_sram_raddr_a2[1]), .CLK(net22266), .Q(sram_raddr_a2[1]) );
  DFFSSRX1_HVT sram_raddr_a2_reg_0_ ( .D(1'b0), .SETB(n100), .RSTB(
        n_sram_raddr_a2[0]), .CLK(net22266), .Q(sram_raddr_a2[0]), .QN(n361)
         );
  DFFSSRX1_HVT sram_raddr_a3_reg_9_ ( .D(1'b0), .SETB(n156), .RSTB(
        n_sram_raddr_a3[9]), .CLK(net23595), .Q(sram_raddr_a3[9]) );
  DFFSSRX1_HVT sram_raddr_a3_reg_8_ ( .D(1'b0), .SETB(n101), .RSTB(
        n_sram_raddr_a3[8]), .CLK(net23595), .Q(sram_raddr_a3[8]) );
  DFFSSRX1_HVT sram_raddr_a3_reg_7_ ( .D(1'b0), .SETB(n138), .RSTB(
        n_sram_raddr_a3[7]), .CLK(net23595), .Q(sram_raddr_a3[7]), .QN(n271)
         );
  DFFSSRX1_HVT sram_raddr_a3_reg_6_ ( .D(1'b0), .SETB(n141), .RSTB(
        n_sram_raddr_a3[6]), .CLK(net23595), .Q(sram_raddr_a3[6]), .QN(n310)
         );
  DFFSSRX1_HVT sram_raddr_a3_reg_5_ ( .D(1'b0), .SETB(n145), .RSTB(
        n_sram_raddr_a3[5]), .CLK(net23595), .Q(sram_raddr_a3[5]), .QN(n289)
         );
  DFFSSRX1_HVT sram_raddr_a3_reg_4_ ( .D(1'b0), .SETB(n134), .RSTB(
        n_sram_raddr_a3[4]), .CLK(net23595), .Q(sram_raddr_a3[4]), .QN(n171)
         );
  DFFSSRX1_HVT sram_raddr_a3_reg_3_ ( .D(1'b0), .SETB(n138), .RSTB(
        n_sram_raddr_a3[3]), .CLK(net23595), .Q(sram_raddr_a3[3]), .QN(n205)
         );
  DFFSSRX1_HVT sram_raddr_a3_reg_2_ ( .D(1'b0), .SETB(n143), .RSTB(
        n_sram_raddr_a3[2]), .CLK(net23595), .Q(sram_raddr_a3[2]), .QN(n164)
         );
  DFFSSRX1_HVT sram_raddr_a3_reg_1_ ( .D(1'b0), .SETB(n146), .RSTB(
        n_sram_raddr_a3[1]), .CLK(net23595), .Q(sram_raddr_a3[1]) );
  DFFSSRX1_HVT sram_raddr_a3_reg_0_ ( .D(1'b0), .SETB(n134), .RSTB(
        n_sram_raddr_a3[0]), .CLK(net23595), .Q(sram_raddr_a3[0]), .QN(n360)
         );
  DFFSSRX1_HVT sram_raddr_a4_reg_9_ ( .D(1'b0), .SETB(n137), .RSTB(
        n_sram_raddr_a4[9]), .CLK(net21376), .Q(sram_raddr_a4[9]) );
  DFFSSRX1_HVT sram_raddr_a4_reg_8_ ( .D(1'b0), .SETB(n142), .RSTB(
        n_sram_raddr_a4[8]), .CLK(net21376), .Q(sram_raddr_a4[8]) );
  DFFSSRX1_HVT sram_raddr_a4_reg_7_ ( .D(1'b0), .SETB(n112), .RSTB(
        n_sram_raddr_a4[7]), .CLK(net21376), .Q(sram_raddr_a4[7]), .QN(n272)
         );
  DFFSSRX1_HVT sram_raddr_a4_reg_6_ ( .D(1'b0), .SETB(n133), .RSTB(
        n_sram_raddr_a4[6]), .CLK(net21376), .Q(sram_raddr_a4[6]), .QN(n317)
         );
  DFFSSRX1_HVT sram_raddr_a4_reg_5_ ( .D(1'b0), .SETB(n137), .RSTB(
        n_sram_raddr_a4[5]), .CLK(net21376), .Q(sram_raddr_a4[5]), .QN(n270)
         );
  DFFSSRX1_HVT sram_raddr_a4_reg_4_ ( .D(1'b0), .SETB(n100), .RSTB(
        n_sram_raddr_a4[4]), .CLK(net21376), .Q(sram_raddr_a4[4]), .QN(n311)
         );
  DFFSSRX1_HVT sram_raddr_a4_reg_3_ ( .D(1'b0), .SETB(n100), .RSTB(
        n_sram_raddr_a4[3]), .CLK(net21376), .Q(sram_raddr_a4[3]), .QN(n210)
         );
  DFFSSRX1_HVT sram_raddr_a4_reg_2_ ( .D(1'b0), .SETB(n101), .RSTB(
        n_sram_raddr_a4[2]), .CLK(net21376), .Q(sram_raddr_a4[2]), .QN(n174)
         );
  DFFSSRX1_HVT sram_raddr_a4_reg_1_ ( .D(1'b0), .SETB(n139), .RSTB(
        n_sram_raddr_a4[1]), .CLK(net21376), .Q(sram_raddr_a4[1]), .QN(n358)
         );
  DFFSSRX1_HVT sram_raddr_a4_reg_0_ ( .D(1'b0), .SETB(n143), .RSTB(
        n_sram_raddr_a4[0]), .CLK(net21376), .Q(sram_raddr_a4[0]), .QN(n212)
         );
  DFFSSRX1_HVT sram_raddr_a5_reg_9_ ( .D(1'b0), .SETB(n146), .RSTB(
        n_sram_raddr_a5[9]), .CLK(net22703), .Q(sram_raddr_a5[9]) );
  DFFSSRX1_HVT sram_raddr_a5_reg_8_ ( .D(1'b0), .SETB(n135), .RSTB(
        n_sram_raddr_a5[8]), .CLK(net22703), .Q(sram_raddr_a5[8]) );
  DFFSSRX1_HVT sram_raddr_a5_reg_7_ ( .D(1'b0), .SETB(n139), .RSTB(
        n_sram_raddr_a5[7]), .CLK(net22703), .Q(sram_raddr_a5[7]) );
  DFFSSRX1_HVT sram_raddr_a5_reg_6_ ( .D(1'b0), .SETB(n144), .RSTB(
        n_sram_raddr_a5[6]), .CLK(net22703), .Q(sram_raddr_a5[6]), .QN(n330)
         );
  DFFSSRX1_HVT sram_raddr_a5_reg_5_ ( .D(1'b0), .SETB(n147), .RSTB(
        n_sram_raddr_a5[5]), .CLK(net22703), .Q(sram_raddr_a5[5]), .QN(n327)
         );
  DFFSSRX1_HVT sram_raddr_a5_reg_4_ ( .D(1'b0), .SETB(n135), .RSTB(
        n_sram_raddr_a5[4]), .CLK(net22703), .Q(sram_raddr_a5[4]), .QN(n301)
         );
  DFFSSRX1_HVT sram_raddr_a5_reg_3_ ( .D(1'b0), .SETB(n137), .RSTB(
        n_sram_raddr_a5[3]), .CLK(net22703), .Q(sram_raddr_a5[3]), .QN(n201)
         );
  DFFSSRX1_HVT sram_raddr_a5_reg_2_ ( .D(1'b0), .SETB(n142), .RSTB(
        n_sram_raddr_a5[2]), .CLK(net22703), .Q(sram_raddr_a5[2]), .QN(n316)
         );
  DFFSSRX1_HVT sram_raddr_a5_reg_1_ ( .D(1'b0), .SETB(n133), .RSTB(
        n_sram_raddr_a5[1]), .CLK(net22703), .Q(sram_raddr_a5[1]) );
  DFFSSRX1_HVT sram_raddr_a5_reg_0_ ( .D(1'b0), .SETB(n133), .RSTB(
        n_sram_raddr_a5[0]), .CLK(net22703), .Q(sram_raddr_a5[0]), .QN(n373)
         );
  DFFSSRX1_HVT sram_raddr_a6_reg_9_ ( .D(1'b0), .SETB(n112), .RSTB(
        n_sram_raddr_a6[9]), .CLK(net24033), .Q(sram_raddr_a6[9]) );
  DFFSSRX1_HVT sram_raddr_a6_reg_8_ ( .D(1'b0), .SETB(n113), .RSTB(
        n_sram_raddr_a6[8]), .CLK(net24033), .Q(sram_raddr_a6[8]) );
  DFFSSRX1_HVT sram_raddr_a6_reg_7_ ( .D(1'b0), .SETB(n114), .RSTB(
        n_sram_raddr_a6[7]), .CLK(net24033), .Q(sram_raddr_a6[7]) );
  DFFSSRX1_HVT sram_raddr_a6_reg_6_ ( .D(1'b0), .SETB(n111), .RSTB(
        n_sram_raddr_a6[6]), .CLK(net24033), .Q(sram_raddr_a6[6]) );
  DFFSSRX1_HVT sram_raddr_a6_reg_5_ ( .D(1'b0), .SETB(n136), .RSTB(
        n_sram_raddr_a6[5]), .CLK(net24033), .Q(sram_raddr_a6[5]) );
  DFFSSRX1_HVT sram_raddr_a6_reg_4_ ( .D(1'b0), .SETB(n144), .RSTB(
        n_sram_raddr_a6[4]), .CLK(net24033), .Q(sram_raddr_a6[4]), .QN(n383)
         );
  DFFSSRX1_HVT sram_raddr_a6_reg_3_ ( .D(1'b0), .SETB(n147), .RSTB(
        n_sram_raddr_a6[3]), .CLK(net24033), .Q(sram_raddr_a6[3]) );
  DFFSSRX1_HVT sram_raddr_a6_reg_2_ ( .D(1'b0), .SETB(n132), .RSTB(
        n_sram_raddr_a6[2]), .CLK(net24033), .Q(sram_raddr_a6[2]), .QN(n337)
         );
  DFFSSRX1_HVT sram_raddr_a6_reg_1_ ( .D(1'b0), .SETB(n136), .RSTB(
        n_sram_raddr_a6[1]), .CLK(net24033), .Q(sram_raddr_a6[1]) );
  DFFSSRX1_HVT sram_raddr_a6_reg_0_ ( .D(1'b0), .SETB(n141), .RSTB(
        n_sram_raddr_a6[0]), .CLK(net24033), .Q(sram_raddr_a6[0]), .QN(n228)
         );
  DFFSSRX1_HVT sram_raddr_b7_reg_9_ ( .D(1'b0), .SETB(n145), .RSTB(
        n_sram_raddr_b7[9]), .CLK(net24567), .Q(sram_raddr_b7[9]), .QN(n281)
         );
  DFFSSRX1_HVT sram_raddr_b7_reg_8_ ( .D(1'b0), .SETB(n132), .RSTB(
        n_sram_raddr_b7[8]), .CLK(net24567), .Q(sram_raddr_b7[8]), .QN(n280)
         );
  DFFSSRX1_HVT sram_raddr_b7_reg_7_ ( .D(1'b0), .SETB(n137), .RSTB(
        n_sram_raddr_b7[7]), .CLK(net24567), .Q(sram_raddr_b7[7]), .QN(n198)
         );
  DFFSSRX1_HVT sram_raddr_b7_reg_6_ ( .D(1'b0), .SETB(n141), .RSTB(
        n_sram_raddr_b7[6]), .CLK(net24567), .Q(sram_raddr_b7[6]) );
  DFFSSRX1_HVT sram_raddr_b7_reg_5_ ( .D(1'b0), .SETB(n145), .RSTB(
        n_sram_raddr_b7[5]), .CLK(net24567), .Q(sram_raddr_b7[5]), .QN(n255)
         );
  DFFSSRX1_HVT sram_raddr_b7_reg_4_ ( .D(1'b0), .SETB(n132), .RSTB(
        n_sram_raddr_b7[4]), .CLK(net24567), .Q(sram_raddr_b7[4]) );
  DFFSSRX1_HVT sram_raddr_b7_reg_3_ ( .D(1'b0), .SETB(n100), .RSTB(
        n_sram_raddr_b7[3]), .CLK(net24567), .Q(sram_raddr_b7[3]), .QN(n304)
         );
  DFFSSRX1_HVT sram_raddr_b7_reg_2_ ( .D(1'b0), .SETB(n100), .RSTB(
        n_sram_raddr_b7[2]), .CLK(net24567), .Q(sram_raddr_b7[2]), .QN(n257)
         );
  DFFSSRX1_HVT sram_raddr_b7_reg_1_ ( .D(1'b0), .SETB(n156), .RSTB(
        n_sram_raddr_b7[1]), .CLK(net24567), .Q(sram_raddr_b7[1]) );
  DFFSSRX1_HVT sram_raddr_b7_reg_0_ ( .D(1'b0), .SETB(n101), .RSTB(
        n_sram_raddr_b7[0]), .CLK(net24567), .Q(sram_raddr_b7[0]), .QN(n308)
         );
  DFFSSRX1_HVT sram_raddr_b8_reg_9_ ( .D(1'b0), .SETB(n138), .RSTB(
        n_sram_raddr_b8[9]), .CLK(net25082), .Q(sram_raddr_b8[9]), .QN(n288)
         );
  DFFSSRX1_HVT sram_raddr_b8_reg_8_ ( .D(1'b0), .SETB(n141), .RSTB(
        n_sram_raddr_b8[8]), .CLK(net25082), .Q(sram_raddr_b8[8]), .QN(n260)
         );
  DFFSSRX1_HVT sram_raddr_b8_reg_7_ ( .D(1'b0), .SETB(n145), .RSTB(
        n_sram_raddr_b8[7]), .CLK(net25082), .Q(sram_raddr_b8[7]), .QN(n189)
         );
  DFFSSRX1_HVT sram_raddr_b8_reg_6_ ( .D(1'b0), .SETB(n134), .RSTB(
        n_sram_raddr_b8[6]), .CLK(net25082), .Q(sram_raddr_b8[6]) );
  DFFSSRX1_HVT sram_raddr_b8_reg_5_ ( .D(1'b0), .SETB(n138), .RSTB(
        n_sram_raddr_b8[5]), .CLK(net25082), .Q(sram_raddr_b8[5]), .QN(n256)
         );
  DFFSSRX1_HVT sram_raddr_b8_reg_4_ ( .D(1'b0), .SETB(n143), .RSTB(
        n_sram_raddr_b8[4]), .CLK(net25082), .Q(sram_raddr_b8[4]), .QN(n208)
         );
  DFFSSRX1_HVT sram_raddr_b8_reg_3_ ( .D(1'b0), .SETB(n146), .RSTB(
        n_sram_raddr_b8[3]), .CLK(net25082), .Q(sram_raddr_b8[3]), .QN(n305)
         );
  DFFSSRX1_HVT sram_raddr_b8_reg_2_ ( .D(1'b0), .SETB(n134), .RSTB(
        n_sram_raddr_b8[2]), .CLK(net25082), .Q(sram_raddr_b8[2]), .QN(n170)
         );
  DFFSSRX1_HVT sram_raddr_b8_reg_1_ ( .D(1'b0), .SETB(n137), .RSTB(
        n_sram_raddr_b8[1]), .CLK(net25082), .Q(sram_raddr_b8[1]) );
  DFFSSRX1_HVT sram_raddr_b8_reg_0_ ( .D(1'b0), .SETB(n143), .RSTB(
        n_sram_raddr_b8[0]), .CLK(net25082), .Q(sram_raddr_b8[0]), .QN(n309)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_9_ ( .D(1'b0), .SETB(n146), .RSTB(
        n_sram_raddr_b0[9]), .CLK(net25597), .Q(sram_raddr_b0[9]), .QN(n325)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_8_ ( .D(1'b0), .SETB(n134), .RSTB(
        n_sram_raddr_b0[8]), .CLK(net25597), .Q(sram_raddr_b0[8]), .QN(n314)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_7_ ( .D(1'b0), .SETB(n101), .RSTB(
        n_sram_raddr_b0[7]), .CLK(net25597), .Q(sram_raddr_b0[7]), .QN(n211)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_6_ ( .D(1'b0), .SETB(n100), .RSTB(
        n_sram_raddr_b0[6]), .CLK(net25597), .Q(sram_raddr_b0[6]), .QN(n262)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_5_ ( .D(1'b0), .SETB(n142), .RSTB(
        n_sram_raddr_b0[5]), .CLK(net25597), .Q(sram_raddr_b0[5]), .QN(n196)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_4_ ( .D(1'b0), .SETB(n101), .RSTB(
        n_sram_raddr_b0[4]), .CLK(net25597), .Q(sram_raddr_b0[4]), .QN(n251)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_3_ ( .D(1'b0), .SETB(n139), .RSTB(
        n_sram_raddr_b0[3]), .CLK(net25597), .Q(sram_raddr_b0[3]), .QN(n306)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_2_ ( .D(1'b0), .SETB(n143), .RSTB(
        n_sram_raddr_b0[2]), .CLK(net25597), .Q(sram_raddr_b0[2]), .QN(n259)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_1_ ( .D(1'b0), .SETB(n146), .RSTB(
        n_sram_raddr_b0[1]), .CLK(net25597), .Q(sram_raddr_b0[1]), .QN(n239)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_0_ ( .D(1'b0), .SETB(n135), .RSTB(
        n_sram_raddr_b0[0]), .CLK(net25597), .Q(sram_raddr_b0[0]), .QN(n184)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_9_ ( .D(1'b0), .SETB(n139), .RSTB(
        n_sram_raddr_b1[9]), .CLK(net26112), .Q(sram_raddr_b1[9]), .QN(n286)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_8_ ( .D(1'b0), .SETB(n144), .RSTB(
        n_sram_raddr_b1[8]), .CLK(net26112), .Q(sram_raddr_b1[8]), .QN(n191)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_7_ ( .D(1'b0), .SETB(n147), .RSTB(
        n_sram_raddr_b1[7]), .CLK(net26112), .Q(sram_raddr_b1[7]), .QN(n244)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_6_ ( .D(1'b0), .SETB(n135), .RSTB(
        n_sram_raddr_b1[6]), .CLK(net26112), .Q(sram_raddr_b1[6]), .QN(n266)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_5_ ( .D(1'b0), .SETB(n136), .RSTB(
        n_sram_raddr_b1[5]), .CLK(net26112), .Q(sram_raddr_b1[5]), .QN(n195)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_4_ ( .D(1'b0), .SETB(n144), .RSTB(
        n_sram_raddr_b1[4]), .CLK(net26112), .Q(sram_raddr_b1[4]), .QN(n250)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_3_ ( .D(1'b0), .SETB(n147), .RSTB(
        n_sram_raddr_b1[3]), .CLK(net26112), .Q(sram_raddr_b1[3]), .QN(n248)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_2_ ( .D(1'b0), .SETB(n135), .RSTB(
        n_sram_raddr_b1[2]), .CLK(net26112), .Q(sram_raddr_b1[2]), .QN(n188)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_1_ ( .D(1'b0), .SETB(n112), .RSTB(
        n_sram_raddr_b1[1]), .CLK(net26112), .Q(sram_raddr_b1[1]), .QN(n331)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_0_ ( .D(1'b0), .SETB(n113), .RSTB(
        n_sram_raddr_b1[0]), .CLK(net26112), .Q(sram_raddr_b1[0]), .QN(n175)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_9_ ( .D(1'b0), .SETB(n114), .RSTB(
        n_sram_raddr_b2[9]), .CLK(net26627), .Q(sram_raddr_b2[9]), .QN(n287)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_8_ ( .D(1'b0), .SETB(n111), .RSTB(
        n_sram_raddr_b2[8]), .CLK(net26627), .Q(sram_raddr_b2[8]), .QN(n192)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_7_ ( .D(1'b0), .SETB(n136), .RSTB(
        n_sram_raddr_b2[7]), .CLK(net26627), .Q(sram_raddr_b2[7]), .QN(n245)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_6_ ( .D(1'b0), .SETB(n144), .RSTB(
        n_sram_raddr_b2[6]), .CLK(net26627), .Q(sram_raddr_b2[6]), .QN(n267)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_5_ ( .D(1'b0), .SETB(n147), .RSTB(
        n_sram_raddr_b2[5]), .CLK(net26627), .Q(sram_raddr_b2[5]), .QN(n203)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_4_ ( .D(1'b0), .SETB(n132), .RSTB(
        n_sram_raddr_b2[4]), .CLK(net26627), .Q(sram_raddr_b2[4]), .QN(n297)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_3_ ( .D(1'b0), .SETB(n136), .RSTB(
        n_sram_raddr_b2[3]), .CLK(net26627), .Q(sram_raddr_b2[3]) );
  DFFSSRX1_HVT sram_raddr_b2_reg_2_ ( .D(1'b0), .SETB(n141), .RSTB(
        n_sram_raddr_b2[2]), .CLK(net26627), .Q(sram_raddr_b2[2]), .QN(n264)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_1_ ( .D(1'b0), .SETB(n145), .RSTB(
        n_sram_raddr_b2[1]), .CLK(net26627), .Q(sram_raddr_b2[1]), .QN(n238)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_0_ ( .D(1'b0), .SETB(n132), .RSTB(
        n_sram_raddr_b2[0]), .CLK(net26627), .Q(sram_raddr_b2[0]), .QN(n168)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_9_ ( .D(1'b0), .SETB(n138), .RSTB(
        n_sram_raddr_b3[9]), .CLK(net27142), .Q(sram_raddr_b3[9]), .QN(n279)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_8_ ( .D(1'b0), .SETB(n141), .RSTB(
        n_sram_raddr_b3[8]), .CLK(net27142), .Q(sram_raddr_b3[8]), .QN(n186)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_7_ ( .D(1'b0), .SETB(n145), .RSTB(
        n_sram_raddr_b3[7]), .CLK(net27142), .Q(sram_raddr_b3[7]), .QN(n243)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_6_ ( .D(1'b0), .SETB(n132), .RSTB(
        n_sram_raddr_b3[6]), .CLK(net27142), .Q(sram_raddr_b3[6]) );
  DFFSSRX1_HVT sram_raddr_b3_reg_5_ ( .D(1'b0), .SETB(n100), .RSTB(
        n_sram_raddr_b3[5]), .CLK(net27142), .Q(sram_raddr_b3[5]), .QN(n190)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_4_ ( .D(1'b0), .SETB(n100), .RSTB(
        n_sram_raddr_b3[4]), .CLK(net27142), .Q(sram_raddr_b3[4]), .QN(n253)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_3_ ( .D(1'b0), .SETB(n156), .RSTB(
        n_sram_raddr_b3[3]), .CLK(net27142), .Q(sram_raddr_b3[3]), .QN(n307)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_2_ ( .D(1'b0), .SETB(n101), .RSTB(
        n_sram_raddr_b3[2]), .CLK(net27142), .Q(sram_raddr_b3[2]), .QN(n249)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_1_ ( .D(1'b0), .SETB(n138), .RSTB(
        n_sram_raddr_b3[1]), .CLK(net27142), .Q(sram_raddr_b3[1]), .QN(n335)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_0_ ( .D(1'b0), .SETB(n141), .RSTB(
        n_sram_raddr_b3[0]), .CLK(net27142), .Q(sram_raddr_b3[0]), .QN(n215)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_9_ ( .D(1'b0), .SETB(n145), .RSTB(
        n_sram_raddr_b4[9]), .CLK(net27657), .Q(sram_raddr_b4[9]), .QN(n261)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_8_ ( .D(1'b0), .SETB(n134), .RSTB(
        n_sram_raddr_b4[8]), .CLK(net27657), .Q(sram_raddr_b4[8]), .QN(n265)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_7_ ( .D(1'b0), .SETB(n138), .RSTB(
        n_sram_raddr_b4[7]), .CLK(net27657), .Q(sram_raddr_b4[7]), .QN(n269)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_6_ ( .D(1'b0), .SETB(n143), .RSTB(
        n_sram_raddr_b4[6]), .CLK(net27657), .Q(sram_raddr_b4[6]), .QN(n263)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_5_ ( .D(1'b0), .SETB(n146), .RSTB(
        n_sram_raddr_b4[5]), .CLK(net27657), .Q(sram_raddr_b4[5]), .QN(n199)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_4_ ( .D(1'b0), .SETB(n134), .RSTB(
        n_sram_raddr_b4[4]), .CLK(net27657), .Q(sram_raddr_b4[4]), .QN(n284)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_3_ ( .D(1'b0), .SETB(n139), .RSTB(
        n_sram_raddr_b4[3]), .CLK(net27657), .Q(sram_raddr_b4[3]), .QN(n293)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_2_ ( .D(1'b0), .SETB(n143), .RSTB(
        n_sram_raddr_b4[2]), .CLK(net27657), .Q(sram_raddr_b4[2]), .QN(n246)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_1_ ( .D(1'b0), .SETB(n146), .RSTB(
        n_sram_raddr_b4[1]), .CLK(net27657), .Q(sram_raddr_b4[1]), .QN(n332)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_0_ ( .D(1'b0), .SETB(n134), .RSTB(
        n_sram_raddr_b4[0]), .CLK(net27657), .Q(sram_raddr_b4[0]), .QN(n206)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_9_ ( .D(1'b0), .SETB(n101), .RSTB(
        n_sram_raddr_b5[9]), .CLK(net28172), .Q(sram_raddr_b5[9]), .QN(n282)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_8_ ( .D(1'b0), .SETB(n100), .RSTB(
        n_sram_raddr_b5[8]), .CLK(net28172), .Q(sram_raddr_b5[8]), .QN(n187)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_7_ ( .D(1'b0), .SETB(n100), .RSTB(
        n_sram_raddr_b5[7]), .CLK(net28172), .Q(sram_raddr_b5[7]), .QN(n303)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_6_ ( .D(1'b0), .SETB(n101), .RSTB(
        n_sram_raddr_b5[6]), .CLK(net28172), .Q(sram_raddr_b5[6]), .QN(n295)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_5_ ( .D(1'b0), .SETB(n139), .RSTB(
        n_sram_raddr_b5[5]), .CLK(net28172), .Q(sram_raddr_b5[5]), .QN(n193)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_4_ ( .D(1'b0), .SETB(n143), .RSTB(
        n_sram_raddr_b5[4]), .CLK(net28172), .Q(sram_raddr_b5[4]), .QN(n252)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_3_ ( .D(1'b0), .SETB(n146), .RSTB(
        n_sram_raddr_b5[3]), .CLK(net28172), .Q(sram_raddr_b5[3]), .QN(n291)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_2_ ( .D(1'b0), .SETB(n135), .RSTB(
        n_sram_raddr_b5[2]), .CLK(net28172), .Q(sram_raddr_b5[2]), .QN(n247)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_1_ ( .D(1'b0), .SETB(n139), .RSTB(
        n_sram_raddr_b5[1]), .CLK(net28172), .Q(sram_raddr_b5[1]), .QN(n333)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_0_ ( .D(1'b0), .SETB(n144), .RSTB(
        n_sram_raddr_b5[0]), .CLK(net28172), .Q(sram_raddr_b5[0]), .QN(n207)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_9_ ( .D(1'b0), .SETB(n147), .RSTB(
        n_sram_raddr_b6[9]), .CLK(net28687), .Q(sram_raddr_b6[9]), .QN(n292)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_8_ ( .D(1'b0), .SETB(n135), .RSTB(
        n_sram_raddr_b6[8]), .CLK(net28687), .Q(sram_raddr_b6[8]), .QN(n258)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_7_ ( .D(1'b0), .SETB(n136), .RSTB(
        n_sram_raddr_b6[7]), .CLK(net28687), .Q(sram_raddr_b6[7]), .QN(n197)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_6_ ( .D(1'b0), .SETB(n144), .RSTB(
        n_sram_raddr_b6[6]), .CLK(net28687), .Q(sram_raddr_b6[6]) );
  DFFSSRX1_HVT sram_raddr_b6_reg_5_ ( .D(1'b0), .SETB(n147), .RSTB(
        n_sram_raddr_b6[5]), .CLK(net28687), .Q(sram_raddr_b6[5]), .QN(n254)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_4_ ( .D(1'b0), .SETB(n135), .RSTB(
        n_sram_raddr_b6[4]), .CLK(net28687), .Q(sram_raddr_b6[4]), .QN(n298)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_3_ ( .D(1'b0), .SETB(n112), .RSTB(
        n_sram_raddr_b6[3]), .CLK(net28687), .Q(sram_raddr_b6[3]), .QN(n202)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_2_ ( .D(1'b0), .SETB(n113), .RSTB(
        n_sram_raddr_b6[2]), .CLK(net28687), .Q(sram_raddr_b6[2]), .QN(n169)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_1_ ( .D(1'b0), .SETB(n114), .RSTB(
        n_sram_raddr_b6[1]), .CLK(net28687), .Q(sram_raddr_b6[1]) );
  DFFSSRX1_HVT sram_raddr_b6_reg_0_ ( .D(1'b0), .SETB(n111), .RSTB(
        n_sram_raddr_b6[0]), .CLK(net28687), .Q(sram_raddr_b6[0]), .QN(n322)
         );
  DFFSSRX1_HVT delay_sram_write_enable_b0_reg ( .D(n_sram_write_enable_b0), 
        .SETB(n105), .RSTB(1'b1), .CLK(clk), .Q(delay_sram_write_enable_b0) );
  DFFSSRX1_HVT delay_sram_write_enable_b1_reg ( .D(n_sram_write_enable_b1), 
        .SETB(n107), .RSTB(1'b1), .CLK(clk), .Q(delay_sram_write_enable_b1) );
  DFFSSRX1_HVT delay_sram_write_enable_b2_reg ( .D(n_sram_write_enable_b2), 
        .SETB(n106), .RSTB(1'b1), .CLK(clk), .Q(delay_sram_write_enable_b2) );
  DFFSSRX1_HVT delay_sram_write_enable_b3_reg ( .D(n_sram_write_enable_b3), 
        .SETB(n105), .RSTB(1'b1), .CLK(clk), .Q(delay_sram_write_enable_b3) );
  DFFSSRX1_HVT delay_sram_write_enable_b4_reg ( .D(n_sram_write_enable_b4), 
        .SETB(n107), .RSTB(1'b1), .CLK(clk), .Q(delay_sram_write_enable_b4) );
  DFFSSRX1_HVT delay_sram_write_enable_b5_reg ( .D(n_sram_write_enable_b5), 
        .SETB(n106), .RSTB(1'b1), .CLK(clk), .Q(delay_sram_write_enable_b5) );
  DFFSSRX1_HVT delay_sram_write_enable_b6_reg ( .D(n_sram_write_enable_b6), 
        .SETB(n105), .RSTB(1'b1), .CLK(clk), .Q(delay_sram_write_enable_b6) );
  DFFSSRX1_HVT delay_sram_write_enable_b7_reg ( .D(n_sram_write_enable_b7), 
        .SETB(n107), .RSTB(1'b1), .CLK(clk), .Q(delay_sram_write_enable_b7) );
  DFFSSRX1_HVT delay2_sram_write_enable_b7_reg ( .D(delay_sram_write_enable_b7), .SETB(n107), .RSTB(1'b1), .CLK(clk), .Q(delay2_sram_write_enable_b7) );
  DFFSSRX1_HVT sram_write_enable_b7_reg ( .D(delay2_sram_write_enable_b7), 
        .SETB(n107), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b7) );
  DFFSSRX1_HVT delay_sram_write_enable_b8_reg ( .D(n_sram_write_enable_b8), 
        .SETB(n107), .RSTB(1'b1), .CLK(clk), .Q(delay_sram_write_enable_b8) );
  DFFSSRX1_HVT delay2_sram_write_enable_b8_reg ( .D(delay_sram_write_enable_b8), .SETB(n107), .RSTB(1'b1), .CLK(clk), .Q(delay2_sram_write_enable_b8) );
  DFFSSRX1_HVT sram_write_enable_b8_reg ( .D(delay2_sram_write_enable_b8), 
        .SETB(n107), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b8) );
  DFFSSRX1_HVT delay2_sram_write_enable_b0_reg ( .D(delay_sram_write_enable_b0), .SETB(n106), .RSTB(1'b1), .CLK(clk), .Q(delay2_sram_write_enable_b0) );
  DFFSSRX1_HVT sram_write_enable_b0_reg ( .D(delay2_sram_write_enable_b0), 
        .SETB(n105), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b0) );
  DFFSSRX1_HVT delay2_sram_write_enable_b1_reg ( .D(delay_sram_write_enable_b1), .SETB(n106), .RSTB(1'b1), .CLK(clk), .Q(delay2_sram_write_enable_b1) );
  DFFSSRX1_HVT sram_write_enable_b1_reg ( .D(delay2_sram_write_enable_b1), 
        .SETB(n107), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b1) );
  DFFSSRX1_HVT delay2_sram_write_enable_b2_reg ( .D(delay_sram_write_enable_b2), .SETB(n105), .RSTB(1'b1), .CLK(clk), .Q(delay2_sram_write_enable_b2) );
  DFFSSRX1_HVT sram_write_enable_b2_reg ( .D(delay2_sram_write_enable_b2), 
        .SETB(n106), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b2) );
  DFFSSRX1_HVT delay2_sram_write_enable_b3_reg ( .D(delay_sram_write_enable_b3), .SETB(n105), .RSTB(1'b1), .CLK(clk), .Q(delay2_sram_write_enable_b3) );
  DFFSSRX1_HVT sram_write_enable_b3_reg ( .D(delay2_sram_write_enable_b3), 
        .SETB(n107), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b3) );
  DFFSSRX1_HVT delay2_sram_write_enable_b4_reg ( .D(delay_sram_write_enable_b4), .SETB(n106), .RSTB(1'b1), .CLK(clk), .Q(delay2_sram_write_enable_b4) );
  DFFSSRX1_HVT sram_write_enable_b4_reg ( .D(delay2_sram_write_enable_b4), 
        .SETB(n105), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b4) );
  DFFSSRX1_HVT delay2_sram_write_enable_b5_reg ( .D(delay_sram_write_enable_b5), .SETB(n106), .RSTB(1'b1), .CLK(clk), .Q(delay2_sram_write_enable_b5) );
  DFFSSRX1_HVT sram_write_enable_b5_reg ( .D(delay2_sram_write_enable_b5), 
        .SETB(n107), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b5) );
  DFFSSRX1_HVT delay2_sram_write_enable_b6_reg ( .D(delay_sram_write_enable_b6), .SETB(n105), .RSTB(1'b1), .CLK(clk), .Q(delay2_sram_write_enable_b6) );
  DFFSSRX1_HVT sram_write_enable_b6_reg ( .D(delay2_sram_write_enable_b6), 
        .SETB(n106), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b6) );
  DFFSSRX1_HVT delay_sram_write_enable_d3_reg ( .D(n_sram_write_enable_d3), 
        .SETB(n105), .RSTB(1'b1), .CLK(clk), .Q(delay_sram_write_enable_d3) );
  DFFSSRX1_HVT delay_sram_write_enable_d4_reg ( .D(n_sram_write_enable_d4), 
        .SETB(n107), .RSTB(1'b1), .CLK(clk), .Q(delay_sram_write_enable_d4) );
  DFFSSRX1_HVT sram_write_enable_d3_reg ( .D(delay_sram_write_enable_d3), 
        .SETB(n106), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_d3) );
  DFFSSRX1_HVT sram_write_enable_d4_reg ( .D(delay_sram_write_enable_d4), 
        .SETB(n105), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_d4) );
  DFFSSRX1_HVT delay_sram_write_enable_c0_reg ( .D(n_sram_write_enable_c0), 
        .SETB(n106), .RSTB(1'b1), .CLK(clk), .Q(delay_sram_write_enable_c0) );
  DFFSSRX1_HVT sram_write_enable_c0_reg ( .D(delay_sram_write_enable_c0), 
        .SETB(n107), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_c0) );
  DFFSSRX1_HVT delay_sram_write_enable_c1_reg ( .D(n_sram_write_enable_c1), 
        .SETB(n105), .RSTB(1'b1), .CLK(clk), .Q(delay_sram_write_enable_c1) );
  DFFSSRX1_HVT sram_write_enable_c1_reg ( .D(delay_sram_write_enable_c1), 
        .SETB(n106), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_c1) );
  DFFSSRX1_HVT delay_sram_write_enable_c2_reg ( .D(n_sram_write_enable_c2), 
        .SETB(n105), .RSTB(1'b1), .CLK(clk), .Q(delay_sram_write_enable_c2) );
  DFFSSRX1_HVT sram_write_enable_c2_reg ( .D(delay_sram_write_enable_c2), 
        .SETB(n107), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_c2) );
  DFFSSRX1_HVT delay_sram_write_enable_c3_reg ( .D(n_sram_write_enable_c3), 
        .SETB(n106), .RSTB(1'b1), .CLK(clk), .Q(delay_sram_write_enable_c3) );
  DFFSSRX1_HVT sram_write_enable_c3_reg ( .D(delay_sram_write_enable_c3), 
        .SETB(n105), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_c3) );
  DFFSSRX1_HVT delay_sram_write_enable_c4_reg ( .D(n_sram_write_enable_c4), 
        .SETB(n106), .RSTB(1'b1), .CLK(clk), .Q(delay_sram_write_enable_c4) );
  DFFSSRX1_HVT sram_write_enable_c4_reg ( .D(delay_sram_write_enable_c4), 
        .SETB(n107), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_c4) );
  DFFSSRX1_HVT delay_sram_write_enable_d0_reg ( .D(n_sram_write_enable_d0), 
        .SETB(n105), .RSTB(1'b1), .CLK(clk), .Q(delay_sram_write_enable_d0) );
  DFFSSRX1_HVT sram_write_enable_d0_reg ( .D(delay_sram_write_enable_d0), 
        .SETB(n106), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_d0) );
  DFFSSRX1_HVT delay_sram_write_enable_d1_reg ( .D(n_sram_write_enable_d1), 
        .SETB(n105), .RSTB(1'b1), .CLK(clk), .Q(delay_sram_write_enable_d1) );
  DFFSSRX1_HVT sram_write_enable_d1_reg ( .D(delay_sram_write_enable_d1), 
        .SETB(n107), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_d1) );
  DFFSSRX1_HVT delay_sram_write_enable_d2_reg ( .D(n_sram_write_enable_d2), 
        .SETB(n106), .RSTB(1'b1), .CLK(clk), .Q(delay_sram_write_enable_d2) );
  DFFSSRX1_HVT sram_write_enable_d2_reg ( .D(delay_sram_write_enable_d2), 
        .SETB(n106), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_d2) );
  AO221X1_HVT U3 ( .A1(1'b1), .A2(n1604), .A3(n230), .A4(n362), .A5(n80), .Y(
        n82) );
  AO222X1_HVT U4 ( .A1(sram_raddr_b0[3]), .A2(n162), .A3(n43), .A4(n781), .A5(
        1'b1), .A6(n49), .Y(n_sram_raddr_b0[3]) );
  AO221X1_HVT U5 ( .A1(1'b1), .A2(n1974), .A3(n1972), .A4(n1363), .A5(n74), 
        .Y(n76) );
  AO221X1_HVT U6 ( .A1(1'b1), .A2(n1868), .A3(n1867), .A4(n1827), .A5(n50), 
        .Y(n_sram_raddr_a3[8]) );
  AO221X1_HVT U7 ( .A1(1'b1), .A2(n1916), .A3(n1913), .A4(n94), .A5(n39), .Y(
        n_sram_raddr_a4[8]) );
  AO221X1_HVT U8 ( .A1(1'b1), .A2(n1963), .A3(n1962), .A4(n94), .A5(n32), .Y(
        n_sram_raddr_a5[8]) );
  AO221X1_HVT U9 ( .A1(1'b1), .A2(n1133), .A3(n1263), .A4(sram_raddr_b4[4]), 
        .A5(n27), .Y(n29) );
  AO221X1_HVT U10 ( .A1(1'b1), .A2(n1081), .A3(n1074), .A4(n197), .A5(n4), .Y(
        n6) );
  OA221X1_HVT U11 ( .A1(1'b0), .A2(n1543), .A3(col[2]), .A4(n1542), .A5(n1541), 
        .Y(net19704) );
  OA221X1_HVT U12 ( .A1(1'b0), .A2(n129), .A3(addr_change[0]), .A4(
        addr_change[1]), .A5(n1535), .Y(net20009) );
  OA221X1_HVT U13 ( .A1(1'b0), .A2(n1522), .A3(n1510), .A4(
        delay1_sram_waddr_d[8]), .A5(n1509), .Y(net19978) );
  OA221X1_HVT U14 ( .A1(1'b0), .A2(n1507), .A3(n1495), .A4(
        delay1_sram_waddr_c[8]), .A5(n1494), .Y(net19962) );
  OA21X1_HVT U15 ( .A1(sram_raddr_b0[2]), .A2(sram_raddr_b0[3]), .A3(n150), 
        .Y(n43) );
  OA221X1_HVT U16 ( .A1(1'b0), .A2(n998), .A3(sram_raddr_b0[6]), .A4(n800), 
        .A5(n809), .Y(n1071) );
  OA221X1_HVT U17 ( .A1(1'b0), .A2(n1533), .A3(addr_change[3]), .A4(n70), .A5(
        n1532), .Y(net20007) );
  OA221X1_HVT U18 ( .A1(1'b0), .A2(n1522), .A3(n1512), .A4(
        delay1_sram_waddr_d[7]), .A5(n1511), .Y(net19979) );
  OA221X1_HVT U19 ( .A1(1'b0), .A2(n1507), .A3(n1497), .A4(
        delay1_sram_waddr_c[7]), .A5(n1496), .Y(net19963) );
  OA221X1_HVT U20 ( .A1(1'b0), .A2(n1528), .A3(channel_cnt[1]), .A4(
        channel_cnt[0]), .A5(n1527), .Y(net19997) );
  OA221X1_HVT U21 ( .A1(1'b0), .A2(n1522), .A3(n1514), .A4(
        delay1_sram_waddr_d[6]), .A5(n1513), .Y(net19980) );
  OA221X1_HVT U22 ( .A1(1'b0), .A2(n1507), .A3(n1499), .A4(
        delay1_sram_waddr_c[6]), .A5(n1498), .Y(net19964) );
  OA221X1_HVT U23 ( .A1(1'b0), .A2(n1522), .A3(n1516), .A4(
        delay1_sram_waddr_d[5]), .A5(n1515), .Y(net19981) );
  OA221X1_HVT U24 ( .A1(1'b0), .A2(n1507), .A3(n1501), .A4(
        delay1_sram_waddr_c[5]), .A5(n1500), .Y(net19965) );
  OA221X1_HVT U25 ( .A1(1'b0), .A2(n1522), .A3(n1518), .A4(
        delay1_sram_waddr_d[4]), .A5(n1517), .Y(net19982) );
  OA221X1_HVT U26 ( .A1(1'b0), .A2(n1507), .A3(n1503), .A4(
        delay1_sram_waddr_c[4]), .A5(n1502), .Y(net19966) );
  OA221X1_HVT U27 ( .A1(1'b0), .A2(n1522), .A3(delay1_sram_waddr_d[3]), .A4(
        n24), .A5(n1519), .Y(net19983) );
  OA221X1_HVT U28 ( .A1(1'b0), .A2(n1507), .A3(delay1_sram_waddr_c[3]), .A4(
        n23), .A5(n1504), .Y(net19967) );
  OA221X1_HVT U29 ( .A1(1'b0), .A2(n99), .A3(sram_raddr_b2[8]), .A4(n1339), 
        .A5(n739), .Y(n744) );
  OA221X1_HVT U30 ( .A1(1'b0), .A2(n1522), .A3(delay1_sram_waddr_d[2]), .A4(
        n11), .A5(n1520), .Y(net19984) );
  OA221X1_HVT U31 ( .A1(1'b0), .A2(n1507), .A3(delay1_sram_waddr_c[2]), .A4(n9), .A5(n1505), .Y(net19968) );
  OA221X1_HVT U32 ( .A1(1'b0), .A2(n1296), .A3(sram_raddr_b1[8]), .A4(n1339), 
        .A5(n647), .Y(n652) );
  INVX1_HVT U33 ( .A(n1811), .Y(n96) );
  NAND2X2_HVT U34 ( .A1(n1296), .A2(n1339), .Y(n1270) );
  NAND2X2_HVT U35 ( .A1(n493), .A2(n1334), .Y(n1443) );
  OAI21X1_HVT U37 ( .A1(n1800), .A2(n1796), .A3(n1881), .Y(n1930) );
  NAND2X0_HVT U38 ( .A1(n1076), .A2(n1096), .Y(n2) );
  AO221X1_HVT U39 ( .A1(n1078), .A2(n243), .A3(n1078), .A4(n1073), .A5(n155), 
        .Y(n3) );
  AND3X1_HVT U40 ( .A1(n1080), .A2(sram_raddr_b6[7]), .A3(n124), .Y(n4) );
  NAND4X0_HVT U42 ( .A1(n1075), .A2(n2), .A3(n3), .A4(n6), .Y(n7) );
  AO222X1_HVT U43 ( .A1(n7), .A2(n129), .A3(n197), .A4(n1090), .A5(
        sram_raddr_b6[7]), .A6(n1087), .Y(n_sram_raddr_b6[7]) );
  INVX0_HVT U45 ( .A(n1506), .Y(n9) );
  INVX0_HVT U47 ( .A(n1521), .Y(n11) );
  NAND2X0_HVT U49 ( .A1(n1096), .A2(n1097), .Y(n13) );
  AO22X1_HVT U50 ( .A1(n124), .A2(n1092), .A3(n258), .A4(n1091), .Y(n14) );
  AO22X1_HVT U51 ( .A1(n292), .A2(n1093), .A3(sram_raddr_b6[9]), .A4(n14), .Y(
        n15) );
  INVX0_HVT U52 ( .A(n1094), .Y(n16) );
  AO221X1_HVT U53 ( .A1(n1094), .A2(n279), .A3(n16), .A4(sram_raddr_b3[9]), 
        .A5(n110), .Y(n17) );
  NAND4X0_HVT U54 ( .A1(n1095), .A2(n13), .A3(n15), .A4(n17), .Y(n18) );
  AND3X1_HVT U55 ( .A1(sram_raddr_b6[8]), .A2(n1090), .A3(sram_raddr_b6[7]), 
        .Y(n19) );
  AO222X1_HVT U56 ( .A1(n18), .A2(n130), .A3(sram_raddr_b6[9]), .A4(n1098), 
        .A5(n292), .A6(n19), .Y(n_sram_raddr_b6[9]) );
  AO21X1_HVT U57 ( .A1(sram_raddr_a3[8]), .A2(n1866), .A3(n1869), .Y(n20) );
  AO222X1_HVT U58 ( .A1(n20), .A2(n1945), .A3(n1871), .A4(n1867), .A5(
        sram_raddr_a6[8]), .A6(n109), .Y(n21) );
  OR2X1_HVT U59 ( .A1(n1868), .A2(n21), .Y(n_sram_raddr_a6[8]) );
  INVX0_HVT U61 ( .A(n1505), .Y(n23) );
  INVX0_HVT U62 ( .A(n1520), .Y(n24) );
  NAND2X0_HVT U64 ( .A1(n875), .A2(n882), .Y(n26) );
  AO22X1_HVT U65 ( .A1(n873), .A2(n910), .A3(n1183), .A4(n26), .Y(n27) );
  INVX0_HVT U67 ( .A(n26), .Y(n30) );
  AO222X1_HVT U68 ( .A1(n29), .A2(n130), .A3(n30), .A4(n150), .A5(
        sram_raddr_b4[4]), .A6(n161), .Y(n_sram_raddr_b4[4]) );
  AO22X1_HVT U70 ( .A1(n1967), .A2(sram_raddr_a5[8]), .A3(n1830), .A4(n1826), 
        .Y(n32) );
  NAND2X0_HVT U73 ( .A1(sram_raddr_b3[2]), .A2(n1263), .Y(n35) );
  NAND4X0_HVT U74 ( .A1(n1023), .A2(n770), .A3(n767), .A4(n35), .Y(n36) );
  AO21X1_HVT U75 ( .A1(n768), .A2(n825), .A3(n36), .Y(n37) );
  AO222X1_HVT U76 ( .A1(n37), .A2(n130), .A3(sram_raddr_b3[2]), .A4(n162), 
        .A5(n249), .A6(n103), .Y(n_sram_raddr_b3[2]) );
  AO22X1_HVT U78 ( .A1(n1920), .A2(sram_raddr_a4[8]), .A3(n1787), .A4(n1784), 
        .Y(n39) );
  NAND4X0_HVT U81 ( .A1(state[0]), .A2(n1109), .A3(n232), .A4(n177), .Y(n42)
         );
  AO21X1_HVT U82 ( .A1(n1363), .A2(n42), .A3(n159), .Y(net19836) );
  AO21X1_HVT U83 ( .A1(n123), .A2(n505), .A3(n306), .Y(n44) );
  NAND2X0_HVT U84 ( .A1(n259), .A2(n1077), .Y(n45) );
  NAND4X0_HVT U85 ( .A1(n306), .A2(n688), .A3(n511), .A4(n45), .Y(n46) );
  NAND3X0_HVT U86 ( .A1(n775), .A2(n44), .A3(n46), .Y(n48) );
  OA221X1_HVT U87 ( .A1(n48), .A2(n771), .A3(n48), .A4(n1239), .A5(n119), .Y(
        n49) );
  AO22X1_HVT U88 ( .A1(n109), .A2(sram_raddr_a3[8]), .A3(n1751), .A4(n1748), 
        .Y(n50) );
  INVX0_HVT U92 ( .A(n1484), .Y(n54) );
  OA21X1_HVT U93 ( .A1(delay1_sram_waddr_b[2]), .A2(n54), .A3(n1488), .Y(n55)
         );
  AO21X1_HVT U94 ( .A1(n1485), .A2(delay1_sram_waddr_b[2]), .A3(n1483), .Y(n56) );
  AO22X1_HVT U95 ( .A1(n1482), .A2(n55), .A3(n1487), .A4(n56), .Y(net19945) );
  INVX0_HVT U97 ( .A(n1546), .Y(n58) );
  NAND3X0_HVT U98 ( .A1(n179), .A2(row[3]), .A3(n58), .Y(n457) );
  AND3X1_HVT U99 ( .A1(n250), .A2(n124), .A3(n867), .Y(n59) );
  OA22X1_HVT U100 ( .A1(n59), .A2(n846), .A3(n658), .A4(n614), .Y(n60) );
  OA22X1_HVT U101 ( .A1(n195), .A2(n60), .A3(n879), .A4(n154), .Y(n61) );
  NAND3X0_HVT U102 ( .A1(n878), .A2(n616), .A3(n61), .Y(n62) );
  NAND2X0_HVT U103 ( .A1(n622), .A2(n195), .Y(n63) );
  AND2X1_HVT U104 ( .A1(n63), .A2(n623), .Y(n64) );
  AO222X1_HVT U105 ( .A1(n62), .A2(n130), .A3(sram_raddr_b1[5]), .A4(n160), 
        .A5(n102), .A6(n64), .Y(n_sram_raddr_b1[5]) );
  NAND2X0_HVT U106 ( .A1(n1951), .A2(sram_raddr_a5[6]), .Y(n65) );
  NAND2X0_HVT U107 ( .A1(n1954), .A2(n65), .Y(n66) );
  AO222X1_HVT U108 ( .A1(n66), .A2(n1945), .A3(n1965), .A4(n1952), .A5(
        sram_raddr_a8[6]), .A6(n1967), .Y(n67) );
  OR2X1_HVT U109 ( .A1(n1953), .A2(n67), .Y(n_sram_raddr_a8[6]) );
  AND3X1_HVT U112 ( .A1(addr_change[0]), .A2(addr_change[2]), .A3(
        addr_change[1]), .Y(n70) );
  INVX0_HVT U114 ( .A(n464), .Y(n72) );
  NAND3X0_HVT U115 ( .A1(n1972), .A2(n1977), .A3(n72), .Y(n73) );
  INVX0_HVT U116 ( .A(n1973), .Y(n74) );
  NAND3X0_HVT U118 ( .A1(n1730), .A2(n73), .A3(n76), .Y(n_box_sel_1_) );
  OA22X1_HVT U121 ( .A1(n230), .A2(n1895), .A3(n115), .A4(n1757), .Y(n79) );
  INVX0_HVT U122 ( .A(n1640), .Y(n80) );
  NAND3X0_HVT U124 ( .A1(n79), .A2(n1756), .A3(n82), .Y(n_sram_raddr_a1[1]) );
  AO21X1_HVT U125 ( .A1(sram_raddr_a5[8]), .A2(n1961), .A3(n1964), .Y(n83) );
  AO222X1_HVT U126 ( .A1(n83), .A2(n95), .A3(n1965), .A4(n1962), .A5(
        sram_raddr_a8[8]), .A6(n1967), .Y(n84) );
  OR2X1_HVT U127 ( .A1(n1963), .A2(n84), .Y(n_sram_raddr_a8[8]) );
  AND2X1_HVT U131 ( .A1(n1476), .A2(n1488), .Y(n88) );
  AO21X1_HVT U132 ( .A1(delay1_sram_waddr_b[3]), .A2(n1479), .A3(
        delay1_sram_waddr_b[4]), .Y(n89) );
  AO221X1_HVT U133 ( .A1(delay1_sram_waddr_b[4]), .A2(delay1_sram_waddr_b[3]), 
        .A3(delay1_sram_waddr_b[4]), .A4(n1478), .A5(n1477), .Y(n90) );
  AO22X1_HVT U134 ( .A1(n88), .A2(n89), .A3(n1487), .A4(n90), .Y(net19939) );
  AO21X1_HVT U135 ( .A1(channel_cnt[2]), .A2(n1526), .A3(channel_cnt[3]), .Y(
        n91) );
  AND3X1_HVT U136 ( .A1(n1528), .A2(n1525), .A3(n91), .Y(net19995) );
  NAND4X0_HVT U138 ( .A1(weight_cnt[2]), .A2(n275), .A3(n227), .A4(n354), .Y(
        n93) );
  NOR3X0_HVT U139 ( .A1(conv1_done), .A2(n469), .A3(n93), .Y(n_conv1_done) );
  INVX8_HVT U140 ( .A(srstn), .Y(n104) );
  INVX8_HVT U141 ( .A(n104), .Y(n107) );
  INVX8_HVT U142 ( .A(n104), .Y(n105) );
  INVX4_HVT U143 ( .A(n104), .Y(n106) );
  INVX1_HVT U144 ( .A(n106), .Y(n156) );
  INVX1_HVT U145 ( .A(n1924), .Y(n94) );
  AOI22X1_HVT U146 ( .A1(n1872), .A2(n1871), .A3(n1945), .A4(n1870), .Y(n1873)
         );
  INVX0_HVT U147 ( .A(n1961), .Y(n1955) );
  INVX1_HVT U148 ( .A(n161), .Y(n99) );
  INVX1_HVT U149 ( .A(n1239), .Y(n110) );
  INVX2_HVT U150 ( .A(n116), .Y(n95) );
  INVX0_HVT U151 ( .A(n117), .Y(n129) );
  INVX0_HVT U152 ( .A(n1364), .Y(n1420) );
  INVX1_HVT U153 ( .A(n1339), .Y(n103) );
  INVX2_HVT U154 ( .A(n156), .Y(n97) );
  INVX1_HVT U155 ( .A(n117), .Y(n1536) );
  INVX1_HVT U156 ( .A(n1419), .Y(n1423) );
  INVX1_HVT U157 ( .A(n1241), .Y(n1238) );
  OAI221X1_HVT U158 ( .A1(n486), .A2(n179), .A3(n486), .A4(n234), .A5(n598), 
        .Y(n1301) );
  INVX1_HVT U159 ( .A(n1042), .Y(n1040) );
  INVX1_HVT U160 ( .A(n1537), .Y(n98) );
  INVX0_HVT U161 ( .A(n1367), .Y(n1370) );
  INVX0_HVT U162 ( .A(n1969), .Y(n386) );
  INVX0_HVT U163 ( .A(n1833), .Y(n398) );
  INVX0_HVT U164 ( .A(n1754), .Y(n403) );
  INVX0_HVT U165 ( .A(n1371), .Y(n1372) );
  INVX0_HVT U166 ( .A(n996), .Y(n1008) );
  INVX0_HVT U167 ( .A(n652), .Y(n650) );
  INVX0_HVT U168 ( .A(n1494), .Y(n1493) );
  INVX0_HVT U169 ( .A(n839), .Y(n840) );
  INVX0_HVT U170 ( .A(n744), .Y(n742) );
  INVX0_HVT U171 ( .A(n1509), .Y(n1508) );
  INVX0_HVT U172 ( .A(n722), .Y(n707) );
  INVX0_HVT U173 ( .A(n1790), .Y(n400) );
  INVX0_HVT U174 ( .A(n1596), .Y(n1597) );
  INVX0_HVT U175 ( .A(n1922), .Y(n389) );
  INVX0_HVT U176 ( .A(n1705), .Y(n1706) );
  INVX0_HVT U177 ( .A(n1874), .Y(n392) );
  INVX0_HVT U178 ( .A(n612), .Y(n607) );
  INVX0_HVT U179 ( .A(n523), .Y(n514) );
  INVX0_HVT U180 ( .A(n1640), .Y(n1613) );
  INVX0_HVT U181 ( .A(n1925), .Y(n1926) );
  INVX0_HVT U182 ( .A(n1918), .Y(n1894) );
  INVX0_HVT U183 ( .A(n642), .Y(n659) );
  NOR2X1_HVT U184 ( .A1(n1961), .A2(sram_raddr_a5[8]), .Y(n1964) );
  INVX0_HVT U185 ( .A(n1590), .Y(n1557) );
  INVX0_HVT U186 ( .A(n981), .Y(n982) );
  INVX0_HVT U187 ( .A(n1707), .Y(n1708) );
  INVX0_HVT U188 ( .A(n1434), .Y(n1422) );
  INVX0_HVT U189 ( .A(n1698), .Y(n1670) );
  INVX0_HVT U190 ( .A(n628), .Y(n658) );
  INVX0_HVT U191 ( .A(n1592), .Y(n1593) );
  INVX0_HVT U192 ( .A(n1719), .Y(n405) );
  INVX1_HVT U193 ( .A(n1742), .Y(n108) );
  INVX0_HVT U194 ( .A(n733), .Y(n751) );
  INVX0_HVT U195 ( .A(n999), .Y(n1000) );
  INVX0_HVT U196 ( .A(n1305), .Y(n1306) );
  INVX0_HVT U197 ( .A(n917), .Y(n918) );
  INVX0_HVT U198 ( .A(n1700), .Y(n1701) );
  INVX1_HVT U199 ( .A(n154), .Y(n1239) );
  INVX0_HVT U200 ( .A(n1646), .Y(n1647) );
  INVX0_HVT U201 ( .A(n831), .Y(n832) );
  INVX1_HVT U202 ( .A(n140), .Y(n113) );
  INVX1_HVT U203 ( .A(n131), .Y(n112) );
  INVX1_HVT U204 ( .A(n131), .Y(n111) );
  INVX1_HVT U205 ( .A(n97), .Y(n114) );
  INVX0_HVT U206 ( .A(n1648), .Y(n1649) );
  INVX0_HVT U207 ( .A(n1598), .Y(n1599) );
  INVX1_HVT U208 ( .A(n98), .Y(n119) );
  INVX0_HVT U209 ( .A(n1702), .Y(n1703) );
  NOR2X1_HVT U210 ( .A1(n1462), .A2(n1461), .Y(n1466) );
  INVX1_HVT U211 ( .A(n1945), .Y(n115) );
  INVX0_HVT U212 ( .A(n1433), .Y(net19715) );
  INVX1_HVT U213 ( .A(n1945), .Y(n116) );
  INVX0_HVT U214 ( .A(n1408), .Y(n1404) );
  INVX0_HVT U215 ( .A(n544), .Y(n546) );
  INVX1_HVT U216 ( .A(n1210), .Y(n121) );
  INVX1_HVT U217 ( .A(n1210), .Y(n120) );
  INVX1_HVT U218 ( .A(n1210), .Y(n122) );
  INVX0_HVT U219 ( .A(n647), .Y(n638) );
  INVX0_HVT U220 ( .A(n739), .Y(n729) );
  INVX2_HVT U221 ( .A(n140), .Y(n100) );
  INVX2_HVT U222 ( .A(n131), .Y(n101) );
  INVX0_HVT U223 ( .A(n1853), .Y(n1855) );
  INVX0_HVT U224 ( .A(n1096), .Y(n1045) );
  INVX2_HVT U225 ( .A(n1339), .Y(n102) );
  INVX0_HVT U226 ( .A(n1194), .Y(n846) );
  NOR2X1_HVT U227 ( .A1(n1912), .A2(sram_raddr_a4[8]), .Y(n1917) );
  INVX0_HVT U228 ( .A(n1642), .Y(n1643) );
  INVX0_HVT U229 ( .A(n1876), .Y(n1884) );
  INVX0_HVT U230 ( .A(n879), .Y(n880) );
  INVX0_HVT U231 ( .A(n1226), .Y(n1288) );
  INVX0_HVT U232 ( .A(n1583), .Y(n1584) );
  INVX0_HVT U233 ( .A(n1078), .Y(n1079) );
  INVX0_HVT U234 ( .A(n631), .Y(n617) );
  AND2X1_HVT U235 ( .A1(n1544), .A2(n178), .Y(n1811) );
  INVX0_HVT U236 ( .A(n1341), .Y(n478) );
  INVX1_HVT U237 ( .A(n117), .Y(n128) );
  NOR2X1_HVT U238 ( .A1(n271), .A2(n1582), .Y(n1594) );
  INVX0_HVT U239 ( .A(n1686), .Y(n1692) );
  NOR2X1_HVT U240 ( .A1(n272), .A2(n1632), .Y(n1644) );
  NOR2X0_HVT U241 ( .A1(conv1_weight_done), .A2(n1735), .Y(n1945) );
  NOR2X1_HVT U242 ( .A1(n1414), .A2(sram_raddr_weight[5]), .Y(n1417) );
  INVX0_HVT U243 ( .A(n1196), .Y(n1202) );
  INVX1_HVT U244 ( .A(n117), .Y(n127) );
  AND3X1_HVT U245 ( .A1(n490), .A2(n237), .A3(n183), .Y(n998) );
  INVX1_HVT U246 ( .A(n1296), .Y(n161) );
  INVX1_HVT U247 ( .A(n1339), .Y(n148) );
  AND4X1_HVT U248 ( .A1(row[0]), .A2(n490), .A3(n489), .A4(n167), .Y(n1304) );
  INVX1_HVT U249 ( .A(n1296), .Y(n160) );
  INVX1_HVT U250 ( .A(n1339), .Y(n150) );
  INVX1_HVT U251 ( .A(n1339), .Y(n149) );
  INVX1_HVT U252 ( .A(n156), .Y(n131) );
  INVX1_HVT U253 ( .A(n156), .Y(n140) );
  INVX0_HVT U254 ( .A(n1633), .Y(n1634) );
  INVX0_HVT U255 ( .A(n1354), .Y(n1357) );
  INVX0_HVT U256 ( .A(n1577), .Y(n1578) );
  INVX0_HVT U257 ( .A(n976), .Y(n968) );
  INVX0_HVT U258 ( .A(n1274), .Y(n1262) );
  INVX0_HVT U259 ( .A(n1907), .Y(n1911) );
  INVX0_HVT U260 ( .A(n1923), .Y(n1957) );
  INVX0_HVT U261 ( .A(n893), .Y(n884) );
  NOR2X1_HVT U262 ( .A1(n1866), .A2(sram_raddr_a3[8]), .Y(n1869) );
  INVX0_HVT U263 ( .A(n1301), .Y(n125) );
  INVX0_HVT U264 ( .A(n491), .Y(n490) );
  INVX0_HVT U265 ( .A(n1687), .Y(n1694) );
  INVX0_HVT U266 ( .A(n636), .Y(n648) );
  NOR2X1_HVT U267 ( .A1(n98), .A2(addr_change[0]), .Y(net20010) );
  INVX0_HVT U268 ( .A(n1467), .Y(n1468) );
  INVX0_HVT U269 ( .A(n603), .Y(n604) );
  INVX0_HVT U270 ( .A(n515), .Y(n516) );
  INVX0_HVT U271 ( .A(n904), .Y(n419) );
  INVX0_HVT U272 ( .A(n608), .Y(n609) );
  INVX0_HVT U273 ( .A(n1976), .Y(n1971) );
  INVX0_HVT U274 ( .A(n464), .Y(n1974) );
  INVX0_HVT U275 ( .A(n1975), .Y(n1978) );
  INVX0_HVT U276 ( .A(n1525), .Y(n1524) );
  INVX0_HVT U277 ( .A(n549), .Y(n558) );
  INVX0_HVT U278 ( .A(n693), .Y(n694) );
  INVX0_HVT U279 ( .A(n1127), .Y(n1129) );
  INVX0_HVT U280 ( .A(n727), .Y(n740) );
  INVX0_HVT U281 ( .A(n1017), .Y(n472) );
  INVX0_HVT U282 ( .A(n1134), .Y(n1138) );
  INVX0_HVT U283 ( .A(n965), .Y(n966) );
  INVX0_HVT U284 ( .A(n698), .Y(n699) );
  INVX0_HVT U285 ( .A(n1934), .Y(n1939) );
  INVX1_HVT U286 ( .A(n1537), .Y(n118) );
  INVX1_HVT U287 ( .A(n1537), .Y(n117) );
  INVX0_HVT U288 ( .A(n1554), .Y(n1559) );
  INVX0_HVT U289 ( .A(n1726), .Y(n1729) );
  INVX0_HVT U290 ( .A(n1125), .Y(n1124) );
  INVX0_HVT U291 ( .A(n1532), .Y(n1531) );
  INVX0_HVT U292 ( .A(n1552), .Y(n1553) );
  INVX0_HVT U293 ( .A(n506), .Y(n500) );
  INVX0_HVT U294 ( .A(n1273), .Y(n408) );
  INVX0_HVT U295 ( .A(n503), .Y(n498) );
  INVX0_HVT U296 ( .A(n1527), .Y(n1526) );
  INVX0_HVT U297 ( .A(n536), .Y(n783) );
  INVX0_HVT U298 ( .A(n1345), .Y(n1346) );
  INVX0_HVT U299 ( .A(n1441), .Y(n1738) );
  INVX0_HVT U300 ( .A(n681), .Y(n676) );
  INVX0_HVT U301 ( .A(n1541), .Y(n1361) );
  INVX0_HVT U302 ( .A(n1765), .Y(n1766) );
  INVX0_HVT U303 ( .A(n1609), .Y(n1610) );
  INVX0_HVT U304 ( .A(n1843), .Y(n1844) );
  INVX0_HVT U305 ( .A(n1166), .Y(n411) );
  INVX0_HVT U306 ( .A(n622), .Y(n869) );
  INVX0_HVT U307 ( .A(n1431), .Y(n1418) );
  INVX0_HVT U308 ( .A(n592), .Y(n586) );
  INVX0_HVT U309 ( .A(n1072), .Y(n415) );
  INVX0_HVT U310 ( .A(n1660), .Y(n1661) );
  INVX0_HVT U311 ( .A(n1449), .Y(n1451) );
  INVX0_HVT U312 ( .A(n1333), .Y(n1739) );
  INVX0_HVT U313 ( .A(mode[0]), .Y(n461) );
  INVX0_HVT U314 ( .A(mode[1]), .Y(n463) );
  AND3X1_HVT U315 ( .A1(state[0]), .A2(state[1]), .A3(n1445), .Y(n1537) );
  INVX0_HVT U316 ( .A(n1742), .Y(n109) );
  INVX1_HVT U317 ( .A(n131), .Y(n133) );
  INVX1_HVT U318 ( .A(n97), .Y(n137) );
  INVX1_HVT U319 ( .A(n140), .Y(n142) );
  AND2X1_HVT U320 ( .A1(mode[1]), .A2(n461), .Y(n1324) );
  INVX1_HVT U321 ( .A(n1301), .Y(n126) );
  INVX1_HVT U322 ( .A(n118), .Y(n130) );
  INVX0_HVT U323 ( .A(n1301), .Y(n123) );
  INVX0_HVT U324 ( .A(n1301), .Y(n124) );
  INVX2_HVT U325 ( .A(n131), .Y(n132) );
  INVX2_HVT U326 ( .A(n131), .Y(n134) );
  INVX2_HVT U327 ( .A(n131), .Y(n135) );
  INVX2_HVT U328 ( .A(n97), .Y(n136) );
  INVX2_HVT U329 ( .A(n97), .Y(n138) );
  INVX2_HVT U330 ( .A(n97), .Y(n139) );
  INVX2_HVT U331 ( .A(n140), .Y(n141) );
  INVX2_HVT U332 ( .A(n140), .Y(n143) );
  INVX2_HVT U333 ( .A(n140), .Y(n144) );
  INVX2_HVT U334 ( .A(n97), .Y(n145) );
  INVX2_HVT U335 ( .A(n97), .Y(n146) );
  INVX2_HVT U336 ( .A(n97), .Y(n147) );
  INVX1_HVT U337 ( .A(n1811), .Y(n151) );
  INVX1_HVT U338 ( .A(n998), .Y(n152) );
  INVX1_HVT U339 ( .A(n998), .Y(n153) );
  INVX1_HVT U340 ( .A(n1304), .Y(n154) );
  INVX1_HVT U341 ( .A(n1304), .Y(n155) );
  INVX1_HVT U342 ( .A(n105), .Y(n157) );
  INVX2_HVT U343 ( .A(n107), .Y(n158) );
  INVX2_HVT U344 ( .A(srstn), .Y(n159) );
  OAI21X1_HVT U345 ( .A1(n1546), .A2(n491), .A3(n1523), .Y(n1296) );
  INVX0_HVT U346 ( .A(n1296), .Y(n162) );
  INVX1_HVT U347 ( .A(n1363), .Y(n1979) );
  OR2X1_HVT U348 ( .A1(n493), .A2(n492), .Y(n1339) );
  INVX1_HVT U349 ( .A(n1249), .Y(n1284) );
  INVX1_HVT U350 ( .A(n1895), .Y(n1920) );
  NOR2X0_HVT U351 ( .A1(n232), .A2(n1109), .Y(n1445) );
  OR3X1_HVT U352 ( .A1(row[0]), .A2(n489), .A3(n491), .Y(n1210) );
  INVX1_HVT U353 ( .A(n126), .Y(n1263) );
  OA221X1_HVT U354 ( .A1(n1539), .A2(n1135), .A3(n1539), .A4(
        addr_col_sel_cnt[0]), .A5(n1538), .Y(n1895) );
  NAND4X0_HVT U355 ( .A1(state[0]), .A2(state[1]), .A3(n1108), .A4(n1109), .Y(
        n1363) );
  INVX1_HVT U356 ( .A(n1461), .Y(n1488) );
  INVX1_HVT U357 ( .A(n1458), .Y(n1487) );
  INVX1_HVT U358 ( .A(n1360), .Y(n1543) );
  INVX1_HVT U359 ( .A(n1142), .Y(n1183) );
  INVX1_HVT U360 ( .A(n1052), .Y(n1077) );
  OA221X1_HVT U361 ( .A1(n1539), .A2(n1136), .A3(n1539), .A4(
        addr_col_sel_cnt[1]), .A5(n1538), .Y(n1805) );
  OAI21X1_HVT U362 ( .A1(n178), .A2(n1334), .A3(n1342), .Y(n_conv1_weight_done) );
  INVX1_HVT U363 ( .A(mem_sel), .Y(n1492) );
  AO221X1_HVT U364 ( .A1(sram_raddr_a2[4]), .A2(n1810), .A3(n283), .A4(n1806), 
        .A5(n96), .Y(n1942) );
  AO221X1_HVT U365 ( .A1(n1815), .A2(n1812), .A3(n1815), .A4(n300), .A5(n96), 
        .Y(n1948) );
  AO221X1_HVT U366 ( .A1(sram_raddr_a1[6]), .A2(n1779), .A3(n294), .A4(n1774), 
        .A5(n96), .Y(n1904) );
  AO221X1_HVT U367 ( .A1(sram_raddr_a1[4]), .A2(n1766), .A3(n200), .A4(n1765), 
        .A5(n151), .Y(n1891) );
  AO221X1_HVT U368 ( .A1(n1783), .A2(n1780), .A3(n1783), .A4(n273), .A5(n96), 
        .Y(n1909) );
  AO221X1_HVT U369 ( .A1(sram_raddr_a0[5]), .A2(n1729), .A3(n299), .A4(n1726), 
        .A5(n151), .Y(n1851) );
  AO221X1_HVT U370 ( .A1(sram_raddr_a0[7]), .A2(n1746), .A3(n274), .A4(n1743), 
        .A5(n96), .Y(n1864) );
  AO221X1_HVT U371 ( .A1(n1726), .A2(n1721), .A3(n1726), .A4(n290), .A5(n151), 
        .Y(n1846) );
  INVX2_HVT U372 ( .A(n96), .Y(n1881) );
  OAI21X1_HVT U373 ( .A1(sram_raddr_a4[4]), .A2(n1615), .A3(n1622), .Y(n1764)
         );
  INVX1_HVT U374 ( .A(n1443), .Y(n1435) );
  OAI21X1_HVT U375 ( .A1(sram_raddr_a4[6]), .A2(n1626), .A3(n1632), .Y(n1773)
         );
  OAI21X1_HVT U376 ( .A1(sram_raddr_a3[6]), .A2(n1575), .A3(n1582), .Y(n1734)
         );
  OAI21X1_HVT U377 ( .A1(n724), .A2(n189), .A3(n733), .Y(n1280) );
  OAI21X1_HVT U378 ( .A1(n633), .A2(n198), .A3(n642), .Y(n1177) );
  OAI21X1_HVT U379 ( .A1(n1376), .A2(n320), .A3(n1375), .Y(n1379) );
  NAND2X0_HVT U380 ( .A1(n151), .A2(n1876), .Y(n1640) );
  AOI221X1_HVT U381 ( .A1(n1590), .A2(n172), .A3(n1590), .A4(n1558), .A5(n109), 
        .Y(n1566) );
  NAND2X0_HVT U382 ( .A1(n96), .A2(n1853), .Y(n1590) );
  AO22X1_HVT U383 ( .A1(write_col[1]), .A2(n1324), .A3(write_row[0]), .A4(
        n1329), .Y(n484) );
  AND2X1_HVT U384 ( .A1(n129), .A2(n1530), .Y(n1533) );
  AO21X1_HVT U385 ( .A1(n1454), .A2(n1453), .A3(n1489), .Y(n1461) );
  NAND2X0_HVT U386 ( .A1(n119), .A2(n1420), .Y(n1434) );
  NAND2X0_HVT U387 ( .A1(n129), .A2(n1364), .Y(n1433) );
  NAND4X0_HVT U388 ( .A1(addr_row_sel_cnt[0]), .A2(n1137), .A3(n1545), .A4(
        n1979), .Y(n1735) );
  AND2X1_HVT U389 ( .A1(n1329), .A2(write_enable), .Y(n1447) );
  INVX1_HVT U390 ( .A(n1336), .Y(n1523) );
  NAND2X0_HVT U391 ( .A1(channel_cnt[1]), .A2(channel_cnt[0]), .Y(n1527) );
  NAND2X0_HVT U392 ( .A1(row[1]), .A2(row[0]), .Y(n1546) );
  INVX2_HVT U393 ( .A(n1805), .Y(n1967) );
  INVX1_HVT U394 ( .A(n1653), .Y(n1545) );
  NAND2X0_HVT U395 ( .A1(col[1]), .A2(col[0]), .Y(n486) );
  INVX1_HVT U396 ( .A(n493), .Y(n1528) );
  AND2X1_HVT U397 ( .A1(n127), .A2(mem_sel), .Y(n1522) );
  AND2X1_HVT U398 ( .A1(n1537), .A2(n1492), .Y(n1507) );
  NAND3X0_HVT U399 ( .A1(n488), .A2(n179), .A3(n234), .Y(n491) );
  AND3X1_HVT U400 ( .A1(n1542), .A2(n163), .A3(n167), .Y(n488) );
  NOR4X1_HVT U401 ( .A1(delay2_addr_change_2_), .A2(n1152), .A3(n357), .A4(
        n1325), .Y(n1328) );
  INVX1_HVT U402 ( .A(n484), .Y(n485) );
  NOR4X1_HVT U403 ( .A1(channel_cnt[1]), .A2(channel_cnt[4]), .A3(
        conv2_weight_done), .A4(n470), .Y(n471) );
  INVX1_HVT U404 ( .A(n1472), .Y(n1477) );
  INVX1_HVT U405 ( .A(n1478), .Y(n1483) );
  INVX1_HVT U406 ( .A(n1511), .Y(n1510) );
  INVX1_HVT U407 ( .A(n1513), .Y(n1512) );
  INVX1_HVT U408 ( .A(n1515), .Y(n1514) );
  INVX1_HVT U409 ( .A(n1517), .Y(n1516) );
  INVX1_HVT U410 ( .A(n1519), .Y(n1518) );
  INVX1_HVT U411 ( .A(n1496), .Y(n1495) );
  INVX1_HVT U412 ( .A(n1498), .Y(n1497) );
  INVX1_HVT U413 ( .A(n1500), .Y(n1499) );
  INVX1_HVT U414 ( .A(n1502), .Y(n1501) );
  INVX1_HVT U415 ( .A(n1504), .Y(n1503) );
  INVX1_HVT U416 ( .A(n1469), .Y(n1465) );
  INVX1_HVT U417 ( .A(n1476), .Y(n1473) );
  INVX1_HVT U418 ( .A(n1482), .Y(n1479) );
  INVX1_HVT U419 ( .A(n1830), .Y(n1804) );
  NAND2X0_HVT U420 ( .A1(n1924), .A2(n1923), .Y(n1965) );
  INVX1_HVT U421 ( .A(n1946), .Y(n1950) );
  INVX1_HVT U422 ( .A(n1828), .Y(n1829) );
  INVX1_HVT U423 ( .A(n1825), .Y(n1824) );
  INVX1_HVT U424 ( .A(n1820), .Y(n1819) );
  INVX1_HVT U425 ( .A(n1806), .Y(n1810) );
  INVX1_HVT U426 ( .A(n1787), .Y(n1778) );
  INVX1_HVT U427 ( .A(n1605), .Y(n1606) );
  INVX1_HVT U428 ( .A(n1751), .Y(n1741) );
  INVX1_HVT U429 ( .A(n1896), .Y(n1901) );
  INVX1_HVT U430 ( .A(n1785), .Y(n1786) );
  INVX1_HVT U431 ( .A(n1774), .Y(n1779) );
  INVX1_HVT U432 ( .A(n1749), .Y(n1750) );
  INVX1_HVT U433 ( .A(n1743), .Y(n1746) );
  INVX1_HVT U434 ( .A(n1856), .Y(n1861) );
  INVX1_HVT U435 ( .A(n1827), .Y(n1924) );
  INVX1_HVT U436 ( .A(n1051), .Y(n1038) );
  INVX1_HVT U437 ( .A(n1074), .Y(n1066) );
  INVX1_HVT U438 ( .A(n1285), .Y(n1286) );
  INVX1_HVT U439 ( .A(n1178), .Y(n1182) );
  INVX1_HVT U440 ( .A(n1184), .Y(n1185) );
  INVX1_HVT U441 ( .A(n1193), .Y(n1208) );
  INVX1_HVT U442 ( .A(n1140), .Y(n1141) );
  INVX1_HVT U443 ( .A(n1159), .Y(n1170) );
  INVX1_HVT U444 ( .A(n1248), .Y(n1235) );
  NAND2X0_HVT U445 ( .A1(n1210), .A2(n1127), .Y(n1198) );
  INVX1_HVT U446 ( .A(n629), .Y(n630) );
  INVX1_HVT U447 ( .A(n644), .Y(n663) );
  INVX1_HVT U448 ( .A(n905), .Y(n906) );
  INVX1_HVT U449 ( .A(n820), .Y(n821) );
  INVX1_HVT U450 ( .A(n815), .Y(n819) );
  INVX1_HVT U451 ( .A(n882), .Y(n1126) );
  INVX1_HVT U452 ( .A(n896), .Y(n897) );
  INVX1_HVT U453 ( .A(n964), .Y(n1240) );
  INVX1_HVT U454 ( .A(n736), .Y(n755) );
  INVX1_HVT U455 ( .A(n985), .Y(n986) );
  INVX1_HVT U456 ( .A(n1020), .Y(n1081) );
  INVX1_HVT U457 ( .A(n1362), .Y(n1092) );
  INVX1_HVT U458 ( .A(n566), .Y(n519) );
  INVX1_HVT U459 ( .A(n613), .Y(n618) );
  INVX1_HVT U460 ( .A(n601), .Y(n602) );
  NAND2X0_HVT U461 ( .A1(col[0]), .A2(n125), .Y(n1194) );
  INVX1_HVT U462 ( .A(n1614), .Y(n1615) );
  INVX1_HVT U463 ( .A(n1608), .Y(n1627) );
  INVX1_HVT U464 ( .A(n870), .Y(n868) );
  INVX1_HVT U465 ( .A(n910), .Y(n920) );
  INVX1_HVT U466 ( .A(n1672), .Y(n1671) );
  INVX1_HVT U467 ( .A(n1677), .Y(n1678) );
  INVX1_HVT U468 ( .A(n1673), .Y(n1674) );
  INVX1_HVT U469 ( .A(n1688), .Y(n1690) );
  INVX1_HVT U470 ( .A(n953), .Y(n951) );
  INVX1_HVT U471 ( .A(n992), .Y(n1005) );
  INVX1_HVT U472 ( .A(n688), .Y(n734) );
  INVX1_HVT U473 ( .A(n704), .Y(n952) );
  INVX1_HVT U474 ( .A(n702), .Y(n710) );
  INVX1_HVT U475 ( .A(n721), .Y(n750) );
  INVX1_HVT U476 ( .A(n719), .Y(n706) );
  INVX1_HVT U477 ( .A(n697), .Y(n712) );
  INVX1_HVT U478 ( .A(n797), .Y(n1041) );
  INVX1_HVT U479 ( .A(n524), .Y(n532) );
  INVX1_HVT U480 ( .A(n520), .Y(n521) );
  INVX1_HVT U481 ( .A(n825), .Y(n837) );
  NAND3X0_HVT U482 ( .A1(n163), .A2(n167), .A3(n268), .Y(n1249) );
  INVX1_HVT U483 ( .A(n784), .Y(n782) );
  INVX1_HVT U484 ( .A(n1380), .Y(n1382) );
  INVX1_HVT U485 ( .A(n1397), .Y(n1391) );
  INVX1_HVT U486 ( .A(n1395), .Y(n1398) );
  INVX1_HVT U487 ( .A(n1413), .Y(n1416) );
  NOR4X1_HVT U488 ( .A1(sram_raddr_weight[11]), .A2(sram_raddr_weight[9]), 
        .A3(sram_raddr_weight[10]), .A4(n1394), .Y(n1387) );
  INVX1_HVT U489 ( .A(n1568), .Y(n1567) );
  INVX1_HVT U490 ( .A(n1563), .Y(n1570) );
  AND2X1_HVT U491 ( .A1(mode[0]), .A2(n463), .Y(n1329) );
  INVX1_HVT U492 ( .A(n1489), .Y(n1448) );
  NAND2X0_HVT U493 ( .A1(n105), .A2(n1540), .Y(net28264) );
  NOR4X1_HVT U494 ( .A1(n1527), .A2(n233), .A3(channel_cnt[3]), .A4(
        channel_cnt[2]), .Y(n492) );
  INVX1_HVT U495 ( .A(n1535), .Y(n1534) );
  INVX1_HVT U496 ( .A(n486), .Y(n1542) );
  OAI221X1_HVT U497 ( .A1(n703), .A2(n1304), .A3(n703), .A4(n962), .A5(n127), 
        .Y(n185) );
  AOI222X1_HVT U498 ( .A1(sram_raddr_b6[6]), .A2(n1066), .A3(sram_raddr_b6[6]), 
        .A4(n1263), .A5(n1066), .A6(n1065), .Y(n216) );
  OAI222X1_HVT U499 ( .A1(sram_raddr_weight[5]), .A2(n1416), .A3(
        sram_raddr_weight[5]), .A4(n1443), .A5(n372), .A6(n1415), .Y(n217) );
  OAI221X1_HVT U500 ( .A1(n881), .A2(n910), .A3(n881), .A4(n880), .A5(n127), 
        .Y(n218) );
  OAI221X1_HVT U501 ( .A1(sram_raddr_b5[5]), .A2(n1240), .A3(n193), .A4(n964), 
        .A5(n148), .Y(n219) );
  AOI22X1_HVT U502 ( .A1(n1239), .A2(n1019), .A3(n1018), .A4(n1096), .Y(n220)
         );
  AOI22X1_HVT U503 ( .A1(n1759), .A2(n1787), .A3(sram_raddr_a4[2]), .A4(n1920), 
        .Y(n221) );
  AOI22X1_HVT U504 ( .A1(sram_raddr_b8[1]), .A2(n1226), .A3(n1214), .A4(n1310), 
        .Y(n222) );
  AOI22X1_HVT U505 ( .A1(n95), .A2(n164), .A3(n1837), .A4(n1871), .Y(n223) );
  AOI22X1_HVT U506 ( .A1(n95), .A2(sram_raddr_a3[1]), .A3(n1836), .A4(n1871), 
        .Y(n224) );
  AOI22X1_HVT U507 ( .A1(sram_raddr_a7[2]), .A2(n1920), .A3(n1882), .A4(n1918), 
        .Y(n225) );
  AOI22X1_HVT U508 ( .A1(sram_raddr_b7[1]), .A2(n1194), .A3(n1102), .A4(n1198), 
        .Y(n226) );
  AOI22X1_HVT U509 ( .A1(sram_raddr_a2[9]), .A2(n1711), .A3(n1710), .A4(n1709), 
        .Y(n240) );
  AOI22X1_HVT U510 ( .A1(sram_raddr_a1[9]), .A2(n1652), .A3(n1651), .A4(n1650), 
        .Y(n241) );
  AOI22X1_HVT U511 ( .A1(sram_raddr_a0[9]), .A2(n1602), .A3(n1601), .A4(n1600), 
        .Y(n242) );
  OAI221X1_HVT U512 ( .A1(sram_raddr_a1[2]), .A2(n1604), .A3(sram_raddr_a1[2]), 
        .A4(n1640), .A5(n1607), .Y(n340) );
  OAI221X1_HVT U513 ( .A1(n963), .A2(n992), .A3(n963), .A4(n962), .A5(n128), 
        .Y(n341) );
  AOI22X1_HVT U514 ( .A1(n1716), .A2(n1751), .A3(sram_raddr_a3[2]), .A4(n108), 
        .Y(n342) );
  AOI22X1_HVT U515 ( .A1(sram_raddr_a8[2]), .A2(n1967), .A3(n1931), .A4(n1965), 
        .Y(n343) );
  AOI22X1_HVT U516 ( .A1(sram_raddr_a8[9]), .A2(n1967), .A3(n1966), .A4(n1965), 
        .Y(n344) );
  AOI22X1_HVT U517 ( .A1(sram_raddr_a7[9]), .A2(n1920), .A3(n1919), .A4(n1918), 
        .Y(n345) );
  NAND2X0_HVT U518 ( .A1(n94), .A2(n1882), .Y(n346) );
  NAND2X0_HVT U519 ( .A1(n1881), .A2(n204), .Y(n347) );
  AO221X1_HVT U520 ( .A1(n172), .A2(n1558), .A3(n172), .A4(n1557), .A5(n1566), 
        .Y(n348) );
  NAND2X0_HVT U521 ( .A1(n436), .A2(n437), .Y(n349) );
  NAND2X0_HVT U522 ( .A1(n448), .A2(n449), .Y(n350) );
  NAND2X0_HVT U523 ( .A1(n430), .A2(n431), .Y(n351) );
  NAND2X0_HVT U524 ( .A1(n1945), .A2(n1968), .Y(n387) );
  NAND3X0_HVT U525 ( .A1(n344), .A2(n386), .A3(n387), .Y(n_sram_raddr_a8[9])
         );
  NAND2X0_HVT U526 ( .A1(n95), .A2(n1932), .Y(n388) );
  NAND3X0_HVT U527 ( .A1(n343), .A2(n1930), .A3(n388), .Y(n_sram_raddr_a8[2])
         );
  NAND2X0_HVT U528 ( .A1(n95), .A2(n1921), .Y(n390) );
  NAND3X0_HVT U529 ( .A1(n345), .A2(n389), .A3(n390), .Y(n_sram_raddr_a7[9])
         );
  NAND2X0_HVT U530 ( .A1(n95), .A2(n174), .Y(n391) );
  NAND3X0_HVT U531 ( .A1(n225), .A2(n396), .A3(n391), .Y(n_sram_raddr_a7[2])
         );
  NAND2X0_HVT U532 ( .A1(sram_raddr_a6[9]), .A2(n109), .Y(n393) );
  NAND3X0_HVT U533 ( .A1(n1873), .A2(n392), .A3(n393), .Y(n_sram_raddr_a6[9])
         );
  NAND2X0_HVT U534 ( .A1(sram_raddr_a6[2]), .A2(n109), .Y(n394) );
  NAND3X0_HVT U535 ( .A1(n223), .A2(n347), .A3(n394), .Y(n_sram_raddr_a6[2])
         );
  NAND2X0_HVT U536 ( .A1(sram_raddr_a6[1]), .A2(n108), .Y(n395) );
  NAND3X0_HVT U537 ( .A1(n224), .A2(n1835), .A3(n395), .Y(n_sram_raddr_a6[1])
         );
  NAND2X0_HVT U538 ( .A1(n1881), .A2(n165), .Y(n396) );
  NAND3X0_HVT U539 ( .A1(n221), .A2(n346), .A3(n396), .Y(n_sram_raddr_a4[2])
         );
  NAND2X0_HVT U540 ( .A1(n1837), .A2(n94), .Y(n397) );
  NAND3X0_HVT U541 ( .A1(n342), .A2(n347), .A3(n397), .Y(n_sram_raddr_a3[2])
         );
  NAND2X0_HVT U542 ( .A1(n95), .A2(n1831), .Y(n399) );
  NAND3X0_HVT U543 ( .A1(n240), .A2(n398), .A3(n399), .Y(n_sram_raddr_a2[9])
         );
  NAND2X0_HVT U544 ( .A1(n1945), .A2(n1788), .Y(n401) );
  NAND3X0_HVT U545 ( .A1(n241), .A2(n400), .A3(n401), .Y(n_sram_raddr_a1[9])
         );
  NAND2X0_HVT U546 ( .A1(n1945), .A2(n1759), .Y(n402) );
  NAND3X0_HVT U547 ( .A1(n346), .A2(n340), .A3(n402), .Y(n_sram_raddr_a1[2])
         );
  NAND2X0_HVT U548 ( .A1(n1945), .A2(n1752), .Y(n404) );
  NAND3X0_HVT U549 ( .A1(n242), .A2(n403), .A3(n404), .Y(n_sram_raddr_a0[9])
         );
  NAND2X0_HVT U550 ( .A1(n1945), .A2(n1717), .Y(n406) );
  NAND3X0_HVT U551 ( .A1(n405), .A2(n348), .A3(n406), .Y(n_sram_raddr_a0[3])
         );
  NAND2X0_HVT U552 ( .A1(n1417), .A2(n127), .Y(n407) );
  NAND3X0_HVT U553 ( .A1(n217), .A2(n1431), .A3(n407), .Y(net19857) );
  NAND2X0_HVT U554 ( .A1(n256), .A2(n1258), .Y(n409) );
  NAND3X0_HVT U555 ( .A1(n103), .A2(n408), .A3(n409), .Y(n1259) );
  NAND2X0_HVT U556 ( .A1(n1239), .A2(n1215), .Y(n410) );
  NAND3X0_HVT U557 ( .A1(n222), .A2(n1213), .A3(n410), .Y(n1216) );
  NAND2X0_HVT U558 ( .A1(n255), .A2(n1156), .Y(n412) );
  NAND3X0_HVT U559 ( .A1(n103), .A2(n411), .A3(n412), .Y(n1157) );
  NAND2X0_HVT U560 ( .A1(n1239), .A2(n1103), .Y(n413) );
  NAND3X0_HVT U561 ( .A1(n226), .A2(n1101), .A3(n413), .Y(n1104) );
  NAND2X0_HVT U562 ( .A1(n1067), .A2(n1096), .Y(n414) );
  NAND3X0_HVT U563 ( .A1(n216), .A2(n351), .A3(n414), .Y(n1070) );
  NAND2X0_HVT U564 ( .A1(n254), .A2(n1061), .Y(n416) );
  NAND3X0_HVT U565 ( .A1(n103), .A2(n415), .A3(n416), .Y(n1062) );
  NAND2X0_HVT U566 ( .A1(sram_raddr_b6[1]), .A2(n1020), .Y(n417) );
  NAND3X0_HVT U567 ( .A1(n220), .A2(n1016), .A3(n417), .Y(n1021) );
  NAND2X0_HVT U568 ( .A1(sram_raddr_b5[5]), .A2(n160), .Y(n418) );
  NAND3X0_HVT U569 ( .A1(n219), .A2(n341), .A3(n418), .Y(n_sram_raddr_b5[5])
         );
  NAND2X0_HVT U570 ( .A1(n263), .A2(n883), .Y(n420) );
  NAND3X0_HVT U571 ( .A1(n103), .A2(n419), .A3(n420), .Y(n891) );
  NAND2X0_HVT U572 ( .A1(sram_raddr_b4[5]), .A2(n161), .Y(n421) );
  NAND3X0_HVT U573 ( .A1(n349), .A2(n218), .A3(n421), .Y(n_sram_raddr_b4[5])
         );
  NAND2X0_HVT U574 ( .A1(n267), .A2(n716), .Y(n422) );
  NAND3X0_HVT U575 ( .A1(n103), .A2(n727), .A3(n422), .Y(n717) );
  NAND2X0_HVT U576 ( .A1(sram_raddr_b2[5]), .A2(n162), .Y(n423) );
  NAND3X0_HVT U577 ( .A1(n350), .A2(n185), .A3(n423), .Y(n_sram_raddr_b2[5])
         );
  NAND2X0_HVT U578 ( .A1(n266), .A2(n623), .Y(n424) );
  NAND3X0_HVT U579 ( .A1(n103), .A2(n636), .A3(n424), .Y(n624) );
  NAND2X0_HVT U580 ( .A1(n262), .A2(n537), .Y(n425) );
  NAND3X0_HVT U581 ( .A1(n103), .A2(n549), .A3(n425), .Y(n538) );
  AND2X1_HVT U582 ( .A1(n456), .A2(n457), .Y(n1827) );
  AND2X1_HVT U583 ( .A1(n1521), .A2(n1522), .Y(n426) );
  OR2X1_HVT U584 ( .A1(delay1_sram_waddr_d[1]), .A2(delay1_sram_waddr_d[0]), 
        .Y(n427) );
  AND2X1_HVT U585 ( .A1(n426), .A2(n427), .Y(net19985) );
  AND2X1_HVT U586 ( .A1(n1506), .A2(n1507), .Y(n428) );
  OR2X1_HVT U587 ( .A1(delay1_sram_waddr_c[1]), .A2(delay1_sram_waddr_c[0]), 
        .Y(n429) );
  AND2X1_HVT U588 ( .A1(n428), .A2(n429), .Y(net19969) );
  AND2X1_HVT U589 ( .A1(n1073), .A2(n1304), .Y(n430) );
  OR2X1_HVT U590 ( .A1(n1064), .A2(sram_raddr_b3[6]), .Y(n431) );
  AND2X1_HVT U591 ( .A1(n1003), .A2(n1006), .Y(n432) );
  OR2X1_HVT U592 ( .A1(n1004), .A2(n1005), .Y(n433) );
  AND2X1_HVT U593 ( .A1(n432), .A2(n433), .Y(n1007) );
  AND2X1_HVT U594 ( .A1(n934), .A2(n936), .Y(n434) );
  OR2X1_HVT U595 ( .A1(n935), .A2(n1005), .Y(n435) );
  AND2X1_HVT U596 ( .A1(n434), .A2(n435), .Y(n937) );
  AND2X1_HVT U597 ( .A1(n883), .A2(n149), .Y(n436) );
  OR2X1_HVT U598 ( .A1(n1126), .A2(sram_raddr_b4[5]), .Y(n437) );
  AND2X1_HVT U599 ( .A1(n852), .A2(n854), .Y(n438) );
  OR2X1_HVT U600 ( .A1(n853), .A2(n920), .Y(n439) );
  AND2X1_HVT U601 ( .A1(n438), .A2(n439), .Y(n855) );
  AND2X1_HVT U602 ( .A1(n835), .A2(n838), .Y(n440) );
  OR2X1_HVT U603 ( .A1(n836), .A2(n837), .Y(n441) );
  AND2X1_HVT U604 ( .A1(n440), .A2(n441), .Y(n841) );
  AND2X1_HVT U605 ( .A1(n793), .A2(n795), .Y(n442) );
  OR2X1_HVT U606 ( .A1(n794), .A2(n837), .Y(n443) );
  AND2X1_HVT U607 ( .A1(n442), .A2(n443), .Y(n796) );
  AND2X1_HVT U608 ( .A1(n792), .A2(n1058), .Y(n444) );
  OR2X1_HVT U609 ( .A1(n1052), .A2(n804), .Y(n445) );
  AND2X1_HVT U610 ( .A1(n444), .A2(n445), .Y(n795) );
  AND2X1_HVT U611 ( .A1(n971), .A2(n714), .Y(n446) );
  OR2X1_HVT U612 ( .A1(n969), .A2(n154), .Y(n447) );
  AND2X1_HVT U613 ( .A1(n446), .A2(n447), .Y(n715) );
  AND2X1_HVT U614 ( .A1(n716), .A2(n102), .Y(n448) );
  OR2X1_HVT U615 ( .A1(n952), .A2(sram_raddr_b2[5]), .Y(n449) );
  AND2X1_HVT U616 ( .A1(n887), .A2(n620), .Y(n450) );
  OR2X1_HVT U617 ( .A1(n888), .A2(n154), .Y(n451) );
  AND2X1_HVT U618 ( .A1(n450), .A2(n451), .Y(n621) );
  AND2X1_HVT U619 ( .A1(n861), .A2(n594), .Y(n452) );
  OR2X1_HVT U620 ( .A1(n858), .A2(n155), .Y(n453) );
  AND2X1_HVT U621 ( .A1(n452), .A2(n453), .Y(n595) );
  AND2X1_HVT U622 ( .A1(n801), .A2(n534), .Y(n454) );
  OR2X1_HVT U623 ( .A1(n802), .A2(n154), .Y(n455) );
  AND2X1_HVT U624 ( .A1(n454), .A2(n455), .Y(n535) );
  AND2X1_HVT U625 ( .A1(n276), .A2(n1547), .Y(n456) );
  AND2X1_HVT U626 ( .A1(n456), .A2(n457), .Y(n458) );
  AO21X1_HVT U627 ( .A1(n463), .A2(n461), .A3(n158), .Y(N2888) );
  NAND3X0_HVT U628 ( .A1(col[3]), .A2(n1542), .A3(n167), .Y(n1653) );
  AND2X1_HVT U629 ( .A1(n1979), .A2(n1653), .Y(n1970) );
  AND3X1_HVT U630 ( .A1(n1970), .A2(n1135), .A3(n1136), .Y(
        n_addr_col_sel_cnt[0]) );
  AND3X1_HVT U631 ( .A1(n1135), .A2(n1970), .A3(addr_col_sel_cnt[0]), .Y(
        n_addr_col_sel_cnt[1]) );
  AND4X1_HVT U632 ( .A1(n1137), .A2(n1545), .A3(n1979), .A4(n276), .Y(n1544)
         );
  AO21X1_HVT U633 ( .A1(addr_row_sel_cnt[0]), .A2(n1970), .A3(n1544), .Y(
        n_addr_row_sel_cnt_0_) );
  AO22X1_HVT U634 ( .A1(col[1]), .A2(n1324), .A3(n1329), .A4(data_sel_col[1]), 
        .Y(n1972) );
  AO22X1_HVT U635 ( .A1(row[0]), .A2(n1324), .A3(n1329), .A4(data_sel_row[0]), 
        .Y(n1975) );
  AO22X1_HVT U636 ( .A1(row[1]), .A2(n1324), .A3(n1329), .A4(data_sel_row[1]), 
        .Y(n1976) );
  OAI221X1_HVT U637 ( .A1(n1972), .A2(n1975), .A3(n1972), .A4(n1976), .A5(
        n1979), .Y(n1730) );
  NAND4X0_HVT U638 ( .A1(n1109), .A2(n166), .A3(n177), .A4(n232), .Y(n493) );
  NAND3X0_HVT U639 ( .A1(n98), .A2(n493), .A3(n1363), .Y(n1973) );
  AO22X1_HVT U640 ( .A1(col[0]), .A2(n1324), .A3(n1329), .A4(data_sel_col[0]), 
        .Y(n464) );
  NAND2X0_HVT U641 ( .A1(n117), .A2(n493), .Y(n1977) );
  NAND3X0_HVT U642 ( .A1(n1979), .A2(n464), .A3(n1972), .Y(n1723) );
  NAND4X0_HVT U643 ( .A1(weight_cnt[4]), .A2(n176), .A3(n213), .A4(n324), .Y(
        n469) );
  NAND4X0_HVT U644 ( .A1(state[1]), .A2(n1108), .A3(n1109), .A4(n166), .Y(
        n1334) );
  AO22X1_HVT U645 ( .A1(row[1]), .A2(col[3]), .A3(n237), .A4(n163), .Y(n489)
         );
  NAND2X0_HVT U646 ( .A1(row[1]), .A2(col[3]), .Y(n476) );
  OA221X1_HVT U647 ( .A1(n183), .A2(n167), .A3(n183), .A4(n489), .A5(n476), 
        .Y(n467) );
  AO21X1_HVT U648 ( .A1(n183), .A2(n167), .A3(n486), .Y(n474) );
  NAND3X0_HVT U649 ( .A1(row[0]), .A2(n167), .A3(n489), .Y(n465) );
  NAND2X0_HVT U650 ( .A1(row[0]), .A2(col[2]), .Y(n473) );
  OA22X1_HVT U651 ( .A1(n474), .A2(n465), .A3(n476), .A4(n473), .Y(n466) );
  AO221X1_HVT U652 ( .A1(n179), .A2(n467), .A3(n179), .A4(n466), .A5(n234), 
        .Y(n477) );
  OR2X1_HVT U653 ( .A1(n1363), .A2(n477), .Y(n1342) );
  NAND4X0_HVT U654 ( .A1(weight_cnt[1]), .A2(weight_cnt[5]), .A3(n367), .A4(
        n227), .Y(n468) );
  NOR3X0_HVT U655 ( .A1(conv_done), .A2(n469), .A3(n468), .Y(n_conv_done) );
  AND2X1_HVT U656 ( .A1(n1979), .A2(n178), .Y(n1654) );
  NAND2X0_HVT U657 ( .A1(n1284), .A2(n194), .Y(n1017) );
  NOR2X0_HVT U658 ( .A1(n493), .A2(channel_cnt[0]), .Y(net19998) );
  OR2X1_HVT U659 ( .A1(channel_cnt[2]), .A2(channel_cnt[3]), .Y(n470) );
  AO22X1_HVT U660 ( .A1(n1654), .A2(n472), .A3(net19998), .A4(n471), .Y(
        n_load_data_enable) );
  AO21X1_HVT U661 ( .A1(n474), .A2(n473), .A3(n489), .Y(n475) );
  NAND4X0_HVT U662 ( .A1(n476), .A2(n475), .A3(n179), .A4(n234), .Y(n1364) );
  NAND2X0_HVT U663 ( .A1(n1979), .A2(n477), .Y(n1341) );
  OA22X1_HVT U664 ( .A1(n488), .A2(n1434), .A3(n1545), .A4(n1341), .Y(n1360)
         );
  NAND2X0_HVT U665 ( .A1(n1435), .A2(n1360), .Y(n479) );
  AO22X1_HVT U666 ( .A1(n1545), .A2(n478), .A3(n488), .A4(n1422), .Y(n481) );
  AO22X1_HVT U667 ( .A1(row[0]), .A2(n479), .A3(n183), .A4(n481), .Y(n_row[0])
         );
  AND2X1_HVT U668 ( .A1(row[0]), .A2(n481), .Y(n480) );
  AO21X1_HVT U669 ( .A1(n1546), .A2(n481), .A3(n479), .Y(n482) );
  OA21X1_HVT U670 ( .A1(row[1]), .A2(n480), .A3(n482), .Y(n_row[1]) );
  OA222X1_HVT U671 ( .A1(row[2]), .A2(row[1]), .A3(row[2]), .A4(n480), .A5(
        n179), .A6(n482), .Y(n_row[2]) );
  AND3X1_HVT U672 ( .A1(row[0]), .A2(row[1]), .A3(n481), .Y(n483) );
  AO22X1_HVT U673 ( .A1(row[2]), .A2(n483), .A3(row[3]), .A4(n482), .Y(
        n_row[3]) );
  AND3X1_HVT U674 ( .A1(n1447), .A2(write_col[0]), .A3(n484), .Y(
        n_sram_bytemask_b[0]) );
  AND3X1_HVT U675 ( .A1(n1447), .A2(n352), .A3(n484), .Y(n_sram_bytemask_b[1])
         );
  AND3X1_HVT U676 ( .A1(write_col[0]), .A2(n1447), .A3(n485), .Y(
        n_sram_bytemask_b[2]) );
  AND3X1_HVT U677 ( .A1(n1447), .A2(n485), .A3(n352), .Y(n_sram_bytemask_b[3])
         );
  AND4X1_HVT U678 ( .A1(write_col[0]), .A2(n1324), .A3(n1492), .A4(n484), .Y(
        n_sram_bytemask_c[0]) );
  AND4X1_HVT U679 ( .A1(n1324), .A2(n352), .A3(n1492), .A4(n484), .Y(
        n_sram_bytemask_c[1]) );
  AND4X1_HVT U680 ( .A1(write_col[0]), .A2(n1324), .A3(n485), .A4(n1492), .Y(
        n_sram_bytemask_c[2]) );
  AND4X1_HVT U681 ( .A1(n1324), .A2(n485), .A3(n352), .A4(n1492), .Y(
        n_sram_bytemask_c[3]) );
  AND4X1_HVT U682 ( .A1(mem_sel), .A2(write_col[0]), .A3(n1324), .A4(n484), 
        .Y(n_sram_bytemask_d[0]) );
  AND4X1_HVT U683 ( .A1(mem_sel), .A2(n1324), .A3(n352), .A4(n484), .Y(
        n_sram_bytemask_d[1]) );
  AND4X1_HVT U684 ( .A1(write_col[0]), .A2(mem_sel), .A3(n1324), .A4(n485), 
        .Y(n_sram_bytemask_d[2]) );
  AND4X1_HVT U685 ( .A1(mem_sel), .A2(n1324), .A3(n485), .A4(n352), .Y(
        n_sram_bytemask_d[3]) );
  AO22X1_HVT U686 ( .A1(col[1]), .A2(n194), .A3(n268), .A4(col[0]), .Y(n1362)
         );
  AND2X1_HVT U687 ( .A1(n163), .A2(n167), .Y(n598) );
  NAND2X0_HVT U688 ( .A1(n1092), .A2(n123), .Y(n1020) );
  NAND2X0_HVT U689 ( .A1(n152), .A2(n1017), .Y(n566) );
  OA22X1_HVT U690 ( .A1(n1210), .A2(sram_raddr_b6[0]), .A3(n155), .A4(
        sram_raddr_b3[0]), .Y(n1014) );
  OAI221X1_HVT U691 ( .A1(n184), .A2(n1081), .A3(sram_raddr_b0[0]), .A4(n519), 
        .A5(n1014), .Y(n494) );
  NAND2X0_HVT U692 ( .A1(n1528), .A2(n492), .Y(n1336) );
  AO22X1_HVT U693 ( .A1(n127), .A2(n494), .A3(sram_raddr_b0[0]), .A4(n1270), 
        .Y(n_sram_raddr_b0[0]) );
  NAND2X0_HVT U694 ( .A1(sram_raddr_b3[0]), .A2(sram_raddr_b3[1]), .Y(n506) );
  NAND2X0_HVT U695 ( .A1(n215), .A2(n335), .Y(n1042) );
  NAND2X0_HVT U696 ( .A1(n506), .A2(n1042), .Y(n1019) );
  OA22X1_HVT U697 ( .A1(n1081), .A2(n239), .A3(n110), .A4(n1019), .Y(n496) );
  NAND2X0_HVT U698 ( .A1(sram_raddr_b6[1]), .A2(sram_raddr_b6[0]), .Y(n503) );
  OA21X1_HVT U699 ( .A1(sram_raddr_b6[1]), .A2(sram_raddr_b6[0]), .A3(n503), 
        .Y(n1018) );
  NAND2X0_HVT U700 ( .A1(n121), .A2(n1018), .Y(n764) );
  NAND2X0_HVT U701 ( .A1(sram_raddr_b0[0]), .A2(sram_raddr_b0[1]), .Y(n762) );
  NAND2X0_HVT U702 ( .A1(n184), .A2(n239), .Y(n784) );
  NAND3X0_HVT U703 ( .A1(n566), .A2(n762), .A3(n784), .Y(n495) );
  NAND3X0_HVT U704 ( .A1(n496), .A2(n764), .A3(n495), .Y(n497) );
  AO22X1_HVT U705 ( .A1(n119), .A2(n497), .A3(sram_raddr_b0[1]), .A4(n1270), 
        .Y(n_sram_raddr_b0[1]) );
  NAND3X0_HVT U706 ( .A1(n163), .A2(n167), .A3(n1362), .Y(n1052) );
  NAND2X0_HVT U707 ( .A1(n259), .A2(n762), .Y(n511) );
  OA22X1_HVT U708 ( .A1(sram_raddr_b0[2]), .A2(n1052), .A3(n519), .A4(n511), 
        .Y(n505) );
  AO22X1_HVT U709 ( .A1(sram_raddr_b6[2]), .A2(n498), .A3(n169), .A4(n503), 
        .Y(n1025) );
  NAND2X0_HVT U710 ( .A1(n120), .A2(n1025), .Y(n767) );
  AO221X1_HVT U711 ( .A1(n125), .A2(n519), .A3(n125), .A4(n762), .A5(n259), 
        .Y(n499) );
  NAND3X0_HVT U712 ( .A1(n505), .A2(n767), .A3(n499), .Y(n501) );
  AO22X1_HVT U713 ( .A1(sram_raddr_b3[2]), .A2(n500), .A3(n249), .A4(n506), 
        .Y(n768) );
  OA221X1_HVT U714 ( .A1(n501), .A2(n1239), .A3(n501), .A4(n768), .A5(n128), 
        .Y(n502) );
  AO221X1_HVT U715 ( .A1(sram_raddr_b0[2]), .A2(n161), .A3(n259), .A4(n149), 
        .A5(n502), .Y(n_sram_raddr_b0[2]) );
  NAND2X0_HVT U717 ( .A1(n169), .A2(n503), .Y(n504) );
  NAND2X0_HVT U718 ( .A1(sram_raddr_b6[3]), .A2(n504), .Y(n508) );
  OA21X1_HVT U719 ( .A1(sram_raddr_b6[3]), .A2(n504), .A3(n508), .Y(n1029) );
  NAND2X0_HVT U720 ( .A1(n122), .A2(n1029), .Y(n775) );
  NAND4X0_HVT U721 ( .A1(col[1]), .A2(n163), .A3(n167), .A4(n194), .Y(n1209)
         );
  NAND2X0_HVT U722 ( .A1(n152), .A2(n1209), .Y(n721) );
  NAND2X0_HVT U723 ( .A1(n750), .A2(n1249), .Y(n688) );
  NAND2X0_HVT U724 ( .A1(n249), .A2(n506), .Y(n507) );
  NAND2X0_HVT U725 ( .A1(sram_raddr_b3[3]), .A2(n507), .Y(n509) );
  OA21X1_HVT U726 ( .A1(sram_raddr_b3[3]), .A2(n507), .A3(n509), .Y(n771) );
  NAND2X0_HVT U728 ( .A1(sram_raddr_b0[3]), .A2(sram_raddr_b0[2]), .Y(n781) );
  NAND2X0_HVT U729 ( .A1(n298), .A2(n508), .Y(n524) );
  OA21X1_HVT U730 ( .A1(n508), .A2(n298), .A3(n524), .Y(n1044) );
  NAND2X0_HVT U731 ( .A1(n253), .A2(n509), .Y(n520) );
  OA21X1_HVT U732 ( .A1(n509), .A2(n253), .A3(n520), .Y(n780) );
  OA22X1_HVT U733 ( .A1(n1044), .A2(n1210), .A3(n780), .A4(n154), .Y(n787) );
  NAND2X0_HVT U734 ( .A1(n251), .A2(n781), .Y(n510) );
  NAND3X0_HVT U735 ( .A1(sram_raddr_b0[4]), .A2(sram_raddr_b0[3]), .A3(
        sram_raddr_b0[2]), .Y(n536) );
  NAND2X0_HVT U736 ( .A1(n510), .A2(n536), .Y(n515) );
  NAND2X0_HVT U737 ( .A1(sram_raddr_b0[3]), .A2(n511), .Y(n512) );
  AND2X1_HVT U738 ( .A1(n251), .A2(n512), .Y(n529) );
  AO22X1_HVT U739 ( .A1(n1077), .A2(n515), .A3(n529), .A4(n566), .Y(n523) );
  AO221X1_HVT U740 ( .A1(n126), .A2(n519), .A3(n126), .A4(n512), .A5(n251), 
        .Y(n513) );
  NAND3X0_HVT U741 ( .A1(n787), .A2(n514), .A3(n513), .Y(n517) );
  AO222X1_HVT U742 ( .A1(n517), .A2(n129), .A3(n148), .A4(n516), .A5(
        sram_raddr_b0[4]), .A6(n162), .Y(n_sram_raddr_b0[4]) );
  AND3X1_HVT U743 ( .A1(n124), .A2(n251), .A3(n781), .Y(n518) );
  OA22X1_HVT U744 ( .A1(n519), .A2(n529), .A3(n1081), .A4(n518), .Y(n522) );
  NAND2X0_HVT U745 ( .A1(n521), .A2(n190), .Y(n531) );
  OA21X1_HVT U746 ( .A1(n521), .A2(n190), .A3(n531), .Y(n794) );
  OA22X1_HVT U747 ( .A1(n522), .A2(n196), .A3(n794), .A4(n155), .Y(n525) );
  NAND3X0_HVT U748 ( .A1(n196), .A2(n536), .A3(n523), .Y(n530) );
  AO22X1_HVT U749 ( .A1(sram_raddr_b6[5]), .A2(n524), .A3(n254), .A4(n532), 
        .Y(n1054) );
  NAND2X0_HVT U750 ( .A1(n120), .A2(n1054), .Y(n793) );
  NAND3X0_HVT U751 ( .A1(n525), .A2(n530), .A3(n793), .Y(n526) );
  AO22X1_HVT U752 ( .A1(n1537), .A2(n526), .A3(sram_raddr_b0[5]), .A4(n162), 
        .Y(n528) );
  NAND4X0_HVT U753 ( .A1(sram_raddr_b0[5]), .A2(sram_raddr_b0[4]), .A3(
        sram_raddr_b0[3]), .A4(sram_raddr_b0[2]), .Y(n537) );
  NAND2X0_HVT U754 ( .A1(n196), .A2(n536), .Y(n527) );
  OA222X1_HVT U755 ( .A1(n528), .A2(n149), .A3(n528), .A4(n537), .A5(n528), 
        .A6(n527), .Y(n_sram_raddr_b0[5]) );
  NAND3X0_HVT U756 ( .A1(n196), .A2(n251), .A3(n781), .Y(n540) );
  NAND2X0_HVT U757 ( .A1(n529), .A2(n196), .Y(n541) );
  AOI22X1_HVT U758 ( .A1(n1077), .A2(n540), .A3(n566), .A4(n541), .Y(n542) );
  OA222X1_HVT U759 ( .A1(n262), .A2(n123), .A3(n262), .A4(n530), .A5(
        sram_raddr_b0[6]), .A6(n542), .Y(n534) );
  NAND2X0_HVT U760 ( .A1(sram_raddr_b3[6]), .A2(n531), .Y(n543) );
  OAI21X1_HVT U761 ( .A1(sram_raddr_b3[6]), .A2(n531), .A3(n543), .Y(n802) );
  NAND2X0_HVT U762 ( .A1(n532), .A2(n254), .Y(n533) );
  NAND2X0_HVT U763 ( .A1(sram_raddr_b6[6]), .A2(n533), .Y(n544) );
  OA21X1_HVT U764 ( .A1(sram_raddr_b6[6]), .A2(n533), .A3(n544), .Y(n1067) );
  NAND2X0_HVT U765 ( .A1(n120), .A2(n1067), .Y(n801) );
  OA22X1_HVT U766 ( .A1(n535), .A2(n98), .A3(n262), .A4(n1296), .Y(n539) );
  NAND3X0_HVT U767 ( .A1(sram_raddr_b0[6]), .A2(sram_raddr_b0[5]), .A3(n783), 
        .Y(n549) );
  NAND2X0_HVT U768 ( .A1(n539), .A2(n538), .Y(n_sram_raddr_b0[6]) );
  NAND2X0_HVT U769 ( .A1(sram_raddr_b0[6]), .A2(n540), .Y(n563) );
  NAND2X0_HVT U770 ( .A1(sram_raddr_b0[6]), .A2(n541), .Y(n562) );
  AO22X1_HVT U771 ( .A1(n1077), .A2(n563), .A3(n566), .A4(n562), .Y(n553) );
  NAND2X0_HVT U772 ( .A1(n553), .A2(n211), .Y(n548) );
  OA21X1_HVT U773 ( .A1(n542), .A2(n262), .A3(n125), .Y(n554) );
  NAND2X0_HVT U774 ( .A1(n243), .A2(n543), .Y(n571) );
  OA21X1_HVT U775 ( .A1(n543), .A2(n243), .A3(n571), .Y(n810) );
  OA22X1_HVT U776 ( .A1(n554), .A2(n211), .A3(n810), .A4(n155), .Y(n547) );
  AND2X1_HVT U777 ( .A1(n197), .A2(n544), .Y(n567) );
  AO21X1_HVT U778 ( .A1(n546), .A2(sram_raddr_b6[7]), .A3(n567), .Y(n1076) );
  NAND2X0_HVT U779 ( .A1(n121), .A2(n1076), .Y(n812) );
  NAND3X0_HVT U780 ( .A1(n548), .A2(n547), .A3(n812), .Y(n552) );
  NAND2X0_HVT U781 ( .A1(n211), .A2(n549), .Y(n551) );
  NAND2X0_HVT U782 ( .A1(sram_raddr_b0[7]), .A2(n558), .Y(n557) );
  AND2X1_HVT U783 ( .A1(n103), .A2(n557), .Y(n550) );
  AO222X1_HVT U784 ( .A1(n552), .A2(n129), .A3(n551), .A4(n550), .A5(n162), 
        .A6(sram_raddr_b0[7]), .Y(n_sram_raddr_b0[7]) );
  HADDX1_HVT U785 ( .A0(sram_raddr_b6[8]), .B0(n567), .SO(n1086) );
  NAND2X0_HVT U786 ( .A1(n121), .A2(n1086), .Y(n824) );
  NAND3X0_HVT U787 ( .A1(n314), .A2(n211), .A3(n553), .Y(n570) );
  AO221X1_HVT U788 ( .A1(n554), .A2(n734), .A3(n554), .A4(n211), .A5(n314), 
        .Y(n556) );
  HADDX1_HVT U789 ( .A0(n186), .B0(n571), .SO(n826) );
  NAND2X0_HVT U790 ( .A1(n1304), .A2(n826), .Y(n555) );
  NAND4X0_HVT U791 ( .A1(n824), .A2(n570), .A3(n556), .A4(n555), .Y(n560) );
  AO221X1_HVT U792 ( .A1(n102), .A2(n314), .A3(n148), .A4(n557), .A5(n162), 
        .Y(n561) );
  NAND3X0_HVT U793 ( .A1(sram_raddr_b0[7]), .A2(n149), .A3(n558), .Y(n574) );
  NAND2X0_HVT U794 ( .A1(n314), .A2(n574), .Y(n559) );
  AO22X1_HVT U795 ( .A1(n1536), .A2(n560), .A3(n561), .A4(n559), .Y(
        n_sram_raddr_b0[8]) );
  NAND2X0_HVT U796 ( .A1(sram_raddr_b0[9]), .A2(n561), .Y(n577) );
  NAND3X0_HVT U797 ( .A1(n314), .A2(n211), .A3(n562), .Y(n565) );
  NAND4X0_HVT U798 ( .A1(n124), .A2(n314), .A3(n211), .A4(n563), .Y(n564) );
  AOI22X1_HVT U799 ( .A1(n566), .A2(n565), .A3(n1020), .A4(n564), .Y(n569) );
  NAND2X0_HVT U800 ( .A1(n567), .A2(n258), .Y(n568) );
  HADDX1_HVT U801 ( .A0(n568), .B0(n292), .SO(n1097) );
  NAND2X0_HVT U802 ( .A1(n120), .A2(n1097), .Y(n835) );
  OA221X1_HVT U803 ( .A1(sram_raddr_b0[9]), .A2(n570), .A3(n325), .A4(n569), 
        .A5(n835), .Y(n573) );
  OR2X1_HVT U804 ( .A1(n571), .A2(sram_raddr_b3[8]), .Y(n572) );
  HADDX1_HVT U805 ( .A0(sram_raddr_b3[9]), .B0(n572), .SO(n836) );
  AO221X1_HVT U806 ( .A1(n573), .A2(n110), .A3(n573), .A4(n836), .A5(n98), .Y(
        n576) );
  OR3X1_HVT U807 ( .A1(sram_raddr_b0[9]), .A2(n574), .A3(n314), .Y(n575) );
  NAND3X0_HVT U808 ( .A1(n577), .A2(n576), .A3(n575), .Y(n_sram_raddr_b0[9])
         );
  NAND2X0_HVT U809 ( .A1(col[0]), .A2(n1284), .Y(n1127) );
  NAND2X0_HVT U810 ( .A1(n152), .A2(n1127), .Y(n628) );
  AO22X1_HVT U811 ( .A1(n122), .A2(n308), .A3(n1304), .A4(n206), .Y(n578) );
  AO221X1_HVT U812 ( .A1(sram_raddr_b1[0]), .A2(n1194), .A3(n175), .A4(n628), 
        .A5(n578), .Y(n579) );
  AO22X1_HVT U813 ( .A1(n130), .A2(n579), .A3(sram_raddr_b1[0]), .A4(n1270), 
        .Y(n_sram_raddr_b1[0]) );
  NAND2X0_HVT U814 ( .A1(sram_raddr_b4[0]), .A2(sram_raddr_b4[1]), .Y(n583) );
  NAND2X0_HVT U815 ( .A1(n206), .A2(n332), .Y(n1125) );
  NAND2X0_HVT U816 ( .A1(n583), .A2(n1125), .Y(n1103) );
  OA22X1_HVT U817 ( .A1(n846), .A2(n331), .A3(n155), .A4(n1103), .Y(n581) );
  NAND2X0_HVT U818 ( .A1(sram_raddr_b7[1]), .A2(sram_raddr_b7[0]), .Y(n592) );
  OA21X1_HVT U819 ( .A1(sram_raddr_b7[1]), .A2(sram_raddr_b7[0]), .A3(n592), 
        .Y(n1102) );
  NAND2X0_HVT U820 ( .A1(n122), .A2(n1102), .Y(n849) );
  NAND2X0_HVT U821 ( .A1(sram_raddr_b1[0]), .A2(sram_raddr_b1[1]), .Y(n847) );
  NAND2X0_HVT U822 ( .A1(n175), .A2(n331), .Y(n870) );
  NAND3X0_HVT U823 ( .A1(n628), .A2(n847), .A3(n870), .Y(n580) );
  NAND3X0_HVT U824 ( .A1(n581), .A2(n849), .A3(n580), .Y(n582) );
  AO22X1_HVT U825 ( .A1(n119), .A2(n582), .A3(sram_raddr_b1[1]), .A4(n1270), 
        .Y(n_sram_raddr_b1[1]) );
  NAND3X0_HVT U826 ( .A1(sram_raddr_b1[0]), .A2(sram_raddr_b1[1]), .A3(n628), 
        .Y(n585) );
  NAND2X0_HVT U827 ( .A1(n188), .A2(n585), .Y(n589) );
  NAND2X0_HVT U828 ( .A1(n246), .A2(n583), .Y(n591) );
  OA21X1_HVT U829 ( .A1(n583), .A2(n246), .A3(n591), .Y(n853) );
  OA22X1_HVT U830 ( .A1(n734), .A2(n589), .A3(n853), .A4(n155), .Y(n584) );
  OA221X1_HVT U831 ( .A1(n188), .A2(n126), .A3(n188), .A4(n585), .A5(n584), 
        .Y(n587) );
  AO22X1_HVT U832 ( .A1(sram_raddr_b7[2]), .A2(n586), .A3(n257), .A4(n592), 
        .Y(n1110) );
  NAND2X0_HVT U833 ( .A1(n121), .A2(n1110), .Y(n852) );
  AOI21X1_HVT U834 ( .A1(n587), .A2(n852), .A3(n98), .Y(n588) );
  AO221X1_HVT U835 ( .A1(sram_raddr_b1[2]), .A2(n161), .A3(n188), .A4(n150), 
        .A5(n588), .Y(n_sram_raddr_b1[2]) );
  HADDX1_HVT U836 ( .A0(n248), .B0(n589), .SO(n590) );
  OA22X1_HVT U837 ( .A1(n123), .A2(n248), .A3(n734), .A4(n590), .Y(n594) );
  NAND2X0_HVT U838 ( .A1(sram_raddr_b4[3]), .A2(n591), .Y(n603) );
  OAI21X1_HVT U839 ( .A1(sram_raddr_b4[3]), .A2(n591), .A3(n603), .Y(n858) );
  NAND2X0_HVT U840 ( .A1(n257), .A2(n592), .Y(n593) );
  NAND2X0_HVT U841 ( .A1(sram_raddr_b7[3]), .A2(n593), .Y(n601) );
  OA21X1_HVT U842 ( .A1(sram_raddr_b7[3]), .A2(n593), .A3(n601), .Y(n1113) );
  NAND2X0_HVT U843 ( .A1(n120), .A2(n1113), .Y(n861) );
  OA22X1_HVT U844 ( .A1(n595), .A2(n98), .A3(n99), .A4(n248), .Y(n597) );
  AO221X1_HVT U845 ( .A1(sram_raddr_b1[3]), .A2(sram_raddr_b1[2]), .A3(n248), 
        .A4(n188), .A5(n1339), .Y(n596) );
  NAND2X0_HVT U846 ( .A1(n597), .A2(n596), .Y(n_sram_raddr_b1[3]) );
  NAND2X0_HVT U847 ( .A1(n598), .A2(n194), .Y(n1142) );
  NAND3X0_HVT U848 ( .A1(sram_raddr_b1[4]), .A2(sram_raddr_b1[3]), .A3(
        sram_raddr_b1[2]), .Y(n622) );
  NAND2X0_HVT U849 ( .A1(sram_raddr_b1[3]), .A2(sram_raddr_b1[2]), .Y(n867) );
  NAND2X0_HVT U850 ( .A1(n250), .A2(n867), .Y(n599) );
  NAND2X0_HVT U851 ( .A1(n622), .A2(n599), .Y(n608) );
  AO21X1_HVT U852 ( .A1(n188), .A2(n847), .A3(n248), .Y(n600) );
  AND2X1_HVT U853 ( .A1(n250), .A2(n600), .Y(n614) );
  AO22X1_HVT U854 ( .A1(n1183), .A2(n608), .A3(n614), .A4(n628), .Y(n612) );
  AO221X1_HVT U855 ( .A1(n125), .A2(n658), .A3(n126), .A4(n600), .A5(n250), 
        .Y(n606) );
  OR2X1_HVT U856 ( .A1(sram_raddr_b7[4]), .A2(n602), .Y(n613) );
  AO21X1_HVT U857 ( .A1(n602), .A2(sram_raddr_b7[4]), .A3(n618), .Y(n1128) );
  NAND2X0_HVT U858 ( .A1(n121), .A2(n1128), .Y(n872) );
  AND2X1_HVT U859 ( .A1(n284), .A2(n603), .Y(n611) );
  AO21X1_HVT U860 ( .A1(n604), .A2(sram_raddr_b4[4]), .A3(n611), .Y(n873) );
  NAND2X0_HVT U861 ( .A1(n1304), .A2(n873), .Y(n605) );
  NAND4X0_HVT U862 ( .A1(n607), .A2(n606), .A3(n872), .A4(n605), .Y(n610) );
  AO222X1_HVT U863 ( .A1(n610), .A2(n127), .A3(n150), .A4(n609), .A5(n161), 
        .A6(sram_raddr_b1[4]), .Y(n_sram_raddr_b1[4]) );
  NAND2X0_HVT U864 ( .A1(n611), .A2(n199), .Y(n631) );
  OA21X1_HVT U865 ( .A1(n611), .A2(n199), .A3(n631), .Y(n879) );
  NAND3X0_HVT U866 ( .A1(n195), .A2(n622), .A3(n612), .Y(n616) );
  AO22X1_HVT U867 ( .A1(sram_raddr_b7[5]), .A2(n613), .A3(n255), .A4(n618), 
        .Y(n1147) );
  NAND2X0_HVT U868 ( .A1(n122), .A2(n1147), .Y(n878) );
  NAND4X0_HVT U869 ( .A1(sram_raddr_b1[5]), .A2(sram_raddr_b1[4]), .A3(
        sram_raddr_b1[3]), .A4(sram_raddr_b1[2]), .Y(n623) );
  NAND2X0_HVT U870 ( .A1(n614), .A2(n195), .Y(n627) );
  NAND3X0_HVT U871 ( .A1(n195), .A2(n250), .A3(n867), .Y(n626) );
  AO21X1_HVT U872 ( .A1(n1183), .A2(n626), .A3(n628), .Y(n629) );
  NAND2X0_HVT U873 ( .A1(n627), .A2(n629), .Y(n615) );
  OA222X1_HVT U874 ( .A1(n266), .A2(n125), .A3(n266), .A4(n616), .A5(
        sram_raddr_b1[6]), .A6(n615), .Y(n620) );
  AO22X1_HVT U875 ( .A1(sram_raddr_b4[6]), .A2(n631), .A3(n263), .A4(n617), 
        .Y(n888) );
  NAND2X0_HVT U876 ( .A1(n618), .A2(n255), .Y(n619) );
  NAND2X0_HVT U877 ( .A1(sram_raddr_b7[6]), .A2(n619), .Y(n633) );
  OA21X1_HVT U878 ( .A1(sram_raddr_b7[6]), .A2(n619), .A3(n633), .Y(n1161) );
  NAND2X0_HVT U879 ( .A1(n122), .A2(n1161), .Y(n887) );
  OA22X1_HVT U880 ( .A1(n621), .A2(n117), .A3(n99), .A4(n266), .Y(n625) );
  NAND3X0_HVT U881 ( .A1(sram_raddr_b1[6]), .A2(sram_raddr_b1[5]), .A3(n869), 
        .Y(n636) );
  NAND2X0_HVT U882 ( .A1(n625), .A2(n624), .Y(n_sram_raddr_b1[6]) );
  NAND2X0_HVT U883 ( .A1(sram_raddr_b1[6]), .A2(n626), .Y(n654) );
  NAND2X0_HVT U884 ( .A1(sram_raddr_b1[6]), .A2(n627), .Y(n656) );
  AO22X1_HVT U885 ( .A1(n1183), .A2(n654), .A3(n628), .A4(n656), .Y(n641) );
  NAND2X0_HVT U886 ( .A1(n641), .A2(n244), .Y(n635) );
  OA21X1_HVT U887 ( .A1(n630), .A2(n656), .A3(n123), .Y(n643) );
  NAND2X0_HVT U888 ( .A1(sram_raddr_b4[6]), .A2(n631), .Y(n632) );
  NAND2X0_HVT U889 ( .A1(n269), .A2(n632), .Y(n644) );
  OA21X1_HVT U890 ( .A1(n632), .A2(n269), .A3(n644), .Y(n895) );
  OA22X1_HVT U891 ( .A1(n643), .A2(n244), .A3(n895), .A4(n155), .Y(n634) );
  NAND2X0_HVT U892 ( .A1(n198), .A2(n633), .Y(n642) );
  NAND2X0_HVT U893 ( .A1(n122), .A2(n1177), .Y(n899) );
  NAND3X0_HVT U894 ( .A1(n635), .A2(n634), .A3(n899), .Y(n640) );
  NAND2X0_HVT U895 ( .A1(n244), .A2(n636), .Y(n639) );
  NAND2X0_HVT U896 ( .A1(sram_raddr_b1[7]), .A2(n648), .Y(n637) );
  NAND2X0_HVT U897 ( .A1(n150), .A2(n637), .Y(n647) );
  AO222X1_HVT U898 ( .A1(n640), .A2(n128), .A3(n639), .A4(n638), .A5(
        sram_raddr_b1[7]), .A6(n160), .Y(n_sram_raddr_b1[7]) );
  NAND3X0_HVT U899 ( .A1(n244), .A2(n191), .A3(n641), .Y(n662) );
  AO22X1_HVT U900 ( .A1(sram_raddr_b7[8]), .A2(n642), .A3(n280), .A4(n659), 
        .Y(n1190) );
  NAND2X0_HVT U901 ( .A1(n121), .A2(n1190), .Y(n908) );
  AO221X1_HVT U902 ( .A1(n643), .A2(n734), .A3(n643), .A4(n244), .A5(n191), 
        .Y(n646) );
  AO22X1_HVT U903 ( .A1(sram_raddr_b4[8]), .A2(n644), .A3(n265), .A4(n663), 
        .Y(n909) );
  NAND2X0_HVT U904 ( .A1(n1239), .A2(n909), .Y(n645) );
  NAND4X0_HVT U905 ( .A1(n662), .A2(n908), .A3(n646), .A4(n645), .Y(n651) );
  NAND3X0_HVT U906 ( .A1(n148), .A2(sram_raddr_b1[7]), .A3(n648), .Y(n653) );
  NAND2X0_HVT U907 ( .A1(n191), .A2(n653), .Y(n649) );
  AO22X1_HVT U908 ( .A1(n119), .A2(n651), .A3(n650), .A4(n649), .Y(
        n_sram_raddr_b1[8]) );
  AO222X1_HVT U909 ( .A1(n286), .A2(n191), .A3(n286), .A4(n653), .A5(
        sram_raddr_b1[9]), .A6(n652), .Y(n667) );
  AND2X1_HVT U910 ( .A1(n244), .A2(n191), .Y(n657) );
  OA221X1_HVT U911 ( .A1(col[0]), .A2(n657), .A3(col[0]), .A4(n654), .A5(n124), 
        .Y(n655) );
  OA221X1_HVT U912 ( .A1(n658), .A2(n657), .A3(n658), .A4(n656), .A5(n655), 
        .Y(n661) );
  NAND2X0_HVT U913 ( .A1(n659), .A2(n280), .Y(n660) );
  HADDX1_HVT U914 ( .A0(n281), .B0(n660), .SO(n1199) );
  NAND2X0_HVT U915 ( .A1(n122), .A2(n1199), .Y(n922) );
  OA221X1_HVT U916 ( .A1(sram_raddr_b1[9]), .A2(n662), .A3(n286), .A4(n661), 
        .A5(n922), .Y(n665) );
  NAND2X0_HVT U917 ( .A1(n663), .A2(n265), .Y(n664) );
  HADDX1_HVT U918 ( .A0(sram_raddr_b4[9]), .B0(n664), .SO(n919) );
  AO221X1_HVT U919 ( .A1(n665), .A2(n155), .A3(n665), .A4(n919), .A5(n117), 
        .Y(n666) );
  NAND2X0_HVT U920 ( .A1(n667), .A2(n666), .Y(n_sram_raddr_b1[9]) );
  NAND2X0_HVT U921 ( .A1(col[1]), .A2(n124), .Y(n1226) );
  AO22X1_HVT U922 ( .A1(n121), .A2(n309), .A3(n1239), .A4(n207), .Y(n668) );
  AO221X1_HVT U923 ( .A1(sram_raddr_b2[0]), .A2(n1226), .A3(n168), .A4(n721), 
        .A5(n668), .Y(n669) );
  AO22X1_HVT U924 ( .A1(n119), .A2(n669), .A3(sram_raddr_b2[0]), .A4(n1270), 
        .Y(n_sram_raddr_b2[0]) );
  NAND2X0_HVT U925 ( .A1(sram_raddr_b5[0]), .A2(sram_raddr_b5[1]), .Y(n673) );
  NAND2X0_HVT U926 ( .A1(n207), .A2(n333), .Y(n1241) );
  NAND2X0_HVT U927 ( .A1(n673), .A2(n1241), .Y(n1215) );
  OA22X1_HVT U928 ( .A1(n1288), .A2(n238), .A3(n154), .A4(n1215), .Y(n671) );
  NAND2X0_HVT U929 ( .A1(sram_raddr_b8[1]), .A2(sram_raddr_b8[0]), .Y(n681) );
  OA21X1_HVT U930 ( .A1(sram_raddr_b8[1]), .A2(sram_raddr_b8[0]), .A3(n681), 
        .Y(n1214) );
  NAND2X0_HVT U931 ( .A1(n121), .A2(n1214), .Y(n931) );
  NAND2X0_HVT U932 ( .A1(sram_raddr_b2[0]), .A2(sram_raddr_b2[1]), .Y(n930) );
  NAND2X0_HVT U933 ( .A1(n168), .A2(n238), .Y(n953) );
  NAND3X0_HVT U934 ( .A1(n721), .A2(n930), .A3(n953), .Y(n670) );
  NAND3X0_HVT U935 ( .A1(n671), .A2(n931), .A3(n670), .Y(n672) );
  AO22X1_HVT U936 ( .A1(n129), .A2(n672), .A3(sram_raddr_b2[1]), .A4(n1270), 
        .Y(n_sram_raddr_b2[1]) );
  NAND3X0_HVT U937 ( .A1(sram_raddr_b2[0]), .A2(sram_raddr_b2[1]), .A3(n721), 
        .Y(n675) );
  NAND2X0_HVT U938 ( .A1(n264), .A2(n675), .Y(n679) );
  NAND2X0_HVT U939 ( .A1(n247), .A2(n673), .Y(n683) );
  OA21X1_HVT U940 ( .A1(n673), .A2(n247), .A3(n683), .Y(n935) );
  OA22X1_HVT U941 ( .A1(n734), .A2(n679), .A3(n935), .A4(n155), .Y(n674) );
  OA221X1_HVT U942 ( .A1(n264), .A2(n126), .A3(n264), .A4(n675), .A5(n674), 
        .Y(n677) );
  AO22X1_HVT U943 ( .A1(sram_raddr_b8[2]), .A2(n676), .A3(n170), .A4(n681), 
        .Y(n1220) );
  NAND2X0_HVT U944 ( .A1(n122), .A2(n1220), .Y(n934) );
  AOI21X1_HVT U945 ( .A1(n677), .A2(n934), .A3(n117), .Y(n678) );
  AO221X1_HVT U946 ( .A1(sram_raddr_b2[2]), .A2(n162), .A3(n264), .A4(n150), 
        .A5(n678), .Y(n_sram_raddr_b2[2]) );
  HADDX1_HVT U947 ( .A0(sram_raddr_b2[3]), .B0(n679), .SO(n680) );
  AO22X1_HVT U948 ( .A1(sram_raddr_b2[3]), .A2(n1263), .A3(n680), .A4(n688), 
        .Y(n687) );
  NAND2X0_HVT U949 ( .A1(n170), .A2(n681), .Y(n682) );
  NAND2X0_HVT U950 ( .A1(sram_raddr_b8[3]), .A2(n682), .Y(n690) );
  OA21X1_HVT U951 ( .A1(sram_raddr_b8[3]), .A2(n682), .A3(n690), .Y(n1223) );
  NAND2X0_HVT U952 ( .A1(sram_raddr_b5[3]), .A2(n683), .Y(n689) );
  OA21X1_HVT U953 ( .A1(sram_raddr_b5[3]), .A2(n683), .A3(n689), .Y(n939) );
  AO22X1_HVT U954 ( .A1(n120), .A2(n1223), .A3(n1304), .A4(n939), .Y(n686) );
  NAND2X0_HVT U955 ( .A1(sram_raddr_b2[3]), .A2(sram_raddr_b2[2]), .Y(n950) );
  OA21X1_HVT U956 ( .A1(sram_raddr_b2[3]), .A2(sram_raddr_b2[2]), .A3(n950), 
        .Y(n684) );
  AO22X1_HVT U957 ( .A1(n162), .A2(sram_raddr_b2[3]), .A3(n150), .A4(n684), 
        .Y(n685) );
  AO221X1_HVT U958 ( .A1(n130), .A2(n687), .A3(n128), .A4(n686), .A5(n685), 
        .Y(n_sram_raddr_b2[3]) );
  NAND3X0_HVT U959 ( .A1(sram_raddr_b2[3]), .A2(sram_raddr_b2[0]), .A3(
        sram_raddr_b2[1]), .Y(n705) );
  OA221X1_HVT U960 ( .A1(n1284), .A2(n950), .A3(n1284), .A4(n705), .A5(n688), 
        .Y(n696) );
  NAND3X0_HVT U961 ( .A1(sram_raddr_b2[4]), .A2(sram_raddr_b2[3]), .A3(
        sram_raddr_b2[2]), .Y(n704) );
  NAND2X0_HVT U962 ( .A1(n297), .A2(n950), .Y(n698) );
  NAND2X0_HVT U963 ( .A1(n704), .A2(n698), .Y(n693) );
  NAND2X0_HVT U964 ( .A1(n696), .A2(n693), .Y(n692) );
  NAND2X0_HVT U965 ( .A1(n252), .A2(n689), .Y(n702) );
  OA21X1_HVT U966 ( .A1(n689), .A2(n252), .A3(n702), .Y(n949) );
  OA221X1_HVT U967 ( .A1(n750), .A2(n950), .A3(n750), .A4(n705), .A5(n124), 
        .Y(n700) );
  OA22X1_HVT U968 ( .A1(n949), .A2(n155), .A3(n700), .A4(n297), .Y(n691) );
  NAND2X0_HVT U969 ( .A1(n208), .A2(n690), .Y(n697) );
  OAI21X1_HVT U970 ( .A1(n690), .A2(n208), .A3(n697), .Y(n1236) );
  NAND2X0_HVT U971 ( .A1(n122), .A2(n1236), .Y(n954) );
  NAND3X0_HVT U972 ( .A1(n692), .A2(n691), .A3(n954), .Y(n695) );
  AO222X1_HVT U973 ( .A1(n695), .A2(n127), .A3(n149), .A4(n694), .A5(n161), 
        .A6(sram_raddr_b2[4]), .Y(n_sram_raddr_b2[4]) );
  NAND3X0_HVT U974 ( .A1(n203), .A2(n297), .A3(n950), .Y(n719) );
  NAND2X0_HVT U975 ( .A1(n706), .A2(n696), .Y(n709) );
  AO22X1_HVT U976 ( .A1(sram_raddr_b8[5]), .A2(n697), .A3(n256), .A4(n712), 
        .Y(n1251) );
  NAND2X0_HVT U977 ( .A1(n122), .A2(n1251), .Y(n960) );
  AO221X1_HVT U978 ( .A1(n700), .A2(n734), .A3(n700), .A4(n699), .A5(n203), 
        .Y(n701) );
  NAND3X0_HVT U979 ( .A1(n709), .A2(n960), .A3(n701), .Y(n703) );
  AO22X1_HVT U980 ( .A1(sram_raddr_b5[5]), .A2(n702), .A3(n193), .A4(n710), 
        .Y(n962) );
  NAND4X0_HVT U981 ( .A1(sram_raddr_b2[5]), .A2(sram_raddr_b2[4]), .A3(
        sram_raddr_b2[3]), .A4(sram_raddr_b2[2]), .Y(n716) );
  NAND2X0_HVT U982 ( .A1(n706), .A2(n705), .Y(n720) );
  OA21X1_HVT U983 ( .A1(n706), .A2(n1249), .A3(n750), .Y(n722) );
  NAND2X0_HVT U984 ( .A1(n720), .A2(n707), .Y(n708) );
  OA222X1_HVT U985 ( .A1(n267), .A2(n125), .A3(n267), .A4(n709), .A5(
        sram_raddr_b2[6]), .A6(n708), .Y(n714) );
  NAND2X0_HVT U986 ( .A1(n710), .A2(n193), .Y(n711) );
  NAND2X0_HVT U987 ( .A1(sram_raddr_b5[6]), .A2(n711), .Y(n723) );
  OAI21X1_HVT U988 ( .A1(sram_raddr_b5[6]), .A2(n711), .A3(n723), .Y(n969) );
  NAND2X0_HVT U989 ( .A1(n712), .A2(n256), .Y(n713) );
  NAND2X0_HVT U990 ( .A1(sram_raddr_b8[6]), .A2(n713), .Y(n724) );
  OA21X1_HVT U991 ( .A1(sram_raddr_b8[6]), .A2(n713), .A3(n724), .Y(n1261) );
  NAND2X0_HVT U992 ( .A1(n122), .A2(n1261), .Y(n971) );
  OA22X1_HVT U993 ( .A1(n715), .A2(n98), .A3(n99), .A4(n267), .Y(n718) );
  NAND3X0_HVT U994 ( .A1(sram_raddr_b2[6]), .A2(sram_raddr_b2[5]), .A3(n952), 
        .Y(n727) );
  NAND2X0_HVT U995 ( .A1(n718), .A2(n717), .Y(n_sram_raddr_b2[6]) );
  NAND2X0_HVT U996 ( .A1(sram_raddr_b2[6]), .A2(n719), .Y(n746) );
  NAND2X0_HVT U997 ( .A1(sram_raddr_b2[6]), .A2(n720), .Y(n748) );
  AO22X1_HVT U998 ( .A1(n1284), .A2(n746), .A3(n721), .A4(n748), .Y(n732) );
  NAND2X0_HVT U999 ( .A1(n732), .A2(n245), .Y(n726) );
  OA21X1_HVT U1000 ( .A1(n722), .A2(n748), .A3(n123), .Y(n735) );
  NAND2X0_HVT U1001 ( .A1(n303), .A2(n723), .Y(n736) );
  OA21X1_HVT U1002 ( .A1(n723), .A2(n303), .A3(n736), .Y(n981) );
  OA22X1_HVT U1003 ( .A1(n735), .A2(n245), .A3(n981), .A4(n154), .Y(n725) );
  NAND2X0_HVT U1004 ( .A1(n189), .A2(n724), .Y(n733) );
  NAND2X0_HVT U1005 ( .A1(n122), .A2(n1280), .Y(n979) );
  NAND3X0_HVT U1006 ( .A1(n726), .A2(n725), .A3(n979), .Y(n731) );
  NAND2X0_HVT U1007 ( .A1(n245), .A2(n727), .Y(n730) );
  NAND2X0_HVT U1008 ( .A1(sram_raddr_b2[7]), .A2(n740), .Y(n728) );
  NAND2X0_HVT U1009 ( .A1(n148), .A2(n728), .Y(n739) );
  AO222X1_HVT U1010 ( .A1(n731), .A2(n130), .A3(n730), .A4(n729), .A5(
        sram_raddr_b2[7]), .A6(n161), .Y(n_sram_raddr_b2[7]) );
  NAND3X0_HVT U1011 ( .A1(n245), .A2(n192), .A3(n732), .Y(n754) );
  AO22X1_HVT U1012 ( .A1(sram_raddr_b8[8]), .A2(n733), .A3(n260), .A4(n751), 
        .Y(n1293) );
  NAND2X0_HVT U1013 ( .A1(n120), .A2(n1293), .Y(n989) );
  AO221X1_HVT U1014 ( .A1(n735), .A2(n734), .A3(n735), .A4(n245), .A5(n192), 
        .Y(n738) );
  AO22X1_HVT U1015 ( .A1(sram_raddr_b5[8]), .A2(n736), .A3(n187), .A4(n755), 
        .Y(n991) );
  NAND2X0_HVT U1016 ( .A1(n1239), .A2(n991), .Y(n737) );
  NAND4X0_HVT U1017 ( .A1(n754), .A2(n989), .A3(n738), .A4(n737), .Y(n743) );
  NAND3X0_HVT U1018 ( .A1(n102), .A2(sram_raddr_b2[7]), .A3(n740), .Y(n745) );
  NAND2X0_HVT U1019 ( .A1(n192), .A2(n745), .Y(n741) );
  AO22X1_HVT U1020 ( .A1(n1537), .A2(n743), .A3(n742), .A4(n741), .Y(
        n_sram_raddr_b2[8]) );
  AO222X1_HVT U1021 ( .A1(n287), .A2(n192), .A3(n287), .A4(n745), .A5(
        sram_raddr_b2[9]), .A6(n744), .Y(n759) );
  AND2X1_HVT U1022 ( .A1(n245), .A2(n192), .Y(n749) );
  OA221X1_HVT U1023 ( .A1(n1249), .A2(n749), .A3(n1249), .A4(n746), .A5(n124), 
        .Y(n747) );
  OA221X1_HVT U1024 ( .A1(n750), .A2(n749), .A3(n750), .A4(n748), .A5(n747), 
        .Y(n753) );
  NAND2X0_HVT U1025 ( .A1(n751), .A2(n260), .Y(n752) );
  HADDX1_HVT U1026 ( .A0(n288), .B0(n752), .SO(n1311) );
  NAND2X0_HVT U1027 ( .A1(n121), .A2(n1311), .Y(n1003) );
  OA221X1_HVT U1028 ( .A1(sram_raddr_b2[9]), .A2(n754), .A3(n287), .A4(n753), 
        .A5(n1003), .Y(n757) );
  NAND2X0_HVT U1029 ( .A1(n755), .A2(n187), .Y(n756) );
  HADDX1_HVT U1030 ( .A0(sram_raddr_b5[9]), .B0(n756), .SO(n1004) );
  AO221X1_HVT U1031 ( .A1(n757), .A2(n154), .A3(n757), .A4(n1004), .A5(n118), 
        .Y(n758) );
  NAND2X0_HVT U1032 ( .A1(n759), .A2(n758), .Y(n_sram_raddr_b2[9]) );
  NAND2X0_HVT U1033 ( .A1(n1017), .A2(n155), .Y(n825) );
  AO22X1_HVT U1034 ( .A1(n122), .A2(n322), .A3(n998), .A4(n184), .Y(n760) );
  AO221X1_HVT U1035 ( .A1(sram_raddr_b3[0]), .A2(n1020), .A3(n215), .A4(n825), 
        .A5(n760), .Y(n761) );
  AO22X1_HVT U1036 ( .A1(n119), .A2(n761), .A3(sram_raddr_b3[0]), .A4(n1270), 
        .Y(n_sram_raddr_b3[0]) );
  OA22X1_HVT U1037 ( .A1(n1081), .A2(n335), .A3(n837), .A4(n1019), .Y(n765) );
  NAND2X0_HVT U1038 ( .A1(n762), .A2(n784), .Y(n763) );
  NAND2X0_HVT U1039 ( .A1(n998), .A2(n763), .Y(n1016) );
  NAND3X0_HVT U1040 ( .A1(n765), .A2(n764), .A3(n1016), .Y(n766) );
  AO22X1_HVT U1041 ( .A1(n1537), .A2(n766), .A3(sram_raddr_b3[1]), .A4(n1270), 
        .Y(n_sram_raddr_b3[1]) );
  NAND2X0_HVT U1042 ( .A1(n1077), .A2(n249), .Y(n770) );
  AO221X1_HVT U1043 ( .A1(sram_raddr_b0[2]), .A2(n784), .A3(n259), .A4(n782), 
        .A5(n153), .Y(n1023) );
  NAND2X0_HVT U1044 ( .A1(n102), .A2(n249), .Y(n769) );
  NAND2X0_HVT U1045 ( .A1(n99), .A2(n769), .Y(n779) );
  NAND2X0_HVT U1046 ( .A1(n123), .A2(n770), .Y(n772) );
  AOI22X1_HVT U1047 ( .A1(sram_raddr_b3[3]), .A2(n772), .A3(n771), .A4(n825), 
        .Y(n776) );
  OA222X1_HVT U1048 ( .A1(sram_raddr_b0[3]), .A2(sram_raddr_b0[2]), .A3(
        sram_raddr_b0[3]), .A4(n784), .A5(n782), .A6(n781), .Y(n773) );
  NAND2X0_HVT U1049 ( .A1(n998), .A2(n773), .Y(n1033) );
  NAND3X0_HVT U1050 ( .A1(n1077), .A2(sram_raddr_b3[2]), .A3(n307), .Y(n774)
         );
  NAND4X0_HVT U1051 ( .A1(n776), .A2(n775), .A3(n1033), .A4(n774), .Y(n778) );
  AND2X1_HVT U1052 ( .A1(sram_raddr_b3[2]), .A2(n307), .Y(n777) );
  AO222X1_HVT U1053 ( .A1(n779), .A2(sram_raddr_b3[3]), .A3(n778), .A4(n130), 
        .A5(n777), .A6(n149), .Y(n_sram_raddr_b3[3]) );
  NAND3X0_HVT U1054 ( .A1(sram_raddr_b3[4]), .A2(sram_raddr_b3[3]), .A3(
        sram_raddr_b3[2]), .Y(n797) );
  NAND2X0_HVT U1055 ( .A1(sram_raddr_b3[3]), .A2(sram_raddr_b3[2]), .Y(n1039)
         );
  NAND2X0_HVT U1056 ( .A1(n253), .A2(n1039), .Y(n791) );
  AND2X1_HVT U1057 ( .A1(n797), .A2(n791), .Y(n788) );
  OA22X1_HVT U1058 ( .A1(n126), .A2(n253), .A3(n788), .A4(n1052), .Y(n786) );
  OR2X1_HVT U1059 ( .A1(n780), .A2(n1017), .Y(n785) );
  OA21X1_HVT U1060 ( .A1(n782), .A2(n781), .A3(n251), .Y(n790) );
  OAI221X1_HVT U1061 ( .A1(n790), .A2(n784), .A3(n790), .A4(n783), .A5(n998), 
        .Y(n1046) );
  NAND4X0_HVT U1062 ( .A1(n787), .A2(n786), .A3(n785), .A4(n1046), .Y(n789) );
  AO222X1_HVT U1063 ( .A1(n789), .A2(n129), .A3(n102), .A4(n788), .A5(
        sram_raddr_b3[4]), .A6(n161), .Y(n_sram_raddr_b3[4]) );
  NAND2X0_HVT U1064 ( .A1(n790), .A2(n196), .Y(n800) );
  AO221X1_HVT U1065 ( .A1(n800), .A2(n790), .A3(n800), .A4(n196), .A5(n152), 
        .Y(n1058) );
  NAND3X0_HVT U1066 ( .A1(n190), .A2(n253), .A3(n1039), .Y(n804) );
  OAI221X1_HVT U1067 ( .A1(n1263), .A2(n1362), .A3(n1263), .A4(n791), .A5(
        sram_raddr_b3[5]), .Y(n792) );
  OA22X1_HVT U1068 ( .A1(n796), .A2(n98), .A3(n190), .A4(n99), .Y(n799) );
  AO221X1_HVT U1069 ( .A1(sram_raddr_b3[5]), .A2(n1041), .A3(n190), .A4(n797), 
        .A5(n1339), .Y(n798) );
  NAND2X0_HVT U1070 ( .A1(n799), .A2(n798), .Y(n_sram_raddr_b3[5]) );
  NAND2X0_HVT U1071 ( .A1(sram_raddr_b0[6]), .A2(n800), .Y(n809) );
  NAND2X0_HVT U1072 ( .A1(sram_raddr_b3[6]), .A2(n804), .Y(n822) );
  AO22X1_HVT U1073 ( .A1(n1077), .A2(n822), .A3(sram_raddr_b3[6]), .A4(n1263), 
        .Y(n805) );
  OAI21X1_HVT U1074 ( .A1(n837), .A2(n802), .A3(n801), .Y(n803) );
  AO221X1_HVT U1075 ( .A1(n805), .A2(sram_raddr_b3[6]), .A3(n805), .A4(n804), 
        .A5(n803), .Y(n808) );
  NAND3X0_HVT U1076 ( .A1(sram_raddr_b3[6]), .A2(sram_raddr_b3[5]), .A3(n1041), 
        .Y(n815) );
  OA221X1_HVT U1077 ( .A1(sram_raddr_b3[6]), .A2(sram_raddr_b3[5]), .A3(
        sram_raddr_b3[6]), .A4(n1041), .A5(n815), .Y(n806) );
  AO22X1_HVT U1078 ( .A1(sram_raddr_b3[6]), .A2(n161), .A3(n103), .A4(n806), 
        .Y(n807) );
  AO221X1_HVT U1079 ( .A1(n128), .A2(n1071), .A3(n127), .A4(n808), .A5(n807), 
        .Y(n_sram_raddr_b3[6]) );
  NAND2X0_HVT U1080 ( .A1(n211), .A2(n809), .Y(n820) );
  AO221X1_HVT U1081 ( .A1(n820), .A2(n211), .A3(n820), .A4(n809), .A5(n153), 
        .Y(n1075) );
  OA21X1_HVT U1082 ( .A1(n837), .A2(n810), .A3(n1075), .Y(n814) );
  NAND3X0_HVT U1083 ( .A1(n1077), .A2(n243), .A3(n822), .Y(n813) );
  AO221X1_HVT U1084 ( .A1(n126), .A2(n1092), .A3(n126), .A4(n822), .A5(n243), 
        .Y(n811) );
  NAND4X0_HVT U1085 ( .A1(n814), .A2(n813), .A3(n812), .A4(n811), .Y(n817) );
  NAND3X0_HVT U1086 ( .A1(sram_raddr_b3[7]), .A2(n819), .A3(n99), .Y(n818) );
  OA221X1_HVT U1087 ( .A1(sram_raddr_b3[7]), .A2(n150), .A3(sram_raddr_b3[7]), 
        .A4(n819), .A5(n818), .Y(n816) );
  AO22X1_HVT U1088 ( .A1(n128), .A2(n817), .A3(n816), .A4(n1270), .Y(
        n_sram_raddr_b3[7]) );
  OA22X1_HVT U1089 ( .A1(n186), .A2(n818), .A3(n162), .A4(n150), .Y(n839) );
  AND3X1_HVT U1090 ( .A1(sram_raddr_b3[7]), .A2(n149), .A3(n819), .Y(n829) );
  NAND4X0_HVT U1091 ( .A1(n1077), .A2(n243), .A3(n186), .A4(n822), .Y(n834) );
  NAND2X0_HVT U1092 ( .A1(n821), .A2(n314), .Y(n831) );
  AO221X1_HVT U1093 ( .A1(n831), .A2(n821), .A3(n831), .A4(n314), .A5(n153), 
        .Y(n1084) );
  AND3X1_HVT U1094 ( .A1(n124), .A2(n243), .A3(n822), .Y(n830) );
  OR3X1_HVT U1095 ( .A1(n1081), .A2(n830), .A3(n186), .Y(n823) );
  NAND4X0_HVT U1096 ( .A1(n824), .A2(n834), .A3(n1084), .A4(n823), .Y(n827) );
  OA221X1_HVT U1097 ( .A1(n827), .A2(n826), .A3(n827), .A4(n825), .A5(n127), 
        .Y(n828) );
  AO221X1_HVT U1098 ( .A1(n839), .A2(sram_raddr_b3[8]), .A3(n839), .A4(n829), 
        .A5(n828), .Y(n_sram_raddr_b3[8]) );
  NAND3X0_HVT U1099 ( .A1(n279), .A2(n829), .A3(sram_raddr_b3[8]), .Y(n843) );
  AO22X1_HVT U1100 ( .A1(n1092), .A2(n124), .A3(n830), .A4(n186), .Y(n833) );
  AO221X1_HVT U1101 ( .A1(sram_raddr_b0[9]), .A2(n832), .A3(n325), .A4(n831), 
        .A5(n152), .Y(n1095) );
  OA221X1_HVT U1102 ( .A1(sram_raddr_b3[9]), .A2(n834), .A3(n279), .A4(n833), 
        .A5(n1095), .Y(n838) );
  OA22X1_HVT U1103 ( .A1(n841), .A2(n98), .A3(n279), .A4(n840), .Y(n842) );
  NAND2X0_HVT U1104 ( .A1(n843), .A2(n842), .Y(n_sram_raddr_b3[9]) );
  NAND2X0_HVT U1105 ( .A1(n155), .A2(n1127), .Y(n910) );
  AO22X1_HVT U1106 ( .A1(n120), .A2(n308), .A3(n998), .A4(n175), .Y(n844) );
  AO221X1_HVT U1107 ( .A1(sram_raddr_b4[0]), .A2(n1194), .A3(n206), .A4(n910), 
        .A5(n844), .Y(n845) );
  AO22X1_HVT U1108 ( .A1(n119), .A2(n845), .A3(sram_raddr_b4[0]), .A4(n1270), 
        .Y(n_sram_raddr_b4[0]) );
  OA22X1_HVT U1109 ( .A1(n920), .A2(n1103), .A3(n846), .A4(n332), .Y(n850) );
  NAND2X0_HVT U1110 ( .A1(n847), .A2(n870), .Y(n848) );
  NAND2X0_HVT U1111 ( .A1(n998), .A2(n848), .Y(n1101) );
  NAND3X0_HVT U1112 ( .A1(n850), .A2(n849), .A3(n1101), .Y(n851) );
  AO22X1_HVT U1113 ( .A1(n1537), .A2(n851), .A3(sram_raddr_b4[1]), .A4(n1270), 
        .Y(n_sram_raddr_b4[1]) );
  AO221X1_HVT U1114 ( .A1(sram_raddr_b1[2]), .A2(n870), .A3(n188), .A4(n868), 
        .A5(n153), .Y(n1106) );
  OA221X1_HVT U1115 ( .A1(sram_raddr_b4[2]), .A2(n1142), .A3(n246), .A4(n125), 
        .A5(n1106), .Y(n854) );
  OA22X1_HVT U1116 ( .A1(n855), .A2(n118), .A3(n1296), .A4(n246), .Y(n856) );
  NAND2X0_HVT U1117 ( .A1(n149), .A2(n246), .Y(n863) );
  NAND2X0_HVT U1118 ( .A1(n856), .A2(n863), .Y(n_sram_raddr_b4[2]) );
  OA21X1_HVT U1119 ( .A1(sram_raddr_b4[2]), .A2(n1142), .A3(n125), .Y(n857) );
  OA22X1_HVT U1120 ( .A1(n920), .A2(n858), .A3(n857), .A4(n293), .Y(n862) );
  OA222X1_HVT U1121 ( .A1(sram_raddr_b1[3]), .A2(sram_raddr_b1[2]), .A3(
        sram_raddr_b1[3]), .A4(n870), .A5(n868), .A6(n867), .Y(n859) );
  NAND2X0_HVT U1122 ( .A1(n998), .A2(n859), .Y(n1117) );
  NAND3X0_HVT U1123 ( .A1(sram_raddr_b4[2]), .A2(n1183), .A3(n293), .Y(n860)
         );
  NAND4X0_HVT U1124 ( .A1(n862), .A2(n861), .A3(n1117), .A4(n860), .Y(n866) );
  NAND2X0_HVT U1125 ( .A1(n99), .A2(n863), .Y(n865) );
  AND2X1_HVT U1126 ( .A1(sram_raddr_b4[2]), .A2(n293), .Y(n864) );
  AO222X1_HVT U1127 ( .A1(n866), .A2(n128), .A3(n865), .A4(sram_raddr_b4[3]), 
        .A5(n864), .A6(n150), .Y(n_sram_raddr_b4[3]) );
  OA21X1_HVT U1128 ( .A1(n868), .A2(n867), .A3(n250), .Y(n874) );
  OAI221X1_HVT U1129 ( .A1(n874), .A2(n870), .A3(n874), .A4(n869), .A5(n998), 
        .Y(n871) );
  NAND2X0_HVT U1130 ( .A1(n872), .A2(n871), .Y(n1133) );
  NAND3X0_HVT U1131 ( .A1(sram_raddr_b4[4]), .A2(sram_raddr_b4[3]), .A3(
        sram_raddr_b4[2]), .Y(n882) );
  NAND2X0_HVT U1132 ( .A1(sram_raddr_b4[3]), .A2(sram_raddr_b4[2]), .Y(n1123)
         );
  NAND2X0_HVT U1133 ( .A1(n284), .A2(n1123), .Y(n875) );
  NAND2X0_HVT U1134 ( .A1(n874), .A2(n195), .Y(n893) );
  AO221X1_HVT U1135 ( .A1(n893), .A2(n874), .A3(n893), .A4(n195), .A5(n153), 
        .Y(n1151) );
  AND3X1_HVT U1136 ( .A1(n199), .A2(n284), .A3(n1123), .Y(n885) );
  NAND2X0_HVT U1137 ( .A1(n1183), .A2(n885), .Y(n877) );
  OAI221X1_HVT U1138 ( .A1(n1263), .A2(n194), .A3(n1263), .A4(n875), .A5(
        sram_raddr_b4[5]), .Y(n876) );
  NAND4X0_HVT U1139 ( .A1(n878), .A2(n1151), .A3(n877), .A4(n876), .Y(n881) );
  NAND4X0_HVT U1140 ( .A1(sram_raddr_b4[5]), .A2(sram_raddr_b4[4]), .A3(
        sram_raddr_b4[3]), .A4(sram_raddr_b4[2]), .Y(n883) );
  NAND2X0_HVT U1141 ( .A1(sram_raddr_b4[6]), .A2(n161), .Y(n892) );
  AND3X1_HVT U1142 ( .A1(sram_raddr_b4[6]), .A2(sram_raddr_b4[5]), .A3(n1126), 
        .Y(n904) );
  AO221X1_HVT U1143 ( .A1(sram_raddr_b1[6]), .A2(n893), .A3(n266), .A4(n884), 
        .A5(n153), .Y(n1159) );
  OA21X1_HVT U1144 ( .A1(n885), .A2(n263), .A3(n1183), .Y(n896) );
  AO222X1_HVT U1145 ( .A1(n263), .A2(n897), .A3(n263), .A4(n885), .A5(n897), 
        .A6(n123), .Y(n886) );
  AND3X1_HVT U1146 ( .A1(n887), .A2(n1159), .A3(n886), .Y(n889) );
  AO221X1_HVT U1147 ( .A1(n889), .A2(n920), .A3(n889), .A4(n888), .A5(n118), 
        .Y(n890) );
  NAND3X0_HVT U1148 ( .A1(n892), .A2(n891), .A3(n890), .Y(n_sram_raddr_b4[6])
         );
  NAND2X0_HVT U1149 ( .A1(sram_raddr_b1[6]), .A2(n893), .Y(n894) );
  NAND2X0_HVT U1150 ( .A1(n244), .A2(n894), .Y(n905) );
  AO221X1_HVT U1151 ( .A1(n905), .A2(n894), .A3(n905), .A4(n244), .A5(n153), 
        .Y(n1174) );
  OA21X1_HVT U1152 ( .A1(n920), .A2(n895), .A3(n1174), .Y(n900) );
  NAND2X0_HVT U1153 ( .A1(n896), .A2(n269), .Y(n913) );
  NAND3X0_HVT U1154 ( .A1(sram_raddr_b4[7]), .A2(n1194), .A3(n897), .Y(n898)
         );
  NAND4X0_HVT U1155 ( .A1(n900), .A2(n913), .A3(n899), .A4(n898), .Y(n902) );
  NAND3X0_HVT U1156 ( .A1(sram_raddr_b4[7]), .A2(n904), .A3(n99), .Y(n903) );
  OA221X1_HVT U1157 ( .A1(sram_raddr_b4[7]), .A2(n102), .A3(sram_raddr_b4[7]), 
        .A4(n904), .A5(n903), .Y(n901) );
  AO22X1_HVT U1158 ( .A1(n119), .A2(n902), .A3(n901), .A4(n1270), .Y(
        n_sram_raddr_b4[7]) );
  OA22X1_HVT U1159 ( .A1(n160), .A2(n150), .A3(n903), .A4(n265), .Y(n924) );
  AND3X1_HVT U1160 ( .A1(n148), .A2(sram_raddr_b4[7]), .A3(n904), .Y(n925) );
  OR2X1_HVT U1161 ( .A1(n913), .A2(sram_raddr_b4[8]), .Y(n914) );
  NAND2X0_HVT U1162 ( .A1(n906), .A2(n191), .Y(n917) );
  AO221X1_HVT U1163 ( .A1(n917), .A2(n906), .A3(n917), .A4(n191), .A5(n153), 
        .Y(n1189) );
  NAND3X0_HVT U1164 ( .A1(sram_raddr_b4[8]), .A2(n1194), .A3(n913), .Y(n907)
         );
  NAND4X0_HVT U1165 ( .A1(n914), .A2(n908), .A3(n1189), .A4(n907), .Y(n911) );
  OA221X1_HVT U1166 ( .A1(n911), .A2(n910), .A3(n911), .A4(n909), .A5(n128), 
        .Y(n912) );
  AO221X1_HVT U1167 ( .A1(n924), .A2(sram_raddr_b4[8]), .A3(n924), .A4(n925), 
        .A5(n912), .Y(n_sram_raddr_b4[8]) );
  NAND2X0_HVT U1168 ( .A1(n1194), .A2(n913), .Y(n916) );
  NAND2X0_HVT U1169 ( .A1(sram_raddr_b4[8]), .A2(n1183), .Y(n915) );
  OA222X1_HVT U1170 ( .A1(n261), .A2(n916), .A3(n261), .A4(n915), .A5(
        sram_raddr_b4[9]), .A6(n914), .Y(n923) );
  AO221X1_HVT U1171 ( .A1(sram_raddr_b1[9]), .A2(n918), .A3(n286), .A4(n917), 
        .A5(n153), .Y(n1193) );
  OR2X1_HVT U1172 ( .A1(n920), .A2(n919), .Y(n921) );
  NAND4X0_HVT U1173 ( .A1(n923), .A2(n922), .A3(n1193), .A4(n921), .Y(n927) );
  OA222X1_HVT U1174 ( .A1(sram_raddr_b4[9]), .A2(sram_raddr_b4[8]), .A3(
        sram_raddr_b4[9]), .A4(n925), .A5(n924), .A6(n261), .Y(n926) );
  AO21X1_HVT U1175 ( .A1(n129), .A2(n927), .A3(n926), .Y(n_sram_raddr_b4[9])
         );
  NAND2X0_HVT U1176 ( .A1(n1209), .A2(n110), .Y(n992) );
  AO22X1_HVT U1177 ( .A1(n121), .A2(n309), .A3(n998), .A4(n168), .Y(n928) );
  AO221X1_HVT U1178 ( .A1(sram_raddr_b5[0]), .A2(n1226), .A3(n207), .A4(n992), 
        .A5(n928), .Y(n929) );
  AO22X1_HVT U1179 ( .A1(n127), .A2(n929), .A3(sram_raddr_b5[0]), .A4(n1270), 
        .Y(n_sram_raddr_b5[0]) );
  OA22X1_HVT U1180 ( .A1(n1005), .A2(n1215), .A3(n1288), .A4(n333), .Y(n932)
         );
  AO21X1_HVT U1181 ( .A1(n930), .A2(n953), .A3(n153), .Y(n1213) );
  NAND3X0_HVT U1182 ( .A1(n932), .A2(n931), .A3(n1213), .Y(n933) );
  AO22X1_HVT U1183 ( .A1(n1537), .A2(n933), .A3(sram_raddr_b5[1]), .A4(n1270), 
        .Y(n_sram_raddr_b5[1]) );
  AO221X1_HVT U1184 ( .A1(sram_raddr_b2[2]), .A2(n953), .A3(n264), .A4(n951), 
        .A5(n152), .Y(n1219) );
  OA221X1_HVT U1185 ( .A1(sram_raddr_b5[2]), .A2(n1249), .A3(n247), .A4(n125), 
        .A5(n1219), .Y(n936) );
  OA22X1_HVT U1186 ( .A1(n937), .A2(n98), .A3(n99), .A4(n247), .Y(n938) );
  NAND2X0_HVT U1187 ( .A1(n103), .A2(n247), .Y(n944) );
  NAND2X0_HVT U1188 ( .A1(n938), .A2(n944), .Y(n_sram_raddr_b5[2]) );
  AOI22X1_HVT U1189 ( .A1(n122), .A2(n1223), .A3(n939), .A4(n992), .Y(n943) );
  AO221X1_HVT U1190 ( .A1(n123), .A2(sram_raddr_b5[2]), .A3(n125), .A4(n1249), 
        .A5(n291), .Y(n942) );
  OA222X1_HVT U1191 ( .A1(sram_raddr_b2[3]), .A2(sram_raddr_b2[2]), .A3(
        sram_raddr_b2[3]), .A4(n953), .A5(n951), .A6(n950), .Y(n940) );
  NAND2X0_HVT U1192 ( .A1(n998), .A2(n940), .Y(n1229) );
  NAND3X0_HVT U1193 ( .A1(n1284), .A2(sram_raddr_b5[2]), .A3(n291), .Y(n941)
         );
  NAND4X0_HVT U1194 ( .A1(n943), .A2(n942), .A3(n1229), .A4(n941), .Y(n947) );
  NAND2X0_HVT U1195 ( .A1(n99), .A2(n944), .Y(n946) );
  AND2X1_HVT U1196 ( .A1(sram_raddr_b5[2]), .A2(n291), .Y(n945) );
  AO222X1_HVT U1197 ( .A1(n947), .A2(n129), .A3(n946), .A4(sram_raddr_b5[3]), 
        .A5(n945), .A6(n103), .Y(n_sram_raddr_b5[3]) );
  NAND3X0_HVT U1198 ( .A1(sram_raddr_b5[4]), .A2(sram_raddr_b5[3]), .A3(
        sram_raddr_b5[2]), .Y(n964) );
  NAND2X0_HVT U1199 ( .A1(sram_raddr_b5[3]), .A2(sram_raddr_b5[2]), .Y(n1237)
         );
  NAND2X0_HVT U1200 ( .A1(n252), .A2(n1237), .Y(n948) );
  AND2X1_HVT U1201 ( .A1(n964), .A2(n948), .Y(n956) );
  OA22X1_HVT U1202 ( .A1(n1005), .A2(n949), .A3(n956), .A4(n1249), .Y(n955) );
  OA21X1_HVT U1203 ( .A1(n951), .A2(n950), .A3(n297), .Y(n959) );
  OAI221X1_HVT U1204 ( .A1(n959), .A2(n953), .A3(n959), .A4(n952), .A5(n998), 
        .Y(n1244) );
  NAND3X0_HVT U1205 ( .A1(n955), .A2(n954), .A3(n1244), .Y(n957) );
  AO21X1_HVT U1206 ( .A1(n130), .A2(n1263), .A3(n160), .Y(n1540) );
  AO222X1_HVT U1207 ( .A1(n957), .A2(n130), .A3(n1540), .A4(sram_raddr_b5[4]), 
        .A5(n956), .A6(n148), .Y(n_sram_raddr_b5[4]) );
  OA221X1_HVT U1208 ( .A1(col[1]), .A2(n252), .A3(col[1]), .A4(n1237), .A5(
        n124), .Y(n958) );
  NAND3X0_HVT U1209 ( .A1(n193), .A2(n252), .A3(n1237), .Y(n965) );
  OA22X1_HVT U1210 ( .A1(n958), .A2(n193), .A3(n1249), .A4(n965), .Y(n961) );
  NAND2X0_HVT U1211 ( .A1(n959), .A2(n203), .Y(n976) );
  AO221X1_HVT U1212 ( .A1(n976), .A2(n959), .A3(n976), .A4(n203), .A5(n153), 
        .Y(n1255) );
  NAND3X0_HVT U1213 ( .A1(n961), .A2(n960), .A3(n1255), .Y(n963) );
  NAND2X0_HVT U1214 ( .A1(sram_raddr_b5[6]), .A2(n965), .Y(n987) );
  NAND2X0_HVT U1215 ( .A1(n1284), .A2(n987), .Y(n967) );
  AO222X1_HVT U1216 ( .A1(n967), .A2(n295), .A3(n967), .A4(n126), .A5(n295), 
        .A6(n966), .Y(n972) );
  AO221X1_HVT U1217 ( .A1(sram_raddr_b2[6]), .A2(n976), .A3(n267), .A4(n968), 
        .A5(n153), .Y(n1269) );
  OR2X1_HVT U1218 ( .A1(n1005), .A2(n969), .Y(n970) );
  NAND4X0_HVT U1219 ( .A1(n972), .A2(n971), .A3(n1269), .A4(n970), .Y(n975) );
  AND4X1_HVT U1220 ( .A1(sram_raddr_b5[5]), .A2(sram_raddr_b5[4]), .A3(
        sram_raddr_b5[3]), .A4(sram_raddr_b5[2]), .Y(n973) );
  OAI221X1_HVT U1221 ( .A1(n1339), .A2(sram_raddr_b5[6]), .A3(n1339), .A4(n973), .A5(n99), .Y(n993) );
  AO21X1_HVT U1222 ( .A1(n148), .A2(n973), .A3(sram_raddr_b5[6]), .Y(n974) );
  AO22X1_HVT U1223 ( .A1(n119), .A2(n975), .A3(n993), .A4(n974), .Y(
        n_sram_raddr_b5[6]) );
  AND4X1_HVT U1224 ( .A1(n103), .A2(sram_raddr_b5[6]), .A3(sram_raddr_b5[5]), 
        .A4(n1240), .Y(n1009) );
  NAND3X0_HVT U1225 ( .A1(n1284), .A2(n303), .A3(n987), .Y(n980) );
  NAND2X0_HVT U1226 ( .A1(sram_raddr_b2[6]), .A2(n976), .Y(n977) );
  NAND2X0_HVT U1227 ( .A1(n245), .A2(n977), .Y(n985) );
  AO221X1_HVT U1228 ( .A1(n985), .A2(n977), .A3(n985), .A4(n245), .A5(n153), 
        .Y(n1278) );
  AO221X1_HVT U1229 ( .A1(n123), .A2(col[1]), .A3(n123), .A4(n987), .A5(n303), 
        .Y(n978) );
  NAND4X0_HVT U1230 ( .A1(n980), .A2(n979), .A3(n1278), .A4(n978), .Y(n983) );
  OA221X1_HVT U1231 ( .A1(n983), .A2(n992), .A3(n983), .A4(n982), .A5(n128), 
        .Y(n984) );
  AO221X1_HVT U1232 ( .A1(sram_raddr_b5[7]), .A2(n993), .A3(n303), .A4(n1009), 
        .A5(n984), .Y(n_sram_raddr_b5[7]) );
  NAND4X0_HVT U1233 ( .A1(n1284), .A2(n303), .A3(n187), .A4(n987), .Y(n1002)
         );
  NAND2X0_HVT U1234 ( .A1(n986), .A2(n192), .Y(n999) );
  AO221X1_HVT U1235 ( .A1(n999), .A2(n986), .A3(n999), .A4(n192), .A5(n153), 
        .Y(n1291) );
  AND3X1_HVT U1236 ( .A1(n124), .A2(n303), .A3(n987), .Y(n997) );
  OR3X1_HVT U1237 ( .A1(n1288), .A2(n997), .A3(n187), .Y(n988) );
  NAND4X0_HVT U1238 ( .A1(n1002), .A2(n989), .A3(n1291), .A4(n988), .Y(n990)
         );
  AO21X1_HVT U1239 ( .A1(n992), .A2(n991), .A3(n990), .Y(n995) );
  AO221X1_HVT U1240 ( .A1(n149), .A2(n187), .A3(n102), .A4(n303), .A5(n993), 
        .Y(n996) );
  AO21X1_HVT U1241 ( .A1(sram_raddr_b5[7]), .A2(n1009), .A3(sram_raddr_b5[8]), 
        .Y(n994) );
  AO22X1_HVT U1242 ( .A1(n1537), .A2(n995), .A3(n996), .A4(n994), .Y(
        n_sram_raddr_b5[8]) );
  AO22X1_HVT U1243 ( .A1(col[1]), .A2(n124), .A3(n997), .A4(n187), .Y(n1001)
         );
  AO221X1_HVT U1244 ( .A1(sram_raddr_b2[9]), .A2(n1000), .A3(n287), .A4(n999), 
        .A5(n153), .Y(n1308) );
  OA221X1_HVT U1245 ( .A1(sram_raddr_b5[9]), .A2(n1002), .A3(n282), .A4(n1001), 
        .A5(n1308), .Y(n1006) );
  OA22X1_HVT U1246 ( .A1(n1008), .A2(n282), .A3(n1007), .A4(n118), .Y(n1011)
         );
  NAND4X0_HVT U1247 ( .A1(sram_raddr_b5[8]), .A2(sram_raddr_b5[7]), .A3(n1009), 
        .A4(n282), .Y(n1010) );
  NAND2X0_HVT U1248 ( .A1(n1011), .A2(n1010), .Y(n_sram_raddr_b5[9]) );
  AO22X1_HVT U1249 ( .A1(sram_raddr_b6[0]), .A2(n1081), .A3(n322), .A4(n1017), 
        .Y(n1013) );
  NAND2X0_HVT U1250 ( .A1(n998), .A2(n184), .Y(n1012) );
  NAND3X0_HVT U1251 ( .A1(n1014), .A2(n1013), .A3(n1012), .Y(n1015) );
  AO22X1_HVT U1252 ( .A1(n130), .A2(n1015), .A3(sram_raddr_b6[0]), .A4(n1270), 
        .Y(n_sram_raddr_b6[0]) );
  NAND2X0_HVT U1253 ( .A1(n1210), .A2(n1017), .Y(n1096) );
  AO22X1_HVT U1254 ( .A1(n119), .A2(n1021), .A3(sram_raddr_b6[1]), .A4(n1270), 
        .Y(n_sram_raddr_b6[1]) );
  AO22X1_HVT U1255 ( .A1(sram_raddr_b6[2]), .A2(n123), .A3(n169), .A4(n1052), 
        .Y(n1024) );
  AO221X1_HVT U1256 ( .A1(sram_raddr_b3[2]), .A2(n1042), .A3(n249), .A4(n1040), 
        .A5(n154), .Y(n1022) );
  NAND3X0_HVT U1257 ( .A1(n1024), .A2(n1023), .A3(n1022), .Y(n1026) );
  OA221X1_HVT U1258 ( .A1(n1026), .A2(n1096), .A3(n1026), .A4(n1025), .A5(n130), .Y(n1027) );
  AO221X1_HVT U1259 ( .A1(sram_raddr_b6[2]), .A2(n160), .A3(n169), .A4(n149), 
        .A5(n1027), .Y(n_sram_raddr_b6[2]) );
  NAND2X0_HVT U1260 ( .A1(n102), .A2(n169), .Y(n1028) );
  NAND2X0_HVT U1261 ( .A1(n99), .A2(n1028), .Y(n1037) );
  OA222X1_HVT U1262 ( .A1(sram_raddr_b3[3]), .A2(sram_raddr_b3[2]), .A3(
        sram_raddr_b3[3]), .A4(n1042), .A5(n1040), .A6(n1039), .Y(n1030) );
  AOI22X1_HVT U1263 ( .A1(n1304), .A2(n1030), .A3(n1029), .A4(n1096), .Y(n1034) );
  AO221X1_HVT U1264 ( .A1(n126), .A2(sram_raddr_b6[2]), .A3(n126), .A4(n1052), 
        .A5(n202), .Y(n1032) );
  NAND3X0_HVT U1265 ( .A1(sram_raddr_b6[2]), .A2(n1077), .A3(n202), .Y(n1031)
         );
  NAND4X0_HVT U1266 ( .A1(n1034), .A2(n1033), .A3(n1032), .A4(n1031), .Y(n1036) );
  AND2X1_HVT U1267 ( .A1(sram_raddr_b6[2]), .A2(n202), .Y(n1035) );
  AO222X1_HVT U1268 ( .A1(n1037), .A2(sram_raddr_b6[3]), .A3(n1036), .A4(n129), 
        .A5(n1035), .A6(n102), .Y(n_sram_raddr_b6[3]) );
  NAND3X0_HVT U1269 ( .A1(sram_raddr_b6[4]), .A2(sram_raddr_b6[3]), .A3(
        sram_raddr_b6[2]), .Y(n1061) );
  OA21X1_HVT U1270 ( .A1(n202), .A2(n169), .A3(n298), .Y(n1051) );
  AND2X1_HVT U1271 ( .A1(n1061), .A2(n1038), .Y(n1049) );
  OA22X1_HVT U1272 ( .A1(n126), .A2(n298), .A3(n1049), .A4(n1052), .Y(n1048)
         );
  OA21X1_HVT U1273 ( .A1(n1040), .A2(n1039), .A3(n253), .Y(n1055) );
  AOI21X1_HVT U1274 ( .A1(n1042), .A2(n1041), .A3(n1055), .Y(n1043) );
  OA22X1_HVT U1275 ( .A1(n1045), .A2(n1044), .A3(n1043), .A4(n110), .Y(n1047)
         );
  NAND3X0_HVT U1276 ( .A1(n1048), .A2(n1047), .A3(n1046), .Y(n1050) );
  AO222X1_HVT U1277 ( .A1(n1050), .A2(n129), .A3(n148), .A4(n1049), .A5(
        sram_raddr_b6[4]), .A6(n160), .Y(n_sram_raddr_b6[4]) );
  OA21X1_HVT U1278 ( .A1(n1092), .A2(n1051), .A3(n123), .Y(n1053) );
  NAND2X0_HVT U1279 ( .A1(n1051), .A2(n254), .Y(n1065) );
  OA22X1_HVT U1280 ( .A1(n1053), .A2(n254), .A3(n1052), .A4(n1065), .Y(n1059)
         );
  NAND2X0_HVT U1281 ( .A1(n1096), .A2(n1054), .Y(n1057) );
  NAND2X0_HVT U1282 ( .A1(n1055), .A2(n190), .Y(n1064) );
  AO221X1_HVT U1283 ( .A1(n1064), .A2(n1055), .A3(n1064), .A4(n190), .A5(n154), 
        .Y(n1056) );
  AND4X1_HVT U1284 ( .A1(n1059), .A2(n1058), .A3(n1057), .A4(n1056), .Y(n1060)
         );
  OA22X1_HVT U1285 ( .A1(n1060), .A2(n117), .A3(n254), .A4(n99), .Y(n1063) );
  AND4X1_HVT U1286 ( .A1(sram_raddr_b6[5]), .A2(sram_raddr_b6[4]), .A3(
        sram_raddr_b6[3]), .A4(sram_raddr_b6[2]), .Y(n1072) );
  NAND2X0_HVT U1287 ( .A1(n1063), .A2(n1062), .Y(n_sram_raddr_b6[5]) );
  NAND2X0_HVT U1288 ( .A1(sram_raddr_b3[6]), .A2(n1064), .Y(n1073) );
  NAND2X0_HVT U1289 ( .A1(sram_raddr_b6[6]), .A2(n1065), .Y(n1080) );
  NAND2X0_HVT U1290 ( .A1(n1077), .A2(n1080), .Y(n1074) );
  NAND2X0_HVT U1291 ( .A1(sram_raddr_b6[6]), .A2(n1072), .Y(n1068) );
  AO21X1_HVT U1292 ( .A1(n102), .A2(n1068), .A3(n162), .Y(n1087) );
  OA221X1_HVT U1293 ( .A1(sram_raddr_b6[6]), .A2(n103), .A3(sram_raddr_b6[6]), 
        .A4(n1072), .A5(n1087), .Y(n1069) );
  AO221X1_HVT U1294 ( .A1(n129), .A2(n1071), .A3(n130), .A4(n1070), .A5(n1069), 
        .Y(n_sram_raddr_b6[6]) );
  AND3X1_HVT U1295 ( .A1(sram_raddr_b6[6]), .A2(n103), .A3(n1072), .Y(n1090)
         );
  NAND2X0_HVT U1296 ( .A1(n243), .A2(n1073), .Y(n1078) );
  NAND4X0_HVT U1297 ( .A1(n1077), .A2(n258), .A3(n197), .A4(n1080), .Y(n1093)
         );
  NAND2X0_HVT U1298 ( .A1(n1079), .A2(n186), .Y(n1094) );
  AO221X1_HVT U1299 ( .A1(n1094), .A2(n1079), .A3(n1094), .A4(n186), .A5(n154), 
        .Y(n1083) );
  AND3X1_HVT U1300 ( .A1(n124), .A2(n197), .A3(n1080), .Y(n1091) );
  OR3X1_HVT U1301 ( .A1(n1081), .A2(n1091), .A3(n258), .Y(n1082) );
  NAND4X0_HVT U1302 ( .A1(n1093), .A2(n1084), .A3(n1083), .A4(n1082), .Y(n1085) );
  AO21X1_HVT U1303 ( .A1(n1086), .A2(n1096), .A3(n1085), .Y(n1089) );
  AO221X1_HVT U1304 ( .A1(n149), .A2(n197), .A3(n150), .A4(n258), .A5(n1087), 
        .Y(n1098) );
  AO21X1_HVT U1305 ( .A1(sram_raddr_b6[7]), .A2(n1090), .A3(sram_raddr_b6[8]), 
        .Y(n1088) );
  AO22X1_HVT U1306 ( .A1(n119), .A2(n1089), .A3(n1098), .A4(n1088), .Y(
        n_sram_raddr_b6[8]) );
  AO22X1_HVT U1307 ( .A1(n998), .A2(n175), .A3(n1304), .A4(n206), .Y(n1099) );
  AO221X1_HVT U1308 ( .A1(sram_raddr_b7[0]), .A2(n1194), .A3(n308), .A4(n1198), 
        .A5(n1099), .Y(n1100) );
  AO22X1_HVT U1309 ( .A1(n119), .A2(n1100), .A3(sram_raddr_b7[0]), .A4(n1270), 
        .Y(n_sram_raddr_b7[0]) );
  AO22X1_HVT U1310 ( .A1(n129), .A2(n1104), .A3(sram_raddr_b7[1]), .A4(n1270), 
        .Y(n_sram_raddr_b7[1]) );
  AO22X1_HVT U1311 ( .A1(sram_raddr_b7[2]), .A2(n125), .A3(n257), .A4(n1142), 
        .Y(n1107) );
  AO221X1_HVT U1312 ( .A1(sram_raddr_b4[2]), .A2(n1125), .A3(n246), .A4(n1124), 
        .A5(n154), .Y(n1105) );
  NAND3X0_HVT U1313 ( .A1(n1107), .A2(n1106), .A3(n1105), .Y(n1111) );
  OA221X1_HVT U1314 ( .A1(n1111), .A2(n1198), .A3(n1111), .A4(n1110), .A5(n129), .Y(n1112) );
  AO221X1_HVT U1315 ( .A1(sram_raddr_b7[2]), .A2(n162), .A3(n257), .A4(n148), 
        .A5(n1112), .Y(n_sram_raddr_b7[2]) );
  OA222X1_HVT U1316 ( .A1(sram_raddr_b4[3]), .A2(sram_raddr_b4[2]), .A3(
        sram_raddr_b4[3]), .A4(n1125), .A5(n1124), .A6(n1123), .Y(n1114) );
  AOI22X1_HVT U1317 ( .A1(n1304), .A2(n1114), .A3(n1113), .A4(n1198), .Y(n1118) );
  NAND3X0_HVT U1318 ( .A1(sram_raddr_b7[2]), .A2(n1183), .A3(n304), .Y(n1116)
         );
  AO221X1_HVT U1319 ( .A1(n125), .A2(sram_raddr_b7[2]), .A3(n126), .A4(n1142), 
        .A5(n304), .Y(n1115) );
  NAND4X0_HVT U1320 ( .A1(n1118), .A2(n1117), .A3(n1116), .A4(n1115), .Y(n1122) );
  NAND2X0_HVT U1321 ( .A1(n102), .A2(n257), .Y(n1119) );
  NAND2X0_HVT U1322 ( .A1(n1296), .A2(n1119), .Y(n1121) );
  AND2X1_HVT U1323 ( .A1(sram_raddr_b7[2]), .A2(n304), .Y(n1120) );
  AO222X1_HVT U1324 ( .A1(n1122), .A2(n127), .A3(n1121), .A4(sram_raddr_b7[3]), 
        .A5(n1120), .A6(n148), .Y(n_sram_raddr_b7[3]) );
  NAND3X0_HVT U1325 ( .A1(sram_raddr_b7[4]), .A2(sram_raddr_b7[3]), .A3(
        sram_raddr_b7[2]), .Y(n1156) );
  AO21X1_HVT U1326 ( .A1(sram_raddr_b7[3]), .A2(sram_raddr_b7[2]), .A3(
        sram_raddr_b7[4]), .Y(n1140) );
  NAND2X0_HVT U1327 ( .A1(n1156), .A2(n1140), .Y(n1134) );
  AO22X1_HVT U1328 ( .A1(n1183), .A2(n1134), .A3(sram_raddr_b7[4]), .A4(n1263), 
        .Y(n1132) );
  OA21X1_HVT U1329 ( .A1(n1124), .A2(n1123), .A3(n284), .Y(n1148) );
  AO21X1_HVT U1330 ( .A1(n1126), .A2(n1125), .A3(n1148), .Y(n1130) );
  AO22X1_HVT U1331 ( .A1(n1304), .A2(n1130), .A3(n1129), .A4(n1128), .Y(n1131)
         );
  OR3X1_HVT U1332 ( .A1(n1133), .A2(n1132), .A3(n1131), .Y(n1139) );
  AO222X1_HVT U1333 ( .A1(n1139), .A2(n128), .A3(n102), .A4(n1138), .A5(n162), 
        .A6(sram_raddr_b7[4]), .Y(n_sram_raddr_b7[4]) );
  OA21X1_HVT U1334 ( .A1(col[0]), .A2(n1141), .A3(n123), .Y(n1144) );
  NAND2X0_HVT U1335 ( .A1(n1141), .A2(n255), .Y(n1164) );
  OA22X1_HVT U1336 ( .A1(n1144), .A2(n255), .A3(n1142), .A4(n1164), .Y(n1154)
         );
  NAND2X0_HVT U1337 ( .A1(n1198), .A2(n1147), .Y(n1150) );
  NAND2X0_HVT U1338 ( .A1(n1148), .A2(n199), .Y(n1160) );
  AO221X1_HVT U1339 ( .A1(n1160), .A2(n1148), .A3(n1160), .A4(n199), .A5(n154), 
        .Y(n1149) );
  AND4X1_HVT U1340 ( .A1(n1154), .A2(n1151), .A3(n1150), .A4(n1149), .Y(n1155)
         );
  OA22X1_HVT U1341 ( .A1(n1155), .A2(n117), .A3(n99), .A4(n255), .Y(n1158) );
  AND4X1_HVT U1342 ( .A1(sram_raddr_b7[5]), .A2(sram_raddr_b7[4]), .A3(
        sram_raddr_b7[3]), .A4(sram_raddr_b7[2]), .Y(n1166) );
  NAND2X0_HVT U1343 ( .A1(n1158), .A2(n1157), .Y(n_sram_raddr_b7[5]) );
  NAND2X0_HVT U1344 ( .A1(sram_raddr_b7[6]), .A2(n1164), .Y(n1186) );
  AO22X1_HVT U1345 ( .A1(n1183), .A2(n1186), .A3(sram_raddr_b7[6]), .A4(n1263), 
        .Y(n1165) );
  NAND2X0_HVT U1346 ( .A1(sram_raddr_b4[6]), .A2(n1160), .Y(n1171) );
  OA21X1_HVT U1347 ( .A1(sram_raddr_b4[6]), .A2(n1160), .A3(n1171), .Y(n1162)
         );
  AO22X1_HVT U1348 ( .A1(n1304), .A2(n1162), .A3(n1161), .A4(n1198), .Y(n1163)
         );
  AO221X1_HVT U1349 ( .A1(n1165), .A2(sram_raddr_b7[6]), .A3(n1165), .A4(n1164), .A5(n1163), .Y(n1169) );
  NAND2X0_HVT U1350 ( .A1(sram_raddr_b7[6]), .A2(n1166), .Y(n1178) );
  OA21X1_HVT U1351 ( .A1(sram_raddr_b7[6]), .A2(n1166), .A3(n1178), .Y(n1167)
         );
  AO22X1_HVT U1352 ( .A1(n160), .A2(sram_raddr_b7[6]), .A3(n149), .A4(n1167), 
        .Y(n1168) );
  AO221X1_HVT U1353 ( .A1(n127), .A2(n1170), .A3(n129), .A4(n1169), .A5(n1168), 
        .Y(n_sram_raddr_b7[6]) );
  NAND3X0_HVT U1354 ( .A1(n1183), .A2(n198), .A3(n1186), .Y(n1175) );
  NAND2X0_HVT U1355 ( .A1(n269), .A2(n1171), .Y(n1184) );
  AO221X1_HVT U1356 ( .A1(n1184), .A2(n1171), .A3(n1184), .A4(n269), .A5(n154), 
        .Y(n1173) );
  AO221X1_HVT U1357 ( .A1(n125), .A2(col[0]), .A3(n123), .A4(n1186), .A5(n198), 
        .Y(n1172) );
  NAND4X0_HVT U1358 ( .A1(n1175), .A2(n1174), .A3(n1173), .A4(n1172), .Y(n1176) );
  AO21X1_HVT U1359 ( .A1(n1198), .A2(n1177), .A3(n1176), .Y(n1180) );
  NAND3X0_HVT U1360 ( .A1(sram_raddr_b7[7]), .A2(n1182), .A3(n99), .Y(n1181)
         );
  OA221X1_HVT U1361 ( .A1(sram_raddr_b7[7]), .A2(n149), .A3(sram_raddr_b7[7]), 
        .A4(n1182), .A5(n1181), .Y(n1179) );
  AO22X1_HVT U1362 ( .A1(n1537), .A2(n1180), .A3(n1179), .A4(n1270), .Y(
        n_sram_raddr_b7[7]) );
  OA22X1_HVT U1363 ( .A1(n162), .A2(n102), .A3(n1181), .A4(n280), .Y(n1204) );
  AND3X1_HVT U1364 ( .A1(n102), .A2(sram_raddr_b7[7]), .A3(n1182), .Y(n1205)
         );
  NAND4X0_HVT U1365 ( .A1(n1183), .A2(n280), .A3(n198), .A4(n1186), .Y(n1196)
         );
  NAND2X0_HVT U1366 ( .A1(n1185), .A2(n265), .Y(n1197) );
  AO221X1_HVT U1367 ( .A1(n1197), .A2(n1185), .A3(n1197), .A4(n265), .A5(n155), 
        .Y(n1188) );
  NAND3X0_HVT U1368 ( .A1(n123), .A2(n198), .A3(n1186), .Y(n1195) );
  NAND3X0_HVT U1369 ( .A1(sram_raddr_b7[8]), .A2(n1194), .A3(n1195), .Y(n1187)
         );
  NAND4X0_HVT U1370 ( .A1(n1196), .A2(n1189), .A3(n1188), .A4(n1187), .Y(n1191) );
  OA221X1_HVT U1371 ( .A1(n1191), .A2(n1198), .A3(n1191), .A4(n1190), .A5(n130), .Y(n1192) );
  AO221X1_HVT U1372 ( .A1(n1204), .A2(sram_raddr_b7[8]), .A3(n1204), .A4(n1205), .A5(n1192), .Y(n_sram_raddr_b7[8]) );
  OA21X1_HVT U1373 ( .A1(sram_raddr_b7[8]), .A2(n1195), .A3(n1194), .Y(n1203)
         );
  HADDX1_HVT U1374 ( .A0(n261), .B0(n1197), .SO(n1200) );
  AO22X1_HVT U1375 ( .A1(n1304), .A2(n1200), .A3(n1199), .A4(n1198), .Y(n1201)
         );
  AO221X1_HVT U1376 ( .A1(sram_raddr_b7[9]), .A2(n1203), .A3(n281), .A4(n1202), 
        .A5(n1201), .Y(n1207) );
  OA222X1_HVT U1377 ( .A1(sram_raddr_b7[9]), .A2(sram_raddr_b7[8]), .A3(
        sram_raddr_b7[9]), .A4(n1205), .A5(n1204), .A6(n281), .Y(n1206) );
  AO221X1_HVT U1378 ( .A1(n128), .A2(n1208), .A3(n130), .A4(n1207), .A5(n1206), 
        .Y(n_sram_raddr_b7[9]) );
  NAND2X0_HVT U1379 ( .A1(n1210), .A2(n1209), .Y(n1310) );
  AO22X1_HVT U1380 ( .A1(n998), .A2(n168), .A3(n1304), .A4(n207), .Y(n1211) );
  AO221X1_HVT U1381 ( .A1(sram_raddr_b8[0]), .A2(n1226), .A3(n309), .A4(n1310), 
        .A5(n1211), .Y(n1212) );
  AO22X1_HVT U1382 ( .A1(n119), .A2(n1212), .A3(sram_raddr_b8[0]), .A4(n1270), 
        .Y(n_sram_raddr_b8[0]) );
  AO22X1_HVT U1383 ( .A1(n128), .A2(n1216), .A3(sram_raddr_b8[1]), .A4(n1270), 
        .Y(n_sram_raddr_b8[1]) );
  AO22X1_HVT U1384 ( .A1(sram_raddr_b8[2]), .A2(n125), .A3(n170), .A4(n1249), 
        .Y(n1218) );
  AO221X1_HVT U1385 ( .A1(sram_raddr_b5[2]), .A2(n1241), .A3(n247), .A4(n1238), 
        .A5(n110), .Y(n1217) );
  NAND3X0_HVT U1386 ( .A1(n1219), .A2(n1218), .A3(n1217), .Y(n1221) );
  OA221X1_HVT U1387 ( .A1(n1221), .A2(n1310), .A3(n1221), .A4(n1220), .A5(n127), .Y(n1222) );
  AO221X1_HVT U1388 ( .A1(sram_raddr_b8[2]), .A2(n162), .A3(n170), .A4(n102), 
        .A5(n1222), .Y(n_sram_raddr_b8[2]) );
  OA222X1_HVT U1389 ( .A1(sram_raddr_b5[3]), .A2(sram_raddr_b5[2]), .A3(
        sram_raddr_b5[3]), .A4(n1241), .A5(n1238), .A6(n1237), .Y(n1224) );
  AOI22X1_HVT U1390 ( .A1(n1304), .A2(n1224), .A3(n1223), .A4(n1310), .Y(n1230) );
  NAND2X0_HVT U1391 ( .A1(n125), .A2(sram_raddr_b8[2]), .Y(n1225) );
  NAND3X0_HVT U1392 ( .A1(sram_raddr_b8[3]), .A2(n1226), .A3(n1225), .Y(n1228)
         );
  NAND3X0_HVT U1393 ( .A1(n1284), .A2(sram_raddr_b8[2]), .A3(n305), .Y(n1227)
         );
  NAND4X0_HVT U1394 ( .A1(n1230), .A2(n1229), .A3(n1228), .A4(n1227), .Y(n1234) );
  NAND2X0_HVT U1395 ( .A1(n148), .A2(n170), .Y(n1231) );
  NAND2X0_HVT U1396 ( .A1(n1296), .A2(n1231), .Y(n1233) );
  AND2X1_HVT U1397 ( .A1(sram_raddr_b8[2]), .A2(n305), .Y(n1232) );
  AO222X1_HVT U1398 ( .A1(n1234), .A2(n130), .A3(n1233), .A4(sram_raddr_b8[3]), 
        .A5(n1232), .A6(n102), .Y(n_sram_raddr_b8[3]) );
  NAND3X0_HVT U1399 ( .A1(sram_raddr_b8[4]), .A2(sram_raddr_b8[3]), .A3(
        sram_raddr_b8[2]), .Y(n1258) );
  OA21X1_HVT U1400 ( .A1(n305), .A2(n170), .A3(n208), .Y(n1248) );
  AND2X1_HVT U1401 ( .A1(n1258), .A2(n1235), .Y(n1246) );
  OA22X1_HVT U1402 ( .A1(n125), .A2(n208), .A3(n1246), .A4(n1249), .Y(n1245)
         );
  NAND2X0_HVT U1403 ( .A1(n1310), .A2(n1236), .Y(n1243) );
  OA21X1_HVT U1404 ( .A1(n1238), .A2(n1237), .A3(n252), .Y(n1252) );
  OAI221X1_HVT U1405 ( .A1(n1252), .A2(n1241), .A3(n1252), .A4(n1240), .A5(
        n1304), .Y(n1242) );
  NAND4X0_HVT U1406 ( .A1(n1245), .A2(n1244), .A3(n1243), .A4(n1242), .Y(n1247) );
  AO222X1_HVT U1407 ( .A1(n1247), .A2(n128), .A3(n103), .A4(n1246), .A5(n160), 
        .A6(sram_raddr_b8[4]), .Y(n_sram_raddr_b8[4]) );
  OA21X1_HVT U1408 ( .A1(col[1]), .A2(n1248), .A3(n124), .Y(n1250) );
  NAND2X0_HVT U1409 ( .A1(n1248), .A2(n256), .Y(n1264) );
  OA22X1_HVT U1410 ( .A1(n1250), .A2(n256), .A3(n1249), .A4(n1264), .Y(n1256)
         );
  NAND2X0_HVT U1411 ( .A1(n1310), .A2(n1251), .Y(n1254) );
  NAND2X0_HVT U1412 ( .A1(n1252), .A2(n193), .Y(n1274) );
  AO221X1_HVT U1413 ( .A1(n1274), .A2(n1252), .A3(n1274), .A4(n193), .A5(n155), 
        .Y(n1253) );
  AND4X1_HVT U1414 ( .A1(n1256), .A2(n1255), .A3(n1254), .A4(n1253), .Y(n1257)
         );
  OA22X1_HVT U1415 ( .A1(n1257), .A2(n118), .A3(n1296), .A4(n256), .Y(n1260)
         );
  AND4X1_HVT U1416 ( .A1(sram_raddr_b8[5]), .A2(sram_raddr_b8[4]), .A3(
        sram_raddr_b8[3]), .A4(sram_raddr_b8[2]), .Y(n1273) );
  NAND2X0_HVT U1417 ( .A1(n1260), .A2(n1259), .Y(n_sram_raddr_b8[5]) );
  NAND2X0_HVT U1418 ( .A1(n1261), .A2(n1310), .Y(n1268) );
  AO221X1_HVT U1419 ( .A1(sram_raddr_b5[6]), .A2(n1274), .A3(n295), .A4(n1262), 
        .A5(n155), .Y(n1267) );
  NAND2X0_HVT U1420 ( .A1(sram_raddr_b8[6]), .A2(n1264), .Y(n1287) );
  AND2X1_HVT U1421 ( .A1(n1284), .A2(n1287), .Y(n1265) );
  OAI222X1_HVT U1422 ( .A1(sram_raddr_b8[6]), .A2(n1265), .A3(sram_raddr_b8[6]), .A4(n1264), .A5(n1265), .A6(n1263), .Y(n1266) );
  NAND4X0_HVT U1423 ( .A1(n1269), .A2(n1268), .A3(n1267), .A4(n1266), .Y(n1272) );
  NAND3X0_HVT U1424 ( .A1(sram_raddr_b8[6]), .A2(n1273), .A3(n99), .Y(n1295)
         );
  AND2X1_HVT U1425 ( .A1(n1270), .A2(n1295), .Y(n1283) );
  AO21X1_HVT U1426 ( .A1(n102), .A2(n1273), .A3(sram_raddr_b8[6]), .Y(n1271)
         );
  AO22X1_HVT U1427 ( .A1(n128), .A2(n1272), .A3(n1283), .A4(n1271), .Y(
        n_sram_raddr_b8[6]) );
  AND3X1_HVT U1428 ( .A1(n148), .A2(sram_raddr_b8[6]), .A3(n1273), .Y(n1299)
         );
  NAND3X0_HVT U1429 ( .A1(n1284), .A2(n189), .A3(n1287), .Y(n1279) );
  NAND2X0_HVT U1430 ( .A1(sram_raddr_b5[6]), .A2(n1274), .Y(n1275) );
  NAND2X0_HVT U1431 ( .A1(n303), .A2(n1275), .Y(n1285) );
  AO221X1_HVT U1432 ( .A1(n1285), .A2(n1275), .A3(n1285), .A4(n303), .A5(n110), 
        .Y(n1277) );
  AO221X1_HVT U1433 ( .A1(n123), .A2(col[1]), .A3(n123), .A4(n1287), .A5(n189), 
        .Y(n1276) );
  NAND4X0_HVT U1434 ( .A1(n1279), .A2(n1278), .A3(n1277), .A4(n1276), .Y(n1281) );
  OA221X1_HVT U1435 ( .A1(n1281), .A2(n1310), .A3(n1281), .A4(n1280), .A5(n127), .Y(n1282) );
  AO221X1_HVT U1436 ( .A1(sram_raddr_b8[7]), .A2(n1283), .A3(n189), .A4(n1299), 
        .A5(n1282), .Y(n_sram_raddr_b8[7]) );
  NAND4X0_HVT U1437 ( .A1(n1284), .A2(n189), .A3(n260), .A4(n1287), .Y(n1302)
         );
  NAND2X0_HVT U1438 ( .A1(n1286), .A2(n187), .Y(n1305) );
  AO221X1_HVT U1439 ( .A1(n1305), .A2(n1286), .A3(n1305), .A4(n187), .A5(n110), 
        .Y(n1290) );
  AND3X1_HVT U1440 ( .A1(n124), .A2(n189), .A3(n1287), .Y(n1300) );
  OR3X1_HVT U1441 ( .A1(n1288), .A2(n1300), .A3(n260), .Y(n1289) );
  NAND4X0_HVT U1442 ( .A1(n1302), .A2(n1291), .A3(n1290), .A4(n1289), .Y(n1292) );
  AO21X1_HVT U1443 ( .A1(n1310), .A2(n1293), .A3(n1292), .Y(n1298) );
  NAND2X0_HVT U1444 ( .A1(sram_raddr_b8[8]), .A2(sram_raddr_b8[7]), .Y(n1294)
         );
  OA22X1_HVT U1445 ( .A1(n161), .A2(n150), .A3(n1295), .A4(n1294), .Y(n1315)
         );
  AO21X1_HVT U1446 ( .A1(sram_raddr_b8[7]), .A2(n1299), .A3(sram_raddr_b8[8]), 
        .Y(n1297) );
  AO22X1_HVT U1447 ( .A1(n1537), .A2(n1298), .A3(n1315), .A4(n1297), .Y(
        n_sram_raddr_b8[8]) );
  AND3X1_HVT U1448 ( .A1(sram_raddr_b8[8]), .A2(sram_raddr_b8[7]), .A3(n1299), 
        .Y(n1314) );
  AO22X1_HVT U1449 ( .A1(col[1]), .A2(n124), .A3(n1300), .A4(n260), .Y(n1303)
         );
  AO22X1_HVT U1450 ( .A1(sram_raddr_b8[9]), .A2(n1303), .A3(n288), .A4(n1302), 
        .Y(n1309) );
  AO221X1_HVT U1451 ( .A1(sram_raddr_b5[9]), .A2(n1306), .A3(n282), .A4(n1305), 
        .A5(n155), .Y(n1307) );
  NAND3X0_HVT U1452 ( .A1(n1309), .A2(n1308), .A3(n1307), .Y(n1312) );
  OA221X1_HVT U1453 ( .A1(n1312), .A2(n1311), .A3(n1312), .A4(n1310), .A5(n128), .Y(n1313) );
  AO221X1_HVT U1454 ( .A1(sram_raddr_b8[9]), .A2(n1315), .A3(n288), .A4(n1314), 
        .A5(n1313), .Y(n_sram_raddr_b8[9]) );
  OA221X1_HVT U1455 ( .A1(n1146), .A2(write_col[1]), .A3(n180), .A4(n235), 
        .A5(n1145), .Y(n1322) );
  OR2X1_HVT U1456 ( .A1(n1143), .A2(write_row[2]), .Y(n1316) );
  NAND3X0_HVT U1457 ( .A1(write_row[2]), .A2(n1143), .A3(n302), .Y(n1320) );
  AND4X1_HVT U1458 ( .A1(n1447), .A2(n1316), .A3(n302), .A4(n1320), .Y(n1317)
         );
  NAND2X0_HVT U1459 ( .A1(n1322), .A2(n1317), .Y(n_sram_write_enable_b0) );
  OA221X1_HVT U1460 ( .A1(write_col[1]), .A2(n181), .A3(n235), .A4(n1145), 
        .A5(n1146), .Y(n1323) );
  NAND2X0_HVT U1461 ( .A1(n1317), .A2(n1323), .Y(n_sram_write_enable_b1) );
  NAND3X0_HVT U1462 ( .A1(write_col[1]), .A2(n1146), .A3(n181), .Y(n1449) );
  NAND3X0_HVT U1463 ( .A1(n1145), .A2(n180), .A3(n235), .Y(n1453) );
  NAND2X0_HVT U1464 ( .A1(n1449), .A2(n1453), .Y(n1446) );
  NAND2X0_HVT U1465 ( .A1(n1317), .A2(n1446), .Y(n_sram_write_enable_b2) );
  OR3X1_HVT U1466 ( .A1(n1143), .A2(write_row[2]), .A3(n302), .Y(n1321) );
  NAND2X0_HVT U1467 ( .A1(n1143), .A2(n302), .Y(n1318) );
  AND4X1_HVT U1468 ( .A1(n1447), .A2(n382), .A3(n1321), .A4(n1318), .Y(n1319)
         );
  NAND2X0_HVT U1469 ( .A1(n1322), .A2(n1319), .Y(n_sram_write_enable_b3) );
  NAND2X0_HVT U1470 ( .A1(n1323), .A2(n1319), .Y(n_sram_write_enable_b4) );
  NAND2X0_HVT U1471 ( .A1(n1319), .A2(n1446), .Y(n_sram_write_enable_b5) );
  NAND2X0_HVT U1472 ( .A1(n1321), .A2(n1320), .Y(n1450) );
  NAND3X0_HVT U1473 ( .A1(n1447), .A2(n1322), .A3(n1450), .Y(
        n_sram_write_enable_b6) );
  NAND3X0_HVT U1474 ( .A1(n1447), .A2(n1323), .A3(n1450), .Y(
        n_sram_write_enable_b7) );
  NAND3X0_HVT U1475 ( .A1(n1447), .A2(n1450), .A3(n1446), .Y(
        n_sram_write_enable_b8) );
  AND4X1_HVT U1476 ( .A1(n1324), .A2(n1153), .A3(delay2_write_enable), .A4(
        n1152), .Y(n1326) );
  NAND3X0_HVT U1477 ( .A1(n1326), .A2(n1492), .A3(n353), .Y(
        n_sram_write_enable_c0) );
  NAND3X0_HVT U1478 ( .A1(delay2_addr_change_2_), .A2(n1326), .A3(n1492), .Y(
        n_sram_write_enable_c1) );
  AND4X1_HVT U1479 ( .A1(n1324), .A2(delay2_write_enable), .A3(n1152), .A4(
        n357), .Y(n1327) );
  NAND3X0_HVT U1480 ( .A1(n1327), .A2(n1492), .A3(n353), .Y(
        n_sram_write_enable_c2) );
  NAND3X0_HVT U1481 ( .A1(delay2_addr_change_2_), .A2(n1327), .A3(n1492), .Y(
        n_sram_write_enable_c3) );
  NAND2X0_HVT U1482 ( .A1(n1324), .A2(delay2_write_enable), .Y(n1325) );
  NAND2X0_HVT U1483 ( .A1(n1328), .A2(n1492), .Y(n_sram_write_enable_c4) );
  NAND3X0_HVT U1484 ( .A1(mem_sel), .A2(n1326), .A3(n353), .Y(
        n_sram_write_enable_d0) );
  NAND3X0_HVT U1485 ( .A1(mem_sel), .A2(delay2_addr_change_2_), .A3(n1326), 
        .Y(n_sram_write_enable_d1) );
  NAND3X0_HVT U1486 ( .A1(mem_sel), .A2(n1327), .A3(n353), .Y(
        n_sram_write_enable_d2) );
  NAND3X0_HVT U1487 ( .A1(mem_sel), .A2(delay2_addr_change_2_), .A3(n1327), 
        .Y(n_sram_write_enable_d3) );
  NAND2X0_HVT U1488 ( .A1(mem_sel), .A2(n1328), .Y(n_sram_write_enable_d4) );
  NAND4X0_HVT U1489 ( .A1(state[0]), .A2(n1108), .A3(n1109), .A4(n177), .Y(
        n1333) );
  NAND3X0_HVT U1490 ( .A1(n1445), .A2(n166), .A3(n177), .Y(n1490) );
  NAND2X0_HVT U1491 ( .A1(n1528), .A2(conv_done), .Y(n1338) );
  NAND4X0_HVT U1492 ( .A1(n1108), .A2(n1109), .A3(n1329), .A4(n166), .Y(n1330)
         );
  AND4X1_HVT U1493 ( .A1(n1336), .A2(n1490), .A3(n1338), .A4(n1330), .Y(n1332)
         );
  NAND3X0_HVT U1494 ( .A1(n1979), .A2(n178), .A3(n369), .Y(n1331) );
  NAND4X0_HVT U1495 ( .A1(n1332), .A2(n1334), .A3(n1333), .A4(n1331), .Y(
        n_state[0]) );
  OA22X1_HVT U1496 ( .A1(conv1_done), .A2(n1363), .A3(conv_done), .A4(n1336), 
        .Y(n1335) );
  NAND3X0_HVT U1497 ( .A1(state[0]), .A2(n1445), .A3(n177), .Y(n1441) );
  NAND4X0_HVT U1498 ( .A1(n1335), .A2(n1334), .A3(n1333), .A4(n1441), .Y(
        n_state[1]) );
  OA22X1_HVT U1499 ( .A1(conv_done), .A2(n1336), .A3(n1363), .A4(n369), .Y(
        n1337) );
  NAND2X0_HVT U1500 ( .A1(n1445), .A2(n177), .Y(n1431) );
  NAND2X0_HVT U1501 ( .A1(n1337), .A2(n1431), .Y(n_state[2]) );
  NAND2X0_HVT U1502 ( .A1(state[1]), .A2(n1445), .Y(n1340) );
  NAND3X0_HVT U1503 ( .A1(n1340), .A2(n1339), .A3(n1338), .Y(n_state[3]) );
  NAND3X0_HVT U1504 ( .A1(n1435), .A2(n1434), .A3(n1341), .Y(n1352) );
  NAND2X0_HVT U1505 ( .A1(n1433), .A2(n1342), .Y(n1356) );
  AO22X1_HVT U1506 ( .A1(weight_cnt[0]), .A2(n1352), .A3(n227), .A4(n1356), 
        .Y(n_weight_cnt[0]) );
  AO22X1_HVT U1507 ( .A1(weight_cnt[1]), .A2(n227), .A3(n354), .A4(
        weight_cnt[0]), .Y(n1343) );
  AO22X1_HVT U1508 ( .A1(n1343), .A2(n1356), .A3(weight_cnt[1]), .A4(n1352), 
        .Y(n_weight_cnt[1]) );
  AND3X1_HVT U1509 ( .A1(weight_cnt[1]), .A2(weight_cnt[0]), .A3(n1356), .Y(
        n1349) );
  NAND3X0_HVT U1510 ( .A1(weight_cnt[1]), .A2(weight_cnt[0]), .A3(
        weight_cnt[2]), .Y(n1345) );
  AO21X1_HVT U1511 ( .A1(n1356), .A2(n1345), .A3(n1352), .Y(n1344) );
  OA21X1_HVT U1512 ( .A1(weight_cnt[2]), .A2(n1349), .A3(n1344), .Y(
        n_weight_cnt[2]) );
  AND4X1_HVT U1513 ( .A1(weight_cnt[1]), .A2(weight_cnt[0]), .A3(weight_cnt[2]), .A4(n1356), .Y(n1347) );
  AO22X1_HVT U1514 ( .A1(weight_cnt[3]), .A2(n1344), .A3(n176), .A4(n1347), 
        .Y(n_weight_cnt[3]) );
  NAND3X0_HVT U1515 ( .A1(weight_cnt[3]), .A2(n1346), .A3(weight_cnt[4]), .Y(
        n1351) );
  AO21X1_HVT U1516 ( .A1(n1356), .A2(n1351), .A3(n1352), .Y(n1348) );
  OA221X1_HVT U1517 ( .A1(weight_cnt[4]), .A2(n1347), .A3(weight_cnt[4]), .A4(
        weight_cnt[3]), .A5(n1348), .Y(n_weight_cnt[4]) );
  AND4X1_HVT U1518 ( .A1(weight_cnt[2]), .A2(weight_cnt[3]), .A3(weight_cnt[4]), .A4(n275), .Y(n1350) );
  AO22X1_HVT U1519 ( .A1(n1350), .A2(n1349), .A3(weight_cnt[5]), .A4(n1348), 
        .Y(n_weight_cnt[5]) );
  NOR2X0_HVT U1520 ( .A1(n1351), .A2(n275), .Y(n1353) );
  OR3X1_HVT U1521 ( .A1(n1351), .A2(n275), .A3(n213), .Y(n1354) );
  AO21X1_HVT U1522 ( .A1(n1356), .A2(n1354), .A3(n1352), .Y(n1355) );
  OA221X1_HVT U1523 ( .A1(weight_cnt[6]), .A2(n1353), .A3(weight_cnt[6]), .A4(
        n1356), .A5(n1355), .Y(n_weight_cnt[6]) );
  OA222X1_HVT U1524 ( .A1(weight_cnt[7]), .A2(n1357), .A3(weight_cnt[7]), .A4(
        n1356), .A5(n324), .A6(n1355), .Y(n_weight_cnt[7]) );
  OR3X1_HVT U1525 ( .A1(write_enable), .A2(conv2_weight_done), .A3(
        load_data_enable), .Y(n1359) );
  OR3X1_HVT U1526 ( .A1(conv1_weight_done), .A2(write_enable), .A3(
        load_data_enable), .Y(n1358) );
  AO22X1_HVT U1527 ( .A1(n1528), .A2(n1359), .A3(n1979), .A4(n1358), .Y(
        n_write_enable) );
  NAND2X0_HVT U1528 ( .A1(n1528), .A2(n107), .Y(net19513) );
  NAND3X0_HVT U1529 ( .A1(col[2]), .A2(col[1]), .A3(col[0]), .Y(n1541) );
  OA221X1_HVT U1530 ( .A1(n1361), .A2(col[3]), .A3(n1541), .A4(n163), .A5(
        n1543), .Y(net19699) );
  AND2X1_HVT U1531 ( .A1(n1543), .A2(n1362), .Y(net19709) );
  AND2X1_HVT U1532 ( .A1(n194), .A2(n1543), .Y(net19714) );
  AO221X1_HVT U1533 ( .A1(sram_raddr_weight[4]), .A2(sram_raddr_weight[3]), 
        .A3(sram_raddr_weight[4]), .A4(sram_raddr_weight[2]), .A5(n1364), .Y(
        n1414) );
  NAND2X0_HVT U1534 ( .A1(n1417), .A2(n315), .Y(n1408) );
  OR3X1_HVT U1535 ( .A1(sram_raddr_weight[7]), .A2(sram_raddr_weight[8]), .A3(
        n1408), .Y(n1394) );
  AND2X1_HVT U1536 ( .A1(n1387), .A2(n319), .Y(n1376) );
  NAND2X0_HVT U1537 ( .A1(n1376), .A2(n320), .Y(n1375) );
  OR3X1_HVT U1538 ( .A1(n1375), .A2(n98), .A3(sram_raddr_weight[14]), .Y(n1371) );
  NAND2X0_HVT U1539 ( .A1(n355), .A2(n1371), .Y(n1369) );
  NAND4X0_HVT U1540 ( .A1(sram_raddr_weight[3]), .A2(sram_raddr_weight[2]), 
        .A3(sram_raddr_weight[0]), .A4(sram_raddr_weight[1]), .Y(n1419) );
  NAND2X0_HVT U1541 ( .A1(sram_raddr_weight[4]), .A2(n1423), .Y(n1413) );
  AND2X1_HVT U1542 ( .A1(sram_raddr_weight[5]), .A2(n1416), .Y(n1410) );
  AND2X1_HVT U1543 ( .A1(sram_raddr_weight[6]), .A2(n1410), .Y(n1403) );
  NAND2X0_HVT U1544 ( .A1(sram_raddr_weight[7]), .A2(n1403), .Y(n1395) );
  NAND2X0_HVT U1545 ( .A1(sram_raddr_weight[8]), .A2(n1398), .Y(n1397) );
  NAND4X0_HVT U1546 ( .A1(sram_raddr_weight[11]), .A2(sram_raddr_weight[9]), 
        .A3(sram_raddr_weight[10]), .A4(n1391), .Y(n1380) );
  AND4X1_HVT U1547 ( .A1(sram_raddr_weight[12]), .A2(sram_raddr_weight[13]), 
        .A3(n1382), .A4(n1443), .Y(n1373) );
  NAND2X0_HVT U1548 ( .A1(sram_raddr_weight[14]), .A2(n1373), .Y(n1367) );
  NAND2X0_HVT U1549 ( .A1(sram_raddr_weight[15]), .A2(n1367), .Y(n1366) );
  AO22X1_HVT U1550 ( .A1(n119), .A2(n1375), .A3(n1443), .A4(n1367), .Y(n1374)
         );
  AO21X1_HVT U1551 ( .A1(n127), .A2(sram_raddr_weight[14]), .A3(n1374), .Y(
        n1368) );
  AO221X1_HVT U1552 ( .A1(sram_raddr_weight[15]), .A2(n119), .A3(n355), .A4(
        n1443), .A5(n1368), .Y(n1365) );
  OA222X1_HVT U1553 ( .A1(sram_raddr_weight[16]), .A2(n1369), .A3(
        sram_raddr_weight[16]), .A4(n1366), .A5(n381), .A6(n1365), .Y(net19752) );
  OA22X1_HVT U1554 ( .A1(n1370), .A2(n1369), .A3(n355), .A4(n1368), .Y(
        net19759) );
  AO221X1_HVT U1555 ( .A1(n1374), .A2(sram_raddr_weight[14]), .A3(n1374), .A4(
        n1373), .A5(n1372), .Y(net19766) );
  NAND3X0_HVT U1556 ( .A1(sram_raddr_weight[13]), .A2(sram_raddr_weight[12]), 
        .A3(n1382), .Y(n1377) );
  OA221X1_HVT U1557 ( .A1(sram_raddr_weight[13]), .A2(sram_raddr_weight[12]), 
        .A3(sram_raddr_weight[13]), .A4(n1382), .A5(n1377), .Y(n1378) );
  AO22X1_HVT U1558 ( .A1(n1537), .A2(n1379), .A3(n1378), .A4(n1443), .Y(
        net19773) );
  OR3X1_HVT U1559 ( .A1(sram_raddr_weight[9]), .A2(sram_raddr_weight[10]), 
        .A3(n1394), .Y(n1381) );
  AO22X1_HVT U1560 ( .A1(n130), .A2(n1381), .A3(n1443), .A4(n1380), .Y(n1386)
         );
  AO21X1_HVT U1561 ( .A1(n128), .A2(sram_raddr_weight[11]), .A3(n1386), .Y(
        n1384) );
  AO22X1_HVT U1562 ( .A1(n1537), .A2(n1387), .A3(n1382), .A4(n1443), .Y(n1383)
         );
  AO22X1_HVT U1563 ( .A1(sram_raddr_weight[12]), .A2(n1384), .A3(n319), .A4(
        n1383), .Y(net19780) );
  AND3X1_HVT U1564 ( .A1(sram_raddr_weight[9]), .A2(n1391), .A3(n1443), .Y(
        n1389) );
  AO21X1_HVT U1565 ( .A1(sram_raddr_weight[10]), .A2(n1389), .A3(
        sram_raddr_weight[11]), .Y(n1385) );
  AO22X1_HVT U1566 ( .A1(n127), .A2(n1387), .A3(n1386), .A4(n1385), .Y(
        net19787) );
  NOR3X0_HVT U1567 ( .A1(sram_raddr_weight[9]), .A2(n1394), .A3(n117), .Y(
        n1393) );
  AO22X1_HVT U1568 ( .A1(n129), .A2(n1394), .A3(n1443), .A4(n1397), .Y(n1390)
         );
  AO221X1_HVT U1569 ( .A1(sram_raddr_weight[9]), .A2(n1537), .A3(n296), .A4(
        n1443), .A5(n1390), .Y(n1388) );
  AO222X1_HVT U1570 ( .A1(n356), .A2(n1389), .A3(n356), .A4(n1393), .A5(
        sram_raddr_weight[10]), .A6(n1388), .Y(net19794) );
  OA222X1_HVT U1571 ( .A1(sram_raddr_weight[9]), .A2(n1391), .A3(
        sram_raddr_weight[9]), .A4(n1443), .A5(n296), .A6(n1390), .Y(n1392) );
  OR3X1_HVT U1572 ( .A1(n1393), .A2(n1418), .A3(n1392), .Y(net19808) );
  OR2X1_HVT U1573 ( .A1(n98), .A2(n1394), .Y(n1401) );
  AND2X1_HVT U1574 ( .A1(n1443), .A2(n1395), .Y(n1402) );
  AO221X1_HVT U1575 ( .A1(n119), .A2(sram_raddr_weight[7]), .A3(n1537), .A4(
        n1408), .A5(n1402), .Y(n1396) );
  NAND2X0_HVT U1576 ( .A1(sram_raddr_weight[8]), .A2(n1396), .Y(n1400) );
  NAND3X0_HVT U1577 ( .A1(n1398), .A2(n1443), .A3(n1397), .Y(n1399) );
  NAND4X0_HVT U1578 ( .A1(n1401), .A2(n1431), .A3(n1400), .A4(n1399), .Y(
        net19815) );
  NAND2X0_HVT U1579 ( .A1(n1402), .A2(n1403), .Y(n1407) );
  OA22X1_HVT U1580 ( .A1(n1404), .A2(n98), .A3(n1435), .A4(n1403), .Y(n1405)
         );
  AO222X1_HVT U1581 ( .A1(n318), .A2(n98), .A3(n318), .A4(n1408), .A5(
        sram_raddr_weight[7]), .A6(n1405), .Y(n1406) );
  NAND3X0_HVT U1582 ( .A1(n1407), .A2(n1406), .A3(n1431), .Y(net19843) );
  OA22X1_HVT U1583 ( .A1(n1417), .A2(n118), .A3(n1435), .A4(n1410), .Y(n1409)
         );
  OA22X1_HVT U1584 ( .A1(n1409), .A2(n315), .A3(n98), .A4(n1408), .Y(n1412) );
  NAND3X0_HVT U1585 ( .A1(n1410), .A2(n315), .A3(n1443), .Y(n1411) );
  NAND3X0_HVT U1586 ( .A1(n1412), .A2(n1431), .A3(n1411), .Y(net19850) );
  AO22X1_HVT U1587 ( .A1(n128), .A2(n1414), .A3(n1443), .A4(n1413), .Y(n1415)
         );
  AND3X1_HVT U1588 ( .A1(state[1]), .A2(n1445), .A3(n166), .Y(n1737) );
  NAND2X0_HVT U1589 ( .A1(n1443), .A2(n1419), .Y(n1427) );
  NAND4X0_HVT U1590 ( .A1(n119), .A2(n1420), .A3(n321), .A4(n209), .Y(n1430)
         );
  NAND3X0_HVT U1591 ( .A1(n1433), .A2(n1427), .A3(n1430), .Y(n1425) );
  NAND2X0_HVT U1592 ( .A1(n1420), .A2(n209), .Y(n1426) );
  OR2X1_HVT U1593 ( .A1(sram_raddr_weight[3]), .A2(n1426), .Y(n1421) );
  AO22X1_HVT U1594 ( .A1(n1423), .A2(n1443), .A3(n1422), .A4(n1421), .Y(n1424)
         );
  AND4X1_HVT U1595 ( .A1(n1108), .A2(n1109), .A3(n166), .A4(n177), .Y(n1529)
         );
  AO221X1_HVT U1596 ( .A1(n1445), .A2(n177), .A3(n1445), .A4(n166), .A5(n1529), 
        .Y(n1437) );
  AO221X1_HVT U1597 ( .A1(sram_raddr_weight[4]), .A2(n1425), .A3(n374), .A4(
        n1424), .A5(n1437), .Y(net19871) );
  NAND3X0_HVT U1598 ( .A1(sram_raddr_weight[2]), .A2(sram_raddr_weight[0]), 
        .A3(sram_raddr_weight[1]), .Y(n1428) );
  AOI22X1_HVT U1599 ( .A1(n128), .A2(n1426), .A3(n1443), .A4(n1428), .Y(n1429)
         );
  OA22X1_HVT U1600 ( .A1(n1429), .A2(n321), .A3(n1428), .A4(n1427), .Y(n1432)
         );
  NAND3X0_HVT U1601 ( .A1(n1432), .A2(n1431), .A3(n1430), .Y(net19878) );
  NAND2X0_HVT U1602 ( .A1(sram_raddr_weight[0]), .A2(sram_raddr_weight[1]), 
        .Y(n1436) );
  NAND2X0_HVT U1603 ( .A1(n1443), .A2(n1436), .Y(n1440) );
  NAND2X0_HVT U1604 ( .A1(n1433), .A2(n1440), .Y(n1439) );
  OAI21X1_HVT U1605 ( .A1(n1436), .A2(n1435), .A3(n1434), .Y(n1438) );
  AO221X1_HVT U1606 ( .A1(sram_raddr_weight[2]), .A2(n1439), .A3(n209), .A4(
        n1438), .A5(n1437), .Y(net19885) );
  AO222X1_HVT U1607 ( .A1(n364), .A2(n1440), .A3(n364), .A4(n231), .A5(n1440), 
        .A6(n118), .Y(n1442) );
  NAND2X0_HVT U1608 ( .A1(n1442), .A2(n1441), .Y(net19899) );
  AO21X1_HVT U1609 ( .A1(state[1]), .A2(sram_raddr_weight[0]), .A3(n166), .Y(
        n1444) );
  AO22X1_HVT U1610 ( .A1(n1445), .A2(n1444), .A3(n1443), .A4(n231), .Y(
        net19913) );
  NAND2X0_HVT U1611 ( .A1(write_col[0]), .A2(n1446), .Y(n1489) );
  AO21X1_HVT U1612 ( .A1(n1448), .A2(n1447), .A3(N2888), .Y(net19921) );
  NAND2X0_HVT U1613 ( .A1(write_row[0]), .A2(n1450), .Y(n1454) );
  NAND3X0_HVT U1614 ( .A1(write_col[0]), .A2(n1451), .A3(n1454), .Y(n1458) );
  OR3X1_HVT U1615 ( .A1(delay1_sram_waddr_b[0]), .A2(delay1_sram_waddr_b[1]), 
        .A3(delay1_sram_waddr_b[2]), .Y(n1478) );
  OR3X1_HVT U1616 ( .A1(delay1_sram_waddr_b[4]), .A2(delay1_sram_waddr_b[3]), 
        .A3(n1478), .Y(n1472) );
  OR3X1_HVT U1617 ( .A1(delay1_sram_waddr_b[6]), .A2(delay1_sram_waddr_b[5]), 
        .A3(n1472), .Y(n1467) );
  NOR2X0_HVT U1618 ( .A1(n1467), .A2(delay1_sram_waddr_b[7]), .Y(n1463) );
  NAND2X0_HVT U1619 ( .A1(n1463), .A2(n328), .Y(n1452) );
  HADDX1_HVT U1620 ( .A0(delay1_sram_waddr_b[9]), .B0(n1452), .SO(n1457) );
  NAND3X0_HVT U1621 ( .A1(delay1_sram_waddr_b[0]), .A2(delay1_sram_waddr_b[1]), 
        .A3(delay1_sram_waddr_b[2]), .Y(n1482) );
  NAND3X0_HVT U1622 ( .A1(delay1_sram_waddr_b[4]), .A2(delay1_sram_waddr_b[3]), 
        .A3(n1479), .Y(n1476) );
  NAND3X0_HVT U1623 ( .A1(delay1_sram_waddr_b[6]), .A2(delay1_sram_waddr_b[5]), 
        .A3(n1473), .Y(n1469) );
  AND2X1_HVT U1624 ( .A1(delay1_sram_waddr_b[7]), .A2(n1465), .Y(n1462) );
  NAND2X0_HVT U1625 ( .A1(delay1_sram_waddr_b[8]), .A2(n1462), .Y(n1455) );
  HADDX1_HVT U1626 ( .A0(delay1_sram_waddr_b[9]), .B0(n1455), .SO(n1456) );
  OAI22X1_HVT U1627 ( .A1(n1458), .A2(n1457), .A3(n1461), .A4(n1456), .Y(
        net19924) );
  OAI22X1_HVT U1628 ( .A1(n1463), .A2(n1458), .A3(n1462), .A4(n1461), .Y(n1460) );
  AO22X1_HVT U1629 ( .A1(n1487), .A2(n1463), .A3(n1488), .A4(n1462), .Y(n1459)
         );
  AO22X1_HVT U1630 ( .A1(delay1_sram_waddr_b[8]), .A2(n1460), .A3(n328), .A4(
        n1459), .Y(net19927) );
  OA221X1_HVT U1631 ( .A1(n1463), .A2(delay1_sram_waddr_b[7]), .A3(n1463), 
        .A4(n1467), .A5(n1487), .Y(n1464) );
  AO221X1_HVT U1632 ( .A1(n1466), .A2(delay1_sram_waddr_b[7]), .A3(n1466), 
        .A4(n1465), .A5(n1464), .Y(net19930) );
  AO221X1_HVT U1633 ( .A1(delay1_sram_waddr_b[6]), .A2(delay1_sram_waddr_b[5]), 
        .A3(delay1_sram_waddr_b[6]), .A4(n1472), .A5(n1468), .Y(n1471) );
  OA221X1_HVT U1634 ( .A1(delay1_sram_waddr_b[6]), .A2(delay1_sram_waddr_b[5]), 
        .A3(delay1_sram_waddr_b[6]), .A4(n1473), .A5(n1469), .Y(n1470) );
  AO22X1_HVT U1635 ( .A1(n1487), .A2(n1471), .A3(n1488), .A4(n1470), .Y(
        net19933) );
  AO22X1_HVT U1636 ( .A1(n1487), .A2(n1472), .A3(n1488), .A4(n1476), .Y(n1475)
         );
  AO22X1_HVT U1637 ( .A1(n1487), .A2(n1477), .A3(n1488), .A4(n1473), .Y(n1474)
         );
  AO22X1_HVT U1638 ( .A1(delay1_sram_waddr_b[5]), .A2(n1475), .A3(n365), .A4(
        n1474), .Y(net19936) );
  AO22X1_HVT U1639 ( .A1(n1487), .A2(n1478), .A3(n1488), .A4(n1482), .Y(n1481)
         );
  AO22X1_HVT U1640 ( .A1(n1487), .A2(n1483), .A3(n1488), .A4(n1479), .Y(n1480)
         );
  AO22X1_HVT U1641 ( .A1(delay1_sram_waddr_b[3]), .A2(n1481), .A3(n366), .A4(
        n1480), .Y(net19942) );
  NAND2X0_HVT U1642 ( .A1(delay1_sram_waddr_b[0]), .A2(delay1_sram_waddr_b[1]), 
        .Y(n1484) );
  OR2X1_HVT U1643 ( .A1(delay1_sram_waddr_b[0]), .A2(delay1_sram_waddr_b[1]), 
        .Y(n1485) );
  NAND2X0_HVT U1644 ( .A1(n1485), .A2(n1484), .Y(n1486) );
  MUX21X1_HVT U1645 ( .A1(n1488), .A2(n1487), .S0(n1486), .Y(net19948) );
  NOR2X0_HVT U1646 ( .A1(n1489), .A2(delay1_sram_waddr_b[0]), .Y(net19951) );
  NAND2X0_HVT U1647 ( .A1(addr_change[0]), .A2(addr_change[1]), .Y(n1535) );
  NAND4X0_HVT U1648 ( .A1(addr_change[4]), .A2(n1534), .A3(n182), .A4(n236), 
        .Y(n1530) );
  OR2X1_HVT U1649 ( .A1(n1530), .A2(n118), .Y(n1491) );
  NAND3X0_HVT U1650 ( .A1(n1491), .A2(n106), .A3(n1490), .Y(net19959) );
  NAND4X0_HVT U1651 ( .A1(delay1_sram_waddr_c[0]), .A2(delay1_sram_waddr_c[1]), 
        .A3(delay1_sram_waddr_c[2]), .A4(delay1_sram_waddr_c[3]), .Y(n1504) );
  NAND2X0_HVT U1652 ( .A1(n1503), .A2(delay1_sram_waddr_c[4]), .Y(n1502) );
  NAND2X0_HVT U1653 ( .A1(n1501), .A2(delay1_sram_waddr_c[5]), .Y(n1500) );
  NAND2X0_HVT U1654 ( .A1(n1499), .A2(delay1_sram_waddr_c[6]), .Y(n1498) );
  NAND2X0_HVT U1655 ( .A1(n1497), .A2(delay1_sram_waddr_c[7]), .Y(n1496) );
  NAND2X0_HVT U1656 ( .A1(n1495), .A2(delay1_sram_waddr_c[8]), .Y(n1494) );
  OA221X1_HVT U1657 ( .A1(n1493), .A2(delay1_sram_waddr_c[9]), .A3(n1494), 
        .A4(n384), .A5(n1507), .Y(net19961) );
  NAND3X0_HVT U1658 ( .A1(delay1_sram_waddr_c[0]), .A2(delay1_sram_waddr_c[1]), 
        .A3(delay1_sram_waddr_c[2]), .Y(n1505) );
  NAND2X0_HVT U1659 ( .A1(delay1_sram_waddr_c[0]), .A2(delay1_sram_waddr_c[1]), 
        .Y(n1506) );
  AND2X1_HVT U1660 ( .A1(n1507), .A2(n370), .Y(net19970) );
  NAND4X0_HVT U1661 ( .A1(delay1_sram_waddr_d[0]), .A2(delay1_sram_waddr_d[1]), 
        .A3(delay1_sram_waddr_d[2]), .A4(delay1_sram_waddr_d[3]), .Y(n1519) );
  NAND2X0_HVT U1662 ( .A1(n1518), .A2(delay1_sram_waddr_d[4]), .Y(n1517) );
  NAND2X0_HVT U1663 ( .A1(n1516), .A2(delay1_sram_waddr_d[5]), .Y(n1515) );
  NAND2X0_HVT U1664 ( .A1(n1514), .A2(delay1_sram_waddr_d[6]), .Y(n1513) );
  NAND2X0_HVT U1665 ( .A1(n1512), .A2(delay1_sram_waddr_d[7]), .Y(n1511) );
  NAND2X0_HVT U1666 ( .A1(n1510), .A2(delay1_sram_waddr_d[8]), .Y(n1509) );
  OA221X1_HVT U1667 ( .A1(n1508), .A2(delay1_sram_waddr_d[9]), .A3(n1509), 
        .A4(n385), .A5(n1522), .Y(net19977) );
  NAND3X0_HVT U1668 ( .A1(delay1_sram_waddr_d[0]), .A2(delay1_sram_waddr_d[1]), 
        .A3(delay1_sram_waddr_d[2]), .Y(n1520) );
  NAND2X0_HVT U1669 ( .A1(delay1_sram_waddr_d[0]), .A2(delay1_sram_waddr_d[1]), 
        .Y(n1521) );
  AND2X1_HVT U1670 ( .A1(n1522), .A2(n371), .Y(net19986) );
  NAND2X0_HVT U1671 ( .A1(n1523), .A2(n106), .Y(net19993) );
  NAND3X0_HVT U1672 ( .A1(n1526), .A2(channel_cnt[2]), .A3(channel_cnt[3]), 
        .Y(n1525) );
  OA221X1_HVT U1673 ( .A1(channel_cnt[4]), .A2(n1524), .A3(n233), .A4(n1525), 
        .A5(n1528), .Y(net19994) );
  OA221X1_HVT U1674 ( .A1(n1526), .A2(channel_cnt[2]), .A3(n1527), .A4(n363), 
        .A5(n1528), .Y(net19996) );
  OR3X1_HVT U1675 ( .A1(n127), .A2(n1529), .A3(n157), .Y(net20004) );
  NAND4X0_HVT U1676 ( .A1(addr_change[0]), .A2(addr_change[1]), .A3(
        addr_change[2]), .A4(addr_change[3]), .Y(n1532) );
  OA221X1_HVT U1677 ( .A1(addr_change[4]), .A2(n1531), .A3(n380), .A4(n1532), 
        .A5(n1533), .Y(net20006) );
  OA221X1_HVT U1678 ( .A1(n1534), .A2(addr_change[2]), .A3(n1535), .A4(n182), 
        .A5(n1533), .Y(net20008) );
  NAND3X0_HVT U1679 ( .A1(n1979), .A2(n1653), .A3(n178), .Y(n1539) );
  NAND4X0_HVT U1680 ( .A1(addr_row_sel_cnt[0]), .A2(n1545), .A3(n1654), .A4(
        addr_row_sel_cnt[1]), .Y(n1538) );
  NAND2X0_HVT U1681 ( .A1(n107), .A2(n1920), .Y(net20953) );
  NAND2X0_HVT U1682 ( .A1(n106), .A2(n1967), .Y(net22280) );
  OA221X1_HVT U1683 ( .A1(n1539), .A2(n1136), .A3(n1539), .A4(n1135), .A5(
        n1538), .Y(n1742) );
  NAND2X0_HVT U1684 ( .A1(n105), .A2(n108), .Y(net23610) );
  NAND2X0_HVT U1685 ( .A1(n_addr_col_sel_cnt[0]), .A2(n178), .Y(n1853) );
  AND4X1_HVT U1686 ( .A1(n1545), .A2(n1979), .A3(addr_row_sel_cnt[1]), .A4(
        n178), .Y(n1547) );
  AO22X1_HVT U1687 ( .A1(n1827), .A2(n228), .A3(n95), .A4(n360), .Y(n1548) );
  AO221X1_HVT U1688 ( .A1(sram_raddr_a0[0]), .A2(n108), .A3(n359), .A4(n1590), 
        .A5(n1548), .Y(n_sram_raddr_a0[0]) );
  NAND2X0_HVT U1689 ( .A1(sram_raddr_a6[1]), .A2(sram_raddr_a6[0]), .Y(n1552)
         );
  OA21X1_HVT U1690 ( .A1(sram_raddr_a6[1]), .A2(sram_raddr_a6[0]), .A3(n1552), 
        .Y(n1836) );
  NAND2X0_HVT U1691 ( .A1(n94), .A2(n1836), .Y(n1714) );
  AO221X1_HVT U1692 ( .A1(n1742), .A2(n1557), .A3(n1742), .A4(sram_raddr_a0[0]), .A5(n368), .Y(n1551) );
  NAND3X0_HVT U1693 ( .A1(sram_raddr_a0[0]), .A2(n1590), .A3(n368), .Y(n1550)
         );
  NAND2X0_HVT U1694 ( .A1(sram_raddr_a3[1]), .A2(sram_raddr_a3[0]), .Y(n1554)
         );
  OA21X1_HVT U1695 ( .A1(sram_raddr_a3[1]), .A2(sram_raddr_a3[0]), .A3(n1554), 
        .Y(n1713) );
  NAND2X0_HVT U1696 ( .A1(n95), .A2(n1713), .Y(n1549) );
  NAND4X0_HVT U1697 ( .A1(n1714), .A2(n1551), .A3(n1550), .A4(n1549), .Y(
        n_sram_raddr_a0[1]) );
  NAND3X0_HVT U1698 ( .A1(sram_raddr_a0[2]), .A2(sram_raddr_a0[1]), .A3(
        sram_raddr_a0[0]), .Y(n1558) );
  AO21X1_HVT U1699 ( .A1(n1590), .A2(n1558), .A3(n109), .Y(n1556) );
  AND3X1_HVT U1700 ( .A1(sram_raddr_a0[1]), .A2(sram_raddr_a0[0]), .A3(n1590), 
        .Y(n1562) );
  AO22X1_HVT U1701 ( .A1(n1553), .A2(n337), .A3(n1552), .A4(sram_raddr_a6[2]), 
        .Y(n1837) );
  AO22X1_HVT U1702 ( .A1(sram_raddr_a3[2]), .A2(n1554), .A3(n164), .A4(n1559), 
        .Y(n1716) );
  AO22X1_HVT U1703 ( .A1(n458), .A2(n1837), .A3(n95), .A4(n1716), .Y(n1555) );
  AO221X1_HVT U1704 ( .A1(n1556), .A2(sram_raddr_a0[2]), .A3(n1556), .A4(n1562), .A5(n1555), .Y(n_sram_raddr_a0[2]) );
  NAND4X0_HVT U1705 ( .A1(sram_raddr_a3[2]), .A2(sram_raddr_a3[3]), .A3(
        sram_raddr_a3[1]), .A4(sram_raddr_a3[0]), .Y(n1561) );
  OA221X1_HVT U1706 ( .A1(sram_raddr_a3[3]), .A2(sram_raddr_a3[2]), .A3(
        sram_raddr_a3[3]), .A4(n1559), .A5(n1561), .Y(n1717) );
  AND3X1_HVT U1707 ( .A1(sram_raddr_a6[1]), .A2(sram_raddr_a6[0]), .A3(
        sram_raddr_a6[2]), .Y(n1560) );
  NAND4X0_HVT U1708 ( .A1(sram_raddr_a6[1]), .A2(sram_raddr_a6[0]), .A3(
        sram_raddr_a6[2]), .A4(sram_raddr_a6[3]), .Y(n1563) );
  OA21X1_HVT U1709 ( .A1(n1560), .A2(sram_raddr_a6[3]), .A3(n1563), .Y(n1838)
         );
  AND2X1_HVT U1710 ( .A1(n1827), .A2(n1838), .Y(n1719) );
  OR2X1_HVT U1711 ( .A1(n171), .A2(n1561), .Y(n1568) );
  AO21X1_HVT U1712 ( .A1(n171), .A2(n1561), .A3(n1567), .Y(n1720) );
  OA22X1_HVT U1713 ( .A1(n1566), .A2(n290), .A3(n115), .A4(n1720), .Y(n1564)
         );
  NAND4X0_HVT U1714 ( .A1(sram_raddr_a0[2]), .A2(sram_raddr_a0[3]), .A3(n1562), 
        .A4(n290), .Y(n1565) );
  AO22X1_HVT U1715 ( .A1(n1570), .A2(n383), .A3(n1563), .A4(sram_raddr_a6[4]), 
        .Y(n1842) );
  NAND2X0_HVT U1716 ( .A1(n94), .A2(n1842), .Y(n1722) );
  NAND3X0_HVT U1717 ( .A1(n1564), .A2(n1565), .A3(n1722), .Y(
        n_sram_raddr_a0[4]) );
  AND2X1_HVT U1718 ( .A1(n1566), .A2(n1565), .Y(n1574) );
  AND2X1_HVT U1719 ( .A1(sram_raddr_a3[5]), .A2(n1567), .Y(n1575) );
  AO21X1_HVT U1720 ( .A1(n289), .A2(n1568), .A3(n1575), .Y(n1725) );
  OA22X1_HVT U1721 ( .A1(n1574), .A2(n299), .A3(n116), .A4(n1725), .Y(n1572)
         );
  AND2X1_HVT U1722 ( .A1(sram_raddr_a0[1]), .A2(sram_raddr_a0[0]), .Y(n1569)
         );
  AND4X1_HVT U1723 ( .A1(sram_raddr_a0[4]), .A2(sram_raddr_a0[2]), .A3(
        sram_raddr_a0[3]), .A4(n1569), .Y(n1576) );
  NAND3X0_HVT U1724 ( .A1(n1576), .A2(n1590), .A3(n299), .Y(n1573) );
  AND2X1_HVT U1725 ( .A1(n1570), .A2(sram_raddr_a6[4]), .Y(n1571) );
  NAND2X0_HVT U1726 ( .A1(n1571), .A2(sram_raddr_a6[5]), .Y(n1577) );
  OA21X1_HVT U1727 ( .A1(n1571), .A2(sram_raddr_a6[5]), .A3(n1577), .Y(n1848)
         );
  NAND2X0_HVT U1728 ( .A1(n94), .A2(n1848), .Y(n1727) );
  NAND3X0_HVT U1729 ( .A1(n1572), .A2(n1573), .A3(n1727), .Y(
        n_sram_raddr_a0[5]) );
  AND2X1_HVT U1730 ( .A1(n1574), .A2(n1573), .Y(n1581) );
  NAND2X0_HVT U1731 ( .A1(sram_raddr_a3[6]), .A2(n1575), .Y(n1582) );
  OA22X1_HVT U1732 ( .A1(n1581), .A2(n329), .A3(n116), .A4(n1734), .Y(n1579)
         );
  AND2X1_HVT U1733 ( .A1(sram_raddr_a0[5]), .A2(n1576), .Y(n1585) );
  NAND3X0_HVT U1734 ( .A1(n1585), .A2(n1590), .A3(n329), .Y(n1580) );
  NAND2X0_HVT U1735 ( .A1(n1578), .A2(sram_raddr_a6[6]), .Y(n1583) );
  OA21X1_HVT U1736 ( .A1(n1578), .A2(sram_raddr_a6[6]), .A3(n1583), .Y(n1854)
         );
  NAND2X0_HVT U1737 ( .A1(n458), .A2(n1854), .Y(n1732) );
  NAND3X0_HVT U1738 ( .A1(n1579), .A2(n1580), .A3(n1732), .Y(
        n_sram_raddr_a0[6]) );
  AND2X1_HVT U1739 ( .A1(n1581), .A2(n1580), .Y(n1589) );
  AO21X1_HVT U1740 ( .A1(n271), .A2(n1582), .A3(n1594), .Y(n1740) );
  OA22X1_HVT U1741 ( .A1(n1589), .A2(n274), .A3(n116), .A4(n1740), .Y(n1587)
         );
  NAND2X0_HVT U1742 ( .A1(n1584), .A2(sram_raddr_a6[7]), .Y(n1592) );
  OA21X1_HVT U1743 ( .A1(n1584), .A2(sram_raddr_a6[7]), .A3(n1592), .Y(n1860)
         );
  NAND2X0_HVT U1744 ( .A1(n1827), .A2(n1860), .Y(n1744) );
  AND2X1_HVT U1745 ( .A1(sram_raddr_a0[6]), .A2(n1585), .Y(n1591) );
  NAND3X0_HVT U1746 ( .A1(n1591), .A2(n274), .A3(n1590), .Y(n1586) );
  NAND3X0_HVT U1747 ( .A1(n1587), .A2(n1744), .A3(n1586), .Y(
        n_sram_raddr_a0[7]) );
  NAND2X0_HVT U1748 ( .A1(n274), .A2(n1590), .Y(n1588) );
  NAND2X0_HVT U1749 ( .A1(n1589), .A2(n1588), .Y(n1602) );
  AND3X1_HVT U1750 ( .A1(sram_raddr_a0[7]), .A2(n1591), .A3(n1590), .Y(n1600)
         );
  NAND2X0_HVT U1751 ( .A1(n1593), .A2(sram_raddr_a6[8]), .Y(n1596) );
  OA21X1_HVT U1752 ( .A1(n1593), .A2(sram_raddr_a6[8]), .A3(n1596), .Y(n1867)
         );
  NAND2X0_HVT U1753 ( .A1(sram_raddr_a3[8]), .A2(n1594), .Y(n1598) );
  OA21X1_HVT U1754 ( .A1(sram_raddr_a3[8]), .A2(n1594), .A3(n1598), .Y(n1748)
         );
  AO22X1_HVT U1755 ( .A1(n458), .A2(n1867), .A3(n1945), .A4(n1748), .Y(n1595)
         );
  AO221X1_HVT U1756 ( .A1(sram_raddr_a0[8]), .A2(n1602), .A3(n375), .A4(n1600), 
        .A5(n1595), .Y(n_sram_raddr_a0[8]) );
  HADDX1_HVT U1757 ( .A0(sram_raddr_a6[9]), .B0(n1597), .SO(n1872) );
  AND2X1_HVT U1758 ( .A1(n458), .A2(n1872), .Y(n1754) );
  HADDX1_HVT U1759 ( .A0(sram_raddr_a3[9]), .B0(n1599), .SO(n1752) );
  HADDX1_HVT U1760 ( .A0(sram_raddr_a0[9]), .B0(sram_raddr_a0[8]), .SO(n1601)
         );
  NAND2X0_HVT U1761 ( .A1(n_addr_col_sel_cnt[1]), .A2(n178), .Y(n1876) );
  AO22X1_HVT U1762 ( .A1(n1827), .A2(n278), .A3(n1945), .A4(n212), .Y(n1603)
         );
  AO221X1_HVT U1763 ( .A1(sram_raddr_a1[0]), .A2(n1920), .A3(n362), .A4(n1640), 
        .A5(n1603), .Y(n_sram_raddr_a1[0]) );
  NAND2X0_HVT U1764 ( .A1(sram_raddr_a4[1]), .A2(sram_raddr_a4[0]), .Y(n1605)
         );
  AO21X1_HVT U1765 ( .A1(n358), .A2(n212), .A3(n1606), .Y(n1757) );
  AO22X1_HVT U1766 ( .A1(sram_raddr_a7[1]), .A2(n278), .A3(n214), .A4(
        sram_raddr_a7[0]), .Y(n1877) );
  NAND2X0_HVT U1767 ( .A1(n458), .A2(n1877), .Y(n1756) );
  AND2X1_HVT U1768 ( .A1(sram_raddr_a1[1]), .A2(sram_raddr_a1[0]), .Y(n1604)
         );
  NAND3X0_HVT U1769 ( .A1(sram_raddr_a1[2]), .A2(sram_raddr_a1[1]), .A3(
        sram_raddr_a1[0]), .Y(n1608) );
  AO21X1_HVT U1770 ( .A1(n1640), .A2(n1608), .A3(n1920), .Y(n1607) );
  AO22X1_HVT U1771 ( .A1(sram_raddr_a4[2]), .A2(n1605), .A3(n174), .A4(n1606), 
        .Y(n1759) );
  NAND3X0_HVT U1772 ( .A1(sram_raddr_a7[1]), .A2(sram_raddr_a7[0]), .A3(
        sram_raddr_a7[2]), .Y(n1609) );
  OA221X1_HVT U1773 ( .A1(sram_raddr_a7[2]), .A2(sram_raddr_a7[0]), .A3(
        sram_raddr_a7[2]), .A4(sram_raddr_a7[1]), .A5(n1609), .Y(n1882) );
  NAND4X0_HVT U1774 ( .A1(sram_raddr_a4[2]), .A2(sram_raddr_a4[3]), .A3(
        sram_raddr_a4[1]), .A4(sram_raddr_a4[0]), .Y(n1614) );
  OA221X1_HVT U1775 ( .A1(sram_raddr_a4[3]), .A2(sram_raddr_a4[2]), .A3(
        sram_raddr_a4[3]), .A4(n1606), .A5(n1614), .Y(n1762) );
  AOI22X1_HVT U1776 ( .A1(n95), .A2(n1762), .A3(sram_raddr_a1[3]), .A4(n1607), 
        .Y(n1612) );
  NAND3X0_HVT U1777 ( .A1(n1627), .A2(n1640), .A3(n173), .Y(n1611) );
  AO22X1_HVT U1778 ( .A1(n1610), .A2(n339), .A3(n1609), .A4(sram_raddr_a7[3]), 
        .Y(n1883) );
  NAND2X0_HVT U1779 ( .A1(n458), .A2(n1883), .Y(n1761) );
  NAND3X0_HVT U1780 ( .A1(n1612), .A2(n1611), .A3(n1761), .Y(
        n_sram_raddr_a1[3]) );
  OA221X1_HVT U1781 ( .A1(n1613), .A2(sram_raddr_a1[3]), .A3(n1613), .A4(n1627), .A5(n1895), .Y(n1619) );
  NAND2X0_HVT U1782 ( .A1(sram_raddr_a4[4]), .A2(n1615), .Y(n1622) );
  OA22X1_HVT U1783 ( .A1(n1619), .A2(n200), .A3(n116), .A4(n1764), .Y(n1617)
         );
  NAND4X0_HVT U1784 ( .A1(sram_raddr_a1[3]), .A2(n1627), .A3(n1640), .A4(n200), 
        .Y(n1618) );
  AND4X1_HVT U1785 ( .A1(sram_raddr_a7[1]), .A2(sram_raddr_a7[0]), .A3(
        sram_raddr_a7[2]), .A4(sram_raddr_a7[3]), .Y(n1616) );
  NAND2X0_HVT U1786 ( .A1(n1616), .A2(sram_raddr_a7[4]), .Y(n1621) );
  OA21X1_HVT U1787 ( .A1(n1616), .A2(sram_raddr_a7[4]), .A3(n1621), .Y(n1888)
         );
  NAND2X0_HVT U1788 ( .A1(n1827), .A2(n1888), .Y(n1767) );
  NAND3X0_HVT U1789 ( .A1(n1617), .A2(n1618), .A3(n1767), .Y(
        n_sram_raddr_a1[4]) );
  AND2X1_HVT U1790 ( .A1(n1619), .A2(n1618), .Y(n1625) );
  OR2X1_HVT U1791 ( .A1(n277), .A2(n1625), .Y(n1623) );
  AND3X1_HVT U1792 ( .A1(sram_raddr_a1[4]), .A2(sram_raddr_a1[3]), .A3(n1627), 
        .Y(n1620) );
  NAND3X0_HVT U1793 ( .A1(n1620), .A2(n1640), .A3(n277), .Y(n1624) );
  NOR2X0_HVT U1794 ( .A1(n1621), .A2(n313), .Y(n1628) );
  AO21X1_HVT U1795 ( .A1(n1621), .A2(n313), .A3(n1628), .Y(n1893) );
  NOR2X0_HVT U1796 ( .A1(n270), .A2(n1622), .Y(n1626) );
  AO21X1_HVT U1797 ( .A1(n270), .A2(n1622), .A3(n1626), .Y(n1769) );
  OA22X1_HVT U1798 ( .A1(n1924), .A2(n1893), .A3(n115), .A4(n1769), .Y(n1772)
         );
  NAND3X0_HVT U1799 ( .A1(n1623), .A2(n1624), .A3(n1772), .Y(
        n_sram_raddr_a1[5]) );
  AND2X1_HVT U1800 ( .A1(n1625), .A2(n1624), .Y(n1631) );
  NAND2X0_HVT U1801 ( .A1(sram_raddr_a4[6]), .A2(n1626), .Y(n1632) );
  OA22X1_HVT U1802 ( .A1(n1631), .A2(n294), .A3(n116), .A4(n1773), .Y(n1629)
         );
  AND4X1_HVT U1803 ( .A1(sram_raddr_a1[5]), .A2(sram_raddr_a1[4]), .A3(
        sram_raddr_a1[3]), .A4(n1627), .Y(n1635) );
  NAND3X0_HVT U1804 ( .A1(n1635), .A2(n1640), .A3(n294), .Y(n1630) );
  NAND2X0_HVT U1805 ( .A1(n1628), .A2(sram_raddr_a7[6]), .Y(n1633) );
  OA21X1_HVT U1806 ( .A1(n1628), .A2(sram_raddr_a7[6]), .A3(n1633), .Y(n1900)
         );
  NAND2X0_HVT U1807 ( .A1(n458), .A2(n1900), .Y(n1775) );
  NAND3X0_HVT U1808 ( .A1(n1629), .A2(n1630), .A3(n1775), .Y(
        n_sram_raddr_a1[6]) );
  AND2X1_HVT U1809 ( .A1(n1631), .A2(n1630), .Y(n1639) );
  AO21X1_HVT U1810 ( .A1(n272), .A2(n1632), .A3(n1644), .Y(n1777) );
  OA22X1_HVT U1811 ( .A1(n1639), .A2(n273), .A3(n115), .A4(n1777), .Y(n1637)
         );
  NAND2X0_HVT U1812 ( .A1(n1634), .A2(sram_raddr_a7[7]), .Y(n1642) );
  OA21X1_HVT U1813 ( .A1(n1634), .A2(sram_raddr_a7[7]), .A3(n1642), .Y(n1906)
         );
  NAND2X0_HVT U1814 ( .A1(n94), .A2(n1906), .Y(n1781) );
  AND2X1_HVT U1815 ( .A1(sram_raddr_a1[6]), .A2(n1635), .Y(n1641) );
  NAND3X0_HVT U1816 ( .A1(n1641), .A2(n273), .A3(n1640), .Y(n1636) );
  NAND3X0_HVT U1817 ( .A1(n1637), .A2(n1781), .A3(n1636), .Y(
        n_sram_raddr_a1[7]) );
  NAND2X0_HVT U1818 ( .A1(n273), .A2(n1640), .Y(n1638) );
  NAND2X0_HVT U1819 ( .A1(n1639), .A2(n1638), .Y(n1652) );
  AND3X1_HVT U1820 ( .A1(sram_raddr_a1[7]), .A2(n1641), .A3(n1640), .Y(n1650)
         );
  NAND2X0_HVT U1821 ( .A1(n1643), .A2(sram_raddr_a7[8]), .Y(n1646) );
  OA21X1_HVT U1822 ( .A1(n1643), .A2(sram_raddr_a7[8]), .A3(n1646), .Y(n1913)
         );
  NAND2X0_HVT U1823 ( .A1(sram_raddr_a4[8]), .A2(n1644), .Y(n1648) );
  OA21X1_HVT U1824 ( .A1(sram_raddr_a4[8]), .A2(n1644), .A3(n1648), .Y(n1784)
         );
  AO22X1_HVT U1825 ( .A1(n458), .A2(n1913), .A3(n1945), .A4(n1784), .Y(n1645)
         );
  AO221X1_HVT U1826 ( .A1(sram_raddr_a1[8]), .A2(n1652), .A3(n376), .A4(n1650), 
        .A5(n1645), .Y(n_sram_raddr_a1[8]) );
  HADDX1_HVT U1827 ( .A0(sram_raddr_a7[9]), .B0(n1647), .SO(n1919) );
  AND2X1_HVT U1828 ( .A1(n1827), .A2(n1919), .Y(n1790) );
  HADDX1_HVT U1829 ( .A0(sram_raddr_a4[9]), .B0(n1649), .SO(n1788) );
  HADDX1_HVT U1830 ( .A0(sram_raddr_a1[9]), .B0(sram_raddr_a1[8]), .SO(n1651)
         );
  OA22X1_HVT U1831 ( .A1(sram_raddr_a2[0]), .A2(n96), .A3(sram_raddr_a5[0]), 
        .A4(n115), .Y(n1925) );
  NAND4X0_HVT U1832 ( .A1(n1654), .A2(n1136), .A3(n1653), .A4(
        addr_col_sel_cnt[1]), .Y(n1923) );
  AO22X1_HVT U1833 ( .A1(sram_raddr_a2[0]), .A2(n1805), .A3(n361), .A4(n1923), 
        .Y(n1656) );
  NAND2X0_HVT U1834 ( .A1(n1827), .A2(n229), .Y(n1655) );
  NAND3X0_HVT U1835 ( .A1(n1925), .A2(n1656), .A3(n1655), .Y(
        n_sram_raddr_a2[0]) );
  NAND2X0_HVT U1836 ( .A1(sram_raddr_a2[1]), .A2(sram_raddr_a2[0]), .Y(n1662)
         );
  OA21X1_HVT U1837 ( .A1(sram_raddr_a2[1]), .A2(sram_raddr_a2[0]), .A3(n1662), 
        .Y(n1792) );
  NAND2X0_HVT U1838 ( .A1(n151), .A2(n1923), .Y(n1698) );
  AOI22X1_HVT U1839 ( .A1(sram_raddr_a2[1]), .A2(n1967), .A3(n1792), .A4(n1698), .Y(n1658) );
  NAND2X0_HVT U1840 ( .A1(sram_raddr_a5[1]), .A2(sram_raddr_a5[0]), .Y(n1665)
         );
  OA21X1_HVT U1841 ( .A1(sram_raddr_a5[1]), .A2(sram_raddr_a5[0]), .A3(n1665), 
        .Y(n1793) );
  NAND2X0_HVT U1842 ( .A1(n95), .A2(n1793), .Y(n1657) );
  NAND2X0_HVT U1843 ( .A1(sram_raddr_a8[1]), .A2(sram_raddr_a8[0]), .Y(n1660)
         );
  OA21X1_HVT U1844 ( .A1(sram_raddr_a8[1]), .A2(sram_raddr_a8[0]), .A3(n1660), 
        .Y(n1927) );
  NAND2X0_HVT U1845 ( .A1(n94), .A2(n1927), .Y(n1794) );
  NAND3X0_HVT U1846 ( .A1(n1658), .A2(n1657), .A3(n1794), .Y(
        n_sram_raddr_a2[1]) );
  NAND3X0_HVT U1847 ( .A1(sram_raddr_a5[2]), .A2(sram_raddr_a5[1]), .A3(
        sram_raddr_a5[0]), .Y(n1659) );
  NAND2X0_HVT U1848 ( .A1(n316), .A2(n1665), .Y(n1934) );
  NAND2X0_HVT U1849 ( .A1(n1659), .A2(n1934), .Y(n1932) );
  OA22X1_HVT U1850 ( .A1(n1805), .A2(n334), .A3(n115), .A4(n1932), .Y(n1664)
         );
  AO22X1_HVT U1851 ( .A1(n1661), .A2(n336), .A3(n1660), .A4(sram_raddr_a8[2]), 
        .Y(n1931) );
  NAND2X0_HVT U1852 ( .A1(n94), .A2(n1931), .Y(n1797) );
  AND3X1_HVT U1853 ( .A1(sram_raddr_a2[2]), .A2(sram_raddr_a2[1]), .A3(
        sram_raddr_a2[0]), .Y(n1796) );
  AND2X1_HVT U1854 ( .A1(n334), .A2(n1662), .Y(n1800) );
  OR3X1_HVT U1855 ( .A1(n1670), .A2(n1796), .A3(n1800), .Y(n1663) );
  NAND3X0_HVT U1856 ( .A1(n1664), .A2(n1797), .A3(n1663), .Y(
        n_sram_raddr_a2[2]) );
  OA21X1_HVT U1857 ( .A1(n1670), .A2(n1796), .A3(n1805), .Y(n1666) );
  NAND4X0_HVT U1858 ( .A1(sram_raddr_a5[3]), .A2(sram_raddr_a5[2]), .A3(
        sram_raddr_a5[1]), .A4(sram_raddr_a5[0]), .Y(n1672) );
  AO221X1_HVT U1859 ( .A1(n201), .A2(n316), .A3(n201), .A4(n1665), .A5(n1671), 
        .Y(n1799) );
  OA22X1_HVT U1860 ( .A1(n1666), .A2(n285), .A3(n116), .A4(n1799), .Y(n1669)
         );
  NAND3X0_HVT U1861 ( .A1(n1796), .A2(n1698), .A3(n285), .Y(n1668) );
  AND3X1_HVT U1862 ( .A1(sram_raddr_a8[1]), .A2(sram_raddr_a8[0]), .A3(
        sram_raddr_a8[2]), .Y(n1667) );
  NAND4X0_HVT U1863 ( .A1(sram_raddr_a8[1]), .A2(sram_raddr_a8[0]), .A3(
        sram_raddr_a8[2]), .A4(sram_raddr_a8[3]), .Y(n1673) );
  OA21X1_HVT U1864 ( .A1(n1667), .A2(sram_raddr_a8[3]), .A3(n1673), .Y(n1933)
         );
  NAND2X0_HVT U1865 ( .A1(n1827), .A2(n1933), .Y(n1801) );
  NAND3X0_HVT U1866 ( .A1(n1669), .A2(n1668), .A3(n1801), .Y(
        n_sram_raddr_a2[3]) );
  OA221X1_HVT U1867 ( .A1(n1670), .A2(sram_raddr_a2[3]), .A3(n1670), .A4(n1796), .A5(n1805), .Y(n1681) );
  AND2X1_HVT U1868 ( .A1(sram_raddr_a5[4]), .A2(n1671), .Y(n1676) );
  AO21X1_HVT U1869 ( .A1(n301), .A2(n1672), .A3(n1676), .Y(n1803) );
  OA22X1_HVT U1870 ( .A1(n1681), .A2(n283), .A3(n115), .A4(n1803), .Y(n1675)
         );
  NAND4X0_HVT U1871 ( .A1(sram_raddr_a2[3]), .A2(n1796), .A3(n1698), .A4(n283), 
        .Y(n1680) );
  NAND2X0_HVT U1872 ( .A1(n1674), .A2(sram_raddr_a8[4]), .Y(n1677) );
  OA21X1_HVT U1873 ( .A1(n1674), .A2(sram_raddr_a8[4]), .A3(n1677), .Y(n1938)
         );
  NAND2X0_HVT U1874 ( .A1(n94), .A2(n1938), .Y(n1807) );
  NAND3X0_HVT U1875 ( .A1(n1675), .A2(n1680), .A3(n1807), .Y(
        n_sram_raddr_a2[4]) );
  NAND2X0_HVT U1876 ( .A1(sram_raddr_a5[5]), .A2(n1676), .Y(n1687) );
  OA21X1_HVT U1877 ( .A1(sram_raddr_a5[5]), .A2(n1676), .A3(n1687), .Y(n1809)
         );
  NAND2X0_HVT U1878 ( .A1(n95), .A2(n1809), .Y(n1684) );
  NAND2X0_HVT U1879 ( .A1(n1678), .A2(sram_raddr_a8[5]), .Y(n1686) );
  OA21X1_HVT U1880 ( .A1(n1678), .A2(sram_raddr_a8[5]), .A3(n1686), .Y(n1944)
         );
  NAND2X0_HVT U1881 ( .A1(n94), .A2(n1944), .Y(n1813) );
  AND3X1_HVT U1882 ( .A1(sram_raddr_a2[4]), .A2(sram_raddr_a2[3]), .A3(n1796), 
        .Y(n1679) );
  NAND3X0_HVT U1883 ( .A1(n1679), .A2(n1698), .A3(n300), .Y(n1682) );
  NAND3X0_HVT U1884 ( .A1(n1681), .A2(n1682), .A3(n1680), .Y(n1688) );
  AO21X1_HVT U1885 ( .A1(n300), .A2(n1682), .A3(n1690), .Y(n1683) );
  NAND3X0_HVT U1886 ( .A1(n1684), .A2(n1813), .A3(n1683), .Y(
        n_sram_raddr_a2[5]) );
  AND4X1_HVT U1887 ( .A1(sram_raddr_a2[5]), .A2(sram_raddr_a2[4]), .A3(
        sram_raddr_a2[3]), .A4(n1796), .Y(n1685) );
  AND2X1_HVT U1888 ( .A1(n1685), .A2(n1698), .Y(n1691) );
  AO22X1_HVT U1889 ( .A1(n1692), .A2(n338), .A3(n1686), .A4(sram_raddr_a8[6]), 
        .Y(n1952) );
  AO22X1_HVT U1890 ( .A1(sram_raddr_a5[6]), .A2(n1687), .A3(n330), .A4(n1694), 
        .Y(n1816) );
  AO22X1_HVT U1891 ( .A1(n458), .A2(n1952), .A3(n95), .A4(n1816), .Y(n1818) );
  AO221X1_HVT U1892 ( .A1(sram_raddr_a2[6]), .A2(n1688), .A3(n323), .A4(n1691), 
        .A5(n1818), .Y(n_sram_raddr_a2[6]) );
  NAND2X0_HVT U1893 ( .A1(n1691), .A2(n323), .Y(n1689) );
  NAND2X0_HVT U1894 ( .A1(n1690), .A2(n1689), .Y(n1697) );
  AND2X1_HVT U1895 ( .A1(sram_raddr_a2[6]), .A2(n1691), .Y(n1699) );
  AND2X1_HVT U1896 ( .A1(n1692), .A2(sram_raddr_a8[6]), .Y(n1693) );
  NAND2X0_HVT U1897 ( .A1(n1693), .A2(sram_raddr_a8[7]), .Y(n1700) );
  OA21X1_HVT U1898 ( .A1(n1693), .A2(sram_raddr_a8[7]), .A3(n1700), .Y(n1956)
         );
  AND2X1_HVT U1899 ( .A1(sram_raddr_a5[6]), .A2(n1694), .Y(n1695) );
  NAND2X0_HVT U1900 ( .A1(sram_raddr_a5[7]), .A2(n1695), .Y(n1702) );
  OA21X1_HVT U1901 ( .A1(sram_raddr_a5[7]), .A2(n1695), .A3(n1702), .Y(n1822)
         );
  AO22X1_HVT U1902 ( .A1(n1827), .A2(n1956), .A3(n95), .A4(n1822), .Y(n1696)
         );
  AO221X1_HVT U1903 ( .A1(sram_raddr_a2[7]), .A2(n1697), .A3(n312), .A4(n1699), 
        .A5(n1696), .Y(n_sram_raddr_a2[7]) );
  AO21X1_HVT U1904 ( .A1(n312), .A2(n1698), .A3(n1697), .Y(n1711) );
  AND2X1_HVT U1905 ( .A1(sram_raddr_a2[7]), .A2(n1699), .Y(n1709) );
  NAND2X0_HVT U1906 ( .A1(n1701), .A2(sram_raddr_a8[8]), .Y(n1705) );
  OA21X1_HVT U1907 ( .A1(n1701), .A2(sram_raddr_a8[8]), .A3(n1705), .Y(n1962)
         );
  NAND2X0_HVT U1908 ( .A1(sram_raddr_a5[8]), .A2(n1703), .Y(n1707) );
  OA21X1_HVT U1909 ( .A1(sram_raddr_a5[8]), .A2(n1703), .A3(n1707), .Y(n1826)
         );
  AO22X1_HVT U1910 ( .A1(n458), .A2(n1962), .A3(n1945), .A4(n1826), .Y(n1704)
         );
  AO221X1_HVT U1911 ( .A1(sram_raddr_a2[8]), .A2(n1711), .A3(n326), .A4(n1709), 
        .A5(n1704), .Y(n_sram_raddr_a2[8]) );
  HADDX1_HVT U1912 ( .A0(sram_raddr_a8[9]), .B0(n1706), .SO(n1966) );
  AND2X1_HVT U1913 ( .A1(n458), .A2(n1966), .Y(n1833) );
  HADDX1_HVT U1914 ( .A0(sram_raddr_a5[9]), .B0(n1708), .SO(n1831) );
  HADDX1_HVT U1915 ( .A0(sram_raddr_a2[9]), .B0(sram_raddr_a2[8]), .SO(n1710)
         );
  NAND2X0_HVT U1916 ( .A1(n1853), .A2(n115), .Y(n1751) );
  AO22X1_HVT U1917 ( .A1(n458), .A2(n228), .A3(n1881), .A4(sram_raddr_a0[0]), 
        .Y(n1712) );
  AO221X1_HVT U1918 ( .A1(sram_raddr_a3[0]), .A2(n109), .A3(n360), .A4(n1751), 
        .A5(n1712), .Y(n_sram_raddr_a3[0]) );
  AOI22X1_HVT U1919 ( .A1(n1713), .A2(n1751), .A3(sram_raddr_a3[1]), .A4(n109), 
        .Y(n1715) );
  NAND2X0_HVT U1920 ( .A1(n1881), .A2(sram_raddr_a0[1]), .Y(n1835) );
  NAND3X0_HVT U1921 ( .A1(n1715), .A2(n1714), .A3(n1835), .Y(
        n_sram_raddr_a3[1]) );
  OA221X1_HVT U1922 ( .A1(sram_raddr_a0[2]), .A2(n172), .A3(n204), .A4(
        sram_raddr_a0[3]), .A5(n1881), .Y(n1841) );
  AO22X1_HVT U1923 ( .A1(n1717), .A2(n1751), .A3(sram_raddr_a3[3]), .A4(n108), 
        .Y(n1718) );
  OR3X1_HVT U1924 ( .A1(n1719), .A2(n1841), .A3(n1718), .Y(n_sram_raddr_a3[3])
         );
  OA22X1_HVT U1925 ( .A1(n1742), .A2(n171), .A3(n1741), .A4(n1720), .Y(n1724)
         );
  NAND3X0_HVT U1926 ( .A1(n290), .A2(n204), .A3(n172), .Y(n1726) );
  AND2X1_HVT U1927 ( .A1(n204), .A2(n172), .Y(n1721) );
  NAND3X0_HVT U1928 ( .A1(n1724), .A2(n1722), .A3(n1846), .Y(
        n_sram_raddr_a3[4]) );
  OA22X1_HVT U1929 ( .A1(n1742), .A2(n289), .A3(n1741), .A4(n1725), .Y(n1728)
         );
  NAND3X0_HVT U1930 ( .A1(n1728), .A2(n1727), .A3(n1851), .Y(
        n_sram_raddr_a3[5]) );
  NAND2X0_HVT U1931 ( .A1(n1729), .A2(n299), .Y(n1731) );
  OR2X1_HVT U1932 ( .A1(n1731), .A2(sram_raddr_a0[6]), .Y(n1743) );
  NAND2X0_HVT U1933 ( .A1(sram_raddr_a0[6]), .A2(n1731), .Y(n1733) );
  OA221X1_HVT U1934 ( .A1(n151), .A2(n1743), .A3(n151), .A4(n1733), .A5(n1732), 
        .Y(n1859) );
  OA22X1_HVT U1935 ( .A1(n1742), .A2(n310), .A3(n1741), .A4(n1734), .Y(n1736)
         );
  NAND2X0_HVT U1936 ( .A1(n1859), .A2(n1736), .Y(n_sram_raddr_a3[6]) );
  OA22X1_HVT U1937 ( .A1(n1742), .A2(n271), .A3(n1741), .A4(n1740), .Y(n1745)
         );
  NAND3X0_HVT U1938 ( .A1(n1745), .A2(n1744), .A3(n1864), .Y(
        n_sram_raddr_a3[7]) );
  NAND2X0_HVT U1939 ( .A1(n1746), .A2(n274), .Y(n1747) );
  OR2X1_HVT U1940 ( .A1(n1747), .A2(sram_raddr_a0[8]), .Y(n1749) );
  OA221X1_HVT U1941 ( .A1(n1750), .A2(sram_raddr_a0[8]), .A3(n1750), .A4(n1747), .A5(n1881), .Y(n1868) );
  OA221X1_HVT U1942 ( .A1(sram_raddr_a0[9]), .A2(n1750), .A3(n377), .A4(n1749), 
        .A5(n1881), .Y(n1874) );
  AO22X1_HVT U1943 ( .A1(n1752), .A2(n1751), .A3(sram_raddr_a3[9]), .A4(n109), 
        .Y(n1753) );
  OR3X1_HVT U1944 ( .A1(n1754), .A2(n1874), .A3(n1753), .Y(n_sram_raddr_a3[9])
         );
  NAND2X0_HVT U1945 ( .A1(n116), .A2(n1876), .Y(n1787) );
  AO22X1_HVT U1946 ( .A1(n1827), .A2(n278), .A3(n1881), .A4(sram_raddr_a1[0]), 
        .Y(n1755) );
  AO221X1_HVT U1947 ( .A1(sram_raddr_a4[0]), .A2(n1920), .A3(n212), .A4(n1787), 
        .A5(n1755), .Y(n_sram_raddr_a4[0]) );
  OA21X1_HVT U1948 ( .A1(n230), .A2(n151), .A3(n1756), .Y(n1880) );
  OA22X1_HVT U1949 ( .A1(n1778), .A2(n1757), .A3(n1895), .A4(n358), .Y(n1758)
         );
  NAND2X0_HVT U1950 ( .A1(n1880), .A2(n1758), .Y(n_sram_raddr_a4[1]) );
  AO221X1_HVT U1951 ( .A1(sram_raddr_a1[3]), .A2(n165), .A3(n173), .A4(
        sram_raddr_a1[2]), .A5(n151), .Y(n1760) );
  NAND2X0_HVT U1952 ( .A1(n1761), .A2(n1760), .Y(n1886) );
  AO22X1_HVT U1953 ( .A1(n1762), .A2(n1787), .A3(sram_raddr_a4[3]), .A4(n1920), 
        .Y(n1763) );
  OR2X1_HVT U1954 ( .A1(n1886), .A2(n1763), .Y(n_sram_raddr_a4[3]) );
  OA22X1_HVT U1955 ( .A1(n1895), .A2(n311), .A3(n1778), .A4(n1764), .Y(n1768)
         );
  NAND2X0_HVT U1956 ( .A1(n173), .A2(n165), .Y(n1765) );
  NAND3X0_HVT U1957 ( .A1(n1768), .A2(n1767), .A3(n1891), .Y(
        n_sram_raddr_a4[4]) );
  OA22X1_HVT U1958 ( .A1(n1895), .A2(n270), .A3(n1876), .A4(n1769), .Y(n1771)
         );
  NAND4X0_HVT U1959 ( .A1(n277), .A2(n200), .A3(n173), .A4(n165), .Y(n1774) );
  AND3X1_HVT U1960 ( .A1(n200), .A2(n173), .A3(n165), .Y(n1770) );
  AO221X1_HVT U1961 ( .A1(n1774), .A2(n1770), .A3(n1774), .A4(n277), .A5(n151), 
        .Y(n1898) );
  NAND3X0_HVT U1962 ( .A1(n1772), .A2(n1771), .A3(n1898), .Y(
        n_sram_raddr_a4[5]) );
  OA22X1_HVT U1963 ( .A1(n1895), .A2(n317), .A3(n1778), .A4(n1773), .Y(n1776)
         );
  NAND3X0_HVT U1964 ( .A1(n1776), .A2(n1775), .A3(n1904), .Y(
        n_sram_raddr_a4[6]) );
  OA22X1_HVT U1965 ( .A1(n1895), .A2(n272), .A3(n1778), .A4(n1777), .Y(n1782)
         );
  AND2X1_HVT U1966 ( .A1(n1779), .A2(n294), .Y(n1780) );
  NAND2X0_HVT U1967 ( .A1(n1780), .A2(n273), .Y(n1783) );
  NAND3X0_HVT U1968 ( .A1(n1782), .A2(n1781), .A3(n1909), .Y(
        n_sram_raddr_a4[7]) );
  OR2X1_HVT U1969 ( .A1(n1783), .A2(sram_raddr_a1[8]), .Y(n1785) );
  OA221X1_HVT U1970 ( .A1(n1786), .A2(sram_raddr_a1[8]), .A3(n1786), .A4(n1783), .A5(n1881), .Y(n1916) );
  OA221X1_HVT U1971 ( .A1(sram_raddr_a1[9]), .A2(n1786), .A3(n378), .A4(n1785), 
        .A5(n1881), .Y(n1922) );
  AO22X1_HVT U1972 ( .A1(n1788), .A2(n1787), .A3(sram_raddr_a4[9]), .A4(n1920), 
        .Y(n1789) );
  OR3X1_HVT U1973 ( .A1(n1790), .A2(n1922), .A3(n1789), .Y(n_sram_raddr_a4[9])
         );
  NAND2X0_HVT U1974 ( .A1(n115), .A2(n1923), .Y(n1830) );
  AO22X1_HVT U1975 ( .A1(n458), .A2(n229), .A3(n1881), .A4(n361), .Y(n1791) );
  AO221X1_HVT U1976 ( .A1(sram_raddr_a5[0]), .A2(n1967), .A3(n373), .A4(n1830), 
        .A5(n1791), .Y(n_sram_raddr_a5[0]) );
  AOI22X1_HVT U1977 ( .A1(n1881), .A2(n1792), .A3(n95), .A4(n1793), .Y(n1929)
         );
  AOI22X1_HVT U1978 ( .A1(n1957), .A2(n1793), .A3(sram_raddr_a5[1]), .A4(n1967), .Y(n1795) );
  NAND3X0_HVT U1979 ( .A1(n1929), .A2(n1795), .A3(n1794), .Y(
        n_sram_raddr_a5[1]) );
  OA22X1_HVT U1980 ( .A1(n1804), .A2(n1932), .A3(n1805), .A4(n316), .Y(n1798)
         );
  NAND3X0_HVT U1981 ( .A1(n1798), .A2(n1797), .A3(n1930), .Y(
        n_sram_raddr_a5[2]) );
  OA22X1_HVT U1982 ( .A1(n1804), .A2(n1799), .A3(n1805), .A4(n201), .Y(n1802)
         );
  NAND2X0_HVT U1983 ( .A1(n1800), .A2(n285), .Y(n1806) );
  AO221X1_HVT U1984 ( .A1(n1806), .A2(n1800), .A3(n1806), .A4(n285), .A5(n96), 
        .Y(n1936) );
  NAND3X0_HVT U1985 ( .A1(n1802), .A2(n1801), .A3(n1936), .Y(
        n_sram_raddr_a5[3]) );
  OA22X1_HVT U1986 ( .A1(n1805), .A2(n301), .A3(n1804), .A4(n1803), .Y(n1808)
         );
  NAND3X0_HVT U1987 ( .A1(n1808), .A2(n1807), .A3(n1942), .Y(
        n_sram_raddr_a5[4]) );
  AOI22X1_HVT U1988 ( .A1(n1809), .A2(n1830), .A3(sram_raddr_a5[5]), .A4(n1967), .Y(n1814) );
  AND2X1_HVT U1989 ( .A1(n1810), .A2(n283), .Y(n1812) );
  NAND2X0_HVT U1990 ( .A1(n1812), .A2(n300), .Y(n1815) );
  NAND3X0_HVT U1991 ( .A1(n1814), .A2(n1813), .A3(n1948), .Y(
        n_sram_raddr_a5[5]) );
  OR2X1_HVT U1992 ( .A1(n1815), .A2(sram_raddr_a2[6]), .Y(n1820) );
  OA221X1_HVT U1993 ( .A1(n1819), .A2(sram_raddr_a2[6]), .A3(n1819), .A4(n1815), .A5(n1881), .Y(n1953) );
  AO22X1_HVT U1994 ( .A1(n1957), .A2(n1816), .A3(sram_raddr_a5[6]), .A4(n1967), 
        .Y(n1817) );
  OR3X1_HVT U1995 ( .A1(n1953), .A2(n1818), .A3(n1817), .Y(n_sram_raddr_a5[6])
         );
  NAND2X0_HVT U1996 ( .A1(n1819), .A2(n312), .Y(n1825) );
  AO21X1_HVT U1997 ( .A1(sram_raddr_a2[7]), .A2(n1820), .A3(n1824), .Y(n1821)
         );
  AO22X1_HVT U1998 ( .A1(n458), .A2(n1956), .A3(n1881), .A4(n1821), .Y(n1959)
         );
  AO22X1_HVT U1999 ( .A1(n1822), .A2(n1830), .A3(sram_raddr_a5[7]), .A4(n1967), 
        .Y(n1823) );
  OR2X1_HVT U2000 ( .A1(n1959), .A2(n1823), .Y(n_sram_raddr_a5[7]) );
  NAND2X0_HVT U2001 ( .A1(n1824), .A2(n326), .Y(n1828) );
  OA221X1_HVT U2002 ( .A1(n1829), .A2(sram_raddr_a2[8]), .A3(n1829), .A4(n1825), .A5(n1881), .Y(n1963) );
  OA221X1_HVT U2003 ( .A1(sram_raddr_a2[9]), .A2(n1829), .A3(n379), .A4(n1828), 
        .A5(n1881), .Y(n1969) );
  AO22X1_HVT U2004 ( .A1(n1831), .A2(n1830), .A3(sram_raddr_a5[9]), .A4(n1967), 
        .Y(n1832) );
  OR3X1_HVT U2005 ( .A1(n1833), .A2(n1969), .A3(n1832), .Y(n_sram_raddr_a5[9])
         );
  NAND2X0_HVT U2006 ( .A1(n1924), .A2(n1853), .Y(n1871) );
  AO22X1_HVT U2007 ( .A1(n1881), .A2(sram_raddr_a0[0]), .A3(n95), .A4(
        sram_raddr_a3[0]), .Y(n1834) );
  AO221X1_HVT U2008 ( .A1(sram_raddr_a6[0]), .A2(n108), .A3(n228), .A4(n1871), 
        .A5(n1834), .Y(n_sram_raddr_a6[0]) );
  OA221X1_HVT U2009 ( .A1(sram_raddr_a3[2]), .A2(n205), .A3(n164), .A4(
        sram_raddr_a3[3]), .A5(n1945), .Y(n1840) );
  AO22X1_HVT U2010 ( .A1(sram_raddr_a6[3]), .A2(n108), .A3(n1838), .A4(n1871), 
        .Y(n1839) );
  OR3X1_HVT U2011 ( .A1(n1841), .A2(n1840), .A3(n1839), .Y(n_sram_raddr_a6[3])
         );
  AOI22X1_HVT U2012 ( .A1(sram_raddr_a6[4]), .A2(n108), .A3(n1842), .A4(n1871), 
        .Y(n1847) );
  NAND2X0_HVT U2013 ( .A1(n164), .A2(n205), .Y(n1843) );
  AO221X1_HVT U2014 ( .A1(sram_raddr_a3[4]), .A2(n1844), .A3(n171), .A4(n1843), 
        .A5(n116), .Y(n1845) );
  NAND3X0_HVT U2015 ( .A1(n1847), .A2(n1846), .A3(n1845), .Y(
        n_sram_raddr_a6[4]) );
  AOI22X1_HVT U2016 ( .A1(sram_raddr_a6[5]), .A2(n108), .A3(n1848), .A4(n1871), 
        .Y(n1852) );
  NAND4X0_HVT U2017 ( .A1(n289), .A2(n171), .A3(n164), .A4(n205), .Y(n1856) );
  AND3X1_HVT U2018 ( .A1(n171), .A2(n164), .A3(n205), .Y(n1849) );
  AO221X1_HVT U2019 ( .A1(n1856), .A2(n1849), .A3(n1856), .A4(n289), .A5(n116), 
        .Y(n1850) );
  NAND3X0_HVT U2020 ( .A1(n1852), .A2(n1851), .A3(n1850), .Y(
        n_sram_raddr_a6[5]) );
  AOI22X1_HVT U2021 ( .A1(sram_raddr_a6[6]), .A2(n108), .A3(n1855), .A4(n1854), 
        .Y(n1858) );
  AO221X1_HVT U2022 ( .A1(sram_raddr_a3[6]), .A2(n1861), .A3(n310), .A4(n1856), 
        .A5(n116), .Y(n1857) );
  NAND3X0_HVT U2023 ( .A1(n1859), .A2(n1858), .A3(n1857), .Y(
        n_sram_raddr_a6[6]) );
  AOI22X1_HVT U2024 ( .A1(sram_raddr_a6[7]), .A2(n109), .A3(n1860), .A4(n1871), 
        .Y(n1865) );
  AND2X1_HVT U2025 ( .A1(n1861), .A2(n310), .Y(n1862) );
  NAND2X0_HVT U2026 ( .A1(n1862), .A2(n271), .Y(n1866) );
  AO221X1_HVT U2027 ( .A1(n1866), .A2(n1862), .A3(n1866), .A4(n271), .A5(n115), 
        .Y(n1863) );
  NAND3X0_HVT U2028 ( .A1(n1865), .A2(n1864), .A3(n1863), .Y(
        n_sram_raddr_a6[7]) );
  HADDX1_HVT U2029 ( .A0(sram_raddr_a3[9]), .B0(n1869), .SO(n1870) );
  NAND2X0_HVT U2030 ( .A1(n1924), .A2(n1876), .Y(n1918) );
  AO22X1_HVT U2031 ( .A1(n1881), .A2(sram_raddr_a1[0]), .A3(n1945), .A4(
        sram_raddr_a4[0]), .Y(n1875) );
  AO221X1_HVT U2032 ( .A1(sram_raddr_a7[0]), .A2(n1920), .A3(n278), .A4(n1918), 
        .A5(n1875), .Y(n_sram_raddr_a7[0]) );
  OA22X1_HVT U2033 ( .A1(n1895), .A2(n214), .A3(n115), .A4(n358), .Y(n1879) );
  NAND2X0_HVT U2034 ( .A1(n1884), .A2(n1877), .Y(n1878) );
  NAND3X0_HVT U2035 ( .A1(n1880), .A2(n1879), .A3(n1878), .Y(
        n_sram_raddr_a7[1]) );
  OA221X1_HVT U2036 ( .A1(sram_raddr_a4[2]), .A2(n210), .A3(n174), .A4(
        sram_raddr_a4[3]), .A5(n95), .Y(n1887) );
  AO22X1_HVT U2037 ( .A1(sram_raddr_a7[3]), .A2(n1920), .A3(n1884), .A4(n1883), 
        .Y(n1885) );
  OR3X1_HVT U2038 ( .A1(n1887), .A2(n1886), .A3(n1885), .Y(n_sram_raddr_a7[3])
         );
  AOI22X1_HVT U2039 ( .A1(sram_raddr_a7[4]), .A2(n1920), .A3(n1888), .A4(n1918), .Y(n1892) );
  NAND3X0_HVT U2040 ( .A1(n311), .A2(n174), .A3(n210), .Y(n1896) );
  AND2X1_HVT U2041 ( .A1(n174), .A2(n210), .Y(n1889) );
  AO221X1_HVT U2042 ( .A1(n1896), .A2(n1889), .A3(n1896), .A4(n311), .A5(n116), 
        .Y(n1890) );
  NAND3X0_HVT U2043 ( .A1(n1892), .A2(n1891), .A3(n1890), .Y(
        n_sram_raddr_a7[4]) );
  OA22X1_HVT U2044 ( .A1(n1895), .A2(n313), .A3(n1894), .A4(n1893), .Y(n1899)
         );
  AO221X1_HVT U2045 ( .A1(sram_raddr_a4[5]), .A2(n1901), .A3(n270), .A4(n1896), 
        .A5(n115), .Y(n1897) );
  NAND3X0_HVT U2046 ( .A1(n1899), .A2(n1898), .A3(n1897), .Y(
        n_sram_raddr_a7[5]) );
  AOI22X1_HVT U2047 ( .A1(sram_raddr_a7[6]), .A2(n1920), .A3(n1900), .A4(n1918), .Y(n1905) );
  AND2X1_HVT U2048 ( .A1(n1901), .A2(n270), .Y(n1902) );
  NAND2X0_HVT U2049 ( .A1(n1902), .A2(n317), .Y(n1907) );
  AO221X1_HVT U2050 ( .A1(n1907), .A2(n1902), .A3(n1907), .A4(n317), .A5(n116), 
        .Y(n1903) );
  NAND3X0_HVT U2051 ( .A1(n1905), .A2(n1904), .A3(n1903), .Y(
        n_sram_raddr_a7[6]) );
  AOI22X1_HVT U2052 ( .A1(sram_raddr_a7[7]), .A2(n1920), .A3(n1906), .A4(n1918), .Y(n1910) );
  AO221X1_HVT U2053 ( .A1(sram_raddr_a4[7]), .A2(n1911), .A3(n272), .A4(n1907), 
        .A5(n115), .Y(n1908) );
  NAND3X0_HVT U2054 ( .A1(n1910), .A2(n1909), .A3(n1908), .Y(
        n_sram_raddr_a7[7]) );
  NAND2X0_HVT U2055 ( .A1(n1911), .A2(n272), .Y(n1912) );
  OA221X1_HVT U2056 ( .A1(n1917), .A2(sram_raddr_a4[8]), .A3(n1917), .A4(n1912), .A5(n95), .Y(n1915) );
  AO22X1_HVT U2057 ( .A1(sram_raddr_a7[8]), .A2(n1920), .A3(n1913), .A4(n1918), 
        .Y(n1914) );
  OR3X1_HVT U2058 ( .A1(n1916), .A2(n1915), .A3(n1914), .Y(n_sram_raddr_a7[8])
         );
  HADDX1_HVT U2059 ( .A0(sram_raddr_a4[9]), .B0(n1917), .SO(n1921) );
  AO221X1_HVT U2060 ( .A1(sram_raddr_a8[0]), .A2(n1967), .A3(n229), .A4(n1965), 
        .A5(n1926), .Y(n_sram_raddr_a8[0]) );
  AOI22X1_HVT U2061 ( .A1(sram_raddr_a8[1]), .A2(n1967), .A3(n1927), .A4(n1965), .Y(n1928) );
  NAND2X0_HVT U2062 ( .A1(n1929), .A2(n1928), .Y(n_sram_raddr_a8[1]) );
  AOI22X1_HVT U2063 ( .A1(sram_raddr_a8[3]), .A2(n1967), .A3(n1933), .A4(n1965), .Y(n1937) );
  AO221X1_HVT U2064 ( .A1(sram_raddr_a5[3]), .A2(n1939), .A3(n201), .A4(n1934), 
        .A5(n115), .Y(n1935) );
  NAND3X0_HVT U2065 ( .A1(n1937), .A2(n1936), .A3(n1935), .Y(
        n_sram_raddr_a8[3]) );
  AOI22X1_HVT U2066 ( .A1(sram_raddr_a8[4]), .A2(n1967), .A3(n1938), .A4(n1965), .Y(n1943) );
  AND2X1_HVT U2067 ( .A1(n1939), .A2(n201), .Y(n1940) );
  NAND2X0_HVT U2068 ( .A1(n1940), .A2(n301), .Y(n1946) );
  AO221X1_HVT U2069 ( .A1(n1946), .A2(n1940), .A3(n1946), .A4(n301), .A5(n115), 
        .Y(n1941) );
  NAND3X0_HVT U2070 ( .A1(n1943), .A2(n1942), .A3(n1941), .Y(
        n_sram_raddr_a8[4]) );
  AOI22X1_HVT U2071 ( .A1(sram_raddr_a8[5]), .A2(n1967), .A3(n1944), .A4(n1965), .Y(n1949) );
  AO221X1_HVT U2072 ( .A1(sram_raddr_a5[5]), .A2(n1950), .A3(n327), .A4(n1946), 
        .A5(n115), .Y(n1947) );
  NAND3X0_HVT U2073 ( .A1(n1949), .A2(n1948), .A3(n1947), .Y(
        n_sram_raddr_a8[5]) );
  NAND2X0_HVT U2074 ( .A1(n1950), .A2(n327), .Y(n1951) );
  OR2X1_HVT U2075 ( .A1(n1951), .A2(sram_raddr_a5[6]), .Y(n1954) );
  OR2X1_HVT U2076 ( .A1(n1954), .A2(sram_raddr_a5[7]), .Y(n1961) );
  OA221X1_HVT U2077 ( .A1(n1955), .A2(sram_raddr_a5[7]), .A3(n1955), .A4(n1954), .A5(n95), .Y(n1960) );
  AO22X1_HVT U2078 ( .A1(sram_raddr_a8[7]), .A2(n1967), .A3(n1957), .A4(n1956), 
        .Y(n1958) );
  OR3X1_HVT U2079 ( .A1(n1960), .A2(n1959), .A3(n1958), .Y(n_sram_raddr_a8[7])
         );
  HADDX1_HVT U2080 ( .A0(sram_raddr_a5[9]), .B0(n1964), .SO(n1968) );
  AND2X1_HVT U2081 ( .A1(n1970), .A2(addr_row_sel_cnt[1]), .Y(n487) );
  OA221X1_HVT U2082 ( .A1(n1979), .A2(n1971), .A3(n1979), .A4(n1977), .A5(
        n1975), .Y(n462) );
  AO22X1_HVT U2083 ( .A1(n1974), .A2(n1973), .A3(n1977), .A4(n1972), .Y(n460)
         );
  OA221X1_HVT U2084 ( .A1(n1979), .A2(n1978), .A3(n1979), .A4(n1977), .A5(
        n1976), .Y(n459) );
endmodule


module data_reg ( clk, srstn, mode, box_sel, sram_rdata_a0, sram_rdata_a1, 
        sram_rdata_a2, sram_rdata_a3, sram_rdata_a4, sram_rdata_a5, 
        sram_rdata_a6, sram_rdata_a7, sram_rdata_a8, sram_rdata_b0, 
        sram_rdata_b1, sram_rdata_b2, sram_rdata_b3, sram_rdata_b4, 
        sram_rdata_b5, sram_rdata_b6, sram_rdata_b7, sram_rdata_b8, 
        sram_rdata_weight, conv1_weight, weight, src_window );
  input [1:0] mode;
  input [3:0] box_sel;
  input [31:0] sram_rdata_a0;
  input [31:0] sram_rdata_a1;
  input [31:0] sram_rdata_a2;
  input [31:0] sram_rdata_a3;
  input [31:0] sram_rdata_a4;
  input [31:0] sram_rdata_a5;
  input [31:0] sram_rdata_a6;
  input [31:0] sram_rdata_a7;
  input [31:0] sram_rdata_a8;
  input [31:0] sram_rdata_b0;
  input [31:0] sram_rdata_b1;
  input [31:0] sram_rdata_b2;
  input [31:0] sram_rdata_b3;
  input [31:0] sram_rdata_b4;
  input [31:0] sram_rdata_b5;
  input [31:0] sram_rdata_b6;
  input [31:0] sram_rdata_b7;
  input [31:0] sram_rdata_b8;
  input [99:0] sram_rdata_weight;
  output [99:0] conv1_weight;
  output [99:0] weight;
  output [287:0] src_window;
  input clk, srstn;
  wire   N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52,
         N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66,
         N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80,
         N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94,
         N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139,
         N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161,
         N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172,
         N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183,
         N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194,
         N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205,
         N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216,
         N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227,
         N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238,
         N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249,
         N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260,
         N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271,
         N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282,
         N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293,
         N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304,
         N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315,
         N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326,
         N346, n777, n2, n3, n5, n6, n8, n9, n11, n12, n14, n15, n17, n18, n20,
         n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n3900, n4000, n4100, n4200, n4300, n4400, n4500, n4600,
         n4700, n4800, n4900, n5000, n5100, n5200, n5300, n5400, n5500, n5600,
         n5700, n5800, n5900, n6000, n6100, n6200, n6300, n6400, n6500, n6600,
         n6700, n6800, n6900, n7000, n7100, n7200, n7300, n7400, n7500, n7600,
         n7700, n7800, n7900, n8000, n8100, n8200, n8300, n8400, n8500, n8600,
         n8700, n8800, n8900, n9000, n9100, n9200, n9300, n9400, n9500, n9600,
         n9700, n9800, n9900, n10000, n10100, n10200, n10300, n10400, n10500,
         n10600, n10700, n10800, n10900, n11000, n11100, n11200, n11300,
         n11400, n11500, n11600, n11700, n11800, n11900, n12000, n12100,
         n12200, n12300, n12400, n12500, n12600, n12700, n12800, n12900,
         n13000, n13100, n13200, n13300, n13400, n13500, n13600, n1370, n1380,
         n1390, n1400, n1410, n1420, n1430, n1440, n1450, n1460, n1470, n1480,
         n1490, n1500, n1510, n1520, n1530, n1540, n1550, n1560, n1570, n1580,
         n1590, n1600, n1610, n1620, n1630, n1640, n1650, n1660, n1670, n1680,
         n1690, n1700, n1710, n1720, n1730, n1740, n1750, n1760, n1770, n1780,
         n1790, n1800, n1810, n1820, n1830, n1840, n1850, n1860, n1870, n1880,
         n1890, n1900, n1910, n1920, n1930, n1940, n1950, n1960, n1970, n1980,
         n1990, n2000, n2010, n2020, n2030, n2040, n2050, n2060, n2070, n2080,
         n2090, n2100, n2110, n2120, n2130, n2140, n2150, n2160, n2170, n2180,
         n2190, n2200, n2210, n2220, n2230, n2240, n2250, n2260, n2270, n2280,
         n2290, n2300, n2310, n2320, n2330, n2340, n2350, n2360, n2370, n2380,
         n2390, n2400, n2410, n2420, n2430, n2440, n2450, n2460, n2470, n2480,
         n2490, n2500, n2510, n2520, n2530, n2540, n2550, n2560, n2570, n2580,
         n2590, n2600, n2610, n2620, n2630, n2640, n2650, n2660, n2670, n2680,
         n2690, n2700, n2710, n2720, n2730, n2740, n2750, n2760, n2770, n2780,
         n2790, n2800, n2810, n2820, n2830, n2840, n2850, n2860, n2870, n2880,
         n2890, n2900, n2910, n2920, n2930, n2940, n2950, n2960, n2970, n2980,
         n2990, n3000, n3010, n3020, n3030, n3040, n3050, n3060, n3070, n3080,
         n3090, n3100, n3110, n3120, n3130, n3140, n3150, n3160, n3170, n3180,
         n3190, n3200, n3210, n3220, n3230, n3240, n3250, n3260, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n3460, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n3901, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n4001, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n4101, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n4201, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n4301, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n4401, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n4501, n451, n452, n453, n454, n455, n456, n457, n458, n459, n4601,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n4701, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n4801, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n4901, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n5001, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n5101, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n5201, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n5301, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n5401, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n5501, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n5601, n561, n562, n563, n564, n565, n566, n567, n568, n569, n5701,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n5801, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n5901, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n6001, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n6101, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n6201, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n6301, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n6401, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n6501, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n6601, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n6701, n671, n672, n673, n674, n675, n676, n677, n678, n679, n6801,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n6901, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n7001, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n7101, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n7201, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n7301, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n7401, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n7501, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n7601, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n7701, n771, n772, n773, n774, n775, n778, n779, n7801, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n7901, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n8001, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n8101, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n8201, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n8301, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n8401, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n8501, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n8601, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n8701, n871, n872, n873, n874, n875, n876, n877, n878, n879, n8801,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n8901, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n9001, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n9101, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n9201, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n9301, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n9401, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n9501, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n9601, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n9701, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n9801, n981, n982, n983, n984, n985, n986, n987, n988, n989, n9901,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n10001, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n10101, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n10201, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n10301, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n10401, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n10501, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n10601, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n10701, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n10801, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n10901, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n11001, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n11101, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n11201, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n11301, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n11401, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n11501, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n11601, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n11701, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n11801, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n11901, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n12001, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n12101, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n12201, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n12301, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n12401, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n12501, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n12601, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n12701, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n12801, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n12901, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n13001, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n13101, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n13201, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n13301, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n13401, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n13501, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n13601, n1361,
         n1362;
  wire   [287:0] n_src_aox;
  wire   [31:0] sram_rdata_0;
  wire   [31:0] sram_rdata_1;
  wire   [31:0] sram_rdata_2;
  wire   [31:0] sram_rdata_3;
  wire   [31:0] sram_rdata_4;
  wire   [31:0] sram_rdata_5;
  wire   [31:0] sram_rdata_6;
  wire   [31:0] sram_rdata_7;
  wire   [31:0] sram_rdata_8;

  DFFSSRX1_HVT src_aox_reg_0__7_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[287]), .CLK(clk), .Q(src_window[287]) );
  DFFSSRX1_HVT src_aox_reg_0__6_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[286]), .CLK(clk), .Q(src_window[286]) );
  DFFSSRX1_HVT src_aox_reg_0__5_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[285]), .CLK(clk), .Q(src_window[285]) );
  DFFSSRX1_HVT src_aox_reg_0__4_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[284]), .CLK(clk), .Q(src_window[284]) );
  DFFSSRX1_HVT src_aox_reg_0__3_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[283]), .CLK(clk), .Q(src_window[283]) );
  DFFSSRX1_HVT src_aox_reg_0__2_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[282]), .CLK(clk), .Q(src_window[282]) );
  DFFSSRX1_HVT src_aox_reg_0__1_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[281]), .CLK(clk), .Q(src_window[281]) );
  DFFSSRX1_HVT src_aox_reg_0__0_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[280]), .CLK(clk), .Q(src_window[280]) );
  DFFSSRX1_HVT src_aox_reg_1__7_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[279]), .CLK(clk), .Q(src_window[279]) );
  DFFSSRX1_HVT src_aox_reg_1__6_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[278]), .CLK(clk), .Q(src_window[278]) );
  DFFSSRX1_HVT src_aox_reg_1__5_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[277]), .CLK(clk), .Q(src_window[277]) );
  DFFSSRX1_HVT src_aox_reg_1__4_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[276]), .CLK(clk), .Q(src_window[276]) );
  DFFSSRX1_HVT src_aox_reg_1__3_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[275]), .CLK(clk), .Q(src_window[275]) );
  DFFSSRX1_HVT src_aox_reg_1__2_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[274]), .CLK(clk), .Q(src_window[274]) );
  DFFSSRX1_HVT src_aox_reg_1__1_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[273]), .CLK(clk), .Q(src_window[273]) );
  DFFSSRX1_HVT src_aox_reg_1__0_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[272]), .CLK(clk), .Q(src_window[272]) );
  DFFSSRX1_HVT src_aox_reg_2__7_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[271]), .CLK(clk), .Q(src_window[271]) );
  DFFSSRX1_HVT src_aox_reg_2__6_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[270]), .CLK(clk), .Q(src_window[270]) );
  DFFSSRX1_HVT src_aox_reg_2__5_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[269]), .CLK(clk), .Q(src_window[269]) );
  DFFSSRX1_HVT src_aox_reg_2__4_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[268]), .CLK(clk), .Q(src_window[268]) );
  DFFSSRX1_HVT src_aox_reg_2__3_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[267]), .CLK(clk), .Q(src_window[267]) );
  DFFSSRX1_HVT src_aox_reg_2__2_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[266]), .CLK(clk), .Q(src_window[266]) );
  DFFSSRX1_HVT src_aox_reg_2__1_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[265]), .CLK(clk), .Q(src_window[265]) );
  DFFSSRX1_HVT src_aox_reg_2__0_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[264]), .CLK(clk), .Q(src_window[264]) );
  DFFSSRX1_HVT src_aox_reg_3__7_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[263]), .CLK(clk), .Q(src_window[263]) );
  DFFSSRX1_HVT src_aox_reg_3__6_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[262]), .CLK(clk), .Q(src_window[262]) );
  DFFSSRX1_HVT src_aox_reg_3__5_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[261]), .CLK(clk), .Q(src_window[261]) );
  DFFSSRX1_HVT src_aox_reg_3__4_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[260]), .CLK(clk), .Q(src_window[260]) );
  DFFSSRX1_HVT src_aox_reg_3__3_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[259]), .CLK(clk), .Q(src_window[259]) );
  DFFSSRX1_HVT src_aox_reg_3__2_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[258]), .CLK(clk), .Q(src_window[258]) );
  DFFSSRX1_HVT src_aox_reg_3__1_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[257]), .CLK(clk), .Q(src_window[257]) );
  DFFSSRX1_HVT src_aox_reg_3__0_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[256]), .CLK(clk), .Q(src_window[256]) );
  DFFSSRX1_HVT src_aox_reg_4__7_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[255]), .CLK(clk), .Q(src_window[255]) );
  DFFSSRX1_HVT src_aox_reg_4__6_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[254]), .CLK(clk), .Q(src_window[254]) );
  DFFSSRX1_HVT src_aox_reg_4__5_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[253]), .CLK(clk), .Q(src_window[253]) );
  DFFSSRX1_HVT src_aox_reg_4__4_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[252]), .CLK(clk), .Q(src_window[252]) );
  DFFSSRX1_HVT src_aox_reg_4__3_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[251]), .CLK(clk), .Q(src_window[251]) );
  DFFSSRX1_HVT src_aox_reg_4__2_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[250]), .CLK(clk), .Q(src_window[250]) );
  DFFSSRX1_HVT src_aox_reg_4__1_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[249]), .CLK(clk), .Q(src_window[249]) );
  DFFSSRX1_HVT src_aox_reg_4__0_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[248]), .CLK(clk), .Q(src_window[248]) );
  DFFSSRX1_HVT src_aox_reg_5__7_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[247]), .CLK(clk), .Q(src_window[247]) );
  DFFSSRX1_HVT src_aox_reg_5__6_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[246]), .CLK(clk), .Q(src_window[246]) );
  DFFSSRX1_HVT src_aox_reg_5__5_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[245]), .CLK(clk), .Q(src_window[245]) );
  DFFSSRX1_HVT src_aox_reg_5__4_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[244]), .CLK(clk), .Q(src_window[244]) );
  DFFSSRX1_HVT src_aox_reg_5__3_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[243]), .CLK(clk), .Q(src_window[243]) );
  DFFSSRX1_HVT src_aox_reg_5__2_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[242]), .CLK(clk), .Q(src_window[242]) );
  DFFSSRX1_HVT src_aox_reg_5__1_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[241]), .CLK(clk), .Q(src_window[241]) );
  DFFSSRX1_HVT src_aox_reg_5__0_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[240]), .CLK(clk), .Q(src_window[240]) );
  DFFSSRX1_HVT src_aox_reg_6__7_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[239]), .CLK(clk), .Q(src_window[239]) );
  DFFSSRX1_HVT src_aox_reg_6__6_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[238]), .CLK(clk), .Q(src_window[238]) );
  DFFSSRX1_HVT src_aox_reg_6__5_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[237]), .CLK(clk), .Q(src_window[237]) );
  DFFSSRX1_HVT src_aox_reg_6__4_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[236]), .CLK(clk), .Q(src_window[236]) );
  DFFSSRX1_HVT src_aox_reg_6__3_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[235]), .CLK(clk), .Q(src_window[235]) );
  DFFSSRX1_HVT src_aox_reg_6__2_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[234]), .CLK(clk), .Q(src_window[234]) );
  DFFSSRX1_HVT src_aox_reg_6__1_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[233]), .CLK(clk), .Q(src_window[233]) );
  DFFSSRX1_HVT src_aox_reg_6__0_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[232]), .CLK(clk), .Q(src_window[232]) );
  DFFSSRX1_HVT src_aox_reg_7__7_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[231]), .CLK(clk), .Q(src_window[231]) );
  DFFSSRX1_HVT src_aox_reg_7__6_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[230]), .CLK(clk), .Q(src_window[230]) );
  DFFSSRX1_HVT src_aox_reg_7__5_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[229]), .CLK(clk), .Q(src_window[229]) );
  DFFSSRX1_HVT src_aox_reg_7__4_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[228]), .CLK(clk), .Q(src_window[228]) );
  DFFSSRX1_HVT src_aox_reg_7__3_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[227]), .CLK(clk), .Q(src_window[227]) );
  DFFSSRX1_HVT src_aox_reg_7__2_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[226]), .CLK(clk), .Q(src_window[226]) );
  DFFSSRX1_HVT src_aox_reg_7__1_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[225]), .CLK(clk), .Q(src_window[225]) );
  DFFSSRX1_HVT src_aox_reg_7__0_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[224]), .CLK(clk), .Q(src_window[224]) );
  DFFSSRX1_HVT src_aox_reg_8__7_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[223]), .CLK(clk), .Q(src_window[223]) );
  DFFSSRX1_HVT src_aox_reg_8__6_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[222]), .CLK(clk), .Q(src_window[222]) );
  DFFSSRX1_HVT src_aox_reg_8__5_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[221]), .CLK(clk), .Q(src_window[221]) );
  DFFSSRX1_HVT src_aox_reg_8__4_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[220]), .CLK(clk), .Q(src_window[220]) );
  DFFSSRX1_HVT src_aox_reg_8__3_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[219]), .CLK(clk), .Q(src_window[219]) );
  DFFSSRX1_HVT src_aox_reg_8__2_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[218]), .CLK(clk), .Q(src_window[218]) );
  DFFSSRX1_HVT src_aox_reg_8__1_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[217]), .CLK(clk), .Q(src_window[217]) );
  DFFSSRX1_HVT src_aox_reg_8__0_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[216]), .CLK(clk), .Q(src_window[216]) );
  DFFSSRX1_HVT src_aox_reg_9__7_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[215]), .CLK(clk), .Q(src_window[215]) );
  DFFSSRX1_HVT src_aox_reg_9__6_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[214]), .CLK(clk), .Q(src_window[214]) );
  DFFSSRX1_HVT src_aox_reg_9__5_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[213]), .CLK(clk), .Q(src_window[213]) );
  DFFSSRX1_HVT src_aox_reg_9__4_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[212]), .CLK(clk), .Q(src_window[212]) );
  DFFSSRX1_HVT src_aox_reg_9__3_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[211]), .CLK(clk), .Q(src_window[211]) );
  DFFSSRX1_HVT src_aox_reg_9__2_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[210]), .CLK(clk), .Q(src_window[210]) );
  DFFSSRX1_HVT src_aox_reg_9__1_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[209]), .CLK(clk), .Q(src_window[209]) );
  DFFSSRX1_HVT src_aox_reg_9__0_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[208]), .CLK(clk), .Q(src_window[208]) );
  DFFSSRX1_HVT src_aox_reg_10__7_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[207]), .CLK(clk), .Q(src_window[207]) );
  DFFSSRX1_HVT src_aox_reg_10__6_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[206]), .CLK(clk), .Q(src_window[206]) );
  DFFSSRX1_HVT src_aox_reg_10__5_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[205]), .CLK(clk), .Q(src_window[205]) );
  DFFSSRX1_HVT src_aox_reg_10__4_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[204]), .CLK(clk), .Q(src_window[204]) );
  DFFSSRX1_HVT src_aox_reg_10__3_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[203]), .CLK(clk), .Q(src_window[203]) );
  DFFSSRX1_HVT src_aox_reg_10__2_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[202]), .CLK(clk), .Q(src_window[202]) );
  DFFSSRX1_HVT src_aox_reg_10__1_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[201]), .CLK(clk), .Q(src_window[201]) );
  DFFSSRX1_HVT src_aox_reg_10__0_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[200]), .CLK(clk), .Q(src_window[200]) );
  DFFSSRX1_HVT src_aox_reg_11__7_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[199]), .CLK(clk), .Q(src_window[199]) );
  DFFSSRX1_HVT src_aox_reg_11__6_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[198]), .CLK(clk), .Q(src_window[198]) );
  DFFSSRX1_HVT src_aox_reg_11__5_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[197]), .CLK(clk), .Q(src_window[197]) );
  DFFSSRX1_HVT src_aox_reg_11__4_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[196]), .CLK(clk), .Q(src_window[196]) );
  DFFSSRX1_HVT src_aox_reg_11__3_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[195]), .CLK(clk), .Q(src_window[195]) );
  DFFSSRX1_HVT src_aox_reg_11__2_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[194]), .CLK(clk), .Q(src_window[194]) );
  DFFSSRX1_HVT src_aox_reg_11__1_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[193]), .CLK(clk), .Q(src_window[193]) );
  DFFSSRX1_HVT src_aox_reg_11__0_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[192]), .CLK(clk), .Q(src_window[192]) );
  DFFSSRX1_HVT src_aox_reg_12__7_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[191]), .CLK(clk), .Q(src_window[191]) );
  DFFSSRX1_HVT src_aox_reg_12__6_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[190]), .CLK(clk), .Q(src_window[190]) );
  DFFSSRX1_HVT src_aox_reg_12__5_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[189]), .CLK(clk), .Q(src_window[189]) );
  DFFSSRX1_HVT src_aox_reg_12__4_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[188]), .CLK(clk), .Q(src_window[188]) );
  DFFSSRX1_HVT src_aox_reg_12__3_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[187]), .CLK(clk), .Q(src_window[187]) );
  DFFSSRX1_HVT src_aox_reg_12__2_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[186]), .CLK(clk), .Q(src_window[186]) );
  DFFSSRX1_HVT src_aox_reg_12__1_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[185]), .CLK(clk), .Q(src_window[185]) );
  DFFSSRX1_HVT src_aox_reg_12__0_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[184]), .CLK(clk), .Q(src_window[184]) );
  DFFSSRX1_HVT src_aox_reg_13__7_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[183]), .CLK(clk), .Q(src_window[183]) );
  DFFSSRX1_HVT src_aox_reg_13__6_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[182]), .CLK(clk), .Q(src_window[182]) );
  DFFSSRX1_HVT src_aox_reg_13__5_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[181]), .CLK(clk), .Q(src_window[181]) );
  DFFSSRX1_HVT src_aox_reg_13__4_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[180]), .CLK(clk), .Q(src_window[180]) );
  DFFSSRX1_HVT src_aox_reg_13__3_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[179]), .CLK(clk), .Q(src_window[179]) );
  DFFSSRX1_HVT src_aox_reg_13__2_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[178]), .CLK(clk), .Q(src_window[178]) );
  DFFSSRX1_HVT src_aox_reg_13__1_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[177]), .CLK(clk), .Q(src_window[177]) );
  DFFSSRX1_HVT src_aox_reg_13__0_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[176]), .CLK(clk), .Q(src_window[176]) );
  DFFSSRX1_HVT src_aox_reg_14__7_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[175]), .CLK(clk), .Q(src_window[175]) );
  DFFSSRX1_HVT src_aox_reg_14__6_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[174]), .CLK(clk), .Q(src_window[174]) );
  DFFSSRX1_HVT src_aox_reg_14__5_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[173]), .CLK(clk), .Q(src_window[173]) );
  DFFSSRX1_HVT src_aox_reg_14__4_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[172]), .CLK(clk), .Q(src_window[172]) );
  DFFSSRX1_HVT src_aox_reg_14__3_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[171]), .CLK(clk), .Q(src_window[171]) );
  DFFSSRX1_HVT src_aox_reg_14__2_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[170]), .CLK(clk), .Q(src_window[170]) );
  DFFSSRX1_HVT src_aox_reg_14__1_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[169]), .CLK(clk), .Q(src_window[169]) );
  DFFSSRX1_HVT src_aox_reg_14__0_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[168]), .CLK(clk), .Q(src_window[168]) );
  DFFSSRX1_HVT src_aox_reg_15__7_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[167]), .CLK(clk), .Q(src_window[167]) );
  DFFSSRX1_HVT src_aox_reg_15__6_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[166]), .CLK(clk), .Q(src_window[166]) );
  DFFSSRX1_HVT src_aox_reg_15__5_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[165]), .CLK(clk), .Q(src_window[165]) );
  DFFSSRX1_HVT src_aox_reg_15__4_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[164]), .CLK(clk), .Q(src_window[164]) );
  DFFSSRX1_HVT src_aox_reg_15__3_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[163]), .CLK(clk), .Q(src_window[163]) );
  DFFSSRX1_HVT src_aox_reg_15__2_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[162]), .CLK(clk), .Q(src_window[162]) );
  DFFSSRX1_HVT src_aox_reg_15__1_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[161]), .CLK(clk), .Q(src_window[161]) );
  DFFSSRX1_HVT src_aox_reg_15__0_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[160]), .CLK(clk), .Q(src_window[160]) );
  DFFSSRX1_HVT src_aox_reg_16__7_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[159]), .CLK(clk), .Q(src_window[159]) );
  DFFSSRX1_HVT src_aox_reg_16__6_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[158]), .CLK(clk), .Q(src_window[158]) );
  DFFSSRX1_HVT src_aox_reg_16__5_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[157]), .CLK(clk), .Q(src_window[157]) );
  DFFSSRX1_HVT src_aox_reg_16__4_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[156]), .CLK(clk), .Q(src_window[156]) );
  DFFSSRX1_HVT src_aox_reg_16__3_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[155]), .CLK(clk), .Q(src_window[155]) );
  DFFSSRX1_HVT src_aox_reg_16__2_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[154]), .CLK(clk), .Q(src_window[154]) );
  DFFSSRX1_HVT src_aox_reg_16__1_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[153]), .CLK(clk), .Q(src_window[153]) );
  DFFSSRX1_HVT src_aox_reg_16__0_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[152]), .CLK(clk), .Q(src_window[152]) );
  DFFSSRX1_HVT src_aox_reg_17__7_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[151]), .CLK(clk), .Q(src_window[151]) );
  DFFSSRX1_HVT src_aox_reg_17__6_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[150]), .CLK(clk), .Q(src_window[150]) );
  DFFSSRX1_HVT src_aox_reg_17__5_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[149]), .CLK(clk), .Q(src_window[149]) );
  DFFSSRX1_HVT src_aox_reg_17__4_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[148]), .CLK(clk), .Q(src_window[148]) );
  DFFSSRX1_HVT src_aox_reg_17__3_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[147]), .CLK(clk), .Q(src_window[147]) );
  DFFSSRX1_HVT src_aox_reg_17__2_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[146]), .CLK(clk), .Q(src_window[146]) );
  DFFSSRX1_HVT src_aox_reg_17__1_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[145]), .CLK(clk), .Q(src_window[145]) );
  DFFSSRX1_HVT src_aox_reg_17__0_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[144]), .CLK(clk), .Q(src_window[144]) );
  DFFSSRX1_HVT src_aox_reg_18__7_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[143]), .CLK(clk), .Q(src_window[143]) );
  DFFSSRX1_HVT src_aox_reg_18__6_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[142]), .CLK(clk), .Q(src_window[142]) );
  DFFSSRX1_HVT src_aox_reg_18__5_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[141]), .CLK(clk), .Q(src_window[141]) );
  DFFSSRX1_HVT src_aox_reg_18__4_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[140]), .CLK(clk), .Q(src_window[140]) );
  DFFSSRX1_HVT src_aox_reg_18__3_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[139]), .CLK(clk), .Q(src_window[139]) );
  DFFSSRX1_HVT src_aox_reg_18__2_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[138]), .CLK(clk), .Q(src_window[138]) );
  DFFSSRX1_HVT src_aox_reg_18__1_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[137]), .CLK(clk), .Q(src_window[137]) );
  DFFSSRX1_HVT src_aox_reg_18__0_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[136]), .CLK(clk), .Q(src_window[136]) );
  DFFSSRX1_HVT src_aox_reg_19__7_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[135]), .CLK(clk), .Q(src_window[135]) );
  DFFSSRX1_HVT src_aox_reg_19__6_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[134]), .CLK(clk), .Q(src_window[134]) );
  DFFSSRX1_HVT src_aox_reg_19__5_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[133]), .CLK(clk), .Q(src_window[133]) );
  DFFSSRX1_HVT src_aox_reg_19__4_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[132]), .CLK(clk), .Q(src_window[132]) );
  DFFSSRX1_HVT src_aox_reg_19__3_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[131]), .CLK(clk), .Q(src_window[131]) );
  DFFSSRX1_HVT src_aox_reg_19__2_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[130]), .CLK(clk), .Q(src_window[130]) );
  DFFSSRX1_HVT src_aox_reg_19__1_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[129]), .CLK(clk), .Q(src_window[129]) );
  DFFSSRX1_HVT src_aox_reg_19__0_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[128]), .CLK(clk), .Q(src_window[128]) );
  DFFSSRX1_HVT src_aox_reg_20__7_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[127]), .CLK(clk), .Q(src_window[127]) );
  DFFSSRX1_HVT src_aox_reg_20__6_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[126]), .CLK(clk), .Q(src_window[126]) );
  DFFSSRX1_HVT src_aox_reg_20__5_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[125]), .CLK(clk), .Q(src_window[125]) );
  DFFSSRX1_HVT src_aox_reg_20__4_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[124]), .CLK(clk), .Q(src_window[124]) );
  DFFSSRX1_HVT src_aox_reg_20__3_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[123]), .CLK(clk), .Q(src_window[123]) );
  DFFSSRX1_HVT src_aox_reg_20__2_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[122]), .CLK(clk), .Q(src_window[122]) );
  DFFSSRX1_HVT src_aox_reg_20__1_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[121]), .CLK(clk), .Q(src_window[121]) );
  DFFSSRX1_HVT src_aox_reg_20__0_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[120]), .CLK(clk), .Q(src_window[120]) );
  DFFSSRX1_HVT src_aox_reg_21__7_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[119]), .CLK(clk), .Q(src_window[119]) );
  DFFSSRX1_HVT src_aox_reg_21__6_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[118]), .CLK(clk), .Q(src_window[118]) );
  DFFSSRX1_HVT src_aox_reg_21__5_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[117]), .CLK(clk), .Q(src_window[117]) );
  DFFSSRX1_HVT src_aox_reg_21__4_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[116]), .CLK(clk), .Q(src_window[116]) );
  DFFSSRX1_HVT src_aox_reg_21__3_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[115]), .CLK(clk), .Q(src_window[115]) );
  DFFSSRX1_HVT src_aox_reg_21__2_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[114]), .CLK(clk), .Q(src_window[114]) );
  DFFSSRX1_HVT src_aox_reg_21__1_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[113]), .CLK(clk), .Q(src_window[113]) );
  DFFSSRX1_HVT src_aox_reg_21__0_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[112]), .CLK(clk), .Q(src_window[112]) );
  DFFSSRX1_HVT src_aox_reg_22__7_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[111]), .CLK(clk), .Q(src_window[111]) );
  DFFSSRX1_HVT src_aox_reg_22__6_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[110]), .CLK(clk), .Q(src_window[110]) );
  DFFSSRX1_HVT src_aox_reg_22__5_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[109]), .CLK(clk), .Q(src_window[109]) );
  DFFSSRX1_HVT src_aox_reg_22__4_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[108]), .CLK(clk), .Q(src_window[108]) );
  DFFSSRX1_HVT src_aox_reg_22__3_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[107]), .CLK(clk), .Q(src_window[107]) );
  DFFSSRX1_HVT src_aox_reg_22__2_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[106]), .CLK(clk), .Q(src_window[106]) );
  DFFSSRX1_HVT src_aox_reg_22__1_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[105]), .CLK(clk), .Q(src_window[105]) );
  DFFSSRX1_HVT src_aox_reg_22__0_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[104]), .CLK(clk), .Q(src_window[104]) );
  DFFSSRX1_HVT src_aox_reg_23__7_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[103]), .CLK(clk), .Q(src_window[103]) );
  DFFSSRX1_HVT src_aox_reg_23__6_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[102]), .CLK(clk), .Q(src_window[102]) );
  DFFSSRX1_HVT src_aox_reg_23__5_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[101]), .CLK(clk), .Q(src_window[101]) );
  DFFSSRX1_HVT src_aox_reg_23__4_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[100]), .CLK(clk), .Q(src_window[100]) );
  DFFSSRX1_HVT src_aox_reg_23__3_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[99]), .CLK(clk), .Q(src_window[99]) );
  DFFSSRX1_HVT src_aox_reg_23__2_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[98]), .CLK(clk), .Q(src_window[98]) );
  DFFSSRX1_HVT src_aox_reg_23__1_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[97]), .CLK(clk), .Q(src_window[97]) );
  DFFSSRX1_HVT src_aox_reg_23__0_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[96]), .CLK(clk), .Q(src_window[96]) );
  DFFSSRX1_HVT src_aox_reg_24__7_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[95]), .CLK(clk), .Q(src_window[95]) );
  DFFSSRX1_HVT src_aox_reg_24__6_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[94]), .CLK(clk), .Q(src_window[94]) );
  DFFSSRX1_HVT src_aox_reg_24__5_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[93]), .CLK(clk), .Q(src_window[93]) );
  DFFSSRX1_HVT src_aox_reg_24__4_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[92]), .CLK(clk), .Q(src_window[92]) );
  DFFSSRX1_HVT src_aox_reg_24__3_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[91]), .CLK(clk), .Q(src_window[91]) );
  DFFSSRX1_HVT src_aox_reg_24__2_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[90]), .CLK(clk), .Q(src_window[90]) );
  DFFSSRX1_HVT src_aox_reg_24__1_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[89]), .CLK(clk), .Q(src_window[89]) );
  DFFSSRX1_HVT src_aox_reg_24__0_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[88]), .CLK(clk), .Q(src_window[88]) );
  DFFSSRX1_HVT src_aox_reg_25__7_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[87]), .CLK(clk), .Q(src_window[87]) );
  DFFSSRX1_HVT src_aox_reg_25__6_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[86]), .CLK(clk), .Q(src_window[86]) );
  DFFSSRX1_HVT src_aox_reg_25__5_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[85]), .CLK(clk), .Q(src_window[85]) );
  DFFSSRX1_HVT src_aox_reg_25__4_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[84]), .CLK(clk), .Q(src_window[84]) );
  DFFSSRX1_HVT src_aox_reg_25__3_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[83]), .CLK(clk), .Q(src_window[83]) );
  DFFSSRX1_HVT src_aox_reg_25__2_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[82]), .CLK(clk), .Q(src_window[82]) );
  DFFSSRX1_HVT src_aox_reg_25__1_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[81]), .CLK(clk), .Q(src_window[81]) );
  DFFSSRX1_HVT src_aox_reg_25__0_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[80]), .CLK(clk), .Q(src_window[80]) );
  DFFSSRX1_HVT src_aox_reg_26__7_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[79]), .CLK(clk), .Q(src_window[79]) );
  DFFSSRX1_HVT src_aox_reg_26__6_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[78]), .CLK(clk), .Q(src_window[78]) );
  DFFSSRX1_HVT src_aox_reg_26__5_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[77]), .CLK(clk), .Q(src_window[77]) );
  DFFSSRX1_HVT src_aox_reg_26__4_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[76]), .CLK(clk), .Q(src_window[76]) );
  DFFSSRX1_HVT src_aox_reg_26__3_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[75]), .CLK(clk), .Q(src_window[75]) );
  DFFSSRX1_HVT src_aox_reg_26__2_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[74]), .CLK(clk), .Q(src_window[74]) );
  DFFSSRX1_HVT src_aox_reg_26__1_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[73]), .CLK(clk), .Q(src_window[73]) );
  DFFSSRX1_HVT src_aox_reg_26__0_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[72]), .CLK(clk), .Q(src_window[72]) );
  DFFSSRX1_HVT src_aox_reg_27__7_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[71]), .CLK(clk), .Q(src_window[71]) );
  DFFSSRX1_HVT src_aox_reg_27__6_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[70]), .CLK(clk), .Q(src_window[70]) );
  DFFSSRX1_HVT src_aox_reg_27__5_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[69]), .CLK(clk), .Q(src_window[69]) );
  DFFSSRX1_HVT src_aox_reg_27__4_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[68]), .CLK(clk), .Q(src_window[68]) );
  DFFSSRX1_HVT src_aox_reg_27__3_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[67]), .CLK(clk), .Q(src_window[67]) );
  DFFSSRX1_HVT src_aox_reg_27__2_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[66]), .CLK(clk), .Q(src_window[66]) );
  DFFSSRX1_HVT src_aox_reg_27__1_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[65]), .CLK(clk), .Q(src_window[65]) );
  DFFSSRX1_HVT src_aox_reg_27__0_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[64]), .CLK(clk), .Q(src_window[64]) );
  DFFSSRX1_HVT src_aox_reg_28__7_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[63]), .CLK(clk), .Q(src_window[63]) );
  DFFSSRX1_HVT src_aox_reg_28__6_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[62]), .CLK(clk), .Q(src_window[62]) );
  DFFSSRX1_HVT src_aox_reg_28__5_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[61]), .CLK(clk), .Q(src_window[61]) );
  DFFSSRX1_HVT src_aox_reg_28__4_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[60]), .CLK(clk), .Q(src_window[60]) );
  DFFSSRX1_HVT src_aox_reg_28__3_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[59]), .CLK(clk), .Q(src_window[59]) );
  DFFSSRX1_HVT src_aox_reg_28__2_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[58]), .CLK(clk), .Q(src_window[58]) );
  DFFSSRX1_HVT src_aox_reg_28__1_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[57]), .CLK(clk), .Q(src_window[57]) );
  DFFSSRX1_HVT src_aox_reg_28__0_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[56]), .CLK(clk), .Q(src_window[56]) );
  DFFSSRX1_HVT src_aox_reg_29__7_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[55]), .CLK(clk), .Q(src_window[55]) );
  DFFSSRX1_HVT src_aox_reg_29__6_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[54]), .CLK(clk), .Q(src_window[54]) );
  DFFSSRX1_HVT src_aox_reg_29__5_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[53]), .CLK(clk), .Q(src_window[53]) );
  DFFSSRX1_HVT src_aox_reg_29__4_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[52]), .CLK(clk), .Q(src_window[52]) );
  DFFSSRX1_HVT src_aox_reg_29__3_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[51]), .CLK(clk), .Q(src_window[51]) );
  DFFSSRX1_HVT src_aox_reg_29__2_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[50]), .CLK(clk), .Q(src_window[50]) );
  DFFSSRX1_HVT src_aox_reg_29__1_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[49]), .CLK(clk), .Q(src_window[49]) );
  DFFSSRX1_HVT src_aox_reg_29__0_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[48]), .CLK(clk), .Q(src_window[48]) );
  DFFSSRX1_HVT src_aox_reg_30__7_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[47]), .CLK(clk), .Q(src_window[47]) );
  DFFSSRX1_HVT src_aox_reg_30__6_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[46]), .CLK(clk), .Q(src_window[46]) );
  DFFSSRX1_HVT src_aox_reg_30__5_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[45]), .CLK(clk), .Q(src_window[45]) );
  DFFSSRX1_HVT src_aox_reg_30__4_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[44]), .CLK(clk), .Q(src_window[44]) );
  DFFSSRX1_HVT src_aox_reg_30__3_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[43]), .CLK(clk), .Q(src_window[43]) );
  DFFSSRX1_HVT src_aox_reg_30__2_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[42]), .CLK(clk), .Q(src_window[42]) );
  DFFSSRX1_HVT src_aox_reg_30__1_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[41]), .CLK(clk), .Q(src_window[41]) );
  DFFSSRX1_HVT src_aox_reg_30__0_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[40]), .CLK(clk), .Q(src_window[40]) );
  DFFSSRX1_HVT src_aox_reg_31__7_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[39]), .CLK(clk), .Q(src_window[39]) );
  DFFSSRX1_HVT src_aox_reg_31__6_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[38]), .CLK(clk), .Q(src_window[38]) );
  DFFSSRX1_HVT src_aox_reg_31__5_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[37]), .CLK(clk), .Q(src_window[37]) );
  DFFSSRX1_HVT src_aox_reg_31__4_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[36]), .CLK(clk), .Q(src_window[36]) );
  DFFSSRX1_HVT src_aox_reg_31__3_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[35]), .CLK(clk), .Q(src_window[35]) );
  DFFSSRX1_HVT src_aox_reg_31__2_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[34]), .CLK(clk), .Q(src_window[34]) );
  DFFSSRX1_HVT src_aox_reg_31__1_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[33]), .CLK(clk), .Q(src_window[33]) );
  DFFSSRX1_HVT src_aox_reg_31__0_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[32]), .CLK(clk), .Q(src_window[32]) );
  DFFSSRX1_HVT src_aox_reg_32__7_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[31]), .CLK(clk), .Q(src_window[31]) );
  DFFSSRX1_HVT src_aox_reg_32__6_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[30]), .CLK(clk), .Q(src_window[30]) );
  DFFSSRX1_HVT src_aox_reg_32__5_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[29]), .CLK(clk), .Q(src_window[29]) );
  DFFSSRX1_HVT src_aox_reg_32__4_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[28]), .CLK(clk), .Q(src_window[28]) );
  DFFSSRX1_HVT src_aox_reg_32__3_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[27]), .CLK(clk), .Q(src_window[27]) );
  DFFSSRX1_HVT src_aox_reg_32__2_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[26]), .CLK(clk), .Q(src_window[26]) );
  DFFSSRX1_HVT src_aox_reg_32__1_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[25]), .CLK(clk), .Q(src_window[25]) );
  DFFSSRX1_HVT src_aox_reg_32__0_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[24]), .CLK(clk), .Q(src_window[24]) );
  DFFSSRX1_HVT src_aox_reg_33__7_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[23]), .CLK(clk), .Q(src_window[23]) );
  DFFSSRX1_HVT src_aox_reg_33__6_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[22]), .CLK(clk), .Q(src_window[22]) );
  DFFSSRX1_HVT src_aox_reg_33__5_ ( .D(1'b0), .SETB(n1390), .RSTB(
        n_src_aox[21]), .CLK(clk), .Q(src_window[21]) );
  DFFSSRX1_HVT src_aox_reg_33__4_ ( .D(1'b0), .SETB(n1450), .RSTB(
        n_src_aox[20]), .CLK(clk), .Q(src_window[20]) );
  DFFSSRX1_HVT src_aox_reg_33__3_ ( .D(1'b0), .SETB(n1490), .RSTB(
        n_src_aox[19]), .CLK(clk), .Q(src_window[19]) );
  DFFSSRX1_HVT src_aox_reg_33__2_ ( .D(1'b0), .SETB(n1420), .RSTB(
        n_src_aox[18]), .CLK(clk), .Q(src_window[18]) );
  DFFSSRX1_HVT src_aox_reg_33__1_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[17]), .CLK(clk), .Q(src_window[17]) );
  DFFSSRX1_HVT src_aox_reg_33__0_ ( .D(1'b0), .SETB(n1480), .RSTB(
        n_src_aox[16]), .CLK(clk), .Q(src_window[16]) );
  DFFSSRX1_HVT src_aox_reg_34__7_ ( .D(1'b0), .SETB(n1410), .RSTB(
        n_src_aox[15]), .CLK(clk), .Q(src_window[15]) );
  DFFSSRX1_HVT src_aox_reg_34__6_ ( .D(1'b0), .SETB(n1440), .RSTB(
        n_src_aox[14]), .CLK(clk), .Q(src_window[14]) );
  DFFSSRX1_HVT src_aox_reg_34__5_ ( .D(1'b0), .SETB(n1470), .RSTB(
        n_src_aox[13]), .CLK(clk), .Q(src_window[13]) );
  DFFSSRX1_HVT src_aox_reg_34__4_ ( .D(1'b0), .SETB(n1400), .RSTB(
        n_src_aox[12]), .CLK(clk), .Q(src_window[12]) );
  DFFSSRX1_HVT src_aox_reg_34__3_ ( .D(1'b0), .SETB(n1430), .RSTB(
        n_src_aox[11]), .CLK(clk), .Q(src_window[11]) );
  DFFSSRX1_HVT src_aox_reg_34__2_ ( .D(1'b0), .SETB(n1460), .RSTB(
        n_src_aox[10]), .CLK(clk), .Q(src_window[10]) );
  DFFSSRX1_HVT src_aox_reg_34__1_ ( .D(1'b0), .SETB(n1390), .RSTB(n_src_aox[9]), .CLK(clk), .Q(src_window[9]) );
  DFFSSRX1_HVT src_aox_reg_34__0_ ( .D(1'b0), .SETB(n1450), .RSTB(n_src_aox[8]), .CLK(clk), .Q(src_window[8]) );
  DFFSSRX1_HVT src_aox_reg_35__7_ ( .D(1'b0), .SETB(n1490), .RSTB(n_src_aox[7]), .CLK(clk), .Q(src_window[7]) );
  DFFSSRX1_HVT src_aox_reg_35__6_ ( .D(1'b0), .SETB(n1420), .RSTB(n_src_aox[6]), .CLK(clk), .Q(src_window[6]) );
  DFFSSRX1_HVT src_aox_reg_35__5_ ( .D(1'b0), .SETB(n1440), .RSTB(n_src_aox[5]), .CLK(clk), .Q(src_window[5]) );
  DFFSSRX1_HVT src_aox_reg_35__4_ ( .D(1'b0), .SETB(n1480), .RSTB(n_src_aox[4]), .CLK(clk), .Q(src_window[4]) );
  DFFSSRX1_HVT src_aox_reg_35__3_ ( .D(1'b0), .SETB(n1410), .RSTB(n_src_aox[3]), .CLK(clk), .Q(src_window[3]) );
  DFFSSRX1_HVT src_aox_reg_35__2_ ( .D(1'b0), .SETB(n1430), .RSTB(n_src_aox[2]), .CLK(clk), .Q(src_window[2]) );
  DFFSSRX1_HVT src_aox_reg_35__1_ ( .D(1'b0), .SETB(n1470), .RSTB(n_src_aox[1]), .CLK(clk), .Q(src_window[1]) );
  DFFSSRX1_HVT src_aox_reg_35__0_ ( .D(1'b0), .SETB(n1400), .RSTB(n_src_aox[0]), .CLK(clk), .Q(src_window[0]) );
  DFFSSRX1_HVT conv1_weight_reg_99_ ( .D(1'b0), .SETB(n4800), .RSTB(
        sram_rdata_weight[99]), .CLK(clk), .Q(conv1_weight[99]) );
  DFFSSRX1_HVT weight_reg_99_ ( .D(1'b0), .SETB(n777), .RSTB(conv1_weight[99]), 
        .CLK(clk), .Q(weight[99]) );
  DFFSSRX1_HVT conv1_weight_reg_98_ ( .D(1'b0), .SETB(n34), .RSTB(
        sram_rdata_weight[98]), .CLK(clk), .Q(conv1_weight[98]) );
  DFFSSRX1_HVT weight_reg_98_ ( .D(1'b0), .SETB(n1760), .RSTB(conv1_weight[98]), .CLK(clk), .Q(weight[98]) );
  DFFSSRX1_HVT conv1_weight_reg_97_ ( .D(1'b0), .SETB(n34), .RSTB(
        sram_rdata_weight[97]), .CLK(clk), .Q(conv1_weight[97]) );
  DFFSSRX1_HVT weight_reg_97_ ( .D(1'b0), .SETB(n33), .RSTB(conv1_weight[97]), 
        .CLK(clk), .Q(weight[97]) );
  DFFSSRX1_HVT conv1_weight_reg_96_ ( .D(1'b0), .SETB(n33), .RSTB(
        sram_rdata_weight[96]), .CLK(clk), .Q(conv1_weight[96]) );
  DFFSSRX1_HVT weight_reg_96_ ( .D(1'b0), .SETB(n1760), .RSTB(conv1_weight[96]), .CLK(clk), .Q(weight[96]) );
  DFFSSRX1_HVT conv1_weight_reg_95_ ( .D(1'b0), .SETB(n4800), .RSTB(
        sram_rdata_weight[95]), .CLK(clk), .Q(conv1_weight[95]) );
  DFFSSRX1_HVT weight_reg_95_ ( .D(1'b0), .SETB(n7700), .RSTB(conv1_weight[95]), .CLK(clk), .Q(weight[95]) );
  DFFSSRX1_HVT conv1_weight_reg_94_ ( .D(1'b0), .SETB(n7700), .RSTB(
        sram_rdata_weight[94]), .CLK(clk), .Q(conv1_weight[94]) );
  DFFSSRX1_HVT weight_reg_94_ ( .D(1'b0), .SETB(n1760), .RSTB(conv1_weight[94]), .CLK(clk), .Q(weight[94]) );
  DFFSSRX1_HVT conv1_weight_reg_93_ ( .D(1'b0), .SETB(n34), .RSTB(
        sram_rdata_weight[93]), .CLK(clk), .Q(conv1_weight[93]) );
  DFFSSRX1_HVT weight_reg_93_ ( .D(1'b0), .SETB(n33), .RSTB(conv1_weight[93]), 
        .CLK(clk), .Q(weight[93]) );
  DFFSSRX1_HVT conv1_weight_reg_92_ ( .D(1'b0), .SETB(n33), .RSTB(
        sram_rdata_weight[92]), .CLK(clk), .Q(conv1_weight[92]) );
  DFFSSRX1_HVT weight_reg_92_ ( .D(1'b0), .SETB(n1760), .RSTB(conv1_weight[92]), .CLK(clk), .Q(weight[92]) );
  DFFSSRX1_HVT conv1_weight_reg_91_ ( .D(1'b0), .SETB(n4800), .RSTB(
        sram_rdata_weight[91]), .CLK(clk), .Q(conv1_weight[91]) );
  DFFSSRX1_HVT weight_reg_91_ ( .D(1'b0), .SETB(n7800), .RSTB(conv1_weight[91]), .CLK(clk), .Q(weight[91]) );
  DFFSSRX1_HVT conv1_weight_reg_90_ ( .D(1'b0), .SETB(n7800), .RSTB(
        sram_rdata_weight[90]), .CLK(clk), .Q(conv1_weight[90]) );
  DFFSSRX1_HVT weight_reg_90_ ( .D(1'b0), .SETB(n1760), .RSTB(conv1_weight[90]), .CLK(clk), .Q(weight[90]) );
  DFFSSRX1_HVT conv1_weight_reg_89_ ( .D(1'b0), .SETB(n34), .RSTB(
        sram_rdata_weight[89]), .CLK(clk), .Q(conv1_weight[89]) );
  DFFSSRX1_HVT weight_reg_89_ ( .D(1'b0), .SETB(n4900), .RSTB(conv1_weight[89]), .CLK(clk), .Q(weight[89]) );
  DFFSSRX1_HVT conv1_weight_reg_88_ ( .D(1'b0), .SETB(n4900), .RSTB(
        sram_rdata_weight[88]), .CLK(clk), .Q(conv1_weight[88]) );
  DFFSSRX1_HVT weight_reg_88_ ( .D(1'b0), .SETB(n1760), .RSTB(conv1_weight[88]), .CLK(clk), .Q(weight[88]) );
  DFFSSRX1_HVT conv1_weight_reg_87_ ( .D(1'b0), .SETB(n4800), .RSTB(
        sram_rdata_weight[87]), .CLK(clk), .Q(conv1_weight[87]) );
  DFFSSRX1_HVT weight_reg_87_ ( .D(1'b0), .SETB(n7900), .RSTB(conv1_weight[87]), .CLK(clk), .Q(weight[87]) );
  DFFSSRX1_HVT conv1_weight_reg_86_ ( .D(1'b0), .SETB(n7900), .RSTB(
        sram_rdata_weight[86]), .CLK(clk), .Q(conv1_weight[86]) );
  DFFSSRX1_HVT weight_reg_86_ ( .D(1'b0), .SETB(n1760), .RSTB(conv1_weight[86]), .CLK(clk), .Q(weight[86]) );
  DFFSSRX1_HVT conv1_weight_reg_85_ ( .D(1'b0), .SETB(n34), .RSTB(
        sram_rdata_weight[85]), .CLK(clk), .Q(conv1_weight[85]) );
  DFFSSRX1_HVT weight_reg_85_ ( .D(1'b0), .SETB(n4900), .RSTB(conv1_weight[85]), .CLK(clk), .Q(weight[85]) );
  DFFSSRX1_HVT conv1_weight_reg_84_ ( .D(1'b0), .SETB(n4900), .RSTB(
        sram_rdata_weight[84]), .CLK(clk), .Q(conv1_weight[84]) );
  DFFSSRX1_HVT weight_reg_84_ ( .D(1'b0), .SETB(n1760), .RSTB(conv1_weight[84]), .CLK(clk), .Q(weight[84]) );
  DFFSSRX1_HVT conv1_weight_reg_83_ ( .D(1'b0), .SETB(n4800), .RSTB(
        sram_rdata_weight[83]), .CLK(clk), .Q(conv1_weight[83]) );
  DFFSSRX1_HVT weight_reg_83_ ( .D(1'b0), .SETB(n777), .RSTB(conv1_weight[83]), 
        .CLK(clk), .Q(weight[83]) );
  DFFSSRX1_HVT conv1_weight_reg_82_ ( .D(1'b0), .SETB(n4800), .RSTB(
        sram_rdata_weight[82]), .CLK(clk), .Q(conv1_weight[82]) );
  DFFSSRX1_HVT weight_reg_82_ ( .D(1'b0), .SETB(n1760), .RSTB(conv1_weight[82]), .CLK(clk), .Q(weight[82]) );
  DFFSSRX1_HVT conv1_weight_reg_81_ ( .D(1'b0), .SETB(n34), .RSTB(
        sram_rdata_weight[81]), .CLK(clk), .Q(conv1_weight[81]) );
  DFFSSRX1_HVT weight_reg_81_ ( .D(1'b0), .SETB(n33), .RSTB(conv1_weight[81]), 
        .CLK(clk), .Q(weight[81]) );
  DFFSSRX1_HVT conv1_weight_reg_80_ ( .D(1'b0), .SETB(n33), .RSTB(
        sram_rdata_weight[80]), .CLK(clk), .Q(conv1_weight[80]) );
  DFFSSRX1_HVT weight_reg_80_ ( .D(1'b0), .SETB(n1760), .RSTB(conv1_weight[80]), .CLK(clk), .Q(weight[80]) );
  DFFSSRX1_HVT conv1_weight_reg_79_ ( .D(1'b0), .SETB(n4800), .RSTB(
        sram_rdata_weight[79]), .CLK(clk), .Q(conv1_weight[79]) );
  DFFSSRX1_HVT weight_reg_79_ ( .D(1'b0), .SETB(n7700), .RSTB(conv1_weight[79]), .CLK(clk), .Q(weight[79]) );
  DFFSSRX1_HVT conv1_weight_reg_78_ ( .D(1'b0), .SETB(n7700), .RSTB(
        sram_rdata_weight[78]), .CLK(clk), .Q(conv1_weight[78]) );
  DFFSSRX1_HVT weight_reg_78_ ( .D(1'b0), .SETB(n1760), .RSTB(conv1_weight[78]), .CLK(clk), .Q(weight[78]) );
  DFFSSRX1_HVT conv1_weight_reg_77_ ( .D(1'b0), .SETB(n34), .RSTB(
        sram_rdata_weight[77]), .CLK(clk), .Q(conv1_weight[77]) );
  DFFSSRX1_HVT weight_reg_77_ ( .D(1'b0), .SETB(n33), .RSTB(conv1_weight[77]), 
        .CLK(clk), .Q(weight[77]) );
  DFFSSRX1_HVT conv1_weight_reg_76_ ( .D(1'b0), .SETB(n33), .RSTB(
        sram_rdata_weight[76]), .CLK(clk), .Q(conv1_weight[76]) );
  DFFSSRX1_HVT weight_reg_76_ ( .D(1'b0), .SETB(n1760), .RSTB(conv1_weight[76]), .CLK(clk), .Q(weight[76]) );
  DFFSSRX1_HVT conv1_weight_reg_75_ ( .D(1'b0), .SETB(n4800), .RSTB(
        sram_rdata_weight[75]), .CLK(clk), .Q(conv1_weight[75]) );
  DFFSSRX1_HVT weight_reg_75_ ( .D(1'b0), .SETB(n7800), .RSTB(conv1_weight[75]), .CLK(clk), .Q(weight[75]) );
  DFFSSRX1_HVT conv1_weight_reg_74_ ( .D(1'b0), .SETB(n7800), .RSTB(
        sram_rdata_weight[74]), .CLK(clk), .Q(conv1_weight[74]) );
  DFFSSRX1_HVT weight_reg_74_ ( .D(1'b0), .SETB(n1760), .RSTB(conv1_weight[74]), .CLK(clk), .Q(weight[74]) );
  DFFSSRX1_HVT conv1_weight_reg_73_ ( .D(1'b0), .SETB(n34), .RSTB(
        sram_rdata_weight[73]), .CLK(clk), .Q(conv1_weight[73]) );
  DFFSSRX1_HVT weight_reg_73_ ( .D(1'b0), .SETB(n4900), .RSTB(conv1_weight[73]), .CLK(clk), .Q(weight[73]) );
  DFFSSRX1_HVT conv1_weight_reg_72_ ( .D(1'b0), .SETB(n4900), .RSTB(
        sram_rdata_weight[72]), .CLK(clk), .Q(conv1_weight[72]) );
  DFFSSRX1_HVT weight_reg_72_ ( .D(1'b0), .SETB(n1760), .RSTB(conv1_weight[72]), .CLK(clk), .Q(weight[72]) );
  DFFSSRX1_HVT conv1_weight_reg_71_ ( .D(1'b0), .SETB(n4800), .RSTB(
        sram_rdata_weight[71]), .CLK(clk), .Q(conv1_weight[71]) );
  DFFSSRX1_HVT weight_reg_71_ ( .D(1'b0), .SETB(n7900), .RSTB(conv1_weight[71]), .CLK(clk), .Q(weight[71]) );
  DFFSSRX1_HVT conv1_weight_reg_70_ ( .D(1'b0), .SETB(n7900), .RSTB(
        sram_rdata_weight[70]), .CLK(clk), .Q(conv1_weight[70]) );
  DFFSSRX1_HVT weight_reg_70_ ( .D(1'b0), .SETB(n1760), .RSTB(conv1_weight[70]), .CLK(clk), .Q(weight[70]) );
  DFFSSRX1_HVT conv1_weight_reg_69_ ( .D(1'b0), .SETB(n34), .RSTB(
        sram_rdata_weight[69]), .CLK(clk), .Q(conv1_weight[69]) );
  DFFSSRX1_HVT weight_reg_69_ ( .D(1'b0), .SETB(n4900), .RSTB(conv1_weight[69]), .CLK(clk), .Q(weight[69]) );
  DFFSSRX1_HVT conv1_weight_reg_68_ ( .D(1'b0), .SETB(n4900), .RSTB(
        sram_rdata_weight[68]), .CLK(clk), .Q(conv1_weight[68]) );
  DFFSSRX1_HVT weight_reg_68_ ( .D(1'b0), .SETB(n1760), .RSTB(conv1_weight[68]), .CLK(clk), .Q(weight[68]) );
  DFFSSRX1_HVT conv1_weight_reg_67_ ( .D(1'b0), .SETB(n4800), .RSTB(
        sram_rdata_weight[67]), .CLK(clk), .Q(conv1_weight[67]) );
  DFFSSRX1_HVT weight_reg_67_ ( .D(1'b0), .SETB(n777), .RSTB(conv1_weight[67]), 
        .CLK(clk), .Q(weight[67]) );
  DFFSSRX1_HVT conv1_weight_reg_66_ ( .D(1'b0), .SETB(n1370), .RSTB(
        sram_rdata_weight[66]), .CLK(clk), .Q(conv1_weight[66]) );
  DFFSSRX1_HVT weight_reg_66_ ( .D(1'b0), .SETB(n1760), .RSTB(conv1_weight[66]), .CLK(clk), .Q(weight[66]) );
  DFFSSRX1_HVT conv1_weight_reg_65_ ( .D(1'b0), .SETB(n34), .RSTB(
        sram_rdata_weight[65]), .CLK(clk), .Q(conv1_weight[65]) );
  DFFSSRX1_HVT weight_reg_65_ ( .D(1'b0), .SETB(n33), .RSTB(conv1_weight[65]), 
        .CLK(clk), .Q(weight[65]) );
  DFFSSRX1_HVT conv1_weight_reg_64_ ( .D(1'b0), .SETB(n33), .RSTB(
        sram_rdata_weight[64]), .CLK(clk), .Q(conv1_weight[64]) );
  DFFSSRX1_HVT weight_reg_64_ ( .D(1'b0), .SETB(n1760), .RSTB(conv1_weight[64]), .CLK(clk), .Q(weight[64]) );
  DFFSSRX1_HVT conv1_weight_reg_63_ ( .D(1'b0), .SETB(n4800), .RSTB(
        sram_rdata_weight[63]), .CLK(clk), .Q(conv1_weight[63]) );
  DFFSSRX1_HVT weight_reg_63_ ( .D(1'b0), .SETB(n7700), .RSTB(conv1_weight[63]), .CLK(clk), .Q(weight[63]) );
  DFFSSRX1_HVT conv1_weight_reg_62_ ( .D(1'b0), .SETB(n7700), .RSTB(
        sram_rdata_weight[62]), .CLK(clk), .Q(conv1_weight[62]) );
  DFFSSRX1_HVT weight_reg_62_ ( .D(1'b0), .SETB(n1760), .RSTB(conv1_weight[62]), .CLK(clk), .Q(weight[62]) );
  DFFSSRX1_HVT conv1_weight_reg_61_ ( .D(1'b0), .SETB(n34), .RSTB(
        sram_rdata_weight[61]), .CLK(clk), .Q(conv1_weight[61]) );
  DFFSSRX1_HVT weight_reg_61_ ( .D(1'b0), .SETB(n33), .RSTB(conv1_weight[61]), 
        .CLK(clk), .Q(weight[61]) );
  DFFSSRX1_HVT conv1_weight_reg_60_ ( .D(1'b0), .SETB(n33), .RSTB(
        sram_rdata_weight[60]), .CLK(clk), .Q(conv1_weight[60]) );
  DFFSSRX1_HVT weight_reg_60_ ( .D(1'b0), .SETB(n1760), .RSTB(conv1_weight[60]), .CLK(clk), .Q(weight[60]) );
  DFFSSRX1_HVT conv1_weight_reg_59_ ( .D(1'b0), .SETB(n4800), .RSTB(
        sram_rdata_weight[59]), .CLK(clk), .Q(conv1_weight[59]) );
  DFFSSRX1_HVT weight_reg_59_ ( .D(1'b0), .SETB(n7800), .RSTB(conv1_weight[59]), .CLK(clk), .Q(weight[59]) );
  DFFSSRX1_HVT conv1_weight_reg_58_ ( .D(1'b0), .SETB(n7800), .RSTB(
        sram_rdata_weight[58]), .CLK(clk), .Q(conv1_weight[58]) );
  DFFSSRX1_HVT weight_reg_58_ ( .D(1'b0), .SETB(n1760), .RSTB(conv1_weight[58]), .CLK(clk), .Q(weight[58]) );
  DFFSSRX1_HVT conv1_weight_reg_57_ ( .D(1'b0), .SETB(n34), .RSTB(
        sram_rdata_weight[57]), .CLK(clk), .Q(conv1_weight[57]) );
  DFFSSRX1_HVT weight_reg_57_ ( .D(1'b0), .SETB(n4900), .RSTB(conv1_weight[57]), .CLK(clk), .Q(weight[57]) );
  DFFSSRX1_HVT conv1_weight_reg_56_ ( .D(1'b0), .SETB(n4900), .RSTB(
        sram_rdata_weight[56]), .CLK(clk), .Q(conv1_weight[56]) );
  DFFSSRX1_HVT weight_reg_56_ ( .D(1'b0), .SETB(n7800), .RSTB(conv1_weight[56]), .CLK(clk), .Q(weight[56]) );
  DFFSSRX1_HVT conv1_weight_reg_55_ ( .D(1'b0), .SETB(n4800), .RSTB(
        sram_rdata_weight[55]), .CLK(clk), .Q(conv1_weight[55]) );
  DFFSSRX1_HVT weight_reg_55_ ( .D(1'b0), .SETB(n7900), .RSTB(conv1_weight[55]), .CLK(clk), .Q(weight[55]) );
  DFFSSRX1_HVT conv1_weight_reg_54_ ( .D(1'b0), .SETB(n7900), .RSTB(
        sram_rdata_weight[54]), .CLK(clk), .Q(conv1_weight[54]) );
  DFFSSRX1_HVT weight_reg_54_ ( .D(1'b0), .SETB(n7700), .RSTB(conv1_weight[54]), .CLK(clk), .Q(weight[54]) );
  DFFSSRX1_HVT conv1_weight_reg_53_ ( .D(1'b0), .SETB(n34), .RSTB(
        sram_rdata_weight[53]), .CLK(clk), .Q(conv1_weight[53]) );
  DFFSSRX1_HVT weight_reg_53_ ( .D(1'b0), .SETB(n4900), .RSTB(conv1_weight[53]), .CLK(clk), .Q(weight[53]) );
  DFFSSRX1_HVT conv1_weight_reg_52_ ( .D(1'b0), .SETB(n4900), .RSTB(
        sram_rdata_weight[52]), .CLK(clk), .Q(conv1_weight[52]) );
  DFFSSRX1_HVT weight_reg_52_ ( .D(1'b0), .SETB(n777), .RSTB(conv1_weight[52]), 
        .CLK(clk), .Q(weight[52]) );
  DFFSSRX1_HVT conv1_weight_reg_51_ ( .D(1'b0), .SETB(n4800), .RSTB(
        sram_rdata_weight[51]), .CLK(clk), .Q(conv1_weight[51]) );
  DFFSSRX1_HVT weight_reg_51_ ( .D(1'b0), .SETB(n777), .RSTB(conv1_weight[51]), 
        .CLK(clk), .Q(weight[51]) );
  DFFSSRX1_HVT conv1_weight_reg_50_ ( .D(1'b0), .SETB(n1810), .RSTB(
        sram_rdata_weight[50]), .CLK(clk), .Q(conv1_weight[50]) );
  DFFSSRX1_HVT weight_reg_50_ ( .D(1'b0), .SETB(n7800), .RSTB(conv1_weight[50]), .CLK(clk), .Q(weight[50]) );
  DFFSSRX1_HVT conv1_weight_reg_49_ ( .D(1'b0), .SETB(n34), .RSTB(
        sram_rdata_weight[49]), .CLK(clk), .Q(conv1_weight[49]) );
  DFFSSRX1_HVT weight_reg_49_ ( .D(1'b0), .SETB(n33), .RSTB(conv1_weight[49]), 
        .CLK(clk), .Q(weight[49]) );
  DFFSSRX1_HVT conv1_weight_reg_48_ ( .D(1'b0), .SETB(n33), .RSTB(
        sram_rdata_weight[48]), .CLK(clk), .Q(conv1_weight[48]) );
  DFFSSRX1_HVT weight_reg_48_ ( .D(1'b0), .SETB(n7700), .RSTB(conv1_weight[48]), .CLK(clk), .Q(weight[48]) );
  DFFSSRX1_HVT conv1_weight_reg_47_ ( .D(1'b0), .SETB(n4800), .RSTB(
        sram_rdata_weight[47]), .CLK(clk), .Q(conv1_weight[47]) );
  DFFSSRX1_HVT weight_reg_47_ ( .D(1'b0), .SETB(n7700), .RSTB(conv1_weight[47]), .CLK(clk), .Q(weight[47]) );
  DFFSSRX1_HVT conv1_weight_reg_46_ ( .D(1'b0), .SETB(n7700), .RSTB(
        sram_rdata_weight[46]), .CLK(clk), .Q(conv1_weight[46]) );
  DFFSSRX1_HVT weight_reg_46_ ( .D(1'b0), .SETB(n777), .RSTB(conv1_weight[46]), 
        .CLK(clk), .Q(weight[46]) );
  DFFSSRX1_HVT conv1_weight_reg_45_ ( .D(1'b0), .SETB(n34), .RSTB(
        sram_rdata_weight[45]), .CLK(clk), .Q(conv1_weight[45]) );
  DFFSSRX1_HVT weight_reg_45_ ( .D(1'b0), .SETB(n33), .RSTB(conv1_weight[45]), 
        .CLK(clk), .Q(weight[45]) );
  DFFSSRX1_HVT conv1_weight_reg_44_ ( .D(1'b0), .SETB(n33), .RSTB(
        sram_rdata_weight[44]), .CLK(clk), .Q(conv1_weight[44]) );
  DFFSSRX1_HVT weight_reg_44_ ( .D(1'b0), .SETB(n7900), .RSTB(conv1_weight[44]), .CLK(clk), .Q(weight[44]) );
  DFFSSRX1_HVT conv1_weight_reg_43_ ( .D(1'b0), .SETB(n4800), .RSTB(
        sram_rdata_weight[43]), .CLK(clk), .Q(conv1_weight[43]) );
  DFFSSRX1_HVT weight_reg_43_ ( .D(1'b0), .SETB(n7800), .RSTB(conv1_weight[43]), .CLK(clk), .Q(weight[43]) );
  DFFSSRX1_HVT conv1_weight_reg_42_ ( .D(1'b0), .SETB(n7800), .RSTB(
        sram_rdata_weight[42]), .CLK(clk), .Q(conv1_weight[42]) );
  DFFSSRX1_HVT weight_reg_42_ ( .D(1'b0), .SETB(n7900), .RSTB(conv1_weight[42]), .CLK(clk), .Q(weight[42]) );
  DFFSSRX1_HVT conv1_weight_reg_41_ ( .D(1'b0), .SETB(n34), .RSTB(
        sram_rdata_weight[41]), .CLK(clk), .Q(conv1_weight[41]) );
  DFFSSRX1_HVT weight_reg_41_ ( .D(1'b0), .SETB(n4900), .RSTB(conv1_weight[41]), .CLK(clk), .Q(weight[41]) );
  DFFSSRX1_HVT conv1_weight_reg_40_ ( .D(1'b0), .SETB(n4900), .RSTB(
        sram_rdata_weight[40]), .CLK(clk), .Q(conv1_weight[40]) );
  DFFSSRX1_HVT weight_reg_40_ ( .D(1'b0), .SETB(n7900), .RSTB(conv1_weight[40]), .CLK(clk), .Q(weight[40]) );
  DFFSSRX1_HVT conv1_weight_reg_39_ ( .D(1'b0), .SETB(n4800), .RSTB(
        sram_rdata_weight[39]), .CLK(clk), .Q(conv1_weight[39]) );
  DFFSSRX1_HVT weight_reg_39_ ( .D(1'b0), .SETB(n7900), .RSTB(conv1_weight[39]), .CLK(clk), .Q(weight[39]) );
  DFFSSRX1_HVT conv1_weight_reg_38_ ( .D(1'b0), .SETB(n7900), .RSTB(
        sram_rdata_weight[38]), .CLK(clk), .Q(conv1_weight[38]) );
  DFFSSRX1_HVT weight_reg_38_ ( .D(1'b0), .SETB(n33), .RSTB(conv1_weight[38]), 
        .CLK(clk), .Q(weight[38]) );
  DFFSSRX1_HVT conv1_weight_reg_37_ ( .D(1'b0), .SETB(n34), .RSTB(
        sram_rdata_weight[37]), .CLK(clk), .Q(conv1_weight[37]) );
  DFFSSRX1_HVT weight_reg_37_ ( .D(1'b0), .SETB(n4900), .RSTB(conv1_weight[37]), .CLK(clk), .Q(weight[37]) );
  DFFSSRX1_HVT conv1_weight_reg_36_ ( .D(1'b0), .SETB(n4900), .RSTB(
        sram_rdata_weight[36]), .CLK(clk), .Q(conv1_weight[36]) );
  DFFSSRX1_HVT weight_reg_36_ ( .D(1'b0), .SETB(n4900), .RSTB(conv1_weight[36]), .CLK(clk), .Q(weight[36]) );
  DFFSSRX1_HVT conv1_weight_reg_35_ ( .D(1'b0), .SETB(n4800), .RSTB(
        sram_rdata_weight[35]), .CLK(clk), .Q(conv1_weight[35]) );
  DFFSSRX1_HVT weight_reg_35_ ( .D(1'b0), .SETB(n777), .RSTB(conv1_weight[35]), 
        .CLK(clk), .Q(weight[35]) );
  DFFSSRX1_HVT conv1_weight_reg_34_ ( .D(1'b0), .SETB(n1530), .RSTB(
        sram_rdata_weight[34]), .CLK(clk), .Q(conv1_weight[34]) );
  DFFSSRX1_HVT weight_reg_34_ ( .D(1'b0), .SETB(n1810), .RSTB(conv1_weight[34]), .CLK(clk), .Q(weight[34]) );
  DFFSSRX1_HVT conv1_weight_reg_33_ ( .D(1'b0), .SETB(n1370), .RSTB(
        sram_rdata_weight[33]), .CLK(clk), .Q(conv1_weight[33]) );
  DFFSSRX1_HVT weight_reg_33_ ( .D(1'b0), .SETB(n777), .RSTB(conv1_weight[33]), 
        .CLK(clk), .Q(weight[33]) );
  DFFSSRX1_HVT conv1_weight_reg_32_ ( .D(1'b0), .SETB(n1510), .RSTB(
        sram_rdata_weight[32]), .CLK(clk), .Q(conv1_weight[32]) );
  DFFSSRX1_HVT weight_reg_32_ ( .D(1'b0), .SETB(n1810), .RSTB(conv1_weight[32]), .CLK(clk), .Q(weight[32]) );
  DFFSSRX1_HVT conv1_weight_reg_31_ ( .D(1'b0), .SETB(n13500), .RSTB(
        sram_rdata_weight[31]), .CLK(clk), .Q(conv1_weight[31]) );
  DFFSSRX1_HVT weight_reg_31_ ( .D(1'b0), .SETB(n4900), .RSTB(conv1_weight[31]), .CLK(clk), .Q(weight[31]) );
  DFFSSRX1_HVT conv1_weight_reg_30_ ( .D(1'b0), .SETB(n1500), .RSTB(
        sram_rdata_weight[30]), .CLK(clk), .Q(conv1_weight[30]) );
  DFFSSRX1_HVT weight_reg_30_ ( .D(1'b0), .SETB(n1810), .RSTB(conv1_weight[30]), .CLK(clk), .Q(weight[30]) );
  DFFSSRX1_HVT conv1_weight_reg_29_ ( .D(1'b0), .SETB(n13600), .RSTB(
        sram_rdata_weight[29]), .CLK(clk), .Q(conv1_weight[29]) );
  DFFSSRX1_HVT weight_reg_29_ ( .D(1'b0), .SETB(n34), .RSTB(conv1_weight[29]), 
        .CLK(clk), .Q(weight[29]) );
  DFFSSRX1_HVT conv1_weight_reg_28_ ( .D(1'b0), .SETB(n1530), .RSTB(
        sram_rdata_weight[28]), .CLK(clk), .Q(conv1_weight[28]) );
  DFFSSRX1_HVT weight_reg_28_ ( .D(1'b0), .SETB(n1810), .RSTB(conv1_weight[28]), .CLK(clk), .Q(weight[28]) );
  DFFSSRX1_HVT conv1_weight_reg_27_ ( .D(1'b0), .SETB(n1370), .RSTB(
        sram_rdata_weight[27]), .CLK(clk), .Q(conv1_weight[27]) );
  DFFSSRX1_HVT weight_reg_27_ ( .D(1'b0), .SETB(n33), .RSTB(conv1_weight[27]), 
        .CLK(clk), .Q(weight[27]) );
  DFFSSRX1_HVT conv1_weight_reg_26_ ( .D(1'b0), .SETB(n1510), .RSTB(
        sram_rdata_weight[26]), .CLK(clk), .Q(conv1_weight[26]) );
  DFFSSRX1_HVT weight_reg_26_ ( .D(1'b0), .SETB(n1810), .RSTB(conv1_weight[26]), .CLK(clk), .Q(weight[26]) );
  DFFSSRX1_HVT conv1_weight_reg_25_ ( .D(1'b0), .SETB(n1380), .RSTB(
        sram_rdata_weight[25]), .CLK(clk), .Q(conv1_weight[25]) );
  DFFSSRX1_HVT weight_reg_25_ ( .D(1'b0), .SETB(n33), .RSTB(conv1_weight[25]), 
        .CLK(clk), .Q(weight[25]) );
  DFFSSRX1_HVT conv1_weight_reg_24_ ( .D(1'b0), .SETB(n1520), .RSTB(
        sram_rdata_weight[24]), .CLK(clk), .Q(conv1_weight[24]) );
  DFFSSRX1_HVT weight_reg_24_ ( .D(1'b0), .SETB(n1810), .RSTB(conv1_weight[24]), .CLK(clk), .Q(weight[24]) );
  DFFSSRX1_HVT conv1_weight_reg_23_ ( .D(1'b0), .SETB(n13600), .RSTB(
        sram_rdata_weight[23]), .CLK(clk), .Q(conv1_weight[23]) );
  DFFSSRX1_HVT weight_reg_23_ ( .D(1'b0), .SETB(n4900), .RSTB(conv1_weight[23]), .CLK(clk), .Q(weight[23]) );
  DFFSSRX1_HVT conv1_weight_reg_22_ ( .D(1'b0), .SETB(n1530), .RSTB(
        sram_rdata_weight[22]), .CLK(clk), .Q(conv1_weight[22]) );
  DFFSSRX1_HVT weight_reg_22_ ( .D(1'b0), .SETB(n1810), .RSTB(conv1_weight[22]), .CLK(clk), .Q(weight[22]) );
  DFFSSRX1_HVT conv1_weight_reg_21_ ( .D(1'b0), .SETB(n1370), .RSTB(
        sram_rdata_weight[21]), .CLK(clk), .Q(conv1_weight[21]) );
  DFFSSRX1_HVT weight_reg_21_ ( .D(1'b0), .SETB(n1510), .RSTB(conv1_weight[21]), .CLK(clk), .Q(weight[21]) );
  DFFSSRX1_HVT conv1_weight_reg_20_ ( .D(1'b0), .SETB(n1810), .RSTB(
        sram_rdata_weight[20]), .CLK(clk), .Q(conv1_weight[20]) );
  DFFSSRX1_HVT weight_reg_20_ ( .D(1'b0), .SETB(n13500), .RSTB(
        conv1_weight[20]), .CLK(clk), .Q(weight[20]) );
  DFFSSRX1_HVT conv1_weight_reg_19_ ( .D(1'b0), .SETB(n4800), .RSTB(
        sram_rdata_weight[19]), .CLK(clk), .Q(conv1_weight[19]) );
  DFFSSRX1_HVT weight_reg_19_ ( .D(1'b0), .SETB(n1500), .RSTB(conv1_weight[19]), .CLK(clk), .Q(weight[19]) );
  DFFSSRX1_HVT conv1_weight_reg_18_ ( .D(1'b0), .SETB(n1810), .RSTB(
        sram_rdata_weight[18]), .CLK(clk), .Q(conv1_weight[18]) );
  DFFSSRX1_HVT weight_reg_18_ ( .D(1'b0), .SETB(n13600), .RSTB(
        conv1_weight[18]), .CLK(clk), .Q(weight[18]) );
  DFFSSRX1_HVT conv1_weight_reg_17_ ( .D(1'b0), .SETB(n7700), .RSTB(
        sram_rdata_weight[17]), .CLK(clk), .Q(conv1_weight[17]) );
  DFFSSRX1_HVT weight_reg_17_ ( .D(1'b0), .SETB(n1530), .RSTB(conv1_weight[17]), .CLK(clk), .Q(weight[17]) );
  DFFSSRX1_HVT conv1_weight_reg_16_ ( .D(1'b0), .SETB(n1810), .RSTB(
        sram_rdata_weight[16]), .CLK(clk), .Q(conv1_weight[16]) );
  DFFSSRX1_HVT weight_reg_16_ ( .D(1'b0), .SETB(n1370), .RSTB(conv1_weight[16]), .CLK(clk), .Q(weight[16]) );
  DFFSSRX1_HVT conv1_weight_reg_15_ ( .D(1'b0), .SETB(n7700), .RSTB(
        sram_rdata_weight[15]), .CLK(clk), .Q(conv1_weight[15]) );
  DFFSSRX1_HVT weight_reg_15_ ( .D(1'b0), .SETB(n1510), .RSTB(conv1_weight[15]), .CLK(clk), .Q(weight[15]) );
  DFFSSRX1_HVT conv1_weight_reg_14_ ( .D(1'b0), .SETB(n1810), .RSTB(
        sram_rdata_weight[14]), .CLK(clk), .Q(conv1_weight[14]) );
  DFFSSRX1_HVT weight_reg_14_ ( .D(1'b0), .SETB(n1380), .RSTB(conv1_weight[14]), .CLK(clk), .Q(weight[14]) );
  DFFSSRX1_HVT conv1_weight_reg_13_ ( .D(1'b0), .SETB(n1750), .RSTB(
        sram_rdata_weight[13]), .CLK(clk), .Q(conv1_weight[13]) );
  DFFSSRX1_HVT weight_reg_13_ ( .D(1'b0), .SETB(n1520), .RSTB(conv1_weight[13]), .CLK(clk), .Q(weight[13]) );
  DFFSSRX1_HVT conv1_weight_reg_12_ ( .D(1'b0), .SETB(n1810), .RSTB(
        sram_rdata_weight[12]), .CLK(clk), .Q(conv1_weight[12]) );
  DFFSSRX1_HVT weight_reg_12_ ( .D(1'b0), .SETB(n13600), .RSTB(
        conv1_weight[12]), .CLK(clk), .Q(weight[12]) );
  DFFSSRX1_HVT conv1_weight_reg_11_ ( .D(1'b0), .SETB(n1530), .RSTB(
        sram_rdata_weight[11]), .CLK(clk), .Q(conv1_weight[11]) );
  DFFSSRX1_HVT weight_reg_11_ ( .D(1'b0), .SETB(n1810), .RSTB(conv1_weight[11]), .CLK(clk), .Q(weight[11]) );
  DFFSSRX1_HVT conv1_weight_reg_10_ ( .D(1'b0), .SETB(n1370), .RSTB(
        sram_rdata_weight[10]), .CLK(clk), .Q(conv1_weight[10]) );
  DFFSSRX1_HVT weight_reg_10_ ( .D(1'b0), .SETB(n34), .RSTB(conv1_weight[10]), 
        .CLK(clk), .Q(weight[10]) );
  DFFSSRX1_HVT conv1_weight_reg_9_ ( .D(1'b0), .SETB(n1510), .RSTB(
        sram_rdata_weight[9]), .CLK(clk), .Q(conv1_weight[9]) );
  DFFSSRX1_HVT weight_reg_9_ ( .D(1'b0), .SETB(n1810), .RSTB(conv1_weight[9]), 
        .CLK(clk), .Q(weight[9]) );
  DFFSSRX1_HVT conv1_weight_reg_8_ ( .D(1'b0), .SETB(n13500), .RSTB(
        sram_rdata_weight[8]), .CLK(clk), .Q(conv1_weight[8]) );
  DFFSSRX1_HVT weight_reg_8_ ( .D(1'b0), .SETB(n33), .RSTB(conv1_weight[8]), 
        .CLK(clk), .Q(weight[8]) );
  DFFSSRX1_HVT conv1_weight_reg_7_ ( .D(1'b0), .SETB(n1500), .RSTB(
        sram_rdata_weight[7]), .CLK(clk), .Q(conv1_weight[7]) );
  DFFSSRX1_HVT weight_reg_7_ ( .D(1'b0), .SETB(n1810), .RSTB(conv1_weight[7]), 
        .CLK(clk), .Q(weight[7]) );
  DFFSSRX1_HVT conv1_weight_reg_6_ ( .D(1'b0), .SETB(n13600), .RSTB(
        sram_rdata_weight[6]), .CLK(clk), .Q(conv1_weight[6]) );
  DFFSSRX1_HVT weight_reg_6_ ( .D(1'b0), .SETB(n33), .RSTB(conv1_weight[6]), 
        .CLK(clk), .Q(weight[6]) );
  DFFSSRX1_HVT conv1_weight_reg_5_ ( .D(1'b0), .SETB(n1530), .RSTB(
        sram_rdata_weight[5]), .CLK(clk), .Q(conv1_weight[5]) );
  DFFSSRX1_HVT weight_reg_5_ ( .D(1'b0), .SETB(n1810), .RSTB(conv1_weight[5]), 
        .CLK(clk), .Q(weight[5]) );
  DFFSSRX1_HVT conv1_weight_reg_4_ ( .D(1'b0), .SETB(n1370), .RSTB(
        sram_rdata_weight[4]), .CLK(clk), .Q(conv1_weight[4]) );
  DFFSSRX1_HVT weight_reg_4_ ( .D(1'b0), .SETB(n1750), .RSTB(conv1_weight[4]), 
        .CLK(clk), .Q(weight[4]) );
  DFFSSRX1_HVT conv1_weight_reg_3_ ( .D(1'b0), .SETB(n1510), .RSTB(
        sram_rdata_weight[3]), .CLK(clk), .Q(conv1_weight[3]) );
  DFFSSRX1_HVT weight_reg_3_ ( .D(1'b0), .SETB(n1780), .RSTB(conv1_weight[3]), 
        .CLK(clk), .Q(weight[3]) );
  DFFSSRX1_HVT conv1_weight_reg_2_ ( .D(1'b0), .SETB(n1380), .RSTB(
        sram_rdata_weight[2]), .CLK(clk), .Q(conv1_weight[2]) );
  DFFSSRX1_HVT weight_reg_2_ ( .D(1'b0), .SETB(n1520), .RSTB(conv1_weight[2]), 
        .CLK(clk), .Q(weight[2]) );
  DFFSSRX1_HVT conv1_weight_reg_1_ ( .D(1'b0), .SETB(n1780), .RSTB(
        sram_rdata_weight[1]), .CLK(clk), .Q(conv1_weight[1]) );
  DFFSSRX1_HVT weight_reg_1_ ( .D(1'b0), .SETB(n13500), .RSTB(conv1_weight[1]), 
        .CLK(clk), .Q(weight[1]) );
  DFFSSRX1_HVT conv1_weight_reg_0_ ( .D(1'b0), .SETB(n4800), .RSTB(
        sram_rdata_weight[0]), .CLK(clk), .Q(conv1_weight[0]) );
  DFFSSRX1_HVT weight_reg_0_ ( .D(1'b0), .SETB(n1530), .RSTB(conv1_weight[0]), 
        .CLK(clk), .Q(weight[0]) );
  DFFSSRX1_HVT sram_rdata_8_reg_31_ ( .D(1'b0), .SETB(n1780), .RSTB(N326), 
        .CLK(clk), .Q(sram_rdata_8[31]) );
  DFFSSRX1_HVT sram_rdata_8_reg_30_ ( .D(1'b0), .SETB(n1370), .RSTB(N325), 
        .CLK(clk), .Q(sram_rdata_8[30]) );
  DFFSSRX1_HVT sram_rdata_8_reg_29_ ( .D(1'b0), .SETB(n7800), .RSTB(N324), 
        .CLK(clk), .Q(sram_rdata_8[29]) );
  DFFSSRX1_HVT sram_rdata_8_reg_28_ ( .D(1'b0), .SETB(n1500), .RSTB(N323), 
        .CLK(clk), .Q(sram_rdata_8[28]) );
  DFFSSRX1_HVT sram_rdata_8_reg_27_ ( .D(1'b0), .SETB(n1780), .RSTB(N322), 
        .CLK(clk), .Q(sram_rdata_8[27]) );
  DFFSSRX1_HVT sram_rdata_8_reg_26_ ( .D(1'b0), .SETB(n13500), .RSTB(N321), 
        .CLK(clk), .Q(sram_rdata_8[26]) );
  DFFSSRX1_HVT sram_rdata_8_reg_25_ ( .D(1'b0), .SETB(n7800), .RSTB(N320), 
        .CLK(clk), .Q(sram_rdata_8[25]) );
  DFFSSRX1_HVT sram_rdata_8_reg_24_ ( .D(1'b0), .SETB(n1500), .RSTB(N319), 
        .CLK(clk), .Q(sram_rdata_8[24]) );
  DFFSSRX1_HVT sram_rdata_8_reg_23_ ( .D(1'b0), .SETB(n1780), .RSTB(N318), 
        .CLK(clk), .Q(sram_rdata_8[23]) );
  DFFSSRX1_HVT sram_rdata_8_reg_22_ ( .D(1'b0), .SETB(n1380), .RSTB(N317), 
        .CLK(clk), .Q(sram_rdata_8[22]) );
  DFFSSRX1_HVT sram_rdata_8_reg_21_ ( .D(1'b0), .SETB(n1530), .RSTB(N316), 
        .CLK(clk), .Q(sram_rdata_8[21]) );
  DFFSSRX1_HVT sram_rdata_8_reg_20_ ( .D(1'b0), .SETB(n1780), .RSTB(N315), 
        .CLK(clk), .Q(sram_rdata_8[20]) );
  DFFSSRX1_HVT sram_rdata_8_reg_19_ ( .D(1'b0), .SETB(n1370), .RSTB(N314), 
        .CLK(clk), .Q(sram_rdata_8[19]) );
  DFFSSRX1_HVT sram_rdata_8_reg_18_ ( .D(1'b0), .SETB(n1750), .RSTB(N313), 
        .CLK(clk), .Q(sram_rdata_8[18]) );
  DFFSSRX1_HVT sram_rdata_8_reg_17_ ( .D(1'b0), .SETB(n1520), .RSTB(N312), 
        .CLK(clk), .Q(sram_rdata_8[17]) );
  DFFSSRX1_HVT sram_rdata_8_reg_16_ ( .D(1'b0), .SETB(n1780), .RSTB(N311), 
        .CLK(clk), .Q(sram_rdata_8[16]) );
  DFFSSRX1_HVT sram_rdata_8_reg_15_ ( .D(1'b0), .SETB(n1380), .RSTB(N310), 
        .CLK(clk), .Q(sram_rdata_8[15]) );
  DFFSSRX1_HVT sram_rdata_8_reg_14_ ( .D(1'b0), .SETB(n34), .RSTB(N309), .CLK(
        clk), .Q(sram_rdata_8[14]) );
  DFFSSRX1_HVT sram_rdata_8_reg_13_ ( .D(1'b0), .SETB(n1520), .RSTB(N308), 
        .CLK(clk), .Q(sram_rdata_8[13]) );
  DFFSSRX1_HVT sram_rdata_8_reg_12_ ( .D(1'b0), .SETB(n1780), .RSTB(N307), 
        .CLK(clk), .Q(sram_rdata_8[12]) );
  DFFSSRX1_HVT sram_rdata_8_reg_11_ ( .D(1'b0), .SETB(n13500), .RSTB(N306), 
        .CLK(clk), .Q(sram_rdata_8[11]) );
  DFFSSRX1_HVT sram_rdata_8_reg_10_ ( .D(1'b0), .SETB(n4900), .RSTB(N305), 
        .CLK(clk), .Q(sram_rdata_8[10]) );
  DFFSSRX1_HVT sram_rdata_8_reg_9_ ( .D(1'b0), .SETB(n1530), .RSTB(N304), 
        .CLK(clk), .Q(sram_rdata_8[9]) );
  DFFSSRX1_HVT sram_rdata_8_reg_8_ ( .D(1'b0), .SETB(n1780), .RSTB(N303), 
        .CLK(clk), .Q(sram_rdata_8[8]) );
  DFFSSRX1_HVT sram_rdata_8_reg_7_ ( .D(1'b0), .SETB(n1370), .RSTB(N302), 
        .CLK(clk), .Q(sram_rdata_8[7]) );
  DFFSSRX1_HVT sram_rdata_8_reg_6_ ( .D(1'b0), .SETB(n4900), .RSTB(N301), 
        .CLK(clk), .Q(sram_rdata_8[6]) );
  DFFSSRX1_HVT sram_rdata_8_reg_5_ ( .D(1'b0), .SETB(n1500), .RSTB(N300), 
        .CLK(clk), .Q(sram_rdata_8[5]) );
  DFFSSRX1_HVT sram_rdata_8_reg_4_ ( .D(1'b0), .SETB(n1780), .RSTB(N299), 
        .CLK(clk), .Q(sram_rdata_8[4]) );
  DFFSSRX1_HVT sram_rdata_8_reg_3_ ( .D(1'b0), .SETB(n13500), .RSTB(N298), 
        .CLK(clk), .Q(sram_rdata_8[3]) );
  DFFSSRX1_HVT sram_rdata_8_reg_2_ ( .D(1'b0), .SETB(n1500), .RSTB(N297), 
        .CLK(clk), .Q(sram_rdata_8[2]) );
  DFFSSRX1_HVT sram_rdata_8_reg_1_ ( .D(1'b0), .SETB(n1780), .RSTB(N296), 
        .CLK(clk), .Q(sram_rdata_8[1]) );
  DFFSSRX1_HVT sram_rdata_8_reg_0_ ( .D(1'b0), .SETB(n1380), .RSTB(N295), 
        .CLK(clk), .Q(sram_rdata_8[0]) );
  DFFSSRX1_HVT sram_rdata_0_reg_31_ ( .D(1'b0), .SETB(n1750), .RSTB(N70), 
        .CLK(clk), .Q(sram_rdata_0[31]) );
  DFFSSRX1_HVT sram_rdata_0_reg_30_ ( .D(1'b0), .SETB(n1530), .RSTB(N69), 
        .CLK(clk), .Q(sram_rdata_0[30]) );
  DFFSSRX1_HVT sram_rdata_0_reg_29_ ( .D(1'b0), .SETB(n1780), .RSTB(N68), 
        .CLK(clk), .Q(sram_rdata_0[29]) );
  DFFSSRX1_HVT sram_rdata_0_reg_28_ ( .D(1'b0), .SETB(n1370), .RSTB(N67), 
        .CLK(clk), .Q(sram_rdata_0[28]) );
  DFFSSRX1_HVT sram_rdata_0_reg_27_ ( .D(1'b0), .SETB(n4800), .RSTB(N66), 
        .CLK(clk), .Q(sram_rdata_0[27]) );
  DFFSSRX1_HVT sram_rdata_0_reg_26_ ( .D(1'b0), .SETB(n1520), .RSTB(N65), 
        .CLK(clk), .Q(sram_rdata_0[26]) );
  DFFSSRX1_HVT sram_rdata_0_reg_25_ ( .D(1'b0), .SETB(n1780), .RSTB(N64), 
        .CLK(clk), .Q(sram_rdata_0[25]) );
  DFFSSRX1_HVT sram_rdata_0_reg_24_ ( .D(1'b0), .SETB(n1380), .RSTB(N63), 
        .CLK(clk), .Q(sram_rdata_0[24]) );
  DFFSSRX1_HVT sram_rdata_0_reg_23_ ( .D(1'b0), .SETB(n7900), .RSTB(N62), 
        .CLK(clk), .Q(sram_rdata_0[23]) );
  DFFSSRX1_HVT sram_rdata_0_reg_22_ ( .D(1'b0), .SETB(n1520), .RSTB(N61), 
        .CLK(clk), .Q(sram_rdata_0[22]) );
  DFFSSRX1_HVT sram_rdata_0_reg_21_ ( .D(1'b0), .SETB(n1780), .RSTB(N60), 
        .CLK(clk), .Q(sram_rdata_0[21]) );
  DFFSSRX1_HVT sram_rdata_0_reg_20_ ( .D(1'b0), .SETB(n13500), .RSTB(N59), 
        .CLK(clk), .Q(sram_rdata_0[20]) );
  DFFSSRX1_HVT sram_rdata_0_reg_19_ ( .D(1'b0), .SETB(n7900), .RSTB(N58), 
        .CLK(clk), .Q(sram_rdata_0[19]) );
  DFFSSRX1_HVT sram_rdata_0_reg_18_ ( .D(1'b0), .SETB(n1530), .RSTB(N57), 
        .CLK(clk), .Q(sram_rdata_0[18]) );
  DFFSSRX1_HVT sram_rdata_0_reg_17_ ( .D(1'b0), .SETB(n1780), .RSTB(N56), 
        .CLK(clk), .Q(sram_rdata_0[17]) );
  DFFSSRX1_HVT sram_rdata_0_reg_16_ ( .D(1'b0), .SETB(n1370), .RSTB(N55), 
        .CLK(clk), .Q(sram_rdata_0[16]) );
  DFFSSRX1_HVT sram_rdata_0_reg_15_ ( .D(1'b0), .SETB(n1500), .RSTB(N54), 
        .CLK(clk), .Q(sram_rdata_0[15]) );
  DFFSSRX1_HVT sram_rdata_0_reg_14_ ( .D(1'b0), .SETB(n1780), .RSTB(N53), 
        .CLK(clk), .Q(sram_rdata_0[14]) );
  DFFSSRX1_HVT sram_rdata_0_reg_13_ ( .D(1'b0), .SETB(n13500), .RSTB(N52), 
        .CLK(clk), .Q(sram_rdata_0[13]) );
  DFFSSRX1_HVT sram_rdata_0_reg_12_ ( .D(1'b0), .SETB(n1750), .RSTB(N51), 
        .CLK(clk), .Q(sram_rdata_0[12]) );
  DFFSSRX1_HVT sram_rdata_0_reg_11_ ( .D(1'b0), .SETB(n1500), .RSTB(N50), 
        .CLK(clk), .Q(sram_rdata_0[11]) );
  DFFSSRX1_HVT sram_rdata_0_reg_10_ ( .D(1'b0), .SETB(n1780), .RSTB(N49), 
        .CLK(clk), .Q(sram_rdata_0[10]) );
  DFFSSRX1_HVT sram_rdata_0_reg_9_ ( .D(1'b0), .SETB(n1380), .RSTB(N48), .CLK(
        clk), .Q(sram_rdata_0[9]) );
  DFFSSRX1_HVT sram_rdata_0_reg_8_ ( .D(1'b0), .SETB(n34), .RSTB(N47), .CLK(
        clk), .Q(sram_rdata_0[8]) );
  DFFSSRX1_HVT sram_rdata_0_reg_7_ ( .D(1'b0), .SETB(n1530), .RSTB(N46), .CLK(
        clk), .Q(sram_rdata_0[7]) );
  DFFSSRX1_HVT sram_rdata_0_reg_6_ ( .D(1'b0), .SETB(n1780), .RSTB(N45), .CLK(
        clk), .Q(sram_rdata_0[6]) );
  DFFSSRX1_HVT sram_rdata_0_reg_5_ ( .D(1'b0), .SETB(n1370), .RSTB(N44), .CLK(
        clk), .Q(sram_rdata_0[5]) );
  DFFSSRX1_HVT sram_rdata_0_reg_4_ ( .D(1'b0), .SETB(n4900), .RSTB(N43), .CLK(
        clk), .Q(sram_rdata_0[4]) );
  DFFSSRX1_HVT sram_rdata_0_reg_3_ ( .D(1'b0), .SETB(n1520), .RSTB(N42), .CLK(
        clk), .Q(sram_rdata_0[3]) );
  DFFSSRX1_HVT sram_rdata_0_reg_2_ ( .D(1'b0), .SETB(n1780), .RSTB(N41), .CLK(
        clk), .Q(sram_rdata_0[2]) );
  DFFSSRX1_HVT sram_rdata_0_reg_1_ ( .D(1'b0), .SETB(n1380), .RSTB(N40), .CLK(
        clk), .Q(sram_rdata_0[1]) );
  DFFSSRX1_HVT sram_rdata_0_reg_0_ ( .D(1'b0), .SETB(n1520), .RSTB(N39), .CLK(
        clk), .Q(sram_rdata_0[0]) );
  DFFSSRX1_HVT sram_rdata_1_reg_31_ ( .D(1'b0), .SETB(n1780), .RSTB(N102), 
        .CLK(clk), .Q(sram_rdata_1[31]) );
  DFFSSRX1_HVT sram_rdata_1_reg_30_ ( .D(1'b0), .SETB(n13500), .RSTB(N101), 
        .CLK(clk), .Q(sram_rdata_1[30]) );
  DFFSSRX1_HVT sram_rdata_1_reg_29_ ( .D(1'b0), .SETB(n4900), .RSTB(N100), 
        .CLK(clk), .Q(sram_rdata_1[29]) );
  DFFSSRX1_HVT sram_rdata_1_reg_28_ ( .D(1'b0), .SETB(n1530), .RSTB(N99), 
        .CLK(clk), .Q(sram_rdata_1[28]) );
  DFFSSRX1_HVT sram_rdata_1_reg_27_ ( .D(1'b0), .SETB(n1780), .RSTB(N98), 
        .CLK(clk), .Q(sram_rdata_1[27]) );
  DFFSSRX1_HVT sram_rdata_1_reg_26_ ( .D(1'b0), .SETB(n1370), .RSTB(N97), 
        .CLK(clk), .Q(sram_rdata_1[26]) );
  DFFSSRX1_HVT sram_rdata_1_reg_25_ ( .D(1'b0), .SETB(n1750), .RSTB(N96), 
        .CLK(clk), .Q(sram_rdata_1[25]) );
  DFFSSRX1_HVT sram_rdata_1_reg_24_ ( .D(1'b0), .SETB(n1500), .RSTB(N95), 
        .CLK(clk), .Q(sram_rdata_1[24]) );
  DFFSSRX1_HVT sram_rdata_1_reg_23_ ( .D(1'b0), .SETB(n1780), .RSTB(N94), 
        .CLK(clk), .Q(sram_rdata_1[23]) );
  DFFSSRX1_HVT sram_rdata_1_reg_22_ ( .D(1'b0), .SETB(n13600), .RSTB(N93), 
        .CLK(clk), .Q(sram_rdata_1[22]) );
  DFFSSRX1_HVT sram_rdata_1_reg_21_ ( .D(1'b0), .SETB(n4800), .RSTB(N92), 
        .CLK(clk), .Q(sram_rdata_1[21]) );
  DFFSSRX1_HVT sram_rdata_1_reg_20_ ( .D(1'b0), .SETB(n1510), .RSTB(N91), 
        .CLK(clk), .Q(sram_rdata_1[20]) );
  DFFSSRX1_HVT sram_rdata_1_reg_19_ ( .D(1'b0), .SETB(n1780), .RSTB(N90), 
        .CLK(clk), .Q(sram_rdata_1[19]) );
  DFFSSRX1_HVT sram_rdata_1_reg_18_ ( .D(1'b0), .SETB(n1380), .RSTB(N89), 
        .CLK(clk), .Q(sram_rdata_1[18]) );
  DFFSSRX1_HVT sram_rdata_1_reg_17_ ( .D(1'b0), .SETB(n777), .RSTB(N88), .CLK(
        clk), .Q(sram_rdata_1[17]) );
  DFFSSRX1_HVT sram_rdata_1_reg_16_ ( .D(1'b0), .SETB(n1530), .RSTB(N87), 
        .CLK(clk), .Q(sram_rdata_1[16]) );
  DFFSSRX1_HVT sram_rdata_1_reg_15_ ( .D(1'b0), .SETB(n1780), .RSTB(N86), 
        .CLK(clk), .Q(sram_rdata_1[15]) );
  DFFSSRX1_HVT sram_rdata_1_reg_14_ ( .D(1'b0), .SETB(n1370), .RSTB(N85), 
        .CLK(clk), .Q(sram_rdata_1[14]) );
  DFFSSRX1_HVT sram_rdata_1_reg_13_ ( .D(1'b0), .SETB(n1520), .RSTB(N84), 
        .CLK(clk), .Q(sram_rdata_1[13]) );
  DFFSSRX1_HVT sram_rdata_1_reg_12_ ( .D(1'b0), .SETB(n1780), .RSTB(N83), 
        .CLK(clk), .Q(sram_rdata_1[12]) );
  DFFSSRX1_HVT sram_rdata_1_reg_11_ ( .D(1'b0), .SETB(n13500), .RSTB(N82), 
        .CLK(clk), .Q(sram_rdata_1[11]) );
  DFFSSRX1_HVT sram_rdata_1_reg_10_ ( .D(1'b0), .SETB(n777), .RSTB(N81), .CLK(
        clk), .Q(sram_rdata_1[10]) );
  DFFSSRX1_HVT sram_rdata_1_reg_9_ ( .D(1'b0), .SETB(n1500), .RSTB(N80), .CLK(
        clk), .Q(sram_rdata_1[9]) );
  DFFSSRX1_HVT sram_rdata_1_reg_8_ ( .D(1'b0), .SETB(n1780), .RSTB(N79), .CLK(
        clk), .Q(sram_rdata_1[8]) );
  DFFSSRX1_HVT sram_rdata_1_reg_7_ ( .D(1'b0), .SETB(n13500), .RSTB(N78), 
        .CLK(clk), .Q(sram_rdata_1[7]) );
  DFFSSRX1_HVT sram_rdata_1_reg_6_ ( .D(1'b0), .SETB(n1750), .RSTB(N77), .CLK(
        clk), .Q(sram_rdata_1[6]) );
  DFFSSRX1_HVT sram_rdata_1_reg_5_ ( .D(1'b0), .SETB(n1530), .RSTB(N76), .CLK(
        clk), .Q(sram_rdata_1[5]) );
  DFFSSRX1_HVT sram_rdata_1_reg_4_ ( .D(1'b0), .SETB(n1790), .RSTB(N75), .CLK(
        clk), .Q(sram_rdata_1[4]) );
  DFFSSRX1_HVT sram_rdata_1_reg_3_ ( .D(1'b0), .SETB(n1370), .RSTB(N74), .CLK(
        clk), .Q(sram_rdata_1[3]) );
  DFFSSRX1_HVT sram_rdata_1_reg_2_ ( .D(1'b0), .SETB(n34), .RSTB(N73), .CLK(
        clk), .Q(sram_rdata_1[2]) );
  DFFSSRX1_HVT sram_rdata_1_reg_1_ ( .D(1'b0), .SETB(n1500), .RSTB(N72), .CLK(
        clk), .Q(sram_rdata_1[1]) );
  DFFSSRX1_HVT sram_rdata_1_reg_0_ ( .D(1'b0), .SETB(n1790), .RSTB(N71), .CLK(
        clk), .Q(sram_rdata_1[0]) );
  DFFSSRX1_HVT sram_rdata_2_reg_31_ ( .D(1'b0), .SETB(n1380), .RSTB(N134), 
        .CLK(clk), .Q(sram_rdata_2[31]) );
  DFFSSRX1_HVT sram_rdata_2_reg_30_ ( .D(1'b0), .SETB(n1520), .RSTB(N133), 
        .CLK(clk), .Q(sram_rdata_2[30]) );
  DFFSSRX1_HVT sram_rdata_2_reg_29_ ( .D(1'b0), .SETB(n1790), .RSTB(N132), 
        .CLK(clk), .Q(sram_rdata_2[29]) );
  DFFSSRX1_HVT sram_rdata_2_reg_28_ ( .D(1'b0), .SETB(n1380), .RSTB(N131), 
        .CLK(clk), .Q(sram_rdata_2[28]) );
  DFFSSRX1_HVT sram_rdata_2_reg_27_ ( .D(1'b0), .SETB(n33), .RSTB(N130), .CLK(
        clk), .Q(sram_rdata_2[27]) );
  DFFSSRX1_HVT sram_rdata_2_reg_26_ ( .D(1'b0), .SETB(n1530), .RSTB(N129), 
        .CLK(clk), .Q(sram_rdata_2[26]) );
  DFFSSRX1_HVT sram_rdata_2_reg_25_ ( .D(1'b0), .SETB(n1790), .RSTB(N128), 
        .CLK(clk), .Q(sram_rdata_2[25]) );
  DFFSSRX1_HVT sram_rdata_2_reg_24_ ( .D(1'b0), .SETB(n1370), .RSTB(N127), 
        .CLK(clk), .Q(sram_rdata_2[24]) );
  DFFSSRX1_HVT sram_rdata_2_reg_23_ ( .D(1'b0), .SETB(n33), .RSTB(N126), .CLK(
        clk), .Q(sram_rdata_2[23]) );
  DFFSSRX1_HVT sram_rdata_2_reg_22_ ( .D(1'b0), .SETB(n1520), .RSTB(N125), 
        .CLK(clk), .Q(sram_rdata_2[22]) );
  DFFSSRX1_HVT sram_rdata_2_reg_21_ ( .D(1'b0), .SETB(n1790), .RSTB(N124), 
        .CLK(clk), .Q(sram_rdata_2[21]) );
  DFFSSRX1_HVT sram_rdata_2_reg_20_ ( .D(1'b0), .SETB(n13500), .RSTB(N123), 
        .CLK(clk), .Q(sram_rdata_2[20]) );
  DFFSSRX1_HVT sram_rdata_2_reg_19_ ( .D(1'b0), .SETB(n1750), .RSTB(N122), 
        .CLK(clk), .Q(sram_rdata_2[19]) );
  DFFSSRX1_HVT sram_rdata_2_reg_18_ ( .D(1'b0), .SETB(n1500), .RSTB(N121), 
        .CLK(clk), .Q(sram_rdata_2[18]) );
  DFFSSRX1_HVT sram_rdata_2_reg_17_ ( .D(1'b0), .SETB(n1790), .RSTB(N120), 
        .CLK(clk), .Q(sram_rdata_2[17]) );
  DFFSSRX1_HVT sram_rdata_2_reg_16_ ( .D(1'b0), .SETB(n13600), .RSTB(N119), 
        .CLK(clk), .Q(sram_rdata_2[16]) );
  DFFSSRX1_HVT sram_rdata_2_reg_15_ ( .D(1'b0), .SETB(n4800), .RSTB(N118), 
        .CLK(clk), .Q(sram_rdata_2[15]) );
  DFFSSRX1_HVT sram_rdata_2_reg_14_ ( .D(1'b0), .SETB(n1530), .RSTB(N117), 
        .CLK(clk), .Q(sram_rdata_2[14]) );
  DFFSSRX1_HVT sram_rdata_2_reg_13_ ( .D(1'b0), .SETB(n1790), .RSTB(N116), 
        .CLK(clk), .Q(sram_rdata_2[13]) );
  DFFSSRX1_HVT sram_rdata_2_reg_12_ ( .D(1'b0), .SETB(n1370), .RSTB(N115), 
        .CLK(clk), .Q(sram_rdata_2[12]) );
  DFFSSRX1_HVT sram_rdata_2_reg_11_ ( .D(1'b0), .SETB(n1510), .RSTB(N114), 
        .CLK(clk), .Q(sram_rdata_2[11]) );
  DFFSSRX1_HVT sram_rdata_2_reg_10_ ( .D(1'b0), .SETB(n1790), .RSTB(N113), 
        .CLK(clk), .Q(sram_rdata_2[10]) );
  DFFSSRX1_HVT sram_rdata_2_reg_9_ ( .D(1'b0), .SETB(n1380), .RSTB(N112), 
        .CLK(clk), .Q(sram_rdata_2[9]) );
  DFFSSRX1_HVT sram_rdata_2_reg_8_ ( .D(1'b0), .SETB(n7700), .RSTB(N111), 
        .CLK(clk), .Q(sram_rdata_2[8]) );
  DFFSSRX1_HVT sram_rdata_2_reg_7_ ( .D(1'b0), .SETB(n1520), .RSTB(N110), 
        .CLK(clk), .Q(sram_rdata_2[7]) );
  DFFSSRX1_HVT sram_rdata_2_reg_6_ ( .D(1'b0), .SETB(n1790), .RSTB(N109), 
        .CLK(clk), .Q(sram_rdata_2[6]) );
  DFFSSRX1_HVT sram_rdata_2_reg_5_ ( .D(1'b0), .SETB(n13500), .RSTB(N108), 
        .CLK(clk), .Q(sram_rdata_2[5]) );
  DFFSSRX1_HVT sram_rdata_2_reg_4_ ( .D(1'b0), .SETB(n7700), .RSTB(N107), 
        .CLK(clk), .Q(sram_rdata_2[4]) );
  DFFSSRX1_HVT sram_rdata_2_reg_3_ ( .D(1'b0), .SETB(n1530), .RSTB(N106), 
        .CLK(clk), .Q(sram_rdata_2[3]) );
  DFFSSRX1_HVT sram_rdata_2_reg_2_ ( .D(1'b0), .SETB(n1790), .RSTB(N105), 
        .CLK(clk), .Q(sram_rdata_2[2]) );
  DFFSSRX1_HVT sram_rdata_2_reg_1_ ( .D(1'b0), .SETB(n1370), .RSTB(N104), 
        .CLK(clk), .Q(sram_rdata_2[1]) );
  DFFSSRX1_HVT sram_rdata_2_reg_0_ ( .D(1'b0), .SETB(n1750), .RSTB(N103), 
        .CLK(clk), .Q(sram_rdata_2[0]) );
  DFFSSRX1_HVT sram_rdata_3_reg_31_ ( .D(1'b0), .SETB(n1500), .RSTB(N166), 
        .CLK(clk), .Q(sram_rdata_3[31]) );
  DFFSSRX1_HVT sram_rdata_3_reg_30_ ( .D(1'b0), .SETB(n1790), .RSTB(N165), 
        .CLK(clk), .Q(sram_rdata_3[30]) );
  DFFSSRX1_HVT sram_rdata_3_reg_29_ ( .D(1'b0), .SETB(n13500), .RSTB(N164), 
        .CLK(clk), .Q(sram_rdata_3[29]) );
  DFFSSRX1_HVT sram_rdata_3_reg_28_ ( .D(1'b0), .SETB(n34), .RSTB(N163), .CLK(
        clk), .Q(sram_rdata_3[28]) );
  DFFSSRX1_HVT sram_rdata_3_reg_27_ ( .D(1'b0), .SETB(n1500), .RSTB(N162), 
        .CLK(clk), .Q(sram_rdata_3[27]) );
  DFFSSRX1_HVT sram_rdata_3_reg_26_ ( .D(1'b0), .SETB(n1790), .RSTB(N161), 
        .CLK(clk), .Q(sram_rdata_3[26]) );
  DFFSSRX1_HVT sram_rdata_3_reg_25_ ( .D(1'b0), .SETB(n1380), .RSTB(N160), 
        .CLK(clk), .Q(sram_rdata_3[25]) );
  DFFSSRX1_HVT sram_rdata_3_reg_24_ ( .D(1'b0), .SETB(n1530), .RSTB(N159), 
        .CLK(clk), .Q(sram_rdata_3[24]) );
  DFFSSRX1_HVT sram_rdata_3_reg_23_ ( .D(1'b0), .SETB(n1790), .RSTB(N158), 
        .CLK(clk), .Q(sram_rdata_3[23]) );
  DFFSSRX1_HVT sram_rdata_3_reg_22_ ( .D(1'b0), .SETB(n1370), .RSTB(N157), 
        .CLK(clk), .Q(sram_rdata_3[22]) );
  DFFSSRX1_HVT sram_rdata_3_reg_21_ ( .D(1'b0), .SETB(n33), .RSTB(N156), .CLK(
        clk), .Q(sram_rdata_3[21]) );
  DFFSSRX1_HVT sram_rdata_3_reg_20_ ( .D(1'b0), .SETB(n1520), .RSTB(N155), 
        .CLK(clk), .Q(sram_rdata_3[20]) );
  DFFSSRX1_HVT sram_rdata_3_reg_19_ ( .D(1'b0), .SETB(n1790), .RSTB(N154), 
        .CLK(clk), .Q(sram_rdata_3[19]) );
  DFFSSRX1_HVT sram_rdata_3_reg_18_ ( .D(1'b0), .SETB(n1380), .RSTB(N153), 
        .CLK(clk), .Q(sram_rdata_3[18]) );
  DFFSSRX1_HVT sram_rdata_3_reg_17_ ( .D(1'b0), .SETB(n33), .RSTB(N152), .CLK(
        clk), .Q(sram_rdata_3[17]) );
  DFFSSRX1_HVT sram_rdata_3_reg_16_ ( .D(1'b0), .SETB(n1520), .RSTB(N151), 
        .CLK(clk), .Q(sram_rdata_3[16]) );
  DFFSSRX1_HVT sram_rdata_3_reg_15_ ( .D(1'b0), .SETB(n1790), .RSTB(N150), 
        .CLK(clk), .Q(sram_rdata_3[15]) );
  DFFSSRX1_HVT sram_rdata_3_reg_14_ ( .D(1'b0), .SETB(n13500), .RSTB(N149), 
        .CLK(clk), .Q(sram_rdata_3[14]) );
  DFFSSRX1_HVT sram_rdata_3_reg_13_ ( .D(1'b0), .SETB(n1750), .RSTB(N148), 
        .CLK(clk), .Q(sram_rdata_3[13]) );
  DFFSSRX1_HVT sram_rdata_3_reg_12_ ( .D(1'b0), .SETB(n1530), .RSTB(N147), 
        .CLK(clk), .Q(sram_rdata_3[12]) );
  DFFSSRX1_HVT sram_rdata_3_reg_11_ ( .D(1'b0), .SETB(n1790), .RSTB(N146), 
        .CLK(clk), .Q(sram_rdata_3[11]) );
  DFFSSRX1_HVT sram_rdata_3_reg_10_ ( .D(1'b0), .SETB(n1370), .RSTB(N145), 
        .CLK(clk), .Q(sram_rdata_3[10]) );
  DFFSSRX1_HVT sram_rdata_3_reg_9_ ( .D(1'b0), .SETB(n1500), .RSTB(N144), 
        .CLK(clk), .Q(sram_rdata_3[9]) );
  DFFSSRX1_HVT sram_rdata_3_reg_8_ ( .D(1'b0), .SETB(n1790), .RSTB(N143), 
        .CLK(clk), .Q(sram_rdata_3[8]) );
  DFFSSRX1_HVT sram_rdata_3_reg_7_ ( .D(1'b0), .SETB(n13500), .RSTB(N142), 
        .CLK(clk), .Q(sram_rdata_3[7]) );
  DFFSSRX1_HVT sram_rdata_3_reg_6_ ( .D(1'b0), .SETB(n4800), .RSTB(N141), 
        .CLK(clk), .Q(sram_rdata_3[6]) );
  DFFSSRX1_HVT sram_rdata_3_reg_5_ ( .D(1'b0), .SETB(n1500), .RSTB(N140), 
        .CLK(clk), .Q(sram_rdata_3[5]) );
  DFFSSRX1_HVT sram_rdata_3_reg_4_ ( .D(1'b0), .SETB(n1790), .RSTB(N139), 
        .CLK(clk), .Q(sram_rdata_3[4]) );
  DFFSSRX1_HVT sram_rdata_3_reg_3_ ( .D(1'b0), .SETB(n1380), .RSTB(N138), 
        .CLK(clk), .Q(sram_rdata_3[3]) );
  DFFSSRX1_HVT sram_rdata_3_reg_2_ ( .D(1'b0), .SETB(n7800), .RSTB(N137), 
        .CLK(clk), .Q(sram_rdata_3[2]) );
  DFFSSRX1_HVT sram_rdata_3_reg_1_ ( .D(1'b0), .SETB(n1530), .RSTB(N136), 
        .CLK(clk), .Q(sram_rdata_3[1]) );
  DFFSSRX1_HVT sram_rdata_3_reg_0_ ( .D(1'b0), .SETB(n1790), .RSTB(N135), 
        .CLK(clk), .Q(sram_rdata_3[0]) );
  DFFSSRX1_HVT sram_rdata_4_reg_31_ ( .D(1'b0), .SETB(n1370), .RSTB(N198), 
        .CLK(clk), .Q(sram_rdata_4[31]) );
  DFFSSRX1_HVT sram_rdata_4_reg_30_ ( .D(1'b0), .SETB(n7800), .RSTB(N197), 
        .CLK(clk), .Q(sram_rdata_4[30]) );
  DFFSSRX1_HVT sram_rdata_4_reg_29_ ( .D(1'b0), .SETB(n1520), .RSTB(N196), 
        .CLK(clk), .Q(sram_rdata_4[29]) );
  DFFSSRX1_HVT sram_rdata_4_reg_28_ ( .D(1'b0), .SETB(n1790), .RSTB(N195), 
        .CLK(clk), .Q(sram_rdata_4[28]) );
  DFFSSRX1_HVT sram_rdata_4_reg_27_ ( .D(1'b0), .SETB(n1380), .RSTB(N194), 
        .CLK(clk), .Q(sram_rdata_4[27]) );
  DFFSSRX1_HVT sram_rdata_4_reg_26_ ( .D(1'b0), .SETB(n1750), .RSTB(N193), 
        .CLK(clk), .Q(sram_rdata_4[26]) );
  DFFSSRX1_HVT sram_rdata_4_reg_25_ ( .D(1'b0), .SETB(n1520), .RSTB(N192), 
        .CLK(clk), .Q(sram_rdata_4[25]) );
  DFFSSRX1_HVT sram_rdata_4_reg_24_ ( .D(1'b0), .SETB(n1790), .RSTB(N191), 
        .CLK(clk), .Q(sram_rdata_4[24]) );
  DFFSSRX1_HVT sram_rdata_4_reg_23_ ( .D(1'b0), .SETB(n13500), .RSTB(N190), 
        .CLK(clk), .Q(sram_rdata_4[23]) );
  DFFSSRX1_HVT sram_rdata_4_reg_22_ ( .D(1'b0), .SETB(n1530), .RSTB(N189), 
        .CLK(clk), .Q(sram_rdata_4[22]) );
  DFFSSRX1_HVT sram_rdata_4_reg_21_ ( .D(1'b0), .SETB(n1790), .RSTB(N188), 
        .CLK(clk), .Q(sram_rdata_4[21]) );
  DFFSSRX1_HVT sram_rdata_4_reg_20_ ( .D(1'b0), .SETB(n1370), .RSTB(N187), 
        .CLK(clk), .Q(sram_rdata_4[20]) );
  DFFSSRX1_HVT sram_rdata_4_reg_19_ ( .D(1'b0), .SETB(n34), .RSTB(N186), .CLK(
        clk), .Q(sram_rdata_4[19]) );
  DFFSSRX1_HVT sram_rdata_4_reg_18_ ( .D(1'b0), .SETB(n1500), .RSTB(N185), 
        .CLK(clk), .Q(sram_rdata_4[18]) );
  DFFSSRX1_HVT sram_rdata_4_reg_17_ ( .D(1'b0), .SETB(n1790), .RSTB(N184), 
        .CLK(clk), .Q(sram_rdata_4[17]) );
  DFFSSRX1_HVT sram_rdata_4_reg_16_ ( .D(1'b0), .SETB(n13500), .RSTB(N183), 
        .CLK(clk), .Q(sram_rdata_4[16]) );
  DFFSSRX1_HVT sram_rdata_4_reg_15_ ( .D(1'b0), .SETB(n4900), .RSTB(N182), 
        .CLK(clk), .Q(sram_rdata_4[15]) );
  DFFSSRX1_HVT sram_rdata_4_reg_14_ ( .D(1'b0), .SETB(n1500), .RSTB(N181), 
        .CLK(clk), .Q(sram_rdata_4[14]) );
  DFFSSRX1_HVT sram_rdata_4_reg_13_ ( .D(1'b0), .SETB(n1790), .RSTB(N180), 
        .CLK(clk), .Q(sram_rdata_4[13]) );
  DFFSSRX1_HVT sram_rdata_4_reg_12_ ( .D(1'b0), .SETB(n1380), .RSTB(N179), 
        .CLK(clk), .Q(sram_rdata_4[12]) );
  DFFSSRX1_HVT sram_rdata_4_reg_11_ ( .D(1'b0), .SETB(n4900), .RSTB(N178), 
        .CLK(clk), .Q(sram_rdata_4[11]) );
  DFFSSRX1_HVT sram_rdata_4_reg_10_ ( .D(1'b0), .SETB(n1530), .RSTB(N177), 
        .CLK(clk), .Q(sram_rdata_4[10]) );
  DFFSSRX1_HVT sram_rdata_4_reg_9_ ( .D(1'b0), .SETB(n1790), .RSTB(N176), 
        .CLK(clk), .Q(sram_rdata_4[9]) );
  DFFSSRX1_HVT sram_rdata_4_reg_8_ ( .D(1'b0), .SETB(n1370), .RSTB(N175), 
        .CLK(clk), .Q(sram_rdata_4[8]) );
  DFFSSRX1_HVT sram_rdata_4_reg_7_ ( .D(1'b0), .SETB(n1520), .RSTB(N174), 
        .CLK(clk), .Q(sram_rdata_4[7]) );
  DFFSSRX1_HVT sram_rdata_4_reg_6_ ( .D(1'b0), .SETB(n1800), .RSTB(N173), 
        .CLK(clk), .Q(sram_rdata_4[6]) );
  DFFSSRX1_HVT sram_rdata_4_reg_5_ ( .D(1'b0), .SETB(n1380), .RSTB(N172), 
        .CLK(clk), .Q(sram_rdata_4[5]) );
  DFFSSRX1_HVT sram_rdata_4_reg_4_ ( .D(1'b0), .SETB(n1750), .RSTB(N171), 
        .CLK(clk), .Q(sram_rdata_4[4]) );
  DFFSSRX1_HVT sram_rdata_4_reg_3_ ( .D(1'b0), .SETB(n1520), .RSTB(N170), 
        .CLK(clk), .Q(sram_rdata_4[3]) );
  DFFSSRX1_HVT sram_rdata_4_reg_2_ ( .D(1'b0), .SETB(n1800), .RSTB(N169), 
        .CLK(clk), .Q(sram_rdata_4[2]) );
  DFFSSRX1_HVT sram_rdata_4_reg_1_ ( .D(1'b0), .SETB(n13500), .RSTB(N168), 
        .CLK(clk), .Q(sram_rdata_4[1]) );
  DFFSSRX1_HVT sram_rdata_4_reg_0_ ( .D(1'b0), .SETB(n4800), .RSTB(N167), 
        .CLK(clk), .Q(sram_rdata_4[0]) );
  DFFSSRX1_HVT sram_rdata_5_reg_31_ ( .D(1'b0), .SETB(n1530), .RSTB(N230), 
        .CLK(clk), .Q(sram_rdata_5[31]) );
  DFFSSRX1_HVT sram_rdata_5_reg_30_ ( .D(1'b0), .SETB(n1800), .RSTB(N229), 
        .CLK(clk), .Q(sram_rdata_5[30]) );
  DFFSSRX1_HVT sram_rdata_5_reg_29_ ( .D(1'b0), .SETB(n1370), .RSTB(N228), 
        .CLK(clk), .Q(sram_rdata_5[29]) );
  DFFSSRX1_HVT sram_rdata_5_reg_28_ ( .D(1'b0), .SETB(n7900), .RSTB(N227), 
        .CLK(clk), .Q(sram_rdata_5[28]) );
  DFFSSRX1_HVT sram_rdata_5_reg_27_ ( .D(1'b0), .SETB(n1500), .RSTB(N226), 
        .CLK(clk), .Q(sram_rdata_5[27]) );
  DFFSSRX1_HVT sram_rdata_5_reg_26_ ( .D(1'b0), .SETB(n1800), .RSTB(N225), 
        .CLK(clk), .Q(sram_rdata_5[26]) );
  DFFSSRX1_HVT sram_rdata_5_reg_25_ ( .D(1'b0), .SETB(n13500), .RSTB(N224), 
        .CLK(clk), .Q(sram_rdata_5[25]) );
  DFFSSRX1_HVT sram_rdata_5_reg_24_ ( .D(1'b0), .SETB(n7900), .RSTB(N223), 
        .CLK(clk), .Q(sram_rdata_5[24]) );
  DFFSSRX1_HVT sram_rdata_5_reg_23_ ( .D(1'b0), .SETB(n1500), .RSTB(N222), 
        .CLK(clk), .Q(sram_rdata_5[23]) );
  DFFSSRX1_HVT sram_rdata_5_reg_22_ ( .D(1'b0), .SETB(n1800), .RSTB(N221), 
        .CLK(clk), .Q(sram_rdata_5[22]) );
  DFFSSRX1_HVT sram_rdata_5_reg_21_ ( .D(1'b0), .SETB(n1380), .RSTB(N220), 
        .CLK(clk), .Q(sram_rdata_5[21]) );
  DFFSSRX1_HVT sram_rdata_5_reg_20_ ( .D(1'b0), .SETB(n1530), .RSTB(N219), 
        .CLK(clk), .Q(sram_rdata_5[20]) );
  DFFSSRX1_HVT sram_rdata_5_reg_19_ ( .D(1'b0), .SETB(n1800), .RSTB(N218), 
        .CLK(clk), .Q(sram_rdata_5[19]) );
  DFFSSRX1_HVT sram_rdata_5_reg_18_ ( .D(1'b0), .SETB(n1370), .RSTB(N217), 
        .CLK(clk), .Q(sram_rdata_5[18]) );
  DFFSSRX1_HVT sram_rdata_5_reg_17_ ( .D(1'b0), .SETB(n1750), .RSTB(N216), 
        .CLK(clk), .Q(sram_rdata_5[17]) );
  DFFSSRX1_HVT sram_rdata_5_reg_16_ ( .D(1'b0), .SETB(n1520), .RSTB(N215), 
        .CLK(clk), .Q(sram_rdata_5[16]) );
  DFFSSRX1_HVT sram_rdata_5_reg_15_ ( .D(1'b0), .SETB(n1800), .RSTB(N214), 
        .CLK(clk), .Q(sram_rdata_5[15]) );
  DFFSSRX1_HVT sram_rdata_5_reg_14_ ( .D(1'b0), .SETB(n1380), .RSTB(N213), 
        .CLK(clk), .Q(sram_rdata_5[14]) );
  DFFSSRX1_HVT sram_rdata_5_reg_13_ ( .D(1'b0), .SETB(n34), .RSTB(N212), .CLK(
        clk), .Q(sram_rdata_5[13]) );
  DFFSSRX1_HVT sram_rdata_5_reg_12_ ( .D(1'b0), .SETB(n1520), .RSTB(N211), 
        .CLK(clk), .Q(sram_rdata_5[12]) );
  DFFSSRX1_HVT sram_rdata_5_reg_11_ ( .D(1'b0), .SETB(n1800), .RSTB(N210), 
        .CLK(clk), .Q(sram_rdata_5[11]) );
  DFFSSRX1_HVT sram_rdata_5_reg_10_ ( .D(1'b0), .SETB(n13500), .RSTB(N209), 
        .CLK(clk), .Q(sram_rdata_5[10]) );
  DFFSSRX1_HVT sram_rdata_5_reg_9_ ( .D(1'b0), .SETB(n4900), .RSTB(N208), 
        .CLK(clk), .Q(sram_rdata_5[9]) );
  DFFSSRX1_HVT sram_rdata_5_reg_8_ ( .D(1'b0), .SETB(n1530), .RSTB(N207), 
        .CLK(clk), .Q(sram_rdata_5[8]) );
  DFFSSRX1_HVT sram_rdata_5_reg_7_ ( .D(1'b0), .SETB(n1800), .RSTB(N206), 
        .CLK(clk), .Q(sram_rdata_5[7]) );
  DFFSSRX1_HVT sram_rdata_5_reg_6_ ( .D(1'b0), .SETB(n13600), .RSTB(N205), 
        .CLK(clk), .Q(sram_rdata_5[6]) );
  DFFSSRX1_HVT sram_rdata_5_reg_5_ ( .D(1'b0), .SETB(n1760), .RSTB(N204), 
        .CLK(clk), .Q(sram_rdata_5[5]) );
  DFFSSRX1_HVT sram_rdata_5_reg_4_ ( .D(1'b0), .SETB(n1500), .RSTB(N203), 
        .CLK(clk), .Q(sram_rdata_5[4]) );
  DFFSSRX1_HVT sram_rdata_5_reg_3_ ( .D(1'b0), .SETB(n1800), .RSTB(N202), 
        .CLK(clk), .Q(sram_rdata_5[3]) );
  DFFSSRX1_HVT sram_rdata_5_reg_2_ ( .D(1'b0), .SETB(n13500), .RSTB(N201), 
        .CLK(clk), .Q(sram_rdata_5[2]) );
  DFFSSRX1_HVT sram_rdata_5_reg_1_ ( .D(1'b0), .SETB(n1500), .RSTB(N200), 
        .CLK(clk), .Q(sram_rdata_5[1]) );
  DFFSSRX1_HVT sram_rdata_5_reg_0_ ( .D(1'b0), .SETB(n1800), .RSTB(N199), 
        .CLK(clk), .Q(sram_rdata_5[0]) );
  DFFSSRX1_HVT sram_rdata_6_reg_31_ ( .D(1'b0), .SETB(n1380), .RSTB(N262), 
        .CLK(clk), .Q(sram_rdata_6[31]) );
  DFFSSRX1_HVT sram_rdata_6_reg_30_ ( .D(1'b0), .SETB(n1750), .RSTB(N261), 
        .CLK(clk), .Q(sram_rdata_6[30]) );
  DFFSSRX1_HVT sram_rdata_6_reg_29_ ( .D(1'b0), .SETB(n1510), .RSTB(N260), 
        .CLK(clk), .Q(sram_rdata_6[29]) );
  DFFSSRX1_HVT sram_rdata_6_reg_28_ ( .D(1'b0), .SETB(n1800), .RSTB(N259), 
        .CLK(clk), .Q(sram_rdata_6[28]) );
  DFFSSRX1_HVT sram_rdata_6_reg_27_ ( .D(1'b0), .SETB(n13600), .RSTB(N258), 
        .CLK(clk), .Q(sram_rdata_6[27]) );
  DFFSSRX1_HVT sram_rdata_6_reg_26_ ( .D(1'b0), .SETB(n4800), .RSTB(N257), 
        .CLK(clk), .Q(sram_rdata_6[26]) );
  DFFSSRX1_HVT sram_rdata_6_reg_25_ ( .D(1'b0), .SETB(n1520), .RSTB(N256), 
        .CLK(clk), .Q(sram_rdata_6[25]) );
  DFFSSRX1_HVT sram_rdata_6_reg_24_ ( .D(1'b0), .SETB(n1800), .RSTB(N255), 
        .CLK(clk), .Q(sram_rdata_6[24]) );
  DFFSSRX1_HVT sram_rdata_6_reg_23_ ( .D(1'b0), .SETB(n1380), .RSTB(N254), 
        .CLK(clk), .Q(sram_rdata_6[23]) );
  DFFSSRX1_HVT sram_rdata_6_reg_22_ ( .D(1'b0), .SETB(n777), .RSTB(N253), 
        .CLK(clk), .Q(sram_rdata_6[22]) );
  DFFSSRX1_HVT sram_rdata_6_reg_21_ ( .D(1'b0), .SETB(n1520), .RSTB(N252), 
        .CLK(clk), .Q(sram_rdata_6[21]) );
  DFFSSRX1_HVT sram_rdata_6_reg_20_ ( .D(1'b0), .SETB(n1800), .RSTB(N251), 
        .CLK(clk), .Q(sram_rdata_6[20]) );
  DFFSSRX1_HVT sram_rdata_6_reg_19_ ( .D(1'b0), .SETB(n13500), .RSTB(N250), 
        .CLK(clk), .Q(sram_rdata_6[19]) );
  DFFSSRX1_HVT sram_rdata_6_reg_18_ ( .D(1'b0), .SETB(n1510), .RSTB(N249), 
        .CLK(clk), .Q(sram_rdata_6[18]) );
  DFFSSRX1_HVT sram_rdata_6_reg_17_ ( .D(1'b0), .SETB(n1800), .RSTB(N248), 
        .CLK(clk), .Q(sram_rdata_6[17]) );
  DFFSSRX1_HVT sram_rdata_6_reg_16_ ( .D(1'b0), .SETB(n13600), .RSTB(N247), 
        .CLK(clk), .Q(sram_rdata_6[16]) );
  DFFSSRX1_HVT sram_rdata_6_reg_15_ ( .D(1'b0), .SETB(n1760), .RSTB(N246), 
        .CLK(clk), .Q(sram_rdata_6[15]) );
  DFFSSRX1_HVT sram_rdata_6_reg_14_ ( .D(1'b0), .SETB(n1500), .RSTB(N245), 
        .CLK(clk), .Q(sram_rdata_6[14]) );
  DFFSSRX1_HVT sram_rdata_6_reg_13_ ( .D(1'b0), .SETB(n1800), .RSTB(N244), 
        .CLK(clk), .Q(sram_rdata_6[13]) );
  DFFSSRX1_HVT sram_rdata_6_reg_12_ ( .D(1'b0), .SETB(n13500), .RSTB(N243), 
        .CLK(clk), .Q(sram_rdata_6[12]) );
  DFFSSRX1_HVT sram_rdata_6_reg_11_ ( .D(1'b0), .SETB(n4900), .RSTB(N242), 
        .CLK(clk), .Q(sram_rdata_6[11]) );
  DFFSSRX1_HVT sram_rdata_6_reg_10_ ( .D(1'b0), .SETB(n1500), .RSTB(N241), 
        .CLK(clk), .Q(sram_rdata_6[10]) );
  DFFSSRX1_HVT sram_rdata_6_reg_9_ ( .D(1'b0), .SETB(n1800), .RSTB(N240), 
        .CLK(clk), .Q(sram_rdata_6[9]) );
  DFFSSRX1_HVT sram_rdata_6_reg_8_ ( .D(1'b0), .SETB(n1380), .RSTB(N239), 
        .CLK(clk), .Q(sram_rdata_6[8]) );
  DFFSSRX1_HVT sram_rdata_6_reg_7_ ( .D(1'b0), .SETB(n34), .RSTB(N238), .CLK(
        clk), .Q(sram_rdata_6[7]) );
  DFFSSRX1_HVT sram_rdata_6_reg_6_ ( .D(1'b0), .SETB(n1510), .RSTB(N237), 
        .CLK(clk), .Q(sram_rdata_6[6]) );
  DFFSSRX1_HVT sram_rdata_6_reg_5_ ( .D(1'b0), .SETB(n1800), .RSTB(N236), 
        .CLK(clk), .Q(sram_rdata_6[5]) );
  DFFSSRX1_HVT sram_rdata_6_reg_4_ ( .D(1'b0), .SETB(n13600), .RSTB(N235), 
        .CLK(clk), .Q(sram_rdata_6[4]) );
  DFFSSRX1_HVT sram_rdata_6_reg_3_ ( .D(1'b0), .SETB(n33), .RSTB(N234), .CLK(
        clk), .Q(sram_rdata_6[3]) );
  DFFSSRX1_HVT sram_rdata_6_reg_2_ ( .D(1'b0), .SETB(n1520), .RSTB(N233), 
        .CLK(clk), .Q(sram_rdata_6[2]) );
  DFFSSRX1_HVT sram_rdata_6_reg_1_ ( .D(1'b0), .SETB(n1800), .RSTB(N232), 
        .CLK(clk), .Q(sram_rdata_6[1]) );
  DFFSSRX1_HVT sram_rdata_6_reg_0_ ( .D(1'b0), .SETB(n1380), .RSTB(N231), 
        .CLK(clk), .Q(sram_rdata_6[0]) );
  DFFSSRX1_HVT sram_rdata_7_reg_31_ ( .D(1'b0), .SETB(n1520), .RSTB(N294), 
        .CLK(clk), .Q(sram_rdata_7[31]) );
  DFFSSRX1_HVT sram_rdata_7_reg_30_ ( .D(1'b0), .SETB(n1800), .RSTB(N293), 
        .CLK(clk), .Q(sram_rdata_7[30]) );
  DFFSSRX1_HVT sram_rdata_7_reg_29_ ( .D(1'b0), .SETB(n13500), .RSTB(N292), 
        .CLK(clk), .Q(sram_rdata_7[29]) );
  DFFSSRX1_HVT sram_rdata_7_reg_28_ ( .D(1'b0), .SETB(n1760), .RSTB(N291), 
        .CLK(clk), .Q(sram_rdata_7[28]) );
  DFFSSRX1_HVT sram_rdata_7_reg_27_ ( .D(1'b0), .SETB(n1510), .RSTB(N290), 
        .CLK(clk), .Q(sram_rdata_7[27]) );
  DFFSSRX1_HVT sram_rdata_7_reg_26_ ( .D(1'b0), .SETB(n1800), .RSTB(N289), 
        .CLK(clk), .Q(sram_rdata_7[26]) );
  DFFSSRX1_HVT sram_rdata_7_reg_25_ ( .D(1'b0), .SETB(n13600), .RSTB(N288), 
        .CLK(clk), .Q(sram_rdata_7[25]) );
  DFFSSRX1_HVT sram_rdata_7_reg_24_ ( .D(1'b0), .SETB(n7800), .RSTB(N287), 
        .CLK(clk), .Q(sram_rdata_7[24]) );
  DFFSSRX1_HVT sram_rdata_7_reg_23_ ( .D(1'b0), .SETB(n1500), .RSTB(N286), 
        .CLK(clk), .Q(sram_rdata_7[23]) );
  DFFSSRX1_HVT sram_rdata_7_reg_22_ ( .D(1'b0), .SETB(n1800), .RSTB(N285), 
        .CLK(clk), .Q(sram_rdata_7[22]) );
  DFFSSRX1_HVT sram_rdata_7_reg_21_ ( .D(1'b0), .SETB(n13500), .RSTB(N284), 
        .CLK(clk), .Q(sram_rdata_7[21]) );
  DFFSSRX1_HVT sram_rdata_7_reg_20_ ( .D(1'b0), .SETB(n4800), .RSTB(N283), 
        .CLK(clk), .Q(sram_rdata_7[20]) );
  DFFSSRX1_HVT sram_rdata_7_reg_19_ ( .D(1'b0), .SETB(n1500), .RSTB(N282), 
        .CLK(clk), .Q(sram_rdata_7[19]) );
  DFFSSRX1_HVT sram_rdata_7_reg_18_ ( .D(1'b0), .SETB(n1800), .RSTB(N281), 
        .CLK(clk), .Q(sram_rdata_7[18]) );
  DFFSSRX1_HVT sram_rdata_7_reg_17_ ( .D(1'b0), .SETB(n1380), .RSTB(N280), 
        .CLK(clk), .Q(sram_rdata_7[17]) );
  DFFSSRX1_HVT sram_rdata_7_reg_16_ ( .D(1'b0), .SETB(n1510), .RSTB(N279), 
        .CLK(clk), .Q(sram_rdata_7[16]) );
  DFFSSRX1_HVT sram_rdata_7_reg_15_ ( .D(1'b0), .SETB(n1800), .RSTB(N278), 
        .CLK(clk), .Q(sram_rdata_7[15]) );
  DFFSSRX1_HVT sram_rdata_7_reg_14_ ( .D(1'b0), .SETB(n13600), .RSTB(N277), 
        .CLK(clk), .Q(sram_rdata_7[14]) );
  DFFSSRX1_HVT sram_rdata_7_reg_13_ ( .D(1'b0), .SETB(n7700), .RSTB(N276), 
        .CLK(clk), .Q(sram_rdata_7[13]) );
  DFFSSRX1_HVT sram_rdata_7_reg_12_ ( .D(1'b0), .SETB(n1520), .RSTB(N275), 
        .CLK(clk), .Q(sram_rdata_7[12]) );
  DFFSSRX1_HVT sram_rdata_7_reg_11_ ( .D(1'b0), .SETB(n1800), .RSTB(N274), 
        .CLK(clk), .Q(sram_rdata_7[11]) );
  DFFSSRX1_HVT sram_rdata_7_reg_10_ ( .D(1'b0), .SETB(n1380), .RSTB(N273), 
        .CLK(clk), .Q(sram_rdata_7[10]) );
  DFFSSRX1_HVT sram_rdata_7_reg_9_ ( .D(1'b0), .SETB(n1760), .RSTB(N272), 
        .CLK(clk), .Q(sram_rdata_7[9]) );
  DFFSSRX1_HVT sram_rdata_7_reg_8_ ( .D(1'b0), .SETB(n1520), .RSTB(N271), 
        .CLK(clk), .Q(sram_rdata_7[8]) );
  DFFSSRX1_HVT sram_rdata_7_reg_7_ ( .D(1'b0), .SETB(n1800), .RSTB(N270), 
        .CLK(clk), .Q(sram_rdata_7[7]) );
  DFFSSRX1_HVT sram_rdata_7_reg_6_ ( .D(1'b0), .SETB(n13600), .RSTB(N269), 
        .CLK(clk), .Q(sram_rdata_7[6]) );
  DFFSSRX1_HVT sram_rdata_7_reg_5_ ( .D(1'b0), .SETB(n33), .RSTB(N268), .CLK(
        clk), .Q(sram_rdata_7[5]) );
  DFFSSRX1_HVT sram_rdata_7_reg_4_ ( .D(1'b0), .SETB(n1510), .RSTB(N267), 
        .CLK(clk), .Q(sram_rdata_7[4]) );
  DFFSSRX1_HVT sram_rdata_7_reg_3_ ( .D(1'b0), .SETB(n1800), .RSTB(N266), 
        .CLK(clk), .Q(sram_rdata_7[3]) );
  DFFSSRX1_HVT sram_rdata_7_reg_2_ ( .D(1'b0), .SETB(n13600), .RSTB(N265), 
        .CLK(clk), .Q(sram_rdata_7[2]) );
  DFFSSRX1_HVT sram_rdata_7_reg_1_ ( .D(1'b0), .SETB(n34), .RSTB(N264), .CLK(
        clk), .Q(sram_rdata_7[1]) );
  DFFSSRX1_HVT sram_rdata_7_reg_0_ ( .D(1'b0), .SETB(n1510), .RSTB(N263), 
        .CLK(clk), .Q(sram_rdata_7[0]) );
  AO221X1_HVT U3 ( .A1(1'b1), .A2(n23), .A3(sram_rdata_2[19]), .A4(n6100), 
        .A5(n24), .Y(n_src_aox[259]) );
  AO221X1_HVT U4 ( .A1(1'b1), .A2(n20), .A3(sram_rdata_0[29]), .A4(n13000), 
        .A5(n21), .Y(n_src_aox[253]) );
  AO221X1_HVT U5 ( .A1(1'b1), .A2(n17), .A3(sram_rdata_2[18]), .A4(n10501), 
        .A5(n18), .Y(n_src_aox[258]) );
  AO221X1_HVT U6 ( .A1(1'b1), .A2(n14), .A3(sram_rdata_3[23]), .A4(n12500), 
        .A5(n15), .Y(n_src_aox[151]) );
  AO221X1_HVT U7 ( .A1(1'b1), .A2(n11), .A3(sram_rdata_5[10]), .A4(n1049), 
        .A5(n12), .Y(n_src_aox[122]) );
  AO221X1_HVT U8 ( .A1(1'b1), .A2(n8), .A3(sram_rdata_7[22]), .A4(n1051), .A5(
        n9), .Y(n_src_aox[86]) );
  AO221X1_HVT U9 ( .A1(1'b1), .A2(n5), .A3(sram_rdata_6[12]), .A4(n6200), .A5(
        n6), .Y(n_src_aox[12]) );
  AO221X1_HVT U10 ( .A1(1'b1), .A2(n2), .A3(sram_rdata_6[16]), .A4(n1052), 
        .A5(n3), .Y(n_src_aox[48]) );
  NBUFFX2_HVT U11 ( .A(n1357), .Y(n7600) );
  AO22X1_HVT U13 ( .A1(n1261), .A2(n5000), .A3(n1113), .A4(n1039), .Y(n2) );
  AO22X1_HVT U14 ( .A1(n4400), .A2(sram_rdata_7[16]), .A3(sram_rdata_8[16]), 
        .A4(n4200), .Y(n3) );
  AO22X1_HVT U16 ( .A1(n1189), .A2(n5900), .A3(n1077), .A4(n1041), .Y(n5) );
  AO22X1_HVT U17 ( .A1(n4400), .A2(sram_rdata_7[12]), .A3(sram_rdata_8[12]), 
        .A4(n28), .Y(n6) );
  AO22X1_HVT U19 ( .A1(n1337), .A2(n35), .A3(n1151), .A4(n5300), .Y(n8) );
  AO22X1_HVT U20 ( .A1(n4400), .A2(sram_rdata_8[22]), .A3(sram_rdata_6[22]), 
        .A4(n1354), .Y(n9) );
  AO22X1_HVT U22 ( .A1(n1091), .A2(n35), .A3(n1216), .A4(n5300), .Y(n11) );
  AO22X1_HVT U23 ( .A1(n30), .A2(sram_rdata_3[10]), .A3(sram_rdata_4[10]), 
        .A4(n1354), .Y(n12) );
  AO22X1_HVT U25 ( .A1(n11201), .A2(n5000), .A3(n1274), .A4(n5300), .Y(n14) );
  AO22X1_HVT U26 ( .A1(n4400), .A2(sram_rdata_4[23]), .A3(sram_rdata_5[23]), 
        .A4(n29), .Y(n15) );
  AO22X1_HVT U28 ( .A1(n1296), .A2(n5900), .A3(n1297), .A4(n1039), .Y(n17) );
  AO22X1_HVT U29 ( .A1(n1355), .A2(sram_rdata_0[18]), .A3(sram_rdata_1[18]), 
        .A4(n4100), .Y(n18) );
  AO22X1_HVT U31 ( .A1(n1286), .A2(n5000), .A3(n1287), .A4(n1039), .Y(n20) );
  AO22X1_HVT U32 ( .A1(n1029), .A2(sram_rdata_1[29]), .A3(sram_rdata_2[29]), 
        .A4(n28), .Y(n21) );
  AO22X1_HVT U34 ( .A1(n1298), .A2(n5900), .A3(n1299), .A4(n5300), .Y(n23) );
  AO22X1_HVT U35 ( .A1(n4300), .A2(sram_rdata_0[19]), .A3(sram_rdata_1[19]), 
        .A4(n4200), .Y(n24) );
  NBUFFX2_HVT U36 ( .A(n1162), .Y(n1045) );
  INVX1_HVT U37 ( .A(n1790), .Y(n1740) );
  INVX1_HVT U38 ( .A(srstn), .Y(n777) );
  INVX1_HVT U39 ( .A(n1362), .Y(n3900) );
  AND2X1_HVT U40 ( .A1(mode[1]), .A2(n13601), .Y(n25) );
  INVX2_HVT U41 ( .A(n7500), .Y(n26) );
  INVX2_HVT U42 ( .A(n1700), .Y(n27) );
  INVX2_HVT U43 ( .A(n7500), .Y(n28) );
  INVX2_HVT U44 ( .A(n7500), .Y(n29) );
  INVX1_HVT U45 ( .A(n5800), .Y(n4700) );
  INVX2_HVT U46 ( .A(n7400), .Y(n30) );
  INVX2_HVT U47 ( .A(n7400), .Y(n31) );
  INVX2_HVT U48 ( .A(n7400), .Y(n32) );
  AOI21X1_HVT U49 ( .A1(n13100), .A2(n1361), .A3(n1530), .Y(n1061) );
  INVX2_HVT U50 ( .A(n1740), .Y(n33) );
  INVX2_HVT U51 ( .A(n8000), .Y(n34) );
  AOI21X1_HVT U52 ( .A1(n12500), .A2(n1361), .A3(n1370), .Y(N346) );
  INVX0_HVT U53 ( .A(n1740), .Y(n7900) );
  INVX1_HVT U54 ( .A(n5400), .Y(n8400) );
  INVX1_HVT U55 ( .A(n5400), .Y(n8200) );
  INVX1_HVT U56 ( .A(n5500), .Y(n11800) );
  INVX1_HVT U57 ( .A(n5500), .Y(n11000) );
  AOI21X1_HVT U58 ( .A1(n12700), .A2(n1361), .A3(n1780), .Y(n10601) );
  INVX2_HVT U59 ( .A(n5800), .Y(n35) );
  INVX1_HVT U60 ( .A(n5400), .Y(n10600) );
  INVX1_HVT U61 ( .A(n5400), .Y(n8300) );
  INVX1_HVT U62 ( .A(n5400), .Y(n10700) );
  INVX1_HVT U63 ( .A(n5400), .Y(n10800) );
  INVX1_HVT U64 ( .A(n5400), .Y(n10900) );
  INVX2_HVT U65 ( .A(n5800), .Y(n36) );
  INVX1_HVT U66 ( .A(n5400), .Y(n8100) );
  INVX1_HVT U67 ( .A(n1740), .Y(n1750) );
  INVX1_HVT U68 ( .A(n1770), .Y(n13600) );
  INVX1_HVT U69 ( .A(srstn), .Y(n1510) );
  INVX1_HVT U70 ( .A(n5600), .Y(n9700) );
  INVX1_HVT U71 ( .A(n5700), .Y(n9300) );
  INVX1_HVT U72 ( .A(n1045), .Y(n5400) );
  INVX2_HVT U73 ( .A(n6900), .Y(n37) );
  INVX1_HVT U74 ( .A(n1161), .Y(n5500) );
  INVX1_HVT U75 ( .A(n5700), .Y(n8900) );
  INVX2_HVT U76 ( .A(n6900), .Y(n38) );
  INVX1_HVT U77 ( .A(n1025), .Y(n5600) );
  INVX1_HVT U78 ( .A(n1357), .Y(n5800) );
  INVX1_HVT U79 ( .A(n1024), .Y(n5700) );
  INVX1_HVT U80 ( .A(box_sel[2]), .Y(n1064) );
  INVX1_HVT U81 ( .A(box_sel[3]), .Y(n1063) );
  INVX2_HVT U82 ( .A(n7500), .Y(n4000) );
  INVX0_HVT U83 ( .A(n1700), .Y(n1730) );
  INVX2_HVT U84 ( .A(n7500), .Y(n4100) );
  AND3X2_HVT U85 ( .A1(n1064), .A2(n1063), .A3(n11400), .Y(n1035) );
  INVX2_HVT U86 ( .A(n7500), .Y(n4200) );
  INVX1_HVT U87 ( .A(n25), .Y(n1700) );
  INVX2_HVT U88 ( .A(n7400), .Y(n4300) );
  INVX1_HVT U89 ( .A(n5500), .Y(n11400) );
  INVX2_HVT U90 ( .A(n7400), .Y(n4400) );
  INVX2_HVT U91 ( .A(n7400), .Y(n4500) );
  INVX1_HVT U92 ( .A(n25), .Y(n1059) );
  INVX1_HVT U93 ( .A(n1740), .Y(n7700) );
  INVX1_HVT U94 ( .A(n1740), .Y(n7800) );
  INVX2_HVT U95 ( .A(n5800), .Y(n4600) );
  AND3X2_HVT U96 ( .A1(n1064), .A2(n1063), .A3(n11800), .Y(n1354) );
  INVX1_HVT U97 ( .A(n1700), .Y(n1620) );
  INVX1_HVT U98 ( .A(n1059), .Y(n1580) );
  AND3X2_HVT U99 ( .A1(n1064), .A2(n1063), .A3(n11000), .Y(n1034) );
  INVX2_HVT U100 ( .A(n8000), .Y(n4800) );
  INVX2_HVT U101 ( .A(n1740), .Y(n4900) );
  INVX1_HVT U102 ( .A(n10100), .Y(n10500) );
  INVX1_HVT U103 ( .A(n3900), .Y(n13100) );
  INVX1_HVT U104 ( .A(n10100), .Y(n10300) );
  AND3X2_HVT U105 ( .A1(n1064), .A2(n1063), .A3(n9700), .Y(n1355) );
  INVX1_HVT U106 ( .A(n12400), .Y(n12500) );
  INVX1_HVT U107 ( .A(n5800), .Y(n5900) );
  INVX1_HVT U108 ( .A(n7000), .Y(n7100) );
  INVX1_HVT U109 ( .A(n3900), .Y(n6300) );
  INVX1_HVT U110 ( .A(n10100), .Y(n10400) );
  INVX1_HVT U111 ( .A(n10100), .Y(n10200) );
  AND3X2_HVT U112 ( .A1(n1064), .A2(n1063), .A3(n8900), .Y(n1026) );
  INVX1_HVT U113 ( .A(n3900), .Y(n6200) );
  INVX1_HVT U114 ( .A(n3900), .Y(n12700) );
  AND3X2_HVT U115 ( .A1(n1064), .A2(n1063), .A3(n9300), .Y(n1027) );
  INVX1_HVT U116 ( .A(n10100), .Y(n6400) );
  INVX2_HVT U117 ( .A(n5800), .Y(n5000) );
  INVX2_HVT U118 ( .A(n6900), .Y(n5100) );
  INVX1_HVT U119 ( .A(n1362), .Y(n12400) );
  INVX1_HVT U120 ( .A(n5400), .Y(n5200) );
  INVX2_HVT U121 ( .A(n6900), .Y(n5300) );
  INVX1_HVT U122 ( .A(n1045), .Y(n10100) );
  INVX1_HVT U123 ( .A(n1032), .Y(n7000) );
  DELLN1X2_HVT U124 ( .A(n1161), .Y(n10301) );
  DELLN1X2_HVT U125 ( .A(n1161), .Y(n1031) );
  INVX0_HVT U126 ( .A(mode[0]), .Y(n13601) );
  NBUFFX2_HVT U127 ( .A(n11601), .Y(n1025) );
  DELLN1X2_HVT U128 ( .A(n11601), .Y(n1024) );
  NBUFFX2_HVT U129 ( .A(n1359), .Y(n1041) );
  DELLN1X2_HVT U130 ( .A(n1359), .Y(n1042) );
  DELLN1X2_HVT U131 ( .A(n1359), .Y(n1043) );
  DELLN1X2_HVT U132 ( .A(n1359), .Y(n10401) );
  DELLN1X2_HVT U133 ( .A(n1359), .Y(n1044) );
  DELLN1X2_HVT U134 ( .A(n1359), .Y(n1039) );
  DELLN1X2_HVT U135 ( .A(n1162), .Y(n1046) );
  DELLN1X2_HVT U136 ( .A(n1162), .Y(n1048) );
  DELLN1X2_HVT U137 ( .A(n1162), .Y(n1047) );
  INVX2_HVT U138 ( .A(n1770), .Y(n1370) );
  INVX2_HVT U139 ( .A(n1740), .Y(n1380) );
  INVX2_HVT U140 ( .A(n8000), .Y(n13500) );
  INVX2_HVT U141 ( .A(n1770), .Y(n1530) );
  INVX2_HVT U142 ( .A(n8000), .Y(n1520) );
  INVX2_HVT U143 ( .A(n8000), .Y(n1500) );
  DELLN1X2_HVT U144 ( .A(n1357), .Y(n1057) );
  DELLN1X2_HVT U145 ( .A(n1357), .Y(n1055) );
  DELLN1X2_HVT U146 ( .A(n1357), .Y(n1054) );
  DELLN1X2_HVT U147 ( .A(n1362), .Y(n6000) );
  DELLN1X2_HVT U148 ( .A(n1362), .Y(n6100) );
  DELLN1X2_HVT U149 ( .A(n1362), .Y(n1051) );
  DELLN1X2_HVT U150 ( .A(n1362), .Y(n1053) );
  DELLN1X2_HVT U151 ( .A(n1362), .Y(n1052) );
  INVX2_HVT U152 ( .A(n1059), .Y(n6500) );
  INVX2_HVT U153 ( .A(n1059), .Y(n6600) );
  INVX2_HVT U154 ( .A(n1059), .Y(n1690) );
  INVX2_HVT U155 ( .A(n1059), .Y(n1680) );
  INVX2_HVT U156 ( .A(n1059), .Y(n1670) );
  INVX2_HVT U157 ( .A(n1700), .Y(n6700) );
  INVX2_HVT U158 ( .A(n1700), .Y(n6800) );
  INVX2_HVT U159 ( .A(n1700), .Y(n1720) );
  INVX2_HVT U160 ( .A(n1700), .Y(n1710) );
  DELLN1X2_HVT U161 ( .A(n1362), .Y(n1049) );
  DELLN1X2_HVT U162 ( .A(n1362), .Y(n12200) );
  DELLN1X2_HVT U163 ( .A(n1362), .Y(n12300) );
  DELLN1X2_HVT U164 ( .A(n1362), .Y(n10501) );
  DELLN1X2_HVT U165 ( .A(n1357), .Y(n1058) );
  DELLN1X2_HVT U166 ( .A(n1357), .Y(n1056) );
  INVX0_HVT U167 ( .A(n1041), .Y(n6900) );
  DELLN1X2_HVT U168 ( .A(n1161), .Y(n1032) );
  DELLN1X2_HVT U169 ( .A(n1161), .Y(n1033) );
  INVX0_HVT U170 ( .A(n7000), .Y(n7200) );
  INVX0_HVT U171 ( .A(n7000), .Y(n7300) );
  DELLN1X2_HVT U172 ( .A(n1026), .Y(n1028) );
  INVX0_HVT U173 ( .A(n1355), .Y(n7400) );
  DELLN1X2_HVT U174 ( .A(n1027), .Y(n1029) );
  DELLN1X2_HVT U175 ( .A(n1354), .Y(n1038) );
  DELLN1X2_HVT U176 ( .A(n1035), .Y(n1037) );
  DELLN1X2_HVT U177 ( .A(n1034), .Y(n1036) );
  INVX0_HVT U178 ( .A(n1034), .Y(n7500) );
  INVX2_HVT U179 ( .A(n1740), .Y(n1760) );
  INVX0_HVT U180 ( .A(n1760), .Y(n8000) );
  INVX0_HVT U181 ( .A(n5600), .Y(n8500) );
  INVX0_HVT U182 ( .A(n5600), .Y(n8600) );
  INVX0_HVT U183 ( .A(n5600), .Y(n8700) );
  INVX0_HVT U184 ( .A(n5600), .Y(n8800) );
  INVX0_HVT U185 ( .A(n5700), .Y(n9000) );
  INVX0_HVT U186 ( .A(n5700), .Y(n9100) );
  INVX0_HVT U187 ( .A(n5700), .Y(n9200) );
  INVX0_HVT U188 ( .A(n5700), .Y(n9400) );
  INVX0_HVT U189 ( .A(n5700), .Y(n9500) );
  INVX0_HVT U190 ( .A(n5700), .Y(n9600) );
  INVX0_HVT U191 ( .A(n5600), .Y(n9800) );
  INVX0_HVT U192 ( .A(n5600), .Y(n9900) );
  INVX0_HVT U193 ( .A(n5600), .Y(n10000) );
  INVX0_HVT U194 ( .A(n5500), .Y(n11100) );
  INVX0_HVT U195 ( .A(n5500), .Y(n11200) );
  INVX0_HVT U196 ( .A(n5500), .Y(n11300) );
  INVX0_HVT U197 ( .A(n7000), .Y(n11500) );
  INVX0_HVT U198 ( .A(n7000), .Y(n11600) );
  INVX0_HVT U199 ( .A(n7000), .Y(n11700) );
  INVX0_HVT U200 ( .A(n5500), .Y(n11900) );
  INVX0_HVT U201 ( .A(n5500), .Y(n12000) );
  INVX0_HVT U202 ( .A(n5500), .Y(n12100) );
  INVX0_HVT U203 ( .A(n12400), .Y(n12600) );
  INVX0_HVT U204 ( .A(n3900), .Y(n12800) );
  INVX0_HVT U205 ( .A(n3900), .Y(n12900) );
  INVX0_HVT U206 ( .A(n3900), .Y(n13000) );
  INVX0_HVT U207 ( .A(n3900), .Y(n13200) );
  INVX0_HVT U208 ( .A(n3900), .Y(n13300) );
  INVX0_HVT U209 ( .A(n3900), .Y(n13400) );
  INVX2_HVT U210 ( .A(n1770), .Y(n1800) );
  INVX2_HVT U211 ( .A(n1770), .Y(n1810) );
  INVX2_HVT U212 ( .A(n1770), .Y(n1790) );
  INVX2_HVT U213 ( .A(n1770), .Y(n1780) );
  INVX2_HVT U214 ( .A(N346), .Y(n1390) );
  INVX2_HVT U215 ( .A(N346), .Y(n1400) );
  INVX2_HVT U216 ( .A(N346), .Y(n1410) );
  INVX2_HVT U217 ( .A(N346), .Y(n1420) );
  INVX2_HVT U218 ( .A(n10601), .Y(n1430) );
  INVX2_HVT U219 ( .A(n10601), .Y(n1440) );
  INVX2_HVT U220 ( .A(n10601), .Y(n1450) );
  INVX2_HVT U221 ( .A(n1061), .Y(n1460) );
  INVX2_HVT U222 ( .A(n1061), .Y(n1470) );
  INVX2_HVT U223 ( .A(n1061), .Y(n1480) );
  INVX2_HVT U224 ( .A(n1061), .Y(n1490) );
  INVX2_HVT U225 ( .A(n1620), .Y(n1540) );
  INVX2_HVT U226 ( .A(n1580), .Y(n1550) );
  INVX2_HVT U227 ( .A(n1620), .Y(n1560) );
  INVX2_HVT U228 ( .A(n1580), .Y(n1570) );
  INVX2_HVT U229 ( .A(n1580), .Y(n1590) );
  INVX2_HVT U230 ( .A(n1580), .Y(n1600) );
  INVX2_HVT U231 ( .A(n1580), .Y(n1610) );
  INVX2_HVT U232 ( .A(n1620), .Y(n1630) );
  INVX2_HVT U233 ( .A(n1620), .Y(n1640) );
  INVX2_HVT U234 ( .A(n1620), .Y(n1650) );
  INVX2_HVT U235 ( .A(n1620), .Y(n1660) );
  INVX1_HVT U236 ( .A(n777), .Y(n1770) );
  INVX1_HVT U237 ( .A(box_sel[1]), .Y(n1361) );
  INVX1_HVT U238 ( .A(box_sel[0]), .Y(n1062) );
  AOI22X1_HVT U239 ( .A1(n12600), .A2(sram_rdata_6[0]), .A3(n1058), .A4(n1165), 
        .Y(n1820) );
  AOI22X1_HVT U240 ( .A1(n38), .A2(n1358), .A3(n7600), .A4(n1356), .Y(n1830)
         );
  AOI22X1_HVT U241 ( .A1(n1042), .A2(n1353), .A3(n1056), .A4(n1352), .Y(n1840)
         );
  AOI22X1_HVT U242 ( .A1(n1039), .A2(n1351), .A3(n1055), .A4(n13501), .Y(n1850) );
  AOI22X1_HVT U243 ( .A1(n1042), .A2(n1349), .A3(n35), .A4(n1348), .Y(n1860)
         );
  AOI22X1_HVT U244 ( .A1(n37), .A2(n1347), .A3(n1056), .A4(n1346), .Y(n1870)
         );
  AOI22X1_HVT U245 ( .A1(n1041), .A2(n1345), .A3(n1058), .A4(n1344), .Y(n1880)
         );
  AOI22X1_HVT U246 ( .A1(n10401), .A2(n1343), .A3(n1056), .A4(n1342), .Y(n1890) );
  AOI22X1_HVT U247 ( .A1(n38), .A2(n1341), .A3(n1055), .A4(n13401), .Y(n1900)
         );
  AOI22X1_HVT U248 ( .A1(n1041), .A2(n1339), .A3(n1057), .A4(n1338), .Y(n1910)
         );
  AOI22X1_HVT U249 ( .A1(n1043), .A2(n1337), .A3(n35), .A4(n1336), .Y(n1920)
         );
  AOI22X1_HVT U250 ( .A1(n1039), .A2(n1335), .A3(n5900), .A4(n1334), .Y(n1930)
         );
  AOI22X1_HVT U251 ( .A1(n1042), .A2(n1333), .A3(n1058), .A4(n1332), .Y(n1940)
         );
  AOI22X1_HVT U252 ( .A1(n37), .A2(n1331), .A3(n36), .A4(n13301), .Y(n1950) );
  AOI22X1_HVT U253 ( .A1(n5100), .A2(n1329), .A3(n5000), .A4(n1328), .Y(n1960)
         );
  AOI22X1_HVT U254 ( .A1(n5300), .A2(n1327), .A3(n7600), .A4(n1326), .Y(n1970)
         );
  AOI22X1_HVT U255 ( .A1(n1044), .A2(n1325), .A3(n35), .A4(n1324), .Y(n1980)
         );
  AOI22X1_HVT U256 ( .A1(n1039), .A2(n1323), .A3(n7600), .A4(n1322), .Y(n1990)
         );
  AOI22X1_HVT U257 ( .A1(n1042), .A2(n1321), .A3(n36), .A4(n13201), .Y(n2000)
         );
  AOI22X1_HVT U258 ( .A1(n37), .A2(n1319), .A3(n5000), .A4(n1318), .Y(n2010)
         );
  AOI22X1_HVT U259 ( .A1(n10401), .A2(n1317), .A3(n36), .A4(n1316), .Y(n2020)
         );
  AOI22X1_HVT U260 ( .A1(n1039), .A2(n1315), .A3(n7600), .A4(n1314), .Y(n2030)
         );
  AOI22X1_HVT U261 ( .A1(n5300), .A2(n1313), .A3(n4600), .A4(n1312), .Y(n2040)
         );
  AOI22X1_HVT U262 ( .A1(n37), .A2(n1311), .A3(n5000), .A4(n13101), .Y(n2050)
         );
  AOI22X1_HVT U263 ( .A1(n1039), .A2(n1309), .A3(n1056), .A4(n1308), .Y(n2060)
         );
  AOI22X1_HVT U264 ( .A1(n37), .A2(n1307), .A3(n5000), .A4(n1306), .Y(n2070)
         );
  AOI22X1_HVT U265 ( .A1(n37), .A2(n1305), .A3(n1056), .A4(n1304), .Y(n2080)
         );
  AOI22X1_HVT U266 ( .A1(n1043), .A2(n1303), .A3(n7600), .A4(n1302), .Y(n2090)
         );
  AOI22X1_HVT U267 ( .A1(n1042), .A2(n1301), .A3(n4600), .A4(n13001), .Y(n2100) );
  AOI22X1_HVT U268 ( .A1(n37), .A2(n1295), .A3(n1058), .A4(n1294), .Y(n2110)
         );
  AOI22X1_HVT U269 ( .A1(n5100), .A2(n1293), .A3(n7600), .A4(n1292), .Y(n2120)
         );
  AOI22X1_HVT U270 ( .A1(n5300), .A2(n1291), .A3(n36), .A4(n12901), .Y(n2130)
         );
  AOI22X1_HVT U271 ( .A1(n10401), .A2(n1289), .A3(n35), .A4(n1288), .Y(n2140)
         );
  AOI22X1_HVT U272 ( .A1(n5300), .A2(n1285), .A3(n36), .A4(n1284), .Y(n2150)
         );
  AOI22X1_HVT U273 ( .A1(n38), .A2(n1283), .A3(n4700), .A4(n1282), .Y(n2160)
         );
  AOI22X1_HVT U274 ( .A1(n10401), .A2(n1281), .A3(n1054), .A4(n12801), .Y(
        n2170) );
  AOI22X1_HVT U275 ( .A1(n10401), .A2(n1279), .A3(n5000), .A4(n1278), .Y(n2180) );
  AOI22X1_HVT U276 ( .A1(n5100), .A2(n1277), .A3(n4600), .A4(n1276), .Y(n2190)
         );
  AOI22X1_HVT U277 ( .A1(n1039), .A2(n1275), .A3(n1058), .A4(n1274), .Y(n2200)
         );
  AOI22X1_HVT U278 ( .A1(n1044), .A2(n1273), .A3(n36), .A4(n1272), .Y(n2210)
         );
  AOI22X1_HVT U279 ( .A1(n10401), .A2(n1271), .A3(n1058), .A4(n12701), .Y(
        n2220) );
  AOI22X1_HVT U280 ( .A1(n38), .A2(n1269), .A3(n4700), .A4(n1268), .Y(n2230)
         );
  AOI22X1_HVT U281 ( .A1(n1044), .A2(n1267), .A3(n4700), .A4(n1266), .Y(n2240)
         );
  AOI22X1_HVT U282 ( .A1(n1044), .A2(n1265), .A3(n35), .A4(n1264), .Y(n2250)
         );
  AOI22X1_HVT U283 ( .A1(n1042), .A2(n1263), .A3(n5900), .A4(n1262), .Y(n2260)
         );
  AOI22X1_HVT U284 ( .A1(n1044), .A2(n1261), .A3(n1055), .A4(n12601), .Y(n2270) );
  AOI22X1_HVT U285 ( .A1(n1043), .A2(n1259), .A3(n1057), .A4(n1258), .Y(n2280)
         );
  AOI22X1_HVT U286 ( .A1(n1042), .A2(n1257), .A3(n1057), .A4(n1256), .Y(n2290)
         );
  AOI22X1_HVT U287 ( .A1(n5300), .A2(n1255), .A3(n1056), .A4(n1254), .Y(n2300)
         );
  AOI22X1_HVT U288 ( .A1(n1044), .A2(n1253), .A3(n35), .A4(n1252), .Y(n2310)
         );
  AOI22X1_HVT U289 ( .A1(n1041), .A2(n1251), .A3(n36), .A4(n12501), .Y(n2320)
         );
  AOI22X1_HVT U290 ( .A1(n10401), .A2(n1249), .A3(n1057), .A4(n1248), .Y(n2330) );
  AOI22X1_HVT U291 ( .A1(n10401), .A2(n1247), .A3(n1058), .A4(n1246), .Y(n2340) );
  AOI22X1_HVT U292 ( .A1(n1043), .A2(n1245), .A3(n1054), .A4(n1244), .Y(n2350)
         );
  AOI22X1_HVT U293 ( .A1(n1043), .A2(n1243), .A3(n1056), .A4(n1242), .Y(n2360)
         );
  AOI22X1_HVT U294 ( .A1(n38), .A2(n1241), .A3(n35), .A4(n12401), .Y(n2370) );
  AOI22X1_HVT U295 ( .A1(n1043), .A2(n1239), .A3(n5000), .A4(n1238), .Y(n2380)
         );
  AOI22X1_HVT U296 ( .A1(n1042), .A2(n1237), .A3(n1058), .A4(n1236), .Y(n2390)
         );
  AOI22X1_HVT U297 ( .A1(n5100), .A2(n1235), .A3(n5900), .A4(n1234), .Y(n2400)
         );
  AOI22X1_HVT U298 ( .A1(n1043), .A2(n1233), .A3(n5000), .A4(n1232), .Y(n2410)
         );
  AOI22X1_HVT U299 ( .A1(n1044), .A2(n1231), .A3(n4700), .A4(n12301), .Y(n2420) );
  AOI22X1_HVT U300 ( .A1(n1044), .A2(n1229), .A3(n4600), .A4(n1228), .Y(n2430)
         );
  AOI22X1_HVT U301 ( .A1(n38), .A2(n1227), .A3(n4700), .A4(n1226), .Y(n2440)
         );
  AOI22X1_HVT U302 ( .A1(n1042), .A2(n1225), .A3(n1057), .A4(n1224), .Y(n2450)
         );
  AOI22X1_HVT U303 ( .A1(n1042), .A2(n1223), .A3(n1055), .A4(n1222), .Y(n2460)
         );
  AOI22X1_HVT U304 ( .A1(n10401), .A2(n1221), .A3(n5000), .A4(n12201), .Y(
        n2470) );
  AOI22X1_HVT U305 ( .A1(n10401), .A2(n1219), .A3(n5900), .A4(n1218), .Y(n2480) );
  AOI22X1_HVT U306 ( .A1(n1043), .A2(n1217), .A3(n4600), .A4(n1216), .Y(n2490)
         );
  AOI22X1_HVT U307 ( .A1(n1044), .A2(n1215), .A3(n4700), .A4(n1214), .Y(n2500)
         );
  AOI22X1_HVT U308 ( .A1(n38), .A2(n1213), .A3(n4700), .A4(n1212), .Y(n2510)
         );
  AOI22X1_HVT U309 ( .A1(n38), .A2(n1211), .A3(n1058), .A4(n12101), .Y(n2520)
         );
  AOI22X1_HVT U310 ( .A1(n1041), .A2(n1209), .A3(n36), .A4(n1208), .Y(n2530)
         );
  AOI22X1_HVT U311 ( .A1(n1043), .A2(n1207), .A3(n1057), .A4(n1206), .Y(n2540)
         );
  AOI22X1_HVT U312 ( .A1(n1044), .A2(n1205), .A3(n35), .A4(n1204), .Y(n2550)
         );
  AOI22X1_HVT U313 ( .A1(n37), .A2(n1203), .A3(n5900), .A4(n1202), .Y(n2560)
         );
  AOI22X1_HVT U314 ( .A1(n5100), .A2(n1201), .A3(n7600), .A4(n12001), .Y(n2570) );
  AOI22X1_HVT U315 ( .A1(n1043), .A2(n1199), .A3(n5000), .A4(n1198), .Y(n2580)
         );
  AOI22X1_HVT U316 ( .A1(n5300), .A2(n1197), .A3(n1054), .A4(n1196), .Y(n2590)
         );
  AOI22X1_HVT U317 ( .A1(n1044), .A2(n1195), .A3(n7600), .A4(n1194), .Y(n2600)
         );
  AOI22X1_HVT U318 ( .A1(n10401), .A2(n1193), .A3(n35), .A4(n1192), .Y(n2610)
         );
  AOI22X1_HVT U319 ( .A1(n5100), .A2(n1191), .A3(n1055), .A4(n11901), .Y(n2620) );
  AOI22X1_HVT U320 ( .A1(n1042), .A2(n1189), .A3(n4700), .A4(n1188), .Y(n2630)
         );
  AOI22X1_HVT U321 ( .A1(n1042), .A2(n1187), .A3(n1056), .A4(n1186), .Y(n2640)
         );
  AOI22X1_HVT U322 ( .A1(n37), .A2(n1185), .A3(n1055), .A4(n1184), .Y(n2650)
         );
  AOI22X1_HVT U323 ( .A1(n38), .A2(n1183), .A3(n5900), .A4(n1182), .Y(n2660)
         );
  AOI22X1_HVT U324 ( .A1(n38), .A2(n1181), .A3(n4600), .A4(n11801), .Y(n2670)
         );
  AOI22X1_HVT U325 ( .A1(n37), .A2(n1179), .A3(n36), .A4(n1178), .Y(n2680) );
  AOI22X1_HVT U326 ( .A1(n1044), .A2(n1177), .A3(n7600), .A4(n1176), .Y(n2690)
         );
  AOI22X1_HVT U327 ( .A1(n1043), .A2(n1175), .A3(n36), .A4(n1174), .Y(n2700)
         );
  AOI22X1_HVT U328 ( .A1(n1039), .A2(n1173), .A3(n1058), .A4(n1172), .Y(n2710)
         );
  AOI22X1_HVT U329 ( .A1(n1043), .A2(n1171), .A3(n7600), .A4(n11701), .Y(n2720) );
  AOI22X1_HVT U330 ( .A1(n38), .A2(n1169), .A3(n4600), .A4(n1168), .Y(n2730)
         );
  AOI22X1_HVT U331 ( .A1(n1044), .A2(n1167), .A3(n1057), .A4(n1166), .Y(n2740)
         );
  AOI22X1_HVT U332 ( .A1(n1043), .A2(n1165), .A3(n1054), .A4(n1164), .Y(n2750)
         );
  AOI22X1_HVT U333 ( .A1(n38), .A2(n1356), .A3(n36), .A4(n1163), .Y(n2760) );
  AOI22X1_HVT U334 ( .A1(n37), .A2(n1352), .A3(n1055), .A4(n1159), .Y(n2770)
         );
  AOI22X1_HVT U335 ( .A1(n1044), .A2(n13501), .A3(n1057), .A4(n1158), .Y(n2780) );
  AOI22X1_HVT U336 ( .A1(n1043), .A2(n1348), .A3(n4600), .A4(n1157), .Y(n2790)
         );
  AOI22X1_HVT U337 ( .A1(n38), .A2(n1346), .A3(n5000), .A4(n1156), .Y(n2800)
         );
  AOI22X1_HVT U338 ( .A1(n5100), .A2(n1344), .A3(n4700), .A4(n1155), .Y(n2810)
         );
  AOI22X1_HVT U339 ( .A1(n1043), .A2(n1342), .A3(n36), .A4(n1154), .Y(n2820)
         );
  AOI22X1_HVT U340 ( .A1(n1043), .A2(n13401), .A3(n5900), .A4(n1153), .Y(n2830) );
  AOI22X1_HVT U341 ( .A1(n5100), .A2(n1338), .A3(n4700), .A4(n1152), .Y(n2840)
         );
  AOI22X1_HVT U342 ( .A1(n5100), .A2(n1336), .A3(n4600), .A4(n1151), .Y(n2850)
         );
  AOI22X1_HVT U343 ( .A1(n1359), .A2(n1334), .A3(n1054), .A4(n11501), .Y(n2860) );
  AOI22X1_HVT U344 ( .A1(n5300), .A2(n1332), .A3(n1058), .A4(n1149), .Y(n2870)
         );
  AOI22X1_HVT U345 ( .A1(n38), .A2(n13301), .A3(n1057), .A4(n1148), .Y(n2880)
         );
  AOI22X1_HVT U346 ( .A1(n1039), .A2(n1328), .A3(n1056), .A4(n1147), .Y(n2890)
         );
  AOI22X1_HVT U347 ( .A1(n1359), .A2(n1326), .A3(n1058), .A4(n1146), .Y(n2900)
         );
  AOI22X1_HVT U348 ( .A1(n1044), .A2(n1324), .A3(n4600), .A4(n1145), .Y(n2910)
         );
  AOI22X1_HVT U349 ( .A1(n5100), .A2(n1322), .A3(n1058), .A4(n1144), .Y(n2920)
         );
  AOI22X1_HVT U350 ( .A1(n1044), .A2(n13201), .A3(n4700), .A4(n1143), .Y(n2930) );
  AOI22X1_HVT U351 ( .A1(n1043), .A2(n1318), .A3(n1057), .A4(n1142), .Y(n2940)
         );
  AOI22X1_HVT U352 ( .A1(n38), .A2(n1316), .A3(n5000), .A4(n1141), .Y(n2950)
         );
  AOI22X1_HVT U353 ( .A1(n1044), .A2(n1314), .A3(n1054), .A4(n11401), .Y(n2960) );
  AOI22X1_HVT U354 ( .A1(n10401), .A2(n1312), .A3(n35), .A4(n1139), .Y(n2970)
         );
  AOI22X1_HVT U355 ( .A1(n5100), .A2(n13101), .A3(n1055), .A4(n1138), .Y(n2980) );
  AOI22X1_HVT U356 ( .A1(n38), .A2(n1308), .A3(n1055), .A4(n1137), .Y(n2990)
         );
  AOI22X1_HVT U357 ( .A1(n37), .A2(n1306), .A3(n1054), .A4(n1136), .Y(n3000)
         );
  AOI22X1_HVT U358 ( .A1(n1041), .A2(n1304), .A3(n1057), .A4(n1135), .Y(n3010)
         );
  AOI22X1_HVT U359 ( .A1(n38), .A2(n1302), .A3(n1054), .A4(n1134), .Y(n3020)
         );
  AOI22X1_HVT U360 ( .A1(n5100), .A2(n13001), .A3(n4600), .A4(n1133), .Y(n3030) );
  AOI22X1_HVT U361 ( .A1(n5100), .A2(n1298), .A3(n1057), .A4(n1132), .Y(n3040)
         );
  AOI22X1_HVT U362 ( .A1(n1044), .A2(n1296), .A3(n1058), .A4(n1131), .Y(n3050)
         );
  AOI22X1_HVT U363 ( .A1(n10401), .A2(n1294), .A3(n7600), .A4(n11301), .Y(
        n3060) );
  AOI22X1_HVT U364 ( .A1(n1043), .A2(n1292), .A3(n1056), .A4(n1129), .Y(n3070)
         );
  AOI22X1_HVT U365 ( .A1(n1041), .A2(n12901), .A3(n1058), .A4(n1128), .Y(n3080) );
  AOI22X1_HVT U366 ( .A1(n38), .A2(n1288), .A3(n4600), .A4(n1127), .Y(n3090)
         );
  AOI22X1_HVT U367 ( .A1(n1043), .A2(n1286), .A3(n36), .A4(n1126), .Y(n3100)
         );
  AOI22X1_HVT U368 ( .A1(n1043), .A2(n1284), .A3(n1057), .A4(n1125), .Y(n3110)
         );
  AOI22X1_HVT U369 ( .A1(n10401), .A2(n1282), .A3(n1055), .A4(n1124), .Y(n3120) );
  AOI22X1_HVT U370 ( .A1(n1043), .A2(n12801), .A3(n1054), .A4(n1123), .Y(n3130) );
  AOI22X1_HVT U371 ( .A1(n10401), .A2(n1278), .A3(n1055), .A4(n1122), .Y(n3140) );
  AOI22X1_HVT U372 ( .A1(n1359), .A2(n1276), .A3(n4600), .A4(n1121), .Y(n3150)
         );
  AOI22X1_HVT U373 ( .A1(n1039), .A2(n1272), .A3(n1056), .A4(n1119), .Y(n3160)
         );
  AOI22X1_HVT U374 ( .A1(n37), .A2(n12701), .A3(n7600), .A4(n1118), .Y(n3170)
         );
  AOI22X1_HVT U375 ( .A1(n1042), .A2(n1268), .A3(n4700), .A4(n1117), .Y(n3180)
         );
  AOI22X1_HVT U376 ( .A1(n1041), .A2(n1266), .A3(n1058), .A4(n1116), .Y(n3190)
         );
  AOI22X1_HVT U377 ( .A1(n1043), .A2(n1264), .A3(n4600), .A4(n1115), .Y(n3200)
         );
  AOI22X1_HVT U378 ( .A1(n1043), .A2(n1262), .A3(n5000), .A4(n1114), .Y(n3210)
         );
  AOI22X1_HVT U379 ( .A1(n38), .A2(n12601), .A3(n1056), .A4(n1113), .Y(n3220)
         );
  AOI22X1_HVT U380 ( .A1(n5300), .A2(n1258), .A3(n1054), .A4(n1112), .Y(n3230)
         );
  AOI22X1_HVT U381 ( .A1(n1039), .A2(n1256), .A3(n7600), .A4(n1111), .Y(n3240)
         );
  AOI22X1_HVT U382 ( .A1(n1039), .A2(n1254), .A3(n1057), .A4(n11101), .Y(n3250) );
  AOI22X1_HVT U383 ( .A1(n10401), .A2(n1252), .A3(n35), .A4(n1109), .Y(n3260)
         );
  AOI22X1_HVT U384 ( .A1(n1043), .A2(n12501), .A3(n4700), .A4(n1108), .Y(n327)
         );
  AOI22X1_HVT U385 ( .A1(n1041), .A2(n1248), .A3(n1058), .A4(n1107), .Y(n328)
         );
  AOI22X1_HVT U386 ( .A1(n1044), .A2(n1246), .A3(n1056), .A4(n1106), .Y(n329)
         );
  AOI22X1_HVT U387 ( .A1(n38), .A2(n1244), .A3(n7600), .A4(n1105), .Y(n330) );
  AOI22X1_HVT U388 ( .A1(n1043), .A2(n1242), .A3(n7600), .A4(n1104), .Y(n331)
         );
  AOI22X1_HVT U389 ( .A1(n10401), .A2(n12401), .A3(n35), .A4(n1103), .Y(n332)
         );
  AOI22X1_HVT U390 ( .A1(n10401), .A2(n1238), .A3(n5900), .A4(n1102), .Y(n333)
         );
  AOI22X1_HVT U391 ( .A1(n1041), .A2(n1236), .A3(n7600), .A4(n1101), .Y(n334)
         );
  AOI22X1_HVT U392 ( .A1(n1041), .A2(n1234), .A3(n1056), .A4(n11001), .Y(n335)
         );
  AOI22X1_HVT U393 ( .A1(n1041), .A2(n1232), .A3(n7600), .A4(n1099), .Y(n336)
         );
  AOI22X1_HVT U394 ( .A1(n5300), .A2(n12301), .A3(n1054), .A4(n1098), .Y(n337)
         );
  AOI22X1_HVT U395 ( .A1(n38), .A2(n1228), .A3(n35), .A4(n1097), .Y(n338) );
  AOI22X1_HVT U396 ( .A1(n5300), .A2(n1226), .A3(n36), .A4(n1096), .Y(n339) );
  AOI22X1_HVT U397 ( .A1(n10401), .A2(n1224), .A3(n1056), .A4(n1095), .Y(n340)
         );
  AOI22X1_HVT U398 ( .A1(n1041), .A2(n1222), .A3(n36), .A4(n1094), .Y(n341) );
  AOI22X1_HVT U399 ( .A1(n1044), .A2(n12201), .A3(n1056), .A4(n1093), .Y(n342)
         );
  AOI22X1_HVT U400 ( .A1(n5100), .A2(n1218), .A3(n5900), .A4(n1092), .Y(n343)
         );
  AOI22X1_HVT U401 ( .A1(n10401), .A2(n1214), .A3(n1055), .A4(n10901), .Y(n344) );
  AOI22X1_HVT U402 ( .A1(n10401), .A2(n1212), .A3(n36), .A4(n1089), .Y(n345)
         );
  AOI22X1_HVT U403 ( .A1(n1039), .A2(n12101), .A3(n1057), .A4(n1088), .Y(n3460) );
  AOI22X1_HVT U404 ( .A1(n1041), .A2(n1208), .A3(n1055), .A4(n1087), .Y(n347)
         );
  AOI22X1_HVT U405 ( .A1(n1041), .A2(n1206), .A3(n1055), .A4(n1086), .Y(n348)
         );
  AOI22X1_HVT U406 ( .A1(n1359), .A2(n1204), .A3(n4600), .A4(n1085), .Y(n349)
         );
  AOI22X1_HVT U407 ( .A1(n5300), .A2(n1202), .A3(n1054), .A4(n1084), .Y(n350)
         );
  AOI22X1_HVT U408 ( .A1(n37), .A2(n12001), .A3(n1056), .A4(n1083), .Y(n351)
         );
  AOI22X1_HVT U409 ( .A1(n1044), .A2(n1198), .A3(n7600), .A4(n1082), .Y(n352)
         );
  AOI22X1_HVT U410 ( .A1(n37), .A2(n1196), .A3(n1055), .A4(n1081), .Y(n353) );
  AOI22X1_HVT U411 ( .A1(n37), .A2(n1194), .A3(n7600), .A4(n10801), .Y(n354)
         );
  AOI22X1_HVT U412 ( .A1(n1042), .A2(n1192), .A3(n35), .A4(n1079), .Y(n355) );
  AOI22X1_HVT U413 ( .A1(n1039), .A2(n11901), .A3(n1055), .A4(n1078), .Y(n356)
         );
  AOI22X1_HVT U414 ( .A1(n5300), .A2(n1188), .A3(n36), .A4(n1077), .Y(n357) );
  AOI22X1_HVT U415 ( .A1(n5300), .A2(n1186), .A3(n1054), .A4(n1076), .Y(n358)
         );
  AOI22X1_HVT U416 ( .A1(n1044), .A2(n1184), .A3(n1057), .A4(n1075), .Y(n359)
         );
  AOI22X1_HVT U417 ( .A1(n1042), .A2(n1182), .A3(n1057), .A4(n1074), .Y(n360)
         );
  AOI22X1_HVT U418 ( .A1(n37), .A2(n11801), .A3(n4600), .A4(n1073), .Y(n361)
         );
  AOI22X1_HVT U419 ( .A1(n1042), .A2(n1178), .A3(n1057), .A4(n1072), .Y(n362)
         );
  AOI22X1_HVT U420 ( .A1(n5300), .A2(n1176), .A3(n7600), .A4(n1071), .Y(n363)
         );
  AOI22X1_HVT U421 ( .A1(n10401), .A2(n1174), .A3(n1058), .A4(n10701), .Y(n364) );
  AOI22X1_HVT U422 ( .A1(n5300), .A2(n1172), .A3(n4700), .A4(n1069), .Y(n365)
         );
  AOI22X1_HVT U423 ( .A1(n1359), .A2(n11701), .A3(n36), .A4(n1068), .Y(n366)
         );
  AOI22X1_HVT U424 ( .A1(n37), .A2(n1168), .A3(n4600), .A4(n1067), .Y(n367) );
  AOI22X1_HVT U425 ( .A1(n1039), .A2(n1166), .A3(n1057), .A4(n1066), .Y(n368)
         );
  AOI22X1_HVT U426 ( .A1(n37), .A2(n1164), .A3(n5000), .A4(n1065), .Y(n369) );
  AOI22X1_HVT U427 ( .A1(n10401), .A2(n1163), .A3(n1054), .A4(n1358), .Y(n370)
         );
  AOI22X1_HVT U428 ( .A1(n1042), .A2(n1159), .A3(n1054), .A4(n1353), .Y(n371)
         );
  AOI22X1_HVT U429 ( .A1(n38), .A2(n1158), .A3(n1054), .A4(n1351), .Y(n372) );
  AOI22X1_HVT U430 ( .A1(n1042), .A2(n1157), .A3(n35), .A4(n1349), .Y(n373) );
  AOI22X1_HVT U431 ( .A1(n5100), .A2(n1156), .A3(n1054), .A4(n1347), .Y(n374)
         );
  AOI22X1_HVT U432 ( .A1(n1044), .A2(n1155), .A3(n1056), .A4(n1345), .Y(n375)
         );
  AOI22X1_HVT U433 ( .A1(n1041), .A2(n1154), .A3(n5000), .A4(n1343), .Y(n376)
         );
  AOI22X1_HVT U434 ( .A1(n1041), .A2(n1153), .A3(n1058), .A4(n1341), .Y(n377)
         );
  AOI22X1_HVT U435 ( .A1(n37), .A2(n1152), .A3(n1054), .A4(n1339), .Y(n378) );
  AOI22X1_HVT U436 ( .A1(n1041), .A2(n11501), .A3(n36), .A4(n1335), .Y(n379)
         );
  AOI22X1_HVT U437 ( .A1(n10401), .A2(n1149), .A3(n36), .A4(n1333), .Y(n380)
         );
  AOI22X1_HVT U438 ( .A1(n1044), .A2(n1148), .A3(n1055), .A4(n1331), .Y(n381)
         );
  AOI22X1_HVT U439 ( .A1(n1042), .A2(n1147), .A3(n1055), .A4(n1329), .Y(n382)
         );
  AOI22X1_HVT U440 ( .A1(n1042), .A2(n1146), .A3(n1055), .A4(n1327), .Y(n383)
         );
  AOI22X1_HVT U441 ( .A1(n5100), .A2(n1145), .A3(n35), .A4(n1325), .Y(n384) );
  AOI22X1_HVT U442 ( .A1(n5300), .A2(n1144), .A3(n1057), .A4(n1323), .Y(n385)
         );
  AOI22X1_HVT U443 ( .A1(n5100), .A2(n1143), .A3(n1057), .A4(n1321), .Y(n386)
         );
  AOI22X1_HVT U444 ( .A1(n10401), .A2(n1142), .A3(n4700), .A4(n1319), .Y(n387)
         );
  AOI22X1_HVT U445 ( .A1(n1044), .A2(n1141), .A3(n36), .A4(n1317), .Y(n388) );
  AOI22X1_HVT U446 ( .A1(n1041), .A2(n11401), .A3(n1056), .A4(n1315), .Y(n389)
         );
  AOI22X1_HVT U447 ( .A1(n37), .A2(n1139), .A3(n35), .A4(n1313), .Y(n3901) );
  AOI22X1_HVT U448 ( .A1(n1043), .A2(n1138), .A3(n5000), .A4(n1311), .Y(n391)
         );
  AOI22X1_HVT U449 ( .A1(n5300), .A2(n1137), .A3(n7600), .A4(n1309), .Y(n392)
         );
  AOI22X1_HVT U450 ( .A1(n5300), .A2(n1136), .A3(n1054), .A4(n1307), .Y(n393)
         );
  AOI22X1_HVT U451 ( .A1(n1042), .A2(n1135), .A3(n5900), .A4(n1305), .Y(n394)
         );
  AOI22X1_HVT U452 ( .A1(n1039), .A2(n1134), .A3(n1057), .A4(n1303), .Y(n395)
         );
  AOI22X1_HVT U453 ( .A1(n1042), .A2(n1133), .A3(n35), .A4(n1301), .Y(n396) );
  AOI22X1_HVT U454 ( .A1(n5100), .A2(n1132), .A3(n1055), .A4(n1299), .Y(n397)
         );
  AOI22X1_HVT U455 ( .A1(n37), .A2(n1131), .A3(n4600), .A4(n1297), .Y(n398) );
  AOI22X1_HVT U456 ( .A1(n5100), .A2(n11301), .A3(n36), .A4(n1295), .Y(n399)
         );
  AOI22X1_HVT U457 ( .A1(n5300), .A2(n1129), .A3(n1058), .A4(n1293), .Y(n4001)
         );
  AOI22X1_HVT U458 ( .A1(n1041), .A2(n1128), .A3(n36), .A4(n1291), .Y(n401) );
  AOI22X1_HVT U459 ( .A1(n1042), .A2(n1127), .A3(n4600), .A4(n1289), .Y(n402)
         );
  AOI22X1_HVT U460 ( .A1(n5100), .A2(n1126), .A3(n1055), .A4(n1287), .Y(n403)
         );
  AOI22X1_HVT U461 ( .A1(n1041), .A2(n1125), .A3(n35), .A4(n1285), .Y(n404) );
  AOI22X1_HVT U462 ( .A1(n5100), .A2(n1124), .A3(n5900), .A4(n1283), .Y(n405)
         );
  AOI22X1_HVT U463 ( .A1(n5100), .A2(n1123), .A3(n4700), .A4(n1281), .Y(n406)
         );
  AOI22X1_HVT U464 ( .A1(n38), .A2(n1122), .A3(n1054), .A4(n1279), .Y(n407) );
  AOI22X1_HVT U465 ( .A1(n5100), .A2(n1121), .A3(n4600), .A4(n1277), .Y(n408)
         );
  AOI22X1_HVT U466 ( .A1(n37), .A2(n11201), .A3(n5900), .A4(n1275), .Y(n409)
         );
  AOI22X1_HVT U467 ( .A1(n1039), .A2(n1119), .A3(n1056), .A4(n1273), .Y(n4101)
         );
  AOI22X1_HVT U468 ( .A1(n1041), .A2(n1118), .A3(n5000), .A4(n1271), .Y(n411)
         );
  AOI22X1_HVT U469 ( .A1(n1043), .A2(n1117), .A3(n1058), .A4(n1269), .Y(n412)
         );
  AOI22X1_HVT U470 ( .A1(n1041), .A2(n1116), .A3(n1058), .A4(n1267), .Y(n413)
         );
  AOI22X1_HVT U471 ( .A1(n38), .A2(n1115), .A3(n35), .A4(n1265), .Y(n414) );
  AOI22X1_HVT U472 ( .A1(n1039), .A2(n1114), .A3(n1056), .A4(n1263), .Y(n415)
         );
  AOI22X1_HVT U473 ( .A1(n1039), .A2(n1112), .A3(n1057), .A4(n1259), .Y(n416)
         );
  AOI22X1_HVT U474 ( .A1(n1044), .A2(n1111), .A3(n1056), .A4(n1257), .Y(n417)
         );
  AOI22X1_HVT U475 ( .A1(n37), .A2(n11101), .A3(n1055), .A4(n1255), .Y(n418)
         );
  AOI22X1_HVT U476 ( .A1(n1042), .A2(n1109), .A3(n4600), .A4(n1253), .Y(n419)
         );
  AOI22X1_HVT U477 ( .A1(n5300), .A2(n1108), .A3(n1057), .A4(n1251), .Y(n4201)
         );
  AOI22X1_HVT U478 ( .A1(n10401), .A2(n1107), .A3(n1054), .A4(n1249), .Y(n421)
         );
  AOI22X1_HVT U479 ( .A1(n5100), .A2(n1106), .A3(n36), .A4(n1247), .Y(n422) );
  AOI22X1_HVT U480 ( .A1(n5100), .A2(n1105), .A3(n1055), .A4(n1245), .Y(n423)
         );
  AOI22X1_HVT U481 ( .A1(n1041), .A2(n1104), .A3(n5000), .A4(n1243), .Y(n424)
         );
  AOI22X1_HVT U482 ( .A1(n10401), .A2(n1103), .A3(n4600), .A4(n1241), .Y(n425)
         );
  AOI22X1_HVT U483 ( .A1(n37), .A2(n1102), .A3(n1054), .A4(n1239), .Y(n426) );
  AOI22X1_HVT U484 ( .A1(n38), .A2(n1101), .A3(n1057), .A4(n1237), .Y(n427) );
  AOI22X1_HVT U485 ( .A1(n5300), .A2(n11001), .A3(n1058), .A4(n1235), .Y(n428)
         );
  AOI22X1_HVT U486 ( .A1(n1042), .A2(n1099), .A3(n1056), .A4(n1233), .Y(n429)
         );
  AOI22X1_HVT U487 ( .A1(n1039), .A2(n1098), .A3(n1057), .A4(n1231), .Y(n4301)
         );
  AOI22X1_HVT U488 ( .A1(n5100), .A2(n1097), .A3(n35), .A4(n1229), .Y(n431) );
  AOI22X1_HVT U489 ( .A1(n10401), .A2(n1096), .A3(n1054), .A4(n1227), .Y(n432)
         );
  AOI22X1_HVT U490 ( .A1(n1359), .A2(n1095), .A3(n1055), .A4(n1225), .Y(n433)
         );
  AOI22X1_HVT U491 ( .A1(n1042), .A2(n1094), .A3(n36), .A4(n1223), .Y(n434) );
  AOI22X1_HVT U492 ( .A1(n38), .A2(n1093), .A3(n1056), .A4(n1221), .Y(n435) );
  AOI22X1_HVT U493 ( .A1(n37), .A2(n1092), .A3(n36), .A4(n1219), .Y(n436) );
  AOI22X1_HVT U494 ( .A1(n5100), .A2(n1091), .A3(n35), .A4(n1217), .Y(n437) );
  AOI22X1_HVT U495 ( .A1(n1039), .A2(n10901), .A3(n4700), .A4(n1215), .Y(n438)
         );
  AOI22X1_HVT U496 ( .A1(n1041), .A2(n1089), .A3(n1058), .A4(n1213), .Y(n439)
         );
  AOI22X1_HVT U497 ( .A1(n1359), .A2(n1088), .A3(n1054), .A4(n1211), .Y(n4401)
         );
  AOI22X1_HVT U498 ( .A1(n1043), .A2(n1087), .A3(n7600), .A4(n1209), .Y(n441)
         );
  AOI22X1_HVT U499 ( .A1(n5300), .A2(n1086), .A3(n1054), .A4(n1207), .Y(n442)
         );
  AOI22X1_HVT U500 ( .A1(n1044), .A2(n1085), .A3(n4600), .A4(n1205), .Y(n443)
         );
  AOI22X1_HVT U501 ( .A1(n1042), .A2(n1084), .A3(n1058), .A4(n1203), .Y(n444)
         );
  AOI22X1_HVT U502 ( .A1(n1039), .A2(n1083), .A3(n7600), .A4(n1201), .Y(n445)
         );
  AOI22X1_HVT U503 ( .A1(n5100), .A2(n1082), .A3(n1054), .A4(n1199), .Y(n446)
         );
  AOI22X1_HVT U504 ( .A1(n1044), .A2(n1081), .A3(n7600), .A4(n1197), .Y(n447)
         );
  AOI22X1_HVT U505 ( .A1(n37), .A2(n10801), .A3(n1055), .A4(n1195), .Y(n448)
         );
  AOI22X1_HVT U506 ( .A1(n5300), .A2(n1079), .A3(n4600), .A4(n1193), .Y(n449)
         );
  AOI22X1_HVT U507 ( .A1(n1039), .A2(n1078), .A3(n7600), .A4(n1191), .Y(n4501)
         );
  AOI22X1_HVT U508 ( .A1(n5100), .A2(n1076), .A3(n1056), .A4(n1187), .Y(n451)
         );
  AOI22X1_HVT U509 ( .A1(n1042), .A2(n1075), .A3(n4600), .A4(n1185), .Y(n452)
         );
  AOI22X1_HVT U510 ( .A1(n1039), .A2(n1074), .A3(n1055), .A4(n1183), .Y(n453)
         );
  AOI22X1_HVT U511 ( .A1(n1043), .A2(n1073), .A3(n35), .A4(n1181), .Y(n454) );
  AOI22X1_HVT U512 ( .A1(n38), .A2(n1072), .A3(n5000), .A4(n1179), .Y(n455) );
  AOI22X1_HVT U513 ( .A1(n37), .A2(n1071), .A3(n1056), .A4(n1177), .Y(n456) );
  AOI22X1_HVT U514 ( .A1(n10401), .A2(n10701), .A3(n5000), .A4(n1175), .Y(n457) );
  AOI22X1_HVT U515 ( .A1(n1041), .A2(n1069), .A3(n1058), .A4(n1173), .Y(n458)
         );
  AOI22X1_HVT U516 ( .A1(n37), .A2(n1068), .A3(n7600), .A4(n1171), .Y(n459) );
  AOI22X1_HVT U517 ( .A1(n1042), .A2(n1067), .A3(n4600), .A4(n1169), .Y(n4601)
         );
  AOI22X1_HVT U518 ( .A1(n1044), .A2(n1066), .A3(n5000), .A4(n1167), .Y(n461)
         );
  AOI22X1_HVT U519 ( .A1(sram_rdata_0[0]), .A2(n1354), .A3(sram_rdata_2[0]), 
        .A4(n4300), .Y(n462) );
  AOI22X1_HVT U520 ( .A1(sram_rdata_0[0]), .A2(n1355), .A3(sram_rdata_1[0]), 
        .A4(n29), .Y(n463) );
  AOI22X1_HVT U521 ( .A1(sram_rdata_1[0]), .A2(n1027), .A3(sram_rdata_2[0]), 
        .A4(n1354), .Y(n464) );
  AOI22X1_HVT U522 ( .A1(sram_rdata_3[0]), .A2(n26), .A3(sram_rdata_5[0]), 
        .A4(n4400), .Y(n465) );
  AOI22X1_HVT U523 ( .A1(sram_rdata_3[0]), .A2(n30), .A3(sram_rdata_4[0]), 
        .A4(n26), .Y(n466) );
  AOI22X1_HVT U524 ( .A1(sram_rdata_4[0]), .A2(n1027), .A3(sram_rdata_5[0]), 
        .A4(n1035), .Y(n467) );
  AOI22X1_HVT U525 ( .A1(sram_rdata_6[0]), .A2(n1035), .A3(n32), .A4(
        sram_rdata_8[0]), .Y(n468) );
  AOI22X1_HVT U526 ( .A1(sram_rdata_6[0]), .A2(n4400), .A3(sram_rdata_7[0]), 
        .A4(n1034), .Y(n469) );
  AOI22X1_HVT U527 ( .A1(n4500), .A2(sram_rdata_2[31]), .A3(n28), .A4(
        sram_rdata_0[31]), .Y(n4701) );
  AOI22X1_HVT U528 ( .A1(n1028), .A2(sram_rdata_2[30]), .A3(n1036), .A4(
        sram_rdata_0[30]), .Y(n471) );
  AOI22X1_HVT U529 ( .A1(n4300), .A2(sram_rdata_2[29]), .A3(n28), .A4(
        sram_rdata_0[29]), .Y(n472) );
  AOI22X1_HVT U530 ( .A1(n1355), .A2(sram_rdata_2[28]), .A3(n29), .A4(
        sram_rdata_0[28]), .Y(n473) );
  AOI22X1_HVT U531 ( .A1(n4500), .A2(sram_rdata_2[27]), .A3(n4100), .A4(
        sram_rdata_0[27]), .Y(n474) );
  AOI22X1_HVT U532 ( .A1(n1028), .A2(sram_rdata_2[26]), .A3(n1354), .A4(
        sram_rdata_0[26]), .Y(n475) );
  AOI22X1_HVT U533 ( .A1(n1027), .A2(sram_rdata_2[25]), .A3(n4000), .A4(
        sram_rdata_0[25]), .Y(n476) );
  AOI22X1_HVT U534 ( .A1(n4400), .A2(sram_rdata_2[24]), .A3(n1038), .A4(
        sram_rdata_0[24]), .Y(n477) );
  AOI22X1_HVT U535 ( .A1(n31), .A2(sram_rdata_2[23]), .A3(n4000), .A4(
        sram_rdata_0[23]), .Y(n478) );
  AOI22X1_HVT U536 ( .A1(n1028), .A2(sram_rdata_2[22]), .A3(n1035), .A4(
        sram_rdata_0[22]), .Y(n479) );
  AOI22X1_HVT U537 ( .A1(n32), .A2(sram_rdata_2[21]), .A3(n1036), .A4(
        sram_rdata_0[21]), .Y(n4801) );
  AOI22X1_HVT U538 ( .A1(n1355), .A2(sram_rdata_2[20]), .A3(n4200), .A4(
        sram_rdata_0[20]), .Y(n481) );
  AOI22X1_HVT U539 ( .A1(n4300), .A2(sram_rdata_2[19]), .A3(n4100), .A4(
        sram_rdata_0[19]), .Y(n482) );
  AOI22X1_HVT U540 ( .A1(n4500), .A2(sram_rdata_2[18]), .A3(n1354), .A4(
        sram_rdata_0[18]), .Y(n483) );
  AOI22X1_HVT U541 ( .A1(n1027), .A2(sram_rdata_2[17]), .A3(n4000), .A4(
        sram_rdata_0[17]), .Y(n484) );
  AOI22X1_HVT U542 ( .A1(n30), .A2(sram_rdata_2[16]), .A3(n1035), .A4(
        sram_rdata_0[16]), .Y(n485) );
  AOI22X1_HVT U543 ( .A1(n1029), .A2(sram_rdata_0[31]), .A3(n1034), .A4(
        sram_rdata_1[31]), .Y(n486) );
  AOI22X1_HVT U544 ( .A1(n30), .A2(sram_rdata_0[30]), .A3(n4200), .A4(
        sram_rdata_1[30]), .Y(n487) );
  AOI22X1_HVT U545 ( .A1(n4500), .A2(sram_rdata_0[29]), .A3(n4100), .A4(
        sram_rdata_1[29]), .Y(n488) );
  AOI22X1_HVT U546 ( .A1(n1028), .A2(sram_rdata_0[28]), .A3(n1035), .A4(
        sram_rdata_1[28]), .Y(n489) );
  AOI22X1_HVT U547 ( .A1(n4300), .A2(sram_rdata_0[27]), .A3(n1034), .A4(
        sram_rdata_1[27]), .Y(n4901) );
  AOI22X1_HVT U548 ( .A1(n1355), .A2(sram_rdata_0[26]), .A3(n4200), .A4(
        sram_rdata_1[26]), .Y(n491) );
  AOI22X1_HVT U549 ( .A1(n31), .A2(sram_rdata_0[25]), .A3(n1038), .A4(
        sram_rdata_1[25]), .Y(n492) );
  AOI22X1_HVT U550 ( .A1(n1026), .A2(sram_rdata_0[24]), .A3(n4000), .A4(
        sram_rdata_1[24]), .Y(n493) );
  AOI22X1_HVT U551 ( .A1(n1029), .A2(sram_rdata_0[23]), .A3(n1037), .A4(
        sram_rdata_1[23]), .Y(n494) );
  AOI22X1_HVT U552 ( .A1(n4400), .A2(sram_rdata_0[22]), .A3(n4100), .A4(
        sram_rdata_1[22]), .Y(n495) );
  AOI22X1_HVT U553 ( .A1(n4500), .A2(sram_rdata_0[21]), .A3(n1354), .A4(
        sram_rdata_1[21]), .Y(n496) );
  AOI22X1_HVT U554 ( .A1(n1028), .A2(sram_rdata_0[20]), .A3(n1034), .A4(
        sram_rdata_1[20]), .Y(n497) );
  AOI22X1_HVT U555 ( .A1(n32), .A2(sram_rdata_0[17]), .A3(n1038), .A4(
        sram_rdata_1[17]), .Y(n498) );
  AOI22X1_HVT U556 ( .A1(n32), .A2(sram_rdata_0[16]), .A3(n26), .A4(
        sram_rdata_1[16]), .Y(n499) );
  AOI22X1_HVT U557 ( .A1(n1029), .A2(sram_rdata_1[31]), .A3(n1037), .A4(
        sram_rdata_2[31]), .Y(n5001) );
  AOI22X1_HVT U558 ( .A1(n30), .A2(sram_rdata_1[30]), .A3(n1034), .A4(
        sram_rdata_2[30]), .Y(n501) );
  AOI22X1_HVT U559 ( .A1(n30), .A2(sram_rdata_1[28]), .A3(n4100), .A4(
        sram_rdata_2[28]), .Y(n502) );
  AOI22X1_HVT U560 ( .A1(n31), .A2(sram_rdata_1[27]), .A3(n1354), .A4(
        sram_rdata_2[27]), .Y(n503) );
  AOI22X1_HVT U561 ( .A1(n1026), .A2(sram_rdata_1[26]), .A3(n4000), .A4(
        sram_rdata_2[26]), .Y(n504) );
  AOI22X1_HVT U562 ( .A1(n4300), .A2(sram_rdata_1[25]), .A3(n1035), .A4(
        sram_rdata_2[25]), .Y(n505) );
  AOI22X1_HVT U563 ( .A1(n1355), .A2(sram_rdata_1[24]), .A3(n1034), .A4(
        sram_rdata_2[24]), .Y(n506) );
  AOI22X1_HVT U564 ( .A1(n4500), .A2(sram_rdata_1[23]), .A3(n26), .A4(
        sram_rdata_2[23]), .Y(n507) );
  AOI22X1_HVT U565 ( .A1(n1028), .A2(sram_rdata_1[22]), .A3(n1035), .A4(
        sram_rdata_2[22]), .Y(n508) );
  AOI22X1_HVT U566 ( .A1(n1029), .A2(sram_rdata_1[21]), .A3(n1036), .A4(
        sram_rdata_2[21]), .Y(n509) );
  AOI22X1_HVT U567 ( .A1(n4400), .A2(sram_rdata_1[20]), .A3(n28), .A4(
        sram_rdata_2[20]), .Y(n5101) );
  AOI22X1_HVT U568 ( .A1(n31), .A2(sram_rdata_1[19]), .A3(n4100), .A4(
        sram_rdata_2[19]), .Y(n511) );
  AOI22X1_HVT U569 ( .A1(n1026), .A2(sram_rdata_1[18]), .A3(n4200), .A4(
        sram_rdata_2[18]), .Y(n512) );
  AOI22X1_HVT U570 ( .A1(n4300), .A2(sram_rdata_1[17]), .A3(n29), .A4(
        sram_rdata_2[17]), .Y(n513) );
  AOI22X1_HVT U571 ( .A1(n32), .A2(sram_rdata_1[16]), .A3(n1038), .A4(
        sram_rdata_2[16]), .Y(n514) );
  AOI22X1_HVT U572 ( .A1(n32), .A2(sram_rdata_2[15]), .A3(n26), .A4(
        sram_rdata_0[15]), .Y(n515) );
  AOI22X1_HVT U573 ( .A1(n4400), .A2(sram_rdata_2[14]), .A3(n1037), .A4(
        sram_rdata_0[14]), .Y(n516) );
  AOI22X1_HVT U574 ( .A1(n1029), .A2(sram_rdata_2[13]), .A3(n1034), .A4(
        sram_rdata_0[13]), .Y(n517) );
  AOI22X1_HVT U575 ( .A1(n4400), .A2(sram_rdata_2[12]), .A3(n28), .A4(
        sram_rdata_0[12]), .Y(n518) );
  AOI22X1_HVT U576 ( .A1(n1027), .A2(sram_rdata_2[11]), .A3(n29), .A4(
        sram_rdata_0[11]), .Y(n519) );
  AOI22X1_HVT U577 ( .A1(n4400), .A2(sram_rdata_2[10]), .A3(n1354), .A4(
        sram_rdata_0[10]), .Y(n5201) );
  AOI22X1_HVT U578 ( .A1(n31), .A2(sram_rdata_2[9]), .A3(n4000), .A4(
        sram_rdata_0[9]), .Y(n521) );
  AOI22X1_HVT U579 ( .A1(n1028), .A2(sram_rdata_2[8]), .A3(n1354), .A4(
        sram_rdata_0[8]), .Y(n522) );
  AOI22X1_HVT U580 ( .A1(n32), .A2(sram_rdata_2[7]), .A3(n26), .A4(
        sram_rdata_0[7]), .Y(n523) );
  AOI22X1_HVT U581 ( .A1(n4400), .A2(sram_rdata_2[6]), .A3(n1037), .A4(
        sram_rdata_0[6]), .Y(n524) );
  AOI22X1_HVT U582 ( .A1(n31), .A2(sram_rdata_2[5]), .A3(n1037), .A4(
        sram_rdata_0[5]), .Y(n525) );
  AOI22X1_HVT U583 ( .A1(n1028), .A2(sram_rdata_2[4]), .A3(n1036), .A4(
        sram_rdata_0[4]), .Y(n526) );
  AOI22X1_HVT U584 ( .A1(n1027), .A2(sram_rdata_2[3]), .A3(n4200), .A4(
        sram_rdata_0[3]), .Y(n527) );
  AOI22X1_HVT U585 ( .A1(n4400), .A2(sram_rdata_2[2]), .A3(n1034), .A4(
        sram_rdata_0[2]), .Y(n528) );
  AOI22X1_HVT U586 ( .A1(n31), .A2(sram_rdata_2[1]), .A3(n4200), .A4(
        sram_rdata_0[1]), .Y(n529) );
  AOI22X1_HVT U587 ( .A1(n1026), .A2(sram_rdata_0[15]), .A3(n29), .A4(
        sram_rdata_1[15]), .Y(n5301) );
  AOI22X1_HVT U588 ( .A1(n4300), .A2(sram_rdata_0[14]), .A3(n1038), .A4(
        sram_rdata_1[14]), .Y(n531) );
  AOI22X1_HVT U589 ( .A1(n1355), .A2(sram_rdata_0[13]), .A3(n26), .A4(
        sram_rdata_1[13]), .Y(n532) );
  AOI22X1_HVT U590 ( .A1(n4300), .A2(sram_rdata_0[12]), .A3(n1035), .A4(
        sram_rdata_1[12]), .Y(n533) );
  AOI22X1_HVT U591 ( .A1(n1355), .A2(sram_rdata_0[11]), .A3(n1034), .A4(
        sram_rdata_1[11]), .Y(n534) );
  AOI22X1_HVT U592 ( .A1(n1029), .A2(sram_rdata_0[10]), .A3(n4200), .A4(
        sram_rdata_1[10]), .Y(n535) );
  AOI22X1_HVT U593 ( .A1(n4400), .A2(sram_rdata_0[9]), .A3(n29), .A4(
        sram_rdata_1[9]), .Y(n536) );
  AOI22X1_HVT U594 ( .A1(n1029), .A2(sram_rdata_0[8]), .A3(n1038), .A4(
        sram_rdata_1[8]), .Y(n537) );
  AOI22X1_HVT U595 ( .A1(n30), .A2(sram_rdata_0[7]), .A3(n4000), .A4(
        sram_rdata_1[7]), .Y(n538) );
  AOI22X1_HVT U596 ( .A1(n31), .A2(sram_rdata_0[6]), .A3(n1035), .A4(
        sram_rdata_1[6]), .Y(n539) );
  AOI22X1_HVT U597 ( .A1(n1026), .A2(sram_rdata_0[5]), .A3(n29), .A4(
        sram_rdata_1[5]), .Y(n5401) );
  AOI22X1_HVT U598 ( .A1(n4300), .A2(sram_rdata_0[4]), .A3(n1038), .A4(
        sram_rdata_1[4]), .Y(n541) );
  AOI22X1_HVT U599 ( .A1(n1355), .A2(sram_rdata_0[3]), .A3(n4000), .A4(
        sram_rdata_1[3]), .Y(n542) );
  AOI22X1_HVT U600 ( .A1(n31), .A2(sram_rdata_0[2]), .A3(n1034), .A4(
        sram_rdata_1[2]), .Y(n543) );
  AOI22X1_HVT U601 ( .A1(n1026), .A2(sram_rdata_0[1]), .A3(n28), .A4(
        sram_rdata_1[1]), .Y(n544) );
  AOI22X1_HVT U602 ( .A1(n1027), .A2(sram_rdata_1[15]), .A3(n29), .A4(
        sram_rdata_2[15]), .Y(n545) );
  AOI22X1_HVT U603 ( .A1(n30), .A2(sram_rdata_1[14]), .A3(n1037), .A4(
        sram_rdata_2[14]), .Y(n546) );
  AOI22X1_HVT U604 ( .A1(n4500), .A2(sram_rdata_1[13]), .A3(n1036), .A4(
        sram_rdata_2[13]), .Y(n547) );
  AOI22X1_HVT U605 ( .A1(n1028), .A2(sram_rdata_1[12]), .A3(n1354), .A4(
        sram_rdata_2[12]), .Y(n548) );
  AOI22X1_HVT U606 ( .A1(n32), .A2(sram_rdata_1[11]), .A3(n4000), .A4(
        sram_rdata_2[11]), .Y(n549) );
  AOI22X1_HVT U607 ( .A1(n30), .A2(sram_rdata_1[10]), .A3(n1037), .A4(
        sram_rdata_2[10]), .Y(n5501) );
  AOI22X1_HVT U608 ( .A1(n32), .A2(sram_rdata_1[9]), .A3(n1034), .A4(
        sram_rdata_2[9]), .Y(n551) );
  AOI22X1_HVT U609 ( .A1(n1355), .A2(sram_rdata_1[8]), .A3(n4200), .A4(
        sram_rdata_2[8]), .Y(n552) );
  AOI22X1_HVT U610 ( .A1(n1027), .A2(sram_rdata_1[7]), .A3(n4100), .A4(
        sram_rdata_2[7]), .Y(n553) );
  AOI22X1_HVT U611 ( .A1(n30), .A2(sram_rdata_1[6]), .A3(n1038), .A4(
        sram_rdata_2[6]), .Y(n554) );
  AOI22X1_HVT U612 ( .A1(n1027), .A2(sram_rdata_1[5]), .A3(n4000), .A4(
        sram_rdata_2[5]), .Y(n555) );
  AOI22X1_HVT U613 ( .A1(n4400), .A2(sram_rdata_1[4]), .A3(n1035), .A4(
        sram_rdata_2[4]), .Y(n556) );
  AOI22X1_HVT U614 ( .A1(n4500), .A2(sram_rdata_1[3]), .A3(n1036), .A4(
        sram_rdata_2[3]), .Y(n557) );
  AOI22X1_HVT U615 ( .A1(n1026), .A2(sram_rdata_1[2]), .A3(n28), .A4(
        sram_rdata_2[2]), .Y(n558) );
  AOI22X1_HVT U616 ( .A1(n4300), .A2(sram_rdata_1[1]), .A3(n4100), .A4(
        sram_rdata_2[1]), .Y(n559) );
  AOI22X1_HVT U617 ( .A1(n30), .A2(sram_rdata_5[31]), .A3(n1038), .A4(
        sram_rdata_3[31]), .Y(n5601) );
  AOI22X1_HVT U618 ( .A1(n31), .A2(sram_rdata_5[30]), .A3(n28), .A4(
        sram_rdata_3[30]), .Y(n561) );
  AOI22X1_HVT U619 ( .A1(n1026), .A2(sram_rdata_5[29]), .A3(n4100), .A4(
        sram_rdata_3[29]), .Y(n562) );
  AOI22X1_HVT U620 ( .A1(n1029), .A2(sram_rdata_5[28]), .A3(n1354), .A4(
        sram_rdata_3[28]), .Y(n563) );
  AOI22X1_HVT U621 ( .A1(n30), .A2(sram_rdata_5[27]), .A3(n26), .A4(
        sram_rdata_3[27]), .Y(n564) );
  AOI22X1_HVT U622 ( .A1(n4500), .A2(sram_rdata_5[26]), .A3(n1035), .A4(
        sram_rdata_3[26]), .Y(n565) );
  AOI22X1_HVT U623 ( .A1(n1026), .A2(sram_rdata_5[25]), .A3(n26), .A4(
        sram_rdata_3[25]), .Y(n566) );
  AOI22X1_HVT U624 ( .A1(n32), .A2(sram_rdata_5[24]), .A3(n1035), .A4(
        sram_rdata_3[24]), .Y(n567) );
  AOI22X1_HVT U625 ( .A1(n4400), .A2(sram_rdata_5[23]), .A3(n1036), .A4(
        sram_rdata_3[23]), .Y(n568) );
  AOI22X1_HVT U626 ( .A1(n32), .A2(sram_rdata_5[22]), .A3(n28), .A4(
        sram_rdata_3[22]), .Y(n569) );
  AOI22X1_HVT U627 ( .A1(n1355), .A2(sram_rdata_5[21]), .A3(n4100), .A4(
        sram_rdata_3[21]), .Y(n5701) );
  AOI22X1_HVT U628 ( .A1(n1029), .A2(sram_rdata_5[20]), .A3(n1038), .A4(
        sram_rdata_3[20]), .Y(n571) );
  AOI22X1_HVT U629 ( .A1(n30), .A2(sram_rdata_5[19]), .A3(n4000), .A4(
        sram_rdata_3[19]), .Y(n572) );
  AOI22X1_HVT U630 ( .A1(n1029), .A2(sram_rdata_5[18]), .A3(n1037), .A4(
        sram_rdata_3[18]), .Y(n573) );
  AOI22X1_HVT U631 ( .A1(n4400), .A2(sram_rdata_5[17]), .A3(n1036), .A4(
        sram_rdata_3[17]), .Y(n574) );
  AOI22X1_HVT U632 ( .A1(n31), .A2(sram_rdata_5[16]), .A3(n28), .A4(
        sram_rdata_3[16]), .Y(n575) );
  AOI22X1_HVT U633 ( .A1(n1028), .A2(sram_rdata_3[31]), .A3(n1034), .A4(
        sram_rdata_4[31]), .Y(n576) );
  AOI22X1_HVT U634 ( .A1(n32), .A2(sram_rdata_3[30]), .A3(n4200), .A4(
        sram_rdata_4[30]), .Y(n577) );
  AOI22X1_HVT U635 ( .A1(n1355), .A2(sram_rdata_3[29]), .A3(n4100), .A4(
        sram_rdata_4[29]), .Y(n578) );
  AOI22X1_HVT U636 ( .A1(n4500), .A2(sram_rdata_3[28]), .A3(n29), .A4(
        sram_rdata_4[28]), .Y(n579) );
  AOI22X1_HVT U637 ( .A1(n1028), .A2(sram_rdata_3[27]), .A3(n1038), .A4(
        sram_rdata_4[27]), .Y(n5801) );
  AOI22X1_HVT U638 ( .A1(n1027), .A2(sram_rdata_3[26]), .A3(n26), .A4(
        sram_rdata_4[26]), .Y(n581) );
  AOI22X1_HVT U639 ( .A1(n30), .A2(sram_rdata_3[25]), .A3(n1038), .A4(
        sram_rdata_4[25]), .Y(n582) );
  AOI22X1_HVT U640 ( .A1(n31), .A2(sram_rdata_3[24]), .A3(n4000), .A4(
        sram_rdata_4[24]), .Y(n583) );
  AOI22X1_HVT U641 ( .A1(n1028), .A2(sram_rdata_3[23]), .A3(n1037), .A4(
        sram_rdata_4[23]), .Y(n584) );
  AOI22X1_HVT U642 ( .A1(n4300), .A2(sram_rdata_3[22]), .A3(n1036), .A4(
        sram_rdata_4[22]), .Y(n585) );
  AOI22X1_HVT U643 ( .A1(n1355), .A2(sram_rdata_3[21]), .A3(n4200), .A4(
        sram_rdata_4[21]), .Y(n586) );
  AOI22X1_HVT U644 ( .A1(n4300), .A2(sram_rdata_3[20]), .A3(n29), .A4(
        sram_rdata_4[20]), .Y(n587) );
  AOI22X1_HVT U645 ( .A1(n4500), .A2(sram_rdata_3[19]), .A3(n1038), .A4(
        sram_rdata_4[19]), .Y(n588) );
  AOI22X1_HVT U646 ( .A1(n1027), .A2(sram_rdata_3[18]), .A3(n26), .A4(
        sram_rdata_4[18]), .Y(n589) );
  AOI22X1_HVT U647 ( .A1(n4400), .A2(sram_rdata_3[17]), .A3(n1037), .A4(
        sram_rdata_4[17]), .Y(n5901) );
  AOI22X1_HVT U648 ( .A1(n1029), .A2(sram_rdata_3[16]), .A3(n1036), .A4(
        sram_rdata_4[16]), .Y(n591) );
  AOI22X1_HVT U649 ( .A1(n30), .A2(sram_rdata_4[31]), .A3(n28), .A4(
        sram_rdata_5[31]), .Y(n592) );
  AOI22X1_HVT U650 ( .A1(n31), .A2(sram_rdata_4[30]), .A3(n29), .A4(
        sram_rdata_5[30]), .Y(n593) );
  AOI22X1_HVT U651 ( .A1(n1028), .A2(sram_rdata_4[29]), .A3(n1037), .A4(
        sram_rdata_5[29]), .Y(n594) );
  AOI22X1_HVT U652 ( .A1(n32), .A2(sram_rdata_4[28]), .A3(n1034), .A4(
        sram_rdata_5[28]), .Y(n595) );
  AOI22X1_HVT U653 ( .A1(n1355), .A2(sram_rdata_4[27]), .A3(n4200), .A4(
        sram_rdata_5[27]), .Y(n596) );
  AOI22X1_HVT U654 ( .A1(n4500), .A2(sram_rdata_4[26]), .A3(n1038), .A4(
        sram_rdata_5[26]), .Y(n597) );
  AOI22X1_HVT U655 ( .A1(n1026), .A2(sram_rdata_4[25]), .A3(n26), .A4(
        sram_rdata_5[25]), .Y(n598) );
  AOI22X1_HVT U656 ( .A1(n1029), .A2(sram_rdata_4[24]), .A3(n1035), .A4(
        sram_rdata_5[24]), .Y(n599) );
  AOI22X1_HVT U657 ( .A1(n4500), .A2(sram_rdata_4[22]), .A3(n1354), .A4(
        sram_rdata_5[22]), .Y(n6001) );
  AOI22X1_HVT U658 ( .A1(n1028), .A2(sram_rdata_4[21]), .A3(n1034), .A4(
        sram_rdata_5[21]), .Y(n601) );
  AOI22X1_HVT U659 ( .A1(n4300), .A2(sram_rdata_4[20]), .A3(n4200), .A4(
        sram_rdata_5[20]), .Y(n602) );
  AOI22X1_HVT U660 ( .A1(n1355), .A2(sram_rdata_4[19]), .A3(n4100), .A4(
        sram_rdata_5[19]), .Y(n603) );
  AOI22X1_HVT U661 ( .A1(n32), .A2(sram_rdata_4[18]), .A3(n1354), .A4(
        sram_rdata_5[18]), .Y(n604) );
  AOI22X1_HVT U662 ( .A1(n1355), .A2(sram_rdata_4[17]), .A3(n26), .A4(
        sram_rdata_5[17]), .Y(n605) );
  AOI22X1_HVT U663 ( .A1(n1029), .A2(sram_rdata_4[16]), .A3(n1037), .A4(
        sram_rdata_5[16]), .Y(n606) );
  AOI22X1_HVT U664 ( .A1(n4400), .A2(sram_rdata_5[15]), .A3(n1036), .A4(
        sram_rdata_3[15]), .Y(n607) );
  AOI22X1_HVT U665 ( .A1(n1029), .A2(sram_rdata_5[14]), .A3(n28), .A4(
        sram_rdata_3[14]), .Y(n608) );
  AOI22X1_HVT U666 ( .A1(n30), .A2(sram_rdata_5[13]), .A3(n29), .A4(
        sram_rdata_3[13]), .Y(n609) );
  AOI22X1_HVT U667 ( .A1(n31), .A2(sram_rdata_5[12]), .A3(n1354), .A4(
        sram_rdata_3[12]), .Y(n6101) );
  AOI22X1_HVT U668 ( .A1(n1026), .A2(sram_rdata_5[11]), .A3(n4000), .A4(
        sram_rdata_3[11]), .Y(n611) );
  AOI22X1_HVT U669 ( .A1(n32), .A2(sram_rdata_5[10]), .A3(n1037), .A4(
        sram_rdata_3[10]), .Y(n612) );
  AOI22X1_HVT U670 ( .A1(n30), .A2(sram_rdata_5[9]), .A3(n1036), .A4(
        sram_rdata_3[9]), .Y(n613) );
  AOI22X1_HVT U671 ( .A1(n31), .A2(sram_rdata_5[8]), .A3(n4000), .A4(
        sram_rdata_3[8]), .Y(n614) );
  AOI22X1_HVT U672 ( .A1(n1028), .A2(sram_rdata_5[7]), .A3(n1035), .A4(
        sram_rdata_3[7]), .Y(n615) );
  AOI22X1_HVT U673 ( .A1(n1029), .A2(sram_rdata_5[6]), .A3(n1034), .A4(
        sram_rdata_3[6]), .Y(n616) );
  AOI22X1_HVT U674 ( .A1(n4400), .A2(sram_rdata_5[5]), .A3(n28), .A4(
        sram_rdata_3[5]), .Y(n617) );
  AOI22X1_HVT U675 ( .A1(n4500), .A2(sram_rdata_5[4]), .A3(n4100), .A4(
        sram_rdata_3[4]), .Y(n618) );
  AOI22X1_HVT U676 ( .A1(n1026), .A2(sram_rdata_5[3]), .A3(n28), .A4(
        sram_rdata_3[3]), .Y(n619) );
  AOI22X1_HVT U677 ( .A1(n4300), .A2(sram_rdata_5[2]), .A3(n4100), .A4(
        sram_rdata_3[2]), .Y(n6201) );
  AOI22X1_HVT U678 ( .A1(n4500), .A2(sram_rdata_5[1]), .A3(n1038), .A4(
        sram_rdata_3[1]), .Y(n621) );
  AOI22X1_HVT U679 ( .A1(n32), .A2(sram_rdata_3[15]), .A3(n26), .A4(
        sram_rdata_4[15]), .Y(n622) );
  AOI22X1_HVT U680 ( .A1(n4300), .A2(sram_rdata_3[14]), .A3(n1037), .A4(
        sram_rdata_4[14]), .Y(n623) );
  AOI22X1_HVT U681 ( .A1(n1029), .A2(sram_rdata_3[13]), .A3(n1034), .A4(
        sram_rdata_4[13]), .Y(n624) );
  AOI22X1_HVT U682 ( .A1(n4400), .A2(sram_rdata_3[12]), .A3(n4200), .A4(
        sram_rdata_4[12]), .Y(n625) );
  AOI22X1_HVT U683 ( .A1(n1027), .A2(sram_rdata_3[11]), .A3(n4100), .A4(
        sram_rdata_4[11]), .Y(n626) );
  AOI22X1_HVT U684 ( .A1(n4500), .A2(sram_rdata_3[9]), .A3(n4000), .A4(
        sram_rdata_4[9]), .Y(n627) );
  AOI22X1_HVT U685 ( .A1(n1028), .A2(sram_rdata_3[8]), .A3(n1354), .A4(
        sram_rdata_4[8]), .Y(n628) );
  AOI22X1_HVT U686 ( .A1(n32), .A2(sram_rdata_3[7]), .A3(n4000), .A4(
        sram_rdata_4[7]), .Y(n629) );
  AOI22X1_HVT U687 ( .A1(n31), .A2(sram_rdata_3[6]), .A3(n1037), .A4(
        sram_rdata_4[6]), .Y(n6301) );
  AOI22X1_HVT U688 ( .A1(n31), .A2(sram_rdata_3[5]), .A3(n1037), .A4(
        sram_rdata_4[5]), .Y(n631) );
  AOI22X1_HVT U689 ( .A1(n1028), .A2(sram_rdata_3[4]), .A3(n1034), .A4(
        sram_rdata_4[4]), .Y(n632) );
  AOI22X1_HVT U690 ( .A1(n1029), .A2(sram_rdata_3[3]), .A3(n4200), .A4(
        sram_rdata_4[3]), .Y(n633) );
  AOI22X1_HVT U691 ( .A1(n4400), .A2(sram_rdata_3[2]), .A3(n1034), .A4(
        sram_rdata_4[2]), .Y(n634) );
  AOI22X1_HVT U692 ( .A1(n31), .A2(sram_rdata_3[1]), .A3(n4200), .A4(
        sram_rdata_4[1]), .Y(n635) );
  AOI22X1_HVT U693 ( .A1(n1026), .A2(sram_rdata_4[15]), .A3(n29), .A4(
        sram_rdata_5[15]), .Y(n636) );
  AOI22X1_HVT U694 ( .A1(n32), .A2(sram_rdata_4[14]), .A3(n1038), .A4(
        sram_rdata_5[14]), .Y(n637) );
  AOI22X1_HVT U695 ( .A1(n31), .A2(sram_rdata_4[13]), .A3(n4000), .A4(
        sram_rdata_5[13]), .Y(n638) );
  AOI22X1_HVT U696 ( .A1(n4300), .A2(sram_rdata_4[12]), .A3(n1037), .A4(
        sram_rdata_5[12]), .Y(n639) );
  AOI22X1_HVT U697 ( .A1(n1355), .A2(sram_rdata_4[11]), .A3(n1034), .A4(
        sram_rdata_5[11]), .Y(n6401) );
  AOI22X1_HVT U698 ( .A1(n1029), .A2(sram_rdata_4[10]), .A3(n4200), .A4(
        sram_rdata_5[10]), .Y(n641) );
  AOI22X1_HVT U699 ( .A1(n30), .A2(sram_rdata_4[9]), .A3(n29), .A4(
        sram_rdata_5[9]), .Y(n642) );
  AOI22X1_HVT U700 ( .A1(n1029), .A2(sram_rdata_4[8]), .A3(n1038), .A4(
        sram_rdata_5[8]), .Y(n643) );
  AOI22X1_HVT U701 ( .A1(n30), .A2(sram_rdata_4[7]), .A3(n4000), .A4(
        sram_rdata_5[7]), .Y(n644) );
  AOI22X1_HVT U702 ( .A1(n31), .A2(sram_rdata_4[6]), .A3(n1035), .A4(
        sram_rdata_5[6]), .Y(n645) );
  AOI22X1_HVT U703 ( .A1(n1026), .A2(sram_rdata_4[5]), .A3(n4100), .A4(
        sram_rdata_5[5]), .Y(n646) );
  AOI22X1_HVT U704 ( .A1(n4300), .A2(sram_rdata_4[4]), .A3(n1038), .A4(
        sram_rdata_5[4]), .Y(n647) );
  AOI22X1_HVT U705 ( .A1(n1355), .A2(sram_rdata_4[3]), .A3(n26), .A4(
        sram_rdata_5[3]), .Y(n648) );
  AOI22X1_HVT U706 ( .A1(n4500), .A2(sram_rdata_4[2]), .A3(n1034), .A4(
        sram_rdata_5[2]), .Y(n649) );
  AOI22X1_HVT U707 ( .A1(n1028), .A2(sram_rdata_4[1]), .A3(n28), .A4(
        sram_rdata_5[1]), .Y(n6501) );
  AOI22X1_HVT U708 ( .A1(n1027), .A2(sram_rdata_8[31]), .A3(n29), .A4(
        sram_rdata_6[31]), .Y(n651) );
  AOI22X1_HVT U709 ( .A1(n30), .A2(sram_rdata_8[30]), .A3(n1037), .A4(
        sram_rdata_6[30]), .Y(n652) );
  AOI22X1_HVT U710 ( .A1(n31), .A2(sram_rdata_8[29]), .A3(n1036), .A4(
        sram_rdata_6[29]), .Y(n653) );
  AOI22X1_HVT U711 ( .A1(n1028), .A2(sram_rdata_8[28]), .A3(n1038), .A4(
        sram_rdata_6[28]), .Y(n654) );
  AOI22X1_HVT U712 ( .A1(n32), .A2(sram_rdata_8[27]), .A3(n26), .A4(
        sram_rdata_6[27]), .Y(n655) );
  AOI22X1_HVT U713 ( .A1(n1355), .A2(sram_rdata_8[26]), .A3(n1035), .A4(
        sram_rdata_6[26]), .Y(n656) );
  AOI22X1_HVT U714 ( .A1(n32), .A2(sram_rdata_8[25]), .A3(n1036), .A4(
        sram_rdata_6[25]), .Y(n657) );
  AOI22X1_HVT U715 ( .A1(n1355), .A2(sram_rdata_8[24]), .A3(n28), .A4(
        sram_rdata_6[24]), .Y(n658) );
  AOI22X1_HVT U716 ( .A1(n1027), .A2(sram_rdata_8[23]), .A3(n29), .A4(
        sram_rdata_6[23]), .Y(n659) );
  AOI22X1_HVT U717 ( .A1(n1027), .A2(sram_rdata_8[21]), .A3(n26), .A4(
        sram_rdata_6[21]), .Y(n6601) );
  AOI22X1_HVT U718 ( .A1(n30), .A2(sram_rdata_8[20]), .A3(n1035), .A4(
        sram_rdata_6[20]), .Y(n661) );
  AOI22X1_HVT U719 ( .A1(n4500), .A2(sram_rdata_8[19]), .A3(n1036), .A4(
        sram_rdata_6[19]), .Y(n662) );
  AOI22X1_HVT U720 ( .A1(n1028), .A2(sram_rdata_8[18]), .A3(n28), .A4(
        sram_rdata_6[18]), .Y(n663) );
  AOI22X1_HVT U721 ( .A1(n32), .A2(sram_rdata_8[17]), .A3(n4100), .A4(
        sram_rdata_6[17]), .Y(n664) );
  AOI22X1_HVT U722 ( .A1(n1355), .A2(sram_rdata_8[16]), .A3(n1354), .A4(
        sram_rdata_6[16]), .Y(n665) );
  AOI22X1_HVT U723 ( .A1(n4500), .A2(sram_rdata_6[31]), .A3(n28), .A4(
        sram_rdata_7[31]), .Y(n666) );
  AOI22X1_HVT U724 ( .A1(n1026), .A2(sram_rdata_6[30]), .A3(n4100), .A4(
        sram_rdata_7[30]), .Y(n667) );
  AOI22X1_HVT U725 ( .A1(n1029), .A2(sram_rdata_6[29]), .A3(n1038), .A4(
        sram_rdata_7[29]), .Y(n668) );
  AOI22X1_HVT U726 ( .A1(n30), .A2(sram_rdata_6[28]), .A3(n26), .A4(
        sram_rdata_7[28]), .Y(n669) );
  AOI22X1_HVT U727 ( .A1(n31), .A2(sram_rdata_6[27]), .A3(n1035), .A4(
        sram_rdata_7[27]), .Y(n6701) );
  AOI22X1_HVT U728 ( .A1(n1026), .A2(sram_rdata_6[26]), .A3(n4000), .A4(
        sram_rdata_7[26]), .Y(n671) );
  AOI22X1_HVT U729 ( .A1(n32), .A2(sram_rdata_6[25]), .A3(n1035), .A4(
        sram_rdata_7[25]), .Y(n672) );
  AOI22X1_HVT U730 ( .A1(n31), .A2(sram_rdata_6[24]), .A3(n1036), .A4(
        sram_rdata_7[24]), .Y(n673) );
  AOI22X1_HVT U731 ( .A1(n4300), .A2(sram_rdata_6[23]), .A3(n4200), .A4(
        sram_rdata_7[23]), .Y(n674) );
  AOI22X1_HVT U732 ( .A1(n30), .A2(sram_rdata_6[22]), .A3(n4100), .A4(
        sram_rdata_7[22]), .Y(n675) );
  AOI22X1_HVT U733 ( .A1(n1029), .A2(sram_rdata_6[21]), .A3(n1038), .A4(
        sram_rdata_7[21]), .Y(n676) );
  AOI22X1_HVT U734 ( .A1(n4400), .A2(sram_rdata_6[20]), .A3(n26), .A4(
        sram_rdata_7[20]), .Y(n677) );
  AOI22X1_HVT U735 ( .A1(n1029), .A2(sram_rdata_6[19]), .A3(n1037), .A4(
        sram_rdata_7[19]), .Y(n678) );
  AOI22X1_HVT U736 ( .A1(n4400), .A2(sram_rdata_6[18]), .A3(n1036), .A4(
        sram_rdata_7[18]), .Y(n679) );
  AOI22X1_HVT U737 ( .A1(n31), .A2(sram_rdata_6[17]), .A3(n28), .A4(
        sram_rdata_7[17]), .Y(n6801) );
  AOI22X1_HVT U738 ( .A1(n1028), .A2(sram_rdata_6[16]), .A3(n1036), .A4(
        sram_rdata_7[16]), .Y(n681) );
  AOI22X1_HVT U739 ( .A1(n4300), .A2(sram_rdata_7[31]), .A3(n4200), .A4(
        sram_rdata_8[31]), .Y(n682) );
  AOI22X1_HVT U740 ( .A1(n1355), .A2(sram_rdata_7[30]), .A3(n4100), .A4(
        sram_rdata_8[30]), .Y(n683) );
  AOI22X1_HVT U741 ( .A1(n4500), .A2(sram_rdata_7[29]), .A3(n29), .A4(
        sram_rdata_8[29]), .Y(n684) );
  AOI22X1_HVT U742 ( .A1(n1028), .A2(sram_rdata_7[28]), .A3(n1038), .A4(
        sram_rdata_8[28]), .Y(n685) );
  AOI22X1_HVT U743 ( .A1(n1027), .A2(sram_rdata_7[27]), .A3(n4000), .A4(
        sram_rdata_8[27]), .Y(n686) );
  AOI22X1_HVT U744 ( .A1(n30), .A2(sram_rdata_7[26]), .A3(n1038), .A4(
        sram_rdata_8[26]), .Y(n687) );
  AOI22X1_HVT U745 ( .A1(n4500), .A2(sram_rdata_7[25]), .A3(n26), .A4(
        sram_rdata_8[25]), .Y(n688) );
  AOI22X1_HVT U746 ( .A1(n1028), .A2(sram_rdata_7[24]), .A3(n1035), .A4(
        sram_rdata_8[24]), .Y(n689) );
  AOI22X1_HVT U747 ( .A1(n32), .A2(sram_rdata_7[23]), .A3(n1034), .A4(
        sram_rdata_8[23]), .Y(n6901) );
  AOI22X1_HVT U748 ( .A1(n1355), .A2(sram_rdata_7[22]), .A3(n4200), .A4(
        sram_rdata_8[22]), .Y(n691) );
  AOI22X1_HVT U749 ( .A1(n32), .A2(sram_rdata_7[21]), .A3(n29), .A4(
        sram_rdata_8[21]), .Y(n692) );
  AOI22X1_HVT U750 ( .A1(n1355), .A2(sram_rdata_7[20]), .A3(n1354), .A4(
        sram_rdata_8[20]), .Y(n693) );
  AOI22X1_HVT U751 ( .A1(n1027), .A2(sram_rdata_7[19]), .A3(n4000), .A4(
        sram_rdata_8[19]), .Y(n694) );
  AOI22X1_HVT U752 ( .A1(n30), .A2(sram_rdata_7[18]), .A3(n1037), .A4(
        sram_rdata_8[18]), .Y(n695) );
  AOI22X1_HVT U753 ( .A1(n1029), .A2(sram_rdata_7[17]), .A3(n1036), .A4(
        sram_rdata_8[17]), .Y(n696) );
  AOI22X1_HVT U754 ( .A1(n4500), .A2(sram_rdata_8[15]), .A3(n29), .A4(
        sram_rdata_6[15]), .Y(n697) );
  AOI22X1_HVT U755 ( .A1(n1028), .A2(sram_rdata_8[14]), .A3(n1037), .A4(
        sram_rdata_6[14]), .Y(n698) );
  AOI22X1_HVT U756 ( .A1(n4300), .A2(sram_rdata_8[13]), .A3(n1036), .A4(
        sram_rdata_6[13]), .Y(n699) );
  AOI22X1_HVT U757 ( .A1(n1355), .A2(sram_rdata_8[12]), .A3(n28), .A4(
        sram_rdata_6[12]), .Y(n7001) );
  AOI22X1_HVT U758 ( .A1(n4500), .A2(sram_rdata_8[11]), .A3(n1038), .A4(
        sram_rdata_6[11]), .Y(n701) );
  AOI22X1_HVT U759 ( .A1(n1026), .A2(sram_rdata_8[10]), .A3(n4000), .A4(
        sram_rdata_6[10]), .Y(n702) );
  AOI22X1_HVT U760 ( .A1(n1029), .A2(sram_rdata_8[9]), .A3(n1037), .A4(
        sram_rdata_6[9]), .Y(n703) );
  AOI22X1_HVT U761 ( .A1(n30), .A2(sram_rdata_8[8]), .A3(n29), .A4(
        sram_rdata_6[8]), .Y(n704) );
  AOI22X1_HVT U762 ( .A1(n4500), .A2(sram_rdata_8[7]), .A3(n1354), .A4(
        sram_rdata_6[7]), .Y(n705) );
  AOI22X1_HVT U763 ( .A1(n1028), .A2(sram_rdata_8[6]), .A3(n1036), .A4(
        sram_rdata_6[6]), .Y(n706) );
  AOI22X1_HVT U764 ( .A1(n4300), .A2(sram_rdata_8[5]), .A3(n4200), .A4(
        sram_rdata_6[5]), .Y(n707) );
  AOI22X1_HVT U765 ( .A1(n4300), .A2(sram_rdata_8[4]), .A3(n4100), .A4(
        sram_rdata_6[4]), .Y(n708) );
  AOI22X1_HVT U766 ( .A1(n4300), .A2(sram_rdata_8[3]), .A3(n1354), .A4(
        sram_rdata_6[3]), .Y(n709) );
  AOI22X1_HVT U767 ( .A1(n4500), .A2(sram_rdata_8[2]), .A3(n4000), .A4(
        sram_rdata_6[2]), .Y(n7101) );
  AOI22X1_HVT U768 ( .A1(n1029), .A2(sram_rdata_8[1]), .A3(n1037), .A4(
        sram_rdata_6[1]), .Y(n711) );
  AOI22X1_HVT U769 ( .A1(n4400), .A2(sram_rdata_6[15]), .A3(n1036), .A4(
        sram_rdata_7[15]), .Y(n712) );
  AOI22X1_HVT U770 ( .A1(n1027), .A2(sram_rdata_6[14]), .A3(n4200), .A4(
        sram_rdata_7[14]), .Y(n713) );
  AOI22X1_HVT U771 ( .A1(n30), .A2(sram_rdata_6[13]), .A3(n29), .A4(
        sram_rdata_7[13]), .Y(n714) );
  AOI22X1_HVT U772 ( .A1(n4500), .A2(sram_rdata_6[12]), .A3(n1354), .A4(
        sram_rdata_7[12]), .Y(n715) );
  AOI22X1_HVT U773 ( .A1(n1026), .A2(sram_rdata_6[11]), .A3(n26), .A4(
        sram_rdata_7[11]), .Y(n716) );
  AOI22X1_HVT U774 ( .A1(n4300), .A2(sram_rdata_6[10]), .A3(n1035), .A4(
        sram_rdata_7[10]), .Y(n717) );
  AOI22X1_HVT U775 ( .A1(n4300), .A2(sram_rdata_6[9]), .A3(n1036), .A4(
        sram_rdata_7[9]), .Y(n718) );
  AOI22X1_HVT U776 ( .A1(n31), .A2(sram_rdata_6[8]), .A3(n26), .A4(
        sram_rdata_7[8]), .Y(n719) );
  AOI22X1_HVT U777 ( .A1(n1028), .A2(sram_rdata_6[7]), .A3(n1037), .A4(
        sram_rdata_7[7]), .Y(n7201) );
  AOI22X1_HVT U778 ( .A1(n1029), .A2(sram_rdata_6[6]), .A3(n1036), .A4(
        sram_rdata_7[6]), .Y(n721) );
  AOI22X1_HVT U779 ( .A1(n4400), .A2(sram_rdata_6[5]), .A3(n28), .A4(
        sram_rdata_7[5]), .Y(n722) );
  AOI22X1_HVT U780 ( .A1(n31), .A2(sram_rdata_6[4]), .A3(n4100), .A4(
        sram_rdata_7[4]), .Y(n723) );
  AOI22X1_HVT U781 ( .A1(n1028), .A2(sram_rdata_6[3]), .A3(n28), .A4(
        sram_rdata_7[3]), .Y(n724) );
  AOI22X1_HVT U782 ( .A1(n32), .A2(sram_rdata_6[2]), .A3(n4100), .A4(
        sram_rdata_7[2]), .Y(n725) );
  AOI22X1_HVT U783 ( .A1(n31), .A2(sram_rdata_6[1]), .A3(n1038), .A4(
        sram_rdata_7[1]), .Y(n726) );
  AOI22X1_HVT U784 ( .A1(n32), .A2(sram_rdata_7[15]), .A3(n26), .A4(
        sram_rdata_8[15]), .Y(n727) );
  AOI22X1_HVT U785 ( .A1(n32), .A2(sram_rdata_7[14]), .A3(n1037), .A4(
        sram_rdata_8[14]), .Y(n728) );
  AOI22X1_HVT U786 ( .A1(n1029), .A2(sram_rdata_7[13]), .A3(n1036), .A4(
        sram_rdata_8[13]), .Y(n729) );
  AOI22X1_HVT U787 ( .A1(n1029), .A2(sram_rdata_7[11]), .A3(n29), .A4(
        sram_rdata_8[11]), .Y(n7301) );
  AOI22X1_HVT U788 ( .A1(n4400), .A2(sram_rdata_7[10]), .A3(n1038), .A4(
        sram_rdata_8[10]), .Y(n731) );
  AOI22X1_HVT U789 ( .A1(n31), .A2(sram_rdata_7[9]), .A3(n4000), .A4(
        sram_rdata_8[9]), .Y(n732) );
  AOI22X1_HVT U790 ( .A1(n1028), .A2(sram_rdata_7[8]), .A3(n1354), .A4(
        sram_rdata_8[8]), .Y(n733) );
  AOI22X1_HVT U791 ( .A1(n4300), .A2(sram_rdata_7[7]), .A3(n26), .A4(
        sram_rdata_8[7]), .Y(n734) );
  AOI22X1_HVT U792 ( .A1(n1355), .A2(sram_rdata_7[6]), .A3(n1035), .A4(
        sram_rdata_8[6]), .Y(n735) );
  AOI22X1_HVT U793 ( .A1(n4500), .A2(sram_rdata_7[5]), .A3(n1037), .A4(
        sram_rdata_8[5]), .Y(n736) );
  AOI22X1_HVT U794 ( .A1(n1028), .A2(sram_rdata_7[4]), .A3(n1036), .A4(
        sram_rdata_8[4]), .Y(n737) );
  AOI22X1_HVT U795 ( .A1(n1027), .A2(sram_rdata_7[3]), .A3(n28), .A4(
        sram_rdata_8[3]), .Y(n738) );
  AOI22X1_HVT U796 ( .A1(n30), .A2(sram_rdata_7[2]), .A3(n1034), .A4(
        sram_rdata_8[2]), .Y(n739) );
  AOI22X1_HVT U797 ( .A1(n4500), .A2(sram_rdata_7[1]), .A3(n4200), .A4(
        sram_rdata_8[1]), .Y(n7401) );
  AOI22X1_HVT U798 ( .A1(n1026), .A2(sram_rdata_7[0]), .A3(n29), .A4(
        sram_rdata_8[0]), .Y(n741) );
  NAND2X0_HVT U799 ( .A1(n12300), .A2(sram_rdata_1[31]), .Y(n742) );
  NAND3X0_HVT U800 ( .A1(n1830), .A2(n4701), .A3(n742), .Y(n_src_aox[287]) );
  NAND2X0_HVT U801 ( .A1(n1051), .A2(sram_rdata_1[30]), .Y(n743) );
  NAND3X0_HVT U802 ( .A1(n1840), .A2(n471), .A3(n743), .Y(n_src_aox[286]) );
  NAND2X0_HVT U803 ( .A1(n12900), .A2(sram_rdata_1[29]), .Y(n744) );
  NAND3X0_HVT U804 ( .A1(n1850), .A2(n472), .A3(n744), .Y(n_src_aox[285]) );
  NAND2X0_HVT U805 ( .A1(n1049), .A2(sram_rdata_1[28]), .Y(n745) );
  NAND3X0_HVT U806 ( .A1(n1860), .A2(n473), .A3(n745), .Y(n_src_aox[284]) );
  NAND2X0_HVT U807 ( .A1(n6300), .A2(sram_rdata_1[27]), .Y(n746) );
  NAND3X0_HVT U808 ( .A1(n1870), .A2(n474), .A3(n746), .Y(n_src_aox[283]) );
  NAND2X0_HVT U809 ( .A1(n1049), .A2(sram_rdata_1[26]), .Y(n747) );
  NAND3X0_HVT U810 ( .A1(n1880), .A2(n475), .A3(n747), .Y(n_src_aox[282]) );
  NAND2X0_HVT U811 ( .A1(n1052), .A2(sram_rdata_1[25]), .Y(n748) );
  NAND3X0_HVT U812 ( .A1(n1890), .A2(n476), .A3(n748), .Y(n_src_aox[281]) );
  NAND2X0_HVT U813 ( .A1(n6200), .A2(sram_rdata_1[24]), .Y(n749) );
  NAND3X0_HVT U814 ( .A1(n1900), .A2(n477), .A3(n749), .Y(n_src_aox[280]) );
  NAND2X0_HVT U815 ( .A1(n13300), .A2(sram_rdata_1[23]), .Y(n7501) );
  NAND3X0_HVT U816 ( .A1(n1910), .A2(n478), .A3(n7501), .Y(n_src_aox[279]) );
  NAND2X0_HVT U817 ( .A1(n12500), .A2(sram_rdata_1[22]), .Y(n751) );
  NAND3X0_HVT U818 ( .A1(n1920), .A2(n479), .A3(n751), .Y(n_src_aox[278]) );
  NAND2X0_HVT U819 ( .A1(n13000), .A2(sram_rdata_1[21]), .Y(n752) );
  NAND3X0_HVT U820 ( .A1(n1930), .A2(n4801), .A3(n752), .Y(n_src_aox[277]) );
  NAND2X0_HVT U821 ( .A1(n13400), .A2(sram_rdata_1[20]), .Y(n753) );
  NAND3X0_HVT U822 ( .A1(n1940), .A2(n481), .A3(n753), .Y(n_src_aox[276]) );
  NAND2X0_HVT U823 ( .A1(n12700), .A2(sram_rdata_1[19]), .Y(n754) );
  NAND3X0_HVT U824 ( .A1(n1950), .A2(n482), .A3(n754), .Y(n_src_aox[275]) );
  NAND2X0_HVT U825 ( .A1(n13100), .A2(sram_rdata_1[18]), .Y(n755) );
  NAND3X0_HVT U826 ( .A1(n1960), .A2(n483), .A3(n755), .Y(n_src_aox[274]) );
  NAND2X0_HVT U827 ( .A1(n12200), .A2(sram_rdata_1[17]), .Y(n756) );
  NAND3X0_HVT U828 ( .A1(n1970), .A2(n484), .A3(n756), .Y(n_src_aox[273]) );
  NAND2X0_HVT U829 ( .A1(n1049), .A2(sram_rdata_1[16]), .Y(n757) );
  NAND3X0_HVT U830 ( .A1(n1980), .A2(n485), .A3(n757), .Y(n_src_aox[272]) );
  NAND2X0_HVT U831 ( .A1(n1049), .A2(sram_rdata_2[31]), .Y(n758) );
  NAND3X0_HVT U832 ( .A1(n1990), .A2(n486), .A3(n758), .Y(n_src_aox[271]) );
  NAND2X0_HVT U833 ( .A1(n6000), .A2(sram_rdata_2[30]), .Y(n759) );
  NAND3X0_HVT U834 ( .A1(n2000), .A2(n487), .A3(n759), .Y(n_src_aox[270]) );
  NAND2X0_HVT U835 ( .A1(n1053), .A2(sram_rdata_2[29]), .Y(n7601) );
  NAND3X0_HVT U836 ( .A1(n2010), .A2(n488), .A3(n7601), .Y(n_src_aox[269]) );
  NAND2X0_HVT U837 ( .A1(n12300), .A2(sram_rdata_2[28]), .Y(n761) );
  NAND3X0_HVT U838 ( .A1(n2020), .A2(n489), .A3(n761), .Y(n_src_aox[268]) );
  NAND2X0_HVT U839 ( .A1(n10501), .A2(sram_rdata_2[27]), .Y(n762) );
  NAND3X0_HVT U840 ( .A1(n2030), .A2(n4901), .A3(n762), .Y(n_src_aox[267]) );
  NAND2X0_HVT U841 ( .A1(n12600), .A2(sram_rdata_2[26]), .Y(n763) );
  NAND3X0_HVT U842 ( .A1(n2040), .A2(n491), .A3(n763), .Y(n_src_aox[266]) );
  NAND2X0_HVT U843 ( .A1(n12800), .A2(sram_rdata_2[25]), .Y(n764) );
  NAND3X0_HVT U844 ( .A1(n2050), .A2(n492), .A3(n764), .Y(n_src_aox[265]) );
  NAND2X0_HVT U845 ( .A1(n13200), .A2(sram_rdata_2[24]), .Y(n765) );
  NAND3X0_HVT U846 ( .A1(n2060), .A2(n493), .A3(n765), .Y(n_src_aox[264]) );
  NAND2X0_HVT U847 ( .A1(n6300), .A2(sram_rdata_2[23]), .Y(n766) );
  NAND3X0_HVT U848 ( .A1(n2070), .A2(n494), .A3(n766), .Y(n_src_aox[263]) );
  NAND2X0_HVT U849 ( .A1(n13300), .A2(sram_rdata_2[22]), .Y(n767) );
  NAND3X0_HVT U850 ( .A1(n2080), .A2(n495), .A3(n767), .Y(n_src_aox[262]) );
  NAND2X0_HVT U851 ( .A1(n12300), .A2(sram_rdata_2[21]), .Y(n768) );
  NAND3X0_HVT U852 ( .A1(n2090), .A2(n496), .A3(n768), .Y(n_src_aox[261]) );
  NAND2X0_HVT U853 ( .A1(n1053), .A2(sram_rdata_2[20]), .Y(n769) );
  NAND3X0_HVT U854 ( .A1(n2100), .A2(n497), .A3(n769), .Y(n_src_aox[260]) );
  NAND2X0_HVT U855 ( .A1(n12900), .A2(sram_rdata_2[17]), .Y(n7701) );
  NAND3X0_HVT U856 ( .A1(n2110), .A2(n498), .A3(n7701), .Y(n_src_aox[257]) );
  NAND2X0_HVT U857 ( .A1(n13300), .A2(sram_rdata_2[16]), .Y(n771) );
  NAND3X0_HVT U858 ( .A1(n2120), .A2(n499), .A3(n771), .Y(n_src_aox[256]) );
  NAND2X0_HVT U859 ( .A1(n6300), .A2(sram_rdata_0[31]), .Y(n772) );
  NAND3X0_HVT U860 ( .A1(n2130), .A2(n5001), .A3(n772), .Y(n_src_aox[255]) );
  NAND2X0_HVT U861 ( .A1(n12500), .A2(sram_rdata_0[30]), .Y(n773) );
  NAND3X0_HVT U862 ( .A1(n2140), .A2(n501), .A3(n773), .Y(n_src_aox[254]) );
  NAND2X0_HVT U863 ( .A1(n13400), .A2(sram_rdata_0[28]), .Y(n774) );
  NAND3X0_HVT U864 ( .A1(n2150), .A2(n502), .A3(n774), .Y(n_src_aox[252]) );
  NAND2X0_HVT U865 ( .A1(n10501), .A2(sram_rdata_0[27]), .Y(n775) );
  NAND3X0_HVT U866 ( .A1(n2160), .A2(n503), .A3(n775), .Y(n_src_aox[251]) );
  NAND2X0_HVT U867 ( .A1(n6200), .A2(sram_rdata_0[26]), .Y(n778) );
  NAND3X0_HVT U868 ( .A1(n2170), .A2(n504), .A3(n778), .Y(n_src_aox[250]) );
  NAND2X0_HVT U869 ( .A1(n12700), .A2(sram_rdata_0[25]), .Y(n779) );
  NAND3X0_HVT U870 ( .A1(n2180), .A2(n505), .A3(n779), .Y(n_src_aox[249]) );
  NAND2X0_HVT U871 ( .A1(n10501), .A2(sram_rdata_0[24]), .Y(n7801) );
  NAND3X0_HVT U872 ( .A1(n2190), .A2(n506), .A3(n7801), .Y(n_src_aox[248]) );
  NAND2X0_HVT U873 ( .A1(n10501), .A2(sram_rdata_0[23]), .Y(n781) );
  NAND3X0_HVT U874 ( .A1(n2200), .A2(n507), .A3(n781), .Y(n_src_aox[247]) );
  NAND2X0_HVT U875 ( .A1(n1053), .A2(sram_rdata_0[22]), .Y(n782) );
  NAND3X0_HVT U876 ( .A1(n2210), .A2(n508), .A3(n782), .Y(n_src_aox[246]) );
  NAND2X0_HVT U877 ( .A1(n1051), .A2(sram_rdata_0[21]), .Y(n783) );
  NAND3X0_HVT U878 ( .A1(n2220), .A2(n509), .A3(n783), .Y(n_src_aox[245]) );
  NAND2X0_HVT U879 ( .A1(n12600), .A2(sram_rdata_0[20]), .Y(n784) );
  NAND3X0_HVT U880 ( .A1(n2230), .A2(n5101), .A3(n784), .Y(n_src_aox[244]) );
  NAND2X0_HVT U881 ( .A1(n13100), .A2(sram_rdata_0[19]), .Y(n785) );
  NAND3X0_HVT U882 ( .A1(n2240), .A2(n511), .A3(n785), .Y(n_src_aox[243]) );
  NAND2X0_HVT U883 ( .A1(n13400), .A2(sram_rdata_0[18]), .Y(n786) );
  NAND3X0_HVT U884 ( .A1(n2250), .A2(n512), .A3(n786), .Y(n_src_aox[242]) );
  NAND2X0_HVT U885 ( .A1(n12800), .A2(sram_rdata_0[17]), .Y(n787) );
  NAND3X0_HVT U886 ( .A1(n2260), .A2(n513), .A3(n787), .Y(n_src_aox[241]) );
  NAND2X0_HVT U887 ( .A1(n13200), .A2(sram_rdata_0[16]), .Y(n788) );
  NAND3X0_HVT U888 ( .A1(n2270), .A2(n514), .A3(n788), .Y(n_src_aox[240]) );
  NAND2X0_HVT U889 ( .A1(n12900), .A2(sram_rdata_1[15]), .Y(n789) );
  NAND3X0_HVT U890 ( .A1(n2280), .A2(n515), .A3(n789), .Y(n_src_aox[239]) );
  NAND2X0_HVT U891 ( .A1(n13300), .A2(sram_rdata_1[14]), .Y(n7901) );
  NAND3X0_HVT U892 ( .A1(n2290), .A2(n516), .A3(n7901), .Y(n_src_aox[238]) );
  NAND2X0_HVT U893 ( .A1(n12200), .A2(sram_rdata_1[13]), .Y(n791) );
  NAND3X0_HVT U894 ( .A1(n2300), .A2(n517), .A3(n791), .Y(n_src_aox[237]) );
  NAND2X0_HVT U895 ( .A1(n1052), .A2(sram_rdata_1[12]), .Y(n792) );
  NAND3X0_HVT U896 ( .A1(n2310), .A2(n518), .A3(n792), .Y(n_src_aox[236]) );
  NAND2X0_HVT U897 ( .A1(n6000), .A2(sram_rdata_1[11]), .Y(n793) );
  NAND3X0_HVT U898 ( .A1(n2320), .A2(n519), .A3(n793), .Y(n_src_aox[235]) );
  NAND2X0_HVT U899 ( .A1(n6200), .A2(sram_rdata_1[10]), .Y(n794) );
  NAND3X0_HVT U900 ( .A1(n2330), .A2(n5201), .A3(n794), .Y(n_src_aox[234]) );
  NAND2X0_HVT U901 ( .A1(n6000), .A2(sram_rdata_1[9]), .Y(n795) );
  NAND3X0_HVT U902 ( .A1(n2340), .A2(n521), .A3(n795), .Y(n_src_aox[233]) );
  NAND2X0_HVT U903 ( .A1(n1052), .A2(sram_rdata_1[8]), .Y(n796) );
  NAND3X0_HVT U904 ( .A1(n2350), .A2(n522), .A3(n796), .Y(n_src_aox[232]) );
  NAND2X0_HVT U905 ( .A1(n6000), .A2(sram_rdata_1[7]), .Y(n797) );
  NAND3X0_HVT U906 ( .A1(n2360), .A2(n523), .A3(n797), .Y(n_src_aox[231]) );
  NAND2X0_HVT U907 ( .A1(n6200), .A2(sram_rdata_1[6]), .Y(n798) );
  NAND3X0_HVT U908 ( .A1(n2370), .A2(n524), .A3(n798), .Y(n_src_aox[230]) );
  NAND2X0_HVT U909 ( .A1(n13000), .A2(sram_rdata_1[5]), .Y(n799) );
  NAND3X0_HVT U910 ( .A1(n2380), .A2(n525), .A3(n799), .Y(n_src_aox[229]) );
  NAND2X0_HVT U911 ( .A1(n13400), .A2(sram_rdata_1[4]), .Y(n8001) );
  NAND3X0_HVT U912 ( .A1(n2390), .A2(n526), .A3(n8001), .Y(n_src_aox[228]) );
  NAND2X0_HVT U913 ( .A1(n6000), .A2(sram_rdata_1[3]), .Y(n801) );
  NAND3X0_HVT U914 ( .A1(n2400), .A2(n527), .A3(n801), .Y(n_src_aox[227]) );
  NAND2X0_HVT U915 ( .A1(n12500), .A2(sram_rdata_1[2]), .Y(n802) );
  NAND3X0_HVT U916 ( .A1(n2410), .A2(n528), .A3(n802), .Y(n_src_aox[226]) );
  NAND2X0_HVT U917 ( .A1(n1052), .A2(sram_rdata_1[1]), .Y(n803) );
  NAND3X0_HVT U918 ( .A1(n2420), .A2(n529), .A3(n803), .Y(n_src_aox[225]) );
  NAND2X0_HVT U919 ( .A1(sram_rdata_1[0]), .A2(n12800), .Y(n804) );
  NAND3X0_HVT U920 ( .A1(n2430), .A2(n462), .A3(n804), .Y(n_src_aox[224]) );
  NAND2X0_HVT U921 ( .A1(n6300), .A2(sram_rdata_2[15]), .Y(n805) );
  NAND3X0_HVT U922 ( .A1(n2440), .A2(n5301), .A3(n805), .Y(n_src_aox[223]) );
  NAND2X0_HVT U923 ( .A1(n6300), .A2(sram_rdata_2[14]), .Y(n806) );
  NAND3X0_HVT U924 ( .A1(n2450), .A2(n531), .A3(n806), .Y(n_src_aox[222]) );
  NAND2X0_HVT U925 ( .A1(n1051), .A2(sram_rdata_2[13]), .Y(n807) );
  NAND3X0_HVT U926 ( .A1(n2460), .A2(n532), .A3(n807), .Y(n_src_aox[221]) );
  NAND2X0_HVT U927 ( .A1(n12700), .A2(sram_rdata_2[12]), .Y(n808) );
  NAND3X0_HVT U928 ( .A1(n2470), .A2(n533), .A3(n808), .Y(n_src_aox[220]) );
  NAND2X0_HVT U929 ( .A1(n13100), .A2(sram_rdata_2[11]), .Y(n809) );
  NAND3X0_HVT U930 ( .A1(n2480), .A2(n534), .A3(n809), .Y(n_src_aox[219]) );
  NAND2X0_HVT U931 ( .A1(n12600), .A2(sram_rdata_2[10]), .Y(n8101) );
  NAND3X0_HVT U932 ( .A1(n2490), .A2(n535), .A3(n8101), .Y(n_src_aox[218]) );
  NAND2X0_HVT U933 ( .A1(n12900), .A2(sram_rdata_2[9]), .Y(n811) );
  NAND3X0_HVT U934 ( .A1(n2500), .A2(n536), .A3(n811), .Y(n_src_aox[217]) );
  NAND2X0_HVT U935 ( .A1(n12800), .A2(sram_rdata_2[8]), .Y(n812) );
  NAND3X0_HVT U936 ( .A1(n2510), .A2(n537), .A3(n812), .Y(n_src_aox[216]) );
  NAND2X0_HVT U937 ( .A1(n13200), .A2(sram_rdata_2[7]), .Y(n813) );
  NAND3X0_HVT U938 ( .A1(n2520), .A2(n538), .A3(n813), .Y(n_src_aox[215]) );
  NAND2X0_HVT U939 ( .A1(n1052), .A2(sram_rdata_2[6]), .Y(n814) );
  NAND3X0_HVT U940 ( .A1(n2530), .A2(n539), .A3(n814), .Y(n_src_aox[214]) );
  NAND2X0_HVT U941 ( .A1(n1052), .A2(sram_rdata_2[5]), .Y(n815) );
  NAND3X0_HVT U942 ( .A1(n2540), .A2(n5401), .A3(n815), .Y(n_src_aox[213]) );
  NAND2X0_HVT U943 ( .A1(n12900), .A2(sram_rdata_2[4]), .Y(n816) );
  NAND3X0_HVT U944 ( .A1(n2550), .A2(n541), .A3(n816), .Y(n_src_aox[212]) );
  NAND2X0_HVT U945 ( .A1(n6100), .A2(sram_rdata_2[3]), .Y(n817) );
  NAND3X0_HVT U946 ( .A1(n2560), .A2(n542), .A3(n817), .Y(n_src_aox[211]) );
  NAND2X0_HVT U947 ( .A1(n6100), .A2(sram_rdata_2[2]), .Y(n818) );
  NAND3X0_HVT U948 ( .A1(n2570), .A2(n543), .A3(n818), .Y(n_src_aox[210]) );
  NAND2X0_HVT U949 ( .A1(n6100), .A2(sram_rdata_2[1]), .Y(n819) );
  NAND3X0_HVT U950 ( .A1(n2580), .A2(n544), .A3(n819), .Y(n_src_aox[209]) );
  NAND2X0_HVT U951 ( .A1(sram_rdata_2[0]), .A2(n13200), .Y(n8201) );
  NAND3X0_HVT U952 ( .A1(n2590), .A2(n463), .A3(n8201), .Y(n_src_aox[208]) );
  NAND2X0_HVT U953 ( .A1(n6300), .A2(sram_rdata_0[15]), .Y(n821) );
  NAND3X0_HVT U954 ( .A1(n2600), .A2(n545), .A3(n821), .Y(n_src_aox[207]) );
  NAND2X0_HVT U955 ( .A1(n13300), .A2(sram_rdata_0[14]), .Y(n822) );
  NAND3X0_HVT U956 ( .A1(n2610), .A2(n546), .A3(n822), .Y(n_src_aox[206]) );
  NAND2X0_HVT U957 ( .A1(n13300), .A2(sram_rdata_0[13]), .Y(n823) );
  NAND3X0_HVT U958 ( .A1(n2620), .A2(n547), .A3(n823), .Y(n_src_aox[205]) );
  NAND2X0_HVT U959 ( .A1(n12500), .A2(sram_rdata_0[12]), .Y(n824) );
  NAND3X0_HVT U960 ( .A1(n2630), .A2(n548), .A3(n824), .Y(n_src_aox[204]) );
  NAND2X0_HVT U961 ( .A1(n13000), .A2(sram_rdata_0[11]), .Y(n825) );
  NAND3X0_HVT U962 ( .A1(n2640), .A2(n549), .A3(n825), .Y(n_src_aox[203]) );
  NAND2X0_HVT U963 ( .A1(n13400), .A2(sram_rdata_0[10]), .Y(n826) );
  NAND3X0_HVT U964 ( .A1(n2650), .A2(n5501), .A3(n826), .Y(n_src_aox[202]) );
  NAND2X0_HVT U965 ( .A1(n12700), .A2(sram_rdata_0[9]), .Y(n827) );
  NAND3X0_HVT U966 ( .A1(n2660), .A2(n551), .A3(n827), .Y(n_src_aox[201]) );
  NAND2X0_HVT U967 ( .A1(n13100), .A2(sram_rdata_0[8]), .Y(n828) );
  NAND3X0_HVT U968 ( .A1(n2670), .A2(n552), .A3(n828), .Y(n_src_aox[200]) );
  NAND2X0_HVT U969 ( .A1(n1049), .A2(sram_rdata_0[7]), .Y(n829) );
  NAND3X0_HVT U970 ( .A1(n2680), .A2(n553), .A3(n829), .Y(n_src_aox[199]) );
  NAND2X0_HVT U971 ( .A1(n12300), .A2(sram_rdata_0[6]), .Y(n8301) );
  NAND3X0_HVT U972 ( .A1(n2690), .A2(n554), .A3(n8301), .Y(n_src_aox[198]) );
  NAND2X0_HVT U973 ( .A1(n1053), .A2(sram_rdata_0[5]), .Y(n831) );
  NAND3X0_HVT U974 ( .A1(n2700), .A2(n555), .A3(n831), .Y(n_src_aox[197]) );
  NAND2X0_HVT U975 ( .A1(n6100), .A2(sram_rdata_0[4]), .Y(n832) );
  NAND3X0_HVT U976 ( .A1(n2710), .A2(n556), .A3(n832), .Y(n_src_aox[196]) );
  NAND2X0_HVT U977 ( .A1(n6200), .A2(sram_rdata_0[3]), .Y(n833) );
  NAND3X0_HVT U978 ( .A1(n2720), .A2(n557), .A3(n833), .Y(n_src_aox[195]) );
  NAND2X0_HVT U979 ( .A1(n12300), .A2(sram_rdata_0[2]), .Y(n834) );
  NAND3X0_HVT U980 ( .A1(n2730), .A2(n558), .A3(n834), .Y(n_src_aox[194]) );
  NAND2X0_HVT U981 ( .A1(n6200), .A2(sram_rdata_0[1]), .Y(n835) );
  NAND3X0_HVT U982 ( .A1(n2740), .A2(n559), .A3(n835), .Y(n_src_aox[193]) );
  NAND2X0_HVT U983 ( .A1(sram_rdata_0[0]), .A2(n12600), .Y(n836) );
  NAND3X0_HVT U984 ( .A1(n2750), .A2(n464), .A3(n836), .Y(n_src_aox[192]) );
  NAND2X0_HVT U985 ( .A1(n12600), .A2(sram_rdata_4[31]), .Y(n837) );
  NAND3X0_HVT U986 ( .A1(n2760), .A2(n5601), .A3(n837), .Y(n_src_aox[191]) );
  NAND2X0_HVT U987 ( .A1(n12800), .A2(sram_rdata_4[30]), .Y(n838) );
  NAND3X0_HVT U988 ( .A1(n2770), .A2(n561), .A3(n838), .Y(n_src_aox[190]) );
  NAND2X0_HVT U989 ( .A1(n13200), .A2(sram_rdata_4[29]), .Y(n839) );
  NAND3X0_HVT U990 ( .A1(n2780), .A2(n562), .A3(n839), .Y(n_src_aox[189]) );
  NAND2X0_HVT U991 ( .A1(n1053), .A2(sram_rdata_4[28]), .Y(n8401) );
  NAND3X0_HVT U992 ( .A1(n2790), .A2(n563), .A3(n8401), .Y(n_src_aox[188]) );
  NAND2X0_HVT U993 ( .A1(n13000), .A2(sram_rdata_4[27]), .Y(n841) );
  NAND3X0_HVT U994 ( .A1(n2800), .A2(n564), .A3(n841), .Y(n_src_aox[187]) );
  NAND2X0_HVT U995 ( .A1(n6100), .A2(sram_rdata_4[26]), .Y(n842) );
  NAND3X0_HVT U996 ( .A1(n2810), .A2(n565), .A3(n842), .Y(n_src_aox[186]) );
  NAND2X0_HVT U997 ( .A1(n1053), .A2(sram_rdata_4[25]), .Y(n843) );
  NAND3X0_HVT U998 ( .A1(n2820), .A2(n566), .A3(n843), .Y(n_src_aox[185]) );
  NAND2X0_HVT U999 ( .A1(n1053), .A2(sram_rdata_4[24]), .Y(n844) );
  NAND3X0_HVT U1000 ( .A1(n2830), .A2(n567), .A3(n844), .Y(n_src_aox[184]) );
  NAND2X0_HVT U1001 ( .A1(n12300), .A2(sram_rdata_4[23]), .Y(n845) );
  NAND3X0_HVT U1002 ( .A1(n2840), .A2(n568), .A3(n845), .Y(n_src_aox[183]) );
  NAND2X0_HVT U1003 ( .A1(n12900), .A2(sram_rdata_4[22]), .Y(n846) );
  NAND3X0_HVT U1004 ( .A1(n2850), .A2(n569), .A3(n846), .Y(n_src_aox[182]) );
  NAND2X0_HVT U1005 ( .A1(n13300), .A2(sram_rdata_4[21]), .Y(n847) );
  NAND3X0_HVT U1006 ( .A1(n2860), .A2(n5701), .A3(n847), .Y(n_src_aox[181]) );
  NAND2X0_HVT U1007 ( .A1(n13400), .A2(sram_rdata_4[20]), .Y(n848) );
  NAND3X0_HVT U1008 ( .A1(n2870), .A2(n571), .A3(n848), .Y(n_src_aox[180]) );
  NAND2X0_HVT U1009 ( .A1(n12500), .A2(sram_rdata_4[19]), .Y(n849) );
  NAND3X0_HVT U1010 ( .A1(n2880), .A2(n572), .A3(n849), .Y(n_src_aox[179]) );
  NAND2X0_HVT U1011 ( .A1(n13000), .A2(sram_rdata_4[18]), .Y(n8501) );
  NAND3X0_HVT U1012 ( .A1(n2890), .A2(n573), .A3(n8501), .Y(n_src_aox[178]) );
  NAND2X0_HVT U1013 ( .A1(n13400), .A2(sram_rdata_4[17]), .Y(n851) );
  NAND3X0_HVT U1014 ( .A1(n2900), .A2(n574), .A3(n851), .Y(n_src_aox[177]) );
  NAND2X0_HVT U1015 ( .A1(n6000), .A2(sram_rdata_4[16]), .Y(n852) );
  NAND3X0_HVT U1016 ( .A1(n2910), .A2(n575), .A3(n852), .Y(n_src_aox[176]) );
  NAND2X0_HVT U1017 ( .A1(n1051), .A2(sram_rdata_5[31]), .Y(n853) );
  NAND3X0_HVT U1018 ( .A1(n2920), .A2(n576), .A3(n853), .Y(n_src_aox[175]) );
  NAND2X0_HVT U1019 ( .A1(n12700), .A2(sram_rdata_5[30]), .Y(n854) );
  NAND3X0_HVT U1020 ( .A1(n2930), .A2(n577), .A3(n854), .Y(n_src_aox[174]) );
  NAND2X0_HVT U1021 ( .A1(n12300), .A2(sram_rdata_5[29]), .Y(n855) );
  NAND3X0_HVT U1022 ( .A1(n2940), .A2(n578), .A3(n855), .Y(n_src_aox[173]) );
  NAND2X0_HVT U1023 ( .A1(n1051), .A2(sram_rdata_5[28]), .Y(n856) );
  NAND3X0_HVT U1024 ( .A1(n2950), .A2(n579), .A3(n856), .Y(n_src_aox[172]) );
  NAND2X0_HVT U1025 ( .A1(n6200), .A2(sram_rdata_5[27]), .Y(n857) );
  NAND3X0_HVT U1026 ( .A1(n2960), .A2(n5801), .A3(n857), .Y(n_src_aox[171]) );
  NAND2X0_HVT U1027 ( .A1(n1051), .A2(sram_rdata_5[26]), .Y(n858) );
  NAND3X0_HVT U1028 ( .A1(n2970), .A2(n581), .A3(n858), .Y(n_src_aox[170]) );
  NAND2X0_HVT U1029 ( .A1(n12600), .A2(sram_rdata_5[25]), .Y(n859) );
  NAND3X0_HVT U1030 ( .A1(n2980), .A2(n582), .A3(n859), .Y(n_src_aox[169]) );
  NAND2X0_HVT U1031 ( .A1(n13100), .A2(sram_rdata_5[24]), .Y(n8601) );
  NAND3X0_HVT U1032 ( .A1(n2990), .A2(n583), .A3(n8601), .Y(n_src_aox[168]) );
  NAND2X0_HVT U1033 ( .A1(n12500), .A2(sram_rdata_5[23]), .Y(n861) );
  NAND3X0_HVT U1034 ( .A1(n3000), .A2(n584), .A3(n861), .Y(n_src_aox[167]) );
  NAND2X0_HVT U1035 ( .A1(n12800), .A2(sram_rdata_5[22]), .Y(n862) );
  NAND3X0_HVT U1036 ( .A1(n3010), .A2(n585), .A3(n862), .Y(n_src_aox[166]) );
  NAND2X0_HVT U1037 ( .A1(n13200), .A2(sram_rdata_5[21]), .Y(n863) );
  NAND3X0_HVT U1038 ( .A1(n3020), .A2(n586), .A3(n863), .Y(n_src_aox[165]) );
  NAND2X0_HVT U1039 ( .A1(n12900), .A2(sram_rdata_5[20]), .Y(n864) );
  NAND3X0_HVT U1040 ( .A1(n3030), .A2(n587), .A3(n864), .Y(n_src_aox[164]) );
  NAND2X0_HVT U1041 ( .A1(n13300), .A2(sram_rdata_5[19]), .Y(n865) );
  NAND3X0_HVT U1042 ( .A1(n3040), .A2(n588), .A3(n865), .Y(n_src_aox[163]) );
  NAND2X0_HVT U1043 ( .A1(n1049), .A2(sram_rdata_5[18]), .Y(n866) );
  NAND3X0_HVT U1044 ( .A1(n3050), .A2(n589), .A3(n866), .Y(n_src_aox[162]) );
  NAND2X0_HVT U1045 ( .A1(n6300), .A2(sram_rdata_5[17]), .Y(n867) );
  NAND3X0_HVT U1046 ( .A1(n3060), .A2(n5901), .A3(n867), .Y(n_src_aox[161]) );
  NAND2X0_HVT U1047 ( .A1(n1051), .A2(sram_rdata_5[16]), .Y(n868) );
  NAND3X0_HVT U1048 ( .A1(n3070), .A2(n591), .A3(n868), .Y(n_src_aox[160]) );
  NAND2X0_HVT U1049 ( .A1(n1051), .A2(sram_rdata_3[31]), .Y(n869) );
  NAND3X0_HVT U1050 ( .A1(n3080), .A2(n592), .A3(n869), .Y(n_src_aox[159]) );
  NAND2X0_HVT U1051 ( .A1(n1051), .A2(sram_rdata_3[30]), .Y(n8701) );
  NAND3X0_HVT U1052 ( .A1(n3090), .A2(n593), .A3(n8701), .Y(n_src_aox[158]) );
  NAND2X0_HVT U1053 ( .A1(n6300), .A2(sram_rdata_3[29]), .Y(n871) );
  NAND3X0_HVT U1054 ( .A1(n3100), .A2(n594), .A3(n871), .Y(n_src_aox[157]) );
  NAND2X0_HVT U1055 ( .A1(n1051), .A2(sram_rdata_3[28]), .Y(n872) );
  NAND3X0_HVT U1056 ( .A1(n3110), .A2(n595), .A3(n872), .Y(n_src_aox[156]) );
  NAND2X0_HVT U1057 ( .A1(n13200), .A2(sram_rdata_3[27]), .Y(n873) );
  NAND3X0_HVT U1058 ( .A1(n3120), .A2(n596), .A3(n873), .Y(n_src_aox[155]) );
  NAND2X0_HVT U1059 ( .A1(n13000), .A2(sram_rdata_3[26]), .Y(n874) );
  NAND3X0_HVT U1060 ( .A1(n3130), .A2(n597), .A3(n874), .Y(n_src_aox[154]) );
  NAND2X0_HVT U1061 ( .A1(n13400), .A2(sram_rdata_3[25]), .Y(n875) );
  NAND3X0_HVT U1062 ( .A1(n3140), .A2(n598), .A3(n875), .Y(n_src_aox[153]) );
  NAND2X0_HVT U1063 ( .A1(n6000), .A2(sram_rdata_3[24]), .Y(n876) );
  NAND3X0_HVT U1064 ( .A1(n3150), .A2(n599), .A3(n876), .Y(n_src_aox[152]) );
  NAND2X0_HVT U1065 ( .A1(n1053), .A2(sram_rdata_3[22]), .Y(n877) );
  NAND3X0_HVT U1066 ( .A1(n3160), .A2(n6001), .A3(n877), .Y(n_src_aox[150]) );
  NAND2X0_HVT U1067 ( .A1(n12300), .A2(sram_rdata_3[21]), .Y(n878) );
  NAND3X0_HVT U1068 ( .A1(n3170), .A2(n601), .A3(n878), .Y(n_src_aox[149]) );
  NAND2X0_HVT U1069 ( .A1(n1053), .A2(sram_rdata_3[20]), .Y(n879) );
  NAND3X0_HVT U1070 ( .A1(n3180), .A2(n602), .A3(n879), .Y(n_src_aox[148]) );
  NAND2X0_HVT U1071 ( .A1(n12200), .A2(sram_rdata_3[19]), .Y(n8801) );
  NAND3X0_HVT U1072 ( .A1(n3190), .A2(n603), .A3(n8801), .Y(n_src_aox[147]) );
  NAND2X0_HVT U1073 ( .A1(n12700), .A2(sram_rdata_3[18]), .Y(n881) );
  NAND3X0_HVT U1074 ( .A1(n3200), .A2(n604), .A3(n881), .Y(n_src_aox[146]) );
  NAND2X0_HVT U1075 ( .A1(n13100), .A2(sram_rdata_3[17]), .Y(n882) );
  NAND3X0_HVT U1076 ( .A1(n3210), .A2(n605), .A3(n882), .Y(n_src_aox[145]) );
  NAND2X0_HVT U1077 ( .A1(n12600), .A2(sram_rdata_3[16]), .Y(n883) );
  NAND3X0_HVT U1078 ( .A1(n3220), .A2(n606), .A3(n883), .Y(n_src_aox[144]) );
  NAND2X0_HVT U1079 ( .A1(n1362), .A2(sram_rdata_4[15]), .Y(n884) );
  NAND3X0_HVT U1080 ( .A1(n3230), .A2(n607), .A3(n884), .Y(n_src_aox[143]) );
  NAND2X0_HVT U1081 ( .A1(n12800), .A2(sram_rdata_4[14]), .Y(n885) );
  NAND3X0_HVT U1082 ( .A1(n3240), .A2(n608), .A3(n885), .Y(n_src_aox[142]) );
  NAND2X0_HVT U1083 ( .A1(n13200), .A2(sram_rdata_4[13]), .Y(n886) );
  NAND3X0_HVT U1084 ( .A1(n3250), .A2(n609), .A3(n886), .Y(n_src_aox[141]) );
  NAND2X0_HVT U1085 ( .A1(n6000), .A2(sram_rdata_4[12]), .Y(n887) );
  NAND3X0_HVT U1086 ( .A1(n3260), .A2(n6101), .A3(n887), .Y(n_src_aox[140]) );
  NAND2X0_HVT U1087 ( .A1(n6100), .A2(sram_rdata_4[11]), .Y(n888) );
  NAND3X0_HVT U1088 ( .A1(n327), .A2(n611), .A3(n888), .Y(n_src_aox[139]) );
  NAND2X0_HVT U1089 ( .A1(n12900), .A2(sram_rdata_4[10]), .Y(n889) );
  NAND3X0_HVT U1090 ( .A1(n328), .A2(n612), .A3(n889), .Y(n_src_aox[138]) );
  NAND2X0_HVT U1091 ( .A1(n1049), .A2(sram_rdata_4[9]), .Y(n8901) );
  NAND3X0_HVT U1092 ( .A1(n329), .A2(n613), .A3(n8901), .Y(n_src_aox[137]) );
  NAND2X0_HVT U1093 ( .A1(n1049), .A2(sram_rdata_4[8]), .Y(n891) );
  NAND3X0_HVT U1094 ( .A1(n330), .A2(n614), .A3(n891), .Y(n_src_aox[136]) );
  NAND2X0_HVT U1095 ( .A1(n1051), .A2(sram_rdata_4[7]), .Y(n892) );
  NAND3X0_HVT U1096 ( .A1(n331), .A2(n615), .A3(n892), .Y(n_src_aox[135]) );
  NAND2X0_HVT U1097 ( .A1(n1051), .A2(sram_rdata_4[6]), .Y(n893) );
  NAND3X0_HVT U1098 ( .A1(n332), .A2(n616), .A3(n893), .Y(n_src_aox[134]) );
  NAND2X0_HVT U1099 ( .A1(n12800), .A2(sram_rdata_4[5]), .Y(n894) );
  NAND3X0_HVT U1100 ( .A1(n333), .A2(n617), .A3(n894), .Y(n_src_aox[133]) );
  NAND2X0_HVT U1101 ( .A1(n13300), .A2(sram_rdata_4[4]), .Y(n895) );
  NAND3X0_HVT U1102 ( .A1(n334), .A2(n618), .A3(n895), .Y(n_src_aox[132]) );
  NAND2X0_HVT U1103 ( .A1(n12500), .A2(sram_rdata_4[3]), .Y(n896) );
  NAND3X0_HVT U1104 ( .A1(n335), .A2(n619), .A3(n896), .Y(n_src_aox[131]) );
  NAND2X0_HVT U1105 ( .A1(n13000), .A2(sram_rdata_4[2]), .Y(n897) );
  NAND3X0_HVT U1106 ( .A1(n336), .A2(n6201), .A3(n897), .Y(n_src_aox[130]) );
  NAND2X0_HVT U1107 ( .A1(n13400), .A2(sram_rdata_4[1]), .Y(n898) );
  NAND3X0_HVT U1108 ( .A1(n337), .A2(n621), .A3(n898), .Y(n_src_aox[129]) );
  NAND2X0_HVT U1109 ( .A1(n12700), .A2(sram_rdata_4[0]), .Y(n899) );
  NAND3X0_HVT U1110 ( .A1(n338), .A2(n465), .A3(n899), .Y(n_src_aox[128]) );
  NAND2X0_HVT U1111 ( .A1(n13100), .A2(sram_rdata_5[15]), .Y(n9001) );
  NAND3X0_HVT U1112 ( .A1(n339), .A2(n622), .A3(n9001), .Y(n_src_aox[127]) );
  NAND2X0_HVT U1113 ( .A1(n6200), .A2(sram_rdata_5[14]), .Y(n901) );
  NAND3X0_HVT U1114 ( .A1(n340), .A2(n623), .A3(n901), .Y(n_src_aox[126]) );
  NAND2X0_HVT U1115 ( .A1(n6100), .A2(sram_rdata_5[13]), .Y(n902) );
  NAND3X0_HVT U1116 ( .A1(n341), .A2(n624), .A3(n902), .Y(n_src_aox[125]) );
  NAND2X0_HVT U1117 ( .A1(n6200), .A2(sram_rdata_5[12]), .Y(n903) );
  NAND3X0_HVT U1118 ( .A1(n342), .A2(n625), .A3(n903), .Y(n_src_aox[124]) );
  NAND2X0_HVT U1119 ( .A1(n12200), .A2(sram_rdata_5[11]), .Y(n904) );
  NAND3X0_HVT U1120 ( .A1(n343), .A2(n626), .A3(n904), .Y(n_src_aox[123]) );
  NAND2X0_HVT U1121 ( .A1(n6100), .A2(sram_rdata_5[9]), .Y(n905) );
  NAND3X0_HVT U1122 ( .A1(n344), .A2(n627), .A3(n905), .Y(n_src_aox[121]) );
  NAND2X0_HVT U1123 ( .A1(n1052), .A2(sram_rdata_5[8]), .Y(n906) );
  NAND3X0_HVT U1124 ( .A1(n345), .A2(n628), .A3(n906), .Y(n_src_aox[120]) );
  NAND2X0_HVT U1125 ( .A1(n12600), .A2(sram_rdata_5[7]), .Y(n907) );
  NAND3X0_HVT U1126 ( .A1(n3460), .A2(n629), .A3(n907), .Y(n_src_aox[119]) );
  NAND2X0_HVT U1127 ( .A1(n12800), .A2(sram_rdata_5[6]), .Y(n908) );
  NAND3X0_HVT U1128 ( .A1(n347), .A2(n6301), .A3(n908), .Y(n_src_aox[118]) );
  NAND2X0_HVT U1129 ( .A1(n13200), .A2(sram_rdata_5[5]), .Y(n909) );
  NAND3X0_HVT U1130 ( .A1(n348), .A2(n631), .A3(n909), .Y(n_src_aox[117]) );
  NAND2X0_HVT U1131 ( .A1(n1052), .A2(sram_rdata_5[4]), .Y(n9101) );
  NAND3X0_HVT U1132 ( .A1(n349), .A2(n632), .A3(n9101), .Y(n_src_aox[116]) );
  NAND2X0_HVT U1133 ( .A1(n12600), .A2(sram_rdata_5[3]), .Y(n911) );
  NAND3X0_HVT U1134 ( .A1(n350), .A2(n633), .A3(n911), .Y(n_src_aox[115]) );
  NAND2X0_HVT U1135 ( .A1(n12300), .A2(sram_rdata_5[2]), .Y(n912) );
  NAND3X0_HVT U1136 ( .A1(n351), .A2(n634), .A3(n912), .Y(n_src_aox[114]) );
  NAND2X0_HVT U1137 ( .A1(n6100), .A2(sram_rdata_5[1]), .Y(n913) );
  NAND3X0_HVT U1138 ( .A1(n352), .A2(n635), .A3(n913), .Y(n_src_aox[113]) );
  NAND2X0_HVT U1139 ( .A1(n6000), .A2(sram_rdata_5[0]), .Y(n914) );
  NAND3X0_HVT U1140 ( .A1(n353), .A2(n466), .A3(n914), .Y(n_src_aox[112]) );
  NAND2X0_HVT U1141 ( .A1(n12200), .A2(sram_rdata_3[15]), .Y(n915) );
  NAND3X0_HVT U1142 ( .A1(n354), .A2(n636), .A3(n915), .Y(n_src_aox[111]) );
  NAND2X0_HVT U1143 ( .A1(n12900), .A2(sram_rdata_3[14]), .Y(n916) );
  NAND3X0_HVT U1144 ( .A1(n355), .A2(n637), .A3(n916), .Y(n_src_aox[110]) );
  NAND2X0_HVT U1145 ( .A1(n13300), .A2(sram_rdata_3[13]), .Y(n917) );
  NAND3X0_HVT U1146 ( .A1(n356), .A2(n638), .A3(n917), .Y(n_src_aox[109]) );
  NAND2X0_HVT U1147 ( .A1(n12900), .A2(sram_rdata_3[12]), .Y(n918) );
  NAND3X0_HVT U1148 ( .A1(n357), .A2(n639), .A3(n918), .Y(n_src_aox[108]) );
  NAND2X0_HVT U1149 ( .A1(n12500), .A2(sram_rdata_3[11]), .Y(n919) );
  NAND3X0_HVT U1150 ( .A1(n358), .A2(n6401), .A3(n919), .Y(n_src_aox[107]) );
  NAND2X0_HVT U1151 ( .A1(n13000), .A2(sram_rdata_3[10]), .Y(n9201) );
  NAND3X0_HVT U1152 ( .A1(n359), .A2(n641), .A3(n9201), .Y(n_src_aox[106]) );
  NAND2X0_HVT U1153 ( .A1(n13400), .A2(sram_rdata_3[9]), .Y(n921) );
  NAND3X0_HVT U1154 ( .A1(n360), .A2(n642), .A3(n921), .Y(n_src_aox[105]) );
  NAND2X0_HVT U1155 ( .A1(n10501), .A2(sram_rdata_3[8]), .Y(n922) );
  NAND3X0_HVT U1156 ( .A1(n361), .A2(n643), .A3(n922), .Y(n_src_aox[104]) );
  NAND2X0_HVT U1157 ( .A1(n10501), .A2(sram_rdata_3[7]), .Y(n923) );
  NAND3X0_HVT U1158 ( .A1(n362), .A2(n644), .A3(n923), .Y(n_src_aox[103]) );
  NAND2X0_HVT U1159 ( .A1(n12700), .A2(sram_rdata_3[6]), .Y(n924) );
  NAND3X0_HVT U1160 ( .A1(n363), .A2(n645), .A3(n924), .Y(n_src_aox[102]) );
  NAND2X0_HVT U1161 ( .A1(n6300), .A2(sram_rdata_3[5]), .Y(n925) );
  NAND3X0_HVT U1162 ( .A1(n364), .A2(n646), .A3(n925), .Y(n_src_aox[101]) );
  NAND2X0_HVT U1163 ( .A1(n6300), .A2(sram_rdata_3[4]), .Y(n926) );
  NAND3X0_HVT U1164 ( .A1(n365), .A2(n647), .A3(n926), .Y(n_src_aox[100]) );
  NAND2X0_HVT U1165 ( .A1(n6100), .A2(sram_rdata_3[3]), .Y(n927) );
  NAND3X0_HVT U1166 ( .A1(n366), .A2(n648), .A3(n927), .Y(n_src_aox[99]) );
  NAND2X0_HVT U1167 ( .A1(n6100), .A2(sram_rdata_3[2]), .Y(n928) );
  NAND3X0_HVT U1168 ( .A1(n367), .A2(n649), .A3(n928), .Y(n_src_aox[98]) );
  NAND2X0_HVT U1169 ( .A1(n12600), .A2(sram_rdata_3[1]), .Y(n929) );
  NAND3X0_HVT U1170 ( .A1(n368), .A2(n6501), .A3(n929), .Y(n_src_aox[97]) );
  NAND2X0_HVT U1171 ( .A1(n13100), .A2(sram_rdata_3[0]), .Y(n9301) );
  NAND3X0_HVT U1172 ( .A1(n369), .A2(n467), .A3(n9301), .Y(n_src_aox[96]) );
  NAND2X0_HVT U1173 ( .A1(n13200), .A2(sram_rdata_7[31]), .Y(n931) );
  NAND3X0_HVT U1174 ( .A1(n370), .A2(n651), .A3(n931), .Y(n_src_aox[95]) );
  NAND2X0_HVT U1175 ( .A1(n12800), .A2(sram_rdata_7[30]), .Y(n932) );
  NAND3X0_HVT U1176 ( .A1(n371), .A2(n652), .A3(n932), .Y(n_src_aox[94]) );
  NAND2X0_HVT U1177 ( .A1(n13200), .A2(sram_rdata_7[29]), .Y(n933) );
  NAND3X0_HVT U1178 ( .A1(n372), .A2(n653), .A3(n933), .Y(n_src_aox[93]) );
  NAND2X0_HVT U1179 ( .A1(n12900), .A2(sram_rdata_7[28]), .Y(n934) );
  NAND3X0_HVT U1180 ( .A1(n373), .A2(n654), .A3(n934), .Y(n_src_aox[92]) );
  NAND2X0_HVT U1181 ( .A1(n13300), .A2(sram_rdata_7[27]), .Y(n935) );
  NAND3X0_HVT U1182 ( .A1(n374), .A2(n655), .A3(n935), .Y(n_src_aox[91]) );
  NAND2X0_HVT U1183 ( .A1(n6000), .A2(sram_rdata_7[26]), .Y(n936) );
  NAND3X0_HVT U1184 ( .A1(n375), .A2(n656), .A3(n936), .Y(n_src_aox[90]) );
  NAND2X0_HVT U1185 ( .A1(n10501), .A2(sram_rdata_7[25]), .Y(n937) );
  NAND3X0_HVT U1186 ( .A1(n376), .A2(n657), .A3(n937), .Y(n_src_aox[89]) );
  NAND2X0_HVT U1187 ( .A1(n6000), .A2(sram_rdata_7[24]), .Y(n938) );
  NAND3X0_HVT U1188 ( .A1(n377), .A2(n658), .A3(n938), .Y(n_src_aox[88]) );
  NAND2X0_HVT U1189 ( .A1(n12200), .A2(sram_rdata_7[23]), .Y(n939) );
  NAND3X0_HVT U1190 ( .A1(n378), .A2(n659), .A3(n939), .Y(n_src_aox[87]) );
  NAND2X0_HVT U1191 ( .A1(n10501), .A2(sram_rdata_7[21]), .Y(n9401) );
  NAND3X0_HVT U1192 ( .A1(n379), .A2(n6601), .A3(n9401), .Y(n_src_aox[85]) );
  NAND2X0_HVT U1193 ( .A1(n12300), .A2(sram_rdata_7[20]), .Y(n941) );
  NAND3X0_HVT U1194 ( .A1(n380), .A2(n661), .A3(n941), .Y(n_src_aox[84]) );
  NAND2X0_HVT U1195 ( .A1(n13000), .A2(sram_rdata_7[19]), .Y(n942) );
  NAND3X0_HVT U1196 ( .A1(n381), .A2(n662), .A3(n942), .Y(n_src_aox[83]) );
  NAND2X0_HVT U1197 ( .A1(n13000), .A2(sram_rdata_7[18]), .Y(n943) );
  NAND3X0_HVT U1198 ( .A1(n382), .A2(n663), .A3(n943), .Y(n_src_aox[82]) );
  NAND2X0_HVT U1199 ( .A1(n13400), .A2(sram_rdata_7[17]), .Y(n944) );
  NAND3X0_HVT U1200 ( .A1(n383), .A2(n664), .A3(n944), .Y(n_src_aox[81]) );
  NAND2X0_HVT U1201 ( .A1(n1053), .A2(sram_rdata_7[16]), .Y(n945) );
  NAND3X0_HVT U1202 ( .A1(n384), .A2(n665), .A3(n945), .Y(n_src_aox[80]) );
  NAND2X0_HVT U1203 ( .A1(n12500), .A2(sram_rdata_8[31]), .Y(n946) );
  NAND3X0_HVT U1204 ( .A1(n385), .A2(n666), .A3(n946), .Y(n_src_aox[79]) );
  NAND2X0_HVT U1205 ( .A1(n6000), .A2(sram_rdata_8[30]), .Y(n947) );
  NAND3X0_HVT U1206 ( .A1(n386), .A2(n667), .A3(n947), .Y(n_src_aox[78]) );
  NAND2X0_HVT U1207 ( .A1(n10501), .A2(sram_rdata_8[29]), .Y(n948) );
  NAND3X0_HVT U1208 ( .A1(n387), .A2(n668), .A3(n948), .Y(n_src_aox[77]) );
  NAND2X0_HVT U1209 ( .A1(n6100), .A2(sram_rdata_8[28]), .Y(n949) );
  NAND3X0_HVT U1210 ( .A1(n388), .A2(n669), .A3(n949), .Y(n_src_aox[76]) );
  NAND2X0_HVT U1211 ( .A1(n12200), .A2(sram_rdata_8[27]), .Y(n9501) );
  NAND3X0_HVT U1212 ( .A1(n389), .A2(n6701), .A3(n9501), .Y(n_src_aox[75]) );
  NAND2X0_HVT U1213 ( .A1(n12700), .A2(sram_rdata_8[26]), .Y(n951) );
  NAND3X0_HVT U1214 ( .A1(n3901), .A2(n671), .A3(n951), .Y(n_src_aox[74]) );
  NAND2X0_HVT U1215 ( .A1(n13100), .A2(sram_rdata_8[25]), .Y(n952) );
  NAND3X0_HVT U1216 ( .A1(n391), .A2(n672), .A3(n952), .Y(n_src_aox[73]) );
  NAND2X0_HVT U1217 ( .A1(n12600), .A2(sram_rdata_8[24]), .Y(n953) );
  NAND3X0_HVT U1218 ( .A1(n392), .A2(n673), .A3(n953), .Y(n_src_aox[72]) );
  NAND2X0_HVT U1219 ( .A1(n12800), .A2(sram_rdata_8[23]), .Y(n954) );
  NAND3X0_HVT U1220 ( .A1(n393), .A2(n674), .A3(n954), .Y(n_src_aox[71]) );
  NAND2X0_HVT U1221 ( .A1(n12800), .A2(sram_rdata_8[22]), .Y(n955) );
  NAND3X0_HVT U1222 ( .A1(n394), .A2(n675), .A3(n955), .Y(n_src_aox[70]) );
  NAND2X0_HVT U1223 ( .A1(n13200), .A2(sram_rdata_8[21]), .Y(n956) );
  NAND3X0_HVT U1224 ( .A1(n395), .A2(n676), .A3(n956), .Y(n_src_aox[69]) );
  NAND2X0_HVT U1225 ( .A1(n6200), .A2(sram_rdata_8[20]), .Y(n957) );
  NAND3X0_HVT U1226 ( .A1(n396), .A2(n677), .A3(n957), .Y(n_src_aox[68]) );
  NAND2X0_HVT U1227 ( .A1(n6200), .A2(sram_rdata_8[19]), .Y(n958) );
  NAND3X0_HVT U1228 ( .A1(n397), .A2(n678), .A3(n958), .Y(n_src_aox[67]) );
  NAND2X0_HVT U1229 ( .A1(n12900), .A2(sram_rdata_8[18]), .Y(n959) );
  NAND3X0_HVT U1230 ( .A1(n398), .A2(n679), .A3(n959), .Y(n_src_aox[66]) );
  NAND2X0_HVT U1231 ( .A1(n12300), .A2(sram_rdata_8[17]), .Y(n9601) );
  NAND3X0_HVT U1232 ( .A1(n399), .A2(n6801), .A3(n9601), .Y(n_src_aox[65]) );
  NAND2X0_HVT U1233 ( .A1(n12300), .A2(sram_rdata_8[16]), .Y(n961) );
  NAND3X0_HVT U1234 ( .A1(n4001), .A2(n681), .A3(n961), .Y(n_src_aox[64]) );
  NAND2X0_HVT U1235 ( .A1(n1051), .A2(sram_rdata_6[31]), .Y(n962) );
  NAND3X0_HVT U1236 ( .A1(n401), .A2(n682), .A3(n962), .Y(n_src_aox[63]) );
  NAND2X0_HVT U1237 ( .A1(n1049), .A2(sram_rdata_6[30]), .Y(n963) );
  NAND3X0_HVT U1238 ( .A1(n402), .A2(n683), .A3(n963), .Y(n_src_aox[62]) );
  NAND2X0_HVT U1239 ( .A1(n6300), .A2(sram_rdata_6[29]), .Y(n964) );
  NAND3X0_HVT U1240 ( .A1(n403), .A2(n684), .A3(n964), .Y(n_src_aox[61]) );
  NAND2X0_HVT U1241 ( .A1(n13300), .A2(sram_rdata_6[28]), .Y(n965) );
  NAND3X0_HVT U1242 ( .A1(n404), .A2(n685), .A3(n965), .Y(n_src_aox[60]) );
  NAND2X0_HVT U1243 ( .A1(n12500), .A2(sram_rdata_6[27]), .Y(n966) );
  NAND3X0_HVT U1244 ( .A1(n405), .A2(n686), .A3(n966), .Y(n_src_aox[59]) );
  NAND2X0_HVT U1245 ( .A1(n13000), .A2(sram_rdata_6[26]), .Y(n967) );
  NAND3X0_HVT U1246 ( .A1(n406), .A2(n687), .A3(n967), .Y(n_src_aox[58]) );
  NAND2X0_HVT U1247 ( .A1(n13400), .A2(sram_rdata_6[25]), .Y(n968) );
  NAND3X0_HVT U1248 ( .A1(n407), .A2(n688), .A3(n968), .Y(n_src_aox[57]) );
  NAND2X0_HVT U1249 ( .A1(n12700), .A2(sram_rdata_6[24]), .Y(n969) );
  NAND3X0_HVT U1250 ( .A1(n408), .A2(n689), .A3(n969), .Y(n_src_aox[56]) );
  NAND2X0_HVT U1251 ( .A1(n13100), .A2(sram_rdata_6[23]), .Y(n9701) );
  NAND3X0_HVT U1252 ( .A1(n409), .A2(n6901), .A3(n9701), .Y(n_src_aox[55]) );
  NAND2X0_HVT U1253 ( .A1(n1052), .A2(sram_rdata_6[22]), .Y(n971) );
  NAND3X0_HVT U1254 ( .A1(n4101), .A2(n691), .A3(n971), .Y(n_src_aox[54]) );
  NAND2X0_HVT U1255 ( .A1(n1053), .A2(sram_rdata_6[21]), .Y(n972) );
  NAND3X0_HVT U1256 ( .A1(n411), .A2(n692), .A3(n972), .Y(n_src_aox[53]) );
  NAND2X0_HVT U1257 ( .A1(n1049), .A2(sram_rdata_6[20]), .Y(n973) );
  NAND3X0_HVT U1258 ( .A1(n412), .A2(n693), .A3(n973), .Y(n_src_aox[52]) );
  NAND2X0_HVT U1259 ( .A1(n12200), .A2(sram_rdata_6[19]), .Y(n974) );
  NAND3X0_HVT U1260 ( .A1(n413), .A2(n694), .A3(n974), .Y(n_src_aox[51]) );
  NAND2X0_HVT U1261 ( .A1(n1052), .A2(sram_rdata_6[18]), .Y(n975) );
  NAND3X0_HVT U1262 ( .A1(n414), .A2(n695), .A3(n975), .Y(n_src_aox[50]) );
  NAND2X0_HVT U1263 ( .A1(n1049), .A2(sram_rdata_6[17]), .Y(n976) );
  NAND3X0_HVT U1264 ( .A1(n415), .A2(n696), .A3(n976), .Y(n_src_aox[49]) );
  NAND2X0_HVT U1265 ( .A1(n12600), .A2(sram_rdata_7[15]), .Y(n977) );
  NAND3X0_HVT U1266 ( .A1(n416), .A2(n697), .A3(n977), .Y(n_src_aox[47]) );
  NAND2X0_HVT U1267 ( .A1(n12800), .A2(sram_rdata_7[14]), .Y(n978) );
  NAND3X0_HVT U1268 ( .A1(n417), .A2(n698), .A3(n978), .Y(n_src_aox[46]) );
  NAND2X0_HVT U1269 ( .A1(n13200), .A2(sram_rdata_7[13]), .Y(n979) );
  NAND3X0_HVT U1270 ( .A1(n418), .A2(n699), .A3(n979), .Y(n_src_aox[45]) );
  NAND2X0_HVT U1271 ( .A1(n6100), .A2(sram_rdata_7[12]), .Y(n9801) );
  NAND3X0_HVT U1272 ( .A1(n419), .A2(n7001), .A3(n9801), .Y(n_src_aox[44]) );
  NAND2X0_HVT U1273 ( .A1(n1362), .A2(sram_rdata_7[11]), .Y(n981) );
  NAND3X0_HVT U1274 ( .A1(n4201), .A2(n701), .A3(n981), .Y(n_src_aox[43]) );
  NAND2X0_HVT U1275 ( .A1(n10501), .A2(sram_rdata_7[10]), .Y(n982) );
  NAND3X0_HVT U1276 ( .A1(n421), .A2(n702), .A3(n982), .Y(n_src_aox[42]) );
  NAND2X0_HVT U1277 ( .A1(n6300), .A2(sram_rdata_7[9]), .Y(n983) );
  NAND3X0_HVT U1278 ( .A1(n422), .A2(n703), .A3(n983), .Y(n_src_aox[41]) );
  NAND2X0_HVT U1279 ( .A1(n6300), .A2(sram_rdata_7[8]), .Y(n984) );
  NAND3X0_HVT U1280 ( .A1(n423), .A2(n704), .A3(n984), .Y(n_src_aox[40]) );
  NAND2X0_HVT U1281 ( .A1(n12200), .A2(sram_rdata_7[7]), .Y(n985) );
  NAND3X0_HVT U1282 ( .A1(n424), .A2(n705), .A3(n985), .Y(n_src_aox[39]) );
  NAND2X0_HVT U1283 ( .A1(n12900), .A2(sram_rdata_7[6]), .Y(n986) );
  NAND3X0_HVT U1284 ( .A1(n425), .A2(n706), .A3(n986), .Y(n_src_aox[38]) );
  NAND2X0_HVT U1285 ( .A1(n13300), .A2(sram_rdata_7[5]), .Y(n987) );
  NAND3X0_HVT U1286 ( .A1(n426), .A2(n707), .A3(n987), .Y(n_src_aox[37]) );
  NAND2X0_HVT U1287 ( .A1(n6200), .A2(sram_rdata_7[4]), .Y(n988) );
  NAND3X0_HVT U1288 ( .A1(n427), .A2(n708), .A3(n988), .Y(n_src_aox[36]) );
  NAND2X0_HVT U1289 ( .A1(n12500), .A2(sram_rdata_7[3]), .Y(n989) );
  NAND3X0_HVT U1290 ( .A1(n428), .A2(n709), .A3(n989), .Y(n_src_aox[35]) );
  NAND2X0_HVT U1291 ( .A1(n13000), .A2(sram_rdata_7[2]), .Y(n9901) );
  NAND3X0_HVT U1292 ( .A1(n429), .A2(n7101), .A3(n9901), .Y(n_src_aox[34]) );
  NAND2X0_HVT U1293 ( .A1(n13400), .A2(sram_rdata_7[1]), .Y(n991) );
  NAND3X0_HVT U1294 ( .A1(n4301), .A2(n711), .A3(n991), .Y(n_src_aox[33]) );
  NAND2X0_HVT U1295 ( .A1(n1049), .A2(sram_rdata_7[0]), .Y(n992) );
  NAND3X0_HVT U1296 ( .A1(n431), .A2(n468), .A3(n992), .Y(n_src_aox[32]) );
  NAND2X0_HVT U1297 ( .A1(n1049), .A2(sram_rdata_8[15]), .Y(n993) );
  NAND3X0_HVT U1298 ( .A1(n432), .A2(n712), .A3(n993), .Y(n_src_aox[31]) );
  NAND2X0_HVT U1299 ( .A1(n12700), .A2(sram_rdata_8[14]), .Y(n994) );
  NAND3X0_HVT U1300 ( .A1(n433), .A2(n713), .A3(n994), .Y(n_src_aox[30]) );
  NAND2X0_HVT U1301 ( .A1(n1053), .A2(sram_rdata_8[13]), .Y(n995) );
  NAND3X0_HVT U1302 ( .A1(n434), .A2(n714), .A3(n995), .Y(n_src_aox[29]) );
  NAND2X0_HVT U1303 ( .A1(n12300), .A2(sram_rdata_8[12]), .Y(n996) );
  NAND3X0_HVT U1304 ( .A1(n435), .A2(n715), .A3(n996), .Y(n_src_aox[28]) );
  NAND2X0_HVT U1305 ( .A1(n6000), .A2(sram_rdata_8[11]), .Y(n997) );
  NAND3X0_HVT U1306 ( .A1(n436), .A2(n716), .A3(n997), .Y(n_src_aox[27]) );
  NAND2X0_HVT U1307 ( .A1(n12300), .A2(sram_rdata_8[10]), .Y(n998) );
  NAND3X0_HVT U1308 ( .A1(n437), .A2(n717), .A3(n998), .Y(n_src_aox[26]) );
  NAND2X0_HVT U1309 ( .A1(n12600), .A2(sram_rdata_8[9]), .Y(n999) );
  NAND3X0_HVT U1310 ( .A1(n438), .A2(n718), .A3(n999), .Y(n_src_aox[25]) );
  NAND2X0_HVT U1311 ( .A1(n13100), .A2(sram_rdata_8[8]), .Y(n10001) );
  NAND3X0_HVT U1312 ( .A1(n439), .A2(n719), .A3(n10001), .Y(n_src_aox[24]) );
  NAND2X0_HVT U1313 ( .A1(n1362), .A2(sram_rdata_8[7]), .Y(n1001) );
  NAND3X0_HVT U1314 ( .A1(n4401), .A2(n7201), .A3(n1001), .Y(n_src_aox[23]) );
  NAND2X0_HVT U1315 ( .A1(n12800), .A2(sram_rdata_8[6]), .Y(n1002) );
  NAND3X0_HVT U1316 ( .A1(n441), .A2(n721), .A3(n1002), .Y(n_src_aox[22]) );
  NAND2X0_HVT U1317 ( .A1(n13200), .A2(sram_rdata_8[5]), .Y(n1003) );
  NAND3X0_HVT U1318 ( .A1(n442), .A2(n722), .A3(n1003), .Y(n_src_aox[21]) );
  NAND2X0_HVT U1319 ( .A1(n12900), .A2(sram_rdata_8[4]), .Y(n1004) );
  NAND3X0_HVT U1320 ( .A1(n443), .A2(n723), .A3(n1004), .Y(n_src_aox[20]) );
  NAND2X0_HVT U1321 ( .A1(n13300), .A2(sram_rdata_8[3]), .Y(n1005) );
  NAND3X0_HVT U1322 ( .A1(n444), .A2(n724), .A3(n1005), .Y(n_src_aox[19]) );
  NAND2X0_HVT U1323 ( .A1(n1052), .A2(sram_rdata_8[2]), .Y(n1006) );
  NAND3X0_HVT U1324 ( .A1(n445), .A2(n725), .A3(n1006), .Y(n_src_aox[18]) );
  NAND2X0_HVT U1325 ( .A1(n1053), .A2(sram_rdata_8[1]), .Y(n1007) );
  NAND3X0_HVT U1326 ( .A1(n446), .A2(n726), .A3(n1007), .Y(n_src_aox[17]) );
  NAND2X0_HVT U1327 ( .A1(n10501), .A2(sram_rdata_8[0]), .Y(n1008) );
  NAND3X0_HVT U1328 ( .A1(n447), .A2(n469), .A3(n1008), .Y(n_src_aox[16]) );
  NAND2X0_HVT U1329 ( .A1(n12200), .A2(sram_rdata_6[15]), .Y(n1009) );
  NAND3X0_HVT U1330 ( .A1(n448), .A2(n727), .A3(n1009), .Y(n_src_aox[15]) );
  NAND2X0_HVT U1331 ( .A1(n6200), .A2(sram_rdata_6[14]), .Y(n10101) );
  NAND3X0_HVT U1332 ( .A1(n449), .A2(n728), .A3(n10101), .Y(n_src_aox[14]) );
  NAND2X0_HVT U1333 ( .A1(n1053), .A2(sram_rdata_6[13]), .Y(n1011) );
  NAND3X0_HVT U1334 ( .A1(n4501), .A2(n729), .A3(n1011), .Y(n_src_aox[13]) );
  NAND2X0_HVT U1335 ( .A1(n6300), .A2(sram_rdata_6[11]), .Y(n1012) );
  NAND3X0_HVT U1336 ( .A1(n451), .A2(n7301), .A3(n1012), .Y(n_src_aox[11]) );
  NAND2X0_HVT U1337 ( .A1(n13000), .A2(sram_rdata_6[10]), .Y(n1013) );
  NAND3X0_HVT U1338 ( .A1(n452), .A2(n731), .A3(n1013), .Y(n_src_aox[10]) );
  NAND2X0_HVT U1339 ( .A1(n13400), .A2(sram_rdata_6[9]), .Y(n1014) );
  NAND3X0_HVT U1340 ( .A1(n453), .A2(n732), .A3(n1014), .Y(n_src_aox[9]) );
  NAND2X0_HVT U1341 ( .A1(n6000), .A2(sram_rdata_6[8]), .Y(n1015) );
  NAND3X0_HVT U1342 ( .A1(n454), .A2(n733), .A3(n1015), .Y(n_src_aox[8]) );
  NAND2X0_HVT U1343 ( .A1(n12500), .A2(sram_rdata_6[7]), .Y(n1016) );
  NAND3X0_HVT U1344 ( .A1(n455), .A2(n734), .A3(n1016), .Y(n_src_aox[7]) );
  NAND2X0_HVT U1345 ( .A1(n1052), .A2(sram_rdata_6[6]), .Y(n1017) );
  NAND3X0_HVT U1346 ( .A1(n456), .A2(n735), .A3(n1017), .Y(n_src_aox[6]) );
  NAND2X0_HVT U1347 ( .A1(n10501), .A2(sram_rdata_6[5]), .Y(n1018) );
  NAND3X0_HVT U1348 ( .A1(n457), .A2(n736), .A3(n1018), .Y(n_src_aox[5]) );
  NAND2X0_HVT U1349 ( .A1(n10501), .A2(sram_rdata_6[4]), .Y(n1019) );
  NAND3X0_HVT U1350 ( .A1(n458), .A2(n737), .A3(n1019), .Y(n_src_aox[4]) );
  NAND2X0_HVT U1351 ( .A1(n1052), .A2(sram_rdata_6[3]), .Y(n10201) );
  NAND3X0_HVT U1352 ( .A1(n459), .A2(n738), .A3(n10201), .Y(n_src_aox[3]) );
  NAND2X0_HVT U1353 ( .A1(n12700), .A2(sram_rdata_6[2]), .Y(n1021) );
  NAND3X0_HVT U1354 ( .A1(n4601), .A2(n739), .A3(n1021), .Y(n_src_aox[2]) );
  NAND2X0_HVT U1355 ( .A1(n13100), .A2(sram_rdata_6[1]), .Y(n1022) );
  NAND3X0_HVT U1356 ( .A1(n461), .A2(n7401), .A3(n1022), .Y(n_src_aox[1]) );
  NAND2X0_HVT U1357 ( .A1(n38), .A2(n1065), .Y(n1023) );
  NAND3X0_HVT U1358 ( .A1(n1820), .A2(n741), .A3(n1023), .Y(n_src_aox[0]) );
  AND2X1_HVT U1359 ( .A1(box_sel[1]), .A2(box_sel[0]), .Y(n11601) );
  AND2X1_HVT U1360 ( .A1(box_sel[0]), .A2(n1361), .Y(n1161) );
  AND2X1_HVT U1361 ( .A1(box_sel[2]), .A2(n1063), .Y(n1359) );
  AND2X1_HVT U1362 ( .A1(box_sel[1]), .A2(n1062), .Y(n1162) );
  AO222X1_HVT U1363 ( .A1(n8100), .A2(sram_rdata_0[0]), .A3(n8800), .A4(
        sram_rdata_1[0]), .A5(n11400), .A6(sram_rdata_2[0]), .Y(n1065) );
  AND3X1_HVT U1364 ( .A1(n1064), .A2(n1063), .A3(n1062), .Y(n1362) );
  AND2X1_HVT U1365 ( .A1(box_sel[3]), .A2(n1064), .Y(n1357) );
  AO222X1_HVT U1366 ( .A1(n10600), .A2(sram_rdata_3[0]), .A3(n1032), .A4(
        sram_rdata_5[0]), .A5(sram_rdata_4[0]), .A6(n9600), .Y(n1165) );
  AO222X1_HVT U1367 ( .A1(n10900), .A2(sram_rdata_0[1]), .A3(n1161), .A4(
        sram_rdata_2[1]), .A5(sram_rdata_1[1]), .A6(n9100), .Y(n1066) );
  AO222X1_HVT U1368 ( .A1(n1047), .A2(sram_rdata_3[1]), .A3(n1032), .A4(
        sram_rdata_5[1]), .A5(sram_rdata_4[1]), .A6(n9700), .Y(n1167) );
  AO222X1_HVT U1369 ( .A1(n10500), .A2(sram_rdata_0[2]), .A3(n7200), .A4(
        sram_rdata_2[2]), .A5(sram_rdata_1[2]), .A6(n8500), .Y(n1067) );
  AO222X1_HVT U1370 ( .A1(n1048), .A2(sram_rdata_3[2]), .A3(n11600), .A4(
        sram_rdata_5[2]), .A5(sram_rdata_4[2]), .A6(n1024), .Y(n1169) );
  AO222X1_HVT U1371 ( .A1(n8100), .A2(sram_rdata_0[3]), .A3(n7300), .A4(
        sram_rdata_2[3]), .A5(sram_rdata_1[3]), .A6(n8500), .Y(n1068) );
  AO222X1_HVT U1372 ( .A1(n1047), .A2(sram_rdata_3[3]), .A3(n11600), .A4(
        sram_rdata_5[3]), .A5(sram_rdata_4[3]), .A6(n1024), .Y(n1171) );
  AO222X1_HVT U1373 ( .A1(n10600), .A2(sram_rdata_0[4]), .A3(n11200), .A4(
        sram_rdata_2[4]), .A5(sram_rdata_1[4]), .A6(n1025), .Y(n1069) );
  AO222X1_HVT U1374 ( .A1(n1048), .A2(sram_rdata_3[4]), .A3(n11800), .A4(
        sram_rdata_5[4]), .A5(sram_rdata_4[4]), .A6(n1025), .Y(n1173) );
  AO222X1_HVT U1375 ( .A1(n10500), .A2(sram_rdata_0[5]), .A3(n11500), .A4(
        sram_rdata_2[5]), .A5(sram_rdata_1[5]), .A6(n9300), .Y(n10701) );
  AO222X1_HVT U1376 ( .A1(n1048), .A2(sram_rdata_3[5]), .A3(n11100), .A4(
        sram_rdata_5[5]), .A5(sram_rdata_4[5]), .A6(n9200), .Y(n1175) );
  AO222X1_HVT U1377 ( .A1(n6400), .A2(sram_rdata_0[6]), .A3(n11800), .A4(
        sram_rdata_2[6]), .A5(sram_rdata_1[6]), .A6(n9800), .Y(n1071) );
  AO222X1_HVT U1378 ( .A1(n10700), .A2(sram_rdata_3[6]), .A3(n1032), .A4(
        sram_rdata_5[6]), .A5(sram_rdata_4[6]), .A6(n9300), .Y(n1177) );
  AO222X1_HVT U1379 ( .A1(n10800), .A2(sram_rdata_0[7]), .A3(n7300), .A4(
        sram_rdata_2[7]), .A5(sram_rdata_1[7]), .A6(n9000), .Y(n1072) );
  AO222X1_HVT U1380 ( .A1(n8100), .A2(sram_rdata_3[7]), .A3(n1032), .A4(
        sram_rdata_5[7]), .A5(sram_rdata_4[7]), .A6(n9700), .Y(n1179) );
  AO222X1_HVT U1381 ( .A1(n10400), .A2(sram_rdata_0[8]), .A3(n7200), .A4(
        sram_rdata_2[8]), .A5(sram_rdata_1[8]), .A6(n1024), .Y(n1073) );
  AO222X1_HVT U1382 ( .A1(n5200), .A2(sram_rdata_3[8]), .A3(n1161), .A4(
        sram_rdata_5[8]), .A5(sram_rdata_4[8]), .A6(n8500), .Y(n1181) );
  AO222X1_HVT U1383 ( .A1(n8100), .A2(sram_rdata_0[9]), .A3(n1033), .A4(
        sram_rdata_2[9]), .A5(sram_rdata_1[9]), .A6(n8700), .Y(n1074) );
  AO222X1_HVT U1384 ( .A1(n1045), .A2(sram_rdata_3[9]), .A3(n11500), .A4(
        sram_rdata_5[9]), .A5(sram_rdata_4[9]), .A6(n8600), .Y(n1183) );
  AO222X1_HVT U1385 ( .A1(n10900), .A2(sram_rdata_0[10]), .A3(n11300), .A4(
        sram_rdata_2[10]), .A5(sram_rdata_1[10]), .A6(n1024), .Y(n1075) );
  AO222X1_HVT U1386 ( .A1(n8100), .A2(sram_rdata_3[10]), .A3(n12100), .A4(
        sram_rdata_5[10]), .A5(sram_rdata_4[10]), .A6(n8800), .Y(n1185) );
  AO222X1_HVT U1387 ( .A1(n10300), .A2(sram_rdata_0[11]), .A3(n11500), .A4(
        sram_rdata_2[11]), .A5(sram_rdata_1[11]), .A6(n9600), .Y(n1076) );
  AO222X1_HVT U1388 ( .A1(n10800), .A2(sram_rdata_3[11]), .A3(n11200), .A4(
        sram_rdata_5[11]), .A5(sram_rdata_4[11]), .A6(n9200), .Y(n1187) );
  AO222X1_HVT U1389 ( .A1(n1048), .A2(sram_rdata_0[12]), .A3(n12100), .A4(
        sram_rdata_2[12]), .A5(sram_rdata_1[12]), .A6(n10000), .Y(n1077) );
  AO222X1_HVT U1390 ( .A1(n1045), .A2(sram_rdata_3[12]), .A3(n1161), .A4(
        sram_rdata_5[12]), .A5(sram_rdata_4[12]), .A6(n9300), .Y(n1189) );
  AO222X1_HVT U1391 ( .A1(n10700), .A2(sram_rdata_0[13]), .A3(n7300), .A4(
        sram_rdata_2[13]), .A5(sram_rdata_1[13]), .A6(n8900), .Y(n1078) );
  AO222X1_HVT U1392 ( .A1(n6400), .A2(sram_rdata_3[13]), .A3(n10301), .A4(
        sram_rdata_5[13]), .A5(sram_rdata_4[13]), .A6(n9900), .Y(n1191) );
  AO222X1_HVT U1393 ( .A1(n10400), .A2(sram_rdata_0[14]), .A3(n1031), .A4(
        sram_rdata_2[14]), .A5(sram_rdata_1[14]), .A6(n9200), .Y(n1079) );
  AO222X1_HVT U1394 ( .A1(n8100), .A2(sram_rdata_3[14]), .A3(n1031), .A4(
        sram_rdata_5[14]), .A5(sram_rdata_4[14]), .A6(n8700), .Y(n1193) );
  AO222X1_HVT U1395 ( .A1(n1048), .A2(sram_rdata_0[15]), .A3(n1031), .A4(
        sram_rdata_2[15]), .A5(sram_rdata_1[15]), .A6(n9200), .Y(n10801) );
  AO222X1_HVT U1396 ( .A1(n8200), .A2(sram_rdata_3[15]), .A3(n11500), .A4(
        sram_rdata_5[15]), .A5(sram_rdata_4[15]), .A6(n1025), .Y(n1195) );
  AO222X1_HVT U1397 ( .A1(n10700), .A2(sram_rdata_2[0]), .A3(n1025), .A4(
        sram_rdata_0[0]), .A5(n11000), .A6(sram_rdata_1[0]), .Y(n1081) );
  AO222X1_HVT U1398 ( .A1(n8400), .A2(sram_rdata_5[0]), .A3(n11000), .A4(
        sram_rdata_4[0]), .A5(sram_rdata_3[0]), .A6(n10000), .Y(n1197) );
  AO222X1_HVT U1399 ( .A1(n10500), .A2(sram_rdata_2[1]), .A3(n12100), .A4(
        sram_rdata_1[1]), .A5(sram_rdata_0[1]), .A6(n1024), .Y(n1082) );
  AO222X1_HVT U1400 ( .A1(n8400), .A2(sram_rdata_5[1]), .A3(n11700), .A4(
        sram_rdata_4[1]), .A5(sram_rdata_3[1]), .A6(n9500), .Y(n1199) );
  AO222X1_HVT U1401 ( .A1(n8300), .A2(sram_rdata_2[2]), .A3(n11300), .A4(
        sram_rdata_1[2]), .A5(sram_rdata_0[2]), .A6(n9000), .Y(n1083) );
  AO222X1_HVT U1402 ( .A1(n8300), .A2(sram_rdata_5[2]), .A3(n12100), .A4(
        sram_rdata_4[2]), .A5(sram_rdata_3[2]), .A6(n9700), .Y(n1201) );
  AO222X1_HVT U1403 ( .A1(n10800), .A2(sram_rdata_2[3]), .A3(n10301), .A4(
        sram_rdata_1[3]), .A5(sram_rdata_0[3]), .A6(n9600), .Y(n1084) );
  AO222X1_HVT U1404 ( .A1(n1047), .A2(sram_rdata_5[3]), .A3(n11800), .A4(
        sram_rdata_4[3]), .A5(sram_rdata_3[3]), .A6(n8900), .Y(n1203) );
  AO222X1_HVT U1405 ( .A1(n10400), .A2(sram_rdata_2[4]), .A3(n1033), .A4(
        sram_rdata_1[4]), .A5(sram_rdata_0[4]), .A6(n9900), .Y(n1085) );
  AO222X1_HVT U1406 ( .A1(n10900), .A2(sram_rdata_5[4]), .A3(n1161), .A4(
        sram_rdata_4[4]), .A5(sram_rdata_3[4]), .A6(n9500), .Y(n1205) );
  AO222X1_HVT U1407 ( .A1(n1048), .A2(sram_rdata_2[5]), .A3(n11100), .A4(
        sram_rdata_1[5]), .A5(sram_rdata_0[5]), .A6(n8800), .Y(n1086) );
  AO222X1_HVT U1408 ( .A1(n8200), .A2(sram_rdata_5[5]), .A3(n10301), .A4(
        sram_rdata_4[5]), .A5(sram_rdata_3[5]), .A6(n1024), .Y(n1207) );
  AO222X1_HVT U1409 ( .A1(n10900), .A2(sram_rdata_2[6]), .A3(n11500), .A4(
        sram_rdata_1[6]), .A5(sram_rdata_0[6]), .A6(n9200), .Y(n1087) );
  AO222X1_HVT U1410 ( .A1(n8100), .A2(sram_rdata_5[6]), .A3(n11000), .A4(
        sram_rdata_4[6]), .A5(sram_rdata_3[6]), .A6(n9700), .Y(n1209) );
  AO222X1_HVT U1411 ( .A1(n10300), .A2(sram_rdata_2[7]), .A3(n11800), .A4(
        sram_rdata_1[7]), .A5(sram_rdata_0[7]), .A6(n1025), .Y(n1088) );
  AO222X1_HVT U1412 ( .A1(n8300), .A2(sram_rdata_5[7]), .A3(n11400), .A4(
        sram_rdata_4[7]), .A5(sram_rdata_3[7]), .A6(n9600), .Y(n1211) );
  AO222X1_HVT U1413 ( .A1(n1045), .A2(sram_rdata_2[8]), .A3(n11200), .A4(
        sram_rdata_1[8]), .A5(sram_rdata_0[8]), .A6(n9000), .Y(n1089) );
  AO222X1_HVT U1414 ( .A1(n10900), .A2(sram_rdata_5[8]), .A3(n12100), .A4(
        sram_rdata_4[8]), .A5(sram_rdata_3[8]), .A6(n9700), .Y(n1213) );
  AO222X1_HVT U1415 ( .A1(n10900), .A2(sram_rdata_2[9]), .A3(n1032), .A4(
        sram_rdata_1[9]), .A5(sram_rdata_0[9]), .A6(n9400), .Y(n10901) );
  AO222X1_HVT U1416 ( .A1(n1046), .A2(sram_rdata_5[9]), .A3(n1161), .A4(
        sram_rdata_4[9]), .A5(sram_rdata_3[9]), .A6(n9100), .Y(n1215) );
  AO222X1_HVT U1417 ( .A1(n10500), .A2(sram_rdata_2[10]), .A3(n7300), .A4(
        sram_rdata_1[10]), .A5(sram_rdata_0[10]), .A6(n10000), .Y(n1091) );
  AO222X1_HVT U1418 ( .A1(n6400), .A2(sram_rdata_5[10]), .A3(n7300), .A4(
        sram_rdata_4[10]), .A5(sram_rdata_3[10]), .A6(n8500), .Y(n1217) );
  AO222X1_HVT U1419 ( .A1(n8200), .A2(sram_rdata_2[11]), .A3(n1031), .A4(
        sram_rdata_1[11]), .A5(sram_rdata_0[11]), .A6(n9700), .Y(n1092) );
  AO222X1_HVT U1420 ( .A1(n6400), .A2(sram_rdata_5[11]), .A3(n1161), .A4(
        sram_rdata_4[11]), .A5(sram_rdata_3[11]), .A6(n8800), .Y(n1219) );
  AO222X1_HVT U1421 ( .A1(n10600), .A2(sram_rdata_2[12]), .A3(n11500), .A4(
        sram_rdata_1[12]), .A5(sram_rdata_0[12]), .A6(n10000), .Y(n1093) );
  AO222X1_HVT U1422 ( .A1(n1046), .A2(sram_rdata_5[12]), .A3(n11100), .A4(
        sram_rdata_4[12]), .A5(sram_rdata_3[12]), .A6(n8500), .Y(n1221) );
  AO222X1_HVT U1423 ( .A1(n10300), .A2(sram_rdata_2[13]), .A3(n12000), .A4(
        sram_rdata_1[13]), .A5(sram_rdata_0[13]), .A6(n9900), .Y(n1094) );
  AO222X1_HVT U1424 ( .A1(n1047), .A2(sram_rdata_5[13]), .A3(n11400), .A4(
        sram_rdata_4[13]), .A5(sram_rdata_3[13]), .A6(n9600), .Y(n1223) );
  AO222X1_HVT U1425 ( .A1(n1045), .A2(sram_rdata_2[14]), .A3(n11000), .A4(
        sram_rdata_1[14]), .A5(sram_rdata_0[14]), .A6(n8900), .Y(n1095) );
  AO222X1_HVT U1426 ( .A1(n1046), .A2(sram_rdata_5[14]), .A3(n12000), .A4(
        sram_rdata_4[14]), .A5(sram_rdata_3[14]), .A6(n9800), .Y(n1225) );
  AO222X1_HVT U1427 ( .A1(n10900), .A2(sram_rdata_2[15]), .A3(n1032), .A4(
        sram_rdata_1[15]), .A5(sram_rdata_0[15]), .A6(n9600), .Y(n1096) );
  AO222X1_HVT U1428 ( .A1(n1046), .A2(sram_rdata_5[15]), .A3(n7300), .A4(
        sram_rdata_4[15]), .A5(sram_rdata_3[15]), .A6(n9200), .Y(n1227) );
  AO222X1_HVT U1429 ( .A1(n10400), .A2(sram_rdata_1[0]), .A3(n1024), .A4(
        sram_rdata_2[0]), .A5(n11800), .A6(sram_rdata_0[0]), .Y(n1097) );
  AO222X1_HVT U1430 ( .A1(n8400), .A2(sram_rdata_4[0]), .A3(n1032), .A4(
        sram_rdata_3[0]), .A5(n8600), .A6(sram_rdata_5[0]), .Y(n1229) );
  AO222X1_HVT U1431 ( .A1(n6400), .A2(sram_rdata_1[1]), .A3(n1031), .A4(
        sram_rdata_0[1]), .A5(n8800), .A6(sram_rdata_2[1]), .Y(n1098) );
  AO222X1_HVT U1432 ( .A1(n1048), .A2(sram_rdata_4[1]), .A3(n7300), .A4(
        sram_rdata_3[1]), .A5(n8700), .A6(sram_rdata_5[1]), .Y(n1231) );
  AO222X1_HVT U1433 ( .A1(n10800), .A2(sram_rdata_1[2]), .A3(n11300), .A4(
        sram_rdata_0[2]), .A5(n9300), .A6(sram_rdata_2[2]), .Y(n1099) );
  AO222X1_HVT U1434 ( .A1(n1045), .A2(sram_rdata_4[2]), .A3(n11400), .A4(
        sram_rdata_3[2]), .A5(n9000), .A6(sram_rdata_5[2]), .Y(n1233) );
  AO222X1_HVT U1435 ( .A1(n10400), .A2(sram_rdata_1[3]), .A3(n11200), .A4(
        sram_rdata_0[3]), .A5(n9900), .A6(sram_rdata_2[3]), .Y(n11001) );
  AO222X1_HVT U1436 ( .A1(n1162), .A2(sram_rdata_4[3]), .A3(n12100), .A4(
        sram_rdata_3[3]), .A5(n9500), .A6(sram_rdata_5[3]), .Y(n1235) );
  AO222X1_HVT U1437 ( .A1(n8400), .A2(sram_rdata_1[4]), .A3(n11400), .A4(
        sram_rdata_0[4]), .A5(n9000), .A6(sram_rdata_2[4]), .Y(n1101) );
  AO222X1_HVT U1438 ( .A1(n5200), .A2(sram_rdata_4[4]), .A3(n11100), .A4(
        sram_rdata_3[4]), .A5(n9700), .A6(sram_rdata_5[4]), .Y(n1237) );
  AO222X1_HVT U1439 ( .A1(n10700), .A2(sram_rdata_1[5]), .A3(n12000), .A4(
        sram_rdata_0[5]), .A5(n8600), .A6(sram_rdata_2[5]), .Y(n1102) );
  AO222X1_HVT U1440 ( .A1(n6400), .A2(sram_rdata_4[5]), .A3(n1033), .A4(
        sram_rdata_3[5]), .A5(n8700), .A6(sram_rdata_5[5]), .Y(n1239) );
  AO222X1_HVT U1441 ( .A1(n10200), .A2(sram_rdata_1[6]), .A3(n7100), .A4(
        sram_rdata_0[6]), .A5(n9000), .A6(sram_rdata_2[6]), .Y(n1103) );
  AO222X1_HVT U1442 ( .A1(n6400), .A2(sram_rdata_4[6]), .A3(n1031), .A4(
        sram_rdata_3[6]), .A5(n11601), .A6(sram_rdata_5[6]), .Y(n1241) );
  AO222X1_HVT U1443 ( .A1(n1047), .A2(sram_rdata_1[7]), .A3(n7200), .A4(
        sram_rdata_0[7]), .A5(n9300), .A6(sram_rdata_2[7]), .Y(n1104) );
  AO222X1_HVT U1444 ( .A1(n10200), .A2(sram_rdata_4[7]), .A3(n1032), .A4(
        sram_rdata_3[7]), .A5(n8500), .A6(sram_rdata_5[7]), .Y(n1243) );
  AO222X1_HVT U1445 ( .A1(n10600), .A2(sram_rdata_1[8]), .A3(n1032), .A4(
        sram_rdata_0[8]), .A5(n9500), .A6(sram_rdata_2[8]), .Y(n1105) );
  AO222X1_HVT U1446 ( .A1(n1045), .A2(sram_rdata_4[8]), .A3(n11600), .A4(
        sram_rdata_3[8]), .A5(n9200), .A6(sram_rdata_5[8]), .Y(n1245) );
  AO222X1_HVT U1447 ( .A1(n10300), .A2(sram_rdata_1[9]), .A3(n11000), .A4(
        sram_rdata_0[9]), .A5(n9900), .A6(sram_rdata_2[9]), .Y(n1106) );
  AO222X1_HVT U1448 ( .A1(n1046), .A2(sram_rdata_4[9]), .A3(n12000), .A4(
        sram_rdata_3[9]), .A5(n9400), .A6(sram_rdata_5[9]), .Y(n1247) );
  AO222X1_HVT U1449 ( .A1(n8200), .A2(sram_rdata_1[10]), .A3(n11600), .A4(
        sram_rdata_0[10]), .A5(n9100), .A6(sram_rdata_2[10]), .Y(n1107) );
  AO222X1_HVT U1450 ( .A1(n8300), .A2(sram_rdata_4[10]), .A3(n11300), .A4(
        sram_rdata_3[10]), .A5(n9800), .A6(sram_rdata_5[10]), .Y(n1249) );
  AO222X1_HVT U1451 ( .A1(n10700), .A2(sram_rdata_1[11]), .A3(n11900), .A4(
        sram_rdata_0[11]), .A5(n8700), .A6(sram_rdata_2[11]), .Y(n1108) );
  AO222X1_HVT U1452 ( .A1(n8100), .A2(sram_rdata_4[11]), .A3(n11500), .A4(
        sram_rdata_3[11]), .A5(n8600), .A6(sram_rdata_5[11]), .Y(n1251) );
  AO222X1_HVT U1453 ( .A1(n10300), .A2(sram_rdata_1[12]), .A3(n1032), .A4(
        sram_rdata_0[12]), .A5(n8500), .A6(sram_rdata_2[12]), .Y(n1109) );
  AO222X1_HVT U1454 ( .A1(n1048), .A2(sram_rdata_4[12]), .A3(n10301), .A4(
        sram_rdata_3[12]), .A5(n8700), .A6(sram_rdata_5[12]), .Y(n1253) );
  AO222X1_HVT U1455 ( .A1(n5200), .A2(sram_rdata_1[13]), .A3(n12100), .A4(
        sram_rdata_0[13]), .A5(n8600), .A6(sram_rdata_2[13]), .Y(n11101) );
  AO222X1_HVT U1456 ( .A1(n1046), .A2(sram_rdata_4[13]), .A3(n11800), .A4(
        sram_rdata_3[13]), .A5(n8500), .A6(sram_rdata_5[13]), .Y(n1255) );
  AO222X1_HVT U1457 ( .A1(n10600), .A2(sram_rdata_1[14]), .A3(n11500), .A4(
        sram_rdata_0[14]), .A5(n9500), .A6(sram_rdata_2[14]), .Y(n1111) );
  AO222X1_HVT U1458 ( .A1(n5200), .A2(sram_rdata_4[14]), .A3(n11700), .A4(
        sram_rdata_3[14]), .A5(n8900), .A6(sram_rdata_5[14]), .Y(n1257) );
  AO222X1_HVT U1459 ( .A1(n10300), .A2(sram_rdata_1[15]), .A3(n11000), .A4(
        sram_rdata_0[15]), .A5(n9800), .A6(sram_rdata_2[15]), .Y(n1112) );
  AO222X1_HVT U1460 ( .A1(n8400), .A2(sram_rdata_4[15]), .A3(n11900), .A4(
        sram_rdata_3[15]), .A5(n9600), .A6(sram_rdata_5[15]), .Y(n1259) );
  AO222X1_HVT U1461 ( .A1(n8300), .A2(sram_rdata_0[16]), .A3(n11400), .A4(
        sram_rdata_2[16]), .A5(sram_rdata_1[16]), .A6(n9900), .Y(n1113) );
  AO222X1_HVT U1462 ( .A1(n10800), .A2(sram_rdata_3[16]), .A3(n11200), .A4(
        sram_rdata_5[16]), .A5(sram_rdata_4[16]), .A6(n1025), .Y(n1261) );
  AO222X1_HVT U1463 ( .A1(n10900), .A2(sram_rdata_0[17]), .A3(n11900), .A4(
        sram_rdata_2[17]), .A5(sram_rdata_1[17]), .A6(n1024), .Y(n1114) );
  AO222X1_HVT U1464 ( .A1(n6400), .A2(sram_rdata_3[17]), .A3(n1031), .A4(
        sram_rdata_5[17]), .A5(sram_rdata_4[17]), .A6(n1025), .Y(n1263) );
  AO222X1_HVT U1465 ( .A1(n10200), .A2(sram_rdata_0[18]), .A3(n7200), .A4(
        sram_rdata_2[18]), .A5(sram_rdata_1[18]), .A6(n9800), .Y(n1115) );
  AO222X1_HVT U1466 ( .A1(n10900), .A2(sram_rdata_3[18]), .A3(n10301), .A4(
        sram_rdata_5[18]), .A5(sram_rdata_4[18]), .A6(n8500), .Y(n1265) );
  AO222X1_HVT U1467 ( .A1(n10400), .A2(sram_rdata_0[19]), .A3(n1033), .A4(
        sram_rdata_2[19]), .A5(sram_rdata_1[19]), .A6(n9500), .Y(n1116) );
  AO222X1_HVT U1468 ( .A1(n8200), .A2(sram_rdata_3[19]), .A3(n7100), .A4(
        sram_rdata_5[19]), .A5(sram_rdata_4[19]), .A6(n9600), .Y(n1267) );
  AO222X1_HVT U1469 ( .A1(n10800), .A2(sram_rdata_0[20]), .A3(n11000), .A4(
        sram_rdata_2[20]), .A5(sram_rdata_1[20]), .A6(n9100), .Y(n1117) );
  AO222X1_HVT U1470 ( .A1(n5200), .A2(sram_rdata_3[20]), .A3(n11600), .A4(
        sram_rdata_5[20]), .A5(sram_rdata_4[20]), .A6(n9900), .Y(n1269) );
  AO222X1_HVT U1471 ( .A1(n10400), .A2(sram_rdata_0[21]), .A3(n11000), .A4(
        sram_rdata_2[21]), .A5(sram_rdata_1[21]), .A6(n9300), .Y(n1118) );
  AO222X1_HVT U1472 ( .A1(n8100), .A2(sram_rdata_3[21]), .A3(n11900), .A4(
        sram_rdata_5[21]), .A5(sram_rdata_4[21]), .A6(n9200), .Y(n1271) );
  AO222X1_HVT U1473 ( .A1(n1046), .A2(sram_rdata_0[22]), .A3(n11500), .A4(
        sram_rdata_2[22]), .A5(sram_rdata_1[22]), .A6(n10000), .Y(n1119) );
  AO222X1_HVT U1474 ( .A1(n1046), .A2(sram_rdata_3[22]), .A3(n11300), .A4(
        sram_rdata_5[22]), .A5(sram_rdata_4[22]), .A6(n1024), .Y(n1273) );
  AO222X1_HVT U1475 ( .A1(n10700), .A2(sram_rdata_0[23]), .A3(n12000), .A4(
        sram_rdata_2[23]), .A5(sram_rdata_1[23]), .A6(n8600), .Y(n11201) );
  AO222X1_HVT U1476 ( .A1(n1047), .A2(sram_rdata_3[23]), .A3(n7100), .A4(
        sram_rdata_5[23]), .A5(sram_rdata_4[23]), .A6(n8600), .Y(n1275) );
  AO222X1_HVT U1477 ( .A1(n10300), .A2(sram_rdata_0[24]), .A3(n1161), .A4(
        sram_rdata_2[24]), .A5(sram_rdata_1[24]), .A6(n8700), .Y(n1121) );
  AO222X1_HVT U1478 ( .A1(n8400), .A2(sram_rdata_3[24]), .A3(n7100), .A4(
        sram_rdata_5[24]), .A5(sram_rdata_4[24]), .A6(n10000), .Y(n1277) );
  AO222X1_HVT U1479 ( .A1(n8200), .A2(sram_rdata_0[25]), .A3(n12000), .A4(
        sram_rdata_2[25]), .A5(sram_rdata_1[25]), .A6(n8500), .Y(n1122) );
  AO222X1_HVT U1480 ( .A1(n10900), .A2(sram_rdata_3[25]), .A3(n7200), .A4(
        sram_rdata_5[25]), .A5(sram_rdata_4[25]), .A6(n9500), .Y(n1279) );
  AO222X1_HVT U1481 ( .A1(n10600), .A2(sram_rdata_0[26]), .A3(n10301), .A4(
        sram_rdata_2[26]), .A5(sram_rdata_1[26]), .A6(n9100), .Y(n1123) );
  AO222X1_HVT U1482 ( .A1(n8400), .A2(sram_rdata_3[26]), .A3(n11700), .A4(
        sram_rdata_5[26]), .A5(sram_rdata_4[26]), .A6(n9800), .Y(n1281) );
  AO222X1_HVT U1483 ( .A1(n10200), .A2(sram_rdata_0[27]), .A3(n11100), .A4(
        sram_rdata_2[27]), .A5(sram_rdata_1[27]), .A6(n9400), .Y(n1124) );
  AO222X1_HVT U1484 ( .A1(n8100), .A2(sram_rdata_3[27]), .A3(n11900), .A4(
        sram_rdata_5[27]), .A5(sram_rdata_4[27]), .A6(n8900), .Y(n1283) );
  AO222X1_HVT U1485 ( .A1(n5200), .A2(sram_rdata_0[28]), .A3(n11600), .A4(
        sram_rdata_2[28]), .A5(sram_rdata_1[28]), .A6(n9800), .Y(n1125) );
  AO222X1_HVT U1486 ( .A1(n8200), .A2(sram_rdata_3[28]), .A3(n11000), .A4(
        sram_rdata_5[28]), .A5(sram_rdata_4[28]), .A6(n9600), .Y(n1285) );
  AO222X1_HVT U1487 ( .A1(n10900), .A2(sram_rdata_0[29]), .A3(n11800), .A4(
        sram_rdata_2[29]), .A5(sram_rdata_1[29]), .A6(n1025), .Y(n1126) );
  AO222X1_HVT U1488 ( .A1(n8200), .A2(sram_rdata_3[29]), .A3(n12000), .A4(
        sram_rdata_5[29]), .A5(sram_rdata_4[29]), .A6(n8600), .Y(n1287) );
  AO222X1_HVT U1489 ( .A1(n10400), .A2(sram_rdata_0[30]), .A3(n7200), .A4(
        sram_rdata_2[30]), .A5(sram_rdata_1[30]), .A6(n1025), .Y(n1127) );
  AO222X1_HVT U1490 ( .A1(n5200), .A2(sram_rdata_3[30]), .A3(n1161), .A4(
        sram_rdata_5[30]), .A5(sram_rdata_4[30]), .A6(n8700), .Y(n1289) );
  AO222X1_HVT U1491 ( .A1(n10800), .A2(sram_rdata_0[31]), .A3(n1031), .A4(
        sram_rdata_2[31]), .A5(sram_rdata_1[31]), .A6(n1025), .Y(n1128) );
  AO222X1_HVT U1492 ( .A1(n10700), .A2(sram_rdata_3[31]), .A3(n10301), .A4(
        sram_rdata_5[31]), .A5(sram_rdata_4[31]), .A6(n9500), .Y(n1291) );
  AO222X1_HVT U1493 ( .A1(n10800), .A2(sram_rdata_2[16]), .A3(n1032), .A4(
        sram_rdata_1[16]), .A5(sram_rdata_0[16]), .A6(n9000), .Y(n1129) );
  AO222X1_HVT U1494 ( .A1(n8200), .A2(sram_rdata_5[16]), .A3(n11600), .A4(
        sram_rdata_4[16]), .A5(sram_rdata_3[16]), .A6(n9800), .Y(n1293) );
  AO222X1_HVT U1495 ( .A1(n10300), .A2(sram_rdata_2[17]), .A3(n11300), .A4(
        sram_rdata_1[17]), .A5(sram_rdata_0[17]), .A6(n9500), .Y(n11301) );
  AO222X1_HVT U1496 ( .A1(n10800), .A2(sram_rdata_5[17]), .A3(n12100), .A4(
        sram_rdata_4[17]), .A5(sram_rdata_3[17]), .A6(n9000), .Y(n1295) );
  AO222X1_HVT U1497 ( .A1(n10600), .A2(sram_rdata_2[18]), .A3(n11500), .A4(
        sram_rdata_1[18]), .A5(sram_rdata_0[18]), .A6(n9700), .Y(n1131) );
  AO222X1_HVT U1498 ( .A1(n1047), .A2(sram_rdata_5[18]), .A3(n11200), .A4(
        sram_rdata_4[18]), .A5(sram_rdata_3[18]), .A6(n1024), .Y(n1297) );
  AO222X1_HVT U1499 ( .A1(n10600), .A2(sram_rdata_2[19]), .A3(n11900), .A4(
        sram_rdata_1[19]), .A5(sram_rdata_0[19]), .A6(n1025), .Y(n1132) );
  AO222X1_HVT U1500 ( .A1(n8300), .A2(sram_rdata_5[19]), .A3(n1032), .A4(
        sram_rdata_4[19]), .A5(sram_rdata_3[19]), .A6(n9000), .Y(n1299) );
  AO222X1_HVT U1501 ( .A1(n10400), .A2(sram_rdata_2[20]), .A3(n1031), .A4(
        sram_rdata_1[20]), .A5(sram_rdata_0[20]), .A6(n1024), .Y(n1133) );
  AO222X1_HVT U1502 ( .A1(n8300), .A2(sram_rdata_5[20]), .A3(n10301), .A4(
        sram_rdata_4[20]), .A5(sram_rdata_3[20]), .A6(n9100), .Y(n1301) );
  AO222X1_HVT U1503 ( .A1(n6400), .A2(sram_rdata_2[21]), .A3(n1033), .A4(
        sram_rdata_1[21]), .A5(sram_rdata_0[21]), .A6(n9900), .Y(n1134) );
  AO222X1_HVT U1504 ( .A1(n8200), .A2(sram_rdata_5[21]), .A3(n10301), .A4(
        sram_rdata_4[21]), .A5(sram_rdata_3[21]), .A6(n9400), .Y(n1303) );
  AO222X1_HVT U1505 ( .A1(n10800), .A2(sram_rdata_2[22]), .A3(n11900), .A4(
        sram_rdata_1[22]), .A5(sram_rdata_0[22]), .A6(n9000), .Y(n1135) );
  AO222X1_HVT U1506 ( .A1(n10700), .A2(sram_rdata_5[22]), .A3(n11700), .A4(
        sram_rdata_4[22]), .A5(sram_rdata_3[22]), .A6(n10000), .Y(n1305) );
  AO222X1_HVT U1507 ( .A1(n10200), .A2(sram_rdata_2[23]), .A3(n11200), .A4(
        sram_rdata_1[23]), .A5(sram_rdata_0[23]), .A6(n9500), .Y(n1136) );
  AO222X1_HVT U1508 ( .A1(n8100), .A2(sram_rdata_5[23]), .A3(n11800), .A4(
        sram_rdata_4[23]), .A5(sram_rdata_3[23]), .A6(n9100), .Y(n1307) );
  AO222X1_HVT U1509 ( .A1(n1045), .A2(sram_rdata_2[24]), .A3(n11400), .A4(
        sram_rdata_1[24]), .A5(sram_rdata_0[24]), .A6(n9700), .Y(n1137) );
  AO222X1_HVT U1510 ( .A1(n5200), .A2(sram_rdata_5[24]), .A3(n11100), .A4(
        sram_rdata_4[24]), .A5(sram_rdata_3[24]), .A6(n1024), .Y(n1309) );
  AO222X1_HVT U1511 ( .A1(n10800), .A2(sram_rdata_2[25]), .A3(n11800), .A4(
        sram_rdata_1[25]), .A5(sram_rdata_0[25]), .A6(n8600), .Y(n1138) );
  AO222X1_HVT U1512 ( .A1(n10600), .A2(sram_rdata_5[25]), .A3(n1031), .A4(
        sram_rdata_4[25]), .A5(sram_rdata_3[25]), .A6(n1024), .Y(n1311) );
  AO222X1_HVT U1513 ( .A1(n10200), .A2(sram_rdata_2[26]), .A3(n7100), .A4(
        sram_rdata_1[26]), .A5(sram_rdata_0[26]), .A6(n8800), .Y(n1139) );
  AO222X1_HVT U1514 ( .A1(n8300), .A2(sram_rdata_5[26]), .A3(n7200), .A4(
        sram_rdata_4[26]), .A5(sram_rdata_3[26]), .A6(n8600), .Y(n1313) );
  AO222X1_HVT U1515 ( .A1(n1047), .A2(sram_rdata_2[27]), .A3(n7200), .A4(
        sram_rdata_1[27]), .A5(sram_rdata_0[27]), .A6(n8600), .Y(n11401) );
  AO222X1_HVT U1516 ( .A1(n1046), .A2(sram_rdata_5[27]), .A3(n7100), .A4(
        sram_rdata_4[27]), .A5(sram_rdata_3[27]), .A6(n9500), .Y(n1315) );
  AO222X1_HVT U1517 ( .A1(n10900), .A2(sram_rdata_2[28]), .A3(n11000), .A4(
        sram_rdata_1[28]), .A5(sram_rdata_0[28]), .A6(n9000), .Y(n1141) );
  AO222X1_HVT U1518 ( .A1(n8300), .A2(sram_rdata_5[28]), .A3(n11700), .A4(
        sram_rdata_4[28]), .A5(sram_rdata_3[28]), .A6(n10000), .Y(n1317) );
  AO222X1_HVT U1519 ( .A1(n10300), .A2(sram_rdata_2[29]), .A3(n11300), .A4(
        sram_rdata_1[29]), .A5(sram_rdata_0[29]), .A6(n9400), .Y(n1142) );
  AO222X1_HVT U1520 ( .A1(n1046), .A2(sram_rdata_5[29]), .A3(n12100), .A4(
        sram_rdata_4[29]), .A5(sram_rdata_3[29]), .A6(n9200), .Y(n1319) );
  AO222X1_HVT U1521 ( .A1(n8400), .A2(sram_rdata_2[30]), .A3(n11700), .A4(
        sram_rdata_1[30]), .A5(sram_rdata_0[30]), .A6(n9900), .Y(n1143) );
  AO222X1_HVT U1522 ( .A1(n8200), .A2(sram_rdata_5[30]), .A3(n11200), .A4(
        sram_rdata_4[30]), .A5(sram_rdata_3[30]), .A6(n1025), .Y(n1321) );
  AO222X1_HVT U1523 ( .A1(n10700), .A2(sram_rdata_2[31]), .A3(n12100), .A4(
        sram_rdata_1[31]), .A5(sram_rdata_0[31]), .A6(n8700), .Y(n1144) );
  AO222X1_HVT U1524 ( .A1(n8400), .A2(sram_rdata_5[31]), .A3(n1033), .A4(
        sram_rdata_4[31]), .A5(sram_rdata_3[31]), .A6(n9900), .Y(n1323) );
  AO222X1_HVT U1525 ( .A1(n10200), .A2(sram_rdata_1[16]), .A3(n1032), .A4(
        sram_rdata_0[16]), .A5(n8900), .A6(sram_rdata_2[16]), .Y(n1145) );
  AO222X1_HVT U1526 ( .A1(n8100), .A2(sram_rdata_4[16]), .A3(n11100), .A4(
        sram_rdata_3[16]), .A5(n10000), .A6(sram_rdata_5[16]), .Y(n1325) );
  AO222X1_HVT U1527 ( .A1(n8200), .A2(sram_rdata_1[17]), .A3(n1031), .A4(
        sram_rdata_0[17]), .A5(n9600), .A6(sram_rdata_2[17]), .Y(n1146) );
  AO222X1_HVT U1528 ( .A1(n1047), .A2(sram_rdata_4[17]), .A3(n11300), .A4(
        sram_rdata_3[17]), .A5(n8900), .A6(sram_rdata_5[17]), .Y(n1327) );
  AO222X1_HVT U1529 ( .A1(n10800), .A2(sram_rdata_1[18]), .A3(n11700), .A4(
        sram_rdata_0[18]), .A5(n9400), .A6(sram_rdata_2[18]), .Y(n1147) );
  AO222X1_HVT U1530 ( .A1(n6400), .A2(sram_rdata_4[18]), .A3(n11700), .A4(
        sram_rdata_3[18]), .A5(n9100), .A6(sram_rdata_5[18]), .Y(n1329) );
  AO222X1_HVT U1531 ( .A1(n10500), .A2(sram_rdata_1[19]), .A3(n11300), .A4(
        sram_rdata_0[19]), .A5(n11601), .A6(sram_rdata_2[19]), .Y(n1148) );
  AO222X1_HVT U1532 ( .A1(n8100), .A2(sram_rdata_4[19]), .A3(n11900), .A4(
        sram_rdata_3[19]), .A5(n10000), .A6(sram_rdata_5[19]), .Y(n1331) );
  AO222X1_HVT U1533 ( .A1(n1046), .A2(sram_rdata_1[20]), .A3(n11400), .A4(
        sram_rdata_0[20]), .A5(n9500), .A6(sram_rdata_2[20]), .Y(n1149) );
  AO222X1_HVT U1534 ( .A1(n5200), .A2(sram_rdata_4[20]), .A3(n11200), .A4(
        sram_rdata_3[20]), .A5(n9200), .A6(sram_rdata_5[20]), .Y(n1333) );
  AO222X1_HVT U1535 ( .A1(n10700), .A2(sram_rdata_1[21]), .A3(n11800), .A4(
        sram_rdata_0[21]), .A5(n9900), .A6(sram_rdata_2[21]), .Y(n11501) );
  AO222X1_HVT U1536 ( .A1(n1048), .A2(sram_rdata_4[21]), .A3(n11500), .A4(
        sram_rdata_3[21]), .A5(n9500), .A6(sram_rdata_5[21]), .Y(n1335) );
  AO222X1_HVT U1537 ( .A1(n10300), .A2(sram_rdata_1[22]), .A3(n1033), .A4(
        sram_rdata_0[22]), .A5(n9100), .A6(sram_rdata_2[22]), .Y(n1151) );
  AO222X1_HVT U1538 ( .A1(n6400), .A2(sram_rdata_4[22]), .A3(n7200), .A4(
        sram_rdata_3[22]), .A5(n9800), .A6(sram_rdata_5[22]), .Y(n1337) );
  AO222X1_HVT U1539 ( .A1(n8300), .A2(sram_rdata_1[23]), .A3(n7100), .A4(
        sram_rdata_0[23]), .A5(n8800), .A6(sram_rdata_2[23]), .Y(n1152) );
  AO222X1_HVT U1540 ( .A1(n10700), .A2(sram_rdata_4[23]), .A3(n7200), .A4(
        sram_rdata_3[23]), .A5(n1024), .A6(sram_rdata_5[23]), .Y(n1339) );
  AO222X1_HVT U1541 ( .A1(n10900), .A2(sram_rdata_1[24]), .A3(n1033), .A4(
        sram_rdata_0[24]), .A5(n8600), .A6(sram_rdata_2[24]), .Y(n1153) );
  AO222X1_HVT U1542 ( .A1(n1045), .A2(sram_rdata_4[24]), .A3(n11500), .A4(
        sram_rdata_3[24]), .A5(n9200), .A6(sram_rdata_5[24]), .Y(n1341) );
  AO222X1_HVT U1543 ( .A1(n10200), .A2(sram_rdata_1[25]), .A3(n11200), .A4(
        sram_rdata_0[25]), .A5(n8700), .A6(sram_rdata_2[25]), .Y(n1154) );
  AO222X1_HVT U1544 ( .A1(n1047), .A2(sram_rdata_4[25]), .A3(n12100), .A4(
        sram_rdata_3[25]), .A5(n11601), .A6(sram_rdata_5[25]), .Y(n1343) );
  AO222X1_HVT U1545 ( .A1(n10300), .A2(sram_rdata_1[26]), .A3(n11400), .A4(
        sram_rdata_0[26]), .A5(n9400), .A6(sram_rdata_2[26]), .Y(n1155) );
  AO222X1_HVT U1546 ( .A1(n8300), .A2(sram_rdata_4[26]), .A3(n11100), .A4(
        sram_rdata_3[26]), .A5(n9000), .A6(sram_rdata_5[26]), .Y(n1345) );
  AO222X1_HVT U1547 ( .A1(n10700), .A2(sram_rdata_1[27]), .A3(n12100), .A4(
        sram_rdata_0[27]), .A5(n10000), .A6(sram_rdata_2[27]), .Y(n1156) );
  AO222X1_HVT U1548 ( .A1(n8200), .A2(sram_rdata_4[27]), .A3(n11200), .A4(
        sram_rdata_3[27]), .A5(n9300), .A6(sram_rdata_5[27]), .Y(n1347) );
  AO222X1_HVT U1549 ( .A1(n10400), .A2(sram_rdata_1[28]), .A3(n1033), .A4(
        sram_rdata_0[28]), .A5(n9100), .A6(sram_rdata_2[28]), .Y(n1157) );
  AO222X1_HVT U1550 ( .A1(n8400), .A2(sram_rdata_4[28]), .A3(n10301), .A4(
        sram_rdata_3[28]), .A5(n10000), .A6(sram_rdata_5[28]), .Y(n1349) );
  AO222X1_HVT U1551 ( .A1(n1045), .A2(sram_rdata_1[29]), .A3(n1161), .A4(
        sram_rdata_0[29]), .A5(n8800), .A6(sram_rdata_2[29]), .Y(n1158) );
  AO222X1_HVT U1552 ( .A1(n8300), .A2(sram_rdata_4[29]), .A3(n7300), .A4(
        sram_rdata_3[29]), .A5(n9100), .A6(sram_rdata_5[29]), .Y(n1351) );
  AO222X1_HVT U1553 ( .A1(n10900), .A2(sram_rdata_1[30]), .A3(n11200), .A4(
        sram_rdata_0[30]), .A5(n8500), .A6(sram_rdata_2[30]), .Y(n1159) );
  AO222X1_HVT U1554 ( .A1(n1046), .A2(sram_rdata_4[30]), .A3(n11600), .A4(
        sram_rdata_3[30]), .A5(n8700), .A6(sram_rdata_5[30]), .Y(n1353) );
  AO222X1_HVT U1555 ( .A1(n10300), .A2(sram_rdata_1[31]), .A3(n11100), .A4(
        sram_rdata_0[31]), .A5(n8700), .A6(sram_rdata_2[31]), .Y(n1163) );
  AO222X1_HVT U1556 ( .A1(n1047), .A2(sram_rdata_4[31]), .A3(n11800), .A4(
        sram_rdata_3[31]), .A5(n8600), .A6(sram_rdata_5[31]), .Y(n1358) );
  AO222X1_HVT U1557 ( .A1(n1045), .A2(sram_rdata_6[0]), .A3(n11600), .A4(
        sram_rdata_8[0]), .A5(sram_rdata_7[0]), .A6(n8800), .Y(n1164) );
  AO222X1_HVT U1558 ( .A1(n5200), .A2(sram_rdata_6[1]), .A3(n11100), .A4(
        sram_rdata_8[1]), .A5(n9300), .A6(sram_rdata_7[1]), .Y(n1166) );
  AO222X1_HVT U1559 ( .A1(n10900), .A2(sram_rdata_6[2]), .A3(n12000), .A4(
        sram_rdata_8[2]), .A5(n8900), .A6(sram_rdata_7[2]), .Y(n1168) );
  AO222X1_HVT U1560 ( .A1(n10300), .A2(sram_rdata_6[3]), .A3(n12100), .A4(
        sram_rdata_8[3]), .A5(n9700), .A6(sram_rdata_7[3]), .Y(n11701) );
  AO222X1_HVT U1561 ( .A1(n10200), .A2(sram_rdata_6[4]), .A3(n1033), .A4(
        sram_rdata_8[4]), .A5(n9600), .A6(sram_rdata_7[4]), .Y(n1172) );
  AO222X1_HVT U1562 ( .A1(n6400), .A2(sram_rdata_6[5]), .A3(n12100), .A4(
        sram_rdata_8[5]), .A5(n9200), .A6(sram_rdata_7[5]), .Y(n1174) );
  AO222X1_HVT U1563 ( .A1(n8200), .A2(sram_rdata_6[6]), .A3(n7100), .A4(
        sram_rdata_8[6]), .A5(n9700), .A6(sram_rdata_7[6]), .Y(n1176) );
  AO222X1_HVT U1564 ( .A1(n10500), .A2(sram_rdata_6[7]), .A3(n7200), .A4(
        sram_rdata_8[7]), .A5(n8700), .A6(sram_rdata_7[7]), .Y(n1178) );
  AO222X1_HVT U1565 ( .A1(n10800), .A2(sram_rdata_6[8]), .A3(n10301), .A4(
        sram_rdata_8[8]), .A5(n8800), .A6(sram_rdata_7[8]), .Y(n11801) );
  AO222X1_HVT U1566 ( .A1(n10600), .A2(sram_rdata_6[9]), .A3(n11400), .A4(
        sram_rdata_8[9]), .A5(n8500), .A6(sram_rdata_7[9]), .Y(n1182) );
  AO222X1_HVT U1567 ( .A1(n10300), .A2(sram_rdata_6[10]), .A3(n11200), .A4(
        sram_rdata_8[10]), .A5(n8700), .A6(sram_rdata_7[10]), .Y(n1184) );
  AO222X1_HVT U1568 ( .A1(n8400), .A2(sram_rdata_6[11]), .A3(n12000), .A4(
        sram_rdata_8[11]), .A5(n11601), .A6(sram_rdata_7[11]), .Y(n1186) );
  AO222X1_HVT U1569 ( .A1(n1047), .A2(sram_rdata_6[12]), .A3(n11700), .A4(
        sram_rdata_8[12]), .A5(n8600), .A6(sram_rdata_7[12]), .Y(n1188) );
  AO222X1_HVT U1570 ( .A1(n1047), .A2(sram_rdata_6[13]), .A3(n11100), .A4(
        sram_rdata_8[13]), .A5(n9400), .A6(sram_rdata_7[13]), .Y(n11901) );
  AO222X1_HVT U1571 ( .A1(n10700), .A2(sram_rdata_6[14]), .A3(n12000), .A4(
        sram_rdata_8[14]), .A5(n9200), .A6(sram_rdata_7[14]), .Y(n1192) );
  AO222X1_HVT U1572 ( .A1(n1162), .A2(sram_rdata_6[15]), .A3(n1033), .A4(
        sram_rdata_8[15]), .A5(n9700), .A6(sram_rdata_7[15]), .Y(n1194) );
  AO222X1_HVT U1573 ( .A1(n10200), .A2(sram_rdata_8[0]), .A3(n10301), .A4(
        sram_rdata_7[0]), .A5(sram_rdata_6[0]), .A6(n9400), .Y(n1196) );
  AO222X1_HVT U1574 ( .A1(n8200), .A2(sram_rdata_8[1]), .A3(n7300), .A4(
        sram_rdata_7[1]), .A5(n9400), .A6(sram_rdata_6[1]), .Y(n1198) );
  AO222X1_HVT U1575 ( .A1(n10500), .A2(sram_rdata_8[2]), .A3(n7300), .A4(
        sram_rdata_7[2]), .A5(n9000), .A6(sram_rdata_6[2]), .Y(n12001) );
  AO222X1_HVT U1576 ( .A1(n5200), .A2(sram_rdata_8[3]), .A3(n1161), .A4(
        sram_rdata_7[3]), .A5(n10000), .A6(sram_rdata_6[3]), .Y(n1202) );
  AO222X1_HVT U1577 ( .A1(n10700), .A2(sram_rdata_8[4]), .A3(n1033), .A4(
        sram_rdata_7[4]), .A5(n8800), .A6(sram_rdata_6[4]), .Y(n1204) );
  AO222X1_HVT U1578 ( .A1(n5200), .A2(sram_rdata_8[5]), .A3(n11400), .A4(
        sram_rdata_7[5]), .A5(n8800), .A6(sram_rdata_6[5]), .Y(n1206) );
  AO222X1_HVT U1579 ( .A1(n10200), .A2(sram_rdata_8[6]), .A3(n11000), .A4(
        sram_rdata_7[6]), .A5(n8600), .A6(sram_rdata_6[6]), .Y(n1208) );
  AO222X1_HVT U1580 ( .A1(n10300), .A2(sram_rdata_8[7]), .A3(n11900), .A4(
        sram_rdata_7[7]), .A5(n9600), .A6(sram_rdata_6[7]), .Y(n12101) );
  AO222X1_HVT U1581 ( .A1(n8400), .A2(sram_rdata_8[8]), .A3(n11700), .A4(
        sram_rdata_7[8]), .A5(n8900), .A6(sram_rdata_6[8]), .Y(n1212) );
  AO222X1_HVT U1582 ( .A1(n8300), .A2(sram_rdata_8[9]), .A3(n11100), .A4(
        sram_rdata_7[9]), .A5(n8700), .A6(sram_rdata_6[9]), .Y(n1214) );
  AO222X1_HVT U1583 ( .A1(n10600), .A2(sram_rdata_8[10]), .A3(n12000), .A4(
        sram_rdata_7[10]), .A5(n9300), .A6(sram_rdata_6[10]), .Y(n1216) );
  AO222X1_HVT U1584 ( .A1(n1048), .A2(sram_rdata_8[11]), .A3(n7300), .A4(
        sram_rdata_7[11]), .A5(n8900), .A6(sram_rdata_6[11]), .Y(n1218) );
  AO222X1_HVT U1585 ( .A1(n10500), .A2(sram_rdata_8[12]), .A3(n11100), .A4(
        sram_rdata_7[12]), .A5(n9700), .A6(sram_rdata_6[12]), .Y(n12201) );
  AO222X1_HVT U1586 ( .A1(n1047), .A2(sram_rdata_8[13]), .A3(n7200), .A4(
        sram_rdata_7[13]), .A5(n9300), .A6(sram_rdata_6[13]), .Y(n1222) );
  AO222X1_HVT U1587 ( .A1(n10300), .A2(sram_rdata_8[14]), .A3(n10301), .A4(
        sram_rdata_7[14]), .A5(n9100), .A6(sram_rdata_6[14]), .Y(n1224) );
  AO222X1_HVT U1588 ( .A1(n5200), .A2(sram_rdata_8[15]), .A3(n7300), .A4(
        sram_rdata_7[15]), .A5(n9700), .A6(sram_rdata_6[15]), .Y(n1226) );
  AO222X1_HVT U1589 ( .A1(n10600), .A2(sram_rdata_7[0]), .A3(n1161), .A4(
        sram_rdata_6[0]), .A5(n8500), .A6(sram_rdata_8[0]), .Y(n1228) );
  AO222X1_HVT U1590 ( .A1(n8400), .A2(sram_rdata_7[1]), .A3(n11600), .A4(
        sram_rdata_6[1]), .A5(sram_rdata_8[1]), .A6(n1025), .Y(n12301) );
  AO222X1_HVT U1591 ( .A1(n10200), .A2(sram_rdata_7[2]), .A3(n11000), .A4(
        sram_rdata_6[2]), .A5(sram_rdata_8[2]), .A6(n9500), .Y(n1232) );
  AO222X1_HVT U1592 ( .A1(n8300), .A2(sram_rdata_7[3]), .A3(n11900), .A4(
        sram_rdata_6[3]), .A5(sram_rdata_8[3]), .A6(n9200), .Y(n1234) );
  AO222X1_HVT U1593 ( .A1(n8400), .A2(sram_rdata_7[4]), .A3(n11500), .A4(
        sram_rdata_6[4]), .A5(sram_rdata_8[4]), .A6(n10000), .Y(n1236) );
  AO222X1_HVT U1594 ( .A1(n1046), .A2(sram_rdata_7[5]), .A3(n11300), .A4(
        sram_rdata_6[5]), .A5(sram_rdata_8[5]), .A6(n9400), .Y(n1238) );
  AO222X1_HVT U1595 ( .A1(n10800), .A2(sram_rdata_7[6]), .A3(n11900), .A4(
        sram_rdata_6[6]), .A5(sram_rdata_8[6]), .A6(n9100), .Y(n12401) );
  AO222X1_HVT U1596 ( .A1(n1046), .A2(sram_rdata_7[7]), .A3(n11700), .A4(
        sram_rdata_6[7]), .A5(sram_rdata_8[7]), .A6(n9900), .Y(n1242) );
  AO222X1_HVT U1597 ( .A1(n10500), .A2(sram_rdata_7[8]), .A3(n1032), .A4(
        sram_rdata_6[8]), .A5(sram_rdata_8[8]), .A6(n1025), .Y(n1244) );
  AO222X1_HVT U1598 ( .A1(n1047), .A2(sram_rdata_7[9]), .A3(n1031), .A4(
        sram_rdata_6[9]), .A5(sram_rdata_8[9]), .A6(n9600), .Y(n1246) );
  AO222X1_HVT U1599 ( .A1(n8300), .A2(sram_rdata_7[10]), .A3(n11600), .A4(
        sram_rdata_6[10]), .A5(sram_rdata_8[10]), .A6(n9800), .Y(n1248) );
  AO222X1_HVT U1600 ( .A1(n1047), .A2(sram_rdata_7[11]), .A3(n12000), .A4(
        sram_rdata_6[11]), .A5(sram_rdata_8[11]), .A6(n1025), .Y(n12501) );
  AO222X1_HVT U1601 ( .A1(n10900), .A2(sram_rdata_7[12]), .A3(n7100), .A4(
        sram_rdata_6[12]), .A5(sram_rdata_8[12]), .A6(n1025), .Y(n1252) );
  AO222X1_HVT U1602 ( .A1(n5200), .A2(sram_rdata_7[13]), .A3(n11600), .A4(
        sram_rdata_6[13]), .A5(sram_rdata_8[13]), .A6(n9500), .Y(n1254) );
  AO222X1_HVT U1603 ( .A1(n10500), .A2(sram_rdata_7[14]), .A3(n11000), .A4(
        sram_rdata_6[14]), .A5(sram_rdata_8[14]), .A6(n9400), .Y(n1256) );
  AO222X1_HVT U1604 ( .A1(n6400), .A2(sram_rdata_7[15]), .A3(n12000), .A4(
        sram_rdata_6[15]), .A5(sram_rdata_8[15]), .A6(n8900), .Y(n1258) );
  AO222X1_HVT U1605 ( .A1(n8400), .A2(sram_rdata_6[16]), .A3(n11700), .A4(
        sram_rdata_8[16]), .A5(n9800), .A6(sram_rdata_7[16]), .Y(n12601) );
  AO222X1_HVT U1606 ( .A1(n8100), .A2(sram_rdata_6[17]), .A3(n11300), .A4(
        sram_rdata_8[17]), .A5(n8800), .A6(sram_rdata_7[17]), .Y(n1262) );
  AO222X1_HVT U1607 ( .A1(n10600), .A2(sram_rdata_6[18]), .A3(n11800), .A4(
        sram_rdata_8[18]), .A5(n11601), .A6(sram_rdata_7[18]), .Y(n1264) );
  AO222X1_HVT U1608 ( .A1(n1162), .A2(sram_rdata_6[19]), .A3(n7100), .A4(
        sram_rdata_8[19]), .A5(n9000), .A6(sram_rdata_7[19]), .Y(n1266) );
  AO222X1_HVT U1609 ( .A1(n10500), .A2(sram_rdata_6[20]), .A3(n1031), .A4(
        sram_rdata_8[20]), .A5(n9400), .A6(sram_rdata_7[20]), .Y(n1268) );
  AO222X1_HVT U1610 ( .A1(n8100), .A2(sram_rdata_6[21]), .A3(n1033), .A4(
        sram_rdata_8[21]), .A5(n9300), .A6(sram_rdata_7[21]), .Y(n12701) );
  AO222X1_HVT U1611 ( .A1(n6400), .A2(sram_rdata_6[22]), .A3(n7300), .A4(
        sram_rdata_8[22]), .A5(n9200), .A6(sram_rdata_7[22]), .Y(n1272) );
  AO222X1_HVT U1612 ( .A1(n6400), .A2(sram_rdata_6[23]), .A3(n7300), .A4(
        sram_rdata_8[23]), .A5(n10000), .A6(sram_rdata_7[23]), .Y(n1274) );
  AO222X1_HVT U1613 ( .A1(n10800), .A2(sram_rdata_6[24]), .A3(n7200), .A4(
        sram_rdata_8[24]), .A5(n9600), .A6(sram_rdata_7[24]), .Y(n1276) );
  AO222X1_HVT U1614 ( .A1(n10400), .A2(sram_rdata_6[25]), .A3(n11400), .A4(
        sram_rdata_8[25]), .A5(n9100), .A6(sram_rdata_7[25]), .Y(n1278) );
  AO222X1_HVT U1615 ( .A1(n10500), .A2(sram_rdata_6[26]), .A3(n11200), .A4(
        sram_rdata_8[26]), .A5(n9800), .A6(sram_rdata_7[26]), .Y(n12801) );
  AO222X1_HVT U1616 ( .A1(n1048), .A2(sram_rdata_6[27]), .A3(n11900), .A4(
        sram_rdata_8[27]), .A5(n8800), .A6(sram_rdata_7[27]), .Y(n1282) );
  AO222X1_HVT U1617 ( .A1(n1048), .A2(sram_rdata_6[28]), .A3(n11600), .A4(
        sram_rdata_8[28]), .A5(n8500), .A6(sram_rdata_7[28]), .Y(n1284) );
  AO222X1_HVT U1618 ( .A1(n1048), .A2(sram_rdata_6[29]), .A3(n11100), .A4(
        sram_rdata_8[29]), .A5(n8500), .A6(sram_rdata_7[29]), .Y(n1286) );
  AO222X1_HVT U1619 ( .A1(n10700), .A2(sram_rdata_6[30]), .A3(n11900), .A4(
        sram_rdata_8[30]), .A5(n8800), .A6(sram_rdata_7[30]), .Y(n1288) );
  AO222X1_HVT U1620 ( .A1(n10200), .A2(sram_rdata_6[31]), .A3(n11900), .A4(
        sram_rdata_8[31]), .A5(n9100), .A6(sram_rdata_7[31]), .Y(n12901) );
  AO222X1_HVT U1621 ( .A1(n10400), .A2(sram_rdata_8[16]), .A3(n1033), .A4(
        sram_rdata_7[16]), .A5(n8600), .A6(sram_rdata_6[16]), .Y(n1292) );
  AO222X1_HVT U1622 ( .A1(n6400), .A2(sram_rdata_8[17]), .A3(n11700), .A4(
        sram_rdata_7[17]), .A5(n9600), .A6(sram_rdata_6[17]), .Y(n1294) );
  AO222X1_HVT U1623 ( .A1(n1046), .A2(sram_rdata_8[18]), .A3(n11300), .A4(
        sram_rdata_7[18]), .A5(n9000), .A6(sram_rdata_6[18]), .Y(n1296) );
  AO222X1_HVT U1624 ( .A1(n10200), .A2(sram_rdata_8[19]), .A3(n11600), .A4(
        sram_rdata_7[19]), .A5(n9900), .A6(sram_rdata_6[19]), .Y(n1298) );
  AO222X1_HVT U1625 ( .A1(n10600), .A2(sram_rdata_8[20]), .A3(n11900), .A4(
        sram_rdata_7[20]), .A5(n9400), .A6(sram_rdata_6[20]), .Y(n13001) );
  AO222X1_HVT U1626 ( .A1(n1045), .A2(sram_rdata_8[21]), .A3(n11700), .A4(
        sram_rdata_7[21]), .A5(n8900), .A6(sram_rdata_6[21]), .Y(n1302) );
  AO222X1_HVT U1627 ( .A1(n10500), .A2(sram_rdata_8[22]), .A3(n11300), .A4(
        sram_rdata_7[22]), .A5(n9900), .A6(sram_rdata_6[22]), .Y(n1304) );
  AO222X1_HVT U1628 ( .A1(n1045), .A2(sram_rdata_8[23]), .A3(n11800), .A4(
        sram_rdata_7[23]), .A5(n8500), .A6(sram_rdata_6[23]), .Y(n1306) );
  AO222X1_HVT U1629 ( .A1(n8300), .A2(sram_rdata_8[24]), .A3(n11500), .A4(
        sram_rdata_7[24]), .A5(n9500), .A6(sram_rdata_6[24]), .Y(n1308) );
  AO222X1_HVT U1630 ( .A1(n1045), .A2(sram_rdata_8[25]), .A3(n11300), .A4(
        sram_rdata_7[25]), .A5(n9900), .A6(sram_rdata_6[25]), .Y(n13101) );
  AO222X1_HVT U1631 ( .A1(n10800), .A2(sram_rdata_8[26]), .A3(n12000), .A4(
        sram_rdata_7[26]), .A5(n9000), .A6(sram_rdata_6[26]), .Y(n1312) );
  AO222X1_HVT U1632 ( .A1(n1048), .A2(sram_rdata_8[27]), .A3(n1033), .A4(
        sram_rdata_7[27]), .A5(n8800), .A6(sram_rdata_6[27]), .Y(n1314) );
  AO222X1_HVT U1633 ( .A1(n10500), .A2(sram_rdata_8[28]), .A3(n1031), .A4(
        sram_rdata_7[28]), .A5(n11601), .A6(sram_rdata_6[28]), .Y(n1316) );
  AO222X1_HVT U1634 ( .A1(n1048), .A2(sram_rdata_8[29]), .A3(n10301), .A4(
        sram_rdata_7[29]), .A5(n9600), .A6(sram_rdata_6[29]), .Y(n1318) );
  AO222X1_HVT U1635 ( .A1(n10400), .A2(sram_rdata_8[30]), .A3(n7100), .A4(
        sram_rdata_7[30]), .A5(n8900), .A6(sram_rdata_6[30]), .Y(n13201) );
  AO222X1_HVT U1636 ( .A1(n10400), .A2(sram_rdata_8[31]), .A3(n11200), .A4(
        sram_rdata_7[31]), .A5(n9800), .A6(sram_rdata_6[31]), .Y(n1322) );
  AO222X1_HVT U1637 ( .A1(n10700), .A2(sram_rdata_7[16]), .A3(n7200), .A4(
        sram_rdata_6[16]), .A5(sram_rdata_8[16]), .A6(n9900), .Y(n1324) );
  AO222X1_HVT U1638 ( .A1(n1046), .A2(sram_rdata_7[17]), .A3(n11700), .A4(
        sram_rdata_6[17]), .A5(sram_rdata_8[17]), .A6(n9300), .Y(n1326) );
  AO222X1_HVT U1639 ( .A1(n10400), .A2(sram_rdata_7[18]), .A3(n11100), .A4(
        sram_rdata_6[18]), .A5(sram_rdata_8[18]), .A6(n8900), .Y(n1328) );
  AO222X1_HVT U1640 ( .A1(n5200), .A2(sram_rdata_7[19]), .A3(n12100), .A4(
        sram_rdata_6[19]), .A5(sram_rdata_8[19]), .A6(n9800), .Y(n13301) );
  AO222X1_HVT U1641 ( .A1(n10500), .A2(sram_rdata_7[20]), .A3(n11600), .A4(
        sram_rdata_6[20]), .A5(sram_rdata_8[20]), .A6(n1024), .Y(n1332) );
  AO222X1_HVT U1642 ( .A1(n1048), .A2(sram_rdata_7[21]), .A3(n11000), .A4(
        sram_rdata_6[21]), .A5(sram_rdata_8[21]), .A6(n9400), .Y(n1334) );
  AO222X1_HVT U1643 ( .A1(n10600), .A2(sram_rdata_7[22]), .A3(n11800), .A4(
        sram_rdata_6[22]), .A5(sram_rdata_8[22]), .A6(n1024), .Y(n1336) );
  AO222X1_HVT U1644 ( .A1(n10500), .A2(sram_rdata_7[23]), .A3(n10301), .A4(
        sram_rdata_6[23]), .A5(sram_rdata_8[23]), .A6(n9800), .Y(n1338) );
  AO222X1_HVT U1645 ( .A1(n10200), .A2(sram_rdata_7[24]), .A3(n11800), .A4(
        sram_rdata_6[24]), .A5(sram_rdata_8[24]), .A6(n9700), .Y(n13401) );
  AO222X1_HVT U1646 ( .A1(n8400), .A2(sram_rdata_7[25]), .A3(n1031), .A4(
        sram_rdata_6[25]), .A5(sram_rdata_8[25]), .A6(n8700), .Y(n1342) );
  AO222X1_HVT U1647 ( .A1(n8200), .A2(sram_rdata_7[26]), .A3(n7200), .A4(
        sram_rdata_6[26]), .A5(sram_rdata_8[26]), .A6(n9400), .Y(n1344) );
  AO222X1_HVT U1648 ( .A1(n5200), .A2(sram_rdata_7[27]), .A3(n1161), .A4(
        sram_rdata_6[27]), .A5(sram_rdata_8[27]), .A6(n9200), .Y(n1346) );
  AO222X1_HVT U1649 ( .A1(n10600), .A2(sram_rdata_7[28]), .A3(n7300), .A4(
        sram_rdata_6[28]), .A5(sram_rdata_8[28]), .A6(n9800), .Y(n1348) );
  AO222X1_HVT U1650 ( .A1(n8100), .A2(sram_rdata_7[29]), .A3(n11500), .A4(
        sram_rdata_6[29]), .A5(sram_rdata_8[29]), .A6(n9300), .Y(n13501) );
  AO222X1_HVT U1651 ( .A1(n10400), .A2(sram_rdata_7[30]), .A3(n11300), .A4(
        sram_rdata_6[30]), .A5(sram_rdata_8[30]), .A6(n9100), .Y(n1352) );
  AO222X1_HVT U1652 ( .A1(n10200), .A2(sram_rdata_7[31]), .A3(n12000), .A4(
        sram_rdata_6[31]), .A5(sram_rdata_8[31]), .A6(n10000), .Y(n1356) );
  AO22X1_HVT U1653 ( .A1(n1730), .A2(sram_rdata_b1[29]), .A3(n1590), .A4(
        sram_rdata_a1[29]), .Y(N100) );
  AO22X1_HVT U1654 ( .A1(n6700), .A2(sram_rdata_b1[30]), .A3(n1640), .A4(
        sram_rdata_a1[30]), .Y(N101) );
  AO22X1_HVT U1655 ( .A1(n6500), .A2(sram_rdata_b1[31]), .A3(n1550), .A4(
        sram_rdata_a1[31]), .Y(N102) );
  AO22X1_HVT U1656 ( .A1(n1670), .A2(sram_rdata_b2[0]), .A3(n1550), .A4(
        sram_rdata_a2[0]), .Y(N103) );
  AO22X1_HVT U1657 ( .A1(n1720), .A2(sram_rdata_b2[1]), .A3(n1650), .A4(
        sram_rdata_a2[1]), .Y(N104) );
  AO22X1_HVT U1658 ( .A1(n6800), .A2(sram_rdata_b2[2]), .A3(n1550), .A4(
        sram_rdata_a2[2]), .Y(N105) );
  AO22X1_HVT U1659 ( .A1(n6600), .A2(sram_rdata_b2[3]), .A3(n1590), .A4(
        sram_rdata_a2[3]), .Y(N106) );
  AO22X1_HVT U1660 ( .A1(n1680), .A2(sram_rdata_b2[4]), .A3(n1590), .A4(
        sram_rdata_a2[4]), .Y(N107) );
  AO22X1_HVT U1661 ( .A1(n6700), .A2(sram_rdata_b2[5]), .A3(n1560), .A4(
        sram_rdata_a2[5]), .Y(N108) );
  AO22X1_HVT U1662 ( .A1(n27), .A2(sram_rdata_b2[6]), .A3(n1600), .A4(
        sram_rdata_a2[6]), .Y(N109) );
  AO22X1_HVT U1663 ( .A1(n1710), .A2(sram_rdata_b2[7]), .A3(n1640), .A4(
        sram_rdata_a2[7]), .Y(N110) );
  AO22X1_HVT U1664 ( .A1(n6500), .A2(sram_rdata_b2[8]), .A3(n1640), .A4(
        sram_rdata_a2[8]), .Y(N111) );
  AO22X1_HVT U1665 ( .A1(n1710), .A2(sram_rdata_b2[9]), .A3(n1590), .A4(
        sram_rdata_a2[9]), .Y(N112) );
  AO22X1_HVT U1666 ( .A1(n1710), .A2(sram_rdata_b2[10]), .A3(n1630), .A4(
        sram_rdata_a2[10]), .Y(N113) );
  AO22X1_HVT U1667 ( .A1(n1670), .A2(sram_rdata_b2[11]), .A3(n1570), .A4(
        sram_rdata_a2[11]), .Y(N114) );
  AO22X1_HVT U1668 ( .A1(n1670), .A2(sram_rdata_b2[12]), .A3(n1570), .A4(
        sram_rdata_a2[12]), .Y(N115) );
  AO22X1_HVT U1669 ( .A1(n27), .A2(sram_rdata_b2[13]), .A3(n1660), .A4(
        sram_rdata_a2[13]), .Y(N116) );
  AO22X1_HVT U1670 ( .A1(n6800), .A2(sram_rdata_b2[14]), .A3(n1560), .A4(
        sram_rdata_a2[14]), .Y(N117) );
  AO22X1_HVT U1671 ( .A1(n6600), .A2(sram_rdata_b2[15]), .A3(n1600), .A4(
        sram_rdata_a2[15]), .Y(N118) );
  AO22X1_HVT U1672 ( .A1(n1720), .A2(sram_rdata_b2[16]), .A3(n1600), .A4(
        sram_rdata_a2[16]), .Y(N119) );
  AO22X1_HVT U1673 ( .A1(n25), .A2(sram_rdata_b2[17]), .A3(n1560), .A4(
        sram_rdata_a2[17]), .Y(N120) );
  AO22X1_HVT U1674 ( .A1(n25), .A2(sram_rdata_b2[18]), .A3(n1570), .A4(
        sram_rdata_a2[18]), .Y(N121) );
  AO22X1_HVT U1675 ( .A1(n1690), .A2(sram_rdata_b2[19]), .A3(n1650), .A4(
        sram_rdata_a2[19]), .Y(N122) );
  AO22X1_HVT U1676 ( .A1(n1690), .A2(sram_rdata_b2[20]), .A3(n1640), .A4(
        sram_rdata_a2[20]), .Y(N123) );
  AO22X1_HVT U1677 ( .A1(n1710), .A2(sram_rdata_b2[21]), .A3(n1550), .A4(
        sram_rdata_a2[21]), .Y(N124) );
  AO22X1_HVT U1678 ( .A1(n1730), .A2(sram_rdata_b2[22]), .A3(n1610), .A4(
        sram_rdata_a2[22]), .Y(N125) );
  AO22X1_HVT U1679 ( .A1(n1680), .A2(sram_rdata_b2[23]), .A3(n1650), .A4(
        sram_rdata_a2[23]), .Y(N126) );
  AO22X1_HVT U1680 ( .A1(n1670), .A2(sram_rdata_b2[24]), .A3(n1650), .A4(
        sram_rdata_a2[24]), .Y(N127) );
  AO22X1_HVT U1681 ( .A1(n1720), .A2(sram_rdata_b2[25]), .A3(n1640), .A4(
        sram_rdata_a2[25]), .Y(N128) );
  AO22X1_HVT U1682 ( .A1(n6700), .A2(sram_rdata_b2[26]), .A3(n1570), .A4(
        sram_rdata_a2[26]), .Y(N129) );
  AO22X1_HVT U1683 ( .A1(n6500), .A2(sram_rdata_b2[27]), .A3(n1540), .A4(
        sram_rdata_a2[27]), .Y(N130) );
  AO22X1_HVT U1684 ( .A1(n1680), .A2(sram_rdata_b2[28]), .A3(n1540), .A4(
        sram_rdata_a2[28]), .Y(N131) );
  AO22X1_HVT U1685 ( .A1(n1730), .A2(sram_rdata_b2[29]), .A3(n1600), .A4(
        sram_rdata_a2[29]), .Y(N132) );
  AO22X1_HVT U1686 ( .A1(n1730), .A2(sram_rdata_b2[30]), .A3(n1630), .A4(
        sram_rdata_a2[30]), .Y(N133) );
  AO22X1_HVT U1687 ( .A1(n1690), .A2(sram_rdata_b2[31]), .A3(n1600), .A4(
        sram_rdata_a2[31]), .Y(N134) );
  AO22X1_HVT U1688 ( .A1(n6800), .A2(sram_rdata_b3[0]), .A3(n1660), .A4(
        sram_rdata_a3[0]), .Y(N135) );
  AO22X1_HVT U1689 ( .A1(n6800), .A2(sram_rdata_b3[1]), .A3(n1540), .A4(
        sram_rdata_a3[1]), .Y(N136) );
  AO22X1_HVT U1690 ( .A1(n1720), .A2(sram_rdata_b3[2]), .A3(n1570), .A4(
        sram_rdata_a3[2]), .Y(N137) );
  AO22X1_HVT U1691 ( .A1(n1680), .A2(sram_rdata_b3[3]), .A3(n1570), .A4(
        sram_rdata_a3[3]), .Y(N138) );
  AO22X1_HVT U1692 ( .A1(n6600), .A2(sram_rdata_b3[4]), .A3(n1610), .A4(
        sram_rdata_a3[4]), .Y(N139) );
  AO22X1_HVT U1693 ( .A1(n1720), .A2(sram_rdata_b3[5]), .A3(n1590), .A4(
        sram_rdata_a3[5]), .Y(N140) );
  AO22X1_HVT U1694 ( .A1(n27), .A2(sram_rdata_b3[6]), .A3(n1610), .A4(
        sram_rdata_a3[6]), .Y(N141) );
  AO22X1_HVT U1695 ( .A1(n6600), .A2(sram_rdata_b3[7]), .A3(n1660), .A4(
        sram_rdata_a3[7]), .Y(N142) );
  AO22X1_HVT U1696 ( .A1(n1680), .A2(sram_rdata_b3[8]), .A3(n1660), .A4(
        sram_rdata_a3[8]), .Y(N143) );
  AO22X1_HVT U1697 ( .A1(n27), .A2(sram_rdata_b3[9]), .A3(n1630), .A4(
        sram_rdata_a3[9]), .Y(N144) );
  AO22X1_HVT U1698 ( .A1(n6800), .A2(sram_rdata_b3[10]), .A3(n1570), .A4(
        sram_rdata_a3[10]), .Y(N145) );
  AO22X1_HVT U1699 ( .A1(n6600), .A2(sram_rdata_b3[11]), .A3(n1550), .A4(
        sram_rdata_a3[11]), .Y(N146) );
  AO22X1_HVT U1700 ( .A1(n1690), .A2(sram_rdata_b3[12]), .A3(n1540), .A4(
        sram_rdata_a3[12]), .Y(N147) );
  AO22X1_HVT U1701 ( .A1(n27), .A2(sram_rdata_b3[13]), .A3(n1640), .A4(
        sram_rdata_a3[13]), .Y(N148) );
  AO22X1_HVT U1702 ( .A1(n1720), .A2(sram_rdata_b3[14]), .A3(n1650), .A4(
        sram_rdata_a3[14]), .Y(N149) );
  AO22X1_HVT U1703 ( .A1(n1680), .A2(sram_rdata_b3[15]), .A3(n1590), .A4(
        sram_rdata_a3[15]), .Y(N150) );
  AO22X1_HVT U1704 ( .A1(n6800), .A2(sram_rdata_b3[16]), .A3(n1560), .A4(
        sram_rdata_a3[16]), .Y(N151) );
  AO22X1_HVT U1705 ( .A1(n6700), .A2(sram_rdata_b3[17]), .A3(n1540), .A4(
        sram_rdata_a3[17]), .Y(N152) );
  AO22X1_HVT U1706 ( .A1(n1710), .A2(sram_rdata_b3[18]), .A3(n1630), .A4(
        sram_rdata_a3[18]), .Y(N153) );
  AO22X1_HVT U1707 ( .A1(n1670), .A2(sram_rdata_b3[19]), .A3(n1590), .A4(
        sram_rdata_a3[19]), .Y(N154) );
  AO22X1_HVT U1708 ( .A1(n6500), .A2(sram_rdata_b3[20]), .A3(n1610), .A4(
        sram_rdata_a3[20]), .Y(N155) );
  AO22X1_HVT U1709 ( .A1(n25), .A2(sram_rdata_b3[21]), .A3(n1540), .A4(
        sram_rdata_a3[21]), .Y(N156) );
  AO22X1_HVT U1710 ( .A1(n1580), .A2(sram_rdata_b3[22]), .A3(n1550), .A4(
        sram_rdata_a3[22]), .Y(N157) );
  AO22X1_HVT U1711 ( .A1(n1720), .A2(sram_rdata_b3[23]), .A3(n1630), .A4(
        sram_rdata_a3[23]), .Y(N158) );
  AO22X1_HVT U1712 ( .A1(n1690), .A2(sram_rdata_b3[24]), .A3(n1540), .A4(
        sram_rdata_a3[24]), .Y(N159) );
  AO22X1_HVT U1713 ( .A1(n6800), .A2(sram_rdata_b3[25]), .A3(n1600), .A4(
        sram_rdata_a3[25]), .Y(N160) );
  AO22X1_HVT U1714 ( .A1(n25), .A2(sram_rdata_b3[26]), .A3(n1590), .A4(
        sram_rdata_a3[26]), .Y(N161) );
  AO22X1_HVT U1715 ( .A1(n1690), .A2(sram_rdata_b3[27]), .A3(n1640), .A4(
        sram_rdata_a3[27]), .Y(N162) );
  AO22X1_HVT U1716 ( .A1(n6600), .A2(sram_rdata_b3[28]), .A3(n1660), .A4(
        sram_rdata_a3[28]), .Y(N163) );
  AO22X1_HVT U1717 ( .A1(n1730), .A2(sram_rdata_b3[29]), .A3(n1660), .A4(
        sram_rdata_a3[29]), .Y(N164) );
  AO22X1_HVT U1718 ( .A1(n1710), .A2(sram_rdata_b3[30]), .A3(n1550), .A4(
        sram_rdata_a3[30]), .Y(N165) );
  AO22X1_HVT U1719 ( .A1(n1670), .A2(sram_rdata_b3[31]), .A3(n1570), .A4(
        sram_rdata_a3[31]), .Y(N166) );
  AO22X1_HVT U1720 ( .A1(n1690), .A2(sram_rdata_b4[0]), .A3(n1560), .A4(
        sram_rdata_a4[0]), .Y(N167) );
  AO22X1_HVT U1721 ( .A1(n1710), .A2(sram_rdata_b4[1]), .A3(n1600), .A4(
        sram_rdata_a4[1]), .Y(N168) );
  AO22X1_HVT U1722 ( .A1(n25), .A2(sram_rdata_b4[2]), .A3(n1650), .A4(
        sram_rdata_a4[2]), .Y(N169) );
  AO22X1_HVT U1723 ( .A1(n1690), .A2(sram_rdata_b4[3]), .A3(n1590), .A4(
        sram_rdata_a4[3]), .Y(N170) );
  AO22X1_HVT U1724 ( .A1(n1670), .A2(sram_rdata_b4[4]), .A3(n1640), .A4(
        sram_rdata_a4[4]), .Y(N171) );
  AO22X1_HVT U1725 ( .A1(n6800), .A2(sram_rdata_b4[5]), .A3(n1560), .A4(
        sram_rdata_a4[5]), .Y(N172) );
  AO22X1_HVT U1726 ( .A1(n27), .A2(sram_rdata_b4[6]), .A3(n1550), .A4(
        sram_rdata_a4[6]), .Y(N173) );
  AO22X1_HVT U1727 ( .A1(n6600), .A2(sram_rdata_b4[7]), .A3(n1560), .A4(
        sram_rdata_a4[7]), .Y(N174) );
  AO22X1_HVT U1728 ( .A1(n6600), .A2(sram_rdata_b4[8]), .A3(n1640), .A4(
        sram_rdata_a4[8]), .Y(N175) );
  AO22X1_HVT U1729 ( .A1(n6700), .A2(sram_rdata_b4[9]), .A3(n1059), .A4(
        sram_rdata_a4[9]), .Y(N176) );
  AO22X1_HVT U1730 ( .A1(n1720), .A2(sram_rdata_b4[10]), .A3(n1570), .A4(
        sram_rdata_a4[10]), .Y(N177) );
  AO22X1_HVT U1731 ( .A1(n1680), .A2(sram_rdata_b4[11]), .A3(n1630), .A4(
        sram_rdata_a4[11]), .Y(N178) );
  AO22X1_HVT U1732 ( .A1(n6500), .A2(sram_rdata_b4[12]), .A3(n1630), .A4(
        sram_rdata_a4[12]), .Y(N179) );
  AO22X1_HVT U1733 ( .A1(n27), .A2(sram_rdata_b4[13]), .A3(n1650), .A4(
        sram_rdata_a4[13]), .Y(N180) );
  AO22X1_HVT U1734 ( .A1(n6700), .A2(sram_rdata_b4[14]), .A3(n1600), .A4(
        sram_rdata_a4[14]), .Y(N181) );
  AO22X1_HVT U1735 ( .A1(n6500), .A2(sram_rdata_b4[15]), .A3(n1570), .A4(
        sram_rdata_a4[15]), .Y(N182) );
  AO22X1_HVT U1736 ( .A1(n27), .A2(sram_rdata_b4[16]), .A3(n1570), .A4(
        sram_rdata_a4[16]), .Y(N183) );
  AO22X1_HVT U1737 ( .A1(n1720), .A2(sram_rdata_b4[17]), .A3(n1660), .A4(
        sram_rdata_a4[17]), .Y(N184) );
  AO22X1_HVT U1738 ( .A1(n1720), .A2(sram_rdata_b4[18]), .A3(n1630), .A4(
        sram_rdata_a4[18]), .Y(N185) );
  AO22X1_HVT U1739 ( .A1(n1680), .A2(sram_rdata_b4[19]), .A3(n1610), .A4(
        sram_rdata_a4[19]), .Y(N186) );
  AO22X1_HVT U1740 ( .A1(n1680), .A2(sram_rdata_b4[20]), .A3(n1540), .A4(
        sram_rdata_a4[20]), .Y(N187) );
  AO22X1_HVT U1741 ( .A1(n6700), .A2(sram_rdata_b4[21]), .A3(n1560), .A4(
        sram_rdata_a4[21]), .Y(N188) );
  AO22X1_HVT U1742 ( .A1(n1730), .A2(sram_rdata_b4[22]), .A3(n1660), .A4(
        sram_rdata_a4[22]), .Y(N189) );
  AO22X1_HVT U1743 ( .A1(n1690), .A2(sram_rdata_b4[23]), .A3(n1600), .A4(
        sram_rdata_a4[23]), .Y(N190) );
  AO22X1_HVT U1744 ( .A1(n6500), .A2(sram_rdata_b4[24]), .A3(n1660), .A4(
        sram_rdata_a4[24]), .Y(N191) );
  AO22X1_HVT U1745 ( .A1(n1710), .A2(sram_rdata_b4[25]), .A3(n1550), .A4(
        sram_rdata_a4[25]), .Y(N192) );
  AO22X1_HVT U1746 ( .A1(n1710), .A2(sram_rdata_b4[26]), .A3(n1560), .A4(
        sram_rdata_a4[26]), .Y(N193) );
  AO22X1_HVT U1747 ( .A1(n1670), .A2(sram_rdata_b4[27]), .A3(n1640), .A4(
        sram_rdata_a4[27]), .Y(N194) );
  AO22X1_HVT U1748 ( .A1(n1670), .A2(sram_rdata_b4[28]), .A3(n1600), .A4(
        sram_rdata_a4[28]), .Y(N195) );
  AO22X1_HVT U1749 ( .A1(n1730), .A2(sram_rdata_b4[29]), .A3(n1610), .A4(
        sram_rdata_a4[29]), .Y(N196) );
  AO22X1_HVT U1750 ( .A1(n6800), .A2(sram_rdata_b4[30]), .A3(n1059), .A4(
        sram_rdata_a4[30]), .Y(N197) );
  AO22X1_HVT U1751 ( .A1(n6600), .A2(sram_rdata_b4[31]), .A3(n1630), .A4(
        sram_rdata_a4[31]), .Y(N198) );
  AO22X1_HVT U1752 ( .A1(n6700), .A2(sram_rdata_b5[0]), .A3(n1630), .A4(
        sram_rdata_a5[0]), .Y(N199) );
  AO22X1_HVT U1753 ( .A1(n25), .A2(sram_rdata_b5[1]), .A3(n1640), .A4(
        sram_rdata_a5[1]), .Y(N200) );
  AO22X1_HVT U1754 ( .A1(n1710), .A2(sram_rdata_b5[2]), .A3(n1540), .A4(
        sram_rdata_a5[2]), .Y(N201) );
  AO22X1_HVT U1755 ( .A1(n1670), .A2(sram_rdata_b5[3]), .A3(n1550), .A4(
        sram_rdata_a5[3]), .Y(N202) );
  AO22X1_HVT U1756 ( .A1(n1690), .A2(sram_rdata_b5[4]), .A3(n1540), .A4(
        sram_rdata_a5[4]), .Y(N203) );
  AO22X1_HVT U1757 ( .A1(n1710), .A2(sram_rdata_b5[5]), .A3(n1590), .A4(
        sram_rdata_a5[5]), .Y(N204) );
  AO22X1_HVT U1758 ( .A1(n27), .A2(sram_rdata_b5[6]), .A3(n1630), .A4(
        sram_rdata_a5[6]), .Y(N205) );
  AO22X1_HVT U1759 ( .A1(n6500), .A2(sram_rdata_b5[7]), .A3(n1600), .A4(
        sram_rdata_a5[7]), .Y(N206) );
  AO22X1_HVT U1760 ( .A1(n1670), .A2(sram_rdata_b5[8]), .A3(n1640), .A4(
        sram_rdata_a5[8]), .Y(N207) );
  AO22X1_HVT U1761 ( .A1(n1720), .A2(sram_rdata_b5[9]), .A3(n1570), .A4(
        sram_rdata_a5[9]), .Y(N208) );
  AO22X1_HVT U1762 ( .A1(n6700), .A2(sram_rdata_b5[10]), .A3(n1540), .A4(
        sram_rdata_a5[10]), .Y(N209) );
  AO22X1_HVT U1763 ( .A1(n6500), .A2(sram_rdata_b5[11]), .A3(n1560), .A4(
        sram_rdata_a5[11]), .Y(N210) );
  AO22X1_HVT U1764 ( .A1(n1680), .A2(sram_rdata_b5[12]), .A3(n1590), .A4(
        sram_rdata_a5[12]), .Y(N211) );
  AO22X1_HVT U1765 ( .A1(n27), .A2(sram_rdata_b5[13]), .A3(n1600), .A4(
        sram_rdata_a5[13]), .Y(N212) );
  AO22X1_HVT U1766 ( .A1(n1730), .A2(sram_rdata_b5[14]), .A3(n1610), .A4(
        sram_rdata_a5[14]), .Y(N213) );
  AO22X1_HVT U1767 ( .A1(n1690), .A2(sram_rdata_b5[15]), .A3(n1640), .A4(
        sram_rdata_a5[15]), .Y(N214) );
  AO22X1_HVT U1768 ( .A1(n6700), .A2(sram_rdata_b5[16]), .A3(n1640), .A4(
        sram_rdata_a5[16]), .Y(N215) );
  AO22X1_HVT U1769 ( .A1(n6800), .A2(sram_rdata_b5[17]), .A3(n1650), .A4(
        sram_rdata_a5[17]), .Y(N216) );
  AO22X1_HVT U1770 ( .A1(n6700), .A2(sram_rdata_b5[18]), .A3(n1590), .A4(
        sram_rdata_a5[18]), .Y(N217) );
  AO22X1_HVT U1771 ( .A1(n6500), .A2(sram_rdata_b5[19]), .A3(n1550), .A4(
        sram_rdata_a5[19]), .Y(N218) );
  AO22X1_HVT U1772 ( .A1(n6600), .A2(sram_rdata_b5[20]), .A3(n1550), .A4(
        sram_rdata_a5[20]), .Y(N219) );
  AO22X1_HVT U1773 ( .A1(n1720), .A2(sram_rdata_b5[21]), .A3(n1640), .A4(
        sram_rdata_a5[21]), .Y(N220) );
  AO22X1_HVT U1774 ( .A1(n1580), .A2(sram_rdata_b5[22]), .A3(n1650), .A4(
        sram_rdata_a5[22]), .Y(N221) );
  AO22X1_HVT U1775 ( .A1(n1710), .A2(sram_rdata_b5[23]), .A3(n1600), .A4(
        sram_rdata_a5[23]), .Y(N222) );
  AO22X1_HVT U1776 ( .A1(n1680), .A2(sram_rdata_b5[24]), .A3(n1560), .A4(
        sram_rdata_a5[24]), .Y(N223) );
  AO22X1_HVT U1777 ( .A1(n27), .A2(sram_rdata_b5[25]), .A3(n1550), .A4(
        sram_rdata_a5[25]), .Y(N224) );
  AO22X1_HVT U1778 ( .A1(n6800), .A2(sram_rdata_b5[26]), .A3(n1650), .A4(
        sram_rdata_a5[26]), .Y(N225) );
  AO22X1_HVT U1779 ( .A1(n6600), .A2(sram_rdata_b5[27]), .A3(n1590), .A4(
        sram_rdata_a5[27]), .Y(N226) );
  AO22X1_HVT U1780 ( .A1(n1690), .A2(sram_rdata_b5[28]), .A3(n1650), .A4(
        sram_rdata_a5[28]), .Y(N227) );
  AO22X1_HVT U1781 ( .A1(n1730), .A2(sram_rdata_b5[29]), .A3(n1560), .A4(
        sram_rdata_a5[29]), .Y(N228) );
  AO22X1_HVT U1782 ( .A1(n25), .A2(sram_rdata_b5[30]), .A3(n1540), .A4(
        sram_rdata_a5[30]), .Y(N229) );
  AO22X1_HVT U1783 ( .A1(n1690), .A2(sram_rdata_b5[31]), .A3(n1650), .A4(
        sram_rdata_a5[31]), .Y(N230) );
  AO22X1_HVT U1784 ( .A1(n1680), .A2(sram_rdata_b6[0]), .A3(n1610), .A4(
        sram_rdata_a6[0]), .Y(N231) );
  AO22X1_HVT U1785 ( .A1(n6700), .A2(sram_rdata_b6[1]), .A3(n1610), .A4(
        sram_rdata_a6[1]), .Y(N232) );
  AO22X1_HVT U1786 ( .A1(n1720), .A2(sram_rdata_b6[2]), .A3(n1610), .A4(
        sram_rdata_a6[2]), .Y(N233) );
  AO22X1_HVT U1787 ( .A1(n1680), .A2(sram_rdata_b6[3]), .A3(n1660), .A4(
        sram_rdata_a6[3]), .Y(N234) );
  AO22X1_HVT U1788 ( .A1(n6500), .A2(sram_rdata_b6[4]), .A3(n1650), .A4(
        sram_rdata_a6[4]), .Y(N235) );
  AO22X1_HVT U1789 ( .A1(n25), .A2(sram_rdata_b6[5]), .A3(n1660), .A4(
        sram_rdata_a6[5]), .Y(N236) );
  AO22X1_HVT U1790 ( .A1(n6800), .A2(sram_rdata_b6[6]), .A3(n1570), .A4(
        sram_rdata_a6[6]), .Y(N237) );
  AO22X1_HVT U1791 ( .A1(n6600), .A2(sram_rdata_b6[7]), .A3(n1570), .A4(
        sram_rdata_a6[7]), .Y(N238) );
  AO22X1_HVT U1792 ( .A1(n1690), .A2(sram_rdata_b6[8]), .A3(n1560), .A4(
        sram_rdata_a6[8]), .Y(N239) );
  AO22X1_HVT U1793 ( .A1(n6800), .A2(sram_rdata_b6[9]), .A3(n1610), .A4(
        sram_rdata_a6[9]), .Y(N240) );
  AO22X1_HVT U1794 ( .A1(n27), .A2(sram_rdata_b6[10]), .A3(n1650), .A4(
        sram_rdata_a6[10]), .Y(N241) );
  AO22X1_HVT U1795 ( .A1(n6500), .A2(sram_rdata_b6[11]), .A3(n1610), .A4(
        sram_rdata_a6[11]), .Y(N242) );
  AO22X1_HVT U1796 ( .A1(n6600), .A2(sram_rdata_b6[12]), .A3(n1660), .A4(
        sram_rdata_a6[12]), .Y(N243) );
  AO22X1_HVT U1797 ( .A1(n27), .A2(sram_rdata_b6[13]), .A3(n1570), .A4(
        sram_rdata_a6[13]), .Y(N244) );
  AO22X1_HVT U1798 ( .A1(n1720), .A2(sram_rdata_b6[14]), .A3(n1560), .A4(
        sram_rdata_a6[14]), .Y(N245) );
  AO22X1_HVT U1799 ( .A1(n1680), .A2(sram_rdata_b6[15]), .A3(n1570), .A4(
        sram_rdata_a6[15]), .Y(N246) );
  AO22X1_HVT U1800 ( .A1(n1690), .A2(sram_rdata_b6[16]), .A3(n1610), .A4(
        sram_rdata_a6[16]), .Y(N247) );
  AO22X1_HVT U1801 ( .A1(n1710), .A2(sram_rdata_b6[17]), .A3(n1590), .A4(
        sram_rdata_a6[17]), .Y(N248) );
  AO22X1_HVT U1802 ( .A1(n1710), .A2(sram_rdata_b6[18]), .A3(n1590), .A4(
        sram_rdata_a6[18]), .Y(N249) );
  AO22X1_HVT U1803 ( .A1(n1670), .A2(sram_rdata_b6[19]), .A3(n1660), .A4(
        sram_rdata_a6[19]), .Y(N250) );
  AO22X1_HVT U1804 ( .A1(n1670), .A2(sram_rdata_b6[20]), .A3(n1650), .A4(
        sram_rdata_a6[20]), .Y(N251) );
  AO22X1_HVT U1805 ( .A1(n6800), .A2(sram_rdata_b6[21]), .A3(n1630), .A4(
        sram_rdata_a6[21]), .Y(N252) );
  AO22X1_HVT U1806 ( .A1(n25), .A2(sram_rdata_b6[22]), .A3(n1600), .A4(
        sram_rdata_a6[22]), .Y(N253) );
  AO22X1_HVT U1807 ( .A1(n1690), .A2(sram_rdata_b6[23]), .A3(n1570), .A4(
        sram_rdata_a6[23]), .Y(N254) );
  AO22X1_HVT U1808 ( .A1(n6600), .A2(sram_rdata_b6[24]), .A3(n1540), .A4(
        sram_rdata_a6[24]), .Y(N255) );
  AO22X1_HVT U1809 ( .A1(n6700), .A2(sram_rdata_b6[25]), .A3(n1650), .A4(
        sram_rdata_a6[25]), .Y(N256) );
  AO22X1_HVT U1810 ( .A1(n1730), .A2(sram_rdata_b6[26]), .A3(n1630), .A4(
        sram_rdata_a6[26]), .Y(N257) );
  AO22X1_HVT U1811 ( .A1(n27), .A2(sram_rdata_b6[27]), .A3(n1630), .A4(
        sram_rdata_a6[27]), .Y(N258) );
  AO22X1_HVT U1812 ( .A1(n6500), .A2(sram_rdata_b6[28]), .A3(n1540), .A4(
        sram_rdata_a6[28]), .Y(N259) );
  AO22X1_HVT U1813 ( .A1(n1730), .A2(sram_rdata_b6[29]), .A3(n1570), .A4(
        sram_rdata_a6[29]), .Y(N260) );
  AO22X1_HVT U1814 ( .A1(n1710), .A2(sram_rdata_b6[30]), .A3(n1630), .A4(
        sram_rdata_a6[30]), .Y(N261) );
  AO22X1_HVT U1815 ( .A1(n1670), .A2(sram_rdata_b6[31]), .A3(n1540), .A4(
        sram_rdata_a6[31]), .Y(N262) );
  AO22X1_HVT U1816 ( .A1(n27), .A2(sram_rdata_b7[0]), .A3(n1590), .A4(
        sram_rdata_a7[0]), .Y(N263) );
  AO22X1_HVT U1817 ( .A1(n1720), .A2(sram_rdata_b7[1]), .A3(n1550), .A4(
        sram_rdata_a7[1]), .Y(N264) );
  AO22X1_HVT U1818 ( .A1(n6700), .A2(sram_rdata_b7[2]), .A3(n1540), .A4(
        sram_rdata_a7[2]), .Y(N265) );
  AO22X1_HVT U1819 ( .A1(n6500), .A2(sram_rdata_b7[3]), .A3(n1660), .A4(
        sram_rdata_a7[3]), .Y(N266) );
  AO22X1_HVT U1820 ( .A1(n1680), .A2(sram_rdata_b7[4]), .A3(n1600), .A4(
        sram_rdata_a7[4]), .Y(N267) );
  AO22X1_HVT U1821 ( .A1(n6700), .A2(sram_rdata_b7[5]), .A3(n1610), .A4(
        sram_rdata_a7[5]), .Y(N268) );
  AO22X1_HVT U1822 ( .A1(n1720), .A2(sram_rdata_b7[6]), .A3(n1550), .A4(
        sram_rdata_a7[6]), .Y(N269) );
  AO22X1_HVT U1823 ( .A1(n1680), .A2(sram_rdata_b7[7]), .A3(n1640), .A4(
        sram_rdata_a7[7]), .Y(N270) );
  AO22X1_HVT U1824 ( .A1(n6500), .A2(sram_rdata_b7[8]), .A3(n1630), .A4(
        sram_rdata_a7[8]), .Y(N271) );
  AO22X1_HVT U1825 ( .A1(n1710), .A2(sram_rdata_b7[9]), .A3(n1650), .A4(
        sram_rdata_a7[9]), .Y(N272) );
  AO22X1_HVT U1826 ( .A1(n27), .A2(sram_rdata_b7[10]), .A3(n1560), .A4(
        sram_rdata_a7[10]), .Y(N273) );
  AO22X1_HVT U1827 ( .A1(n6700), .A2(sram_rdata_b7[11]), .A3(n1540), .A4(
        sram_rdata_a7[11]), .Y(N274) );
  AO22X1_HVT U1828 ( .A1(n1670), .A2(sram_rdata_b7[12]), .A3(n1560), .A4(
        sram_rdata_a7[12]), .Y(N275) );
  AO22X1_HVT U1829 ( .A1(n27), .A2(sram_rdata_b7[13]), .A3(n1610), .A4(
        sram_rdata_a7[13]), .Y(N276) );
  AO22X1_HVT U1830 ( .A1(n6700), .A2(sram_rdata_b7[14]), .A3(n1660), .A4(
        sram_rdata_a7[14]), .Y(N277) );
  AO22X1_HVT U1831 ( .A1(n6500), .A2(sram_rdata_b7[15]), .A3(n1600), .A4(
        sram_rdata_a7[15]), .Y(N278) );
  AO22X1_HVT U1832 ( .A1(n6500), .A2(sram_rdata_b7[16]), .A3(n1650), .A4(
        sram_rdata_a7[16]), .Y(N279) );
  AO22X1_HVT U1833 ( .A1(n25), .A2(sram_rdata_b7[17]), .A3(n1550), .A4(
        sram_rdata_a7[17]), .Y(N280) );
  AO22X1_HVT U1834 ( .A1(n6800), .A2(sram_rdata_b7[18]), .A3(n1540), .A4(
        sram_rdata_a7[18]), .Y(N281) );
  AO22X1_HVT U1835 ( .A1(n6600), .A2(sram_rdata_b7[19]), .A3(n1570), .A4(
        sram_rdata_a7[19]), .Y(N282) );
  AO22X1_HVT U1836 ( .A1(n1690), .A2(sram_rdata_b7[20]), .A3(n1590), .A4(
        sram_rdata_a7[20]), .Y(N283) );
  AO22X1_HVT U1837 ( .A1(n1710), .A2(sram_rdata_b7[21]), .A3(n1600), .A4(
        sram_rdata_a7[21]), .Y(N284) );
  AO22X1_HVT U1838 ( .A1(n1710), .A2(sram_rdata_b7[22]), .A3(n1590), .A4(
        sram_rdata_a7[22]), .Y(N285) );
  AO22X1_HVT U1839 ( .A1(n1670), .A2(sram_rdata_b7[23]), .A3(n1640), .A4(
        sram_rdata_a7[23]), .Y(N286) );
  AO22X1_HVT U1840 ( .A1(n1670), .A2(sram_rdata_b7[24]), .A3(n1630), .A4(
        sram_rdata_a7[24]), .Y(N287) );
  AO22X1_HVT U1841 ( .A1(n1720), .A2(sram_rdata_b7[25]), .A3(n1640), .A4(
        sram_rdata_a7[25]), .Y(N288) );
  AO22X1_HVT U1842 ( .A1(n1580), .A2(sram_rdata_b7[26]), .A3(n1590), .A4(
        sram_rdata_a7[26]), .Y(N289) );
  AO22X1_HVT U1843 ( .A1(n6600), .A2(sram_rdata_b7[27]), .A3(n1540), .A4(
        sram_rdata_a7[27]), .Y(N290) );
  AO22X1_HVT U1844 ( .A1(n1680), .A2(sram_rdata_b7[28]), .A3(n1540), .A4(
        sram_rdata_a7[28]), .Y(N291) );
  AO22X1_HVT U1845 ( .A1(n1730), .A2(sram_rdata_b7[29]), .A3(n1660), .A4(
        sram_rdata_a7[29]), .Y(N292) );
  AO22X1_HVT U1846 ( .A1(n6800), .A2(sram_rdata_b7[30]), .A3(n1660), .A4(
        sram_rdata_a7[30]), .Y(N293) );
  AO22X1_HVT U1847 ( .A1(n6600), .A2(sram_rdata_b7[31]), .A3(n1590), .A4(
        sram_rdata_a7[31]), .Y(N294) );
  AO22X1_HVT U1848 ( .A1(n27), .A2(sram_rdata_b8[0]), .A3(n1550), .A4(
        sram_rdata_a8[0]), .Y(N295) );
  AO22X1_HVT U1849 ( .A1(n6800), .A2(sram_rdata_b8[1]), .A3(n1550), .A4(
        sram_rdata_a8[1]), .Y(N296) );
  AO22X1_HVT U1850 ( .A1(n1730), .A2(sram_rdata_b8[2]), .A3(n1660), .A4(
        sram_rdata_a8[2]), .Y(N297) );
  AO22X1_HVT U1851 ( .A1(n1690), .A2(sram_rdata_b8[3]), .A3(n1560), .A4(
        sram_rdata_a8[3]), .Y(N298) );
  AO22X1_HVT U1852 ( .A1(n6600), .A2(sram_rdata_b8[4]), .A3(n1630), .A4(
        sram_rdata_a8[4]), .Y(N299) );
  AO22X1_HVT U1853 ( .A1(n1720), .A2(sram_rdata_b8[5]), .A3(n1540), .A4(
        sram_rdata_a8[5]), .Y(N300) );
  AO22X1_HVT U1854 ( .A1(n6700), .A2(sram_rdata_b8[6]), .A3(n1560), .A4(
        sram_rdata_a8[6]), .Y(N301) );
  AO22X1_HVT U1855 ( .A1(n6500), .A2(sram_rdata_b8[7]), .A3(n1640), .A4(
        sram_rdata_a8[7]), .Y(N302) );
  AO22X1_HVT U1856 ( .A1(n1680), .A2(sram_rdata_b8[8]), .A3(n1560), .A4(
        sram_rdata_a8[8]), .Y(N303) );
  AO22X1_HVT U1857 ( .A1(n1620), .A2(sram_rdata_b8[9]), .A3(n1610), .A4(
        sram_rdata_a8[9]), .Y(N304) );
  AO22X1_HVT U1858 ( .A1(n27), .A2(sram_rdata_b8[10]), .A3(n1610), .A4(
        sram_rdata_a8[10]), .Y(N305) );
  AO22X1_HVT U1859 ( .A1(n6700), .A2(sram_rdata_b8[11]), .A3(n1630), .A4(
        sram_rdata_a8[11]), .Y(N306) );
  AO22X1_HVT U1860 ( .A1(n1690), .A2(sram_rdata_b8[12]), .A3(n1640), .A4(
        sram_rdata_a8[12]), .Y(N307) );
  AO22X1_HVT U1861 ( .A1(n27), .A2(sram_rdata_b8[13]), .A3(n1640), .A4(
        sram_rdata_a8[13]), .Y(N308) );
  AO22X1_HVT U1862 ( .A1(n25), .A2(sram_rdata_b8[14]), .A3(n1550), .A4(
        sram_rdata_a8[14]), .Y(N309) );
  AO22X1_HVT U1863 ( .A1(n1690), .A2(sram_rdata_b8[15]), .A3(n1550), .A4(
        sram_rdata_a8[15]), .Y(N310) );
  AO22X1_HVT U1864 ( .A1(n1680), .A2(sram_rdata_b8[16]), .A3(n1550), .A4(
        sram_rdata_a8[16]), .Y(N311) );
  AO22X1_HVT U1865 ( .A1(n6700), .A2(sram_rdata_b8[17]), .A3(n1600), .A4(
        sram_rdata_a8[17]), .Y(N312) );
  AO22X1_HVT U1866 ( .A1(n1720), .A2(sram_rdata_b8[18]), .A3(n1630), .A4(
        sram_rdata_a8[18]), .Y(N313) );
  AO22X1_HVT U1867 ( .A1(n1680), .A2(sram_rdata_b8[19]), .A3(n1600), .A4(
        sram_rdata_a8[19]), .Y(N314) );
  AO22X1_HVT U1868 ( .A1(n6500), .A2(sram_rdata_b8[20]), .A3(n1640), .A4(
        sram_rdata_a8[20]), .Y(N315) );
  AO22X1_HVT U1869 ( .A1(n25), .A2(sram_rdata_b8[21]), .A3(n1570), .A4(
        sram_rdata_a8[21]), .Y(N316) );
  AO22X1_HVT U1870 ( .A1(n6800), .A2(sram_rdata_b8[22]), .A3(n1560), .A4(
        sram_rdata_a8[22]), .Y(N317) );
  AO22X1_HVT U1871 ( .A1(n6600), .A2(sram_rdata_b8[23]), .A3(n1550), .A4(
        sram_rdata_a8[23]), .Y(N318) );
  AO22X1_HVT U1872 ( .A1(n1690), .A2(sram_rdata_b8[24]), .A3(n1600), .A4(
        sram_rdata_a8[24]), .Y(N319) );
  AO22X1_HVT U1873 ( .A1(n6800), .A2(sram_rdata_b8[25]), .A3(n1600), .A4(
        sram_rdata_a8[25]), .Y(N320) );
  AO22X1_HVT U1874 ( .A1(n1730), .A2(sram_rdata_b8[26]), .A3(n1610), .A4(
        sram_rdata_a8[26]), .Y(N321) );
  AO22X1_HVT U1875 ( .A1(n27), .A2(sram_rdata_b8[27]), .A3(n1650), .A4(
        sram_rdata_a8[27]), .Y(N322) );
  AO22X1_HVT U1876 ( .A1(n6600), .A2(sram_rdata_b8[28]), .A3(n1660), .A4(
        sram_rdata_a8[28]), .Y(N323) );
  AO22X1_HVT U1877 ( .A1(n1730), .A2(sram_rdata_b8[29]), .A3(n1650), .A4(
        sram_rdata_a8[29]), .Y(N324) );
  AO22X1_HVT U1878 ( .A1(n1720), .A2(sram_rdata_b8[30]), .A3(n1590), .A4(
        sram_rdata_a8[30]), .Y(N325) );
  AO22X1_HVT U1879 ( .A1(n1680), .A2(sram_rdata_b8[31]), .A3(n1570), .A4(
        sram_rdata_a8[31]), .Y(N326) );
  AO22X1_HVT U1880 ( .A1(n1710), .A2(sram_rdata_b0[0]), .A3(n1560), .A4(
        sram_rdata_a0[0]), .Y(N39) );
  AO22X1_HVT U1881 ( .A1(n1710), .A2(sram_rdata_b0[1]), .A3(n1640), .A4(
        sram_rdata_a0[1]), .Y(N40) );
  AO22X1_HVT U1882 ( .A1(n1710), .A2(sram_rdata_b0[2]), .A3(n1650), .A4(
        sram_rdata_a0[2]), .Y(N41) );
  AO22X1_HVT U1883 ( .A1(n1670), .A2(sram_rdata_b0[3]), .A3(n1590), .A4(
        sram_rdata_a0[3]), .Y(N42) );
  AO22X1_HVT U1884 ( .A1(n1670), .A2(sram_rdata_b0[4]), .A3(n1560), .A4(
        sram_rdata_a0[4]), .Y(N43) );
  AO22X1_HVT U1885 ( .A1(n6800), .A2(sram_rdata_b0[5]), .A3(n1570), .A4(
        sram_rdata_a0[5]), .Y(N44) );
  AO22X1_HVT U1886 ( .A1(n25), .A2(sram_rdata_b0[6]), .A3(n1660), .A4(
        sram_rdata_a0[6]), .Y(N45) );
  AO22X1_HVT U1887 ( .A1(n1690), .A2(sram_rdata_b0[7]), .A3(n1610), .A4(
        sram_rdata_a0[7]), .Y(N46) );
  AO22X1_HVT U1888 ( .A1(n6600), .A2(sram_rdata_b0[8]), .A3(n1610), .A4(
        sram_rdata_a0[8]), .Y(N47) );
  AO22X1_HVT U1889 ( .A1(n6700), .A2(sram_rdata_b0[9]), .A3(n1560), .A4(
        sram_rdata_a0[9]), .Y(N48) );
  AO22X1_HVT U1890 ( .A1(n27), .A2(sram_rdata_b0[10]), .A3(n1540), .A4(
        sram_rdata_a0[10]), .Y(N49) );
  AO22X1_HVT U1891 ( .A1(n6800), .A2(sram_rdata_b0[11]), .A3(n1650), .A4(
        sram_rdata_a0[11]), .Y(N50) );
  AO22X1_HVT U1892 ( .A1(n6500), .A2(sram_rdata_b0[12]), .A3(n1660), .A4(
        sram_rdata_a0[12]), .Y(N51) );
  AO22X1_HVT U1893 ( .A1(n27), .A2(sram_rdata_b0[13]), .A3(n1650), .A4(
        sram_rdata_a0[13]), .Y(N52) );
  AO22X1_HVT U1894 ( .A1(n1710), .A2(sram_rdata_b0[14]), .A3(n1610), .A4(
        sram_rdata_a0[14]), .Y(N53) );
  AO22X1_HVT U1895 ( .A1(n1670), .A2(sram_rdata_b0[15]), .A3(n1650), .A4(
        sram_rdata_a0[15]), .Y(N54) );
  AO22X1_HVT U1896 ( .A1(n6600), .A2(sram_rdata_b0[16]), .A3(n1660), .A4(
        sram_rdata_a0[16]), .Y(N55) );
  AO22X1_HVT U1897 ( .A1(n1720), .A2(sram_rdata_b0[17]), .A3(n1660), .A4(
        sram_rdata_a0[17]), .Y(N56) );
  AO22X1_HVT U1898 ( .A1(n6700), .A2(sram_rdata_b0[18]), .A3(n1570), .A4(
        sram_rdata_a0[18]), .Y(N57) );
  AO22X1_HVT U1899 ( .A1(n6500), .A2(sram_rdata_b0[19]), .A3(n1570), .A4(
        sram_rdata_a0[19]), .Y(N58) );
  AO22X1_HVT U1900 ( .A1(n1680), .A2(sram_rdata_b0[20]), .A3(n1560), .A4(
        sram_rdata_a0[20]), .Y(N59) );
  AO22X1_HVT U1901 ( .A1(n6700), .A2(sram_rdata_b0[21]), .A3(n1600), .A4(
        sram_rdata_a0[21]), .Y(N60) );
  AO22X1_HVT U1902 ( .A1(n1720), .A2(sram_rdata_b0[22]), .A3(n1650), .A4(
        sram_rdata_a0[22]), .Y(N61) );
  AO22X1_HVT U1903 ( .A1(n1680), .A2(sram_rdata_b0[23]), .A3(n1590), .A4(
        sram_rdata_a0[23]), .Y(N62) );
  AO22X1_HVT U1904 ( .A1(n6500), .A2(sram_rdata_b0[24]), .A3(n1630), .A4(
        sram_rdata_a0[24]), .Y(N63) );
  AO22X1_HVT U1905 ( .A1(n1710), .A2(sram_rdata_b0[25]), .A3(n1550), .A4(
        sram_rdata_a0[25]), .Y(N64) );
  AO22X1_HVT U1906 ( .A1(n1730), .A2(sram_rdata_b0[26]), .A3(n1540), .A4(
        sram_rdata_a0[26]), .Y(N65) );
  AO22X1_HVT U1907 ( .A1(n6500), .A2(sram_rdata_b0[27]), .A3(n1540), .A4(
        sram_rdata_a0[27]), .Y(N66) );
  AO22X1_HVT U1908 ( .A1(n1670), .A2(sram_rdata_b0[28]), .A3(n1600), .A4(
        sram_rdata_a0[28]), .Y(N67) );
  AO22X1_HVT U1909 ( .A1(n6500), .A2(sram_rdata_b0[29]), .A3(n1590), .A4(
        sram_rdata_a0[29]), .Y(N68) );
  AO22X1_HVT U1910 ( .A1(n6700), .A2(sram_rdata_b0[30]), .A3(n1600), .A4(
        sram_rdata_a0[30]), .Y(N69) );
  AO22X1_HVT U1911 ( .A1(n1730), .A2(sram_rdata_b0[31]), .A3(n1630), .A4(
        sram_rdata_a0[31]), .Y(N70) );
  AO22X1_HVT U1912 ( .A1(n1670), .A2(sram_rdata_b1[0]), .A3(n1660), .A4(
        sram_rdata_a1[0]), .Y(N71) );
  AO22X1_HVT U1913 ( .A1(n25), .A2(sram_rdata_b1[1]), .A3(n1630), .A4(
        sram_rdata_a1[1]), .Y(N72) );
  AO22X1_HVT U1914 ( .A1(n6800), .A2(sram_rdata_b1[2]), .A3(n1600), .A4(
        sram_rdata_a1[2]), .Y(N73) );
  AO22X1_HVT U1915 ( .A1(n6600), .A2(sram_rdata_b1[3]), .A3(n1570), .A4(
        sram_rdata_a1[3]), .Y(N74) );
  AO22X1_HVT U1916 ( .A1(n1690), .A2(sram_rdata_b1[4]), .A3(n1550), .A4(
        sram_rdata_a1[4]), .Y(N75) );
  AO22X1_HVT U1917 ( .A1(n1670), .A2(sram_rdata_b1[5]), .A3(n1660), .A4(
        sram_rdata_a1[5]), .Y(N76) );
  AO22X1_HVT U1918 ( .A1(n1710), .A2(sram_rdata_b1[6]), .A3(n1630), .A4(
        sram_rdata_a1[6]), .Y(N77) );
  AO22X1_HVT U1919 ( .A1(n1710), .A2(sram_rdata_b1[7]), .A3(n1600), .A4(
        sram_rdata_a1[7]), .Y(N78) );
  AO22X1_HVT U1920 ( .A1(n1670), .A2(sram_rdata_b1[8]), .A3(n1540), .A4(
        sram_rdata_a1[8]), .Y(N79) );
  AO22X1_HVT U1921 ( .A1(n6800), .A2(sram_rdata_b1[9]), .A3(n1550), .A4(
        sram_rdata_a1[9]), .Y(N80) );
  AO22X1_HVT U1922 ( .A1(n27), .A2(sram_rdata_b1[10]), .A3(n1640), .A4(
        sram_rdata_a1[10]), .Y(N81) );
  AO22X1_HVT U1923 ( .A1(n1720), .A2(sram_rdata_b1[11]), .A3(n1610), .A4(
        sram_rdata_a1[11]), .Y(N82) );
  AO22X1_HVT U1924 ( .A1(n1680), .A2(sram_rdata_b1[12]), .A3(n1610), .A4(
        sram_rdata_a1[12]), .Y(N83) );
  AO22X1_HVT U1925 ( .A1(n6600), .A2(sram_rdata_b1[13]), .A3(n1570), .A4(
        sram_rdata_a1[13]), .Y(N84) );
  AO22X1_HVT U1926 ( .A1(n6800), .A2(sram_rdata_b1[14]), .A3(n1560), .A4(
        sram_rdata_a1[14]), .Y(N85) );
  AO22X1_HVT U1927 ( .A1(n27), .A2(sram_rdata_b1[15]), .A3(n1630), .A4(
        sram_rdata_a1[15]), .Y(N86) );
  AO22X1_HVT U1928 ( .A1(n1670), .A2(sram_rdata_b1[16]), .A3(n1610), .A4(
        sram_rdata_a1[16]), .Y(N87) );
  AO22X1_HVT U1929 ( .A1(n1690), .A2(sram_rdata_b1[17]), .A3(n1610), .A4(
        sram_rdata_a1[17]), .Y(N88) );
  AO22X1_HVT U1930 ( .A1(n25), .A2(sram_rdata_b1[18]), .A3(n1590), .A4(
        sram_rdata_a1[18]), .Y(N89) );
  AO22X1_HVT U1931 ( .A1(n6800), .A2(sram_rdata_b1[19]), .A3(n1650), .A4(
        sram_rdata_a1[19]), .Y(N90) );
  AO22X1_HVT U1932 ( .A1(n6600), .A2(sram_rdata_b1[20]), .A3(n1640), .A4(
        sram_rdata_a1[20]), .Y(N91) );
  AO22X1_HVT U1933 ( .A1(n1720), .A2(sram_rdata_b1[21]), .A3(n1640), .A4(
        sram_rdata_a1[21]), .Y(N92) );
  AO22X1_HVT U1934 ( .A1(n6700), .A2(sram_rdata_b1[22]), .A3(n1560), .A4(
        sram_rdata_a1[22]), .Y(N93) );
  AO22X1_HVT U1935 ( .A1(n6500), .A2(sram_rdata_b1[23]), .A3(n1550), .A4(
        sram_rdata_a1[23]), .Y(N94) );
  AO22X1_HVT U1936 ( .A1(n1680), .A2(sram_rdata_b1[24]), .A3(n1540), .A4(
        sram_rdata_a1[24]), .Y(N95) );
  AO22X1_HVT U1937 ( .A1(n1580), .A2(sram_rdata_b1[25]), .A3(n1610), .A4(
        sram_rdata_a1[25]), .Y(N96) );
  AO22X1_HVT U1938 ( .A1(n1730), .A2(sram_rdata_b1[26]), .A3(n1630), .A4(
        sram_rdata_a1[26]), .Y(N97) );
  AO22X1_HVT U1939 ( .A1(n1720), .A2(sram_rdata_b1[27]), .A3(n1590), .A4(
        sram_rdata_a1[27]), .Y(N98) );
  AO22X1_HVT U1940 ( .A1(n1690), .A2(sram_rdata_b1[28]), .A3(n1660), .A4(
        sram_rdata_a1[28]), .Y(N99) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_0 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19092, n1;

  AND2X1_HVT main_gate ( .A1(net19092), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n1), .D(EN), .Q(net19092) );
  INVX0_HVT U1 ( .A(CLK), .Y(n1) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_20 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19092, n2;

  AND2X1_HVT main_gate ( .A1(net19092), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19092) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_19 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19092, n2;

  AND2X1_HVT main_gate ( .A1(net19092), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19092) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_18 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19092, n2;

  AND2X1_HVT main_gate ( .A1(net19092), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19092) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_17 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19092, n2;

  AND2X1_HVT main_gate ( .A1(net19092), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19092) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_16 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19092, n2;

  AND2X1_HVT main_gate ( .A1(net19092), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19092) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_15 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19092, n2;

  AND2X1_HVT main_gate ( .A1(net19092), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19092) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_14 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19092, n2;

  AND2X1_HVT main_gate ( .A1(net19092), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19092) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_13 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19092, n2;

  AND2X1_HVT main_gate ( .A1(net19092), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19092) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_12 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19092, n2;

  AND2X1_HVT main_gate ( .A1(net19092), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19092) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_11 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19092, n2;

  AND2X1_HVT main_gate ( .A1(net19092), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19092) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_10 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19092, n2;

  AND2X1_HVT main_gate ( .A1(net19092), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19092) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_9 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19092, n2;

  AND2X1_HVT main_gate ( .A1(net19092), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19092) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_8 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19092, n2;

  AND2X1_HVT main_gate ( .A1(net19092), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19092) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_7 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19092, n2;

  AND2X1_HVT main_gate ( .A1(net19092), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19092) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_6 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19092, n2;

  AND2X1_HVT main_gate ( .A1(net19092), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19092) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_5 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19092, n2;

  AND2X1_HVT main_gate ( .A1(net19092), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19092) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_4 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19092, n2;

  AND2X1_HVT main_gate ( .A1(net19092), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19092) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_3 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19092, n2;

  AND2X1_HVT main_gate ( .A1(net19092), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19092) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_2 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19092, n2;

  AND2X1_HVT main_gate ( .A1(net19092), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19092) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_1 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net19092, n2;

  AND2X1_HVT main_gate ( .A1(net19092), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net19092) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module bias_sel ( clk, srstn, mode, load_conv1_bias_enable, 
        load_conv2_bias0_enable, load_conv2_bias1_enable, sram_rdata_weight, 
        bias_data, conv1_bias_set_5_, conv1_bias_set_4_, conv1_bias_set_3_, 
        conv1_bias_set_2_, conv1_bias_set_1_, conv1_bias_set_0_, set_5_, 
        set_4_, set_3_, set_2_, set_1_, set_0_ );
  input [1:0] mode;
  input [99:0] sram_rdata_weight;
  output [3:0] bias_data;
  input clk, srstn, load_conv1_bias_enable, load_conv2_bias0_enable,
         load_conv2_bias1_enable, conv1_bias_set_5_, conv1_bias_set_4_,
         conv1_bias_set_3_, conv1_bias_set_2_, conv1_bias_set_1_,
         conv1_bias_set_0_, set_5_, set_4_, set_3_, set_2_, set_1_, set_0_;
  wire   net19121, net19124, net19125, net19126, net19127, net19128, net19129,
         net19130, net19131, net19132, net19135, net19140, net19141, net19142,
         net19143, net19144, net19145, net19146, net19147, net19148, net19149,
         net19152, net19157, net19158, net19159, net19160, net19161, net19162,
         net19163, net19164, net19165, net19166, net19169, net19174, net19175,
         net19176, net19177, net19178, net19179, net19180, net19181, net19182,
         net19183, net19186, net19191, net19192, net19193, net19194, net19195,
         net19196, net19197, net19198, net19199, net19200, net19203, net19208,
         net19209, net19210, net19211, net19212, net19213, net19214, net19215,
         net19216, net19217, net19220, net19225, net19226, net19227, net19228,
         net19229, net19230, net19231, net19232, net19233, net19234, net19237,
         net19242, net19243, net19244, net19245, net19246, net19247, net19248,
         net19249, net19250, net19251, net19254, net19259, net19260, net19261,
         net19262, net19263, net19264, net19265, net19266, net19267, net19268,
         net19271, net19275, net19276, net19277, net19278, net19279, net19280,
         net19281, net19282, net19283, net19284, net19285, net19288, net19301,
         net19302, net19303, net19304, net19305, net19306, net19307, net19308,
         net19309, net19310, net19313, net19318, net19319, net19320, net19321,
         net19322, net19323, net19324, net19325, net19326, net19327, net19330,
         net19335, net19336, net19337, net19338, net19339, net19340, net19341,
         net19342, net19343, net19344, net19347, net19352, net19353, net19354,
         net19355, net19356, net19357, net19358, net19359, net19360, net19361,
         net19364, net19369, net19370, net19371, net19372, net19373, net19374,
         net19375, net19376, net19377, net19378, net19381, net19386, net19387,
         net19388, net19389, net19390, net19391, net19392, net19393, net19394,
         net19395, net19398, net19403, net19404, net19405, net19406, net19407,
         net19408, net19409, net19410, net19411, net19412, net19415, net19420,
         net19421, net19422, net19423, net19424, net19425, net19426, net19427,
         net19428, net19429, net19432, net19437, net19438, net19439, net19440,
         net19441, net19442, net19443, net19444, net19445, net19446, net19449,
         net19453, net19454, net19455, net19456, net19457, net19458, net19459,
         net19460, net19461, net19462, net19463, net19466, net19477, net19483,
         net19487, net19491, net19495, net19498, n305, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401;
  wire   [199:0] conv_weight_box;
  wire   [99:0] delay_weight;

  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_0 clk_gate_conv_weight_box_reg_0_ ( 
        .CLK(clk), .EN(net19275), .ENCLK(net19135) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_20 clk_gate_conv_weight_box_reg_2_ ( 
        .CLK(clk), .EN(net19275), .ENCLK(net19152) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_19 clk_gate_conv_weight_box_reg_5_ ( 
        .CLK(clk), .EN(net19275), .ENCLK(net19169) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_18 clk_gate_conv_weight_box_reg_7_ ( 
        .CLK(clk), .EN(net19275), .ENCLK(net19186) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_17 clk_gate_conv_weight_box_reg_10_ ( 
        .CLK(clk), .EN(net19275), .ENCLK(net19203) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_16 clk_gate_conv_weight_box_reg_12_ ( 
        .CLK(clk), .EN(net19275), .ENCLK(net19220) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_15 clk_gate_conv_weight_box_reg_15_ ( 
        .CLK(clk), .EN(net19275), .ENCLK(net19237) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_14 clk_gate_conv_weight_box_reg_17_ ( 
        .CLK(clk), .EN(net19275), .ENCLK(net19254) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_13 clk_gate_conv_weight_box_reg_20_ ( 
        .CLK(clk), .EN(net19275), .ENCLK(net19271) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_12 clk_gate_conv_weight_box_reg_22_ ( 
        .CLK(clk), .EN(net19275), .ENCLK(net19288) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_11 clk_gate_conv_weight_box_reg_25_ ( 
        .CLK(clk), .EN(net19453), .ENCLK(net19313) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_10 clk_gate_conv_weight_box_reg_27_ ( 
        .CLK(clk), .EN(net19453), .ENCLK(net19330) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_9 clk_gate_conv_weight_box_reg_30_ ( 
        .CLK(clk), .EN(net19453), .ENCLK(net19347) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_8 clk_gate_conv_weight_box_reg_32_ ( 
        .CLK(clk), .EN(net19453), .ENCLK(net19364) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_7 clk_gate_conv_weight_box_reg_35_ ( 
        .CLK(clk), .EN(net19453), .ENCLK(net19381) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_6 clk_gate_conv_weight_box_reg_37_ ( 
        .CLK(clk), .EN(net19453), .ENCLK(net19398) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_5 clk_gate_conv_weight_box_reg_40_ ( 
        .CLK(clk), .EN(net19453), .ENCLK(net19415) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_4 clk_gate_conv_weight_box_reg_42_ ( 
        .CLK(clk), .EN(net19453), .ENCLK(net19432) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_3 clk_gate_conv_weight_box_reg_45_ ( 
        .CLK(clk), .EN(net19453), .ENCLK(net19449) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_2 clk_gate_conv_weight_box_reg_47_ ( 
        .CLK(clk), .EN(net19453), .ENCLK(net19466) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_1 clk_gate_bias_data_reg ( .CLK(clk), 
        .EN(net19477), .ENCLK(net19498) );
  DFFSSRX1_HVT delay_weight_reg_99_ ( .D(1'b0), .SETB(n297), .RSTB(
        sram_rdata_weight[99]), .CLK(clk), .Q(delay_weight[99]) );
  DFFSSRX1_HVT delay_weight_reg_98_ ( .D(1'b0), .SETB(n293), .RSTB(
        sram_rdata_weight[98]), .CLK(clk), .Q(delay_weight[98]) );
  DFFSSRX1_HVT delay_weight_reg_97_ ( .D(1'b0), .SETB(n303), .RSTB(
        sram_rdata_weight[97]), .CLK(clk), .Q(delay_weight[97]) );
  DFFSSRX1_HVT delay_weight_reg_96_ ( .D(1'b0), .SETB(n298), .RSTB(
        sram_rdata_weight[96]), .CLK(clk), .Q(delay_weight[96]) );
  DFFSSRX1_HVT delay_weight_reg_95_ ( .D(1'b0), .SETB(n294), .RSTB(
        sram_rdata_weight[95]), .CLK(clk), .Q(delay_weight[95]) );
  DFFSSRX1_HVT delay_weight_reg_94_ ( .D(1'b0), .SETB(n306), .RSTB(
        sram_rdata_weight[94]), .CLK(clk), .Q(delay_weight[94]) );
  DFFSSRX1_HVT delay_weight_reg_93_ ( .D(1'b0), .SETB(n299), .RSTB(
        sram_rdata_weight[93]), .CLK(clk), .Q(delay_weight[93]) );
  DFFSSRX1_HVT delay_weight_reg_92_ ( .D(1'b0), .SETB(n295), .RSTB(
        sram_rdata_weight[92]), .CLK(clk), .Q(delay_weight[92]) );
  DFFSSRX1_HVT delay_weight_reg_91_ ( .D(1'b0), .SETB(n301), .RSTB(
        sram_rdata_weight[91]), .CLK(clk), .Q(delay_weight[91]) );
  DFFSSRX1_HVT delay_weight_reg_90_ ( .D(1'b0), .SETB(n296), .RSTB(
        sram_rdata_weight[90]), .CLK(clk), .Q(delay_weight[90]) );
  DFFSSRX1_HVT delay_weight_reg_89_ ( .D(1'b0), .SETB(n295), .RSTB(
        sram_rdata_weight[89]), .CLK(clk), .Q(delay_weight[89]) );
  DFFSSRX1_HVT delay_weight_reg_88_ ( .D(1'b0), .SETB(n302), .RSTB(
        sram_rdata_weight[88]), .CLK(clk), .Q(delay_weight[88]) );
  DFFSSRX1_HVT delay_weight_reg_87_ ( .D(1'b0), .SETB(n297), .RSTB(
        sram_rdata_weight[87]), .CLK(clk), .Q(delay_weight[87]) );
  DFFSSRX1_HVT delay_weight_reg_86_ ( .D(1'b0), .SETB(n293), .RSTB(
        sram_rdata_weight[86]), .CLK(clk), .Q(delay_weight[86]) );
  DFFSSRX1_HVT delay_weight_reg_85_ ( .D(1'b0), .SETB(n303), .RSTB(
        sram_rdata_weight[85]), .CLK(clk), .Q(delay_weight[85]) );
  DFFSSRX1_HVT delay_weight_reg_84_ ( .D(1'b0), .SETB(n298), .RSTB(
        sram_rdata_weight[84]), .CLK(clk), .Q(delay_weight[84]) );
  DFFSSRX1_HVT delay_weight_reg_83_ ( .D(1'b0), .SETB(n294), .RSTB(
        sram_rdata_weight[83]), .CLK(clk), .Q(delay_weight[83]) );
  DFFSSRX1_HVT delay_weight_reg_82_ ( .D(1'b0), .SETB(n306), .RSTB(
        sram_rdata_weight[82]), .CLK(clk), .Q(delay_weight[82]) );
  DFFSSRX1_HVT delay_weight_reg_81_ ( .D(1'b0), .SETB(n299), .RSTB(
        sram_rdata_weight[81]), .CLK(clk), .Q(delay_weight[81]) );
  DFFSSRX1_HVT delay_weight_reg_80_ ( .D(1'b0), .SETB(n295), .RSTB(
        sram_rdata_weight[80]), .CLK(clk), .Q(delay_weight[80]) );
  DFFSSRX1_HVT delay_weight_reg_79_ ( .D(1'b0), .SETB(n301), .RSTB(
        sram_rdata_weight[79]), .CLK(clk), .Q(delay_weight[79]) );
  DFFSSRX1_HVT delay_weight_reg_78_ ( .D(1'b0), .SETB(n296), .RSTB(
        sram_rdata_weight[78]), .CLK(clk), .Q(delay_weight[78]) );
  DFFSSRX1_HVT delay_weight_reg_77_ ( .D(1'b0), .SETB(n294), .RSTB(
        sram_rdata_weight[77]), .CLK(clk), .Q(delay_weight[77]) );
  DFFSSRX1_HVT delay_weight_reg_76_ ( .D(1'b0), .SETB(n302), .RSTB(
        sram_rdata_weight[76]), .CLK(clk), .Q(delay_weight[76]) );
  DFFSSRX1_HVT delay_weight_reg_75_ ( .D(1'b0), .SETB(n297), .RSTB(
        sram_rdata_weight[75]), .CLK(clk), .Q(delay_weight[75]) );
  DFFSSRX1_HVT delay_weight_reg_74_ ( .D(1'b0), .SETB(n293), .RSTB(
        sram_rdata_weight[74]), .CLK(clk), .Q(delay_weight[74]) );
  DFFSSRX1_HVT delay_weight_reg_73_ ( .D(1'b0), .SETB(n303), .RSTB(
        sram_rdata_weight[73]), .CLK(clk), .Q(delay_weight[73]) );
  DFFSSRX1_HVT delay_weight_reg_72_ ( .D(1'b0), .SETB(n298), .RSTB(
        sram_rdata_weight[72]), .CLK(clk), .Q(delay_weight[72]) );
  DFFSSRX1_HVT delay_weight_reg_71_ ( .D(1'b0), .SETB(n294), .RSTB(
        sram_rdata_weight[71]), .CLK(clk), .Q(delay_weight[71]) );
  DFFSSRX1_HVT delay_weight_reg_70_ ( .D(1'b0), .SETB(n306), .RSTB(
        sram_rdata_weight[70]), .CLK(clk), .Q(delay_weight[70]) );
  DFFSSRX1_HVT delay_weight_reg_69_ ( .D(1'b0), .SETB(n299), .RSTB(
        sram_rdata_weight[69]), .CLK(clk), .Q(delay_weight[69]) );
  DFFSSRX1_HVT delay_weight_reg_68_ ( .D(1'b0), .SETB(n295), .RSTB(
        sram_rdata_weight[68]), .CLK(clk), .Q(delay_weight[68]) );
  DFFSSRX1_HVT delay_weight_reg_67_ ( .D(1'b0), .SETB(n301), .RSTB(
        sram_rdata_weight[67]), .CLK(clk), .Q(delay_weight[67]) );
  DFFSSRX1_HVT delay_weight_reg_66_ ( .D(1'b0), .SETB(n296), .RSTB(
        sram_rdata_weight[66]), .CLK(clk), .Q(delay_weight[66]) );
  DFFSSRX1_HVT delay_weight_reg_65_ ( .D(1'b0), .SETB(n297), .RSTB(
        sram_rdata_weight[65]), .CLK(clk), .Q(delay_weight[65]) );
  DFFSSRX1_HVT delay_weight_reg_64_ ( .D(1'b0), .SETB(n302), .RSTB(
        sram_rdata_weight[64]), .CLK(clk), .Q(delay_weight[64]) );
  DFFSSRX1_HVT delay_weight_reg_63_ ( .D(1'b0), .SETB(n297), .RSTB(
        sram_rdata_weight[63]), .CLK(clk), .Q(delay_weight[63]) );
  DFFSSRX1_HVT delay_weight_reg_62_ ( .D(1'b0), .SETB(n293), .RSTB(
        sram_rdata_weight[62]), .CLK(clk), .Q(delay_weight[62]) );
  DFFSSRX1_HVT delay_weight_reg_61_ ( .D(1'b0), .SETB(n303), .RSTB(
        sram_rdata_weight[61]), .CLK(clk), .Q(delay_weight[61]) );
  DFFSSRX1_HVT delay_weight_reg_60_ ( .D(1'b0), .SETB(n298), .RSTB(
        sram_rdata_weight[60]), .CLK(clk), .Q(delay_weight[60]) );
  DFFSSRX1_HVT delay_weight_reg_59_ ( .D(1'b0), .SETB(n294), .RSTB(
        sram_rdata_weight[59]), .CLK(clk), .Q(delay_weight[59]) );
  DFFSSRX1_HVT delay_weight_reg_58_ ( .D(1'b0), .SETB(n306), .RSTB(
        sram_rdata_weight[58]), .CLK(clk), .Q(delay_weight[58]) );
  DFFSSRX1_HVT delay_weight_reg_57_ ( .D(1'b0), .SETB(n299), .RSTB(
        sram_rdata_weight[57]), .CLK(clk), .Q(delay_weight[57]) );
  DFFSSRX1_HVT delay_weight_reg_56_ ( .D(1'b0), .SETB(n295), .RSTB(
        sram_rdata_weight[56]), .CLK(clk), .Q(delay_weight[56]) );
  DFFSSRX1_HVT delay_weight_reg_55_ ( .D(1'b0), .SETB(n301), .RSTB(
        sram_rdata_weight[55]), .CLK(clk), .Q(delay_weight[55]) );
  DFFSSRX1_HVT delay_weight_reg_54_ ( .D(1'b0), .SETB(n296), .RSTB(
        sram_rdata_weight[54]), .CLK(clk), .Q(delay_weight[54]) );
  DFFSSRX1_HVT delay_weight_reg_53_ ( .D(1'b0), .SETB(n293), .RSTB(
        sram_rdata_weight[53]), .CLK(clk), .Q(delay_weight[53]) );
  DFFSSRX1_HVT delay_weight_reg_52_ ( .D(1'b0), .SETB(n302), .RSTB(
        sram_rdata_weight[52]), .CLK(clk), .Q(delay_weight[52]) );
  DFFSSRX1_HVT delay_weight_reg_51_ ( .D(1'b0), .SETB(n297), .RSTB(
        sram_rdata_weight[51]), .CLK(clk), .Q(delay_weight[51]) );
  DFFSSRX1_HVT delay_weight_reg_50_ ( .D(1'b0), .SETB(n293), .RSTB(
        sram_rdata_weight[50]), .CLK(clk), .Q(delay_weight[50]) );
  DFFSSRX1_HVT delay_weight_reg_49_ ( .D(1'b0), .SETB(n303), .RSTB(
        sram_rdata_weight[49]), .CLK(clk), .Q(delay_weight[49]) );
  DFFSSRX1_HVT delay_weight_reg_48_ ( .D(1'b0), .SETB(n298), .RSTB(
        sram_rdata_weight[48]), .CLK(clk), .Q(delay_weight[48]) );
  DFFSSRX1_HVT delay_weight_reg_47_ ( .D(1'b0), .SETB(n294), .RSTB(
        sram_rdata_weight[47]), .CLK(clk), .Q(delay_weight[47]) );
  DFFSSRX1_HVT delay_weight_reg_46_ ( .D(1'b0), .SETB(n306), .RSTB(
        sram_rdata_weight[46]), .CLK(clk), .Q(delay_weight[46]) );
  DFFSSRX1_HVT delay_weight_reg_45_ ( .D(1'b0), .SETB(n299), .RSTB(
        sram_rdata_weight[45]), .CLK(clk), .Q(delay_weight[45]) );
  DFFSSRX1_HVT delay_weight_reg_44_ ( .D(1'b0), .SETB(n295), .RSTB(
        sram_rdata_weight[44]), .CLK(clk), .Q(delay_weight[44]) );
  DFFSSRX1_HVT delay_weight_reg_43_ ( .D(1'b0), .SETB(n301), .RSTB(
        sram_rdata_weight[43]), .CLK(clk), .Q(delay_weight[43]) );
  DFFSSRX1_HVT delay_weight_reg_42_ ( .D(1'b0), .SETB(n296), .RSTB(
        sram_rdata_weight[42]), .CLK(clk), .Q(delay_weight[42]) );
  DFFSSRX1_HVT delay_weight_reg_41_ ( .D(1'b0), .SETB(n295), .RSTB(
        sram_rdata_weight[41]), .CLK(clk), .Q(delay_weight[41]) );
  DFFSSRX1_HVT delay_weight_reg_40_ ( .D(1'b0), .SETB(n302), .RSTB(
        sram_rdata_weight[40]), .CLK(clk), .Q(delay_weight[40]) );
  DFFSSRX1_HVT delay_weight_reg_39_ ( .D(1'b0), .SETB(n297), .RSTB(
        sram_rdata_weight[39]), .CLK(clk), .Q(delay_weight[39]) );
  DFFSSRX1_HVT delay_weight_reg_38_ ( .D(1'b0), .SETB(n293), .RSTB(
        sram_rdata_weight[38]), .CLK(clk), .Q(delay_weight[38]) );
  DFFSSRX1_HVT delay_weight_reg_37_ ( .D(1'b0), .SETB(n303), .RSTB(
        sram_rdata_weight[37]), .CLK(clk), .Q(delay_weight[37]) );
  DFFSSRX1_HVT delay_weight_reg_36_ ( .D(1'b0), .SETB(n298), .RSTB(
        sram_rdata_weight[36]), .CLK(clk), .Q(delay_weight[36]) );
  DFFSSRX1_HVT delay_weight_reg_35_ ( .D(1'b0), .SETB(n294), .RSTB(
        sram_rdata_weight[35]), .CLK(clk), .Q(delay_weight[35]) );
  DFFSSRX1_HVT delay_weight_reg_34_ ( .D(1'b0), .SETB(n306), .RSTB(
        sram_rdata_weight[34]), .CLK(clk), .Q(delay_weight[34]) );
  DFFSSRX1_HVT delay_weight_reg_33_ ( .D(1'b0), .SETB(n299), .RSTB(
        sram_rdata_weight[33]), .CLK(clk), .Q(delay_weight[33]) );
  DFFSSRX1_HVT delay_weight_reg_32_ ( .D(1'b0), .SETB(n295), .RSTB(
        sram_rdata_weight[32]), .CLK(clk), .Q(delay_weight[32]) );
  DFFSSRX1_HVT delay_weight_reg_31_ ( .D(1'b0), .SETB(n301), .RSTB(
        sram_rdata_weight[31]), .CLK(clk), .Q(delay_weight[31]) );
  DFFSSRX1_HVT delay_weight_reg_30_ ( .D(1'b0), .SETB(n296), .RSTB(
        sram_rdata_weight[30]), .CLK(clk), .Q(delay_weight[30]) );
  DFFSSRX1_HVT delay_weight_reg_29_ ( .D(1'b0), .SETB(n294), .RSTB(
        sram_rdata_weight[29]), .CLK(clk), .Q(delay_weight[29]) );
  DFFSSRX1_HVT delay_weight_reg_28_ ( .D(1'b0), .SETB(n302), .RSTB(
        sram_rdata_weight[28]), .CLK(clk), .Q(delay_weight[28]) );
  DFFSSRX1_HVT delay_weight_reg_27_ ( .D(1'b0), .SETB(n297), .RSTB(
        sram_rdata_weight[27]), .CLK(clk), .Q(delay_weight[27]) );
  DFFSSRX1_HVT delay_weight_reg_26_ ( .D(1'b0), .SETB(n293), .RSTB(
        sram_rdata_weight[26]), .CLK(clk), .Q(delay_weight[26]) );
  DFFSSRX1_HVT delay_weight_reg_25_ ( .D(1'b0), .SETB(n303), .RSTB(
        sram_rdata_weight[25]), .CLK(clk), .Q(delay_weight[25]) );
  DFFSSRX1_HVT delay_weight_reg_24_ ( .D(1'b0), .SETB(n298), .RSTB(
        sram_rdata_weight[24]), .CLK(clk), .Q(delay_weight[24]) );
  DFFSSRX1_HVT delay_weight_reg_23_ ( .D(1'b0), .SETB(n294), .RSTB(
        sram_rdata_weight[23]), .CLK(clk), .Q(delay_weight[23]) );
  DFFSSRX1_HVT delay_weight_reg_22_ ( .D(1'b0), .SETB(n306), .RSTB(
        sram_rdata_weight[22]), .CLK(clk), .Q(delay_weight[22]) );
  DFFSSRX1_HVT delay_weight_reg_21_ ( .D(1'b0), .SETB(n299), .RSTB(
        sram_rdata_weight[21]), .CLK(clk), .Q(delay_weight[21]) );
  DFFSSRX1_HVT delay_weight_reg_20_ ( .D(1'b0), .SETB(n295), .RSTB(
        sram_rdata_weight[20]), .CLK(clk), .Q(delay_weight[20]) );
  DFFSSRX1_HVT delay_weight_reg_19_ ( .D(1'b0), .SETB(n301), .RSTB(
        sram_rdata_weight[19]), .CLK(clk), .Q(delay_weight[19]) );
  DFFSSRX1_HVT delay_weight_reg_18_ ( .D(1'b0), .SETB(n296), .RSTB(
        sram_rdata_weight[18]), .CLK(clk), .Q(delay_weight[18]) );
  DFFSSRX1_HVT delay_weight_reg_17_ ( .D(1'b0), .SETB(n298), .RSTB(
        sram_rdata_weight[17]), .CLK(clk), .Q(delay_weight[17]) );
  DFFSSRX1_HVT delay_weight_reg_16_ ( .D(1'b0), .SETB(n302), .RSTB(
        sram_rdata_weight[16]), .CLK(clk), .Q(delay_weight[16]) );
  DFFSSRX1_HVT delay_weight_reg_15_ ( .D(1'b0), .SETB(n297), .RSTB(
        sram_rdata_weight[15]), .CLK(clk), .Q(delay_weight[15]) );
  DFFSSRX1_HVT delay_weight_reg_14_ ( .D(1'b0), .SETB(n293), .RSTB(
        sram_rdata_weight[14]), .CLK(clk), .Q(delay_weight[14]) );
  DFFSSRX1_HVT delay_weight_reg_13_ ( .D(1'b0), .SETB(n303), .RSTB(
        sram_rdata_weight[13]), .CLK(clk), .Q(delay_weight[13]) );
  DFFSSRX1_HVT delay_weight_reg_12_ ( .D(1'b0), .SETB(n298), .RSTB(
        sram_rdata_weight[12]), .CLK(clk), .Q(delay_weight[12]) );
  DFFSSRX1_HVT delay_weight_reg_11_ ( .D(1'b0), .SETB(n294), .RSTB(
        sram_rdata_weight[11]), .CLK(clk), .Q(delay_weight[11]) );
  DFFSSRX1_HVT delay_weight_reg_10_ ( .D(1'b0), .SETB(n306), .RSTB(
        sram_rdata_weight[10]), .CLK(clk), .Q(delay_weight[10]) );
  DFFSSRX1_HVT delay_weight_reg_9_ ( .D(1'b0), .SETB(n299), .RSTB(
        sram_rdata_weight[9]), .CLK(clk), .Q(delay_weight[9]) );
  DFFSSRX1_HVT delay_weight_reg_8_ ( .D(1'b0), .SETB(n295), .RSTB(
        sram_rdata_weight[8]), .CLK(clk), .Q(delay_weight[8]) );
  DFFSSRX1_HVT delay_weight_reg_7_ ( .D(1'b0), .SETB(n301), .RSTB(
        sram_rdata_weight[7]), .CLK(clk), .Q(delay_weight[7]) );
  DFFSSRX1_HVT delay_weight_reg_6_ ( .D(1'b0), .SETB(n296), .RSTB(
        sram_rdata_weight[6]), .CLK(clk), .Q(delay_weight[6]) );
  DFFSSRX1_HVT delay_weight_reg_5_ ( .D(1'b0), .SETB(n298), .RSTB(
        sram_rdata_weight[5]), .CLK(clk), .Q(delay_weight[5]) );
  DFFSSRX1_HVT delay_weight_reg_4_ ( .D(1'b0), .SETB(n302), .RSTB(
        sram_rdata_weight[4]), .CLK(clk), .Q(delay_weight[4]) );
  DFFSSRX1_HVT delay_weight_reg_3_ ( .D(1'b0), .SETB(n297), .RSTB(
        sram_rdata_weight[3]), .CLK(clk), .Q(delay_weight[3]) );
  DFFSSRX1_HVT delay_weight_reg_2_ ( .D(1'b0), .SETB(n293), .RSTB(
        sram_rdata_weight[2]), .CLK(clk), .Q(delay_weight[2]) );
  DFFSSRX1_HVT delay_weight_reg_1_ ( .D(1'b0), .SETB(n303), .RSTB(
        sram_rdata_weight[1]), .CLK(clk), .Q(delay_weight[1]) );
  DFFSSRX1_HVT delay_weight_reg_0_ ( .D(1'b0), .SETB(n302), .RSTB(
        sram_rdata_weight[0]), .CLK(clk), .Q(delay_weight[0]) );
  DFFSSRX1_HVT conv_weight_box_reg_0__3_ ( .D(1'b0), .SETB(n303), .RSTB(
        net19121), .CLK(net19135), .Q(conv_weight_box[199]) );
  DFFSSRX1_HVT conv_weight_box_reg_0__2_ ( .D(1'b0), .SETB(n293), .RSTB(
        net19124), .CLK(net19135), .Q(conv_weight_box[198]) );
  DFFSSRX1_HVT conv_weight_box_reg_0__1_ ( .D(1'b0), .SETB(n297), .RSTB(
        net19125), .CLK(net19135), .Q(conv_weight_box[197]) );
  DFFSSRX1_HVT conv_weight_box_reg_0__0_ ( .D(1'b0), .SETB(n302), .RSTB(
        net19126), .CLK(net19135), .Q(conv_weight_box[196]) );
  DFFSSRX1_HVT conv_weight_box_reg_1__3_ ( .D(1'b0), .SETB(n305), .RSTB(
        net19127), .CLK(net19135), .Q(conv_weight_box[195]) );
  DFFSSRX1_HVT conv_weight_box_reg_1__2_ ( .D(1'b0), .SETB(n296), .RSTB(
        net19128), .CLK(net19135), .Q(conv_weight_box[194]) );
  DFFSSRX1_HVT conv_weight_box_reg_1__1_ ( .D(1'b0), .SETB(n301), .RSTB(
        net19129), .CLK(net19135), .Q(conv_weight_box[193]) );
  DFFSSRX1_HVT conv_weight_box_reg_1__0_ ( .D(1'b0), .SETB(n295), .RSTB(
        net19130), .CLK(net19135), .Q(conv_weight_box[192]) );
  DFFSSRX1_HVT conv_weight_box_reg_2__3_ ( .D(1'b0), .SETB(n299), .RSTB(
        net19131), .CLK(net19135), .Q(conv_weight_box[191]) );
  DFFSSRX1_HVT conv_weight_box_reg_2__2_ ( .D(1'b0), .SETB(n306), .RSTB(
        net19132), .CLK(net19135), .Q(conv_weight_box[190]) );
  DFFSSRX1_HVT conv_weight_box_reg_2__1_ ( .D(1'b0), .SETB(n294), .RSTB(
        net19140), .CLK(net19152), .Q(conv_weight_box[189]) );
  DFFSSRX1_HVT conv_weight_box_reg_2__0_ ( .D(1'b0), .SETB(n298), .RSTB(
        net19141), .CLK(net19152), .Q(conv_weight_box[188]) );
  DFFSSRX1_HVT conv_weight_box_reg_3__3_ ( .D(1'b0), .SETB(n303), .RSTB(
        net19142), .CLK(net19152), .Q(conv_weight_box[187]) );
  DFFSSRX1_HVT conv_weight_box_reg_3__2_ ( .D(1'b0), .SETB(n293), .RSTB(
        net19143), .CLK(net19152), .Q(conv_weight_box[186]) );
  DFFSSRX1_HVT conv_weight_box_reg_3__1_ ( .D(1'b0), .SETB(n297), .RSTB(
        net19144), .CLK(net19152), .Q(conv_weight_box[185]) );
  DFFSSRX1_HVT conv_weight_box_reg_3__0_ ( .D(1'b0), .SETB(n302), .RSTB(
        net19145), .CLK(net19152), .Q(conv_weight_box[184]) );
  DFFSSRX1_HVT conv_weight_box_reg_4__3_ ( .D(1'b0), .SETB(n305), .RSTB(
        net19146), .CLK(net19152), .Q(conv_weight_box[183]) );
  DFFSSRX1_HVT conv_weight_box_reg_4__2_ ( .D(1'b0), .SETB(n296), .RSTB(
        net19147), .CLK(net19152), .Q(conv_weight_box[182]) );
  DFFSSRX1_HVT conv_weight_box_reg_4__1_ ( .D(1'b0), .SETB(n301), .RSTB(
        net19148), .CLK(net19152), .Q(conv_weight_box[181]) );
  DFFSSRX1_HVT conv_weight_box_reg_4__0_ ( .D(1'b0), .SETB(n295), .RSTB(
        net19149), .CLK(net19152), .Q(conv_weight_box[180]) );
  DFFSSRX1_HVT conv_weight_box_reg_5__3_ ( .D(1'b0), .SETB(n299), .RSTB(
        net19157), .CLK(net19169), .Q(conv_weight_box[179]) );
  DFFSSRX1_HVT conv_weight_box_reg_5__2_ ( .D(1'b0), .SETB(n306), .RSTB(
        net19158), .CLK(net19169), .Q(conv_weight_box[178]) );
  DFFSSRX1_HVT conv_weight_box_reg_5__1_ ( .D(1'b0), .SETB(n294), .RSTB(
        net19159), .CLK(net19169), .Q(conv_weight_box[177]) );
  DFFSSRX1_HVT conv_weight_box_reg_5__0_ ( .D(1'b0), .SETB(n298), .RSTB(
        net19160), .CLK(net19169), .Q(conv_weight_box[176]) );
  DFFSSRX1_HVT conv_weight_box_reg_6__3_ ( .D(1'b0), .SETB(n303), .RSTB(
        net19161), .CLK(net19169), .Q(conv_weight_box[175]) );
  DFFSSRX1_HVT conv_weight_box_reg_6__2_ ( .D(1'b0), .SETB(n293), .RSTB(
        net19162), .CLK(net19169), .Q(conv_weight_box[174]) );
  DFFSSRX1_HVT conv_weight_box_reg_6__1_ ( .D(1'b0), .SETB(n297), .RSTB(
        net19163), .CLK(net19169), .Q(conv_weight_box[173]) );
  DFFSSRX1_HVT conv_weight_box_reg_6__0_ ( .D(1'b0), .SETB(n302), .RSTB(
        net19164), .CLK(net19169), .Q(conv_weight_box[172]) );
  DFFSSRX1_HVT conv_weight_box_reg_7__3_ ( .D(1'b0), .SETB(n305), .RSTB(
        net19165), .CLK(net19169), .Q(conv_weight_box[171]) );
  DFFSSRX1_HVT conv_weight_box_reg_7__2_ ( .D(1'b0), .SETB(n296), .RSTB(
        net19166), .CLK(net19169), .Q(conv_weight_box[170]) );
  DFFSSRX1_HVT conv_weight_box_reg_7__1_ ( .D(1'b0), .SETB(n301), .RSTB(
        net19174), .CLK(net19186), .Q(conv_weight_box[169]) );
  DFFSSRX1_HVT conv_weight_box_reg_7__0_ ( .D(1'b0), .SETB(n295), .RSTB(
        net19175), .CLK(net19186), .Q(conv_weight_box[168]) );
  DFFSSRX1_HVT conv_weight_box_reg_8__3_ ( .D(1'b0), .SETB(n299), .RSTB(
        net19176), .CLK(net19186), .Q(conv_weight_box[167]) );
  DFFSSRX1_HVT conv_weight_box_reg_8__2_ ( .D(1'b0), .SETB(n306), .RSTB(
        net19177), .CLK(net19186), .Q(conv_weight_box[166]) );
  DFFSSRX1_HVT conv_weight_box_reg_8__1_ ( .D(1'b0), .SETB(n294), .RSTB(
        net19178), .CLK(net19186), .Q(conv_weight_box[165]) );
  DFFSSRX1_HVT conv_weight_box_reg_8__0_ ( .D(1'b0), .SETB(n298), .RSTB(
        net19179), .CLK(net19186), .Q(conv_weight_box[164]) );
  DFFSSRX1_HVT conv_weight_box_reg_9__3_ ( .D(1'b0), .SETB(n303), .RSTB(
        net19180), .CLK(net19186), .Q(conv_weight_box[163]) );
  DFFSSRX1_HVT conv_weight_box_reg_9__2_ ( .D(1'b0), .SETB(n293), .RSTB(
        net19181), .CLK(net19186), .Q(conv_weight_box[162]) );
  DFFSSRX1_HVT conv_weight_box_reg_9__1_ ( .D(1'b0), .SETB(n297), .RSTB(
        net19182), .CLK(net19186), .Q(conv_weight_box[161]) );
  DFFSSRX1_HVT conv_weight_box_reg_9__0_ ( .D(1'b0), .SETB(n302), .RSTB(
        net19183), .CLK(net19186), .Q(conv_weight_box[160]) );
  DFFSSRX1_HVT conv_weight_box_reg_10__3_ ( .D(1'b0), .SETB(n305), .RSTB(
        net19191), .CLK(net19203), .Q(conv_weight_box[159]) );
  DFFSSRX1_HVT conv_weight_box_reg_10__2_ ( .D(1'b0), .SETB(n296), .RSTB(
        net19192), .CLK(net19203), .Q(conv_weight_box[158]) );
  DFFSSRX1_HVT conv_weight_box_reg_10__1_ ( .D(1'b0), .SETB(n301), .RSTB(
        net19193), .CLK(net19203), .Q(conv_weight_box[157]) );
  DFFSSRX1_HVT conv_weight_box_reg_10__0_ ( .D(1'b0), .SETB(n295), .RSTB(
        net19194), .CLK(net19203), .Q(conv_weight_box[156]) );
  DFFSSRX1_HVT conv_weight_box_reg_11__3_ ( .D(1'b0), .SETB(n299), .RSTB(
        net19195), .CLK(net19203), .Q(conv_weight_box[155]) );
  DFFSSRX1_HVT conv_weight_box_reg_11__2_ ( .D(1'b0), .SETB(n306), .RSTB(
        net19196), .CLK(net19203), .Q(conv_weight_box[154]) );
  DFFSSRX1_HVT conv_weight_box_reg_11__1_ ( .D(1'b0), .SETB(n294), .RSTB(
        net19197), .CLK(net19203), .Q(conv_weight_box[153]) );
  DFFSSRX1_HVT conv_weight_box_reg_11__0_ ( .D(1'b0), .SETB(n298), .RSTB(
        net19198), .CLK(net19203), .Q(conv_weight_box[152]) );
  DFFSSRX1_HVT conv_weight_box_reg_12__3_ ( .D(1'b0), .SETB(n303), .RSTB(
        net19199), .CLK(net19203), .Q(conv_weight_box[151]) );
  DFFSSRX1_HVT conv_weight_box_reg_12__2_ ( .D(1'b0), .SETB(n293), .RSTB(
        net19200), .CLK(net19203), .Q(conv_weight_box[150]) );
  DFFSSRX1_HVT conv_weight_box_reg_12__1_ ( .D(1'b0), .SETB(n297), .RSTB(
        net19208), .CLK(net19220), .Q(conv_weight_box[149]) );
  DFFSSRX1_HVT conv_weight_box_reg_12__0_ ( .D(1'b0), .SETB(n302), .RSTB(
        net19209), .CLK(net19220), .Q(conv_weight_box[148]) );
  DFFSSRX1_HVT conv_weight_box_reg_13__3_ ( .D(1'b0), .SETB(n305), .RSTB(
        net19210), .CLK(net19220), .Q(conv_weight_box[147]) );
  DFFSSRX1_HVT conv_weight_box_reg_13__2_ ( .D(1'b0), .SETB(n296), .RSTB(
        net19211), .CLK(net19220), .Q(conv_weight_box[146]) );
  DFFSSRX1_HVT conv_weight_box_reg_13__1_ ( .D(1'b0), .SETB(n301), .RSTB(
        net19212), .CLK(net19220), .Q(conv_weight_box[145]) );
  DFFSSRX1_HVT conv_weight_box_reg_13__0_ ( .D(1'b0), .SETB(n295), .RSTB(
        net19213), .CLK(net19220), .Q(conv_weight_box[144]) );
  DFFSSRX1_HVT conv_weight_box_reg_14__3_ ( .D(1'b0), .SETB(n299), .RSTB(
        net19214), .CLK(net19220), .Q(conv_weight_box[143]) );
  DFFSSRX1_HVT conv_weight_box_reg_14__2_ ( .D(1'b0), .SETB(n306), .RSTB(
        net19215), .CLK(net19220), .Q(conv_weight_box[142]) );
  DFFSSRX1_HVT conv_weight_box_reg_14__1_ ( .D(1'b0), .SETB(n294), .RSTB(
        net19216), .CLK(net19220), .Q(conv_weight_box[141]) );
  DFFSSRX1_HVT conv_weight_box_reg_14__0_ ( .D(1'b0), .SETB(n298), .RSTB(
        net19217), .CLK(net19220), .Q(conv_weight_box[140]) );
  DFFSSRX1_HVT conv_weight_box_reg_15__3_ ( .D(1'b0), .SETB(n303), .RSTB(
        net19225), .CLK(net19237), .Q(conv_weight_box[139]) );
  DFFSSRX1_HVT conv_weight_box_reg_15__2_ ( .D(1'b0), .SETB(n293), .RSTB(
        net19226), .CLK(net19237), .Q(conv_weight_box[138]) );
  DFFSSRX1_HVT conv_weight_box_reg_15__1_ ( .D(1'b0), .SETB(n297), .RSTB(
        net19227), .CLK(net19237), .Q(conv_weight_box[137]) );
  DFFSSRX1_HVT conv_weight_box_reg_15__0_ ( .D(1'b0), .SETB(n302), .RSTB(
        net19228), .CLK(net19237), .Q(conv_weight_box[136]) );
  DFFSSRX1_HVT conv_weight_box_reg_16__3_ ( .D(1'b0), .SETB(n305), .RSTB(
        net19229), .CLK(net19237), .Q(conv_weight_box[135]) );
  DFFSSRX1_HVT conv_weight_box_reg_16__2_ ( .D(1'b0), .SETB(n296), .RSTB(
        net19230), .CLK(net19237), .Q(conv_weight_box[134]) );
  DFFSSRX1_HVT conv_weight_box_reg_16__1_ ( .D(1'b0), .SETB(n301), .RSTB(
        net19231), .CLK(net19237), .Q(conv_weight_box[133]) );
  DFFSSRX1_HVT conv_weight_box_reg_16__0_ ( .D(1'b0), .SETB(n295), .RSTB(
        net19232), .CLK(net19237), .Q(conv_weight_box[132]) );
  DFFSSRX1_HVT conv_weight_box_reg_17__3_ ( .D(1'b0), .SETB(n299), .RSTB(
        net19233), .CLK(net19237), .Q(conv_weight_box[131]) );
  DFFSSRX1_HVT conv_weight_box_reg_17__2_ ( .D(1'b0), .SETB(n306), .RSTB(
        net19234), .CLK(net19237), .Q(conv_weight_box[130]) );
  DFFSSRX1_HVT conv_weight_box_reg_17__1_ ( .D(1'b0), .SETB(n294), .RSTB(
        net19242), .CLK(net19254), .Q(conv_weight_box[129]) );
  DFFSSRX1_HVT conv_weight_box_reg_17__0_ ( .D(1'b0), .SETB(n298), .RSTB(
        net19243), .CLK(net19254), .Q(conv_weight_box[128]) );
  DFFSSRX1_HVT conv_weight_box_reg_18__3_ ( .D(1'b0), .SETB(n303), .RSTB(
        net19244), .CLK(net19254), .Q(conv_weight_box[127]) );
  DFFSSRX1_HVT conv_weight_box_reg_18__2_ ( .D(1'b0), .SETB(n293), .RSTB(
        net19245), .CLK(net19254), .Q(conv_weight_box[126]) );
  DFFSSRX1_HVT conv_weight_box_reg_18__1_ ( .D(1'b0), .SETB(n297), .RSTB(
        net19246), .CLK(net19254), .Q(conv_weight_box[125]) );
  DFFSSRX1_HVT conv_weight_box_reg_18__0_ ( .D(1'b0), .SETB(n302), .RSTB(
        net19247), .CLK(net19254), .Q(conv_weight_box[124]) );
  DFFSSRX1_HVT conv_weight_box_reg_19__3_ ( .D(1'b0), .SETB(n305), .RSTB(
        net19248), .CLK(net19254), .Q(conv_weight_box[123]) );
  DFFSSRX1_HVT conv_weight_box_reg_19__2_ ( .D(1'b0), .SETB(n296), .RSTB(
        net19249), .CLK(net19254), .Q(conv_weight_box[122]) );
  DFFSSRX1_HVT conv_weight_box_reg_19__1_ ( .D(1'b0), .SETB(n301), .RSTB(
        net19250), .CLK(net19254), .Q(conv_weight_box[121]) );
  DFFSSRX1_HVT conv_weight_box_reg_19__0_ ( .D(1'b0), .SETB(n295), .RSTB(
        net19251), .CLK(net19254), .Q(conv_weight_box[120]) );
  DFFSSRX1_HVT conv_weight_box_reg_20__3_ ( .D(1'b0), .SETB(n299), .RSTB(
        net19259), .CLK(net19271), .Q(conv_weight_box[119]) );
  DFFSSRX1_HVT conv_weight_box_reg_20__2_ ( .D(1'b0), .SETB(n306), .RSTB(
        net19260), .CLK(net19271), .Q(conv_weight_box[118]) );
  DFFSSRX1_HVT conv_weight_box_reg_20__1_ ( .D(1'b0), .SETB(n294), .RSTB(
        net19261), .CLK(net19271), .Q(conv_weight_box[117]) );
  DFFSSRX1_HVT conv_weight_box_reg_20__0_ ( .D(1'b0), .SETB(n298), .RSTB(
        net19262), .CLK(net19271), .Q(conv_weight_box[116]) );
  DFFSSRX1_HVT conv_weight_box_reg_21__3_ ( .D(1'b0), .SETB(n303), .RSTB(
        net19263), .CLK(net19271), .Q(conv_weight_box[115]) );
  DFFSSRX1_HVT conv_weight_box_reg_21__2_ ( .D(1'b0), .SETB(n293), .RSTB(
        net19264), .CLK(net19271), .Q(conv_weight_box[114]) );
  DFFSSRX1_HVT conv_weight_box_reg_21__1_ ( .D(1'b0), .SETB(n297), .RSTB(
        net19265), .CLK(net19271), .Q(conv_weight_box[113]) );
  DFFSSRX1_HVT conv_weight_box_reg_21__0_ ( .D(1'b0), .SETB(n302), .RSTB(
        net19266), .CLK(net19271), .Q(conv_weight_box[112]) );
  DFFSSRX1_HVT conv_weight_box_reg_22__3_ ( .D(1'b0), .SETB(n301), .RSTB(
        net19267), .CLK(net19271), .Q(conv_weight_box[111]) );
  DFFSSRX1_HVT conv_weight_box_reg_22__2_ ( .D(1'b0), .SETB(n296), .RSTB(
        net19268), .CLK(net19271), .Q(conv_weight_box[110]) );
  DFFSSRX1_HVT conv_weight_box_reg_22__1_ ( .D(1'b0), .SETB(n301), .RSTB(
        net19276), .CLK(net19288), .Q(conv_weight_box[109]) );
  DFFSSRX1_HVT conv_weight_box_reg_22__0_ ( .D(1'b0), .SETB(n295), .RSTB(
        net19277), .CLK(net19288), .Q(conv_weight_box[108]) );
  DFFSSRX1_HVT conv_weight_box_reg_23__3_ ( .D(1'b0), .SETB(n299), .RSTB(
        net19278), .CLK(net19288), .Q(conv_weight_box[107]) );
  DFFSSRX1_HVT conv_weight_box_reg_23__2_ ( .D(1'b0), .SETB(n306), .RSTB(
        net19279), .CLK(net19288), .Q(conv_weight_box[106]) );
  DFFSSRX1_HVT conv_weight_box_reg_23__1_ ( .D(1'b0), .SETB(n294), .RSTB(
        net19280), .CLK(net19288), .Q(conv_weight_box[105]) );
  DFFSSRX1_HVT conv_weight_box_reg_23__0_ ( .D(1'b0), .SETB(n298), .RSTB(
        net19281), .CLK(net19288), .Q(conv_weight_box[104]) );
  DFFSSRX1_HVT conv_weight_box_reg_24__3_ ( .D(1'b0), .SETB(n303), .RSTB(
        net19282), .CLK(net19288), .Q(conv_weight_box[103]) );
  DFFSSRX1_HVT conv_weight_box_reg_24__2_ ( .D(1'b0), .SETB(n293), .RSTB(
        net19283), .CLK(net19288), .Q(conv_weight_box[102]) );
  DFFSSRX1_HVT conv_weight_box_reg_24__1_ ( .D(1'b0), .SETB(n297), .RSTB(
        net19284), .CLK(net19288), .Q(conv_weight_box[101]) );
  DFFSSRX1_HVT conv_weight_box_reg_24__0_ ( .D(1'b0), .SETB(n302), .RSTB(
        net19285), .CLK(net19288), .Q(conv_weight_box[100]) );
  DFFSSRX1_HVT conv_weight_box_reg_25__3_ ( .D(1'b0), .SETB(n306), .RSTB(
        net19301), .CLK(net19313), .Q(conv_weight_box[99]) );
  DFFSSRX1_HVT conv_weight_box_reg_25__2_ ( .D(1'b0), .SETB(n296), .RSTB(
        net19302), .CLK(net19313), .Q(conv_weight_box[98]) );
  DFFSSRX1_HVT conv_weight_box_reg_25__1_ ( .D(1'b0), .SETB(n301), .RSTB(
        net19303), .CLK(net19313), .Q(conv_weight_box[97]) );
  DFFSSRX1_HVT conv_weight_box_reg_25__0_ ( .D(1'b0), .SETB(n295), .RSTB(
        net19304), .CLK(net19313), .Q(conv_weight_box[96]) );
  DFFSSRX1_HVT conv_weight_box_reg_26__3_ ( .D(1'b0), .SETB(n299), .RSTB(
        net19305), .CLK(net19313), .Q(conv_weight_box[95]) );
  DFFSSRX1_HVT conv_weight_box_reg_26__2_ ( .D(1'b0), .SETB(n306), .RSTB(
        net19306), .CLK(net19313), .Q(conv_weight_box[94]) );
  DFFSSRX1_HVT conv_weight_box_reg_26__1_ ( .D(1'b0), .SETB(n294), .RSTB(
        net19307), .CLK(net19313), .Q(conv_weight_box[93]) );
  DFFSSRX1_HVT conv_weight_box_reg_26__0_ ( .D(1'b0), .SETB(n298), .RSTB(
        net19308), .CLK(net19313), .Q(conv_weight_box[92]) );
  DFFSSRX1_HVT conv_weight_box_reg_27__3_ ( .D(1'b0), .SETB(n303), .RSTB(
        net19309), .CLK(net19313), .Q(conv_weight_box[91]) );
  DFFSSRX1_HVT conv_weight_box_reg_27__2_ ( .D(1'b0), .SETB(n293), .RSTB(
        net19310), .CLK(net19313), .Q(conv_weight_box[90]) );
  DFFSSRX1_HVT conv_weight_box_reg_27__1_ ( .D(1'b0), .SETB(n297), .RSTB(
        net19318), .CLK(net19330), .Q(conv_weight_box[89]) );
  DFFSSRX1_HVT conv_weight_box_reg_27__0_ ( .D(1'b0), .SETB(n302), .RSTB(
        net19319), .CLK(net19330), .Q(conv_weight_box[88]) );
  DFFSSRX1_HVT conv_weight_box_reg_28__3_ ( .D(1'b0), .SETB(n296), .RSTB(
        net19320), .CLK(net19330), .Q(conv_weight_box[87]) );
  DFFSSRX1_HVT conv_weight_box_reg_28__2_ ( .D(1'b0), .SETB(n296), .RSTB(
        net19321), .CLK(net19330), .Q(conv_weight_box[86]) );
  DFFSSRX1_HVT conv_weight_box_reg_28__1_ ( .D(1'b0), .SETB(n301), .RSTB(
        net19322), .CLK(net19330), .Q(conv_weight_box[85]) );
  DFFSSRX1_HVT conv_weight_box_reg_28__0_ ( .D(1'b0), .SETB(n295), .RSTB(
        net19323), .CLK(net19330), .Q(conv_weight_box[84]) );
  DFFSSRX1_HVT conv_weight_box_reg_29__3_ ( .D(1'b0), .SETB(n299), .RSTB(
        net19324), .CLK(net19330), .Q(conv_weight_box[83]) );
  DFFSSRX1_HVT conv_weight_box_reg_29__2_ ( .D(1'b0), .SETB(n306), .RSTB(
        net19325), .CLK(net19330), .Q(conv_weight_box[82]) );
  DFFSSRX1_HVT conv_weight_box_reg_29__1_ ( .D(1'b0), .SETB(n294), .RSTB(
        net19326), .CLK(net19330), .Q(conv_weight_box[81]) );
  DFFSSRX1_HVT conv_weight_box_reg_29__0_ ( .D(1'b0), .SETB(n298), .RSTB(
        net19327), .CLK(net19330), .Q(conv_weight_box[80]) );
  DFFSSRX1_HVT conv_weight_box_reg_30__3_ ( .D(1'b0), .SETB(n303), .RSTB(
        net19335), .CLK(net19347), .Q(conv_weight_box[79]) );
  DFFSSRX1_HVT conv_weight_box_reg_30__2_ ( .D(1'b0), .SETB(n293), .RSTB(
        net19336), .CLK(net19347), .Q(conv_weight_box[78]) );
  DFFSSRX1_HVT conv_weight_box_reg_30__1_ ( .D(1'b0), .SETB(n297), .RSTB(
        net19337), .CLK(net19347), .Q(conv_weight_box[77]) );
  DFFSSRX1_HVT conv_weight_box_reg_30__0_ ( .D(1'b0), .SETB(n302), .RSTB(
        net19338), .CLK(net19347), .Q(conv_weight_box[76]) );
  DFFSSRX1_HVT conv_weight_box_reg_31__3_ ( .D(1'b0), .SETB(n299), .RSTB(
        net19339), .CLK(net19347), .Q(conv_weight_box[75]) );
  DFFSSRX1_HVT conv_weight_box_reg_31__2_ ( .D(1'b0), .SETB(n296), .RSTB(
        net19340), .CLK(net19347), .Q(conv_weight_box[74]) );
  DFFSSRX1_HVT conv_weight_box_reg_31__1_ ( .D(1'b0), .SETB(n301), .RSTB(
        net19341), .CLK(net19347), .Q(conv_weight_box[73]) );
  DFFSSRX1_HVT conv_weight_box_reg_31__0_ ( .D(1'b0), .SETB(n295), .RSTB(
        net19342), .CLK(net19347), .Q(conv_weight_box[72]) );
  DFFSSRX1_HVT conv_weight_box_reg_32__3_ ( .D(1'b0), .SETB(n299), .RSTB(
        net19343), .CLK(net19347), .Q(conv_weight_box[71]) );
  DFFSSRX1_HVT conv_weight_box_reg_32__2_ ( .D(1'b0), .SETB(n306), .RSTB(
        net19344), .CLK(net19347), .Q(conv_weight_box[70]) );
  DFFSSRX1_HVT conv_weight_box_reg_32__1_ ( .D(1'b0), .SETB(n294), .RSTB(
        net19352), .CLK(net19364), .Q(conv_weight_box[69]) );
  DFFSSRX1_HVT conv_weight_box_reg_32__0_ ( .D(1'b0), .SETB(n298), .RSTB(
        net19353), .CLK(net19364), .Q(conv_weight_box[68]) );
  DFFSSRX1_HVT conv_weight_box_reg_33__3_ ( .D(1'b0), .SETB(n303), .RSTB(
        net19354), .CLK(net19364), .Q(conv_weight_box[67]) );
  DFFSSRX1_HVT conv_weight_box_reg_33__2_ ( .D(1'b0), .SETB(n293), .RSTB(
        net19355), .CLK(net19364), .Q(conv_weight_box[66]) );
  DFFSSRX1_HVT conv_weight_box_reg_33__1_ ( .D(1'b0), .SETB(n297), .RSTB(
        net19356), .CLK(net19364), .Q(conv_weight_box[65]) );
  DFFSSRX1_HVT conv_weight_box_reg_33__0_ ( .D(1'b0), .SETB(n302), .RSTB(
        net19357), .CLK(net19364), .Q(conv_weight_box[64]) );
  DFFSSRX1_HVT conv_weight_box_reg_34__3_ ( .D(1'b0), .SETB(n302), .RSTB(
        net19358), .CLK(net19364), .Q(conv_weight_box[63]) );
  DFFSSRX1_HVT conv_weight_box_reg_34__2_ ( .D(1'b0), .SETB(n296), .RSTB(
        net19359), .CLK(net19364), .Q(conv_weight_box[62]) );
  DFFSSRX1_HVT conv_weight_box_reg_34__1_ ( .D(1'b0), .SETB(n301), .RSTB(
        net19360), .CLK(net19364), .Q(conv_weight_box[61]) );
  DFFSSRX1_HVT conv_weight_box_reg_34__0_ ( .D(1'b0), .SETB(n295), .RSTB(
        net19361), .CLK(net19364), .Q(conv_weight_box[60]) );
  DFFSSRX1_HVT conv_weight_box_reg_35__3_ ( .D(1'b0), .SETB(n299), .RSTB(
        net19369), .CLK(net19381), .Q(conv_weight_box[59]) );
  DFFSSRX1_HVT conv_weight_box_reg_35__2_ ( .D(1'b0), .SETB(n306), .RSTB(
        net19370), .CLK(net19381), .Q(conv_weight_box[58]) );
  DFFSSRX1_HVT conv_weight_box_reg_35__1_ ( .D(1'b0), .SETB(n294), .RSTB(
        net19371), .CLK(net19381), .Q(conv_weight_box[57]) );
  DFFSSRX1_HVT conv_weight_box_reg_35__0_ ( .D(1'b0), .SETB(n298), .RSTB(
        net19372), .CLK(net19381), .Q(conv_weight_box[56]) );
  DFFSSRX1_HVT conv_weight_box_reg_36__3_ ( .D(1'b0), .SETB(n303), .RSTB(
        net19373), .CLK(net19381), .Q(conv_weight_box[55]) );
  DFFSSRX1_HVT conv_weight_box_reg_36__2_ ( .D(1'b0), .SETB(n293), .RSTB(
        net19374), .CLK(net19381), .Q(conv_weight_box[54]) );
  DFFSSRX1_HVT conv_weight_box_reg_36__1_ ( .D(1'b0), .SETB(n297), .RSTB(
        net19375), .CLK(net19381), .Q(conv_weight_box[53]) );
  DFFSSRX1_HVT conv_weight_box_reg_36__0_ ( .D(1'b0), .SETB(n302), .RSTB(
        net19376), .CLK(net19381), .Q(conv_weight_box[52]) );
  DFFSSRX1_HVT conv_weight_box_reg_37__3_ ( .D(1'b0), .SETB(n303), .RSTB(
        net19377), .CLK(net19381), .Q(conv_weight_box[51]) );
  DFFSSRX1_HVT conv_weight_box_reg_37__2_ ( .D(1'b0), .SETB(n296), .RSTB(
        net19378), .CLK(net19381), .Q(conv_weight_box[50]) );
  DFFSSRX1_HVT conv_weight_box_reg_37__1_ ( .D(1'b0), .SETB(n301), .RSTB(
        net19386), .CLK(net19398), .Q(conv_weight_box[49]) );
  DFFSSRX1_HVT conv_weight_box_reg_37__0_ ( .D(1'b0), .SETB(n295), .RSTB(
        net19387), .CLK(net19398), .Q(conv_weight_box[48]) );
  DFFSSRX1_HVT conv_weight_box_reg_38__3_ ( .D(1'b0), .SETB(n299), .RSTB(
        net19388), .CLK(net19398), .Q(conv_weight_box[47]) );
  DFFSSRX1_HVT conv_weight_box_reg_38__2_ ( .D(1'b0), .SETB(n306), .RSTB(
        net19389), .CLK(net19398), .Q(conv_weight_box[46]) );
  DFFSSRX1_HVT conv_weight_box_reg_38__1_ ( .D(1'b0), .SETB(n294), .RSTB(
        net19390), .CLK(net19398), .Q(conv_weight_box[45]) );
  DFFSSRX1_HVT conv_weight_box_reg_38__0_ ( .D(1'b0), .SETB(n298), .RSTB(
        net19391), .CLK(net19398), .Q(conv_weight_box[44]) );
  DFFSSRX1_HVT conv_weight_box_reg_39__3_ ( .D(1'b0), .SETB(n303), .RSTB(
        net19392), .CLK(net19398), .Q(conv_weight_box[43]) );
  DFFSSRX1_HVT conv_weight_box_reg_39__2_ ( .D(1'b0), .SETB(n293), .RSTB(
        net19393), .CLK(net19398), .Q(conv_weight_box[42]) );
  DFFSSRX1_HVT conv_weight_box_reg_39__1_ ( .D(1'b0), .SETB(n297), .RSTB(
        net19394), .CLK(net19398), .Q(conv_weight_box[41]) );
  DFFSSRX1_HVT conv_weight_box_reg_39__0_ ( .D(1'b0), .SETB(n302), .RSTB(
        net19395), .CLK(net19398), .Q(conv_weight_box[40]) );
  DFFSSRX1_HVT conv_weight_box_reg_40__3_ ( .D(1'b0), .SETB(n301), .RSTB(
        net19403), .CLK(net19415), .Q(conv_weight_box[39]) );
  DFFSSRX1_HVT conv_weight_box_reg_40__2_ ( .D(1'b0), .SETB(n296), .RSTB(
        net19404), .CLK(net19415), .Q(conv_weight_box[38]) );
  DFFSSRX1_HVT conv_weight_box_reg_40__1_ ( .D(1'b0), .SETB(n301), .RSTB(
        net19405), .CLK(net19415), .Q(conv_weight_box[37]) );
  DFFSSRX1_HVT conv_weight_box_reg_40__0_ ( .D(1'b0), .SETB(n295), .RSTB(
        net19406), .CLK(net19415), .Q(conv_weight_box[36]) );
  DFFSSRX1_HVT conv_weight_box_reg_41__3_ ( .D(1'b0), .SETB(n299), .RSTB(
        net19407), .CLK(net19415), .Q(conv_weight_box[35]) );
  DFFSSRX1_HVT conv_weight_box_reg_41__2_ ( .D(1'b0), .SETB(n306), .RSTB(
        net19408), .CLK(net19415), .Q(conv_weight_box[34]) );
  DFFSSRX1_HVT conv_weight_box_reg_41__1_ ( .D(1'b0), .SETB(n294), .RSTB(
        net19409), .CLK(net19415), .Q(conv_weight_box[33]) );
  DFFSSRX1_HVT conv_weight_box_reg_41__0_ ( .D(1'b0), .SETB(n298), .RSTB(
        net19410), .CLK(net19415), .Q(conv_weight_box[32]) );
  DFFSSRX1_HVT conv_weight_box_reg_42__3_ ( .D(1'b0), .SETB(n303), .RSTB(
        net19411), .CLK(net19415), .Q(conv_weight_box[31]) );
  DFFSSRX1_HVT conv_weight_box_reg_42__2_ ( .D(1'b0), .SETB(n293), .RSTB(
        net19412), .CLK(net19415), .Q(conv_weight_box[30]) );
  DFFSSRX1_HVT conv_weight_box_reg_42__1_ ( .D(1'b0), .SETB(n297), .RSTB(
        net19420), .CLK(net19432), .Q(conv_weight_box[29]) );
  DFFSSRX1_HVT conv_weight_box_reg_42__0_ ( .D(1'b0), .SETB(n302), .RSTB(
        net19421), .CLK(net19432), .Q(conv_weight_box[28]) );
  DFFSSRX1_HVT conv_weight_box_reg_43__3_ ( .D(1'b0), .SETB(n306), .RSTB(
        net19422), .CLK(net19432), .Q(conv_weight_box[27]) );
  DFFSSRX1_HVT conv_weight_box_reg_43__2_ ( .D(1'b0), .SETB(n296), .RSTB(
        net19423), .CLK(net19432), .Q(conv_weight_box[26]) );
  DFFSSRX1_HVT conv_weight_box_reg_43__1_ ( .D(1'b0), .SETB(n301), .RSTB(
        net19424), .CLK(net19432), .Q(conv_weight_box[25]) );
  DFFSSRX1_HVT conv_weight_box_reg_43__0_ ( .D(1'b0), .SETB(n295), .RSTB(
        net19425), .CLK(net19432), .Q(conv_weight_box[24]) );
  DFFSSRX1_HVT conv_weight_box_reg_44__3_ ( .D(1'b0), .SETB(n299), .RSTB(
        net19426), .CLK(net19432), .Q(conv_weight_box[23]) );
  DFFSSRX1_HVT conv_weight_box_reg_44__2_ ( .D(1'b0), .SETB(n306), .RSTB(
        net19427), .CLK(net19432), .Q(conv_weight_box[22]) );
  DFFSSRX1_HVT conv_weight_box_reg_44__1_ ( .D(1'b0), .SETB(n294), .RSTB(
        net19428), .CLK(net19432), .Q(conv_weight_box[21]) );
  DFFSSRX1_HVT conv_weight_box_reg_44__0_ ( .D(1'b0), .SETB(n298), .RSTB(
        net19429), .CLK(net19432), .Q(conv_weight_box[20]) );
  DFFSSRX1_HVT conv_weight_box_reg_45__3_ ( .D(1'b0), .SETB(n303), .RSTB(
        net19437), .CLK(net19449), .Q(conv_weight_box[19]) );
  DFFSSRX1_HVT conv_weight_box_reg_45__2_ ( .D(1'b0), .SETB(n293), .RSTB(
        net19438), .CLK(net19449), .Q(conv_weight_box[18]) );
  DFFSSRX1_HVT conv_weight_box_reg_45__1_ ( .D(1'b0), .SETB(n297), .RSTB(
        net19439), .CLK(net19449), .Q(conv_weight_box[17]) );
  DFFSSRX1_HVT conv_weight_box_reg_45__0_ ( .D(1'b0), .SETB(n302), .RSTB(
        net19440), .CLK(net19449), .Q(conv_weight_box[16]) );
  DFFSSRX1_HVT conv_weight_box_reg_46__3_ ( .D(1'b0), .SETB(n296), .RSTB(
        net19441), .CLK(net19449), .Q(conv_weight_box[15]) );
  DFFSSRX1_HVT conv_weight_box_reg_46__2_ ( .D(1'b0), .SETB(n296), .RSTB(
        net19442), .CLK(net19449), .Q(conv_weight_box[14]) );
  DFFSSRX1_HVT conv_weight_box_reg_46__1_ ( .D(1'b0), .SETB(n301), .RSTB(
        net19443), .CLK(net19449), .Q(conv_weight_box[13]) );
  DFFSSRX1_HVT conv_weight_box_reg_46__0_ ( .D(1'b0), .SETB(n295), .RSTB(
        net19444), .CLK(net19449), .Q(conv_weight_box[12]) );
  DFFSSRX1_HVT conv_weight_box_reg_47__3_ ( .D(1'b0), .SETB(n299), .RSTB(
        net19445), .CLK(net19449), .Q(conv_weight_box[11]) );
  DFFSSRX1_HVT conv_weight_box_reg_47__2_ ( .D(1'b0), .SETB(n306), .RSTB(
        net19446), .CLK(net19449), .Q(conv_weight_box[10]) );
  DFFSSRX1_HVT conv_weight_box_reg_47__1_ ( .D(1'b0), .SETB(n294), .RSTB(
        net19454), .CLK(net19466), .Q(conv_weight_box[9]) );
  DFFSSRX1_HVT conv_weight_box_reg_47__0_ ( .D(1'b0), .SETB(n298), .RSTB(
        net19455), .CLK(net19466), .Q(conv_weight_box[8]) );
  DFFSSRX1_HVT conv_weight_box_reg_48__3_ ( .D(1'b0), .SETB(n303), .RSTB(
        net19456), .CLK(net19466), .Q(conv_weight_box[7]) );
  DFFSSRX1_HVT conv_weight_box_reg_48__2_ ( .D(1'b0), .SETB(n293), .RSTB(
        net19457), .CLK(net19466), .Q(conv_weight_box[6]) );
  DFFSSRX1_HVT conv_weight_box_reg_48__1_ ( .D(1'b0), .SETB(n297), .RSTB(
        net19458), .CLK(net19466), .Q(conv_weight_box[5]) );
  DFFSSRX1_HVT conv_weight_box_reg_48__0_ ( .D(1'b0), .SETB(n302), .RSTB(
        net19459), .CLK(net19466), .Q(conv_weight_box[4]) );
  DFFSSRX1_HVT conv_weight_box_reg_49__3_ ( .D(1'b0), .SETB(n299), .RSTB(
        net19460), .CLK(net19466), .Q(conv_weight_box[3]) );
  DFFSSRX1_HVT conv_weight_box_reg_49__2_ ( .D(1'b0), .SETB(n296), .RSTB(
        net19461), .CLK(net19466), .Q(conv_weight_box[2]) );
  DFFSSRX1_HVT conv_weight_box_reg_49__1_ ( .D(1'b0), .SETB(n301), .RSTB(
        net19462), .CLK(net19466), .Q(conv_weight_box[1]) );
  DFFSSRX1_HVT conv_weight_box_reg_49__0_ ( .D(1'b0), .SETB(n295), .RSTB(
        net19463), .CLK(net19466), .Q(conv_weight_box[0]) );
  DFFSSRX1_HVT bias_data_reg_3_ ( .D(1'b0), .SETB(n299), .RSTB(net19483), 
        .CLK(net19498), .Q(bias_data[3]) );
  DFFSSRX1_HVT bias_data_reg_2_ ( .D(1'b0), .SETB(n306), .RSTB(net19487), 
        .CLK(net19498), .Q(bias_data[2]) );
  DFFSSRX1_HVT bias_data_reg_1_ ( .D(1'b0), .SETB(n294), .RSTB(net19491), 
        .CLK(net19498), .Q(bias_data[1]) );
  DFFSSRX1_HVT bias_data_reg_0_ ( .D(1'b0), .SETB(n298), .RSTB(net19495), 
        .CLK(net19498), .Q(bias_data[0]) );
  AO22X1_HVT U3 ( .A1(conv_weight_box[8]), .A2(n346), .A3(conv_weight_box[12]), 
        .A4(n347), .Y(n1) );
  AO22X1_HVT U4 ( .A1(conv_weight_box[84]), .A2(n348), .A3(conv_weight_box[80]), .A4(n349), .Y(n2) );
  AO22X1_HVT U5 ( .A1(conv_weight_box[20]), .A2(n350), .A3(conv_weight_box[72]), .A4(n351), .Y(n3) );
  AO22X1_HVT U6 ( .A1(conv_weight_box[68]), .A2(n352), .A3(conv_weight_box[64]), .A4(n353), .Y(n4) );
  NOR4X0_HVT U7 ( .A1(n1), .A2(n2), .A3(n3), .A4(n4), .Y(n5) );
  AO22X1_HVT U8 ( .A1(n369), .A2(conv_weight_box[96]), .A3(n367), .A4(
        conv_weight_box[112]), .Y(n6) );
  AO22X1_HVT U9 ( .A1(conv_weight_box[32]), .A2(n363), .A3(conv_weight_box[48]), .A4(n361), .Y(n7) );
  AO22X1_HVT U10 ( .A1(n362), .A2(conv_weight_box[192]), .A3(
        conv_weight_box[176]), .A4(n360), .Y(n8) );
  AO22X1_HVT U11 ( .A1(n364), .A2(conv_weight_box[160]), .A3(n365), .A4(
        conv_weight_box[144]), .Y(n9) );
  NOR4X0_HVT U12 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .Y(n10) );
  AO22X1_HVT U13 ( .A1(n369), .A2(conv_weight_box[100]), .A3(n367), .A4(
        conv_weight_box[116]), .Y(n11) );
  AO22X1_HVT U14 ( .A1(conv_weight_box[36]), .A2(n363), .A3(
        conv_weight_box[52]), .A4(n361), .Y(n12) );
  AO22X1_HVT U15 ( .A1(n362), .A2(conv_weight_box[196]), .A3(
        conv_weight_box[180]), .A4(n360), .Y(n13) );
  AO22X1_HVT U16 ( .A1(n364), .A2(conv_weight_box[164]), .A3(n365), .A4(
        conv_weight_box[148]), .Y(n14) );
  NOR4X0_HVT U17 ( .A1(n11), .A2(n12), .A3(n13), .A4(n14), .Y(n15) );
  OA22X1_HVT U18 ( .A1(n10), .A2(n344), .A3(n15), .A4(n345), .Y(n16) );
  AO22X1_HVT U19 ( .A1(conv_weight_box[76]), .A2(n358), .A3(
        conv_weight_box[128]), .A4(n359), .Y(n17) );
  AO22X1_HVT U20 ( .A1(conv_weight_box[132]), .A2(n354), .A3(
        conv_weight_box[16]), .A4(n355), .Y(n18) );
  AO22X1_HVT U21 ( .A1(conv_weight_box[4]), .A2(n356), .A3(conv_weight_box[0]), 
        .A4(n357), .Y(n19) );
  AO22X1_HVT U22 ( .A1(n368), .A2(conv_weight_box[124]), .A3(n369), .A4(
        conv_weight_box[92]), .Y(n20) );
  AO22X1_HVT U23 ( .A1(n366), .A2(conv_weight_box[60]), .A3(n367), .A4(
        conv_weight_box[108]), .Y(n21) );
  AO22X1_HVT U24 ( .A1(n364), .A2(conv_weight_box[156]), .A3(n365), .A4(
        conv_weight_box[140]), .Y(n22) );
  OR3X1_HVT U25 ( .A1(n20), .A2(n21), .A3(n22), .Y(n23) );
  AO22X1_HVT U26 ( .A1(n362), .A2(conv_weight_box[188]), .A3(
        conv_weight_box[28]), .A4(n363), .Y(n24) );
  AO22X1_HVT U27 ( .A1(conv_weight_box[172]), .A2(n360), .A3(
        conv_weight_box[44]), .A4(n361), .Y(n25) );
  OR3X1_HVT U28 ( .A1(n23), .A2(n24), .A3(n25), .Y(n26) );
  AO22X1_HVT U29 ( .A1(n368), .A2(conv_weight_box[120]), .A3(n369), .A4(
        conv_weight_box[88]), .Y(n27) );
  AO22X1_HVT U30 ( .A1(n366), .A2(conv_weight_box[56]), .A3(n367), .A4(
        conv_weight_box[104]), .Y(n28) );
  AO22X1_HVT U31 ( .A1(n364), .A2(conv_weight_box[152]), .A3(n365), .A4(
        conv_weight_box[136]), .Y(n29) );
  OR3X1_HVT U32 ( .A1(n27), .A2(n28), .A3(n29), .Y(n30) );
  AO22X1_HVT U33 ( .A1(n362), .A2(conv_weight_box[184]), .A3(
        conv_weight_box[24]), .A4(n363), .Y(n31) );
  AO22X1_HVT U34 ( .A1(conv_weight_box[168]), .A2(n360), .A3(
        conv_weight_box[40]), .A4(n361), .Y(n32) );
  OR3X1_HVT U35 ( .A1(n30), .A2(n31), .A3(n32), .Y(n33) );
  AO22X1_HVT U36 ( .A1(n371), .A2(n26), .A3(n370), .A4(n33), .Y(n34) );
  NOR4X0_HVT U37 ( .A1(n17), .A2(n18), .A3(n19), .A4(n34), .Y(n35) );
  NAND3X0_HVT U38 ( .A1(n5), .A2(n16), .A3(n35), .Y(n36) );
  AO22X1_HVT U39 ( .A1(conv_weight_box[8]), .A2(n374), .A3(conv_weight_box[12]), .A4(n375), .Y(n37) );
  AO22X1_HVT U40 ( .A1(conv_weight_box[84]), .A2(n376), .A3(
        conv_weight_box[80]), .A4(n377), .Y(n38) );
  AO22X1_HVT U41 ( .A1(conv_weight_box[20]), .A2(n378), .A3(
        conv_weight_box[72]), .A4(n379), .Y(n39) );
  AO22X1_HVT U42 ( .A1(conv_weight_box[68]), .A2(n380), .A3(
        conv_weight_box[64]), .A4(n381), .Y(n40) );
  NOR4X0_HVT U43 ( .A1(n37), .A2(n38), .A3(n39), .A4(n40), .Y(n41) );
  AO22X1_HVT U44 ( .A1(n397), .A2(conv_weight_box[96]), .A3(n395), .A4(
        conv_weight_box[112]), .Y(n42) );
  AO22X1_HVT U45 ( .A1(conv_weight_box[32]), .A2(n391), .A3(
        conv_weight_box[48]), .A4(n389), .Y(n43) );
  AO22X1_HVT U46 ( .A1(conv_weight_box[192]), .A2(n390), .A3(
        conv_weight_box[176]), .A4(n388), .Y(n44) );
  AO22X1_HVT U47 ( .A1(n392), .A2(conv_weight_box[160]), .A3(n393), .A4(
        conv_weight_box[144]), .Y(n45) );
  NOR4X0_HVT U48 ( .A1(n42), .A2(n43), .A3(n44), .A4(n45), .Y(n46) );
  AO22X1_HVT U49 ( .A1(n397), .A2(conv_weight_box[100]), .A3(n395), .A4(
        conv_weight_box[116]), .Y(n47) );
  AO22X1_HVT U50 ( .A1(n391), .A2(conv_weight_box[36]), .A3(n389), .A4(
        conv_weight_box[52]), .Y(n48) );
  AO22X1_HVT U51 ( .A1(n390), .A2(conv_weight_box[196]), .A3(n388), .A4(
        conv_weight_box[180]), .Y(n49) );
  AO22X1_HVT U52 ( .A1(n392), .A2(conv_weight_box[164]), .A3(n393), .A4(
        conv_weight_box[148]), .Y(n50) );
  NOR4X0_HVT U53 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .Y(n51) );
  OA22X1_HVT U54 ( .A1(n46), .A2(n372), .A3(n51), .A4(n373), .Y(n52) );
  AO22X1_HVT U55 ( .A1(conv_weight_box[76]), .A2(n386), .A3(
        conv_weight_box[128]), .A4(n387), .Y(n53) );
  AO22X1_HVT U56 ( .A1(conv_weight_box[132]), .A2(n382), .A3(
        conv_weight_box[16]), .A4(n383), .Y(n54) );
  AO22X1_HVT U57 ( .A1(conv_weight_box[4]), .A2(n384), .A3(conv_weight_box[0]), 
        .A4(n385), .Y(n55) );
  AO22X1_HVT U58 ( .A1(n396), .A2(conv_weight_box[124]), .A3(n397), .A4(
        conv_weight_box[92]), .Y(n56) );
  AO22X1_HVT U59 ( .A1(n394), .A2(conv_weight_box[60]), .A3(n395), .A4(
        conv_weight_box[108]), .Y(n57) );
  AO22X1_HVT U60 ( .A1(n392), .A2(conv_weight_box[156]), .A3(n393), .A4(
        conv_weight_box[140]), .Y(n58) );
  OR3X1_HVT U61 ( .A1(n56), .A2(n57), .A3(n58), .Y(n59) );
  AO22X1_HVT U62 ( .A1(n391), .A2(conv_weight_box[28]), .A3(n390), .A4(
        conv_weight_box[188]), .Y(n60) );
  AO22X1_HVT U63 ( .A1(n389), .A2(conv_weight_box[44]), .A3(n388), .A4(
        conv_weight_box[172]), .Y(n61) );
  OR3X1_HVT U64 ( .A1(n59), .A2(n60), .A3(n61), .Y(n62) );
  AO22X1_HVT U65 ( .A1(n396), .A2(conv_weight_box[120]), .A3(n397), .A4(
        conv_weight_box[88]), .Y(n63) );
  AO22X1_HVT U66 ( .A1(n394), .A2(conv_weight_box[56]), .A3(n395), .A4(
        conv_weight_box[104]), .Y(n64) );
  AO22X1_HVT U67 ( .A1(n392), .A2(conv_weight_box[152]), .A3(n393), .A4(
        conv_weight_box[136]), .Y(n65) );
  OR3X1_HVT U68 ( .A1(n63), .A2(n64), .A3(n65), .Y(n66) );
  AO22X1_HVT U69 ( .A1(n391), .A2(conv_weight_box[24]), .A3(n390), .A4(
        conv_weight_box[184]), .Y(n67) );
  AO22X1_HVT U70 ( .A1(n389), .A2(conv_weight_box[40]), .A3(n388), .A4(
        conv_weight_box[168]), .Y(n68) );
  OR3X1_HVT U71 ( .A1(n66), .A2(n67), .A3(n68), .Y(n69) );
  AO22X1_HVT U72 ( .A1(n399), .A2(n62), .A3(n398), .A4(n69), .Y(n70) );
  NOR4X0_HVT U73 ( .A1(n53), .A2(n54), .A3(n55), .A4(n70), .Y(n71) );
  NAND3X0_HVT U74 ( .A1(n41), .A2(n52), .A3(n71), .Y(n72) );
  AO22X1_HVT U75 ( .A1(n401), .A2(n36), .A3(n400), .A4(n72), .Y(net19495) );
  AO22X1_HVT U76 ( .A1(conv_weight_box[9]), .A2(n346), .A3(conv_weight_box[13]), .A4(n347), .Y(n73) );
  AO22X1_HVT U77 ( .A1(conv_weight_box[85]), .A2(n348), .A3(
        conv_weight_box[81]), .A4(n349), .Y(n74) );
  AO22X1_HVT U78 ( .A1(conv_weight_box[21]), .A2(n350), .A3(
        conv_weight_box[73]), .A4(n351), .Y(n75) );
  AO22X1_HVT U79 ( .A1(conv_weight_box[69]), .A2(n352), .A3(
        conv_weight_box[65]), .A4(n353), .Y(n76) );
  NOR4X0_HVT U80 ( .A1(n73), .A2(n74), .A3(n75), .A4(n76), .Y(n77) );
  AO22X1_HVT U81 ( .A1(n369), .A2(conv_weight_box[97]), .A3(n367), .A4(
        conv_weight_box[113]), .Y(n78) );
  AO22X1_HVT U82 ( .A1(conv_weight_box[33]), .A2(n363), .A3(
        conv_weight_box[49]), .A4(n361), .Y(n79) );
  AO22X1_HVT U83 ( .A1(n362), .A2(conv_weight_box[193]), .A3(
        conv_weight_box[177]), .A4(n360), .Y(n80) );
  AO22X1_HVT U84 ( .A1(n364), .A2(conv_weight_box[161]), .A3(n365), .A4(
        conv_weight_box[145]), .Y(n81) );
  NOR4X0_HVT U85 ( .A1(n78), .A2(n79), .A3(n80), .A4(n81), .Y(n82) );
  AO22X1_HVT U86 ( .A1(n369), .A2(conv_weight_box[101]), .A3(n367), .A4(
        conv_weight_box[117]), .Y(n83) );
  AO22X1_HVT U87 ( .A1(conv_weight_box[37]), .A2(n363), .A3(
        conv_weight_box[53]), .A4(n361), .Y(n84) );
  AO22X1_HVT U88 ( .A1(n362), .A2(conv_weight_box[197]), .A3(
        conv_weight_box[181]), .A4(n360), .Y(n85) );
  AO22X1_HVT U89 ( .A1(n364), .A2(conv_weight_box[165]), .A3(n365), .A4(
        conv_weight_box[149]), .Y(n86) );
  NOR4X0_HVT U90 ( .A1(n83), .A2(n84), .A3(n85), .A4(n86), .Y(n87) );
  OA22X1_HVT U91 ( .A1(n82), .A2(n344), .A3(n87), .A4(n345), .Y(n88) );
  AO22X1_HVT U92 ( .A1(conv_weight_box[77]), .A2(n358), .A3(
        conv_weight_box[129]), .A4(n359), .Y(n89) );
  AO22X1_HVT U93 ( .A1(conv_weight_box[133]), .A2(n354), .A3(
        conv_weight_box[17]), .A4(n355), .Y(n90) );
  AO22X1_HVT U94 ( .A1(conv_weight_box[5]), .A2(n356), .A3(conv_weight_box[1]), 
        .A4(n357), .Y(n91) );
  AO22X1_HVT U95 ( .A1(n368), .A2(conv_weight_box[125]), .A3(n369), .A4(
        conv_weight_box[93]), .Y(n92) );
  AO22X1_HVT U96 ( .A1(n366), .A2(conv_weight_box[61]), .A3(n367), .A4(
        conv_weight_box[109]), .Y(n93) );
  AO22X1_HVT U97 ( .A1(n364), .A2(conv_weight_box[157]), .A3(n365), .A4(
        conv_weight_box[141]), .Y(n94) );
  OR3X1_HVT U98 ( .A1(n92), .A2(n93), .A3(n94), .Y(n95) );
  AO22X1_HVT U99 ( .A1(n362), .A2(conv_weight_box[189]), .A3(
        conv_weight_box[29]), .A4(n363), .Y(n96) );
  AO22X1_HVT U100 ( .A1(conv_weight_box[173]), .A2(n360), .A3(
        conv_weight_box[45]), .A4(n361), .Y(n97) );
  OR3X1_HVT U101 ( .A1(n95), .A2(n96), .A3(n97), .Y(n98) );
  AO22X1_HVT U102 ( .A1(n368), .A2(conv_weight_box[121]), .A3(n369), .A4(
        conv_weight_box[89]), .Y(n99) );
  AO22X1_HVT U103 ( .A1(n366), .A2(conv_weight_box[57]), .A3(n367), .A4(
        conv_weight_box[105]), .Y(n100) );
  AO22X1_HVT U104 ( .A1(n364), .A2(conv_weight_box[153]), .A3(n365), .A4(
        conv_weight_box[137]), .Y(n101) );
  OR3X1_HVT U105 ( .A1(n99), .A2(n100), .A3(n101), .Y(n102) );
  AO22X1_HVT U106 ( .A1(n362), .A2(conv_weight_box[185]), .A3(
        conv_weight_box[25]), .A4(n363), .Y(n103) );
  AO22X1_HVT U107 ( .A1(conv_weight_box[169]), .A2(n360), .A3(
        conv_weight_box[41]), .A4(n361), .Y(n104) );
  OR3X1_HVT U108 ( .A1(n102), .A2(n103), .A3(n104), .Y(n105) );
  AO22X1_HVT U109 ( .A1(n371), .A2(n98), .A3(n370), .A4(n105), .Y(n106) );
  NOR4X0_HVT U110 ( .A1(n89), .A2(n90), .A3(n91), .A4(n106), .Y(n107) );
  NAND3X0_HVT U111 ( .A1(n77), .A2(n88), .A3(n107), .Y(n108) );
  AO22X1_HVT U112 ( .A1(conv_weight_box[9]), .A2(n374), .A3(
        conv_weight_box[13]), .A4(n375), .Y(n109) );
  AO22X1_HVT U113 ( .A1(conv_weight_box[85]), .A2(n376), .A3(
        conv_weight_box[81]), .A4(n377), .Y(n110) );
  AO22X1_HVT U114 ( .A1(conv_weight_box[21]), .A2(n378), .A3(
        conv_weight_box[73]), .A4(n379), .Y(n111) );
  AO22X1_HVT U115 ( .A1(conv_weight_box[69]), .A2(n380), .A3(
        conv_weight_box[65]), .A4(n381), .Y(n112) );
  NOR4X0_HVT U116 ( .A1(n109), .A2(n110), .A3(n111), .A4(n112), .Y(n113) );
  AO22X1_HVT U117 ( .A1(n397), .A2(conv_weight_box[97]), .A3(n395), .A4(
        conv_weight_box[113]), .Y(n114) );
  AO22X1_HVT U118 ( .A1(conv_weight_box[33]), .A2(n391), .A3(
        conv_weight_box[49]), .A4(n389), .Y(n115) );
  AO22X1_HVT U119 ( .A1(conv_weight_box[193]), .A2(n390), .A3(
        conv_weight_box[177]), .A4(n388), .Y(n116) );
  AO22X1_HVT U120 ( .A1(n392), .A2(conv_weight_box[161]), .A3(n393), .A4(
        conv_weight_box[145]), .Y(n117) );
  NOR4X0_HVT U121 ( .A1(n114), .A2(n115), .A3(n116), .A4(n117), .Y(n118) );
  AO22X1_HVT U122 ( .A1(n397), .A2(conv_weight_box[101]), .A3(n395), .A4(
        conv_weight_box[117]), .Y(n119) );
  AO22X1_HVT U123 ( .A1(n391), .A2(conv_weight_box[37]), .A3(n389), .A4(
        conv_weight_box[53]), .Y(n120) );
  AO22X1_HVT U124 ( .A1(n390), .A2(conv_weight_box[197]), .A3(n388), .A4(
        conv_weight_box[181]), .Y(n121) );
  AO22X1_HVT U125 ( .A1(n392), .A2(conv_weight_box[165]), .A3(n393), .A4(
        conv_weight_box[149]), .Y(n122) );
  NOR4X0_HVT U126 ( .A1(n119), .A2(n120), .A3(n121), .A4(n122), .Y(n123) );
  OA22X1_HVT U127 ( .A1(n118), .A2(n372), .A3(n123), .A4(n373), .Y(n124) );
  AO22X1_HVT U128 ( .A1(conv_weight_box[77]), .A2(n386), .A3(
        conv_weight_box[129]), .A4(n387), .Y(n125) );
  AO22X1_HVT U129 ( .A1(conv_weight_box[133]), .A2(n382), .A3(
        conv_weight_box[17]), .A4(n383), .Y(n126) );
  AO22X1_HVT U130 ( .A1(conv_weight_box[5]), .A2(n384), .A3(conv_weight_box[1]), .A4(n385), .Y(n127) );
  AO22X1_HVT U131 ( .A1(n396), .A2(conv_weight_box[125]), .A3(n397), .A4(
        conv_weight_box[93]), .Y(n128) );
  AO22X1_HVT U132 ( .A1(n394), .A2(conv_weight_box[61]), .A3(n395), .A4(
        conv_weight_box[109]), .Y(n129) );
  AO22X1_HVT U133 ( .A1(n392), .A2(conv_weight_box[157]), .A3(n393), .A4(
        conv_weight_box[141]), .Y(n130) );
  OR3X1_HVT U134 ( .A1(n128), .A2(n129), .A3(n130), .Y(n131) );
  AO22X1_HVT U135 ( .A1(n391), .A2(conv_weight_box[29]), .A3(n390), .A4(
        conv_weight_box[189]), .Y(n132) );
  AO22X1_HVT U136 ( .A1(n389), .A2(conv_weight_box[45]), .A3(n388), .A4(
        conv_weight_box[173]), .Y(n133) );
  OR3X1_HVT U137 ( .A1(n131), .A2(n132), .A3(n133), .Y(n134) );
  AO22X1_HVT U138 ( .A1(n396), .A2(conv_weight_box[121]), .A3(n397), .A4(
        conv_weight_box[89]), .Y(n135) );
  AO22X1_HVT U139 ( .A1(n394), .A2(conv_weight_box[57]), .A3(n395), .A4(
        conv_weight_box[105]), .Y(n136) );
  AO22X1_HVT U140 ( .A1(n392), .A2(conv_weight_box[153]), .A3(n393), .A4(
        conv_weight_box[137]), .Y(n137) );
  OR3X1_HVT U141 ( .A1(n135), .A2(n136), .A3(n137), .Y(n138) );
  AO22X1_HVT U142 ( .A1(n391), .A2(conv_weight_box[25]), .A3(n390), .A4(
        conv_weight_box[185]), .Y(n139) );
  AO22X1_HVT U143 ( .A1(n389), .A2(conv_weight_box[41]), .A3(n388), .A4(
        conv_weight_box[169]), .Y(n140) );
  OR3X1_HVT U144 ( .A1(n138), .A2(n139), .A3(n140), .Y(n141) );
  AO22X1_HVT U145 ( .A1(n399), .A2(n134), .A3(n398), .A4(n141), .Y(n142) );
  NOR4X0_HVT U146 ( .A1(n125), .A2(n126), .A3(n127), .A4(n142), .Y(n143) );
  NAND3X0_HVT U147 ( .A1(n113), .A2(n124), .A3(n143), .Y(n144) );
  AO22X1_HVT U148 ( .A1(n401), .A2(n108), .A3(n400), .A4(n144), .Y(net19491)
         );
  AO22X1_HVT U149 ( .A1(conv_weight_box[10]), .A2(n346), .A3(
        conv_weight_box[14]), .A4(n347), .Y(n145) );
  AO22X1_HVT U150 ( .A1(conv_weight_box[86]), .A2(n348), .A3(
        conv_weight_box[82]), .A4(n349), .Y(n146) );
  AO22X1_HVT U151 ( .A1(conv_weight_box[22]), .A2(n350), .A3(
        conv_weight_box[74]), .A4(n351), .Y(n147) );
  AO22X1_HVT U152 ( .A1(conv_weight_box[70]), .A2(n352), .A3(
        conv_weight_box[66]), .A4(n353), .Y(n148) );
  NOR4X0_HVT U153 ( .A1(n145), .A2(n146), .A3(n147), .A4(n148), .Y(n149) );
  AO22X1_HVT U154 ( .A1(n369), .A2(conv_weight_box[98]), .A3(n367), .A4(
        conv_weight_box[114]), .Y(n150) );
  AO22X1_HVT U155 ( .A1(conv_weight_box[34]), .A2(n363), .A3(
        conv_weight_box[50]), .A4(n361), .Y(n151) );
  AO22X1_HVT U156 ( .A1(n362), .A2(conv_weight_box[194]), .A3(
        conv_weight_box[178]), .A4(n360), .Y(n152) );
  AO22X1_HVT U157 ( .A1(n364), .A2(conv_weight_box[162]), .A3(n365), .A4(
        conv_weight_box[146]), .Y(n153) );
  NOR4X0_HVT U158 ( .A1(n150), .A2(n151), .A3(n152), .A4(n153), .Y(n154) );
  AO22X1_HVT U159 ( .A1(n369), .A2(conv_weight_box[102]), .A3(n367), .A4(
        conv_weight_box[118]), .Y(n155) );
  AO22X1_HVT U160 ( .A1(conv_weight_box[38]), .A2(n363), .A3(
        conv_weight_box[54]), .A4(n361), .Y(n156) );
  AO22X1_HVT U161 ( .A1(n362), .A2(conv_weight_box[198]), .A3(
        conv_weight_box[182]), .A4(n360), .Y(n157) );
  AO22X1_HVT U162 ( .A1(n364), .A2(conv_weight_box[166]), .A3(n365), .A4(
        conv_weight_box[150]), .Y(n158) );
  NOR4X0_HVT U163 ( .A1(n155), .A2(n156), .A3(n157), .A4(n158), .Y(n159) );
  OA22X1_HVT U164 ( .A1(n154), .A2(n344), .A3(n159), .A4(n345), .Y(n160) );
  AO22X1_HVT U165 ( .A1(conv_weight_box[78]), .A2(n358), .A3(
        conv_weight_box[130]), .A4(n359), .Y(n161) );
  AO22X1_HVT U166 ( .A1(conv_weight_box[134]), .A2(n354), .A3(
        conv_weight_box[18]), .A4(n355), .Y(n162) );
  AO22X1_HVT U167 ( .A1(conv_weight_box[6]), .A2(n356), .A3(conv_weight_box[2]), .A4(n357), .Y(n163) );
  AO22X1_HVT U168 ( .A1(n368), .A2(conv_weight_box[126]), .A3(n369), .A4(
        conv_weight_box[94]), .Y(n164) );
  AO22X1_HVT U169 ( .A1(n366), .A2(conv_weight_box[62]), .A3(n367), .A4(
        conv_weight_box[110]), .Y(n165) );
  AO22X1_HVT U170 ( .A1(n364), .A2(conv_weight_box[158]), .A3(n365), .A4(
        conv_weight_box[142]), .Y(n166) );
  OR3X1_HVT U171 ( .A1(n164), .A2(n165), .A3(n166), .Y(n167) );
  AO22X1_HVT U172 ( .A1(n362), .A2(conv_weight_box[190]), .A3(
        conv_weight_box[30]), .A4(n363), .Y(n168) );
  AO22X1_HVT U173 ( .A1(conv_weight_box[174]), .A2(n360), .A3(
        conv_weight_box[46]), .A4(n361), .Y(n169) );
  OR3X1_HVT U174 ( .A1(n167), .A2(n168), .A3(n169), .Y(n170) );
  AO22X1_HVT U175 ( .A1(n368), .A2(conv_weight_box[122]), .A3(n369), .A4(
        conv_weight_box[90]), .Y(n171) );
  AO22X1_HVT U176 ( .A1(n366), .A2(conv_weight_box[58]), .A3(n367), .A4(
        conv_weight_box[106]), .Y(n172) );
  AO22X1_HVT U177 ( .A1(n364), .A2(conv_weight_box[154]), .A3(n365), .A4(
        conv_weight_box[138]), .Y(n173) );
  OR3X1_HVT U178 ( .A1(n171), .A2(n172), .A3(n173), .Y(n174) );
  AO22X1_HVT U179 ( .A1(n362), .A2(conv_weight_box[186]), .A3(
        conv_weight_box[26]), .A4(n363), .Y(n175) );
  AO22X1_HVT U180 ( .A1(conv_weight_box[170]), .A2(n360), .A3(
        conv_weight_box[42]), .A4(n361), .Y(n176) );
  OR3X1_HVT U181 ( .A1(n174), .A2(n175), .A3(n176), .Y(n177) );
  AO22X1_HVT U182 ( .A1(n371), .A2(n170), .A3(n370), .A4(n177), .Y(n178) );
  NOR4X0_HVT U183 ( .A1(n161), .A2(n162), .A3(n163), .A4(n178), .Y(n179) );
  NAND3X0_HVT U184 ( .A1(n149), .A2(n160), .A3(n179), .Y(n180) );
  AO22X1_HVT U185 ( .A1(conv_weight_box[10]), .A2(n374), .A3(
        conv_weight_box[14]), .A4(n375), .Y(n181) );
  AO22X1_HVT U186 ( .A1(conv_weight_box[86]), .A2(n376), .A3(
        conv_weight_box[82]), .A4(n377), .Y(n182) );
  AO22X1_HVT U187 ( .A1(conv_weight_box[22]), .A2(n378), .A3(
        conv_weight_box[74]), .A4(n379), .Y(n183) );
  AO22X1_HVT U188 ( .A1(conv_weight_box[70]), .A2(n380), .A3(
        conv_weight_box[66]), .A4(n381), .Y(n184) );
  NOR4X0_HVT U189 ( .A1(n181), .A2(n182), .A3(n183), .A4(n184), .Y(n185) );
  AO22X1_HVT U190 ( .A1(n397), .A2(conv_weight_box[98]), .A3(n395), .A4(
        conv_weight_box[114]), .Y(n186) );
  AO22X1_HVT U191 ( .A1(conv_weight_box[34]), .A2(n391), .A3(
        conv_weight_box[50]), .A4(n389), .Y(n187) );
  AO22X1_HVT U192 ( .A1(conv_weight_box[194]), .A2(n390), .A3(
        conv_weight_box[178]), .A4(n388), .Y(n188) );
  AO22X1_HVT U193 ( .A1(n392), .A2(conv_weight_box[162]), .A3(n393), .A4(
        conv_weight_box[146]), .Y(n189) );
  NOR4X0_HVT U194 ( .A1(n186), .A2(n187), .A3(n188), .A4(n189), .Y(n190) );
  AO22X1_HVT U195 ( .A1(n397), .A2(conv_weight_box[102]), .A3(n395), .A4(
        conv_weight_box[118]), .Y(n191) );
  AO22X1_HVT U196 ( .A1(n391), .A2(conv_weight_box[38]), .A3(n389), .A4(
        conv_weight_box[54]), .Y(n192) );
  AO22X1_HVT U197 ( .A1(n390), .A2(conv_weight_box[198]), .A3(n388), .A4(
        conv_weight_box[182]), .Y(n193) );
  AO22X1_HVT U198 ( .A1(n392), .A2(conv_weight_box[166]), .A3(n393), .A4(
        conv_weight_box[150]), .Y(n194) );
  NOR4X0_HVT U199 ( .A1(n191), .A2(n192), .A3(n193), .A4(n194), .Y(n195) );
  OA22X1_HVT U200 ( .A1(n190), .A2(n372), .A3(n195), .A4(n373), .Y(n196) );
  AO22X1_HVT U201 ( .A1(conv_weight_box[78]), .A2(n386), .A3(
        conv_weight_box[130]), .A4(n387), .Y(n197) );
  AO22X1_HVT U202 ( .A1(conv_weight_box[134]), .A2(n382), .A3(
        conv_weight_box[18]), .A4(n383), .Y(n198) );
  AO22X1_HVT U203 ( .A1(conv_weight_box[6]), .A2(n384), .A3(conv_weight_box[2]), .A4(n385), .Y(n199) );
  AO22X1_HVT U204 ( .A1(n396), .A2(conv_weight_box[126]), .A3(n397), .A4(
        conv_weight_box[94]), .Y(n200) );
  AO22X1_HVT U205 ( .A1(n394), .A2(conv_weight_box[62]), .A3(n395), .A4(
        conv_weight_box[110]), .Y(n201) );
  AO22X1_HVT U206 ( .A1(n392), .A2(conv_weight_box[158]), .A3(n393), .A4(
        conv_weight_box[142]), .Y(n202) );
  OR3X1_HVT U207 ( .A1(n200), .A2(n201), .A3(n202), .Y(n203) );
  AO22X1_HVT U208 ( .A1(n391), .A2(conv_weight_box[30]), .A3(n390), .A4(
        conv_weight_box[190]), .Y(n204) );
  AO22X1_HVT U209 ( .A1(n389), .A2(conv_weight_box[46]), .A3(n388), .A4(
        conv_weight_box[174]), .Y(n205) );
  OR3X1_HVT U210 ( .A1(n203), .A2(n204), .A3(n205), .Y(n206) );
  AO22X1_HVT U211 ( .A1(n396), .A2(conv_weight_box[122]), .A3(n397), .A4(
        conv_weight_box[90]), .Y(n207) );
  AO22X1_HVT U212 ( .A1(n394), .A2(conv_weight_box[58]), .A3(n395), .A4(
        conv_weight_box[106]), .Y(n208) );
  AO22X1_HVT U213 ( .A1(n392), .A2(conv_weight_box[154]), .A3(n393), .A4(
        conv_weight_box[138]), .Y(n209) );
  OR3X1_HVT U214 ( .A1(n207), .A2(n208), .A3(n209), .Y(n210) );
  AO22X1_HVT U215 ( .A1(n391), .A2(conv_weight_box[26]), .A3(n390), .A4(
        conv_weight_box[186]), .Y(n211) );
  AO22X1_HVT U216 ( .A1(n389), .A2(conv_weight_box[42]), .A3(n388), .A4(
        conv_weight_box[170]), .Y(n212) );
  OR3X1_HVT U217 ( .A1(n210), .A2(n211), .A3(n212), .Y(n213) );
  AO22X1_HVT U218 ( .A1(n399), .A2(n206), .A3(n398), .A4(n213), .Y(n214) );
  NOR4X0_HVT U219 ( .A1(n197), .A2(n198), .A3(n199), .A4(n214), .Y(n215) );
  NAND3X0_HVT U220 ( .A1(n185), .A2(n196), .A3(n215), .Y(n216) );
  AO22X1_HVT U221 ( .A1(n401), .A2(n180), .A3(n400), .A4(n216), .Y(net19487)
         );
  AO22X1_HVT U222 ( .A1(conv_weight_box[11]), .A2(n346), .A3(
        conv_weight_box[15]), .A4(n347), .Y(n217) );
  AO22X1_HVT U223 ( .A1(conv_weight_box[87]), .A2(n348), .A3(
        conv_weight_box[83]), .A4(n349), .Y(n218) );
  AO22X1_HVT U224 ( .A1(conv_weight_box[23]), .A2(n350), .A3(
        conv_weight_box[75]), .A4(n351), .Y(n219) );
  AO22X1_HVT U225 ( .A1(conv_weight_box[71]), .A2(n352), .A3(
        conv_weight_box[67]), .A4(n353), .Y(n220) );
  NOR4X0_HVT U226 ( .A1(n217), .A2(n218), .A3(n219), .A4(n220), .Y(n221) );
  AO22X1_HVT U227 ( .A1(conv_weight_box[99]), .A2(n369), .A3(
        conv_weight_box[115]), .A4(n367), .Y(n222) );
  AO22X1_HVT U228 ( .A1(conv_weight_box[35]), .A2(n363), .A3(
        conv_weight_box[51]), .A4(n361), .Y(n223) );
  AO22X1_HVT U229 ( .A1(conv_weight_box[179]), .A2(n360), .A3(
        conv_weight_box[195]), .A4(n362), .Y(n224) );
  AO22X1_HVT U230 ( .A1(n365), .A2(conv_weight_box[147]), .A3(
        conv_weight_box[163]), .A4(n364), .Y(n225) );
  NOR4X0_HVT U231 ( .A1(n222), .A2(n223), .A3(n224), .A4(n225), .Y(n226) );
  AO22X1_HVT U232 ( .A1(conv_weight_box[103]), .A2(n369), .A3(
        conv_weight_box[119]), .A4(n367), .Y(n227) );
  AO22X1_HVT U233 ( .A1(conv_weight_box[39]), .A2(n363), .A3(
        conv_weight_box[55]), .A4(n361), .Y(n228) );
  AO22X1_HVT U234 ( .A1(conv_weight_box[183]), .A2(n360), .A3(
        conv_weight_box[199]), .A4(n362), .Y(n229) );
  AO22X1_HVT U235 ( .A1(n365), .A2(conv_weight_box[151]), .A3(
        conv_weight_box[167]), .A4(n364), .Y(n230) );
  NOR4X0_HVT U236 ( .A1(n227), .A2(n228), .A3(n229), .A4(n230), .Y(n231) );
  OA22X1_HVT U237 ( .A1(n226), .A2(n344), .A3(n231), .A4(n345), .Y(n232) );
  AO22X1_HVT U238 ( .A1(conv_weight_box[79]), .A2(n358), .A3(
        conv_weight_box[131]), .A4(n359), .Y(n233) );
  AO22X1_HVT U239 ( .A1(conv_weight_box[135]), .A2(n354), .A3(
        conv_weight_box[19]), .A4(n355), .Y(n234) );
  AO22X1_HVT U240 ( .A1(conv_weight_box[7]), .A2(n356), .A3(conv_weight_box[3]), .A4(n357), .Y(n235) );
  AO22X1_HVT U241 ( .A1(n368), .A2(conv_weight_box[127]), .A3(
        conv_weight_box[95]), .A4(n369), .Y(n236) );
  AO22X1_HVT U242 ( .A1(n366), .A2(conv_weight_box[63]), .A3(
        conv_weight_box[111]), .A4(n367), .Y(n237) );
  AO22X1_HVT U243 ( .A1(n365), .A2(conv_weight_box[143]), .A3(
        conv_weight_box[159]), .A4(n364), .Y(n238) );
  OR3X1_HVT U244 ( .A1(n236), .A2(n237), .A3(n238), .Y(n239) );
  AO22X1_HVT U245 ( .A1(conv_weight_box[191]), .A2(n362), .A3(
        conv_weight_box[31]), .A4(n363), .Y(n240) );
  AO22X1_HVT U246 ( .A1(conv_weight_box[175]), .A2(n360), .A3(
        conv_weight_box[47]), .A4(n361), .Y(n241) );
  OR3X1_HVT U247 ( .A1(n239), .A2(n240), .A3(n241), .Y(n242) );
  AO22X1_HVT U248 ( .A1(n368), .A2(conv_weight_box[123]), .A3(
        conv_weight_box[91]), .A4(n369), .Y(n243) );
  AO22X1_HVT U249 ( .A1(n366), .A2(conv_weight_box[59]), .A3(
        conv_weight_box[107]), .A4(n367), .Y(n244) );
  AO22X1_HVT U250 ( .A1(n365), .A2(conv_weight_box[139]), .A3(
        conv_weight_box[155]), .A4(n364), .Y(n245) );
  OR3X1_HVT U251 ( .A1(n243), .A2(n244), .A3(n245), .Y(n246) );
  AO22X1_HVT U252 ( .A1(conv_weight_box[187]), .A2(n362), .A3(
        conv_weight_box[27]), .A4(n363), .Y(n247) );
  AO22X1_HVT U253 ( .A1(conv_weight_box[171]), .A2(n360), .A3(
        conv_weight_box[43]), .A4(n361), .Y(n248) );
  OR3X1_HVT U254 ( .A1(n246), .A2(n247), .A3(n248), .Y(n249) );
  AO22X1_HVT U255 ( .A1(n371), .A2(n242), .A3(n370), .A4(n249), .Y(n250) );
  NOR4X0_HVT U256 ( .A1(n233), .A2(n234), .A3(n235), .A4(n250), .Y(n251) );
  NAND3X0_HVT U257 ( .A1(n221), .A2(n232), .A3(n251), .Y(n252) );
  AO22X1_HVT U258 ( .A1(conv_weight_box[11]), .A2(n374), .A3(
        conv_weight_box[15]), .A4(n375), .Y(n253) );
  AO22X1_HVT U259 ( .A1(conv_weight_box[87]), .A2(n376), .A3(
        conv_weight_box[83]), .A4(n377), .Y(n254) );
  AO22X1_HVT U260 ( .A1(conv_weight_box[23]), .A2(n378), .A3(
        conv_weight_box[75]), .A4(n379), .Y(n255) );
  AO22X1_HVT U261 ( .A1(conv_weight_box[71]), .A2(n380), .A3(
        conv_weight_box[67]), .A4(n381), .Y(n256) );
  NOR4X0_HVT U262 ( .A1(n253), .A2(n254), .A3(n255), .A4(n256), .Y(n257) );
  AO22X1_HVT U263 ( .A1(conv_weight_box[99]), .A2(n397), .A3(
        conv_weight_box[115]), .A4(n395), .Y(n258) );
  AO22X1_HVT U264 ( .A1(conv_weight_box[35]), .A2(n391), .A3(
        conv_weight_box[51]), .A4(n389), .Y(n259) );
  AO22X1_HVT U265 ( .A1(conv_weight_box[179]), .A2(n388), .A3(
        conv_weight_box[195]), .A4(n390), .Y(n260) );
  AO22X1_HVT U266 ( .A1(conv_weight_box[163]), .A2(n392), .A3(
        conv_weight_box[147]), .A4(n393), .Y(n261) );
  NOR4X0_HVT U267 ( .A1(n258), .A2(n259), .A3(n260), .A4(n261), .Y(n262) );
  AO22X1_HVT U268 ( .A1(n397), .A2(conv_weight_box[103]), .A3(n395), .A4(
        conv_weight_box[119]), .Y(n263) );
  AO22X1_HVT U269 ( .A1(n391), .A2(conv_weight_box[39]), .A3(n389), .A4(
        conv_weight_box[55]), .Y(n264) );
  AO22X1_HVT U270 ( .A1(n388), .A2(conv_weight_box[183]), .A3(n390), .A4(
        conv_weight_box[199]), .Y(n265) );
  AO22X1_HVT U271 ( .A1(n392), .A2(conv_weight_box[167]), .A3(n393), .A4(
        conv_weight_box[151]), .Y(n266) );
  NOR4X0_HVT U272 ( .A1(n263), .A2(n264), .A3(n265), .A4(n266), .Y(n267) );
  OA22X1_HVT U273 ( .A1(n262), .A2(n372), .A3(n267), .A4(n373), .Y(n268) );
  AO22X1_HVT U274 ( .A1(conv_weight_box[79]), .A2(n386), .A3(
        conv_weight_box[131]), .A4(n387), .Y(n269) );
  AO22X1_HVT U275 ( .A1(conv_weight_box[135]), .A2(n382), .A3(
        conv_weight_box[19]), .A4(n383), .Y(n270) );
  AO22X1_HVT U276 ( .A1(conv_weight_box[7]), .A2(n384), .A3(conv_weight_box[3]), .A4(n385), .Y(n271) );
  AO22X1_HVT U277 ( .A1(n396), .A2(conv_weight_box[127]), .A3(n397), .A4(
        conv_weight_box[95]), .Y(n272) );
  AO22X1_HVT U278 ( .A1(n394), .A2(conv_weight_box[63]), .A3(n395), .A4(
        conv_weight_box[111]), .Y(n273) );
  AO22X1_HVT U279 ( .A1(n392), .A2(conv_weight_box[159]), .A3(n393), .A4(
        conv_weight_box[143]), .Y(n274) );
  OR3X1_HVT U280 ( .A1(n272), .A2(n273), .A3(n274), .Y(n275) );
  AO22X1_HVT U281 ( .A1(n391), .A2(conv_weight_box[31]), .A3(n390), .A4(
        conv_weight_box[191]), .Y(n276) );
  AO22X1_HVT U282 ( .A1(n389), .A2(conv_weight_box[47]), .A3(n388), .A4(
        conv_weight_box[175]), .Y(n277) );
  OR3X1_HVT U283 ( .A1(n275), .A2(n276), .A3(n277), .Y(n278) );
  AO22X1_HVT U284 ( .A1(n396), .A2(conv_weight_box[123]), .A3(n397), .A4(
        conv_weight_box[91]), .Y(n279) );
  AO22X1_HVT U285 ( .A1(n394), .A2(conv_weight_box[59]), .A3(n395), .A4(
        conv_weight_box[107]), .Y(n280) );
  AO22X1_HVT U286 ( .A1(n392), .A2(conv_weight_box[155]), .A3(n393), .A4(
        conv_weight_box[139]), .Y(n281) );
  OR3X1_HVT U287 ( .A1(n279), .A2(n280), .A3(n281), .Y(n282) );
  AO22X1_HVT U288 ( .A1(n391), .A2(conv_weight_box[27]), .A3(n390), .A4(
        conv_weight_box[187]), .Y(n283) );
  AO22X1_HVT U289 ( .A1(n389), .A2(conv_weight_box[43]), .A3(n388), .A4(
        conv_weight_box[171]), .Y(n284) );
  OR3X1_HVT U290 ( .A1(n282), .A2(n283), .A3(n284), .Y(n285) );
  AO22X1_HVT U291 ( .A1(n399), .A2(n278), .A3(n398), .A4(n285), .Y(n286) );
  NOR4X0_HVT U292 ( .A1(n269), .A2(n270), .A3(n271), .A4(n286), .Y(n287) );
  NAND3X0_HVT U293 ( .A1(n257), .A2(n268), .A3(n287), .Y(n288) );
  AO22X1_HVT U294 ( .A1(n401), .A2(n252), .A3(n400), .A4(n288), .Y(net19483)
         );
  INVX4_HVT U295 ( .A(srstn), .Y(n305) );
  INVX1_HVT U296 ( .A(n316), .Y(n289) );
  NAND2X0_HVT U297 ( .A1(load_conv2_bias1_enable), .A2(n317), .Y(n319) );
  INVX1_HVT U298 ( .A(n372), .Y(n343) );
  INVX1_HVT U299 ( .A(n344), .Y(n331) );
  INVX0_HVT U300 ( .A(mode[1]), .Y(n315) );
  INVX1_HVT U301 ( .A(n316), .Y(n290) );
  INVX0_HVT U302 ( .A(n319), .Y(n308) );
  AOI22X1_HVT U303 ( .A1(n317), .A2(load_conv2_bias0_enable), .A3(mode[0]), 
        .A4(n315), .Y(n316) );
  NOR2X1_HVT U304 ( .A1(load_conv1_bias_enable), .A2(n320), .Y(n401) );
  INVX0_HVT U305 ( .A(n345), .Y(n328) );
  INVX0_HVT U306 ( .A(n373), .Y(n340) );
  OR2X1_HVT U307 ( .A1(n315), .A2(mode[0]), .Y(n332) );
  INVX1_HVT U308 ( .A(n305), .Y(n292) );
  INVX1_HVT U309 ( .A(n305), .Y(n300) );
  INVX1_HVT U310 ( .A(n319), .Y(n291) );
  INVX2_HVT U311 ( .A(n292), .Y(n293) );
  INVX2_HVT U312 ( .A(n292), .Y(n294) );
  INVX2_HVT U313 ( .A(n292), .Y(n295) );
  INVX2_HVT U314 ( .A(n300), .Y(n296) );
  INVX2_HVT U315 ( .A(n292), .Y(n297) );
  INVX2_HVT U316 ( .A(n292), .Y(n298) );
  INVX2_HVT U317 ( .A(n300), .Y(n299) );
  INVX2_HVT U318 ( .A(n300), .Y(n301) );
  INVX2_HVT U319 ( .A(n300), .Y(n302) );
  INVX2_HVT U320 ( .A(n300), .Y(n303) );
  INVX2_HVT U321 ( .A(n300), .Y(n306) );
  INVX2_HVT U322 ( .A(n319), .Y(n307) );
  INVX2_HVT U323 ( .A(n319), .Y(n309) );
  INVX2_HVT U324 ( .A(n319), .Y(n310) );
  INVX2_HVT U325 ( .A(n316), .Y(n311) );
  INVX2_HVT U326 ( .A(n316), .Y(n312) );
  INVX2_HVT U327 ( .A(n316), .Y(n313) );
  INVX1_HVT U328 ( .A(n332), .Y(n317) );
  AND2X1_HVT U329 ( .A1(set_4_), .A2(n339), .Y(n396) );
  AND2X1_HVT U330 ( .A1(set_5_), .A2(n339), .Y(n394) );
  INVX1_HVT U331 ( .A(set_0_), .Y(n341) );
  INVX1_HVT U332 ( .A(set_1_), .Y(n333) );
  INVX1_HVT U333 ( .A(set_4_), .Y(n338) );
  INVX1_HVT U334 ( .A(set_5_), .Y(n342) );
  AND3X1_HVT U335 ( .A1(set_5_), .A2(set_3_), .A3(n337), .Y(n391) );
  AND3X1_HVT U336 ( .A1(set_2_), .A2(set_5_), .A3(n336), .Y(n389) );
  AND3X1_HVT U337 ( .A1(set_2_), .A2(set_4_), .A3(n336), .Y(n395) );
  INVX1_HVT U338 ( .A(set_3_), .Y(n336) );
  AND3X1_HVT U339 ( .A1(set_3_), .A2(set_4_), .A3(n337), .Y(n397) );
  INVX1_HVT U340 ( .A(set_2_), .Y(n337) );
  AND2X1_HVT U341 ( .A1(conv1_bias_set_4_), .A2(n327), .Y(n368) );
  AND2X1_HVT U342 ( .A1(conv1_bias_set_5_), .A2(n327), .Y(n366) );
  INVX1_HVT U343 ( .A(conv1_bias_set_0_), .Y(n329) );
  INVX1_HVT U344 ( .A(conv1_bias_set_1_), .Y(n321) );
  INVX1_HVT U345 ( .A(conv1_bias_set_4_), .Y(n326) );
  INVX1_HVT U346 ( .A(conv1_bias_set_5_), .Y(n330) );
  AND3X1_HVT U347 ( .A1(conv1_bias_set_5_), .A2(conv1_bias_set_3_), .A3(n325), 
        .Y(n363) );
  AND3X1_HVT U348 ( .A1(conv1_bias_set_2_), .A2(conv1_bias_set_5_), .A3(n324), 
        .Y(n361) );
  AND3X1_HVT U349 ( .A1(conv1_bias_set_2_), .A2(conv1_bias_set_4_), .A3(n324), 
        .Y(n367) );
  INVX1_HVT U350 ( .A(conv1_bias_set_3_), .Y(n324) );
  AND3X1_HVT U351 ( .A1(conv1_bias_set_3_), .A2(conv1_bias_set_4_), .A3(n325), 
        .Y(n369) );
  INVX1_HVT U352 ( .A(conv1_bias_set_2_), .Y(n325) );
  NAND2X0_HVT U353 ( .A1(srstn), .A2(n314), .Y(net19275) );
  INVX1_HVT U354 ( .A(load_conv2_bias0_enable), .Y(n318) );
  NAND2X0_HVT U355 ( .A1(mode[0]), .A2(n315), .Y(n320) );
  AO221X1_HVT U356 ( .A1(n317), .A2(n318), .A3(n332), .A4(n320), .A5(n401), 
        .Y(n314) );
  AND2X1_HVT U357 ( .A1(delay_weight[99]), .A2(n313), .Y(net19121) );
  AND2X1_HVT U358 ( .A1(delay_weight[98]), .A2(n289), .Y(net19124) );
  AND2X1_HVT U359 ( .A1(delay_weight[97]), .A2(n313), .Y(net19125) );
  AND2X1_HVT U360 ( .A1(delay_weight[96]), .A2(n312), .Y(net19126) );
  AND2X1_HVT U361 ( .A1(delay_weight[95]), .A2(n311), .Y(net19127) );
  AND2X1_HVT U362 ( .A1(delay_weight[94]), .A2(n312), .Y(net19128) );
  AND2X1_HVT U363 ( .A1(delay_weight[93]), .A2(n290), .Y(net19129) );
  AND2X1_HVT U364 ( .A1(delay_weight[92]), .A2(n312), .Y(net19130) );
  AND2X1_HVT U365 ( .A1(delay_weight[91]), .A2(n311), .Y(net19131) );
  AND2X1_HVT U366 ( .A1(delay_weight[90]), .A2(n311), .Y(net19132) );
  AND2X1_HVT U367 ( .A1(delay_weight[89]), .A2(n312), .Y(net19140) );
  AND2X1_HVT U368 ( .A1(delay_weight[88]), .A2(n313), .Y(net19141) );
  AND2X1_HVT U369 ( .A1(delay_weight[87]), .A2(n312), .Y(net19142) );
  AND2X1_HVT U370 ( .A1(delay_weight[86]), .A2(n313), .Y(net19143) );
  AND2X1_HVT U371 ( .A1(delay_weight[85]), .A2(n289), .Y(net19144) );
  AND2X1_HVT U372 ( .A1(delay_weight[84]), .A2(n311), .Y(net19145) );
  AND2X1_HVT U373 ( .A1(delay_weight[83]), .A2(n311), .Y(net19146) );
  AND2X1_HVT U374 ( .A1(delay_weight[82]), .A2(n311), .Y(net19147) );
  AND2X1_HVT U375 ( .A1(delay_weight[81]), .A2(n289), .Y(net19148) );
  AND2X1_HVT U376 ( .A1(delay_weight[80]), .A2(n312), .Y(net19149) );
  AND2X1_HVT U377 ( .A1(delay_weight[79]), .A2(n313), .Y(net19157) );
  AND2X1_HVT U378 ( .A1(delay_weight[78]), .A2(n313), .Y(net19158) );
  AND2X1_HVT U379 ( .A1(delay_weight[77]), .A2(n289), .Y(net19159) );
  AND2X1_HVT U380 ( .A1(delay_weight[76]), .A2(n312), .Y(net19160) );
  AND2X1_HVT U381 ( .A1(delay_weight[75]), .A2(n311), .Y(net19161) );
  AND2X1_HVT U382 ( .A1(delay_weight[74]), .A2(n290), .Y(net19162) );
  AND2X1_HVT U383 ( .A1(delay_weight[73]), .A2(n290), .Y(net19163) );
  AND2X1_HVT U384 ( .A1(delay_weight[72]), .A2(n313), .Y(net19164) );
  AND2X1_HVT U385 ( .A1(delay_weight[71]), .A2(n313), .Y(net19165) );
  AND2X1_HVT U386 ( .A1(delay_weight[70]), .A2(n313), .Y(net19166) );
  AND2X1_HVT U387 ( .A1(delay_weight[69]), .A2(n289), .Y(net19174) );
  AND2X1_HVT U388 ( .A1(delay_weight[68]), .A2(n311), .Y(net19175) );
  AND2X1_HVT U389 ( .A1(delay_weight[67]), .A2(n290), .Y(net19176) );
  AND2X1_HVT U390 ( .A1(delay_weight[66]), .A2(n312), .Y(net19177) );
  AND2X1_HVT U391 ( .A1(delay_weight[65]), .A2(n311), .Y(net19178) );
  AND2X1_HVT U392 ( .A1(delay_weight[64]), .A2(n311), .Y(net19179) );
  AND2X1_HVT U393 ( .A1(delay_weight[63]), .A2(n313), .Y(net19180) );
  AND2X1_HVT U394 ( .A1(delay_weight[62]), .A2(n312), .Y(net19181) );
  AND2X1_HVT U395 ( .A1(delay_weight[61]), .A2(n289), .Y(net19182) );
  AND2X1_HVT U396 ( .A1(delay_weight[60]), .A2(n312), .Y(net19183) );
  AND2X1_HVT U397 ( .A1(delay_weight[59]), .A2(n313), .Y(net19191) );
  AND2X1_HVT U398 ( .A1(delay_weight[58]), .A2(n312), .Y(net19192) );
  AND2X1_HVT U399 ( .A1(delay_weight[57]), .A2(n290), .Y(net19193) );
  AND2X1_HVT U400 ( .A1(delay_weight[56]), .A2(n311), .Y(net19194) );
  AND2X1_HVT U401 ( .A1(delay_weight[55]), .A2(n290), .Y(net19195) );
  AND2X1_HVT U402 ( .A1(delay_weight[54]), .A2(n311), .Y(net19196) );
  AND2X1_HVT U403 ( .A1(delay_weight[53]), .A2(n289), .Y(net19197) );
  AND2X1_HVT U404 ( .A1(delay_weight[52]), .A2(n313), .Y(net19198) );
  AND2X1_HVT U405 ( .A1(delay_weight[51]), .A2(n312), .Y(net19199) );
  AND2X1_HVT U406 ( .A1(delay_weight[50]), .A2(n289), .Y(net19200) );
  AND2X1_HVT U407 ( .A1(delay_weight[49]), .A2(n289), .Y(net19208) );
  AND2X1_HVT U408 ( .A1(delay_weight[48]), .A2(n311), .Y(net19209) );
  AND2X1_HVT U409 ( .A1(delay_weight[47]), .A2(n312), .Y(net19210) );
  AND2X1_HVT U410 ( .A1(delay_weight[46]), .A2(n311), .Y(net19211) );
  AND2X1_HVT U411 ( .A1(delay_weight[45]), .A2(n289), .Y(net19212) );
  AND2X1_HVT U412 ( .A1(delay_weight[44]), .A2(n313), .Y(net19213) );
  AND2X1_HVT U413 ( .A1(delay_weight[43]), .A2(n290), .Y(net19214) );
  AND2X1_HVT U414 ( .A1(delay_weight[42]), .A2(n313), .Y(net19215) );
  AND2X1_HVT U415 ( .A1(delay_weight[41]), .A2(n313), .Y(net19216) );
  AND2X1_HVT U416 ( .A1(delay_weight[40]), .A2(n312), .Y(net19217) );
  AND2X1_HVT U417 ( .A1(delay_weight[39]), .A2(n311), .Y(net19225) );
  AND2X1_HVT U418 ( .A1(delay_weight[38]), .A2(n311), .Y(net19226) );
  AND2X1_HVT U419 ( .A1(delay_weight[37]), .A2(n290), .Y(net19227) );
  AND2X1_HVT U420 ( .A1(delay_weight[36]), .A2(n313), .Y(net19228) );
  AND2X1_HVT U421 ( .A1(delay_weight[35]), .A2(n312), .Y(net19229) );
  AND2X1_HVT U422 ( .A1(delay_weight[34]), .A2(n313), .Y(net19230) );
  AND2X1_HVT U423 ( .A1(delay_weight[33]), .A2(n289), .Y(net19231) );
  AND2X1_HVT U424 ( .A1(delay_weight[32]), .A2(n313), .Y(net19232) );
  AND2X1_HVT U425 ( .A1(delay_weight[31]), .A2(n290), .Y(net19233) );
  AND2X1_HVT U426 ( .A1(delay_weight[30]), .A2(n312), .Y(net19234) );
  AND2X1_HVT U427 ( .A1(delay_weight[29]), .A2(n290), .Y(net19242) );
  AND2X1_HVT U428 ( .A1(delay_weight[28]), .A2(n311), .Y(net19243) );
  AND2X1_HVT U429 ( .A1(delay_weight[27]), .A2(n313), .Y(net19244) );
  AND2X1_HVT U430 ( .A1(delay_weight[26]), .A2(n289), .Y(net19245) );
  AND2X1_HVT U431 ( .A1(delay_weight[25]), .A2(n289), .Y(net19246) );
  AND2X1_HVT U432 ( .A1(delay_weight[24]), .A2(n312), .Y(net19247) );
  AND2X1_HVT U433 ( .A1(delay_weight[23]), .A2(n311), .Y(net19248) );
  AND2X1_HVT U434 ( .A1(delay_weight[22]), .A2(n312), .Y(net19249) );
  AND2X1_HVT U435 ( .A1(delay_weight[21]), .A2(n290), .Y(net19250) );
  AND2X1_HVT U436 ( .A1(delay_weight[20]), .A2(n312), .Y(net19251) );
  AND2X1_HVT U437 ( .A1(delay_weight[19]), .A2(n290), .Y(net19259) );
  AND2X1_HVT U438 ( .A1(delay_weight[18]), .A2(n311), .Y(net19260) );
  AND2X1_HVT U439 ( .A1(delay_weight[17]), .A2(n312), .Y(net19261) );
  AND2X1_HVT U440 ( .A1(delay_weight[16]), .A2(n313), .Y(net19262) );
  AND2X1_HVT U441 ( .A1(delay_weight[15]), .A2(n312), .Y(net19263) );
  AND2X1_HVT U442 ( .A1(delay_weight[14]), .A2(n313), .Y(net19264) );
  AND2X1_HVT U443 ( .A1(delay_weight[13]), .A2(n289), .Y(net19265) );
  AND2X1_HVT U444 ( .A1(delay_weight[12]), .A2(n311), .Y(net19266) );
  AND2X1_HVT U445 ( .A1(delay_weight[11]), .A2(n311), .Y(net19267) );
  AND2X1_HVT U446 ( .A1(delay_weight[10]), .A2(n311), .Y(net19268) );
  AND2X1_HVT U447 ( .A1(delay_weight[9]), .A2(n289), .Y(net19276) );
  AND2X1_HVT U448 ( .A1(delay_weight[8]), .A2(n312), .Y(net19277) );
  AND2X1_HVT U449 ( .A1(delay_weight[7]), .A2(n290), .Y(net19278) );
  AND2X1_HVT U450 ( .A1(delay_weight[6]), .A2(n313), .Y(net19279) );
  AND2X1_HVT U451 ( .A1(delay_weight[5]), .A2(n289), .Y(net19280) );
  AND2X1_HVT U452 ( .A1(delay_weight[4]), .A2(n312), .Y(net19281) );
  AND2X1_HVT U453 ( .A1(delay_weight[3]), .A2(n311), .Y(net19282) );
  AND2X1_HVT U454 ( .A1(delay_weight[2]), .A2(n290), .Y(net19283) );
  AND2X1_HVT U455 ( .A1(delay_weight[1]), .A2(n290), .Y(net19284) );
  AND2X1_HVT U456 ( .A1(delay_weight[0]), .A2(n313), .Y(net19285) );
  AO21X1_HVT U457 ( .A1(n291), .A2(n318), .A3(n305), .Y(net19453) );
  AND2X1_HVT U458 ( .A1(delay_weight[99]), .A2(n309), .Y(net19301) );
  AND2X1_HVT U459 ( .A1(delay_weight[98]), .A2(n309), .Y(net19302) );
  AND2X1_HVT U460 ( .A1(delay_weight[97]), .A2(n308), .Y(net19303) );
  AND2X1_HVT U461 ( .A1(delay_weight[96]), .A2(n310), .Y(net19304) );
  AND2X1_HVT U462 ( .A1(delay_weight[95]), .A2(n291), .Y(net19305) );
  AND2X1_HVT U463 ( .A1(delay_weight[94]), .A2(n307), .Y(net19306) );
  AND2X1_HVT U464 ( .A1(delay_weight[93]), .A2(n310), .Y(net19307) );
  AND2X1_HVT U465 ( .A1(delay_weight[92]), .A2(n307), .Y(net19308) );
  AND2X1_HVT U466 ( .A1(delay_weight[91]), .A2(n310), .Y(net19309) );
  AND2X1_HVT U467 ( .A1(delay_weight[90]), .A2(n310), .Y(net19310) );
  AND2X1_HVT U468 ( .A1(delay_weight[89]), .A2(n310), .Y(net19318) );
  AND2X1_HVT U469 ( .A1(delay_weight[88]), .A2(n307), .Y(net19319) );
  AND2X1_HVT U470 ( .A1(delay_weight[87]), .A2(n307), .Y(net19320) );
  AND2X1_HVT U471 ( .A1(delay_weight[86]), .A2(n291), .Y(net19321) );
  AND2X1_HVT U472 ( .A1(delay_weight[85]), .A2(n309), .Y(net19322) );
  AND2X1_HVT U473 ( .A1(delay_weight[84]), .A2(n307), .Y(net19323) );
  AND2X1_HVT U474 ( .A1(delay_weight[83]), .A2(n309), .Y(net19324) );
  AND2X1_HVT U475 ( .A1(delay_weight[82]), .A2(n309), .Y(net19325) );
  AND2X1_HVT U476 ( .A1(delay_weight[81]), .A2(n307), .Y(net19326) );
  AND2X1_HVT U477 ( .A1(delay_weight[80]), .A2(n307), .Y(net19327) );
  AND2X1_HVT U478 ( .A1(delay_weight[79]), .A2(n309), .Y(net19335) );
  AND2X1_HVT U479 ( .A1(delay_weight[78]), .A2(n308), .Y(net19336) );
  AND2X1_HVT U480 ( .A1(delay_weight[77]), .A2(n291), .Y(net19337) );
  AND2X1_HVT U481 ( .A1(delay_weight[76]), .A2(n308), .Y(net19338) );
  AND2X1_HVT U482 ( .A1(delay_weight[75]), .A2(n308), .Y(net19339) );
  AND2X1_HVT U483 ( .A1(delay_weight[74]), .A2(n310), .Y(net19340) );
  AND2X1_HVT U484 ( .A1(delay_weight[73]), .A2(n307), .Y(net19341) );
  AND2X1_HVT U485 ( .A1(delay_weight[72]), .A2(n308), .Y(net19342) );
  AND2X1_HVT U486 ( .A1(delay_weight[71]), .A2(n309), .Y(net19343) );
  AND2X1_HVT U487 ( .A1(delay_weight[70]), .A2(n308), .Y(net19344) );
  AND2X1_HVT U488 ( .A1(delay_weight[69]), .A2(n308), .Y(net19352) );
  AND2X1_HVT U489 ( .A1(delay_weight[68]), .A2(n291), .Y(net19353) );
  AND2X1_HVT U490 ( .A1(delay_weight[67]), .A2(n310), .Y(net19354) );
  AND2X1_HVT U491 ( .A1(delay_weight[66]), .A2(n309), .Y(net19355) );
  AND2X1_HVT U492 ( .A1(delay_weight[65]), .A2(n307), .Y(net19356) );
  AND2X1_HVT U493 ( .A1(delay_weight[64]), .A2(n310), .Y(net19357) );
  AND2X1_HVT U494 ( .A1(delay_weight[63]), .A2(n309), .Y(net19358) );
  AND2X1_HVT U495 ( .A1(delay_weight[62]), .A2(n310), .Y(net19359) );
  AND2X1_HVT U496 ( .A1(delay_weight[61]), .A2(n310), .Y(net19360) );
  AND2X1_HVT U497 ( .A1(delay_weight[60]), .A2(n308), .Y(net19361) );
  AND2X1_HVT U498 ( .A1(delay_weight[59]), .A2(n291), .Y(net19369) );
  AND2X1_HVT U499 ( .A1(delay_weight[58]), .A2(n309), .Y(net19370) );
  AND2X1_HVT U500 ( .A1(delay_weight[57]), .A2(n310), .Y(net19371) );
  AND2X1_HVT U501 ( .A1(delay_weight[56]), .A2(n308), .Y(net19372) );
  AND2X1_HVT U502 ( .A1(delay_weight[55]), .A2(n308), .Y(net19373) );
  AND2X1_HVT U503 ( .A1(delay_weight[54]), .A2(n310), .Y(net19374) );
  AND2X1_HVT U504 ( .A1(delay_weight[53]), .A2(n307), .Y(net19375) );
  AND2X1_HVT U505 ( .A1(delay_weight[52]), .A2(n309), .Y(net19376) );
  AND2X1_HVT U506 ( .A1(delay_weight[51]), .A2(n308), .Y(net19377) );
  AND2X1_HVT U507 ( .A1(delay_weight[50]), .A2(n291), .Y(net19378) );
  AND2X1_HVT U508 ( .A1(delay_weight[49]), .A2(n307), .Y(net19386) );
  AND2X1_HVT U509 ( .A1(delay_weight[48]), .A2(n307), .Y(net19387) );
  AND2X1_HVT U510 ( .A1(delay_weight[47]), .A2(n309), .Y(net19388) );
  AND2X1_HVT U511 ( .A1(delay_weight[46]), .A2(n307), .Y(net19389) );
  AND2X1_HVT U512 ( .A1(delay_weight[45]), .A2(n309), .Y(net19390) );
  AND2X1_HVT U513 ( .A1(delay_weight[44]), .A2(n308), .Y(net19391) );
  AND2X1_HVT U514 ( .A1(delay_weight[43]), .A2(n307), .Y(net19392) );
  AND2X1_HVT U515 ( .A1(delay_weight[42]), .A2(n307), .Y(net19393) );
  AND2X1_HVT U516 ( .A1(delay_weight[41]), .A2(n291), .Y(net19394) );
  AND2X1_HVT U517 ( .A1(delay_weight[40]), .A2(n310), .Y(net19395) );
  AND2X1_HVT U518 ( .A1(delay_weight[39]), .A2(n308), .Y(net19403) );
  AND2X1_HVT U519 ( .A1(delay_weight[38]), .A2(n310), .Y(net19404) );
  AND2X1_HVT U520 ( .A1(delay_weight[37]), .A2(n309), .Y(net19405) );
  AND2X1_HVT U521 ( .A1(delay_weight[36]), .A2(n310), .Y(net19406) );
  AND2X1_HVT U522 ( .A1(delay_weight[35]), .A2(n309), .Y(net19407) );
  AND2X1_HVT U523 ( .A1(delay_weight[34]), .A2(n310), .Y(net19408) );
  AND2X1_HVT U524 ( .A1(delay_weight[33]), .A2(n309), .Y(net19409) );
  AND2X1_HVT U525 ( .A1(delay_weight[32]), .A2(n291), .Y(net19410) );
  AND2X1_HVT U526 ( .A1(delay_weight[31]), .A2(n309), .Y(net19411) );
  AND2X1_HVT U527 ( .A1(delay_weight[30]), .A2(n308), .Y(net19412) );
  AND2X1_HVT U528 ( .A1(delay_weight[29]), .A2(n307), .Y(net19420) );
  AND2X1_HVT U529 ( .A1(delay_weight[28]), .A2(n308), .Y(net19421) );
  AND2X1_HVT U530 ( .A1(delay_weight[27]), .A2(n307), .Y(net19422) );
  AND2X1_HVT U531 ( .A1(delay_weight[26]), .A2(n310), .Y(net19423) );
  AND2X1_HVT U532 ( .A1(delay_weight[25]), .A2(n309), .Y(net19424) );
  AND2X1_HVT U533 ( .A1(delay_weight[24]), .A2(n310), .Y(net19425) );
  AND2X1_HVT U534 ( .A1(delay_weight[23]), .A2(n291), .Y(net19426) );
  AND2X1_HVT U535 ( .A1(delay_weight[22]), .A2(n307), .Y(net19427) );
  AND2X1_HVT U536 ( .A1(delay_weight[21]), .A2(n291), .Y(net19428) );
  AND2X1_HVT U537 ( .A1(delay_weight[20]), .A2(n309), .Y(net19429) );
  AND2X1_HVT U538 ( .A1(delay_weight[19]), .A2(n310), .Y(net19437) );
  AND2X1_HVT U539 ( .A1(delay_weight[18]), .A2(n308), .Y(net19438) );
  AND2X1_HVT U540 ( .A1(delay_weight[17]), .A2(n307), .Y(net19439) );
  AND2X1_HVT U541 ( .A1(delay_weight[16]), .A2(n307), .Y(net19440) );
  AND2X1_HVT U542 ( .A1(delay_weight[15]), .A2(n307), .Y(net19441) );
  AND2X1_HVT U543 ( .A1(delay_weight[14]), .A2(n291), .Y(net19442) );
  AND2X1_HVT U544 ( .A1(delay_weight[13]), .A2(n310), .Y(net19443) );
  AND2X1_HVT U545 ( .A1(delay_weight[12]), .A2(n291), .Y(net19444) );
  AND2X1_HVT U546 ( .A1(delay_weight[11]), .A2(n310), .Y(net19445) );
  AND2X1_HVT U547 ( .A1(delay_weight[10]), .A2(n309), .Y(net19446) );
  AND2X1_HVT U548 ( .A1(delay_weight[9]), .A2(n309), .Y(net19454) );
  AND2X1_HVT U549 ( .A1(delay_weight[8]), .A2(n309), .Y(net19455) );
  AND2X1_HVT U550 ( .A1(delay_weight[7]), .A2(n310), .Y(net19456) );
  AND2X1_HVT U551 ( .A1(delay_weight[6]), .A2(n308), .Y(net19457) );
  AND2X1_HVT U552 ( .A1(delay_weight[5]), .A2(n291), .Y(net19458) );
  AND2X1_HVT U553 ( .A1(delay_weight[4]), .A2(n309), .Y(net19459) );
  AND2X1_HVT U554 ( .A1(delay_weight[3]), .A2(n291), .Y(net19460) );
  AND2X1_HVT U555 ( .A1(delay_weight[2]), .A2(n307), .Y(net19461) );
  AND2X1_HVT U556 ( .A1(delay_weight[1]), .A2(n307), .Y(net19462) );
  AND2X1_HVT U557 ( .A1(delay_weight[0]), .A2(n310), .Y(net19463) );
  NAND3X0_HVT U558 ( .A1(srstn), .A2(n320), .A3(n332), .Y(net19477) );
  AND4X1_HVT U559 ( .A1(conv1_bias_set_2_), .A2(n330), .A3(n324), .A4(n326), 
        .Y(n360) );
  AND4X1_HVT U560 ( .A1(n330), .A2(n325), .A3(n324), .A4(n326), .Y(n362) );
  AND4X1_HVT U561 ( .A1(conv1_bias_set_2_), .A2(conv1_bias_set_3_), .A3(n330), 
        .A4(n326), .Y(n365) );
  AND4X1_HVT U562 ( .A1(conv1_bias_set_3_), .A2(n330), .A3(n325), .A4(n326), 
        .Y(n364) );
  NAND2X0_HVT U563 ( .A1(n321), .A2(n329), .Y(n345) );
  NAND2X0_HVT U564 ( .A1(conv1_bias_set_0_), .A2(n321), .Y(n344) );
  AND2X1_HVT U565 ( .A1(conv1_bias_set_1_), .A2(n329), .Y(n371) );
  AND4X1_HVT U566 ( .A1(n371), .A2(conv1_bias_set_5_), .A3(conv1_bias_set_2_), 
        .A4(conv1_bias_set_3_), .Y(n347) );
  AND3X1_HVT U567 ( .A1(conv1_bias_set_5_), .A2(conv1_bias_set_2_), .A3(
        conv1_bias_set_3_), .Y(n322) );
  AND3X1_HVT U568 ( .A1(conv1_bias_set_1_), .A2(conv1_bias_set_0_), .A3(n322), 
        .Y(n346) );
  AND4X1_HVT U569 ( .A1(conv1_bias_set_2_), .A2(conv1_bias_set_3_), .A3(
        conv1_bias_set_4_), .A4(n331), .Y(n349) );
  AND4X1_HVT U570 ( .A1(conv1_bias_set_2_), .A2(conv1_bias_set_3_), .A3(
        conv1_bias_set_4_), .A4(n328), .Y(n348) );
  AND3X1_HVT U571 ( .A1(conv1_bias_set_2_), .A2(conv1_bias_set_3_), .A3(
        conv1_bias_set_4_), .Y(n323) );
  AND3X1_HVT U572 ( .A1(conv1_bias_set_1_), .A2(conv1_bias_set_0_), .A3(n323), 
        .Y(n351) );
  AND4X1_HVT U573 ( .A1(conv1_bias_set_5_), .A2(conv1_bias_set_2_), .A3(
        conv1_bias_set_3_), .A4(n328), .Y(n350) );
  AND2X1_HVT U574 ( .A1(n325), .A2(n324), .Y(n327) );
  AND3X1_HVT U575 ( .A1(n366), .A2(n331), .A3(n326), .Y(n353) );
  AND3X1_HVT U576 ( .A1(n366), .A2(n328), .A3(n326), .Y(n352) );
  AND4X1_HVT U577 ( .A1(conv1_bias_set_5_), .A2(conv1_bias_set_2_), .A3(
        conv1_bias_set_3_), .A4(n331), .Y(n355) );
  AND3X1_HVT U578 ( .A1(n368), .A2(n328), .A3(n330), .Y(n354) );
  AND3X1_HVT U579 ( .A1(conv1_bias_set_0_), .A2(conv1_bias_set_5_), .A3(
        conv1_bias_set_4_), .Y(n357) );
  AND3X1_HVT U580 ( .A1(conv1_bias_set_5_), .A2(conv1_bias_set_4_), .A3(n329), 
        .Y(n356) );
  AND3X1_HVT U581 ( .A1(n368), .A2(n331), .A3(n330), .Y(n359) );
  AND4X1_HVT U582 ( .A1(n371), .A2(conv1_bias_set_2_), .A3(conv1_bias_set_3_), 
        .A4(conv1_bias_set_4_), .Y(n358) );
  AND2X1_HVT U583 ( .A1(conv1_bias_set_1_), .A2(conv1_bias_set_0_), .Y(n370)
         );
  NOR3X0_HVT U584 ( .A1(load_conv2_bias1_enable), .A2(load_conv2_bias0_enable), 
        .A3(n332), .Y(n400) );
  AND4X1_HVT U585 ( .A1(n342), .A2(n337), .A3(n336), .A4(n338), .Y(n390) );
  AND4X1_HVT U586 ( .A1(set_2_), .A2(n342), .A3(n336), .A4(n338), .Y(n388) );
  AND4X1_HVT U587 ( .A1(set_2_), .A2(set_3_), .A3(n342), .A4(n338), .Y(n393)
         );
  AND4X1_HVT U588 ( .A1(set_3_), .A2(n342), .A3(n337), .A4(n338), .Y(n392) );
  NAND2X0_HVT U589 ( .A1(n333), .A2(n341), .Y(n373) );
  NAND2X0_HVT U590 ( .A1(set_0_), .A2(n333), .Y(n372) );
  AND2X1_HVT U591 ( .A1(set_1_), .A2(n341), .Y(n399) );
  AND4X1_HVT U592 ( .A1(n399), .A2(set_5_), .A3(set_2_), .A4(set_3_), .Y(n375)
         );
  AND3X1_HVT U593 ( .A1(set_5_), .A2(set_2_), .A3(set_3_), .Y(n334) );
  AND3X1_HVT U594 ( .A1(set_1_), .A2(set_0_), .A3(n334), .Y(n374) );
  AND4X1_HVT U595 ( .A1(set_2_), .A2(set_3_), .A3(set_4_), .A4(n343), .Y(n377)
         );
  AND4X1_HVT U596 ( .A1(set_2_), .A2(set_3_), .A3(set_4_), .A4(n340), .Y(n376)
         );
  AND3X1_HVT U597 ( .A1(set_2_), .A2(set_3_), .A3(set_4_), .Y(n335) );
  AND3X1_HVT U598 ( .A1(set_1_), .A2(set_0_), .A3(n335), .Y(n379) );
  AND4X1_HVT U599 ( .A1(set_5_), .A2(set_2_), .A3(set_3_), .A4(n340), .Y(n378)
         );
  AND2X1_HVT U600 ( .A1(n337), .A2(n336), .Y(n339) );
  AND3X1_HVT U601 ( .A1(n394), .A2(n343), .A3(n338), .Y(n381) );
  AND3X1_HVT U602 ( .A1(n394), .A2(n340), .A3(n338), .Y(n380) );
  AND4X1_HVT U603 ( .A1(set_5_), .A2(set_2_), .A3(set_3_), .A4(n343), .Y(n383)
         );
  AND3X1_HVT U604 ( .A1(n396), .A2(n340), .A3(n342), .Y(n382) );
  AND3X1_HVT U605 ( .A1(set_0_), .A2(set_5_), .A3(set_4_), .Y(n385) );
  AND3X1_HVT U606 ( .A1(set_5_), .A2(set_4_), .A3(n341), .Y(n384) );
  AND3X1_HVT U607 ( .A1(n396), .A2(n343), .A3(n342), .Y(n387) );
  AND4X1_HVT U608 ( .A1(n399), .A2(set_2_), .A3(set_3_), .A4(set_4_), .Y(n386)
         );
  AND2X1_HVT U609 ( .A1(set_1_), .A2(set_0_), .Y(n398) );
endmodule


module multiply_compare ( clk, srstn, mode, channel, conv1_sram_rdata_weight, 
        conv2_sram_rdata_weight, src_window, data_out );
  input [1:0] mode;
  input [4:0] channel;
  input [99:0] conv1_sram_rdata_weight;
  input [99:0] conv2_sram_rdata_weight;
  input [287:0] src_window;
  output [31:0] data_out;
  input clk, srstn;
  wire   N5, N7, N9, DP_OP_425J2_127_3477_n3255, DP_OP_425J2_127_3477_n3110,
         DP_OP_425J2_127_3477_n2918, DP_OP_425J2_127_3477_n2917,
         DP_OP_425J2_127_3477_n2916, DP_OP_425J2_127_3477_n2915,
         DP_OP_425J2_127_3477_n2914, DP_OP_425J2_127_3477_n2913,
         DP_OP_425J2_127_3477_n2912, DP_OP_425J2_127_3477_n2911,
         DP_OP_425J2_127_3477_n2910, DP_OP_425J2_127_3477_n2909,
         DP_OP_425J2_127_3477_n2908, DP_OP_425J2_127_3477_n2907,
         DP_OP_425J2_127_3477_n2906, DP_OP_425J2_127_3477_n2905,
         DP_OP_425J2_127_3477_n2904, DP_OP_425J2_127_3477_n2903,
         DP_OP_425J2_127_3477_n2902, DP_OP_425J2_127_3477_n2901,
         DP_OP_425J2_127_3477_n2900, DP_OP_425J2_127_3477_n2899,
         DP_OP_425J2_127_3477_n2898, DP_OP_425J2_127_3477_n2897,
         DP_OP_425J2_127_3477_n2896, DP_OP_425J2_127_3477_n2895,
         DP_OP_425J2_127_3477_n2894, DP_OP_425J2_127_3477_n2893,
         DP_OP_425J2_127_3477_n2892, DP_OP_425J2_127_3477_n2891,
         DP_OP_425J2_127_3477_n2890, DP_OP_425J2_127_3477_n2889,
         DP_OP_425J2_127_3477_n2888, DP_OP_425J2_127_3477_n2887,
         DP_OP_425J2_127_3477_n2886, DP_OP_425J2_127_3477_n2885,
         DP_OP_425J2_127_3477_n2884, DP_OP_425J2_127_3477_n2883,
         DP_OP_425J2_127_3477_n2882, DP_OP_425J2_127_3477_n2881,
         DP_OP_425J2_127_3477_n2880, DP_OP_425J2_127_3477_n2879,
         DP_OP_425J2_127_3477_n2878, DP_OP_425J2_127_3477_n2877,
         DP_OP_425J2_127_3477_n2876, DP_OP_425J2_127_3477_n2875,
         DP_OP_425J2_127_3477_n2874, DP_OP_425J2_127_3477_n2872,
         DP_OP_425J2_127_3477_n2871, DP_OP_425J2_127_3477_n2870,
         DP_OP_425J2_127_3477_n2869, DP_OP_425J2_127_3477_n2868,
         DP_OP_425J2_127_3477_n2865, DP_OP_425J2_127_3477_n2864,
         DP_OP_425J2_127_3477_n2862, DP_OP_425J2_127_3477_n2861,
         DP_OP_425J2_127_3477_n2860, DP_OP_425J2_127_3477_n2859,
         DP_OP_425J2_127_3477_n2858, DP_OP_425J2_127_3477_n2857,
         DP_OP_425J2_127_3477_n2856, DP_OP_425J2_127_3477_n2855,
         DP_OP_425J2_127_3477_n2854, DP_OP_425J2_127_3477_n2853,
         DP_OP_425J2_127_3477_n2852, DP_OP_425J2_127_3477_n2851,
         DP_OP_425J2_127_3477_n2850, DP_OP_425J2_127_3477_n2849,
         DP_OP_425J2_127_3477_n2848, DP_OP_425J2_127_3477_n2847,
         DP_OP_425J2_127_3477_n2846, DP_OP_425J2_127_3477_n2845,
         DP_OP_425J2_127_3477_n2844, DP_OP_425J2_127_3477_n2843,
         DP_OP_425J2_127_3477_n2842, DP_OP_425J2_127_3477_n2841,
         DP_OP_425J2_127_3477_n2840, DP_OP_425J2_127_3477_n2839,
         DP_OP_425J2_127_3477_n2838, DP_OP_425J2_127_3477_n2837,
         DP_OP_425J2_127_3477_n2836, DP_OP_425J2_127_3477_n2835,
         DP_OP_425J2_127_3477_n2834, DP_OP_425J2_127_3477_n2833,
         DP_OP_425J2_127_3477_n2832, DP_OP_425J2_127_3477_n2831,
         DP_OP_425J2_127_3477_n2830, DP_OP_425J2_127_3477_n2829,
         DP_OP_425J2_127_3477_n2828, DP_OP_425J2_127_3477_n2827,
         DP_OP_425J2_127_3477_n2826, DP_OP_425J2_127_3477_n2823,
         DP_OP_425J2_127_3477_n2821, DP_OP_425J2_127_3477_n2820,
         DP_OP_425J2_127_3477_n2818, DP_OP_425J2_127_3477_n2817,
         DP_OP_425J2_127_3477_n2816, DP_OP_425J2_127_3477_n2815,
         DP_OP_425J2_127_3477_n2814, DP_OP_425J2_127_3477_n2813,
         DP_OP_425J2_127_3477_n2812, DP_OP_425J2_127_3477_n2811,
         DP_OP_425J2_127_3477_n2810, DP_OP_425J2_127_3477_n2809,
         DP_OP_425J2_127_3477_n2808, DP_OP_425J2_127_3477_n2807,
         DP_OP_425J2_127_3477_n2806, DP_OP_425J2_127_3477_n2805,
         DP_OP_425J2_127_3477_n2804, DP_OP_425J2_127_3477_n2803,
         DP_OP_425J2_127_3477_n2802, DP_OP_425J2_127_3477_n2801,
         DP_OP_425J2_127_3477_n2800, DP_OP_425J2_127_3477_n2799,
         DP_OP_425J2_127_3477_n2798, DP_OP_425J2_127_3477_n2797,
         DP_OP_425J2_127_3477_n2796, DP_OP_425J2_127_3477_n2795,
         DP_OP_425J2_127_3477_n2794, DP_OP_425J2_127_3477_n2793,
         DP_OP_425J2_127_3477_n2792, DP_OP_425J2_127_3477_n2791,
         DP_OP_425J2_127_3477_n2790, DP_OP_425J2_127_3477_n2789,
         DP_OP_425J2_127_3477_n2788, DP_OP_425J2_127_3477_n2787,
         DP_OP_425J2_127_3477_n2786, DP_OP_425J2_127_3477_n2785,
         DP_OP_425J2_127_3477_n2783, DP_OP_425J2_127_3477_n2780,
         DP_OP_425J2_127_3477_n2779, DP_OP_425J2_127_3477_n2778,
         DP_OP_425J2_127_3477_n2777, DP_OP_425J2_127_3477_n2774,
         DP_OP_425J2_127_3477_n2773, DP_OP_425J2_127_3477_n2772,
         DP_OP_425J2_127_3477_n2771, DP_OP_425J2_127_3477_n2770,
         DP_OP_425J2_127_3477_n2769, DP_OP_425J2_127_3477_n2768,
         DP_OP_425J2_127_3477_n2767, DP_OP_425J2_127_3477_n2766,
         DP_OP_425J2_127_3477_n2765, DP_OP_425J2_127_3477_n2764,
         DP_OP_425J2_127_3477_n2763, DP_OP_425J2_127_3477_n2762,
         DP_OP_425J2_127_3477_n2761, DP_OP_425J2_127_3477_n2760,
         DP_OP_425J2_127_3477_n2759, DP_OP_425J2_127_3477_n2758,
         DP_OP_425J2_127_3477_n2757, DP_OP_425J2_127_3477_n2756,
         DP_OP_425J2_127_3477_n2755, DP_OP_425J2_127_3477_n2754,
         DP_OP_425J2_127_3477_n2753, DP_OP_425J2_127_3477_n2752,
         DP_OP_425J2_127_3477_n2751, DP_OP_425J2_127_3477_n2750,
         DP_OP_425J2_127_3477_n2749, DP_OP_425J2_127_3477_n2748,
         DP_OP_425J2_127_3477_n2747, DP_OP_425J2_127_3477_n2746,
         DP_OP_425J2_127_3477_n2745, DP_OP_425J2_127_3477_n2744,
         DP_OP_425J2_127_3477_n2743, DP_OP_425J2_127_3477_n2741,
         DP_OP_425J2_127_3477_n2740, DP_OP_425J2_127_3477_n2739,
         DP_OP_425J2_127_3477_n2738, DP_OP_425J2_127_3477_n2735,
         DP_OP_425J2_127_3477_n2734, DP_OP_425J2_127_3477_n2732,
         DP_OP_425J2_127_3477_n2730, DP_OP_425J2_127_3477_n2729,
         DP_OP_425J2_127_3477_n2728, DP_OP_425J2_127_3477_n2727,
         DP_OP_425J2_127_3477_n2726, DP_OP_425J2_127_3477_n2725,
         DP_OP_425J2_127_3477_n2724, DP_OP_425J2_127_3477_n2723,
         DP_OP_425J2_127_3477_n2722, DP_OP_425J2_127_3477_n2721,
         DP_OP_425J2_127_3477_n2720, DP_OP_425J2_127_3477_n2719,
         DP_OP_425J2_127_3477_n2718, DP_OP_425J2_127_3477_n2717,
         DP_OP_425J2_127_3477_n2716, DP_OP_425J2_127_3477_n2715,
         DP_OP_425J2_127_3477_n2714, DP_OP_425J2_127_3477_n2713,
         DP_OP_425J2_127_3477_n2712, DP_OP_425J2_127_3477_n2711,
         DP_OP_425J2_127_3477_n2710, DP_OP_425J2_127_3477_n2709,
         DP_OP_425J2_127_3477_n2708, DP_OP_425J2_127_3477_n2707,
         DP_OP_425J2_127_3477_n2706, DP_OP_425J2_127_3477_n2705,
         DP_OP_425J2_127_3477_n2704, DP_OP_425J2_127_3477_n2703,
         DP_OP_425J2_127_3477_n2702, DP_OP_425J2_127_3477_n2701,
         DP_OP_425J2_127_3477_n2700, DP_OP_425J2_127_3477_n2699,
         DP_OP_425J2_127_3477_n2696, DP_OP_425J2_127_3477_n2694,
         DP_OP_425J2_127_3477_n2692, DP_OP_425J2_127_3477_n2691,
         DP_OP_425J2_127_3477_n2690, DP_OP_425J2_127_3477_n2688,
         DP_OP_425J2_127_3477_n2686, DP_OP_425J2_127_3477_n2685,
         DP_OP_425J2_127_3477_n2684, DP_OP_425J2_127_3477_n2683,
         DP_OP_425J2_127_3477_n2682, DP_OP_425J2_127_3477_n2681,
         DP_OP_425J2_127_3477_n2680, DP_OP_425J2_127_3477_n2679,
         DP_OP_425J2_127_3477_n2678, DP_OP_425J2_127_3477_n2677,
         DP_OP_425J2_127_3477_n2676, DP_OP_425J2_127_3477_n2675,
         DP_OP_425J2_127_3477_n2674, DP_OP_425J2_127_3477_n2673,
         DP_OP_425J2_127_3477_n2672, DP_OP_425J2_127_3477_n2671,
         DP_OP_425J2_127_3477_n2670, DP_OP_425J2_127_3477_n2669,
         DP_OP_425J2_127_3477_n2668, DP_OP_425J2_127_3477_n2667,
         DP_OP_425J2_127_3477_n2666, DP_OP_425J2_127_3477_n2665,
         DP_OP_425J2_127_3477_n2664, DP_OP_425J2_127_3477_n2663,
         DP_OP_425J2_127_3477_n2662, DP_OP_425J2_127_3477_n2661,
         DP_OP_425J2_127_3477_n2660, DP_OP_425J2_127_3477_n2659,
         DP_OP_425J2_127_3477_n2658, DP_OP_425J2_127_3477_n2657,
         DP_OP_425J2_127_3477_n2656, DP_OP_425J2_127_3477_n2655,
         DP_OP_425J2_127_3477_n2654, DP_OP_425J2_127_3477_n2652,
         DP_OP_425J2_127_3477_n2650, DP_OP_425J2_127_3477_n2649,
         DP_OP_425J2_127_3477_n2646, DP_OP_425J2_127_3477_n2644,
         DP_OP_425J2_127_3477_n2643, DP_OP_425J2_127_3477_n2642,
         DP_OP_425J2_127_3477_n2641, DP_OP_425J2_127_3477_n2640,
         DP_OP_425J2_127_3477_n2639, DP_OP_425J2_127_3477_n2638,
         DP_OP_425J2_127_3477_n2637, DP_OP_425J2_127_3477_n2636,
         DP_OP_425J2_127_3477_n2635, DP_OP_425J2_127_3477_n2634,
         DP_OP_425J2_127_3477_n2633, DP_OP_425J2_127_3477_n2632,
         DP_OP_425J2_127_3477_n2631, DP_OP_425J2_127_3477_n2630,
         DP_OP_425J2_127_3477_n2629, DP_OP_425J2_127_3477_n2628,
         DP_OP_425J2_127_3477_n2627, DP_OP_425J2_127_3477_n2626,
         DP_OP_425J2_127_3477_n2625, DP_OP_425J2_127_3477_n2624,
         DP_OP_425J2_127_3477_n2623, DP_OP_425J2_127_3477_n2622,
         DP_OP_425J2_127_3477_n2621, DP_OP_425J2_127_3477_n2620,
         DP_OP_425J2_127_3477_n2619, DP_OP_425J2_127_3477_n2618,
         DP_OP_425J2_127_3477_n2617, DP_OP_425J2_127_3477_n2616,
         DP_OP_425J2_127_3477_n2615, DP_OP_425J2_127_3477_n2614,
         DP_OP_425J2_127_3477_n2613, DP_OP_425J2_127_3477_n2612,
         DP_OP_425J2_127_3477_n2611, DP_OP_425J2_127_3477_n2610,
         DP_OP_425J2_127_3477_n2598, DP_OP_425J2_127_3477_n2597,
         DP_OP_425J2_127_3477_n2596, DP_OP_425J2_127_3477_n2595,
         DP_OP_425J2_127_3477_n2594, DP_OP_425J2_127_3477_n2593,
         DP_OP_425J2_127_3477_n2592, DP_OP_425J2_127_3477_n2591,
         DP_OP_425J2_127_3477_n2590, DP_OP_425J2_127_3477_n2589,
         DP_OP_425J2_127_3477_n2588, DP_OP_425J2_127_3477_n2587,
         DP_OP_425J2_127_3477_n2586, DP_OP_425J2_127_3477_n2585,
         DP_OP_425J2_127_3477_n2584, DP_OP_425J2_127_3477_n2583,
         DP_OP_425J2_127_3477_n2582, DP_OP_425J2_127_3477_n2581,
         DP_OP_425J2_127_3477_n2580, DP_OP_425J2_127_3477_n2579,
         DP_OP_425J2_127_3477_n2578, DP_OP_425J2_127_3477_n2577,
         DP_OP_425J2_127_3477_n2576, DP_OP_425J2_127_3477_n2575,
         DP_OP_425J2_127_3477_n2574, DP_OP_425J2_127_3477_n2573,
         DP_OP_425J2_127_3477_n2572, DP_OP_425J2_127_3477_n2571,
         DP_OP_425J2_127_3477_n2570, DP_OP_425J2_127_3477_n2569,
         DP_OP_425J2_127_3477_n2568, DP_OP_425J2_127_3477_n2567,
         DP_OP_425J2_127_3477_n2566, DP_OP_425J2_127_3477_n2565,
         DP_OP_425J2_127_3477_n2564, DP_OP_425J2_127_3477_n2563,
         DP_OP_425J2_127_3477_n2559, DP_OP_425J2_127_3477_n2558,
         DP_OP_425J2_127_3477_n2557, DP_OP_425J2_127_3477_n2555,
         DP_OP_425J2_127_3477_n2554, DP_OP_425J2_127_3477_n2553,
         DP_OP_425J2_127_3477_n2552, DP_OP_425J2_127_3477_n2551,
         DP_OP_425J2_127_3477_n2550, DP_OP_425J2_127_3477_n2549,
         DP_OP_425J2_127_3477_n2548, DP_OP_425J2_127_3477_n2547,
         DP_OP_425J2_127_3477_n2546, DP_OP_425J2_127_3477_n2545,
         DP_OP_425J2_127_3477_n2544, DP_OP_425J2_127_3477_n2543,
         DP_OP_425J2_127_3477_n2542, DP_OP_425J2_127_3477_n2541,
         DP_OP_425J2_127_3477_n2540, DP_OP_425J2_127_3477_n2539,
         DP_OP_425J2_127_3477_n2538, DP_OP_425J2_127_3477_n2537,
         DP_OP_425J2_127_3477_n2536, DP_OP_425J2_127_3477_n2535,
         DP_OP_425J2_127_3477_n2534, DP_OP_425J2_127_3477_n2533,
         DP_OP_425J2_127_3477_n2532, DP_OP_425J2_127_3477_n2531,
         DP_OP_425J2_127_3477_n2530, DP_OP_425J2_127_3477_n2529,
         DP_OP_425J2_127_3477_n2528, DP_OP_425J2_127_3477_n2527,
         DP_OP_425J2_127_3477_n2526, DP_OP_425J2_127_3477_n2525,
         DP_OP_425J2_127_3477_n2524, DP_OP_425J2_127_3477_n2523,
         DP_OP_425J2_127_3477_n2519, DP_OP_425J2_127_3477_n2518,
         DP_OP_425J2_127_3477_n2511, DP_OP_425J2_127_3477_n2510,
         DP_OP_425J2_127_3477_n2509, DP_OP_425J2_127_3477_n2508,
         DP_OP_425J2_127_3477_n2507, DP_OP_425J2_127_3477_n2506,
         DP_OP_425J2_127_3477_n2505, DP_OP_425J2_127_3477_n2504,
         DP_OP_425J2_127_3477_n2503, DP_OP_425J2_127_3477_n2502,
         DP_OP_425J2_127_3477_n2501, DP_OP_425J2_127_3477_n2500,
         DP_OP_425J2_127_3477_n2499, DP_OP_425J2_127_3477_n2498,
         DP_OP_425J2_127_3477_n2497, DP_OP_425J2_127_3477_n2496,
         DP_OP_425J2_127_3477_n2495, DP_OP_425J2_127_3477_n2494,
         DP_OP_425J2_127_3477_n2493, DP_OP_425J2_127_3477_n2492,
         DP_OP_425J2_127_3477_n2491, DP_OP_425J2_127_3477_n2490,
         DP_OP_425J2_127_3477_n2489, DP_OP_425J2_127_3477_n2488,
         DP_OP_425J2_127_3477_n2487, DP_OP_425J2_127_3477_n2486,
         DP_OP_425J2_127_3477_n2485, DP_OP_425J2_127_3477_n2484,
         DP_OP_425J2_127_3477_n2483, DP_OP_425J2_127_3477_n2482,
         DP_OP_425J2_127_3477_n2481, DP_OP_425J2_127_3477_n2480,
         DP_OP_425J2_127_3477_n2479, DP_OP_425J2_127_3477_n2477,
         DP_OP_425J2_127_3477_n2476, DP_OP_425J2_127_3477_n2475,
         DP_OP_425J2_127_3477_n2472, DP_OP_425J2_127_3477_n2469,
         DP_OP_425J2_127_3477_n2466, DP_OP_425J2_127_3477_n2465,
         DP_OP_425J2_127_3477_n2464, DP_OP_425J2_127_3477_n2463,
         DP_OP_425J2_127_3477_n2462, DP_OP_425J2_127_3477_n2461,
         DP_OP_425J2_127_3477_n2460, DP_OP_425J2_127_3477_n2459,
         DP_OP_425J2_127_3477_n2458, DP_OP_425J2_127_3477_n2457,
         DP_OP_425J2_127_3477_n2456, DP_OP_425J2_127_3477_n2455,
         DP_OP_425J2_127_3477_n2454, DP_OP_425J2_127_3477_n2453,
         DP_OP_425J2_127_3477_n2452, DP_OP_425J2_127_3477_n2451,
         DP_OP_425J2_127_3477_n2450, DP_OP_425J2_127_3477_n2449,
         DP_OP_425J2_127_3477_n2448, DP_OP_425J2_127_3477_n2447,
         DP_OP_425J2_127_3477_n2446, DP_OP_425J2_127_3477_n2445,
         DP_OP_425J2_127_3477_n2444, DP_OP_425J2_127_3477_n2443,
         DP_OP_425J2_127_3477_n2442, DP_OP_425J2_127_3477_n2441,
         DP_OP_425J2_127_3477_n2440, DP_OP_425J2_127_3477_n2439,
         DP_OP_425J2_127_3477_n2438, DP_OP_425J2_127_3477_n2437,
         DP_OP_425J2_127_3477_n2436, DP_OP_425J2_127_3477_n2435,
         DP_OP_425J2_127_3477_n2434, DP_OP_425J2_127_3477_n2433,
         DP_OP_425J2_127_3477_n2431, DP_OP_425J2_127_3477_n2430,
         DP_OP_425J2_127_3477_n2429, DP_OP_425J2_127_3477_n2428,
         DP_OP_425J2_127_3477_n2427, DP_OP_425J2_127_3477_n2424,
         DP_OP_425J2_127_3477_n2423, DP_OP_425J2_127_3477_n2422,
         DP_OP_425J2_127_3477_n2421, DP_OP_425J2_127_3477_n2420,
         DP_OP_425J2_127_3477_n2419, DP_OP_425J2_127_3477_n2418,
         DP_OP_425J2_127_3477_n2417, DP_OP_425J2_127_3477_n2416,
         DP_OP_425J2_127_3477_n2415, DP_OP_425J2_127_3477_n2414,
         DP_OP_425J2_127_3477_n2413, DP_OP_425J2_127_3477_n2412,
         DP_OP_425J2_127_3477_n2411, DP_OP_425J2_127_3477_n2410,
         DP_OP_425J2_127_3477_n2409, DP_OP_425J2_127_3477_n2408,
         DP_OP_425J2_127_3477_n2407, DP_OP_425J2_127_3477_n2406,
         DP_OP_425J2_127_3477_n2405, DP_OP_425J2_127_3477_n2404,
         DP_OP_425J2_127_3477_n2403, DP_OP_425J2_127_3477_n2402,
         DP_OP_425J2_127_3477_n2401, DP_OP_425J2_127_3477_n2400,
         DP_OP_425J2_127_3477_n2399, DP_OP_425J2_127_3477_n2398,
         DP_OP_425J2_127_3477_n2397, DP_OP_425J2_127_3477_n2396,
         DP_OP_425J2_127_3477_n2395, DP_OP_425J2_127_3477_n2394,
         DP_OP_425J2_127_3477_n2393, DP_OP_425J2_127_3477_n2392,
         DP_OP_425J2_127_3477_n2391, DP_OP_425J2_127_3477_n2387,
         DP_OP_425J2_127_3477_n2386, DP_OP_425J2_127_3477_n2384,
         DP_OP_425J2_127_3477_n2383, DP_OP_425J2_127_3477_n2382,
         DP_OP_425J2_127_3477_n2381, DP_OP_425J2_127_3477_n2378,
         DP_OP_425J2_127_3477_n2377, DP_OP_425J2_127_3477_n2376,
         DP_OP_425J2_127_3477_n2375, DP_OP_425J2_127_3477_n2374,
         DP_OP_425J2_127_3477_n2373, DP_OP_425J2_127_3477_n2372,
         DP_OP_425J2_127_3477_n2371, DP_OP_425J2_127_3477_n2370,
         DP_OP_425J2_127_3477_n2369, DP_OP_425J2_127_3477_n2368,
         DP_OP_425J2_127_3477_n2367, DP_OP_425J2_127_3477_n2366,
         DP_OP_425J2_127_3477_n2365, DP_OP_425J2_127_3477_n2364,
         DP_OP_425J2_127_3477_n2363, DP_OP_425J2_127_3477_n2362,
         DP_OP_425J2_127_3477_n2361, DP_OP_425J2_127_3477_n2360,
         DP_OP_425J2_127_3477_n2359, DP_OP_425J2_127_3477_n2358,
         DP_OP_425J2_127_3477_n2357, DP_OP_425J2_127_3477_n2356,
         DP_OP_425J2_127_3477_n2355, DP_OP_425J2_127_3477_n2354,
         DP_OP_425J2_127_3477_n2353, DP_OP_425J2_127_3477_n2352,
         DP_OP_425J2_127_3477_n2351, DP_OP_425J2_127_3477_n2350,
         DP_OP_425J2_127_3477_n2349, DP_OP_425J2_127_3477_n2348,
         DP_OP_425J2_127_3477_n2347, DP_OP_425J2_127_3477_n2346,
         DP_OP_425J2_127_3477_n2342, DP_OP_425J2_127_3477_n2341,
         DP_OP_425J2_127_3477_n2340, DP_OP_425J2_127_3477_n2339,
         DP_OP_425J2_127_3477_n2337, DP_OP_425J2_127_3477_n2336,
         DP_OP_425J2_127_3477_n2335, DP_OP_425J2_127_3477_n2334,
         DP_OP_425J2_127_3477_n2333, DP_OP_425J2_127_3477_n2332,
         DP_OP_425J2_127_3477_n2331, DP_OP_425J2_127_3477_n2330,
         DP_OP_425J2_127_3477_n2329, DP_OP_425J2_127_3477_n2328,
         DP_OP_425J2_127_3477_n2327, DP_OP_425J2_127_3477_n2326,
         DP_OP_425J2_127_3477_n2325, DP_OP_425J2_127_3477_n2324,
         DP_OP_425J2_127_3477_n2323, DP_OP_425J2_127_3477_n2322,
         DP_OP_425J2_127_3477_n2321, DP_OP_425J2_127_3477_n2320,
         DP_OP_425J2_127_3477_n2319, DP_OP_425J2_127_3477_n2318,
         DP_OP_425J2_127_3477_n2317, DP_OP_425J2_127_3477_n2316,
         DP_OP_425J2_127_3477_n2315, DP_OP_425J2_127_3477_n2314,
         DP_OP_425J2_127_3477_n2313, DP_OP_425J2_127_3477_n2312,
         DP_OP_425J2_127_3477_n2311, DP_OP_425J2_127_3477_n2310,
         DP_OP_425J2_127_3477_n2309, DP_OP_425J2_127_3477_n2308,
         DP_OP_425J2_127_3477_n2307, DP_OP_425J2_127_3477_n2306,
         DP_OP_425J2_127_3477_n2305, DP_OP_425J2_127_3477_n2304,
         DP_OP_425J2_127_3477_n2302, DP_OP_425J2_127_3477_n2300,
         DP_OP_425J2_127_3477_n2297, DP_OP_425J2_127_3477_n2296,
         DP_OP_425J2_127_3477_n2294, DP_OP_425J2_127_3477_n2293,
         DP_OP_425J2_127_3477_n2292, DP_OP_425J2_127_3477_n2291,
         DP_OP_425J2_127_3477_n2290, DP_OP_425J2_127_3477_n2289,
         DP_OP_425J2_127_3477_n2288, DP_OP_425J2_127_3477_n2287,
         DP_OP_425J2_127_3477_n2286, DP_OP_425J2_127_3477_n2285,
         DP_OP_425J2_127_3477_n2284, DP_OP_425J2_127_3477_n2283,
         DP_OP_425J2_127_3477_n2282, DP_OP_425J2_127_3477_n2281,
         DP_OP_425J2_127_3477_n2280, DP_OP_425J2_127_3477_n2279,
         DP_OP_425J2_127_3477_n2278, DP_OP_425J2_127_3477_n2277,
         DP_OP_425J2_127_3477_n2276, DP_OP_425J2_127_3477_n2275,
         DP_OP_425J2_127_3477_n2274, DP_OP_425J2_127_3477_n2273,
         DP_OP_425J2_127_3477_n2272, DP_OP_425J2_127_3477_n2271,
         DP_OP_425J2_127_3477_n2270, DP_OP_425J2_127_3477_n2269,
         DP_OP_425J2_127_3477_n2268, DP_OP_425J2_127_3477_n2267,
         DP_OP_425J2_127_3477_n2266, DP_OP_425J2_127_3477_n2265,
         DP_OP_425J2_127_3477_n2264, DP_OP_425J2_127_3477_n2263,
         DP_OP_425J2_127_3477_n2262, DP_OP_425J2_127_3477_n2261,
         DP_OP_425J2_127_3477_n2260, DP_OP_425J2_127_3477_n2259,
         DP_OP_425J2_127_3477_n2255, DP_OP_425J2_127_3477_n2252,
         DP_OP_425J2_127_3477_n2250, DP_OP_425J2_127_3477_n2249,
         DP_OP_425J2_127_3477_n2248, DP_OP_425J2_127_3477_n2247,
         DP_OP_425J2_127_3477_n2246, DP_OP_425J2_127_3477_n2245,
         DP_OP_425J2_127_3477_n2244, DP_OP_425J2_127_3477_n2243,
         DP_OP_425J2_127_3477_n2242, DP_OP_425J2_127_3477_n2241,
         DP_OP_425J2_127_3477_n2240, DP_OP_425J2_127_3477_n2239,
         DP_OP_425J2_127_3477_n2238, DP_OP_425J2_127_3477_n2237,
         DP_OP_425J2_127_3477_n2236, DP_OP_425J2_127_3477_n2235,
         DP_OP_425J2_127_3477_n2234, DP_OP_425J2_127_3477_n2233,
         DP_OP_425J2_127_3477_n2232, DP_OP_425J2_127_3477_n2231,
         DP_OP_425J2_127_3477_n2230, DP_OP_425J2_127_3477_n2229,
         DP_OP_425J2_127_3477_n2228, DP_OP_425J2_127_3477_n2227,
         DP_OP_425J2_127_3477_n2226, DP_OP_425J2_127_3477_n2225,
         DP_OP_425J2_127_3477_n2224, DP_OP_425J2_127_3477_n2223,
         DP_OP_425J2_127_3477_n2222, DP_OP_425J2_127_3477_n2221,
         DP_OP_425J2_127_3477_n2220, DP_OP_425J2_127_3477_n2219,
         DP_OP_425J2_127_3477_n2218, DP_OP_425J2_127_3477_n2217,
         DP_OP_425J2_127_3477_n2215, DP_OP_425J2_127_3477_n2214,
         DP_OP_425J2_127_3477_n2213, DP_OP_425J2_127_3477_n2209,
         DP_OP_425J2_127_3477_n2205, DP_OP_425J2_127_3477_n2204,
         DP_OP_425J2_127_3477_n2203, DP_OP_425J2_127_3477_n2202,
         DP_OP_425J2_127_3477_n2201, DP_OP_425J2_127_3477_n2200,
         DP_OP_425J2_127_3477_n2199, DP_OP_425J2_127_3477_n2198,
         DP_OP_425J2_127_3477_n2197, DP_OP_425J2_127_3477_n2196,
         DP_OP_425J2_127_3477_n2195, DP_OP_425J2_127_3477_n2194,
         DP_OP_425J2_127_3477_n2193, DP_OP_425J2_127_3477_n2192,
         DP_OP_425J2_127_3477_n2191, DP_OP_425J2_127_3477_n2190,
         DP_OP_425J2_127_3477_n2189, DP_OP_425J2_127_3477_n2188,
         DP_OP_425J2_127_3477_n2187, DP_OP_425J2_127_3477_n2186,
         DP_OP_425J2_127_3477_n2185, DP_OP_425J2_127_3477_n2184,
         DP_OP_425J2_127_3477_n2183, DP_OP_425J2_127_3477_n2182,
         DP_OP_425J2_127_3477_n2181, DP_OP_425J2_127_3477_n2180,
         DP_OP_425J2_127_3477_n2179, DP_OP_425J2_127_3477_n2178,
         DP_OP_425J2_127_3477_n2177, DP_OP_425J2_127_3477_n2176,
         DP_OP_425J2_127_3477_n2175, DP_OP_425J2_127_3477_n2174,
         DP_OP_425J2_127_3477_n2173, DP_OP_425J2_127_3477_n2172,
         DP_OP_425J2_127_3477_n2169, DP_OP_425J2_127_3477_n2168,
         DP_OP_425J2_127_3477_n2166, DP_OP_425J2_127_3477_n2164,
         DP_OP_425J2_127_3477_n2163, DP_OP_425J2_127_3477_n2162,
         DP_OP_425J2_127_3477_n2161, DP_OP_425J2_127_3477_n2160,
         DP_OP_425J2_127_3477_n2159, DP_OP_425J2_127_3477_n2158,
         DP_OP_425J2_127_3477_n2157, DP_OP_425J2_127_3477_n2156,
         DP_OP_425J2_127_3477_n2155, DP_OP_425J2_127_3477_n2154,
         DP_OP_425J2_127_3477_n2153, DP_OP_425J2_127_3477_n2152,
         DP_OP_425J2_127_3477_n2151, DP_OP_425J2_127_3477_n2150,
         DP_OP_425J2_127_3477_n2149, DP_OP_425J2_127_3477_n2148,
         DP_OP_425J2_127_3477_n2147, DP_OP_425J2_127_3477_n2146,
         DP_OP_425J2_127_3477_n2145, DP_OP_425J2_127_3477_n2144,
         DP_OP_425J2_127_3477_n2143, DP_OP_425J2_127_3477_n2142,
         DP_OP_425J2_127_3477_n2141, DP_OP_425J2_127_3477_n2140,
         DP_OP_425J2_127_3477_n2139, DP_OP_425J2_127_3477_n2138,
         DP_OP_425J2_127_3477_n2137, DP_OP_425J2_127_3477_n2136,
         DP_OP_425J2_127_3477_n2135, DP_OP_425J2_127_3477_n2134,
         DP_OP_425J2_127_3477_n2133, DP_OP_425J2_127_3477_n2132,
         DP_OP_425J2_127_3477_n2131, DP_OP_425J2_127_3477_n2130,
         DP_OP_425J2_127_3477_n2129, DP_OP_425J2_127_3477_n2128,
         DP_OP_425J2_127_3477_n2127, DP_OP_425J2_127_3477_n2126,
         DP_OP_425J2_127_3477_n2122, DP_OP_425J2_127_3477_n2120,
         DP_OP_425J2_127_3477_n2119, DP_OP_425J2_127_3477_n2118,
         DP_OP_425J2_127_3477_n2117, DP_OP_425J2_127_3477_n2116,
         DP_OP_425J2_127_3477_n2115, DP_OP_425J2_127_3477_n2114,
         DP_OP_425J2_127_3477_n2113, DP_OP_425J2_127_3477_n2112,
         DP_OP_425J2_127_3477_n2111, DP_OP_425J2_127_3477_n2110,
         DP_OP_425J2_127_3477_n2109, DP_OP_425J2_127_3477_n2108,
         DP_OP_425J2_127_3477_n2107, DP_OP_425J2_127_3477_n2106,
         DP_OP_425J2_127_3477_n2105, DP_OP_425J2_127_3477_n2104,
         DP_OP_425J2_127_3477_n2103, DP_OP_425J2_127_3477_n2102,
         DP_OP_425J2_127_3477_n2101, DP_OP_425J2_127_3477_n2100,
         DP_OP_425J2_127_3477_n2099, DP_OP_425J2_127_3477_n2098,
         DP_OP_425J2_127_3477_n2097, DP_OP_425J2_127_3477_n2096,
         DP_OP_425J2_127_3477_n2095, DP_OP_425J2_127_3477_n2094,
         DP_OP_425J2_127_3477_n2093, DP_OP_425J2_127_3477_n2092,
         DP_OP_425J2_127_3477_n2091, DP_OP_425J2_127_3477_n2090,
         DP_OP_425J2_127_3477_n2089, DP_OP_425J2_127_3477_n2088,
         DP_OP_425J2_127_3477_n2087, DP_OP_425J2_127_3477_n2086,
         DP_OP_425J2_127_3477_n2084, DP_OP_425J2_127_3477_n2083,
         DP_OP_425J2_127_3477_n2079, DP_OP_425J2_127_3477_n2078,
         DP_OP_425J2_127_3477_n2077, DP_OP_425J2_127_3477_n2075,
         DP_OP_425J2_127_3477_n2074, DP_OP_425J2_127_3477_n2073,
         DP_OP_425J2_127_3477_n2072, DP_OP_425J2_127_3477_n2071,
         DP_OP_425J2_127_3477_n2070, DP_OP_425J2_127_3477_n2069,
         DP_OP_425J2_127_3477_n2068, DP_OP_425J2_127_3477_n2067,
         DP_OP_425J2_127_3477_n2066, DP_OP_425J2_127_3477_n2065,
         DP_OP_425J2_127_3477_n2064, DP_OP_425J2_127_3477_n2063,
         DP_OP_425J2_127_3477_n2062, DP_OP_425J2_127_3477_n2061,
         DP_OP_425J2_127_3477_n2060, DP_OP_425J2_127_3477_n2059,
         DP_OP_425J2_127_3477_n2058, DP_OP_425J2_127_3477_n2057,
         DP_OP_425J2_127_3477_n2056, DP_OP_425J2_127_3477_n2055,
         DP_OP_425J2_127_3477_n2054, DP_OP_425J2_127_3477_n2053,
         DP_OP_425J2_127_3477_n2052, DP_OP_425J2_127_3477_n2051,
         DP_OP_425J2_127_3477_n2050, DP_OP_425J2_127_3477_n2049,
         DP_OP_425J2_127_3477_n2048, DP_OP_425J2_127_3477_n2047,
         DP_OP_425J2_127_3477_n2046, DP_OP_425J2_127_3477_n2045,
         DP_OP_425J2_127_3477_n2044, DP_OP_425J2_127_3477_n2043,
         DP_OP_425J2_127_3477_n2042, DP_OP_425J2_127_3477_n2041,
         DP_OP_425J2_127_3477_n2040, DP_OP_425J2_127_3477_n2039,
         DP_OP_425J2_127_3477_n2033, DP_OP_425J2_127_3477_n2029,
         DP_OP_425J2_127_3477_n2028, DP_OP_425J2_127_3477_n2027,
         DP_OP_425J2_127_3477_n2026, DP_OP_425J2_127_3477_n2025,
         DP_OP_425J2_127_3477_n2024, DP_OP_425J2_127_3477_n2023,
         DP_OP_425J2_127_3477_n2022, DP_OP_425J2_127_3477_n2021,
         DP_OP_425J2_127_3477_n2020, DP_OP_425J2_127_3477_n2019,
         DP_OP_425J2_127_3477_n2018, DP_OP_425J2_127_3477_n2017,
         DP_OP_425J2_127_3477_n2016, DP_OP_425J2_127_3477_n2015,
         DP_OP_425J2_127_3477_n2014, DP_OP_425J2_127_3477_n2013,
         DP_OP_425J2_127_3477_n2012, DP_OP_425J2_127_3477_n2011,
         DP_OP_425J2_127_3477_n2010, DP_OP_425J2_127_3477_n2009,
         DP_OP_425J2_127_3477_n2008, DP_OP_425J2_127_3477_n2007,
         DP_OP_425J2_127_3477_n2006, DP_OP_425J2_127_3477_n2005,
         DP_OP_425J2_127_3477_n2004, DP_OP_425J2_127_3477_n2003,
         DP_OP_425J2_127_3477_n2002, DP_OP_425J2_127_3477_n2001,
         DP_OP_425J2_127_3477_n2000, DP_OP_425J2_127_3477_n1999,
         DP_OP_425J2_127_3477_n1998, DP_OP_425J2_127_3477_n1997,
         DP_OP_425J2_127_3477_n1995, DP_OP_425J2_127_3477_n1992,
         DP_OP_425J2_127_3477_n1991, DP_OP_425J2_127_3477_n1990,
         DP_OP_425J2_127_3477_n1989, DP_OP_425J2_127_3477_n1985,
         DP_OP_425J2_127_3477_n1984, DP_OP_425J2_127_3477_n1983,
         DP_OP_425J2_127_3477_n1982, DP_OP_425J2_127_3477_n1981,
         DP_OP_425J2_127_3477_n1980, DP_OP_425J2_127_3477_n1979,
         DP_OP_425J2_127_3477_n1978, DP_OP_425J2_127_3477_n1977,
         DP_OP_425J2_127_3477_n1976, DP_OP_425J2_127_3477_n1975,
         DP_OP_425J2_127_3477_n1974, DP_OP_425J2_127_3477_n1973,
         DP_OP_425J2_127_3477_n1972, DP_OP_425J2_127_3477_n1971,
         DP_OP_425J2_127_3477_n1970, DP_OP_425J2_127_3477_n1969,
         DP_OP_425J2_127_3477_n1968, DP_OP_425J2_127_3477_n1967,
         DP_OP_425J2_127_3477_n1966, DP_OP_425J2_127_3477_n1965,
         DP_OP_425J2_127_3477_n1964, DP_OP_425J2_127_3477_n1963,
         DP_OP_425J2_127_3477_n1962, DP_OP_425J2_127_3477_n1961,
         DP_OP_425J2_127_3477_n1960, DP_OP_425J2_127_3477_n1959,
         DP_OP_425J2_127_3477_n1958, DP_OP_425J2_127_3477_n1957,
         DP_OP_425J2_127_3477_n1956, DP_OP_425J2_127_3477_n1955,
         DP_OP_425J2_127_3477_n1954, DP_OP_425J2_127_3477_n1953,
         DP_OP_425J2_127_3477_n1951, DP_OP_425J2_127_3477_n1950,
         DP_OP_425J2_127_3477_n1945, DP_OP_425J2_127_3477_n1941,
         DP_OP_425J2_127_3477_n1940, DP_OP_425J2_127_3477_n1939,
         DP_OP_425J2_127_3477_n1938, DP_OP_425J2_127_3477_n1937,
         DP_OP_425J2_127_3477_n1936, DP_OP_425J2_127_3477_n1935,
         DP_OP_425J2_127_3477_n1934, DP_OP_425J2_127_3477_n1933,
         DP_OP_425J2_127_3477_n1932, DP_OP_425J2_127_3477_n1931,
         DP_OP_425J2_127_3477_n1930, DP_OP_425J2_127_3477_n1929,
         DP_OP_425J2_127_3477_n1928, DP_OP_425J2_127_3477_n1927,
         DP_OP_425J2_127_3477_n1926, DP_OP_425J2_127_3477_n1925,
         DP_OP_425J2_127_3477_n1924, DP_OP_425J2_127_3477_n1923,
         DP_OP_425J2_127_3477_n1922, DP_OP_425J2_127_3477_n1921,
         DP_OP_425J2_127_3477_n1920, DP_OP_425J2_127_3477_n1919,
         DP_OP_425J2_127_3477_n1918, DP_OP_425J2_127_3477_n1917,
         DP_OP_425J2_127_3477_n1916, DP_OP_425J2_127_3477_n1915,
         DP_OP_425J2_127_3477_n1914, DP_OP_425J2_127_3477_n1913,
         DP_OP_425J2_127_3477_n1912, DP_OP_425J2_127_3477_n1911,
         DP_OP_425J2_127_3477_n1910, DP_OP_425J2_127_3477_n1907,
         DP_OP_425J2_127_3477_n1905, DP_OP_425J2_127_3477_n1903,
         DP_OP_425J2_127_3477_n1901, DP_OP_425J2_127_3477_n1897,
         DP_OP_425J2_127_3477_n1896, DP_OP_425J2_127_3477_n1895,
         DP_OP_425J2_127_3477_n1894, DP_OP_425J2_127_3477_n1893,
         DP_OP_425J2_127_3477_n1892, DP_OP_425J2_127_3477_n1891,
         DP_OP_425J2_127_3477_n1890, DP_OP_425J2_127_3477_n1889,
         DP_OP_425J2_127_3477_n1888, DP_OP_425J2_127_3477_n1887,
         DP_OP_425J2_127_3477_n1886, DP_OP_425J2_127_3477_n1885,
         DP_OP_425J2_127_3477_n1884, DP_OP_425J2_127_3477_n1883,
         DP_OP_425J2_127_3477_n1882, DP_OP_425J2_127_3477_n1881,
         DP_OP_425J2_127_3477_n1880, DP_OP_425J2_127_3477_n1879,
         DP_OP_425J2_127_3477_n1878, DP_OP_425J2_127_3477_n1877,
         DP_OP_425J2_127_3477_n1876, DP_OP_425J2_127_3477_n1875,
         DP_OP_425J2_127_3477_n1874, DP_OP_425J2_127_3477_n1873,
         DP_OP_425J2_127_3477_n1872, DP_OP_425J2_127_3477_n1871,
         DP_OP_425J2_127_3477_n1870, DP_OP_425J2_127_3477_n1869,
         DP_OP_425J2_127_3477_n1868, DP_OP_425J2_127_3477_n1867,
         DP_OP_425J2_127_3477_n1866, DP_OP_425J2_127_3477_n1864,
         DP_OP_425J2_127_3477_n1863, DP_OP_425J2_127_3477_n1862,
         DP_OP_425J2_127_3477_n1861, DP_OP_425J2_127_3477_n1860,
         DP_OP_425J2_127_3477_n1858, DP_OP_425J2_127_3477_n1855,
         DP_OP_425J2_127_3477_n1854, DP_OP_425J2_127_3477_n1853,
         DP_OP_425J2_127_3477_n1852, DP_OP_425J2_127_3477_n1851,
         DP_OP_425J2_127_3477_n1850, DP_OP_425J2_127_3477_n1849,
         DP_OP_425J2_127_3477_n1848, DP_OP_425J2_127_3477_n1847,
         DP_OP_425J2_127_3477_n1846, DP_OP_425J2_127_3477_n1845,
         DP_OP_425J2_127_3477_n1844, DP_OP_425J2_127_3477_n1843,
         DP_OP_425J2_127_3477_n1842, DP_OP_425J2_127_3477_n1841,
         DP_OP_425J2_127_3477_n1840, DP_OP_425J2_127_3477_n1839,
         DP_OP_425J2_127_3477_n1838, DP_OP_425J2_127_3477_n1837,
         DP_OP_425J2_127_3477_n1836, DP_OP_425J2_127_3477_n1835,
         DP_OP_425J2_127_3477_n1834, DP_OP_425J2_127_3477_n1833,
         DP_OP_425J2_127_3477_n1832, DP_OP_425J2_127_3477_n1831,
         DP_OP_425J2_127_3477_n1830, DP_OP_425J2_127_3477_n1829,
         DP_OP_425J2_127_3477_n1828, DP_OP_425J2_127_3477_n1827,
         DP_OP_425J2_127_3477_n1826, DP_OP_425J2_127_3477_n1825,
         DP_OP_425J2_127_3477_n1824, DP_OP_425J2_127_3477_n1823,
         DP_OP_425J2_127_3477_n1822, DP_OP_425J2_127_3477_n1788,
         DP_OP_425J2_127_3477_n1787, DP_OP_425J2_127_3477_n1786,
         DP_OP_425J2_127_3477_n1785, DP_OP_425J2_127_3477_n1784,
         DP_OP_425J2_127_3477_n1783, DP_OP_425J2_127_3477_n1782,
         DP_OP_425J2_127_3477_n1781, DP_OP_425J2_127_3477_n1780,
         DP_OP_425J2_127_3477_n1779, DP_OP_425J2_127_3477_n1778,
         DP_OP_425J2_127_3477_n1777, DP_OP_425J2_127_3477_n1776,
         DP_OP_425J2_127_3477_n1775, DP_OP_425J2_127_3477_n1774,
         DP_OP_425J2_127_3477_n1773, DP_OP_425J2_127_3477_n1772,
         DP_OP_425J2_127_3477_n1771, DP_OP_425J2_127_3477_n1770,
         DP_OP_425J2_127_3477_n1769, DP_OP_425J2_127_3477_n1768,
         DP_OP_425J2_127_3477_n1767, DP_OP_425J2_127_3477_n1766,
         DP_OP_425J2_127_3477_n1765, DP_OP_425J2_127_3477_n1764,
         DP_OP_425J2_127_3477_n1763, DP_OP_425J2_127_3477_n1762,
         DP_OP_425J2_127_3477_n1761, DP_OP_425J2_127_3477_n1760,
         DP_OP_425J2_127_3477_n1759, DP_OP_425J2_127_3477_n1758,
         DP_OP_425J2_127_3477_n1757, DP_OP_425J2_127_3477_n1756,
         DP_OP_425J2_127_3477_n1755, DP_OP_425J2_127_3477_n1754,
         DP_OP_425J2_127_3477_n1753, DP_OP_425J2_127_3477_n1752,
         DP_OP_425J2_127_3477_n1751, DP_OP_425J2_127_3477_n1750,
         DP_OP_425J2_127_3477_n1749, DP_OP_425J2_127_3477_n1748,
         DP_OP_425J2_127_3477_n1747, DP_OP_425J2_127_3477_n1746,
         DP_OP_425J2_127_3477_n1745, DP_OP_425J2_127_3477_n1744,
         DP_OP_425J2_127_3477_n1743, DP_OP_425J2_127_3477_n1742,
         DP_OP_425J2_127_3477_n1741, DP_OP_425J2_127_3477_n1740,
         DP_OP_425J2_127_3477_n1739, DP_OP_425J2_127_3477_n1738,
         DP_OP_425J2_127_3477_n1737, DP_OP_425J2_127_3477_n1736,
         DP_OP_425J2_127_3477_n1735, DP_OP_425J2_127_3477_n1734,
         DP_OP_425J2_127_3477_n1733, DP_OP_425J2_127_3477_n1732,
         DP_OP_425J2_127_3477_n1731, DP_OP_425J2_127_3477_n1730,
         DP_OP_425J2_127_3477_n1729, DP_OP_425J2_127_3477_n1728,
         DP_OP_425J2_127_3477_n1727, DP_OP_425J2_127_3477_n1726,
         DP_OP_425J2_127_3477_n1725, DP_OP_425J2_127_3477_n1724,
         DP_OP_425J2_127_3477_n1723, DP_OP_425J2_127_3477_n1722,
         DP_OP_425J2_127_3477_n1721, DP_OP_425J2_127_3477_n1720,
         DP_OP_425J2_127_3477_n1719, DP_OP_425J2_127_3477_n1718,
         DP_OP_425J2_127_3477_n1717, DP_OP_425J2_127_3477_n1716,
         DP_OP_425J2_127_3477_n1715, DP_OP_425J2_127_3477_n1714,
         DP_OP_425J2_127_3477_n1713, DP_OP_425J2_127_3477_n1712,
         DP_OP_425J2_127_3477_n1711, DP_OP_425J2_127_3477_n1710,
         DP_OP_425J2_127_3477_n1709, DP_OP_425J2_127_3477_n1708,
         DP_OP_425J2_127_3477_n1707, DP_OP_425J2_127_3477_n1706,
         DP_OP_425J2_127_3477_n1705, DP_OP_425J2_127_3477_n1704,
         DP_OP_425J2_127_3477_n1703, DP_OP_425J2_127_3477_n1702,
         DP_OP_425J2_127_3477_n1701, DP_OP_425J2_127_3477_n1700,
         DP_OP_425J2_127_3477_n1699, DP_OP_425J2_127_3477_n1698,
         DP_OP_425J2_127_3477_n1697, DP_OP_425J2_127_3477_n1696,
         DP_OP_425J2_127_3477_n1695, DP_OP_425J2_127_3477_n1694,
         DP_OP_425J2_127_3477_n1693, DP_OP_425J2_127_3477_n1692,
         DP_OP_425J2_127_3477_n1691, DP_OP_425J2_127_3477_n1690,
         DP_OP_425J2_127_3477_n1689, DP_OP_425J2_127_3477_n1688,
         DP_OP_425J2_127_3477_n1687, DP_OP_425J2_127_3477_n1686,
         DP_OP_425J2_127_3477_n1685, DP_OP_425J2_127_3477_n1684,
         DP_OP_425J2_127_3477_n1683, DP_OP_425J2_127_3477_n1682,
         DP_OP_425J2_127_3477_n1681, DP_OP_425J2_127_3477_n1680,
         DP_OP_425J2_127_3477_n1679, DP_OP_425J2_127_3477_n1678,
         DP_OP_425J2_127_3477_n1677, DP_OP_425J2_127_3477_n1676,
         DP_OP_425J2_127_3477_n1675, DP_OP_425J2_127_3477_n1674,
         DP_OP_425J2_127_3477_n1673, DP_OP_425J2_127_3477_n1672,
         DP_OP_425J2_127_3477_n1671, DP_OP_425J2_127_3477_n1670,
         DP_OP_425J2_127_3477_n1669, DP_OP_425J2_127_3477_n1668,
         DP_OP_425J2_127_3477_n1667, DP_OP_425J2_127_3477_n1666,
         DP_OP_425J2_127_3477_n1665, DP_OP_425J2_127_3477_n1664,
         DP_OP_425J2_127_3477_n1663, DP_OP_425J2_127_3477_n1662,
         DP_OP_425J2_127_3477_n1661, DP_OP_425J2_127_3477_n1660,
         DP_OP_425J2_127_3477_n1659, DP_OP_425J2_127_3477_n1658,
         DP_OP_425J2_127_3477_n1657, DP_OP_425J2_127_3477_n1656,
         DP_OP_425J2_127_3477_n1655, DP_OP_425J2_127_3477_n1654,
         DP_OP_425J2_127_3477_n1653, DP_OP_425J2_127_3477_n1652,
         DP_OP_425J2_127_3477_n1651, DP_OP_425J2_127_3477_n1650,
         DP_OP_425J2_127_3477_n1649, DP_OP_425J2_127_3477_n1648,
         DP_OP_425J2_127_3477_n1647, DP_OP_425J2_127_3477_n1646,
         DP_OP_425J2_127_3477_n1645, DP_OP_425J2_127_3477_n1644,
         DP_OP_425J2_127_3477_n1643, DP_OP_425J2_127_3477_n1642,
         DP_OP_425J2_127_3477_n1641, DP_OP_425J2_127_3477_n1640,
         DP_OP_425J2_127_3477_n1639, DP_OP_425J2_127_3477_n1638,
         DP_OP_425J2_127_3477_n1637, DP_OP_425J2_127_3477_n1636,
         DP_OP_425J2_127_3477_n1635, DP_OP_425J2_127_3477_n1634,
         DP_OP_425J2_127_3477_n1633, DP_OP_425J2_127_3477_n1632,
         DP_OP_425J2_127_3477_n1631, DP_OP_425J2_127_3477_n1630,
         DP_OP_425J2_127_3477_n1629, DP_OP_425J2_127_3477_n1628,
         DP_OP_425J2_127_3477_n1627, DP_OP_425J2_127_3477_n1626,
         DP_OP_425J2_127_3477_n1625, DP_OP_425J2_127_3477_n1624,
         DP_OP_425J2_127_3477_n1623, DP_OP_425J2_127_3477_n1622,
         DP_OP_425J2_127_3477_n1621, DP_OP_425J2_127_3477_n1620,
         DP_OP_425J2_127_3477_n1619, DP_OP_425J2_127_3477_n1618,
         DP_OP_425J2_127_3477_n1617, DP_OP_425J2_127_3477_n1616,
         DP_OP_425J2_127_3477_n1615, DP_OP_425J2_127_3477_n1614,
         DP_OP_425J2_127_3477_n1613, DP_OP_425J2_127_3477_n1612,
         DP_OP_425J2_127_3477_n1611, DP_OP_425J2_127_3477_n1610,
         DP_OP_425J2_127_3477_n1609, DP_OP_425J2_127_3477_n1608,
         DP_OP_425J2_127_3477_n1607, DP_OP_425J2_127_3477_n1606,
         DP_OP_425J2_127_3477_n1605, DP_OP_425J2_127_3477_n1604,
         DP_OP_425J2_127_3477_n1603, DP_OP_425J2_127_3477_n1602,
         DP_OP_425J2_127_3477_n1601, DP_OP_425J2_127_3477_n1600,
         DP_OP_425J2_127_3477_n1599, DP_OP_425J2_127_3477_n1598,
         DP_OP_425J2_127_3477_n1597, DP_OP_425J2_127_3477_n1596,
         DP_OP_425J2_127_3477_n1595, DP_OP_425J2_127_3477_n1594,
         DP_OP_425J2_127_3477_n1593, DP_OP_425J2_127_3477_n1592,
         DP_OP_425J2_127_3477_n1591, DP_OP_425J2_127_3477_n1590,
         DP_OP_425J2_127_3477_n1589, DP_OP_425J2_127_3477_n1588,
         DP_OP_425J2_127_3477_n1587, DP_OP_425J2_127_3477_n1586,
         DP_OP_425J2_127_3477_n1585, DP_OP_425J2_127_3477_n1584,
         DP_OP_425J2_127_3477_n1583, DP_OP_425J2_127_3477_n1582,
         DP_OP_425J2_127_3477_n1581, DP_OP_425J2_127_3477_n1580,
         DP_OP_425J2_127_3477_n1579, DP_OP_425J2_127_3477_n1578,
         DP_OP_425J2_127_3477_n1577, DP_OP_425J2_127_3477_n1576,
         DP_OP_425J2_127_3477_n1575, DP_OP_425J2_127_3477_n1574,
         DP_OP_425J2_127_3477_n1573, DP_OP_425J2_127_3477_n1572,
         DP_OP_425J2_127_3477_n1571, DP_OP_425J2_127_3477_n1570,
         DP_OP_425J2_127_3477_n1569, DP_OP_425J2_127_3477_n1568,
         DP_OP_425J2_127_3477_n1567, DP_OP_425J2_127_3477_n1566,
         DP_OP_425J2_127_3477_n1565, DP_OP_425J2_127_3477_n1564,
         DP_OP_425J2_127_3477_n1563, DP_OP_425J2_127_3477_n1562,
         DP_OP_425J2_127_3477_n1561, DP_OP_425J2_127_3477_n1560,
         DP_OP_425J2_127_3477_n1559, DP_OP_425J2_127_3477_n1558,
         DP_OP_425J2_127_3477_n1557, DP_OP_425J2_127_3477_n1556,
         DP_OP_425J2_127_3477_n1555, DP_OP_425J2_127_3477_n1554,
         DP_OP_425J2_127_3477_n1553, DP_OP_425J2_127_3477_n1552,
         DP_OP_425J2_127_3477_n1551, DP_OP_425J2_127_3477_n1550,
         DP_OP_425J2_127_3477_n1549, DP_OP_425J2_127_3477_n1548,
         DP_OP_425J2_127_3477_n1547, DP_OP_425J2_127_3477_n1546,
         DP_OP_425J2_127_3477_n1545, DP_OP_425J2_127_3477_n1544,
         DP_OP_425J2_127_3477_n1543, DP_OP_425J2_127_3477_n1542,
         DP_OP_425J2_127_3477_n1541, DP_OP_425J2_127_3477_n1540,
         DP_OP_425J2_127_3477_n1539, DP_OP_425J2_127_3477_n1538,
         DP_OP_425J2_127_3477_n1537, DP_OP_425J2_127_3477_n1536,
         DP_OP_425J2_127_3477_n1535, DP_OP_425J2_127_3477_n1534,
         DP_OP_425J2_127_3477_n1533, DP_OP_425J2_127_3477_n1532,
         DP_OP_425J2_127_3477_n1531, DP_OP_425J2_127_3477_n1530,
         DP_OP_425J2_127_3477_n1529, DP_OP_425J2_127_3477_n1528,
         DP_OP_425J2_127_3477_n1527, DP_OP_425J2_127_3477_n1526,
         DP_OP_425J2_127_3477_n1525, DP_OP_425J2_127_3477_n1524,
         DP_OP_425J2_127_3477_n1523, DP_OP_425J2_127_3477_n1522,
         DP_OP_425J2_127_3477_n1521, DP_OP_425J2_127_3477_n1520,
         DP_OP_425J2_127_3477_n1519, DP_OP_425J2_127_3477_n1518,
         DP_OP_425J2_127_3477_n1517, DP_OP_425J2_127_3477_n1516,
         DP_OP_425J2_127_3477_n1515, DP_OP_425J2_127_3477_n1514,
         DP_OP_425J2_127_3477_n1513, DP_OP_425J2_127_3477_n1512,
         DP_OP_425J2_127_3477_n1511, DP_OP_425J2_127_3477_n1510,
         DP_OP_425J2_127_3477_n1509, DP_OP_425J2_127_3477_n1508,
         DP_OP_425J2_127_3477_n1507, DP_OP_425J2_127_3477_n1506,
         DP_OP_425J2_127_3477_n1505, DP_OP_425J2_127_3477_n1504,
         DP_OP_425J2_127_3477_n1503, DP_OP_425J2_127_3477_n1502,
         DP_OP_425J2_127_3477_n1501, DP_OP_425J2_127_3477_n1500,
         DP_OP_425J2_127_3477_n1499, DP_OP_425J2_127_3477_n1498,
         DP_OP_425J2_127_3477_n1497, DP_OP_425J2_127_3477_n1496,
         DP_OP_425J2_127_3477_n1495, DP_OP_425J2_127_3477_n1494,
         DP_OP_425J2_127_3477_n1493, DP_OP_425J2_127_3477_n1492,
         DP_OP_425J2_127_3477_n1491, DP_OP_425J2_127_3477_n1490,
         DP_OP_425J2_127_3477_n1489, DP_OP_425J2_127_3477_n1488,
         DP_OP_425J2_127_3477_n1487, DP_OP_425J2_127_3477_n1486,
         DP_OP_425J2_127_3477_n1485, DP_OP_425J2_127_3477_n1484,
         DP_OP_425J2_127_3477_n1483, DP_OP_425J2_127_3477_n1482,
         DP_OP_425J2_127_3477_n1481, DP_OP_425J2_127_3477_n1480,
         DP_OP_425J2_127_3477_n1479, DP_OP_425J2_127_3477_n1478,
         DP_OP_425J2_127_3477_n1477, DP_OP_425J2_127_3477_n1476,
         DP_OP_425J2_127_3477_n1475, DP_OP_425J2_127_3477_n1474,
         DP_OP_425J2_127_3477_n1473, DP_OP_425J2_127_3477_n1472,
         DP_OP_425J2_127_3477_n1471, DP_OP_425J2_127_3477_n1470,
         DP_OP_425J2_127_3477_n1469, DP_OP_425J2_127_3477_n1468,
         DP_OP_425J2_127_3477_n1467, DP_OP_425J2_127_3477_n1466,
         DP_OP_425J2_127_3477_n1465, DP_OP_425J2_127_3477_n1464,
         DP_OP_425J2_127_3477_n1463, DP_OP_425J2_127_3477_n1462,
         DP_OP_425J2_127_3477_n1461, DP_OP_425J2_127_3477_n1460,
         DP_OP_425J2_127_3477_n1459, DP_OP_425J2_127_3477_n1458,
         DP_OP_425J2_127_3477_n1457, DP_OP_425J2_127_3477_n1456,
         DP_OP_425J2_127_3477_n1455, DP_OP_425J2_127_3477_n1454,
         DP_OP_425J2_127_3477_n1453, DP_OP_425J2_127_3477_n1452,
         DP_OP_425J2_127_3477_n1451, DP_OP_425J2_127_3477_n1450,
         DP_OP_425J2_127_3477_n1449, DP_OP_425J2_127_3477_n1448,
         DP_OP_425J2_127_3477_n1447, DP_OP_425J2_127_3477_n1446,
         DP_OP_425J2_127_3477_n1445, DP_OP_425J2_127_3477_n1444,
         DP_OP_425J2_127_3477_n1443, DP_OP_425J2_127_3477_n1442,
         DP_OP_425J2_127_3477_n1441, DP_OP_425J2_127_3477_n1440,
         DP_OP_425J2_127_3477_n1439, DP_OP_425J2_127_3477_n1438,
         DP_OP_425J2_127_3477_n1437, DP_OP_425J2_127_3477_n1436,
         DP_OP_425J2_127_3477_n1435, DP_OP_425J2_127_3477_n1434,
         DP_OP_425J2_127_3477_n1433, DP_OP_425J2_127_3477_n1432,
         DP_OP_425J2_127_3477_n1431, DP_OP_425J2_127_3477_n1430,
         DP_OP_425J2_127_3477_n1429, DP_OP_425J2_127_3477_n1428,
         DP_OP_425J2_127_3477_n1427, DP_OP_425J2_127_3477_n1426,
         DP_OP_425J2_127_3477_n1425, DP_OP_425J2_127_3477_n1424,
         DP_OP_425J2_127_3477_n1423, DP_OP_425J2_127_3477_n1422,
         DP_OP_425J2_127_3477_n1421, DP_OP_425J2_127_3477_n1420,
         DP_OP_425J2_127_3477_n1419, DP_OP_425J2_127_3477_n1418,
         DP_OP_425J2_127_3477_n1417, DP_OP_425J2_127_3477_n1416,
         DP_OP_425J2_127_3477_n1415, DP_OP_425J2_127_3477_n1414,
         DP_OP_425J2_127_3477_n1413, DP_OP_425J2_127_3477_n1412,
         DP_OP_425J2_127_3477_n1411, DP_OP_425J2_127_3477_n1410,
         DP_OP_425J2_127_3477_n1409, DP_OP_425J2_127_3477_n1408,
         DP_OP_425J2_127_3477_n1407, DP_OP_425J2_127_3477_n1406,
         DP_OP_425J2_127_3477_n1405, DP_OP_425J2_127_3477_n1404,
         DP_OP_425J2_127_3477_n1403, DP_OP_425J2_127_3477_n1402,
         DP_OP_425J2_127_3477_n1401, DP_OP_425J2_127_3477_n1400,
         DP_OP_425J2_127_3477_n1399, DP_OP_425J2_127_3477_n1398,
         DP_OP_425J2_127_3477_n1397, DP_OP_425J2_127_3477_n1396,
         DP_OP_425J2_127_3477_n1395, DP_OP_425J2_127_3477_n1394,
         DP_OP_425J2_127_3477_n1393, DP_OP_425J2_127_3477_n1392,
         DP_OP_425J2_127_3477_n1391, DP_OP_425J2_127_3477_n1390,
         DP_OP_425J2_127_3477_n1389, DP_OP_425J2_127_3477_n1388,
         DP_OP_425J2_127_3477_n1387, DP_OP_425J2_127_3477_n1386,
         DP_OP_425J2_127_3477_n1385, DP_OP_425J2_127_3477_n1384,
         DP_OP_425J2_127_3477_n1383, DP_OP_425J2_127_3477_n1382,
         DP_OP_425J2_127_3477_n1381, DP_OP_425J2_127_3477_n1380,
         DP_OP_425J2_127_3477_n1379, DP_OP_425J2_127_3477_n1378,
         DP_OP_425J2_127_3477_n1377, DP_OP_425J2_127_3477_n1376,
         DP_OP_425J2_127_3477_n1375, DP_OP_425J2_127_3477_n1374,
         DP_OP_425J2_127_3477_n1373, DP_OP_425J2_127_3477_n1372,
         DP_OP_425J2_127_3477_n1371, DP_OP_425J2_127_3477_n1370,
         DP_OP_425J2_127_3477_n1369, DP_OP_425J2_127_3477_n1368,
         DP_OP_425J2_127_3477_n1367, DP_OP_425J2_127_3477_n1366,
         DP_OP_425J2_127_3477_n1365, DP_OP_425J2_127_3477_n1364,
         DP_OP_425J2_127_3477_n1363, DP_OP_425J2_127_3477_n1362,
         DP_OP_425J2_127_3477_n1361, DP_OP_425J2_127_3477_n1360,
         DP_OP_425J2_127_3477_n1359, DP_OP_425J2_127_3477_n1358,
         DP_OP_425J2_127_3477_n1357, DP_OP_425J2_127_3477_n1356,
         DP_OP_425J2_127_3477_n1355, DP_OP_425J2_127_3477_n1354,
         DP_OP_425J2_127_3477_n1353, DP_OP_425J2_127_3477_n1352,
         DP_OP_425J2_127_3477_n1351, DP_OP_425J2_127_3477_n1350,
         DP_OP_425J2_127_3477_n1349, DP_OP_425J2_127_3477_n1348,
         DP_OP_425J2_127_3477_n1347, DP_OP_425J2_127_3477_n1346,
         DP_OP_425J2_127_3477_n1345, DP_OP_425J2_127_3477_n1344,
         DP_OP_425J2_127_3477_n1343, DP_OP_425J2_127_3477_n1342,
         DP_OP_425J2_127_3477_n1341, DP_OP_425J2_127_3477_n1340,
         DP_OP_425J2_127_3477_n1339, DP_OP_425J2_127_3477_n1338,
         DP_OP_425J2_127_3477_n1337, DP_OP_425J2_127_3477_n1336,
         DP_OP_425J2_127_3477_n1335, DP_OP_425J2_127_3477_n1334,
         DP_OP_425J2_127_3477_n1333, DP_OP_425J2_127_3477_n1332,
         DP_OP_425J2_127_3477_n1331, DP_OP_425J2_127_3477_n1330,
         DP_OP_425J2_127_3477_n1329, DP_OP_425J2_127_3477_n1328,
         DP_OP_425J2_127_3477_n1327, DP_OP_425J2_127_3477_n1326,
         DP_OP_425J2_127_3477_n1325, DP_OP_425J2_127_3477_n1324,
         DP_OP_425J2_127_3477_n1323, DP_OP_425J2_127_3477_n1322,
         DP_OP_425J2_127_3477_n1321, DP_OP_425J2_127_3477_n1320,
         DP_OP_425J2_127_3477_n1319, DP_OP_425J2_127_3477_n1318,
         DP_OP_425J2_127_3477_n1317, DP_OP_425J2_127_3477_n1316,
         DP_OP_425J2_127_3477_n1315, DP_OP_425J2_127_3477_n1314,
         DP_OP_425J2_127_3477_n1313, DP_OP_425J2_127_3477_n1312,
         DP_OP_425J2_127_3477_n1311, DP_OP_425J2_127_3477_n1310,
         DP_OP_425J2_127_3477_n1309, DP_OP_425J2_127_3477_n1308,
         DP_OP_425J2_127_3477_n1307, DP_OP_425J2_127_3477_n1306,
         DP_OP_425J2_127_3477_n1305, DP_OP_425J2_127_3477_n1304,
         DP_OP_425J2_127_3477_n1303, DP_OP_425J2_127_3477_n1302,
         DP_OP_425J2_127_3477_n1301, DP_OP_425J2_127_3477_n1300,
         DP_OP_425J2_127_3477_n1299, DP_OP_425J2_127_3477_n1298,
         DP_OP_425J2_127_3477_n1297, DP_OP_425J2_127_3477_n1296,
         DP_OP_425J2_127_3477_n1295, DP_OP_425J2_127_3477_n1294,
         DP_OP_425J2_127_3477_n1293, DP_OP_425J2_127_3477_n1292,
         DP_OP_425J2_127_3477_n1291, DP_OP_425J2_127_3477_n1290,
         DP_OP_425J2_127_3477_n1289, DP_OP_425J2_127_3477_n1288,
         DP_OP_425J2_127_3477_n1287, DP_OP_425J2_127_3477_n1286,
         DP_OP_425J2_127_3477_n1285, DP_OP_425J2_127_3477_n1284,
         DP_OP_425J2_127_3477_n1283, DP_OP_425J2_127_3477_n1282,
         DP_OP_425J2_127_3477_n1281, DP_OP_425J2_127_3477_n1280,
         DP_OP_425J2_127_3477_n1279, DP_OP_425J2_127_3477_n1278,
         DP_OP_425J2_127_3477_n1277, DP_OP_425J2_127_3477_n1276,
         DP_OP_425J2_127_3477_n1275, DP_OP_425J2_127_3477_n1274,
         DP_OP_425J2_127_3477_n1273, DP_OP_425J2_127_3477_n1272,
         DP_OP_425J2_127_3477_n1271, DP_OP_425J2_127_3477_n1270,
         DP_OP_425J2_127_3477_n1269, DP_OP_425J2_127_3477_n1268,
         DP_OP_425J2_127_3477_n1267, DP_OP_425J2_127_3477_n1266,
         DP_OP_425J2_127_3477_n1265, DP_OP_425J2_127_3477_n1264,
         DP_OP_425J2_127_3477_n1263, DP_OP_425J2_127_3477_n1262,
         DP_OP_425J2_127_3477_n1261, DP_OP_425J2_127_3477_n1260,
         DP_OP_425J2_127_3477_n1259, DP_OP_425J2_127_3477_n1258,
         DP_OP_425J2_127_3477_n1257, DP_OP_425J2_127_3477_n1256,
         DP_OP_425J2_127_3477_n1255, DP_OP_425J2_127_3477_n1254,
         DP_OP_425J2_127_3477_n1253, DP_OP_425J2_127_3477_n1252,
         DP_OP_425J2_127_3477_n1251, DP_OP_425J2_127_3477_n1250,
         DP_OP_425J2_127_3477_n1249, DP_OP_425J2_127_3477_n1248,
         DP_OP_425J2_127_3477_n1247, DP_OP_425J2_127_3477_n1246,
         DP_OP_425J2_127_3477_n1245, DP_OP_425J2_127_3477_n1244,
         DP_OP_425J2_127_3477_n1243, DP_OP_425J2_127_3477_n1242,
         DP_OP_425J2_127_3477_n1241, DP_OP_425J2_127_3477_n1240,
         DP_OP_425J2_127_3477_n1239, DP_OP_425J2_127_3477_n1238,
         DP_OP_425J2_127_3477_n1237, DP_OP_425J2_127_3477_n1236,
         DP_OP_425J2_127_3477_n1235, DP_OP_425J2_127_3477_n1234,
         DP_OP_425J2_127_3477_n1233, DP_OP_425J2_127_3477_n1232,
         DP_OP_425J2_127_3477_n1231, DP_OP_425J2_127_3477_n1230,
         DP_OP_425J2_127_3477_n1229, DP_OP_425J2_127_3477_n1228,
         DP_OP_425J2_127_3477_n1227, DP_OP_425J2_127_3477_n1226,
         DP_OP_425J2_127_3477_n1225, DP_OP_425J2_127_3477_n1224,
         DP_OP_425J2_127_3477_n1223, DP_OP_425J2_127_3477_n1222,
         DP_OP_425J2_127_3477_n1221, DP_OP_425J2_127_3477_n1220,
         DP_OP_425J2_127_3477_n1219, DP_OP_425J2_127_3477_n1218,
         DP_OP_425J2_127_3477_n1217, DP_OP_425J2_127_3477_n1216,
         DP_OP_425J2_127_3477_n1215, DP_OP_425J2_127_3477_n1214,
         DP_OP_425J2_127_3477_n1213, DP_OP_425J2_127_3477_n1212,
         DP_OP_425J2_127_3477_n1211, DP_OP_425J2_127_3477_n1210,
         DP_OP_425J2_127_3477_n1209, DP_OP_425J2_127_3477_n1208,
         DP_OP_425J2_127_3477_n1207, DP_OP_425J2_127_3477_n1206,
         DP_OP_425J2_127_3477_n1205, DP_OP_425J2_127_3477_n1204,
         DP_OP_425J2_127_3477_n1203, DP_OP_425J2_127_3477_n1202,
         DP_OP_425J2_127_3477_n1201, DP_OP_425J2_127_3477_n1200,
         DP_OP_425J2_127_3477_n1199, DP_OP_425J2_127_3477_n1198,
         DP_OP_425J2_127_3477_n1197, DP_OP_425J2_127_3477_n1196,
         DP_OP_425J2_127_3477_n1195, DP_OP_425J2_127_3477_n1194,
         DP_OP_425J2_127_3477_n1193, DP_OP_425J2_127_3477_n1192,
         DP_OP_425J2_127_3477_n1191, DP_OP_425J2_127_3477_n1190,
         DP_OP_425J2_127_3477_n1189, DP_OP_425J2_127_3477_n1188,
         DP_OP_425J2_127_3477_n1187, DP_OP_425J2_127_3477_n1186,
         DP_OP_425J2_127_3477_n1185, DP_OP_425J2_127_3477_n1184,
         DP_OP_425J2_127_3477_n1183, DP_OP_425J2_127_3477_n1182,
         DP_OP_425J2_127_3477_n1181, DP_OP_425J2_127_3477_n1180,
         DP_OP_425J2_127_3477_n1179, DP_OP_425J2_127_3477_n1178,
         DP_OP_425J2_127_3477_n1177, DP_OP_425J2_127_3477_n1176,
         DP_OP_425J2_127_3477_n1175, DP_OP_425J2_127_3477_n1174,
         DP_OP_425J2_127_3477_n1173, DP_OP_425J2_127_3477_n1172,
         DP_OP_425J2_127_3477_n1171, DP_OP_425J2_127_3477_n1170,
         DP_OP_425J2_127_3477_n1169, DP_OP_425J2_127_3477_n1168,
         DP_OP_425J2_127_3477_n1167, DP_OP_425J2_127_3477_n1166,
         DP_OP_425J2_127_3477_n1165, DP_OP_425J2_127_3477_n1164,
         DP_OP_425J2_127_3477_n1163, DP_OP_425J2_127_3477_n1162,
         DP_OP_425J2_127_3477_n1161, DP_OP_425J2_127_3477_n1160,
         DP_OP_425J2_127_3477_n1159, DP_OP_425J2_127_3477_n1158,
         DP_OP_425J2_127_3477_n1157, DP_OP_425J2_127_3477_n1156,
         DP_OP_425J2_127_3477_n1155, DP_OP_425J2_127_3477_n1154,
         DP_OP_425J2_127_3477_n1153, DP_OP_425J2_127_3477_n1152,
         DP_OP_425J2_127_3477_n1151, DP_OP_425J2_127_3477_n1150,
         DP_OP_425J2_127_3477_n1149, DP_OP_425J2_127_3477_n1148,
         DP_OP_425J2_127_3477_n1147, DP_OP_425J2_127_3477_n1146,
         DP_OP_425J2_127_3477_n1145, DP_OP_425J2_127_3477_n1144,
         DP_OP_425J2_127_3477_n1143, DP_OP_425J2_127_3477_n1142,
         DP_OP_425J2_127_3477_n1141, DP_OP_425J2_127_3477_n1140,
         DP_OP_425J2_127_3477_n1139, DP_OP_425J2_127_3477_n1138,
         DP_OP_425J2_127_3477_n1137, DP_OP_425J2_127_3477_n1136,
         DP_OP_425J2_127_3477_n1135, DP_OP_425J2_127_3477_n1134,
         DP_OP_425J2_127_3477_n1133, DP_OP_425J2_127_3477_n1132,
         DP_OP_425J2_127_3477_n1131, DP_OP_425J2_127_3477_n1130,
         DP_OP_425J2_127_3477_n1129, DP_OP_425J2_127_3477_n1128,
         DP_OP_425J2_127_3477_n1127, DP_OP_425J2_127_3477_n1126,
         DP_OP_425J2_127_3477_n1125, DP_OP_425J2_127_3477_n1124,
         DP_OP_425J2_127_3477_n1123, DP_OP_425J2_127_3477_n1122,
         DP_OP_425J2_127_3477_n1121, DP_OP_425J2_127_3477_n1120,
         DP_OP_425J2_127_3477_n1119, DP_OP_425J2_127_3477_n1118,
         DP_OP_425J2_127_3477_n1117, DP_OP_425J2_127_3477_n1116,
         DP_OP_425J2_127_3477_n1115, DP_OP_425J2_127_3477_n1114,
         DP_OP_425J2_127_3477_n1113, DP_OP_425J2_127_3477_n1112,
         DP_OP_425J2_127_3477_n1111, DP_OP_425J2_127_3477_n1110,
         DP_OP_425J2_127_3477_n1109, DP_OP_425J2_127_3477_n1108,
         DP_OP_425J2_127_3477_n1107, DP_OP_425J2_127_3477_n1106,
         DP_OP_425J2_127_3477_n1105, DP_OP_425J2_127_3477_n1104,
         DP_OP_425J2_127_3477_n1103, DP_OP_425J2_127_3477_n1102,
         DP_OP_425J2_127_3477_n1101, DP_OP_425J2_127_3477_n1100,
         DP_OP_425J2_127_3477_n1099, DP_OP_425J2_127_3477_n1098,
         DP_OP_425J2_127_3477_n1097, DP_OP_425J2_127_3477_n1096,
         DP_OP_425J2_127_3477_n1095, DP_OP_425J2_127_3477_n1094,
         DP_OP_425J2_127_3477_n1093, DP_OP_425J2_127_3477_n1092,
         DP_OP_425J2_127_3477_n1091, DP_OP_425J2_127_3477_n1090,
         DP_OP_425J2_127_3477_n1089, DP_OP_425J2_127_3477_n1088,
         DP_OP_425J2_127_3477_n1087, DP_OP_425J2_127_3477_n1086,
         DP_OP_425J2_127_3477_n1085, DP_OP_425J2_127_3477_n1084,
         DP_OP_425J2_127_3477_n1083, DP_OP_425J2_127_3477_n1082,
         DP_OP_425J2_127_3477_n1081, DP_OP_425J2_127_3477_n1080,
         DP_OP_425J2_127_3477_n1079, DP_OP_425J2_127_3477_n1078,
         DP_OP_425J2_127_3477_n1077, DP_OP_425J2_127_3477_n1076,
         DP_OP_425J2_127_3477_n1075, DP_OP_425J2_127_3477_n1074,
         DP_OP_425J2_127_3477_n1073, DP_OP_425J2_127_3477_n1072,
         DP_OP_425J2_127_3477_n1071, DP_OP_425J2_127_3477_n1070,
         DP_OP_425J2_127_3477_n1069, DP_OP_425J2_127_3477_n1068,
         DP_OP_425J2_127_3477_n1067, DP_OP_425J2_127_3477_n1066,
         DP_OP_425J2_127_3477_n1065, DP_OP_425J2_127_3477_n1064,
         DP_OP_425J2_127_3477_n1063, DP_OP_425J2_127_3477_n1062,
         DP_OP_425J2_127_3477_n1061, DP_OP_425J2_127_3477_n1060,
         DP_OP_425J2_127_3477_n1059, DP_OP_425J2_127_3477_n1058,
         DP_OP_425J2_127_3477_n1057, DP_OP_425J2_127_3477_n1056,
         DP_OP_425J2_127_3477_n1055, DP_OP_425J2_127_3477_n1054,
         DP_OP_425J2_127_3477_n1053, DP_OP_425J2_127_3477_n1052,
         DP_OP_425J2_127_3477_n1051, DP_OP_425J2_127_3477_n1050,
         DP_OP_425J2_127_3477_n1049, DP_OP_425J2_127_3477_n1048,
         DP_OP_425J2_127_3477_n1047, DP_OP_425J2_127_3477_n1046,
         DP_OP_425J2_127_3477_n1045, DP_OP_425J2_127_3477_n1044,
         DP_OP_425J2_127_3477_n1043, DP_OP_425J2_127_3477_n1042,
         DP_OP_425J2_127_3477_n1041, DP_OP_425J2_127_3477_n1040,
         DP_OP_425J2_127_3477_n1039, DP_OP_425J2_127_3477_n1038,
         DP_OP_425J2_127_3477_n1037, DP_OP_425J2_127_3477_n1036,
         DP_OP_425J2_127_3477_n1035, DP_OP_425J2_127_3477_n1034,
         DP_OP_425J2_127_3477_n1033, DP_OP_425J2_127_3477_n1032,
         DP_OP_425J2_127_3477_n1031, DP_OP_425J2_127_3477_n1030,
         DP_OP_425J2_127_3477_n1029, DP_OP_425J2_127_3477_n1028,
         DP_OP_425J2_127_3477_n1027, DP_OP_425J2_127_3477_n1026,
         DP_OP_425J2_127_3477_n1025, DP_OP_425J2_127_3477_n1024,
         DP_OP_425J2_127_3477_n1023, DP_OP_425J2_127_3477_n1022,
         DP_OP_425J2_127_3477_n1021, DP_OP_425J2_127_3477_n1020,
         DP_OP_425J2_127_3477_n1019, DP_OP_425J2_127_3477_n1018,
         DP_OP_425J2_127_3477_n1017, DP_OP_425J2_127_3477_n1016,
         DP_OP_425J2_127_3477_n1015, DP_OP_425J2_127_3477_n1014,
         DP_OP_425J2_127_3477_n1013, DP_OP_425J2_127_3477_n1012,
         DP_OP_425J2_127_3477_n1011, DP_OP_425J2_127_3477_n1010,
         DP_OP_425J2_127_3477_n1009, DP_OP_425J2_127_3477_n1008,
         DP_OP_425J2_127_3477_n1007, DP_OP_425J2_127_3477_n1006,
         DP_OP_425J2_127_3477_n1005, DP_OP_425J2_127_3477_n1004,
         DP_OP_425J2_127_3477_n1003, DP_OP_425J2_127_3477_n1002,
         DP_OP_425J2_127_3477_n1001, DP_OP_425J2_127_3477_n1000,
         DP_OP_425J2_127_3477_n999, DP_OP_425J2_127_3477_n998,
         DP_OP_425J2_127_3477_n997, DP_OP_425J2_127_3477_n996,
         DP_OP_425J2_127_3477_n995, DP_OP_425J2_127_3477_n994,
         DP_OP_425J2_127_3477_n993, DP_OP_425J2_127_3477_n992,
         DP_OP_425J2_127_3477_n991, DP_OP_425J2_127_3477_n990,
         DP_OP_425J2_127_3477_n989, DP_OP_425J2_127_3477_n988,
         DP_OP_425J2_127_3477_n987, DP_OP_425J2_127_3477_n986,
         DP_OP_425J2_127_3477_n985, DP_OP_425J2_127_3477_n984,
         DP_OP_425J2_127_3477_n983, DP_OP_425J2_127_3477_n982,
         DP_OP_425J2_127_3477_n981, DP_OP_425J2_127_3477_n980,
         DP_OP_425J2_127_3477_n979, DP_OP_425J2_127_3477_n978,
         DP_OP_425J2_127_3477_n977, DP_OP_425J2_127_3477_n976,
         DP_OP_425J2_127_3477_n975, DP_OP_425J2_127_3477_n974,
         DP_OP_425J2_127_3477_n973, DP_OP_425J2_127_3477_n972,
         DP_OP_425J2_127_3477_n971, DP_OP_425J2_127_3477_n970,
         DP_OP_425J2_127_3477_n969, DP_OP_425J2_127_3477_n968,
         DP_OP_425J2_127_3477_n967, DP_OP_425J2_127_3477_n966,
         DP_OP_425J2_127_3477_n965, DP_OP_425J2_127_3477_n964,
         DP_OP_425J2_127_3477_n963, DP_OP_425J2_127_3477_n962,
         DP_OP_425J2_127_3477_n961, DP_OP_425J2_127_3477_n960,
         DP_OP_425J2_127_3477_n959, DP_OP_425J2_127_3477_n958,
         DP_OP_425J2_127_3477_n957, DP_OP_425J2_127_3477_n956,
         DP_OP_425J2_127_3477_n955, DP_OP_425J2_127_3477_n954,
         DP_OP_425J2_127_3477_n953, DP_OP_425J2_127_3477_n952,
         DP_OP_425J2_127_3477_n951, DP_OP_425J2_127_3477_n950,
         DP_OP_425J2_127_3477_n949, DP_OP_425J2_127_3477_n948,
         DP_OP_425J2_127_3477_n947, DP_OP_425J2_127_3477_n946,
         DP_OP_425J2_127_3477_n945, DP_OP_425J2_127_3477_n944,
         DP_OP_425J2_127_3477_n943, DP_OP_425J2_127_3477_n942,
         DP_OP_425J2_127_3477_n941, DP_OP_425J2_127_3477_n940,
         DP_OP_425J2_127_3477_n939, DP_OP_425J2_127_3477_n938,
         DP_OP_425J2_127_3477_n937, DP_OP_425J2_127_3477_n936,
         DP_OP_425J2_127_3477_n935, DP_OP_425J2_127_3477_n934,
         DP_OP_425J2_127_3477_n933, DP_OP_425J2_127_3477_n932,
         DP_OP_425J2_127_3477_n931, DP_OP_425J2_127_3477_n930,
         DP_OP_425J2_127_3477_n929, DP_OP_425J2_127_3477_n928,
         DP_OP_425J2_127_3477_n927, DP_OP_425J2_127_3477_n926,
         DP_OP_425J2_127_3477_n925, DP_OP_425J2_127_3477_n924,
         DP_OP_425J2_127_3477_n923, DP_OP_425J2_127_3477_n922,
         DP_OP_425J2_127_3477_n921, DP_OP_425J2_127_3477_n920,
         DP_OP_425J2_127_3477_n919, DP_OP_425J2_127_3477_n918,
         DP_OP_425J2_127_3477_n917, DP_OP_425J2_127_3477_n916,
         DP_OP_425J2_127_3477_n915, DP_OP_425J2_127_3477_n914,
         DP_OP_425J2_127_3477_n913, DP_OP_425J2_127_3477_n912,
         DP_OP_425J2_127_3477_n911, DP_OP_425J2_127_3477_n910,
         DP_OP_425J2_127_3477_n909, DP_OP_425J2_127_3477_n908,
         DP_OP_425J2_127_3477_n907, DP_OP_425J2_127_3477_n906,
         DP_OP_425J2_127_3477_n905, DP_OP_425J2_127_3477_n904,
         DP_OP_425J2_127_3477_n903, DP_OP_425J2_127_3477_n902,
         DP_OP_425J2_127_3477_n901, DP_OP_425J2_127_3477_n900,
         DP_OP_425J2_127_3477_n899, DP_OP_425J2_127_3477_n898,
         DP_OP_425J2_127_3477_n897, DP_OP_425J2_127_3477_n896,
         DP_OP_425J2_127_3477_n895, DP_OP_425J2_127_3477_n894,
         DP_OP_425J2_127_3477_n893, DP_OP_425J2_127_3477_n892,
         DP_OP_425J2_127_3477_n891, DP_OP_425J2_127_3477_n890,
         DP_OP_425J2_127_3477_n889, DP_OP_425J2_127_3477_n888,
         DP_OP_425J2_127_3477_n887, DP_OP_425J2_127_3477_n886,
         DP_OP_425J2_127_3477_n885, DP_OP_425J2_127_3477_n884,
         DP_OP_425J2_127_3477_n883, DP_OP_425J2_127_3477_n882,
         DP_OP_425J2_127_3477_n881, DP_OP_425J2_127_3477_n880,
         DP_OP_425J2_127_3477_n879, DP_OP_425J2_127_3477_n878,
         DP_OP_425J2_127_3477_n877, DP_OP_425J2_127_3477_n876,
         DP_OP_425J2_127_3477_n875, DP_OP_425J2_127_3477_n874,
         DP_OP_425J2_127_3477_n873, DP_OP_425J2_127_3477_n872,
         DP_OP_425J2_127_3477_n871, DP_OP_425J2_127_3477_n870,
         DP_OP_425J2_127_3477_n869, DP_OP_425J2_127_3477_n868,
         DP_OP_425J2_127_3477_n867, DP_OP_425J2_127_3477_n866,
         DP_OP_425J2_127_3477_n865, DP_OP_425J2_127_3477_n864,
         DP_OP_425J2_127_3477_n863, DP_OP_425J2_127_3477_n862,
         DP_OP_425J2_127_3477_n861, DP_OP_425J2_127_3477_n860,
         DP_OP_425J2_127_3477_n859, DP_OP_425J2_127_3477_n858,
         DP_OP_425J2_127_3477_n857, DP_OP_425J2_127_3477_n856,
         DP_OP_425J2_127_3477_n855, DP_OP_425J2_127_3477_n854,
         DP_OP_425J2_127_3477_n853, DP_OP_425J2_127_3477_n852,
         DP_OP_425J2_127_3477_n851, DP_OP_425J2_127_3477_n850,
         DP_OP_425J2_127_3477_n849, DP_OP_425J2_127_3477_n848,
         DP_OP_425J2_127_3477_n847, DP_OP_425J2_127_3477_n846,
         DP_OP_425J2_127_3477_n845, DP_OP_425J2_127_3477_n844,
         DP_OP_425J2_127_3477_n843, DP_OP_425J2_127_3477_n842,
         DP_OP_425J2_127_3477_n841, DP_OP_425J2_127_3477_n840,
         DP_OP_425J2_127_3477_n839, DP_OP_425J2_127_3477_n838,
         DP_OP_425J2_127_3477_n837, DP_OP_425J2_127_3477_n836,
         DP_OP_425J2_127_3477_n835, DP_OP_425J2_127_3477_n834,
         DP_OP_425J2_127_3477_n833, DP_OP_425J2_127_3477_n832,
         DP_OP_425J2_127_3477_n831, DP_OP_425J2_127_3477_n830,
         DP_OP_425J2_127_3477_n829, DP_OP_425J2_127_3477_n828,
         DP_OP_425J2_127_3477_n827, DP_OP_425J2_127_3477_n826,
         DP_OP_425J2_127_3477_n825, DP_OP_425J2_127_3477_n824,
         DP_OP_425J2_127_3477_n823, DP_OP_425J2_127_3477_n822,
         DP_OP_425J2_127_3477_n821, DP_OP_425J2_127_3477_n820,
         DP_OP_425J2_127_3477_n819, DP_OP_425J2_127_3477_n818,
         DP_OP_425J2_127_3477_n817, DP_OP_425J2_127_3477_n816,
         DP_OP_425J2_127_3477_n815, DP_OP_425J2_127_3477_n814,
         DP_OP_425J2_127_3477_n813, DP_OP_425J2_127_3477_n812,
         DP_OP_425J2_127_3477_n811, DP_OP_425J2_127_3477_n810,
         DP_OP_425J2_127_3477_n809, DP_OP_425J2_127_3477_n808,
         DP_OP_425J2_127_3477_n807, DP_OP_425J2_127_3477_n806,
         DP_OP_425J2_127_3477_n805, DP_OP_425J2_127_3477_n804,
         DP_OP_425J2_127_3477_n803, DP_OP_425J2_127_3477_n802,
         DP_OP_425J2_127_3477_n801, DP_OP_425J2_127_3477_n800,
         DP_OP_425J2_127_3477_n799, DP_OP_425J2_127_3477_n798,
         DP_OP_425J2_127_3477_n797, DP_OP_425J2_127_3477_n796,
         DP_OP_425J2_127_3477_n795, DP_OP_425J2_127_3477_n794,
         DP_OP_425J2_127_3477_n793, DP_OP_425J2_127_3477_n792,
         DP_OP_425J2_127_3477_n791, DP_OP_425J2_127_3477_n790,
         DP_OP_425J2_127_3477_n789, DP_OP_425J2_127_3477_n788,
         DP_OP_425J2_127_3477_n787, DP_OP_425J2_127_3477_n786,
         DP_OP_425J2_127_3477_n785, DP_OP_425J2_127_3477_n784,
         DP_OP_425J2_127_3477_n783, DP_OP_425J2_127_3477_n782,
         DP_OP_425J2_127_3477_n781, DP_OP_425J2_127_3477_n780,
         DP_OP_425J2_127_3477_n779, DP_OP_425J2_127_3477_n778,
         DP_OP_425J2_127_3477_n777, DP_OP_425J2_127_3477_n776,
         DP_OP_425J2_127_3477_n775, DP_OP_425J2_127_3477_n774,
         DP_OP_425J2_127_3477_n773, DP_OP_425J2_127_3477_n772,
         DP_OP_425J2_127_3477_n771, DP_OP_425J2_127_3477_n770,
         DP_OP_425J2_127_3477_n769, DP_OP_425J2_127_3477_n768,
         DP_OP_425J2_127_3477_n767, DP_OP_425J2_127_3477_n766,
         DP_OP_425J2_127_3477_n765, DP_OP_425J2_127_3477_n764,
         DP_OP_425J2_127_3477_n763, DP_OP_425J2_127_3477_n762,
         DP_OP_425J2_127_3477_n761, DP_OP_425J2_127_3477_n760,
         DP_OP_425J2_127_3477_n759, DP_OP_425J2_127_3477_n758,
         DP_OP_425J2_127_3477_n757, DP_OP_425J2_127_3477_n756,
         DP_OP_425J2_127_3477_n755, DP_OP_425J2_127_3477_n754,
         DP_OP_425J2_127_3477_n753, DP_OP_425J2_127_3477_n752,
         DP_OP_425J2_127_3477_n751, DP_OP_425J2_127_3477_n750,
         DP_OP_425J2_127_3477_n749, DP_OP_425J2_127_3477_n748,
         DP_OP_425J2_127_3477_n747, DP_OP_425J2_127_3477_n746,
         DP_OP_425J2_127_3477_n745, DP_OP_425J2_127_3477_n744,
         DP_OP_425J2_127_3477_n743, DP_OP_425J2_127_3477_n742,
         DP_OP_425J2_127_3477_n741, DP_OP_425J2_127_3477_n740,
         DP_OP_425J2_127_3477_n739, DP_OP_425J2_127_3477_n738,
         DP_OP_425J2_127_3477_n737, DP_OP_425J2_127_3477_n736,
         DP_OP_425J2_127_3477_n735, DP_OP_425J2_127_3477_n734,
         DP_OP_425J2_127_3477_n733, DP_OP_425J2_127_3477_n732,
         DP_OP_425J2_127_3477_n731, DP_OP_425J2_127_3477_n730,
         DP_OP_425J2_127_3477_n729, DP_OP_425J2_127_3477_n728,
         DP_OP_425J2_127_3477_n727, DP_OP_425J2_127_3477_n726,
         DP_OP_425J2_127_3477_n725, DP_OP_425J2_127_3477_n724,
         DP_OP_425J2_127_3477_n723, DP_OP_425J2_127_3477_n722,
         DP_OP_425J2_127_3477_n721, DP_OP_425J2_127_3477_n720,
         DP_OP_425J2_127_3477_n719, DP_OP_425J2_127_3477_n718,
         DP_OP_425J2_127_3477_n717, DP_OP_425J2_127_3477_n716,
         DP_OP_425J2_127_3477_n715, DP_OP_425J2_127_3477_n714,
         DP_OP_425J2_127_3477_n713, DP_OP_425J2_127_3477_n712,
         DP_OP_425J2_127_3477_n711, DP_OP_425J2_127_3477_n710,
         DP_OP_425J2_127_3477_n709, DP_OP_425J2_127_3477_n708,
         DP_OP_425J2_127_3477_n707, DP_OP_425J2_127_3477_n706,
         DP_OP_425J2_127_3477_n705, DP_OP_425J2_127_3477_n704,
         DP_OP_425J2_127_3477_n703, DP_OP_425J2_127_3477_n702,
         DP_OP_425J2_127_3477_n701, DP_OP_425J2_127_3477_n700,
         DP_OP_425J2_127_3477_n699, DP_OP_425J2_127_3477_n698,
         DP_OP_425J2_127_3477_n697, DP_OP_425J2_127_3477_n696,
         DP_OP_425J2_127_3477_n695, DP_OP_425J2_127_3477_n694,
         DP_OP_425J2_127_3477_n693, DP_OP_425J2_127_3477_n692,
         DP_OP_425J2_127_3477_n691, DP_OP_425J2_127_3477_n690,
         DP_OP_425J2_127_3477_n689, DP_OP_425J2_127_3477_n688,
         DP_OP_425J2_127_3477_n687, DP_OP_425J2_127_3477_n686,
         DP_OP_425J2_127_3477_n685, DP_OP_425J2_127_3477_n684,
         DP_OP_425J2_127_3477_n683, DP_OP_425J2_127_3477_n682,
         DP_OP_425J2_127_3477_n681, DP_OP_425J2_127_3477_n680,
         DP_OP_425J2_127_3477_n679, DP_OP_425J2_127_3477_n678,
         DP_OP_425J2_127_3477_n677, DP_OP_425J2_127_3477_n676,
         DP_OP_425J2_127_3477_n675, DP_OP_425J2_127_3477_n674,
         DP_OP_425J2_127_3477_n673, DP_OP_425J2_127_3477_n672,
         DP_OP_425J2_127_3477_n671, DP_OP_425J2_127_3477_n670,
         DP_OP_425J2_127_3477_n669, DP_OP_425J2_127_3477_n668,
         DP_OP_425J2_127_3477_n667, DP_OP_425J2_127_3477_n666,
         DP_OP_425J2_127_3477_n665, DP_OP_425J2_127_3477_n664,
         DP_OP_425J2_127_3477_n663, DP_OP_425J2_127_3477_n662,
         DP_OP_425J2_127_3477_n661, DP_OP_425J2_127_3477_n660,
         DP_OP_425J2_127_3477_n659, DP_OP_425J2_127_3477_n658,
         DP_OP_425J2_127_3477_n657, DP_OP_425J2_127_3477_n656,
         DP_OP_425J2_127_3477_n655, DP_OP_425J2_127_3477_n654,
         DP_OP_425J2_127_3477_n653, DP_OP_425J2_127_3477_n652,
         DP_OP_425J2_127_3477_n651, DP_OP_425J2_127_3477_n650,
         DP_OP_425J2_127_3477_n649, DP_OP_425J2_127_3477_n648,
         DP_OP_425J2_127_3477_n647, DP_OP_425J2_127_3477_n646,
         DP_OP_425J2_127_3477_n645, DP_OP_425J2_127_3477_n644,
         DP_OP_425J2_127_3477_n643, DP_OP_425J2_127_3477_n642,
         DP_OP_425J2_127_3477_n641, DP_OP_425J2_127_3477_n640,
         DP_OP_425J2_127_3477_n639, DP_OP_425J2_127_3477_n638,
         DP_OP_425J2_127_3477_n637, DP_OP_425J2_127_3477_n636,
         DP_OP_425J2_127_3477_n635, DP_OP_425J2_127_3477_n634,
         DP_OP_425J2_127_3477_n633, DP_OP_425J2_127_3477_n632,
         DP_OP_425J2_127_3477_n631, DP_OP_425J2_127_3477_n630,
         DP_OP_425J2_127_3477_n629, DP_OP_425J2_127_3477_n628,
         DP_OP_425J2_127_3477_n627, DP_OP_425J2_127_3477_n626,
         DP_OP_425J2_127_3477_n625, DP_OP_425J2_127_3477_n624,
         DP_OP_425J2_127_3477_n623, DP_OP_425J2_127_3477_n622,
         DP_OP_425J2_127_3477_n621, DP_OP_425J2_127_3477_n620,
         DP_OP_425J2_127_3477_n619, DP_OP_425J2_127_3477_n618,
         DP_OP_425J2_127_3477_n617, DP_OP_425J2_127_3477_n616,
         DP_OP_425J2_127_3477_n615, DP_OP_425J2_127_3477_n614,
         DP_OP_425J2_127_3477_n613, DP_OP_425J2_127_3477_n612,
         DP_OP_425J2_127_3477_n611, DP_OP_425J2_127_3477_n610,
         DP_OP_425J2_127_3477_n609, DP_OP_425J2_127_3477_n608,
         DP_OP_425J2_127_3477_n607, DP_OP_425J2_127_3477_n606,
         DP_OP_425J2_127_3477_n605, DP_OP_425J2_127_3477_n604,
         DP_OP_425J2_127_3477_n603, DP_OP_425J2_127_3477_n602,
         DP_OP_425J2_127_3477_n601, DP_OP_425J2_127_3477_n600,
         DP_OP_425J2_127_3477_n599, DP_OP_425J2_127_3477_n598,
         DP_OP_425J2_127_3477_n597, DP_OP_425J2_127_3477_n596,
         DP_OP_425J2_127_3477_n595, DP_OP_425J2_127_3477_n594,
         DP_OP_425J2_127_3477_n593, DP_OP_425J2_127_3477_n592,
         DP_OP_425J2_127_3477_n591, DP_OP_425J2_127_3477_n590,
         DP_OP_425J2_127_3477_n589, DP_OP_425J2_127_3477_n588,
         DP_OP_425J2_127_3477_n587, DP_OP_425J2_127_3477_n586,
         DP_OP_425J2_127_3477_n585, DP_OP_425J2_127_3477_n584,
         DP_OP_425J2_127_3477_n583, DP_OP_425J2_127_3477_n582,
         DP_OP_425J2_127_3477_n581, DP_OP_425J2_127_3477_n580,
         DP_OP_425J2_127_3477_n579, DP_OP_425J2_127_3477_n578,
         DP_OP_425J2_127_3477_n577, DP_OP_425J2_127_3477_n576,
         DP_OP_425J2_127_3477_n575, DP_OP_425J2_127_3477_n574,
         DP_OP_425J2_127_3477_n573, DP_OP_425J2_127_3477_n572,
         DP_OP_425J2_127_3477_n571, DP_OP_425J2_127_3477_n570,
         DP_OP_425J2_127_3477_n569, DP_OP_425J2_127_3477_n568,
         DP_OP_425J2_127_3477_n567, DP_OP_425J2_127_3477_n566,
         DP_OP_425J2_127_3477_n565, DP_OP_425J2_127_3477_n564,
         DP_OP_425J2_127_3477_n563, DP_OP_425J2_127_3477_n562,
         DP_OP_425J2_127_3477_n561, DP_OP_425J2_127_3477_n560,
         DP_OP_425J2_127_3477_n559, DP_OP_425J2_127_3477_n558,
         DP_OP_425J2_127_3477_n557, DP_OP_425J2_127_3477_n556,
         DP_OP_425J2_127_3477_n555, DP_OP_425J2_127_3477_n554,
         DP_OP_425J2_127_3477_n553, DP_OP_425J2_127_3477_n552,
         DP_OP_425J2_127_3477_n551, DP_OP_425J2_127_3477_n550,
         DP_OP_425J2_127_3477_n549, DP_OP_425J2_127_3477_n548,
         DP_OP_425J2_127_3477_n547, DP_OP_425J2_127_3477_n546,
         DP_OP_425J2_127_3477_n545, DP_OP_425J2_127_3477_n544,
         DP_OP_425J2_127_3477_n543, DP_OP_425J2_127_3477_n542,
         DP_OP_425J2_127_3477_n541, DP_OP_425J2_127_3477_n540,
         DP_OP_425J2_127_3477_n539, DP_OP_425J2_127_3477_n538,
         DP_OP_425J2_127_3477_n537, DP_OP_425J2_127_3477_n536,
         DP_OP_425J2_127_3477_n535, DP_OP_425J2_127_3477_n534,
         DP_OP_425J2_127_3477_n533, DP_OP_425J2_127_3477_n532,
         DP_OP_425J2_127_3477_n531, DP_OP_425J2_127_3477_n530,
         DP_OP_425J2_127_3477_n529, DP_OP_425J2_127_3477_n528,
         DP_OP_425J2_127_3477_n527, DP_OP_425J2_127_3477_n526,
         DP_OP_425J2_127_3477_n525, DP_OP_425J2_127_3477_n524,
         DP_OP_425J2_127_3477_n523, DP_OP_425J2_127_3477_n522,
         DP_OP_425J2_127_3477_n521, DP_OP_425J2_127_3477_n520,
         DP_OP_425J2_127_3477_n519, DP_OP_425J2_127_3477_n518,
         DP_OP_425J2_127_3477_n517, DP_OP_425J2_127_3477_n516,
         DP_OP_425J2_127_3477_n515, DP_OP_425J2_127_3477_n514,
         DP_OP_425J2_127_3477_n513, DP_OP_425J2_127_3477_n512,
         DP_OP_425J2_127_3477_n511, DP_OP_425J2_127_3477_n510,
         DP_OP_425J2_127_3477_n509, DP_OP_425J2_127_3477_n508,
         DP_OP_425J2_127_3477_n507, DP_OP_425J2_127_3477_n506,
         DP_OP_425J2_127_3477_n505, DP_OP_425J2_127_3477_n504,
         DP_OP_425J2_127_3477_n503, DP_OP_425J2_127_3477_n502,
         DP_OP_425J2_127_3477_n501, DP_OP_425J2_127_3477_n500,
         DP_OP_425J2_127_3477_n499, DP_OP_425J2_127_3477_n498,
         DP_OP_425J2_127_3477_n497, DP_OP_425J2_127_3477_n496,
         DP_OP_425J2_127_3477_n495, DP_OP_425J2_127_3477_n494,
         DP_OP_425J2_127_3477_n493, DP_OP_425J2_127_3477_n492,
         DP_OP_425J2_127_3477_n491, DP_OP_425J2_127_3477_n490,
         DP_OP_425J2_127_3477_n489, DP_OP_425J2_127_3477_n488,
         DP_OP_425J2_127_3477_n487, DP_OP_425J2_127_3477_n486,
         DP_OP_425J2_127_3477_n485, DP_OP_425J2_127_3477_n484,
         DP_OP_425J2_127_3477_n483, DP_OP_425J2_127_3477_n482,
         DP_OP_425J2_127_3477_n481, DP_OP_425J2_127_3477_n480,
         DP_OP_425J2_127_3477_n479, DP_OP_425J2_127_3477_n478,
         DP_OP_425J2_127_3477_n477, DP_OP_425J2_127_3477_n476,
         DP_OP_425J2_127_3477_n475, DP_OP_425J2_127_3477_n474,
         DP_OP_425J2_127_3477_n473, DP_OP_425J2_127_3477_n472,
         DP_OP_425J2_127_3477_n471, DP_OP_425J2_127_3477_n470,
         DP_OP_425J2_127_3477_n469, DP_OP_425J2_127_3477_n468,
         DP_OP_425J2_127_3477_n467, DP_OP_425J2_127_3477_n466,
         DP_OP_425J2_127_3477_n465, DP_OP_425J2_127_3477_n464,
         DP_OP_425J2_127_3477_n463, DP_OP_425J2_127_3477_n462,
         DP_OP_425J2_127_3477_n461, DP_OP_425J2_127_3477_n460,
         DP_OP_425J2_127_3477_n459, DP_OP_425J2_127_3477_n458,
         DP_OP_425J2_127_3477_n457, DP_OP_425J2_127_3477_n456,
         DP_OP_425J2_127_3477_n455, DP_OP_425J2_127_3477_n454,
         DP_OP_425J2_127_3477_n453, DP_OP_425J2_127_3477_n452,
         DP_OP_425J2_127_3477_n451, DP_OP_425J2_127_3477_n450,
         DP_OP_425J2_127_3477_n449, DP_OP_425J2_127_3477_n448,
         DP_OP_425J2_127_3477_n447, DP_OP_425J2_127_3477_n446,
         DP_OP_425J2_127_3477_n445, DP_OP_425J2_127_3477_n444,
         DP_OP_425J2_127_3477_n443, DP_OP_425J2_127_3477_n442,
         DP_OP_425J2_127_3477_n441, DP_OP_425J2_127_3477_n440,
         DP_OP_425J2_127_3477_n439, DP_OP_425J2_127_3477_n438,
         DP_OP_425J2_127_3477_n437, DP_OP_425J2_127_3477_n436,
         DP_OP_425J2_127_3477_n435, DP_OP_425J2_127_3477_n434,
         DP_OP_425J2_127_3477_n433, DP_OP_425J2_127_3477_n432,
         DP_OP_425J2_127_3477_n431, DP_OP_425J2_127_3477_n430,
         DP_OP_425J2_127_3477_n429, DP_OP_425J2_127_3477_n428,
         DP_OP_425J2_127_3477_n427, DP_OP_425J2_127_3477_n426,
         DP_OP_425J2_127_3477_n425, DP_OP_425J2_127_3477_n424,
         DP_OP_425J2_127_3477_n423, DP_OP_425J2_127_3477_n422,
         DP_OP_425J2_127_3477_n421, DP_OP_425J2_127_3477_n420,
         DP_OP_425J2_127_3477_n419, DP_OP_425J2_127_3477_n418,
         DP_OP_425J2_127_3477_n417, DP_OP_425J2_127_3477_n416,
         DP_OP_425J2_127_3477_n415, DP_OP_425J2_127_3477_n414,
         DP_OP_425J2_127_3477_n413, DP_OP_425J2_127_3477_n412,
         DP_OP_425J2_127_3477_n411, DP_OP_425J2_127_3477_n410,
         DP_OP_425J2_127_3477_n409, DP_OP_425J2_127_3477_n408,
         DP_OP_425J2_127_3477_n407, DP_OP_425J2_127_3477_n406,
         DP_OP_425J2_127_3477_n405, DP_OP_425J2_127_3477_n404,
         DP_OP_425J2_127_3477_n403, DP_OP_425J2_127_3477_n402,
         DP_OP_425J2_127_3477_n401, DP_OP_425J2_127_3477_n400,
         DP_OP_425J2_127_3477_n399, DP_OP_425J2_127_3477_n398,
         DP_OP_425J2_127_3477_n397, DP_OP_425J2_127_3477_n396,
         DP_OP_425J2_127_3477_n395, DP_OP_425J2_127_3477_n394,
         DP_OP_425J2_127_3477_n393, DP_OP_425J2_127_3477_n392,
         DP_OP_425J2_127_3477_n391, DP_OP_425J2_127_3477_n390,
         DP_OP_425J2_127_3477_n389, DP_OP_425J2_127_3477_n388,
         DP_OP_425J2_127_3477_n387, DP_OP_425J2_127_3477_n386,
         DP_OP_425J2_127_3477_n385, DP_OP_425J2_127_3477_n384,
         DP_OP_425J2_127_3477_n383, DP_OP_425J2_127_3477_n382,
         DP_OP_425J2_127_3477_n381, DP_OP_425J2_127_3477_n380,
         DP_OP_425J2_127_3477_n379, DP_OP_425J2_127_3477_n378,
         DP_OP_425J2_127_3477_n377, DP_OP_425J2_127_3477_n376,
         DP_OP_425J2_127_3477_n375, DP_OP_425J2_127_3477_n374,
         DP_OP_425J2_127_3477_n373, DP_OP_425J2_127_3477_n372,
         DP_OP_425J2_127_3477_n371, DP_OP_425J2_127_3477_n370,
         DP_OP_425J2_127_3477_n369, DP_OP_425J2_127_3477_n368,
         DP_OP_425J2_127_3477_n367, DP_OP_425J2_127_3477_n366,
         DP_OP_425J2_127_3477_n365, DP_OP_425J2_127_3477_n364,
         DP_OP_425J2_127_3477_n363, DP_OP_425J2_127_3477_n362,
         DP_OP_425J2_127_3477_n361, DP_OP_425J2_127_3477_n360,
         DP_OP_425J2_127_3477_n359, DP_OP_425J2_127_3477_n358,
         DP_OP_425J2_127_3477_n357, DP_OP_425J2_127_3477_n356,
         DP_OP_425J2_127_3477_n355, DP_OP_425J2_127_3477_n354,
         DP_OP_425J2_127_3477_n353, DP_OP_425J2_127_3477_n352,
         DP_OP_425J2_127_3477_n351, DP_OP_425J2_127_3477_n350,
         DP_OP_425J2_127_3477_n349, DP_OP_425J2_127_3477_n348,
         DP_OP_425J2_127_3477_n347, DP_OP_425J2_127_3477_n346,
         DP_OP_425J2_127_3477_n345, DP_OP_425J2_127_3477_n344,
         DP_OP_425J2_127_3477_n343, DP_OP_425J2_127_3477_n342,
         DP_OP_425J2_127_3477_n341, DP_OP_425J2_127_3477_n340,
         DP_OP_425J2_127_3477_n339, DP_OP_425J2_127_3477_n338,
         DP_OP_425J2_127_3477_n337, DP_OP_425J2_127_3477_n336,
         DP_OP_425J2_127_3477_n335, DP_OP_425J2_127_3477_n334,
         DP_OP_425J2_127_3477_n333, DP_OP_425J2_127_3477_n332,
         DP_OP_425J2_127_3477_n331, DP_OP_425J2_127_3477_n330,
         DP_OP_425J2_127_3477_n329, DP_OP_425J2_127_3477_n328,
         DP_OP_425J2_127_3477_n327, DP_OP_425J2_127_3477_n326,
         DP_OP_425J2_127_3477_n325, DP_OP_425J2_127_3477_n324,
         DP_OP_425J2_127_3477_n323, DP_OP_425J2_127_3477_n322,
         DP_OP_425J2_127_3477_n321, DP_OP_425J2_127_3477_n320,
         DP_OP_425J2_127_3477_n319, DP_OP_425J2_127_3477_n318,
         DP_OP_425J2_127_3477_n317, DP_OP_425J2_127_3477_n316,
         DP_OP_425J2_127_3477_n315, DP_OP_425J2_127_3477_n314,
         DP_OP_425J2_127_3477_n313, DP_OP_425J2_127_3477_n312,
         DP_OP_425J2_127_3477_n311, DP_OP_425J2_127_3477_n310,
         DP_OP_425J2_127_3477_n309, DP_OP_425J2_127_3477_n308,
         DP_OP_425J2_127_3477_n307, DP_OP_425J2_127_3477_n306,
         DP_OP_425J2_127_3477_n305, DP_OP_425J2_127_3477_n304,
         DP_OP_425J2_127_3477_n303, DP_OP_425J2_127_3477_n302,
         DP_OP_425J2_127_3477_n301, DP_OP_425J2_127_3477_n300,
         DP_OP_425J2_127_3477_n299, DP_OP_425J2_127_3477_n298,
         DP_OP_425J2_127_3477_n297, DP_OP_425J2_127_3477_n296,
         DP_OP_425J2_127_3477_n295, DP_OP_425J2_127_3477_n294,
         DP_OP_425J2_127_3477_n293, DP_OP_425J2_127_3477_n292,
         DP_OP_425J2_127_3477_n291, DP_OP_425J2_127_3477_n290,
         DP_OP_425J2_127_3477_n289, DP_OP_425J2_127_3477_n288,
         DP_OP_425J2_127_3477_n287, DP_OP_425J2_127_3477_n286,
         DP_OP_425J2_127_3477_n285, DP_OP_425J2_127_3477_n284,
         DP_OP_425J2_127_3477_n283, DP_OP_425J2_127_3477_n282,
         DP_OP_425J2_127_3477_n281, DP_OP_425J2_127_3477_n280,
         DP_OP_425J2_127_3477_n279, DP_OP_425J2_127_3477_n278,
         DP_OP_425J2_127_3477_n277, DP_OP_425J2_127_3477_n276,
         DP_OP_425J2_127_3477_n275, DP_OP_425J2_127_3477_n274,
         DP_OP_425J2_127_3477_n273, DP_OP_425J2_127_3477_n272,
         DP_OP_425J2_127_3477_n271, DP_OP_425J2_127_3477_n270,
         DP_OP_425J2_127_3477_n269, DP_OP_425J2_127_3477_n268,
         DP_OP_425J2_127_3477_n267, DP_OP_425J2_127_3477_n266,
         DP_OP_425J2_127_3477_n265, DP_OP_425J2_127_3477_n264,
         DP_OP_425J2_127_3477_n263, DP_OP_425J2_127_3477_n262,
         DP_OP_425J2_127_3477_n261, DP_OP_425J2_127_3477_n260,
         DP_OP_425J2_127_3477_n259, DP_OP_425J2_127_3477_n258,
         DP_OP_425J2_127_3477_n257, DP_OP_425J2_127_3477_n256,
         DP_OP_425J2_127_3477_n255, DP_OP_425J2_127_3477_n254,
         DP_OP_425J2_127_3477_n253, DP_OP_425J2_127_3477_n252,
         DP_OP_425J2_127_3477_n251, DP_OP_425J2_127_3477_n250,
         DP_OP_425J2_127_3477_n249, DP_OP_425J2_127_3477_n248,
         DP_OP_425J2_127_3477_n247, DP_OP_425J2_127_3477_n246,
         DP_OP_425J2_127_3477_n245, DP_OP_425J2_127_3477_n244,
         DP_OP_425J2_127_3477_n243, DP_OP_425J2_127_3477_n242,
         DP_OP_425J2_127_3477_n241, DP_OP_425J2_127_3477_n240,
         DP_OP_425J2_127_3477_n239, DP_OP_425J2_127_3477_n238,
         DP_OP_425J2_127_3477_n237, DP_OP_425J2_127_3477_n236,
         DP_OP_425J2_127_3477_n235, DP_OP_425J2_127_3477_n234,
         DP_OP_425J2_127_3477_n233, DP_OP_425J2_127_3477_n232,
         DP_OP_425J2_127_3477_n231, DP_OP_425J2_127_3477_n230,
         DP_OP_425J2_127_3477_n229, DP_OP_425J2_127_3477_n228,
         DP_OP_425J2_127_3477_n227, DP_OP_425J2_127_3477_n226,
         DP_OP_425J2_127_3477_n225, DP_OP_425J2_127_3477_n224,
         DP_OP_425J2_127_3477_n223, DP_OP_425J2_127_3477_n222,
         DP_OP_425J2_127_3477_n221, DP_OP_425J2_127_3477_n220,
         DP_OP_425J2_127_3477_n219, DP_OP_425J2_127_3477_n218,
         DP_OP_425J2_127_3477_n217, DP_OP_425J2_127_3477_n216,
         DP_OP_425J2_127_3477_n215, DP_OP_425J2_127_3477_n214,
         DP_OP_425J2_127_3477_n213, DP_OP_425J2_127_3477_n212,
         DP_OP_425J2_127_3477_n211, DP_OP_425J2_127_3477_n210,
         DP_OP_425J2_127_3477_n209, DP_OP_425J2_127_3477_n208,
         DP_OP_425J2_127_3477_n207, DP_OP_425J2_127_3477_n206,
         DP_OP_425J2_127_3477_n205, DP_OP_425J2_127_3477_n204,
         DP_OP_425J2_127_3477_n203, DP_OP_425J2_127_3477_n202,
         DP_OP_425J2_127_3477_n201, DP_OP_425J2_127_3477_n200,
         DP_OP_425J2_127_3477_n199, DP_OP_425J2_127_3477_n198,
         DP_OP_425J2_127_3477_n197, DP_OP_425J2_127_3477_n196,
         DP_OP_425J2_127_3477_n195, DP_OP_425J2_127_3477_n194,
         DP_OP_425J2_127_3477_n193, DP_OP_425J2_127_3477_n192,
         DP_OP_425J2_127_3477_n191, DP_OP_425J2_127_3477_n190,
         DP_OP_425J2_127_3477_n189, DP_OP_425J2_127_3477_n188,
         DP_OP_425J2_127_3477_n187, DP_OP_425J2_127_3477_n186,
         DP_OP_425J2_127_3477_n185, DP_OP_425J2_127_3477_n184,
         DP_OP_425J2_127_3477_n183, DP_OP_425J2_127_3477_n182,
         DP_OP_425J2_127_3477_n181, DP_OP_425J2_127_3477_n180,
         DP_OP_425J2_127_3477_n179, DP_OP_425J2_127_3477_n178,
         DP_OP_425J2_127_3477_n177, DP_OP_425J2_127_3477_n176,
         DP_OP_425J2_127_3477_n175, DP_OP_425J2_127_3477_n174,
         DP_OP_425J2_127_3477_n173, DP_OP_425J2_127_3477_n172,
         DP_OP_425J2_127_3477_n171, DP_OP_425J2_127_3477_n170,
         DP_OP_425J2_127_3477_n169, DP_OP_425J2_127_3477_n168,
         DP_OP_425J2_127_3477_n167, DP_OP_425J2_127_3477_n166,
         DP_OP_425J2_127_3477_n165, DP_OP_425J2_127_3477_n164,
         DP_OP_425J2_127_3477_n163, DP_OP_425J2_127_3477_n162,
         DP_OP_425J2_127_3477_n161, DP_OP_425J2_127_3477_n160,
         DP_OP_425J2_127_3477_n159, DP_OP_425J2_127_3477_n158,
         DP_OP_425J2_127_3477_n157, DP_OP_425J2_127_3477_n156,
         DP_OP_425J2_127_3477_n155, DP_OP_425J2_127_3477_n154,
         DP_OP_425J2_127_3477_n153, DP_OP_425J2_127_3477_n131,
         DP_OP_425J2_127_3477_n130, DP_OP_425J2_127_3477_n129,
         DP_OP_425J2_127_3477_n128, DP_OP_425J2_127_3477_n127,
         DP_OP_425J2_127_3477_n126, DP_OP_425J2_127_3477_n123,
         DP_OP_425J2_127_3477_n122, DP_OP_425J2_127_3477_n121,
         DP_OP_425J2_127_3477_n120, DP_OP_425J2_127_3477_n119,
         DP_OP_425J2_127_3477_n118, DP_OP_425J2_127_3477_n115,
         DP_OP_425J2_127_3477_n114, DP_OP_425J2_127_3477_n113,
         DP_OP_425J2_127_3477_n112, DP_OP_425J2_127_3477_n111,
         DP_OP_425J2_127_3477_n110, DP_OP_425J2_127_3477_n107,
         DP_OP_425J2_127_3477_n106, DP_OP_425J2_127_3477_n105,
         DP_OP_425J2_127_3477_n104, DP_OP_425J2_127_3477_n103,
         DP_OP_425J2_127_3477_n102, DP_OP_425J2_127_3477_n101,
         DP_OP_425J2_127_3477_n99, DP_OP_425J2_127_3477_n98,
         DP_OP_425J2_127_3477_n95, DP_OP_425J2_127_3477_n94,
         DP_OP_425J2_127_3477_n93, DP_OP_425J2_127_3477_n92,
         DP_OP_425J2_127_3477_n90, DP_OP_425J2_127_3477_n88,
         DP_OP_425J2_127_3477_n87, DP_OP_425J2_127_3477_n86,
         DP_OP_425J2_127_3477_n85, DP_OP_425J2_127_3477_n84,
         DP_OP_425J2_127_3477_n83, DP_OP_425J2_127_3477_n82,
         DP_OP_425J2_127_3477_n80, DP_OP_425J2_127_3477_n79,
         DP_OP_425J2_127_3477_n78, DP_OP_425J2_127_3477_n77,
         DP_OP_425J2_127_3477_n76, DP_OP_425J2_127_3477_n75,
         DP_OP_425J2_127_3477_n74, DP_OP_425J2_127_3477_n73,
         DP_OP_425J2_127_3477_n69, DP_OP_425J2_127_3477_n68,
         DP_OP_425J2_127_3477_n67, DP_OP_425J2_127_3477_n66,
         DP_OP_425J2_127_3477_n65, DP_OP_425J2_127_3477_n64,
         DP_OP_425J2_127_3477_n62, DP_OP_425J2_127_3477_n60,
         DP_OP_425J2_127_3477_n59, DP_OP_425J2_127_3477_n57,
         DP_OP_425J2_127_3477_n56, DP_OP_425J2_127_3477_n55,
         DP_OP_425J2_127_3477_n53, DP_OP_425J2_127_3477_n52,
         DP_OP_425J2_127_3477_n51, DP_OP_425J2_127_3477_n50,
         DP_OP_425J2_127_3477_n46, DP_OP_425J2_127_3477_n45,
         DP_OP_425J2_127_3477_n42, DP_OP_425J2_127_3477_n41,
         DP_OP_425J2_127_3477_n39, DP_OP_425J2_127_3477_n38,
         DP_OP_425J2_127_3477_n37, DP_OP_425J2_127_3477_n36,
         DP_OP_425J2_127_3477_n35, DP_OP_425J2_127_3477_n34,
         DP_OP_425J2_127_3477_n33, DP_OP_425J2_127_3477_n32,
         DP_OP_425J2_127_3477_n31, DP_OP_425J2_127_3477_n30,
         DP_OP_425J2_127_3477_n29, DP_OP_425J2_127_3477_n28,
         DP_OP_425J2_127_3477_n27, DP_OP_425J2_127_3477_n26,
         DP_OP_425J2_127_3477_n25, DP_OP_425J2_127_3477_n24,
         DP_OP_425J2_127_3477_n4, DP_OP_425J2_127_3477_n3,
         DP_OP_425J2_127_3477_n2, DP_OP_424J2_126_3477_n2917,
         DP_OP_424J2_126_3477_n2915, DP_OP_424J2_126_3477_n2912,
         DP_OP_424J2_126_3477_n2910, DP_OP_424J2_126_3477_n2909,
         DP_OP_424J2_126_3477_n2906, DP_OP_424J2_126_3477_n2905,
         DP_OP_424J2_126_3477_n2904, DP_OP_424J2_126_3477_n2903,
         DP_OP_424J2_126_3477_n2902, DP_OP_424J2_126_3477_n2901,
         DP_OP_424J2_126_3477_n2900, DP_OP_424J2_126_3477_n2899,
         DP_OP_424J2_126_3477_n2898, DP_OP_424J2_126_3477_n2897,
         DP_OP_424J2_126_3477_n2896, DP_OP_424J2_126_3477_n2895,
         DP_OP_424J2_126_3477_n2894, DP_OP_424J2_126_3477_n2893,
         DP_OP_424J2_126_3477_n2892, DP_OP_424J2_126_3477_n2891,
         DP_OP_424J2_126_3477_n2890, DP_OP_424J2_126_3477_n2889,
         DP_OP_424J2_126_3477_n2888, DP_OP_424J2_126_3477_n2887,
         DP_OP_424J2_126_3477_n2886, DP_OP_424J2_126_3477_n2885,
         DP_OP_424J2_126_3477_n2884, DP_OP_424J2_126_3477_n2883,
         DP_OP_424J2_126_3477_n2882, DP_OP_424J2_126_3477_n2881,
         DP_OP_424J2_126_3477_n2880, DP_OP_424J2_126_3477_n2879,
         DP_OP_424J2_126_3477_n2878, DP_OP_424J2_126_3477_n2877,
         DP_OP_424J2_126_3477_n2876, DP_OP_424J2_126_3477_n2875,
         DP_OP_424J2_126_3477_n2874, DP_OP_424J2_126_3477_n2873,
         DP_OP_424J2_126_3477_n2869, DP_OP_424J2_126_3477_n2867,
         DP_OP_424J2_126_3477_n2865, DP_OP_424J2_126_3477_n2864,
         DP_OP_424J2_126_3477_n2863, DP_OP_424J2_126_3477_n2862,
         DP_OP_424J2_126_3477_n2861, DP_OP_424J2_126_3477_n2860,
         DP_OP_424J2_126_3477_n2859, DP_OP_424J2_126_3477_n2858,
         DP_OP_424J2_126_3477_n2857, DP_OP_424J2_126_3477_n2856,
         DP_OP_424J2_126_3477_n2855, DP_OP_424J2_126_3477_n2854,
         DP_OP_424J2_126_3477_n2853, DP_OP_424J2_126_3477_n2852,
         DP_OP_424J2_126_3477_n2851, DP_OP_424J2_126_3477_n2850,
         DP_OP_424J2_126_3477_n2849, DP_OP_424J2_126_3477_n2848,
         DP_OP_424J2_126_3477_n2847, DP_OP_424J2_126_3477_n2846,
         DP_OP_424J2_126_3477_n2845, DP_OP_424J2_126_3477_n2844,
         DP_OP_424J2_126_3477_n2843, DP_OP_424J2_126_3477_n2842,
         DP_OP_424J2_126_3477_n2841, DP_OP_424J2_126_3477_n2840,
         DP_OP_424J2_126_3477_n2839, DP_OP_424J2_126_3477_n2838,
         DP_OP_424J2_126_3477_n2837, DP_OP_424J2_126_3477_n2836,
         DP_OP_424J2_126_3477_n2835, DP_OP_424J2_126_3477_n2834,
         DP_OP_424J2_126_3477_n2833, DP_OP_424J2_126_3477_n2832,
         DP_OP_424J2_126_3477_n2831, DP_OP_424J2_126_3477_n2830,
         DP_OP_424J2_126_3477_n2829, DP_OP_424J2_126_3477_n2828,
         DP_OP_424J2_126_3477_n2827, DP_OP_424J2_126_3477_n2826,
         DP_OP_424J2_126_3477_n2825, DP_OP_424J2_126_3477_n2824,
         DP_OP_424J2_126_3477_n2823, DP_OP_424J2_126_3477_n2822,
         DP_OP_424J2_126_3477_n2821, DP_OP_424J2_126_3477_n2820,
         DP_OP_424J2_126_3477_n2819, DP_OP_424J2_126_3477_n2818,
         DP_OP_424J2_126_3477_n2817, DP_OP_424J2_126_3477_n2816,
         DP_OP_424J2_126_3477_n2815, DP_OP_424J2_126_3477_n2814,
         DP_OP_424J2_126_3477_n2813, DP_OP_424J2_126_3477_n2812,
         DP_OP_424J2_126_3477_n2811, DP_OP_424J2_126_3477_n2810,
         DP_OP_424J2_126_3477_n2809, DP_OP_424J2_126_3477_n2808,
         DP_OP_424J2_126_3477_n2807, DP_OP_424J2_126_3477_n2806,
         DP_OP_424J2_126_3477_n2805, DP_OP_424J2_126_3477_n2804,
         DP_OP_424J2_126_3477_n2803, DP_OP_424J2_126_3477_n2802,
         DP_OP_424J2_126_3477_n2801, DP_OP_424J2_126_3477_n2800,
         DP_OP_424J2_126_3477_n2799, DP_OP_424J2_126_3477_n2798,
         DP_OP_424J2_126_3477_n2797, DP_OP_424J2_126_3477_n2796,
         DP_OP_424J2_126_3477_n2795, DP_OP_424J2_126_3477_n2794,
         DP_OP_424J2_126_3477_n2793, DP_OP_424J2_126_3477_n2792,
         DP_OP_424J2_126_3477_n2791, DP_OP_424J2_126_3477_n2790,
         DP_OP_424J2_126_3477_n2789, DP_OP_424J2_126_3477_n2788,
         DP_OP_424J2_126_3477_n2787, DP_OP_424J2_126_3477_n2785,
         DP_OP_424J2_126_3477_n2784, DP_OP_424J2_126_3477_n2783,
         DP_OP_424J2_126_3477_n2777, DP_OP_424J2_126_3477_n2775,
         DP_OP_424J2_126_3477_n2774, DP_OP_424J2_126_3477_n2773,
         DP_OP_424J2_126_3477_n2772, DP_OP_424J2_126_3477_n2771,
         DP_OP_424J2_126_3477_n2770, DP_OP_424J2_126_3477_n2769,
         DP_OP_424J2_126_3477_n2768, DP_OP_424J2_126_3477_n2767,
         DP_OP_424J2_126_3477_n2766, DP_OP_424J2_126_3477_n2765,
         DP_OP_424J2_126_3477_n2764, DP_OP_424J2_126_3477_n2763,
         DP_OP_424J2_126_3477_n2762, DP_OP_424J2_126_3477_n2761,
         DP_OP_424J2_126_3477_n2760, DP_OP_424J2_126_3477_n2759,
         DP_OP_424J2_126_3477_n2758, DP_OP_424J2_126_3477_n2757,
         DP_OP_424J2_126_3477_n2756, DP_OP_424J2_126_3477_n2755,
         DP_OP_424J2_126_3477_n2754, DP_OP_424J2_126_3477_n2753,
         DP_OP_424J2_126_3477_n2752, DP_OP_424J2_126_3477_n2751,
         DP_OP_424J2_126_3477_n2750, DP_OP_424J2_126_3477_n2749,
         DP_OP_424J2_126_3477_n2748, DP_OP_424J2_126_3477_n2747,
         DP_OP_424J2_126_3477_n2746, DP_OP_424J2_126_3477_n2745,
         DP_OP_424J2_126_3477_n2744, DP_OP_424J2_126_3477_n2743,
         DP_OP_424J2_126_3477_n2742, DP_OP_424J2_126_3477_n2741,
         DP_OP_424J2_126_3477_n2740, DP_OP_424J2_126_3477_n2738,
         DP_OP_424J2_126_3477_n2737, DP_OP_424J2_126_3477_n2736,
         DP_OP_424J2_126_3477_n2735, DP_OP_424J2_126_3477_n2734,
         DP_OP_424J2_126_3477_n2733, DP_OP_424J2_126_3477_n2732,
         DP_OP_424J2_126_3477_n2731, DP_OP_424J2_126_3477_n2730,
         DP_OP_424J2_126_3477_n2729, DP_OP_424J2_126_3477_n2728,
         DP_OP_424J2_126_3477_n2727, DP_OP_424J2_126_3477_n2726,
         DP_OP_424J2_126_3477_n2725, DP_OP_424J2_126_3477_n2724,
         DP_OP_424J2_126_3477_n2723, DP_OP_424J2_126_3477_n2722,
         DP_OP_424J2_126_3477_n2721, DP_OP_424J2_126_3477_n2720,
         DP_OP_424J2_126_3477_n2719, DP_OP_424J2_126_3477_n2718,
         DP_OP_424J2_126_3477_n2717, DP_OP_424J2_126_3477_n2716,
         DP_OP_424J2_126_3477_n2715, DP_OP_424J2_126_3477_n2714,
         DP_OP_424J2_126_3477_n2713, DP_OP_424J2_126_3477_n2712,
         DP_OP_424J2_126_3477_n2711, DP_OP_424J2_126_3477_n2710,
         DP_OP_424J2_126_3477_n2709, DP_OP_424J2_126_3477_n2708,
         DP_OP_424J2_126_3477_n2707, DP_OP_424J2_126_3477_n2706,
         DP_OP_424J2_126_3477_n2705, DP_OP_424J2_126_3477_n2704,
         DP_OP_424J2_126_3477_n2703, DP_OP_424J2_126_3477_n2702,
         DP_OP_424J2_126_3477_n2701, DP_OP_424J2_126_3477_n2700,
         DP_OP_424J2_126_3477_n2699, DP_OP_424J2_126_3477_n2698,
         DP_OP_424J2_126_3477_n2697, DP_OP_424J2_126_3477_n2696,
         DP_OP_424J2_126_3477_n2695, DP_OP_424J2_126_3477_n2693,
         DP_OP_424J2_126_3477_n2691, DP_OP_424J2_126_3477_n2689,
         DP_OP_424J2_126_3477_n2686, DP_OP_424J2_126_3477_n2685,
         DP_OP_424J2_126_3477_n2684, DP_OP_424J2_126_3477_n2683,
         DP_OP_424J2_126_3477_n2682, DP_OP_424J2_126_3477_n2681,
         DP_OP_424J2_126_3477_n2680, DP_OP_424J2_126_3477_n2679,
         DP_OP_424J2_126_3477_n2678, DP_OP_424J2_126_3477_n2677,
         DP_OP_424J2_126_3477_n2676, DP_OP_424J2_126_3477_n2675,
         DP_OP_424J2_126_3477_n2674, DP_OP_424J2_126_3477_n2673,
         DP_OP_424J2_126_3477_n2672, DP_OP_424J2_126_3477_n2671,
         DP_OP_424J2_126_3477_n2670, DP_OP_424J2_126_3477_n2669,
         DP_OP_424J2_126_3477_n2668, DP_OP_424J2_126_3477_n2667,
         DP_OP_424J2_126_3477_n2666, DP_OP_424J2_126_3477_n2665,
         DP_OP_424J2_126_3477_n2664, DP_OP_424J2_126_3477_n2663,
         DP_OP_424J2_126_3477_n2662, DP_OP_424J2_126_3477_n2661,
         DP_OP_424J2_126_3477_n2660, DP_OP_424J2_126_3477_n2659,
         DP_OP_424J2_126_3477_n2658, DP_OP_424J2_126_3477_n2657,
         DP_OP_424J2_126_3477_n2656, DP_OP_424J2_126_3477_n2655,
         DP_OP_424J2_126_3477_n2654, DP_OP_424J2_126_3477_n2653,
         DP_OP_424J2_126_3477_n2652, DP_OP_424J2_126_3477_n2651,
         DP_OP_424J2_126_3477_n2650, DP_OP_424J2_126_3477_n2649,
         DP_OP_424J2_126_3477_n2644, DP_OP_424J2_126_3477_n2642,
         DP_OP_424J2_126_3477_n2641, DP_OP_424J2_126_3477_n2640,
         DP_OP_424J2_126_3477_n2639, DP_OP_424J2_126_3477_n2638,
         DP_OP_424J2_126_3477_n2637, DP_OP_424J2_126_3477_n2636,
         DP_OP_424J2_126_3477_n2635, DP_OP_424J2_126_3477_n2634,
         DP_OP_424J2_126_3477_n2633, DP_OP_424J2_126_3477_n2632,
         DP_OP_424J2_126_3477_n2631, DP_OP_424J2_126_3477_n2630,
         DP_OP_424J2_126_3477_n2629, DP_OP_424J2_126_3477_n2628,
         DP_OP_424J2_126_3477_n2627, DP_OP_424J2_126_3477_n2626,
         DP_OP_424J2_126_3477_n2625, DP_OP_424J2_126_3477_n2624,
         DP_OP_424J2_126_3477_n2623, DP_OP_424J2_126_3477_n2622,
         DP_OP_424J2_126_3477_n2621, DP_OP_424J2_126_3477_n2620,
         DP_OP_424J2_126_3477_n2619, DP_OP_424J2_126_3477_n2618,
         DP_OP_424J2_126_3477_n2617, DP_OP_424J2_126_3477_n2616,
         DP_OP_424J2_126_3477_n2615, DP_OP_424J2_126_3477_n2614,
         DP_OP_424J2_126_3477_n2613, DP_OP_424J2_126_3477_n2612,
         DP_OP_424J2_126_3477_n2611, DP_OP_424J2_126_3477_n2610,
         DP_OP_424J2_126_3477_n2609, DP_OP_424J2_126_3477_n2608,
         DP_OP_424J2_126_3477_n2607, DP_OP_424J2_126_3477_n2604,
         DP_OP_424J2_126_3477_n2600, DP_OP_424J2_126_3477_n2598,
         DP_OP_424J2_126_3477_n2597, DP_OP_424J2_126_3477_n2596,
         DP_OP_424J2_126_3477_n2595, DP_OP_424J2_126_3477_n2594,
         DP_OP_424J2_126_3477_n2593, DP_OP_424J2_126_3477_n2592,
         DP_OP_424J2_126_3477_n2591, DP_OP_424J2_126_3477_n2590,
         DP_OP_424J2_126_3477_n2589, DP_OP_424J2_126_3477_n2588,
         DP_OP_424J2_126_3477_n2587, DP_OP_424J2_126_3477_n2586,
         DP_OP_424J2_126_3477_n2585, DP_OP_424J2_126_3477_n2584,
         DP_OP_424J2_126_3477_n2583, DP_OP_424J2_126_3477_n2582,
         DP_OP_424J2_126_3477_n2581, DP_OP_424J2_126_3477_n2580,
         DP_OP_424J2_126_3477_n2579, DP_OP_424J2_126_3477_n2578,
         DP_OP_424J2_126_3477_n2577, DP_OP_424J2_126_3477_n2576,
         DP_OP_424J2_126_3477_n2575, DP_OP_424J2_126_3477_n2574,
         DP_OP_424J2_126_3477_n2573, DP_OP_424J2_126_3477_n2572,
         DP_OP_424J2_126_3477_n2571, DP_OP_424J2_126_3477_n2570,
         DP_OP_424J2_126_3477_n2569, DP_OP_424J2_126_3477_n2568,
         DP_OP_424J2_126_3477_n2567, DP_OP_424J2_126_3477_n2566,
         DP_OP_424J2_126_3477_n2565, DP_OP_424J2_126_3477_n2563,
         DP_OP_424J2_126_3477_n2561, DP_OP_424J2_126_3477_n2559,
         DP_OP_424J2_126_3477_n2557, DP_OP_424J2_126_3477_n2555,
         DP_OP_424J2_126_3477_n2554, DP_OP_424J2_126_3477_n2553,
         DP_OP_424J2_126_3477_n2552, DP_OP_424J2_126_3477_n2551,
         DP_OP_424J2_126_3477_n2550, DP_OP_424J2_126_3477_n2549,
         DP_OP_424J2_126_3477_n2548, DP_OP_424J2_126_3477_n2547,
         DP_OP_424J2_126_3477_n2546, DP_OP_424J2_126_3477_n2545,
         DP_OP_424J2_126_3477_n2544, DP_OP_424J2_126_3477_n2543,
         DP_OP_424J2_126_3477_n2542, DP_OP_424J2_126_3477_n2541,
         DP_OP_424J2_126_3477_n2540, DP_OP_424J2_126_3477_n2539,
         DP_OP_424J2_126_3477_n2538, DP_OP_424J2_126_3477_n2537,
         DP_OP_424J2_126_3477_n2536, DP_OP_424J2_126_3477_n2535,
         DP_OP_424J2_126_3477_n2534, DP_OP_424J2_126_3477_n2533,
         DP_OP_424J2_126_3477_n2532, DP_OP_424J2_126_3477_n2531,
         DP_OP_424J2_126_3477_n2530, DP_OP_424J2_126_3477_n2529,
         DP_OP_424J2_126_3477_n2528, DP_OP_424J2_126_3477_n2527,
         DP_OP_424J2_126_3477_n2526, DP_OP_424J2_126_3477_n2525,
         DP_OP_424J2_126_3477_n2524, DP_OP_424J2_126_3477_n2523,
         DP_OP_424J2_126_3477_n2522, DP_OP_424J2_126_3477_n2521,
         DP_OP_424J2_126_3477_n2520, DP_OP_424J2_126_3477_n2517,
         DP_OP_424J2_126_3477_n2512, DP_OP_424J2_126_3477_n2510,
         DP_OP_424J2_126_3477_n2509, DP_OP_424J2_126_3477_n2508,
         DP_OP_424J2_126_3477_n2507, DP_OP_424J2_126_3477_n2506,
         DP_OP_424J2_126_3477_n2505, DP_OP_424J2_126_3477_n2504,
         DP_OP_424J2_126_3477_n2503, DP_OP_424J2_126_3477_n2502,
         DP_OP_424J2_126_3477_n2501, DP_OP_424J2_126_3477_n2500,
         DP_OP_424J2_126_3477_n2499, DP_OP_424J2_126_3477_n2498,
         DP_OP_424J2_126_3477_n2497, DP_OP_424J2_126_3477_n2496,
         DP_OP_424J2_126_3477_n2495, DP_OP_424J2_126_3477_n2494,
         DP_OP_424J2_126_3477_n2493, DP_OP_424J2_126_3477_n2492,
         DP_OP_424J2_126_3477_n2491, DP_OP_424J2_126_3477_n2490,
         DP_OP_424J2_126_3477_n2489, DP_OP_424J2_126_3477_n2488,
         DP_OP_424J2_126_3477_n2487, DP_OP_424J2_126_3477_n2486,
         DP_OP_424J2_126_3477_n2485, DP_OP_424J2_126_3477_n2484,
         DP_OP_424J2_126_3477_n2483, DP_OP_424J2_126_3477_n2482,
         DP_OP_424J2_126_3477_n2481, DP_OP_424J2_126_3477_n2480,
         DP_OP_424J2_126_3477_n2479, DP_OP_424J2_126_3477_n2478,
         DP_OP_424J2_126_3477_n2475, DP_OP_424J2_126_3477_n2474,
         DP_OP_424J2_126_3477_n2472, DP_OP_424J2_126_3477_n2471,
         DP_OP_424J2_126_3477_n2466, DP_OP_424J2_126_3477_n2465,
         DP_OP_424J2_126_3477_n2464, DP_OP_424J2_126_3477_n2463,
         DP_OP_424J2_126_3477_n2462, DP_OP_424J2_126_3477_n2461,
         DP_OP_424J2_126_3477_n2460, DP_OP_424J2_126_3477_n2459,
         DP_OP_424J2_126_3477_n2458, DP_OP_424J2_126_3477_n2457,
         DP_OP_424J2_126_3477_n2456, DP_OP_424J2_126_3477_n2455,
         DP_OP_424J2_126_3477_n2454, DP_OP_424J2_126_3477_n2453,
         DP_OP_424J2_126_3477_n2452, DP_OP_424J2_126_3477_n2451,
         DP_OP_424J2_126_3477_n2450, DP_OP_424J2_126_3477_n2449,
         DP_OP_424J2_126_3477_n2448, DP_OP_424J2_126_3477_n2447,
         DP_OP_424J2_126_3477_n2446, DP_OP_424J2_126_3477_n2445,
         DP_OP_424J2_126_3477_n2444, DP_OP_424J2_126_3477_n2443,
         DP_OP_424J2_126_3477_n2442, DP_OP_424J2_126_3477_n2441,
         DP_OP_424J2_126_3477_n2440, DP_OP_424J2_126_3477_n2439,
         DP_OP_424J2_126_3477_n2438, DP_OP_424J2_126_3477_n2437,
         DP_OP_424J2_126_3477_n2436, DP_OP_424J2_126_3477_n2435,
         DP_OP_424J2_126_3477_n2432, DP_OP_424J2_126_3477_n2430,
         DP_OP_424J2_126_3477_n2428, DP_OP_424J2_126_3477_n2423,
         DP_OP_424J2_126_3477_n2422, DP_OP_424J2_126_3477_n2421,
         DP_OP_424J2_126_3477_n2420, DP_OP_424J2_126_3477_n2419,
         DP_OP_424J2_126_3477_n2418, DP_OP_424J2_126_3477_n2417,
         DP_OP_424J2_126_3477_n2416, DP_OP_424J2_126_3477_n2415,
         DP_OP_424J2_126_3477_n2414, DP_OP_424J2_126_3477_n2413,
         DP_OP_424J2_126_3477_n2412, DP_OP_424J2_126_3477_n2411,
         DP_OP_424J2_126_3477_n2410, DP_OP_424J2_126_3477_n2409,
         DP_OP_424J2_126_3477_n2408, DP_OP_424J2_126_3477_n2407,
         DP_OP_424J2_126_3477_n2406, DP_OP_424J2_126_3477_n2405,
         DP_OP_424J2_126_3477_n2404, DP_OP_424J2_126_3477_n2403,
         DP_OP_424J2_126_3477_n2402, DP_OP_424J2_126_3477_n2401,
         DP_OP_424J2_126_3477_n2400, DP_OP_424J2_126_3477_n2399,
         DP_OP_424J2_126_3477_n2398, DP_OP_424J2_126_3477_n2397,
         DP_OP_424J2_126_3477_n2396, DP_OP_424J2_126_3477_n2395,
         DP_OP_424J2_126_3477_n2394, DP_OP_424J2_126_3477_n2393,
         DP_OP_424J2_126_3477_n2392, DP_OP_424J2_126_3477_n2391,
         DP_OP_424J2_126_3477_n2390, DP_OP_424J2_126_3477_n2389,
         DP_OP_424J2_126_3477_n2388, DP_OP_424J2_126_3477_n2387,
         DP_OP_424J2_126_3477_n2386, DP_OP_424J2_126_3477_n2385,
         DP_OP_424J2_126_3477_n2384, DP_OP_424J2_126_3477_n2383,
         DP_OP_424J2_126_3477_n2382, DP_OP_424J2_126_3477_n2381,
         DP_OP_424J2_126_3477_n2378, DP_OP_424J2_126_3477_n2377,
         DP_OP_424J2_126_3477_n2376, DP_OP_424J2_126_3477_n2375,
         DP_OP_424J2_126_3477_n2374, DP_OP_424J2_126_3477_n2373,
         DP_OP_424J2_126_3477_n2372, DP_OP_424J2_126_3477_n2371,
         DP_OP_424J2_126_3477_n2370, DP_OP_424J2_126_3477_n2369,
         DP_OP_424J2_126_3477_n2368, DP_OP_424J2_126_3477_n2367,
         DP_OP_424J2_126_3477_n2366, DP_OP_424J2_126_3477_n2365,
         DP_OP_424J2_126_3477_n2364, DP_OP_424J2_126_3477_n2363,
         DP_OP_424J2_126_3477_n2362, DP_OP_424J2_126_3477_n2361,
         DP_OP_424J2_126_3477_n2360, DP_OP_424J2_126_3477_n2359,
         DP_OP_424J2_126_3477_n2358, DP_OP_424J2_126_3477_n2357,
         DP_OP_424J2_126_3477_n2356, DP_OP_424J2_126_3477_n2355,
         DP_OP_424J2_126_3477_n2354, DP_OP_424J2_126_3477_n2353,
         DP_OP_424J2_126_3477_n2352, DP_OP_424J2_126_3477_n2351,
         DP_OP_424J2_126_3477_n2350, DP_OP_424J2_126_3477_n2349,
         DP_OP_424J2_126_3477_n2344, DP_OP_424J2_126_3477_n2342,
         DP_OP_424J2_126_3477_n2341, DP_OP_424J2_126_3477_n2339,
         DP_OP_424J2_126_3477_n2338, DP_OP_424J2_126_3477_n2337,
         DP_OP_424J2_126_3477_n2336, DP_OP_424J2_126_3477_n2335,
         DP_OP_424J2_126_3477_n2334, DP_OP_424J2_126_3477_n2333,
         DP_OP_424J2_126_3477_n2332, DP_OP_424J2_126_3477_n2331,
         DP_OP_424J2_126_3477_n2330, DP_OP_424J2_126_3477_n2329,
         DP_OP_424J2_126_3477_n2328, DP_OP_424J2_126_3477_n2327,
         DP_OP_424J2_126_3477_n2326, DP_OP_424J2_126_3477_n2325,
         DP_OP_424J2_126_3477_n2324, DP_OP_424J2_126_3477_n2323,
         DP_OP_424J2_126_3477_n2322, DP_OP_424J2_126_3477_n2321,
         DP_OP_424J2_126_3477_n2320, DP_OP_424J2_126_3477_n2319,
         DP_OP_424J2_126_3477_n2318, DP_OP_424J2_126_3477_n2317,
         DP_OP_424J2_126_3477_n2316, DP_OP_424J2_126_3477_n2315,
         DP_OP_424J2_126_3477_n2314, DP_OP_424J2_126_3477_n2313,
         DP_OP_424J2_126_3477_n2312, DP_OP_424J2_126_3477_n2311,
         DP_OP_424J2_126_3477_n2310, DP_OP_424J2_126_3477_n2309,
         DP_OP_424J2_126_3477_n2308, DP_OP_424J2_126_3477_n2307,
         DP_OP_424J2_126_3477_n2306, DP_OP_424J2_126_3477_n2304,
         DP_OP_424J2_126_3477_n2302, DP_OP_424J2_126_3477_n2296,
         DP_OP_424J2_126_3477_n2293, DP_OP_424J2_126_3477_n2292,
         DP_OP_424J2_126_3477_n2291, DP_OP_424J2_126_3477_n2290,
         DP_OP_424J2_126_3477_n2289, DP_OP_424J2_126_3477_n2288,
         DP_OP_424J2_126_3477_n2287, DP_OP_424J2_126_3477_n2286,
         DP_OP_424J2_126_3477_n2285, DP_OP_424J2_126_3477_n2284,
         DP_OP_424J2_126_3477_n2283, DP_OP_424J2_126_3477_n2282,
         DP_OP_424J2_126_3477_n2281, DP_OP_424J2_126_3477_n2280,
         DP_OP_424J2_126_3477_n2279, DP_OP_424J2_126_3477_n2278,
         DP_OP_424J2_126_3477_n2277, DP_OP_424J2_126_3477_n2276,
         DP_OP_424J2_126_3477_n2275, DP_OP_424J2_126_3477_n2274,
         DP_OP_424J2_126_3477_n2273, DP_OP_424J2_126_3477_n2272,
         DP_OP_424J2_126_3477_n2271, DP_OP_424J2_126_3477_n2270,
         DP_OP_424J2_126_3477_n2269, DP_OP_424J2_126_3477_n2268,
         DP_OP_424J2_126_3477_n2267, DP_OP_424J2_126_3477_n2266,
         DP_OP_424J2_126_3477_n2265, DP_OP_424J2_126_3477_n2264,
         DP_OP_424J2_126_3477_n2263, DP_OP_424J2_126_3477_n2262,
         DP_OP_424J2_126_3477_n2260, DP_OP_424J2_126_3477_n2258,
         DP_OP_424J2_126_3477_n2249, DP_OP_424J2_126_3477_n2248,
         DP_OP_424J2_126_3477_n2247, DP_OP_424J2_126_3477_n2246,
         DP_OP_424J2_126_3477_n2245, DP_OP_424J2_126_3477_n2244,
         DP_OP_424J2_126_3477_n2243, DP_OP_424J2_126_3477_n2242,
         DP_OP_424J2_126_3477_n2241, DP_OP_424J2_126_3477_n2240,
         DP_OP_424J2_126_3477_n2239, DP_OP_424J2_126_3477_n2238,
         DP_OP_424J2_126_3477_n2237, DP_OP_424J2_126_3477_n2236,
         DP_OP_424J2_126_3477_n2235, DP_OP_424J2_126_3477_n2234,
         DP_OP_424J2_126_3477_n2233, DP_OP_424J2_126_3477_n2232,
         DP_OP_424J2_126_3477_n2231, DP_OP_424J2_126_3477_n2230,
         DP_OP_424J2_126_3477_n2229, DP_OP_424J2_126_3477_n2228,
         DP_OP_424J2_126_3477_n2227, DP_OP_424J2_126_3477_n2226,
         DP_OP_424J2_126_3477_n2225, DP_OP_424J2_126_3477_n2224,
         DP_OP_424J2_126_3477_n2223, DP_OP_424J2_126_3477_n2222,
         DP_OP_424J2_126_3477_n2221, DP_OP_424J2_126_3477_n2220,
         DP_OP_424J2_126_3477_n2219, DP_OP_424J2_126_3477_n2218,
         DP_OP_424J2_126_3477_n2216, DP_OP_424J2_126_3477_n2212,
         DP_OP_424J2_126_3477_n2211, DP_OP_424J2_126_3477_n2205,
         DP_OP_424J2_126_3477_n2204, DP_OP_424J2_126_3477_n2203,
         DP_OP_424J2_126_3477_n2202, DP_OP_424J2_126_3477_n2201,
         DP_OP_424J2_126_3477_n2200, DP_OP_424J2_126_3477_n2199,
         DP_OP_424J2_126_3477_n2198, DP_OP_424J2_126_3477_n2197,
         DP_OP_424J2_126_3477_n2196, DP_OP_424J2_126_3477_n2195,
         DP_OP_424J2_126_3477_n2194, DP_OP_424J2_126_3477_n2193,
         DP_OP_424J2_126_3477_n2192, DP_OP_424J2_126_3477_n2191,
         DP_OP_424J2_126_3477_n2190, DP_OP_424J2_126_3477_n2189,
         DP_OP_424J2_126_3477_n2188, DP_OP_424J2_126_3477_n2187,
         DP_OP_424J2_126_3477_n2186, DP_OP_424J2_126_3477_n2185,
         DP_OP_424J2_126_3477_n2184, DP_OP_424J2_126_3477_n2183,
         DP_OP_424J2_126_3477_n2182, DP_OP_424J2_126_3477_n2181,
         DP_OP_424J2_126_3477_n2180, DP_OP_424J2_126_3477_n2179,
         DP_OP_424J2_126_3477_n2178, DP_OP_424J2_126_3477_n2177,
         DP_OP_424J2_126_3477_n2176, DP_OP_424J2_126_3477_n2175,
         DP_OP_424J2_126_3477_n2174, DP_OP_424J2_126_3477_n2173,
         DP_OP_424J2_126_3477_n2171, DP_OP_424J2_126_3477_n2170,
         DP_OP_424J2_126_3477_n2168, DP_OP_424J2_126_3477_n2164,
         DP_OP_424J2_126_3477_n2163, DP_OP_424J2_126_3477_n2161,
         DP_OP_424J2_126_3477_n2160, DP_OP_424J2_126_3477_n2159,
         DP_OP_424J2_126_3477_n2158, DP_OP_424J2_126_3477_n2157,
         DP_OP_424J2_126_3477_n2156, DP_OP_424J2_126_3477_n2155,
         DP_OP_424J2_126_3477_n2154, DP_OP_424J2_126_3477_n2153,
         DP_OP_424J2_126_3477_n2152, DP_OP_424J2_126_3477_n2151,
         DP_OP_424J2_126_3477_n2150, DP_OP_424J2_126_3477_n2149,
         DP_OP_424J2_126_3477_n2148, DP_OP_424J2_126_3477_n2147,
         DP_OP_424J2_126_3477_n2146, DP_OP_424J2_126_3477_n2145,
         DP_OP_424J2_126_3477_n2144, DP_OP_424J2_126_3477_n2143,
         DP_OP_424J2_126_3477_n2142, DP_OP_424J2_126_3477_n2141,
         DP_OP_424J2_126_3477_n2140, DP_OP_424J2_126_3477_n2139,
         DP_OP_424J2_126_3477_n2138, DP_OP_424J2_126_3477_n2137,
         DP_OP_424J2_126_3477_n2136, DP_OP_424J2_126_3477_n2135,
         DP_OP_424J2_126_3477_n2134, DP_OP_424J2_126_3477_n2133,
         DP_OP_424J2_126_3477_n2132, DP_OP_424J2_126_3477_n2131,
         DP_OP_424J2_126_3477_n2130, DP_OP_424J2_126_3477_n2129,
         DP_OP_424J2_126_3477_n2127, DP_OP_424J2_126_3477_n2126,
         DP_OP_424J2_126_3477_n2125, DP_OP_424J2_126_3477_n2124,
         DP_OP_424J2_126_3477_n2120, DP_OP_424J2_126_3477_n2119,
         DP_OP_424J2_126_3477_n2118, DP_OP_424J2_126_3477_n2117,
         DP_OP_424J2_126_3477_n2116, DP_OP_424J2_126_3477_n2115,
         DP_OP_424J2_126_3477_n2114, DP_OP_424J2_126_3477_n2113,
         DP_OP_424J2_126_3477_n2112, DP_OP_424J2_126_3477_n2111,
         DP_OP_424J2_126_3477_n2110, DP_OP_424J2_126_3477_n2109,
         DP_OP_424J2_126_3477_n2108, DP_OP_424J2_126_3477_n2107,
         DP_OP_424J2_126_3477_n2106, DP_OP_424J2_126_3477_n2105,
         DP_OP_424J2_126_3477_n2104, DP_OP_424J2_126_3477_n2103,
         DP_OP_424J2_126_3477_n2102, DP_OP_424J2_126_3477_n2101,
         DP_OP_424J2_126_3477_n2100, DP_OP_424J2_126_3477_n2099,
         DP_OP_424J2_126_3477_n2098, DP_OP_424J2_126_3477_n2097,
         DP_OP_424J2_126_3477_n2096, DP_OP_424J2_126_3477_n2095,
         DP_OP_424J2_126_3477_n2094, DP_OP_424J2_126_3477_n2093,
         DP_OP_424J2_126_3477_n2092, DP_OP_424J2_126_3477_n2091,
         DP_OP_424J2_126_3477_n2090, DP_OP_424J2_126_3477_n2089,
         DP_OP_424J2_126_3477_n2088, DP_OP_424J2_126_3477_n2087,
         DP_OP_424J2_126_3477_n2086, DP_OP_424J2_126_3477_n2085,
         DP_OP_424J2_126_3477_n2084, DP_OP_424J2_126_3477_n2082,
         DP_OP_424J2_126_3477_n2078, DP_OP_424J2_126_3477_n2077,
         DP_OP_424J2_126_3477_n2074, DP_OP_424J2_126_3477_n2073,
         DP_OP_424J2_126_3477_n2072, DP_OP_424J2_126_3477_n2071,
         DP_OP_424J2_126_3477_n2070, DP_OP_424J2_126_3477_n2069,
         DP_OP_424J2_126_3477_n2068, DP_OP_424J2_126_3477_n2067,
         DP_OP_424J2_126_3477_n2066, DP_OP_424J2_126_3477_n2065,
         DP_OP_424J2_126_3477_n2064, DP_OP_424J2_126_3477_n2063,
         DP_OP_424J2_126_3477_n2062, DP_OP_424J2_126_3477_n2061,
         DP_OP_424J2_126_3477_n2060, DP_OP_424J2_126_3477_n2059,
         DP_OP_424J2_126_3477_n2058, DP_OP_424J2_126_3477_n2057,
         DP_OP_424J2_126_3477_n2056, DP_OP_424J2_126_3477_n2055,
         DP_OP_424J2_126_3477_n2054, DP_OP_424J2_126_3477_n2053,
         DP_OP_424J2_126_3477_n2052, DP_OP_424J2_126_3477_n2051,
         DP_OP_424J2_126_3477_n2050, DP_OP_424J2_126_3477_n2049,
         DP_OP_424J2_126_3477_n2048, DP_OP_424J2_126_3477_n2047,
         DP_OP_424J2_126_3477_n2046, DP_OP_424J2_126_3477_n2045,
         DP_OP_424J2_126_3477_n2044, DP_OP_424J2_126_3477_n2043,
         DP_OP_424J2_126_3477_n2042, DP_OP_424J2_126_3477_n2041,
         DP_OP_424J2_126_3477_n2040, DP_OP_424J2_126_3477_n2039,
         DP_OP_424J2_126_3477_n2038, DP_OP_424J2_126_3477_n2037,
         DP_OP_424J2_126_3477_n2035, DP_OP_424J2_126_3477_n2034,
         DP_OP_424J2_126_3477_n2033, DP_OP_424J2_126_3477_n2032,
         DP_OP_424J2_126_3477_n2029, DP_OP_424J2_126_3477_n2028,
         DP_OP_424J2_126_3477_n2027, DP_OP_424J2_126_3477_n2026,
         DP_OP_424J2_126_3477_n2025, DP_OP_424J2_126_3477_n2024,
         DP_OP_424J2_126_3477_n2023, DP_OP_424J2_126_3477_n2022,
         DP_OP_424J2_126_3477_n2021, DP_OP_424J2_126_3477_n2020,
         DP_OP_424J2_126_3477_n2019, DP_OP_424J2_126_3477_n2018,
         DP_OP_424J2_126_3477_n2017, DP_OP_424J2_126_3477_n2016,
         DP_OP_424J2_126_3477_n2015, DP_OP_424J2_126_3477_n2014,
         DP_OP_424J2_126_3477_n2013, DP_OP_424J2_126_3477_n2012,
         DP_OP_424J2_126_3477_n2011, DP_OP_424J2_126_3477_n2010,
         DP_OP_424J2_126_3477_n2009, DP_OP_424J2_126_3477_n2008,
         DP_OP_424J2_126_3477_n2007, DP_OP_424J2_126_3477_n2006,
         DP_OP_424J2_126_3477_n2005, DP_OP_424J2_126_3477_n2004,
         DP_OP_424J2_126_3477_n2003, DP_OP_424J2_126_3477_n2002,
         DP_OP_424J2_126_3477_n2001, DP_OP_424J2_126_3477_n2000,
         DP_OP_424J2_126_3477_n1999, DP_OP_424J2_126_3477_n1998,
         DP_OP_424J2_126_3477_n1996, DP_OP_424J2_126_3477_n1995,
         DP_OP_424J2_126_3477_n1994, DP_OP_424J2_126_3477_n1988,
         DP_OP_424J2_126_3477_n1986, DP_OP_424J2_126_3477_n1985,
         DP_OP_424J2_126_3477_n1984, DP_OP_424J2_126_3477_n1983,
         DP_OP_424J2_126_3477_n1982, DP_OP_424J2_126_3477_n1981,
         DP_OP_424J2_126_3477_n1980, DP_OP_424J2_126_3477_n1979,
         DP_OP_424J2_126_3477_n1978, DP_OP_424J2_126_3477_n1977,
         DP_OP_424J2_126_3477_n1976, DP_OP_424J2_126_3477_n1975,
         DP_OP_424J2_126_3477_n1974, DP_OP_424J2_126_3477_n1973,
         DP_OP_424J2_126_3477_n1972, DP_OP_424J2_126_3477_n1971,
         DP_OP_424J2_126_3477_n1970, DP_OP_424J2_126_3477_n1969,
         DP_OP_424J2_126_3477_n1968, DP_OP_424J2_126_3477_n1967,
         DP_OP_424J2_126_3477_n1966, DP_OP_424J2_126_3477_n1965,
         DP_OP_424J2_126_3477_n1964, DP_OP_424J2_126_3477_n1963,
         DP_OP_424J2_126_3477_n1962, DP_OP_424J2_126_3477_n1961,
         DP_OP_424J2_126_3477_n1960, DP_OP_424J2_126_3477_n1959,
         DP_OP_424J2_126_3477_n1958, DP_OP_424J2_126_3477_n1957,
         DP_OP_424J2_126_3477_n1956, DP_OP_424J2_126_3477_n1955,
         DP_OP_424J2_126_3477_n1954, DP_OP_424J2_126_3477_n1953,
         DP_OP_424J2_126_3477_n1952, DP_OP_424J2_126_3477_n1950,
         DP_OP_424J2_126_3477_n1949, DP_OP_424J2_126_3477_n1948,
         DP_OP_424J2_126_3477_n1942, DP_OP_424J2_126_3477_n1941,
         DP_OP_424J2_126_3477_n1940, DP_OP_424J2_126_3477_n1939,
         DP_OP_424J2_126_3477_n1938, DP_OP_424J2_126_3477_n1937,
         DP_OP_424J2_126_3477_n1936, DP_OP_424J2_126_3477_n1935,
         DP_OP_424J2_126_3477_n1934, DP_OP_424J2_126_3477_n1933,
         DP_OP_424J2_126_3477_n1932, DP_OP_424J2_126_3477_n1931,
         DP_OP_424J2_126_3477_n1930, DP_OP_424J2_126_3477_n1929,
         DP_OP_424J2_126_3477_n1928, DP_OP_424J2_126_3477_n1927,
         DP_OP_424J2_126_3477_n1926, DP_OP_424J2_126_3477_n1925,
         DP_OP_424J2_126_3477_n1924, DP_OP_424J2_126_3477_n1923,
         DP_OP_424J2_126_3477_n1922, DP_OP_424J2_126_3477_n1921,
         DP_OP_424J2_126_3477_n1920, DP_OP_424J2_126_3477_n1919,
         DP_OP_424J2_126_3477_n1918, DP_OP_424J2_126_3477_n1917,
         DP_OP_424J2_126_3477_n1916, DP_OP_424J2_126_3477_n1915,
         DP_OP_424J2_126_3477_n1914, DP_OP_424J2_126_3477_n1913,
         DP_OP_424J2_126_3477_n1912, DP_OP_424J2_126_3477_n1911,
         DP_OP_424J2_126_3477_n1910, DP_OP_424J2_126_3477_n1909,
         DP_OP_424J2_126_3477_n1908, DP_OP_424J2_126_3477_n1907,
         DP_OP_424J2_126_3477_n1906, DP_OP_424J2_126_3477_n1904,
         DP_OP_424J2_126_3477_n1903, DP_OP_424J2_126_3477_n1901,
         DP_OP_424J2_126_3477_n1898, DP_OP_424J2_126_3477_n1897,
         DP_OP_424J2_126_3477_n1896, DP_OP_424J2_126_3477_n1895,
         DP_OP_424J2_126_3477_n1894, DP_OP_424J2_126_3477_n1893,
         DP_OP_424J2_126_3477_n1892, DP_OP_424J2_126_3477_n1891,
         DP_OP_424J2_126_3477_n1890, DP_OP_424J2_126_3477_n1889,
         DP_OP_424J2_126_3477_n1888, DP_OP_424J2_126_3477_n1887,
         DP_OP_424J2_126_3477_n1886, DP_OP_424J2_126_3477_n1885,
         DP_OP_424J2_126_3477_n1884, DP_OP_424J2_126_3477_n1883,
         DP_OP_424J2_126_3477_n1882, DP_OP_424J2_126_3477_n1881,
         DP_OP_424J2_126_3477_n1880, DP_OP_424J2_126_3477_n1879,
         DP_OP_424J2_126_3477_n1878, DP_OP_424J2_126_3477_n1877,
         DP_OP_424J2_126_3477_n1876, DP_OP_424J2_126_3477_n1875,
         DP_OP_424J2_126_3477_n1874, DP_OP_424J2_126_3477_n1873,
         DP_OP_424J2_126_3477_n1872, DP_OP_424J2_126_3477_n1871,
         DP_OP_424J2_126_3477_n1870, DP_OP_424J2_126_3477_n1869,
         DP_OP_424J2_126_3477_n1868, DP_OP_424J2_126_3477_n1867,
         DP_OP_424J2_126_3477_n1866, DP_OP_424J2_126_3477_n1865,
         DP_OP_424J2_126_3477_n1862, DP_OP_424J2_126_3477_n1858,
         DP_OP_424J2_126_3477_n1857, DP_OP_424J2_126_3477_n1854,
         DP_OP_424J2_126_3477_n1853, DP_OP_424J2_126_3477_n1852,
         DP_OP_424J2_126_3477_n1851, DP_OP_424J2_126_3477_n1850,
         DP_OP_424J2_126_3477_n1849, DP_OP_424J2_126_3477_n1848,
         DP_OP_424J2_126_3477_n1847, DP_OP_424J2_126_3477_n1846,
         DP_OP_424J2_126_3477_n1845, DP_OP_424J2_126_3477_n1844,
         DP_OP_424J2_126_3477_n1843, DP_OP_424J2_126_3477_n1842,
         DP_OP_424J2_126_3477_n1841, DP_OP_424J2_126_3477_n1840,
         DP_OP_424J2_126_3477_n1839, DP_OP_424J2_126_3477_n1838,
         DP_OP_424J2_126_3477_n1837, DP_OP_424J2_126_3477_n1836,
         DP_OP_424J2_126_3477_n1835, DP_OP_424J2_126_3477_n1834,
         DP_OP_424J2_126_3477_n1833, DP_OP_424J2_126_3477_n1832,
         DP_OP_424J2_126_3477_n1831, DP_OP_424J2_126_3477_n1830,
         DP_OP_424J2_126_3477_n1829, DP_OP_424J2_126_3477_n1828,
         DP_OP_424J2_126_3477_n1827, DP_OP_424J2_126_3477_n1826,
         DP_OP_424J2_126_3477_n1825, DP_OP_424J2_126_3477_n1824,
         DP_OP_424J2_126_3477_n1823, DP_OP_424J2_126_3477_n1822,
         DP_OP_424J2_126_3477_n1788, DP_OP_424J2_126_3477_n1787,
         DP_OP_424J2_126_3477_n1786, DP_OP_424J2_126_3477_n1785,
         DP_OP_424J2_126_3477_n1784, DP_OP_424J2_126_3477_n1783,
         DP_OP_424J2_126_3477_n1782, DP_OP_424J2_126_3477_n1781,
         DP_OP_424J2_126_3477_n1780, DP_OP_424J2_126_3477_n1779,
         DP_OP_424J2_126_3477_n1778, DP_OP_424J2_126_3477_n1777,
         DP_OP_424J2_126_3477_n1776, DP_OP_424J2_126_3477_n1775,
         DP_OP_424J2_126_3477_n1774, DP_OP_424J2_126_3477_n1773,
         DP_OP_424J2_126_3477_n1772, DP_OP_424J2_126_3477_n1771,
         DP_OP_424J2_126_3477_n1770, DP_OP_424J2_126_3477_n1769,
         DP_OP_424J2_126_3477_n1768, DP_OP_424J2_126_3477_n1767,
         DP_OP_424J2_126_3477_n1766, DP_OP_424J2_126_3477_n1765,
         DP_OP_424J2_126_3477_n1764, DP_OP_424J2_126_3477_n1763,
         DP_OP_424J2_126_3477_n1762, DP_OP_424J2_126_3477_n1761,
         DP_OP_424J2_126_3477_n1760, DP_OP_424J2_126_3477_n1759,
         DP_OP_424J2_126_3477_n1758, DP_OP_424J2_126_3477_n1757,
         DP_OP_424J2_126_3477_n1756, DP_OP_424J2_126_3477_n1755,
         DP_OP_424J2_126_3477_n1754, DP_OP_424J2_126_3477_n1753,
         DP_OP_424J2_126_3477_n1752, DP_OP_424J2_126_3477_n1751,
         DP_OP_424J2_126_3477_n1750, DP_OP_424J2_126_3477_n1749,
         DP_OP_424J2_126_3477_n1748, DP_OP_424J2_126_3477_n1747,
         DP_OP_424J2_126_3477_n1746, DP_OP_424J2_126_3477_n1745,
         DP_OP_424J2_126_3477_n1744, DP_OP_424J2_126_3477_n1743,
         DP_OP_424J2_126_3477_n1742, DP_OP_424J2_126_3477_n1741,
         DP_OP_424J2_126_3477_n1740, DP_OP_424J2_126_3477_n1739,
         DP_OP_424J2_126_3477_n1738, DP_OP_424J2_126_3477_n1737,
         DP_OP_424J2_126_3477_n1736, DP_OP_424J2_126_3477_n1735,
         DP_OP_424J2_126_3477_n1734, DP_OP_424J2_126_3477_n1733,
         DP_OP_424J2_126_3477_n1732, DP_OP_424J2_126_3477_n1731,
         DP_OP_424J2_126_3477_n1730, DP_OP_424J2_126_3477_n1729,
         DP_OP_424J2_126_3477_n1728, DP_OP_424J2_126_3477_n1727,
         DP_OP_424J2_126_3477_n1726, DP_OP_424J2_126_3477_n1725,
         DP_OP_424J2_126_3477_n1724, DP_OP_424J2_126_3477_n1723,
         DP_OP_424J2_126_3477_n1722, DP_OP_424J2_126_3477_n1721,
         DP_OP_424J2_126_3477_n1720, DP_OP_424J2_126_3477_n1719,
         DP_OP_424J2_126_3477_n1718, DP_OP_424J2_126_3477_n1717,
         DP_OP_424J2_126_3477_n1716, DP_OP_424J2_126_3477_n1715,
         DP_OP_424J2_126_3477_n1714, DP_OP_424J2_126_3477_n1713,
         DP_OP_424J2_126_3477_n1712, DP_OP_424J2_126_3477_n1711,
         DP_OP_424J2_126_3477_n1710, DP_OP_424J2_126_3477_n1709,
         DP_OP_424J2_126_3477_n1708, DP_OP_424J2_126_3477_n1707,
         DP_OP_424J2_126_3477_n1706, DP_OP_424J2_126_3477_n1705,
         DP_OP_424J2_126_3477_n1704, DP_OP_424J2_126_3477_n1703,
         DP_OP_424J2_126_3477_n1702, DP_OP_424J2_126_3477_n1701,
         DP_OP_424J2_126_3477_n1700, DP_OP_424J2_126_3477_n1699,
         DP_OP_424J2_126_3477_n1698, DP_OP_424J2_126_3477_n1697,
         DP_OP_424J2_126_3477_n1696, DP_OP_424J2_126_3477_n1695,
         DP_OP_424J2_126_3477_n1694, DP_OP_424J2_126_3477_n1693,
         DP_OP_424J2_126_3477_n1692, DP_OP_424J2_126_3477_n1691,
         DP_OP_424J2_126_3477_n1690, DP_OP_424J2_126_3477_n1689,
         DP_OP_424J2_126_3477_n1688, DP_OP_424J2_126_3477_n1687,
         DP_OP_424J2_126_3477_n1686, DP_OP_424J2_126_3477_n1685,
         DP_OP_424J2_126_3477_n1684, DP_OP_424J2_126_3477_n1683,
         DP_OP_424J2_126_3477_n1682, DP_OP_424J2_126_3477_n1681,
         DP_OP_424J2_126_3477_n1680, DP_OP_424J2_126_3477_n1679,
         DP_OP_424J2_126_3477_n1678, DP_OP_424J2_126_3477_n1677,
         DP_OP_424J2_126_3477_n1676, DP_OP_424J2_126_3477_n1675,
         DP_OP_424J2_126_3477_n1674, DP_OP_424J2_126_3477_n1673,
         DP_OP_424J2_126_3477_n1672, DP_OP_424J2_126_3477_n1671,
         DP_OP_424J2_126_3477_n1670, DP_OP_424J2_126_3477_n1669,
         DP_OP_424J2_126_3477_n1668, DP_OP_424J2_126_3477_n1667,
         DP_OP_424J2_126_3477_n1666, DP_OP_424J2_126_3477_n1665,
         DP_OP_424J2_126_3477_n1664, DP_OP_424J2_126_3477_n1663,
         DP_OP_424J2_126_3477_n1662, DP_OP_424J2_126_3477_n1661,
         DP_OP_424J2_126_3477_n1660, DP_OP_424J2_126_3477_n1659,
         DP_OP_424J2_126_3477_n1658, DP_OP_424J2_126_3477_n1657,
         DP_OP_424J2_126_3477_n1656, DP_OP_424J2_126_3477_n1655,
         DP_OP_424J2_126_3477_n1654, DP_OP_424J2_126_3477_n1653,
         DP_OP_424J2_126_3477_n1652, DP_OP_424J2_126_3477_n1651,
         DP_OP_424J2_126_3477_n1650, DP_OP_424J2_126_3477_n1649,
         DP_OP_424J2_126_3477_n1648, DP_OP_424J2_126_3477_n1647,
         DP_OP_424J2_126_3477_n1646, DP_OP_424J2_126_3477_n1645,
         DP_OP_424J2_126_3477_n1644, DP_OP_424J2_126_3477_n1643,
         DP_OP_424J2_126_3477_n1642, DP_OP_424J2_126_3477_n1641,
         DP_OP_424J2_126_3477_n1640, DP_OP_424J2_126_3477_n1639,
         DP_OP_424J2_126_3477_n1638, DP_OP_424J2_126_3477_n1637,
         DP_OP_424J2_126_3477_n1636, DP_OP_424J2_126_3477_n1635,
         DP_OP_424J2_126_3477_n1634, DP_OP_424J2_126_3477_n1633,
         DP_OP_424J2_126_3477_n1632, DP_OP_424J2_126_3477_n1631,
         DP_OP_424J2_126_3477_n1630, DP_OP_424J2_126_3477_n1629,
         DP_OP_424J2_126_3477_n1628, DP_OP_424J2_126_3477_n1627,
         DP_OP_424J2_126_3477_n1626, DP_OP_424J2_126_3477_n1625,
         DP_OP_424J2_126_3477_n1624, DP_OP_424J2_126_3477_n1623,
         DP_OP_424J2_126_3477_n1622, DP_OP_424J2_126_3477_n1621,
         DP_OP_424J2_126_3477_n1620, DP_OP_424J2_126_3477_n1619,
         DP_OP_424J2_126_3477_n1618, DP_OP_424J2_126_3477_n1617,
         DP_OP_424J2_126_3477_n1616, DP_OP_424J2_126_3477_n1615,
         DP_OP_424J2_126_3477_n1614, DP_OP_424J2_126_3477_n1613,
         DP_OP_424J2_126_3477_n1612, DP_OP_424J2_126_3477_n1611,
         DP_OP_424J2_126_3477_n1610, DP_OP_424J2_126_3477_n1609,
         DP_OP_424J2_126_3477_n1608, DP_OP_424J2_126_3477_n1607,
         DP_OP_424J2_126_3477_n1606, DP_OP_424J2_126_3477_n1605,
         DP_OP_424J2_126_3477_n1604, DP_OP_424J2_126_3477_n1603,
         DP_OP_424J2_126_3477_n1602, DP_OP_424J2_126_3477_n1601,
         DP_OP_424J2_126_3477_n1600, DP_OP_424J2_126_3477_n1599,
         DP_OP_424J2_126_3477_n1598, DP_OP_424J2_126_3477_n1597,
         DP_OP_424J2_126_3477_n1596, DP_OP_424J2_126_3477_n1595,
         DP_OP_424J2_126_3477_n1594, DP_OP_424J2_126_3477_n1593,
         DP_OP_424J2_126_3477_n1592, DP_OP_424J2_126_3477_n1591,
         DP_OP_424J2_126_3477_n1590, DP_OP_424J2_126_3477_n1589,
         DP_OP_424J2_126_3477_n1588, DP_OP_424J2_126_3477_n1587,
         DP_OP_424J2_126_3477_n1586, DP_OP_424J2_126_3477_n1585,
         DP_OP_424J2_126_3477_n1584, DP_OP_424J2_126_3477_n1583,
         DP_OP_424J2_126_3477_n1582, DP_OP_424J2_126_3477_n1581,
         DP_OP_424J2_126_3477_n1580, DP_OP_424J2_126_3477_n1579,
         DP_OP_424J2_126_3477_n1578, DP_OP_424J2_126_3477_n1577,
         DP_OP_424J2_126_3477_n1576, DP_OP_424J2_126_3477_n1575,
         DP_OP_424J2_126_3477_n1574, DP_OP_424J2_126_3477_n1573,
         DP_OP_424J2_126_3477_n1572, DP_OP_424J2_126_3477_n1571,
         DP_OP_424J2_126_3477_n1570, DP_OP_424J2_126_3477_n1569,
         DP_OP_424J2_126_3477_n1568, DP_OP_424J2_126_3477_n1567,
         DP_OP_424J2_126_3477_n1566, DP_OP_424J2_126_3477_n1565,
         DP_OP_424J2_126_3477_n1564, DP_OP_424J2_126_3477_n1563,
         DP_OP_424J2_126_3477_n1562, DP_OP_424J2_126_3477_n1561,
         DP_OP_424J2_126_3477_n1560, DP_OP_424J2_126_3477_n1559,
         DP_OP_424J2_126_3477_n1558, DP_OP_424J2_126_3477_n1557,
         DP_OP_424J2_126_3477_n1556, DP_OP_424J2_126_3477_n1555,
         DP_OP_424J2_126_3477_n1554, DP_OP_424J2_126_3477_n1553,
         DP_OP_424J2_126_3477_n1552, DP_OP_424J2_126_3477_n1551,
         DP_OP_424J2_126_3477_n1550, DP_OP_424J2_126_3477_n1549,
         DP_OP_424J2_126_3477_n1548, DP_OP_424J2_126_3477_n1547,
         DP_OP_424J2_126_3477_n1546, DP_OP_424J2_126_3477_n1545,
         DP_OP_424J2_126_3477_n1544, DP_OP_424J2_126_3477_n1543,
         DP_OP_424J2_126_3477_n1542, DP_OP_424J2_126_3477_n1541,
         DP_OP_424J2_126_3477_n1540, DP_OP_424J2_126_3477_n1539,
         DP_OP_424J2_126_3477_n1538, DP_OP_424J2_126_3477_n1537,
         DP_OP_424J2_126_3477_n1536, DP_OP_424J2_126_3477_n1535,
         DP_OP_424J2_126_3477_n1534, DP_OP_424J2_126_3477_n1533,
         DP_OP_424J2_126_3477_n1532, DP_OP_424J2_126_3477_n1531,
         DP_OP_424J2_126_3477_n1530, DP_OP_424J2_126_3477_n1529,
         DP_OP_424J2_126_3477_n1528, DP_OP_424J2_126_3477_n1527,
         DP_OP_424J2_126_3477_n1526, DP_OP_424J2_126_3477_n1525,
         DP_OP_424J2_126_3477_n1524, DP_OP_424J2_126_3477_n1523,
         DP_OP_424J2_126_3477_n1522, DP_OP_424J2_126_3477_n1521,
         DP_OP_424J2_126_3477_n1520, DP_OP_424J2_126_3477_n1519,
         DP_OP_424J2_126_3477_n1518, DP_OP_424J2_126_3477_n1517,
         DP_OP_424J2_126_3477_n1516, DP_OP_424J2_126_3477_n1515,
         DP_OP_424J2_126_3477_n1514, DP_OP_424J2_126_3477_n1513,
         DP_OP_424J2_126_3477_n1512, DP_OP_424J2_126_3477_n1511,
         DP_OP_424J2_126_3477_n1510, DP_OP_424J2_126_3477_n1509,
         DP_OP_424J2_126_3477_n1508, DP_OP_424J2_126_3477_n1507,
         DP_OP_424J2_126_3477_n1506, DP_OP_424J2_126_3477_n1505,
         DP_OP_424J2_126_3477_n1504, DP_OP_424J2_126_3477_n1503,
         DP_OP_424J2_126_3477_n1502, DP_OP_424J2_126_3477_n1501,
         DP_OP_424J2_126_3477_n1500, DP_OP_424J2_126_3477_n1499,
         DP_OP_424J2_126_3477_n1498, DP_OP_424J2_126_3477_n1497,
         DP_OP_424J2_126_3477_n1496, DP_OP_424J2_126_3477_n1495,
         DP_OP_424J2_126_3477_n1494, DP_OP_424J2_126_3477_n1493,
         DP_OP_424J2_126_3477_n1492, DP_OP_424J2_126_3477_n1491,
         DP_OP_424J2_126_3477_n1490, DP_OP_424J2_126_3477_n1489,
         DP_OP_424J2_126_3477_n1488, DP_OP_424J2_126_3477_n1487,
         DP_OP_424J2_126_3477_n1486, DP_OP_424J2_126_3477_n1485,
         DP_OP_424J2_126_3477_n1484, DP_OP_424J2_126_3477_n1483,
         DP_OP_424J2_126_3477_n1482, DP_OP_424J2_126_3477_n1481,
         DP_OP_424J2_126_3477_n1480, DP_OP_424J2_126_3477_n1479,
         DP_OP_424J2_126_3477_n1478, DP_OP_424J2_126_3477_n1477,
         DP_OP_424J2_126_3477_n1476, DP_OP_424J2_126_3477_n1475,
         DP_OP_424J2_126_3477_n1474, DP_OP_424J2_126_3477_n1473,
         DP_OP_424J2_126_3477_n1472, DP_OP_424J2_126_3477_n1471,
         DP_OP_424J2_126_3477_n1470, DP_OP_424J2_126_3477_n1469,
         DP_OP_424J2_126_3477_n1468, DP_OP_424J2_126_3477_n1467,
         DP_OP_424J2_126_3477_n1466, DP_OP_424J2_126_3477_n1465,
         DP_OP_424J2_126_3477_n1464, DP_OP_424J2_126_3477_n1463,
         DP_OP_424J2_126_3477_n1462, DP_OP_424J2_126_3477_n1461,
         DP_OP_424J2_126_3477_n1460, DP_OP_424J2_126_3477_n1459,
         DP_OP_424J2_126_3477_n1458, DP_OP_424J2_126_3477_n1457,
         DP_OP_424J2_126_3477_n1456, DP_OP_424J2_126_3477_n1455,
         DP_OP_424J2_126_3477_n1454, DP_OP_424J2_126_3477_n1453,
         DP_OP_424J2_126_3477_n1452, DP_OP_424J2_126_3477_n1451,
         DP_OP_424J2_126_3477_n1450, DP_OP_424J2_126_3477_n1449,
         DP_OP_424J2_126_3477_n1448, DP_OP_424J2_126_3477_n1447,
         DP_OP_424J2_126_3477_n1446, DP_OP_424J2_126_3477_n1445,
         DP_OP_424J2_126_3477_n1444, DP_OP_424J2_126_3477_n1443,
         DP_OP_424J2_126_3477_n1442, DP_OP_424J2_126_3477_n1441,
         DP_OP_424J2_126_3477_n1440, DP_OP_424J2_126_3477_n1439,
         DP_OP_424J2_126_3477_n1438, DP_OP_424J2_126_3477_n1437,
         DP_OP_424J2_126_3477_n1436, DP_OP_424J2_126_3477_n1435,
         DP_OP_424J2_126_3477_n1434, DP_OP_424J2_126_3477_n1433,
         DP_OP_424J2_126_3477_n1432, DP_OP_424J2_126_3477_n1431,
         DP_OP_424J2_126_3477_n1430, DP_OP_424J2_126_3477_n1429,
         DP_OP_424J2_126_3477_n1428, DP_OP_424J2_126_3477_n1427,
         DP_OP_424J2_126_3477_n1426, DP_OP_424J2_126_3477_n1425,
         DP_OP_424J2_126_3477_n1424, DP_OP_424J2_126_3477_n1423,
         DP_OP_424J2_126_3477_n1422, DP_OP_424J2_126_3477_n1421,
         DP_OP_424J2_126_3477_n1420, DP_OP_424J2_126_3477_n1419,
         DP_OP_424J2_126_3477_n1418, DP_OP_424J2_126_3477_n1417,
         DP_OP_424J2_126_3477_n1416, DP_OP_424J2_126_3477_n1415,
         DP_OP_424J2_126_3477_n1414, DP_OP_424J2_126_3477_n1413,
         DP_OP_424J2_126_3477_n1412, DP_OP_424J2_126_3477_n1411,
         DP_OP_424J2_126_3477_n1410, DP_OP_424J2_126_3477_n1409,
         DP_OP_424J2_126_3477_n1408, DP_OP_424J2_126_3477_n1407,
         DP_OP_424J2_126_3477_n1406, DP_OP_424J2_126_3477_n1405,
         DP_OP_424J2_126_3477_n1404, DP_OP_424J2_126_3477_n1403,
         DP_OP_424J2_126_3477_n1402, DP_OP_424J2_126_3477_n1401,
         DP_OP_424J2_126_3477_n1400, DP_OP_424J2_126_3477_n1399,
         DP_OP_424J2_126_3477_n1398, DP_OP_424J2_126_3477_n1397,
         DP_OP_424J2_126_3477_n1396, DP_OP_424J2_126_3477_n1395,
         DP_OP_424J2_126_3477_n1394, DP_OP_424J2_126_3477_n1393,
         DP_OP_424J2_126_3477_n1392, DP_OP_424J2_126_3477_n1391,
         DP_OP_424J2_126_3477_n1390, DP_OP_424J2_126_3477_n1389,
         DP_OP_424J2_126_3477_n1388, DP_OP_424J2_126_3477_n1387,
         DP_OP_424J2_126_3477_n1386, DP_OP_424J2_126_3477_n1385,
         DP_OP_424J2_126_3477_n1384, DP_OP_424J2_126_3477_n1383,
         DP_OP_424J2_126_3477_n1382, DP_OP_424J2_126_3477_n1381,
         DP_OP_424J2_126_3477_n1380, DP_OP_424J2_126_3477_n1379,
         DP_OP_424J2_126_3477_n1378, DP_OP_424J2_126_3477_n1377,
         DP_OP_424J2_126_3477_n1376, DP_OP_424J2_126_3477_n1375,
         DP_OP_424J2_126_3477_n1374, DP_OP_424J2_126_3477_n1373,
         DP_OP_424J2_126_3477_n1372, DP_OP_424J2_126_3477_n1371,
         DP_OP_424J2_126_3477_n1370, DP_OP_424J2_126_3477_n1369,
         DP_OP_424J2_126_3477_n1368, DP_OP_424J2_126_3477_n1367,
         DP_OP_424J2_126_3477_n1366, DP_OP_424J2_126_3477_n1365,
         DP_OP_424J2_126_3477_n1364, DP_OP_424J2_126_3477_n1363,
         DP_OP_424J2_126_3477_n1362, DP_OP_424J2_126_3477_n1361,
         DP_OP_424J2_126_3477_n1360, DP_OP_424J2_126_3477_n1359,
         DP_OP_424J2_126_3477_n1358, DP_OP_424J2_126_3477_n1357,
         DP_OP_424J2_126_3477_n1356, DP_OP_424J2_126_3477_n1355,
         DP_OP_424J2_126_3477_n1354, DP_OP_424J2_126_3477_n1353,
         DP_OP_424J2_126_3477_n1352, DP_OP_424J2_126_3477_n1351,
         DP_OP_424J2_126_3477_n1350, DP_OP_424J2_126_3477_n1349,
         DP_OP_424J2_126_3477_n1348, DP_OP_424J2_126_3477_n1347,
         DP_OP_424J2_126_3477_n1346, DP_OP_424J2_126_3477_n1345,
         DP_OP_424J2_126_3477_n1344, DP_OP_424J2_126_3477_n1343,
         DP_OP_424J2_126_3477_n1342, DP_OP_424J2_126_3477_n1341,
         DP_OP_424J2_126_3477_n1340, DP_OP_424J2_126_3477_n1339,
         DP_OP_424J2_126_3477_n1338, DP_OP_424J2_126_3477_n1337,
         DP_OP_424J2_126_3477_n1336, DP_OP_424J2_126_3477_n1335,
         DP_OP_424J2_126_3477_n1334, DP_OP_424J2_126_3477_n1333,
         DP_OP_424J2_126_3477_n1332, DP_OP_424J2_126_3477_n1331,
         DP_OP_424J2_126_3477_n1330, DP_OP_424J2_126_3477_n1329,
         DP_OP_424J2_126_3477_n1328, DP_OP_424J2_126_3477_n1327,
         DP_OP_424J2_126_3477_n1326, DP_OP_424J2_126_3477_n1325,
         DP_OP_424J2_126_3477_n1324, DP_OP_424J2_126_3477_n1323,
         DP_OP_424J2_126_3477_n1322, DP_OP_424J2_126_3477_n1321,
         DP_OP_424J2_126_3477_n1320, DP_OP_424J2_126_3477_n1319,
         DP_OP_424J2_126_3477_n1318, DP_OP_424J2_126_3477_n1317,
         DP_OP_424J2_126_3477_n1316, DP_OP_424J2_126_3477_n1315,
         DP_OP_424J2_126_3477_n1314, DP_OP_424J2_126_3477_n1313,
         DP_OP_424J2_126_3477_n1312, DP_OP_424J2_126_3477_n1311,
         DP_OP_424J2_126_3477_n1310, DP_OP_424J2_126_3477_n1309,
         DP_OP_424J2_126_3477_n1308, DP_OP_424J2_126_3477_n1307,
         DP_OP_424J2_126_3477_n1306, DP_OP_424J2_126_3477_n1305,
         DP_OP_424J2_126_3477_n1304, DP_OP_424J2_126_3477_n1303,
         DP_OP_424J2_126_3477_n1302, DP_OP_424J2_126_3477_n1301,
         DP_OP_424J2_126_3477_n1300, DP_OP_424J2_126_3477_n1299,
         DP_OP_424J2_126_3477_n1298, DP_OP_424J2_126_3477_n1297,
         DP_OP_424J2_126_3477_n1296, DP_OP_424J2_126_3477_n1295,
         DP_OP_424J2_126_3477_n1294, DP_OP_424J2_126_3477_n1293,
         DP_OP_424J2_126_3477_n1292, DP_OP_424J2_126_3477_n1291,
         DP_OP_424J2_126_3477_n1290, DP_OP_424J2_126_3477_n1289,
         DP_OP_424J2_126_3477_n1288, DP_OP_424J2_126_3477_n1287,
         DP_OP_424J2_126_3477_n1286, DP_OP_424J2_126_3477_n1285,
         DP_OP_424J2_126_3477_n1284, DP_OP_424J2_126_3477_n1283,
         DP_OP_424J2_126_3477_n1282, DP_OP_424J2_126_3477_n1281,
         DP_OP_424J2_126_3477_n1280, DP_OP_424J2_126_3477_n1279,
         DP_OP_424J2_126_3477_n1278, DP_OP_424J2_126_3477_n1277,
         DP_OP_424J2_126_3477_n1276, DP_OP_424J2_126_3477_n1275,
         DP_OP_424J2_126_3477_n1274, DP_OP_424J2_126_3477_n1273,
         DP_OP_424J2_126_3477_n1272, DP_OP_424J2_126_3477_n1271,
         DP_OP_424J2_126_3477_n1270, DP_OP_424J2_126_3477_n1269,
         DP_OP_424J2_126_3477_n1268, DP_OP_424J2_126_3477_n1267,
         DP_OP_424J2_126_3477_n1266, DP_OP_424J2_126_3477_n1265,
         DP_OP_424J2_126_3477_n1264, DP_OP_424J2_126_3477_n1263,
         DP_OP_424J2_126_3477_n1262, DP_OP_424J2_126_3477_n1261,
         DP_OP_424J2_126_3477_n1260, DP_OP_424J2_126_3477_n1259,
         DP_OP_424J2_126_3477_n1258, DP_OP_424J2_126_3477_n1257,
         DP_OP_424J2_126_3477_n1256, DP_OP_424J2_126_3477_n1255,
         DP_OP_424J2_126_3477_n1254, DP_OP_424J2_126_3477_n1253,
         DP_OP_424J2_126_3477_n1252, DP_OP_424J2_126_3477_n1251,
         DP_OP_424J2_126_3477_n1250, DP_OP_424J2_126_3477_n1249,
         DP_OP_424J2_126_3477_n1248, DP_OP_424J2_126_3477_n1247,
         DP_OP_424J2_126_3477_n1246, DP_OP_424J2_126_3477_n1245,
         DP_OP_424J2_126_3477_n1244, DP_OP_424J2_126_3477_n1243,
         DP_OP_424J2_126_3477_n1242, DP_OP_424J2_126_3477_n1241,
         DP_OP_424J2_126_3477_n1240, DP_OP_424J2_126_3477_n1239,
         DP_OP_424J2_126_3477_n1238, DP_OP_424J2_126_3477_n1237,
         DP_OP_424J2_126_3477_n1236, DP_OP_424J2_126_3477_n1235,
         DP_OP_424J2_126_3477_n1234, DP_OP_424J2_126_3477_n1233,
         DP_OP_424J2_126_3477_n1232, DP_OP_424J2_126_3477_n1231,
         DP_OP_424J2_126_3477_n1230, DP_OP_424J2_126_3477_n1229,
         DP_OP_424J2_126_3477_n1228, DP_OP_424J2_126_3477_n1227,
         DP_OP_424J2_126_3477_n1226, DP_OP_424J2_126_3477_n1225,
         DP_OP_424J2_126_3477_n1224, DP_OP_424J2_126_3477_n1223,
         DP_OP_424J2_126_3477_n1222, DP_OP_424J2_126_3477_n1221,
         DP_OP_424J2_126_3477_n1220, DP_OP_424J2_126_3477_n1219,
         DP_OP_424J2_126_3477_n1218, DP_OP_424J2_126_3477_n1217,
         DP_OP_424J2_126_3477_n1216, DP_OP_424J2_126_3477_n1215,
         DP_OP_424J2_126_3477_n1214, DP_OP_424J2_126_3477_n1213,
         DP_OP_424J2_126_3477_n1212, DP_OP_424J2_126_3477_n1211,
         DP_OP_424J2_126_3477_n1210, DP_OP_424J2_126_3477_n1209,
         DP_OP_424J2_126_3477_n1208, DP_OP_424J2_126_3477_n1207,
         DP_OP_424J2_126_3477_n1206, DP_OP_424J2_126_3477_n1205,
         DP_OP_424J2_126_3477_n1204, DP_OP_424J2_126_3477_n1203,
         DP_OP_424J2_126_3477_n1202, DP_OP_424J2_126_3477_n1201,
         DP_OP_424J2_126_3477_n1200, DP_OP_424J2_126_3477_n1199,
         DP_OP_424J2_126_3477_n1198, DP_OP_424J2_126_3477_n1197,
         DP_OP_424J2_126_3477_n1196, DP_OP_424J2_126_3477_n1195,
         DP_OP_424J2_126_3477_n1194, DP_OP_424J2_126_3477_n1193,
         DP_OP_424J2_126_3477_n1192, DP_OP_424J2_126_3477_n1191,
         DP_OP_424J2_126_3477_n1190, DP_OP_424J2_126_3477_n1189,
         DP_OP_424J2_126_3477_n1188, DP_OP_424J2_126_3477_n1187,
         DP_OP_424J2_126_3477_n1186, DP_OP_424J2_126_3477_n1185,
         DP_OP_424J2_126_3477_n1184, DP_OP_424J2_126_3477_n1183,
         DP_OP_424J2_126_3477_n1182, DP_OP_424J2_126_3477_n1181,
         DP_OP_424J2_126_3477_n1180, DP_OP_424J2_126_3477_n1179,
         DP_OP_424J2_126_3477_n1178, DP_OP_424J2_126_3477_n1177,
         DP_OP_424J2_126_3477_n1176, DP_OP_424J2_126_3477_n1175,
         DP_OP_424J2_126_3477_n1174, DP_OP_424J2_126_3477_n1173,
         DP_OP_424J2_126_3477_n1172, DP_OP_424J2_126_3477_n1171,
         DP_OP_424J2_126_3477_n1170, DP_OP_424J2_126_3477_n1169,
         DP_OP_424J2_126_3477_n1168, DP_OP_424J2_126_3477_n1167,
         DP_OP_424J2_126_3477_n1166, DP_OP_424J2_126_3477_n1165,
         DP_OP_424J2_126_3477_n1164, DP_OP_424J2_126_3477_n1163,
         DP_OP_424J2_126_3477_n1162, DP_OP_424J2_126_3477_n1161,
         DP_OP_424J2_126_3477_n1160, DP_OP_424J2_126_3477_n1159,
         DP_OP_424J2_126_3477_n1158, DP_OP_424J2_126_3477_n1157,
         DP_OP_424J2_126_3477_n1156, DP_OP_424J2_126_3477_n1155,
         DP_OP_424J2_126_3477_n1154, DP_OP_424J2_126_3477_n1153,
         DP_OP_424J2_126_3477_n1152, DP_OP_424J2_126_3477_n1151,
         DP_OP_424J2_126_3477_n1150, DP_OP_424J2_126_3477_n1149,
         DP_OP_424J2_126_3477_n1148, DP_OP_424J2_126_3477_n1147,
         DP_OP_424J2_126_3477_n1146, DP_OP_424J2_126_3477_n1145,
         DP_OP_424J2_126_3477_n1144, DP_OP_424J2_126_3477_n1143,
         DP_OP_424J2_126_3477_n1142, DP_OP_424J2_126_3477_n1141,
         DP_OP_424J2_126_3477_n1140, DP_OP_424J2_126_3477_n1139,
         DP_OP_424J2_126_3477_n1138, DP_OP_424J2_126_3477_n1137,
         DP_OP_424J2_126_3477_n1136, DP_OP_424J2_126_3477_n1135,
         DP_OP_424J2_126_3477_n1134, DP_OP_424J2_126_3477_n1133,
         DP_OP_424J2_126_3477_n1132, DP_OP_424J2_126_3477_n1131,
         DP_OP_424J2_126_3477_n1130, DP_OP_424J2_126_3477_n1129,
         DP_OP_424J2_126_3477_n1128, DP_OP_424J2_126_3477_n1127,
         DP_OP_424J2_126_3477_n1126, DP_OP_424J2_126_3477_n1125,
         DP_OP_424J2_126_3477_n1124, DP_OP_424J2_126_3477_n1123,
         DP_OP_424J2_126_3477_n1122, DP_OP_424J2_126_3477_n1121,
         DP_OP_424J2_126_3477_n1120, DP_OP_424J2_126_3477_n1119,
         DP_OP_424J2_126_3477_n1118, DP_OP_424J2_126_3477_n1117,
         DP_OP_424J2_126_3477_n1116, DP_OP_424J2_126_3477_n1115,
         DP_OP_424J2_126_3477_n1114, DP_OP_424J2_126_3477_n1113,
         DP_OP_424J2_126_3477_n1112, DP_OP_424J2_126_3477_n1111,
         DP_OP_424J2_126_3477_n1110, DP_OP_424J2_126_3477_n1109,
         DP_OP_424J2_126_3477_n1108, DP_OP_424J2_126_3477_n1107,
         DP_OP_424J2_126_3477_n1106, DP_OP_424J2_126_3477_n1105,
         DP_OP_424J2_126_3477_n1104, DP_OP_424J2_126_3477_n1103,
         DP_OP_424J2_126_3477_n1102, DP_OP_424J2_126_3477_n1101,
         DP_OP_424J2_126_3477_n1100, DP_OP_424J2_126_3477_n1099,
         DP_OP_424J2_126_3477_n1098, DP_OP_424J2_126_3477_n1097,
         DP_OP_424J2_126_3477_n1096, DP_OP_424J2_126_3477_n1095,
         DP_OP_424J2_126_3477_n1094, DP_OP_424J2_126_3477_n1093,
         DP_OP_424J2_126_3477_n1092, DP_OP_424J2_126_3477_n1091,
         DP_OP_424J2_126_3477_n1090, DP_OP_424J2_126_3477_n1089,
         DP_OP_424J2_126_3477_n1088, DP_OP_424J2_126_3477_n1087,
         DP_OP_424J2_126_3477_n1086, DP_OP_424J2_126_3477_n1085,
         DP_OP_424J2_126_3477_n1084, DP_OP_424J2_126_3477_n1083,
         DP_OP_424J2_126_3477_n1082, DP_OP_424J2_126_3477_n1081,
         DP_OP_424J2_126_3477_n1080, DP_OP_424J2_126_3477_n1079,
         DP_OP_424J2_126_3477_n1078, DP_OP_424J2_126_3477_n1077,
         DP_OP_424J2_126_3477_n1076, DP_OP_424J2_126_3477_n1075,
         DP_OP_424J2_126_3477_n1074, DP_OP_424J2_126_3477_n1073,
         DP_OP_424J2_126_3477_n1072, DP_OP_424J2_126_3477_n1071,
         DP_OP_424J2_126_3477_n1070, DP_OP_424J2_126_3477_n1069,
         DP_OP_424J2_126_3477_n1068, DP_OP_424J2_126_3477_n1067,
         DP_OP_424J2_126_3477_n1066, DP_OP_424J2_126_3477_n1065,
         DP_OP_424J2_126_3477_n1064, DP_OP_424J2_126_3477_n1063,
         DP_OP_424J2_126_3477_n1062, DP_OP_424J2_126_3477_n1061,
         DP_OP_424J2_126_3477_n1060, DP_OP_424J2_126_3477_n1059,
         DP_OP_424J2_126_3477_n1058, DP_OP_424J2_126_3477_n1057,
         DP_OP_424J2_126_3477_n1056, DP_OP_424J2_126_3477_n1055,
         DP_OP_424J2_126_3477_n1054, DP_OP_424J2_126_3477_n1053,
         DP_OP_424J2_126_3477_n1052, DP_OP_424J2_126_3477_n1051,
         DP_OP_424J2_126_3477_n1050, DP_OP_424J2_126_3477_n1049,
         DP_OP_424J2_126_3477_n1048, DP_OP_424J2_126_3477_n1047,
         DP_OP_424J2_126_3477_n1046, DP_OP_424J2_126_3477_n1045,
         DP_OP_424J2_126_3477_n1044, DP_OP_424J2_126_3477_n1043,
         DP_OP_424J2_126_3477_n1042, DP_OP_424J2_126_3477_n1041,
         DP_OP_424J2_126_3477_n1040, DP_OP_424J2_126_3477_n1039,
         DP_OP_424J2_126_3477_n1038, DP_OP_424J2_126_3477_n1037,
         DP_OP_424J2_126_3477_n1036, DP_OP_424J2_126_3477_n1035,
         DP_OP_424J2_126_3477_n1034, DP_OP_424J2_126_3477_n1033,
         DP_OP_424J2_126_3477_n1032, DP_OP_424J2_126_3477_n1031,
         DP_OP_424J2_126_3477_n1030, DP_OP_424J2_126_3477_n1029,
         DP_OP_424J2_126_3477_n1028, DP_OP_424J2_126_3477_n1027,
         DP_OP_424J2_126_3477_n1026, DP_OP_424J2_126_3477_n1025,
         DP_OP_424J2_126_3477_n1024, DP_OP_424J2_126_3477_n1023,
         DP_OP_424J2_126_3477_n1022, DP_OP_424J2_126_3477_n1021,
         DP_OP_424J2_126_3477_n1020, DP_OP_424J2_126_3477_n1019,
         DP_OP_424J2_126_3477_n1018, DP_OP_424J2_126_3477_n1017,
         DP_OP_424J2_126_3477_n1016, DP_OP_424J2_126_3477_n1015,
         DP_OP_424J2_126_3477_n1014, DP_OP_424J2_126_3477_n1013,
         DP_OP_424J2_126_3477_n1012, DP_OP_424J2_126_3477_n1011,
         DP_OP_424J2_126_3477_n1010, DP_OP_424J2_126_3477_n1009,
         DP_OP_424J2_126_3477_n1008, DP_OP_424J2_126_3477_n1007,
         DP_OP_424J2_126_3477_n1006, DP_OP_424J2_126_3477_n1005,
         DP_OP_424J2_126_3477_n1004, DP_OP_424J2_126_3477_n1003,
         DP_OP_424J2_126_3477_n1002, DP_OP_424J2_126_3477_n1001,
         DP_OP_424J2_126_3477_n1000, DP_OP_424J2_126_3477_n999,
         DP_OP_424J2_126_3477_n998, DP_OP_424J2_126_3477_n997,
         DP_OP_424J2_126_3477_n996, DP_OP_424J2_126_3477_n995,
         DP_OP_424J2_126_3477_n994, DP_OP_424J2_126_3477_n993,
         DP_OP_424J2_126_3477_n992, DP_OP_424J2_126_3477_n991,
         DP_OP_424J2_126_3477_n990, DP_OP_424J2_126_3477_n989,
         DP_OP_424J2_126_3477_n988, DP_OP_424J2_126_3477_n987,
         DP_OP_424J2_126_3477_n986, DP_OP_424J2_126_3477_n985,
         DP_OP_424J2_126_3477_n984, DP_OP_424J2_126_3477_n983,
         DP_OP_424J2_126_3477_n982, DP_OP_424J2_126_3477_n981,
         DP_OP_424J2_126_3477_n980, DP_OP_424J2_126_3477_n979,
         DP_OP_424J2_126_3477_n978, DP_OP_424J2_126_3477_n977,
         DP_OP_424J2_126_3477_n976, DP_OP_424J2_126_3477_n975,
         DP_OP_424J2_126_3477_n974, DP_OP_424J2_126_3477_n973,
         DP_OP_424J2_126_3477_n972, DP_OP_424J2_126_3477_n971,
         DP_OP_424J2_126_3477_n970, DP_OP_424J2_126_3477_n969,
         DP_OP_424J2_126_3477_n968, DP_OP_424J2_126_3477_n967,
         DP_OP_424J2_126_3477_n966, DP_OP_424J2_126_3477_n965,
         DP_OP_424J2_126_3477_n964, DP_OP_424J2_126_3477_n963,
         DP_OP_424J2_126_3477_n962, DP_OP_424J2_126_3477_n961,
         DP_OP_424J2_126_3477_n960, DP_OP_424J2_126_3477_n959,
         DP_OP_424J2_126_3477_n958, DP_OP_424J2_126_3477_n957,
         DP_OP_424J2_126_3477_n956, DP_OP_424J2_126_3477_n955,
         DP_OP_424J2_126_3477_n954, DP_OP_424J2_126_3477_n953,
         DP_OP_424J2_126_3477_n952, DP_OP_424J2_126_3477_n951,
         DP_OP_424J2_126_3477_n950, DP_OP_424J2_126_3477_n949,
         DP_OP_424J2_126_3477_n948, DP_OP_424J2_126_3477_n947,
         DP_OP_424J2_126_3477_n946, DP_OP_424J2_126_3477_n945,
         DP_OP_424J2_126_3477_n944, DP_OP_424J2_126_3477_n943,
         DP_OP_424J2_126_3477_n942, DP_OP_424J2_126_3477_n941,
         DP_OP_424J2_126_3477_n940, DP_OP_424J2_126_3477_n939,
         DP_OP_424J2_126_3477_n938, DP_OP_424J2_126_3477_n937,
         DP_OP_424J2_126_3477_n936, DP_OP_424J2_126_3477_n935,
         DP_OP_424J2_126_3477_n934, DP_OP_424J2_126_3477_n933,
         DP_OP_424J2_126_3477_n932, DP_OP_424J2_126_3477_n931,
         DP_OP_424J2_126_3477_n930, DP_OP_424J2_126_3477_n929,
         DP_OP_424J2_126_3477_n928, DP_OP_424J2_126_3477_n927,
         DP_OP_424J2_126_3477_n926, DP_OP_424J2_126_3477_n925,
         DP_OP_424J2_126_3477_n924, DP_OP_424J2_126_3477_n923,
         DP_OP_424J2_126_3477_n922, DP_OP_424J2_126_3477_n921,
         DP_OP_424J2_126_3477_n920, DP_OP_424J2_126_3477_n919,
         DP_OP_424J2_126_3477_n918, DP_OP_424J2_126_3477_n917,
         DP_OP_424J2_126_3477_n916, DP_OP_424J2_126_3477_n915,
         DP_OP_424J2_126_3477_n914, DP_OP_424J2_126_3477_n913,
         DP_OP_424J2_126_3477_n912, DP_OP_424J2_126_3477_n911,
         DP_OP_424J2_126_3477_n910, DP_OP_424J2_126_3477_n909,
         DP_OP_424J2_126_3477_n908, DP_OP_424J2_126_3477_n907,
         DP_OP_424J2_126_3477_n906, DP_OP_424J2_126_3477_n905,
         DP_OP_424J2_126_3477_n904, DP_OP_424J2_126_3477_n903,
         DP_OP_424J2_126_3477_n902, DP_OP_424J2_126_3477_n901,
         DP_OP_424J2_126_3477_n900, DP_OP_424J2_126_3477_n899,
         DP_OP_424J2_126_3477_n898, DP_OP_424J2_126_3477_n897,
         DP_OP_424J2_126_3477_n896, DP_OP_424J2_126_3477_n895,
         DP_OP_424J2_126_3477_n894, DP_OP_424J2_126_3477_n893,
         DP_OP_424J2_126_3477_n892, DP_OP_424J2_126_3477_n891,
         DP_OP_424J2_126_3477_n890, DP_OP_424J2_126_3477_n889,
         DP_OP_424J2_126_3477_n888, DP_OP_424J2_126_3477_n887,
         DP_OP_424J2_126_3477_n886, DP_OP_424J2_126_3477_n885,
         DP_OP_424J2_126_3477_n884, DP_OP_424J2_126_3477_n883,
         DP_OP_424J2_126_3477_n882, DP_OP_424J2_126_3477_n881,
         DP_OP_424J2_126_3477_n880, DP_OP_424J2_126_3477_n879,
         DP_OP_424J2_126_3477_n878, DP_OP_424J2_126_3477_n877,
         DP_OP_424J2_126_3477_n876, DP_OP_424J2_126_3477_n875,
         DP_OP_424J2_126_3477_n874, DP_OP_424J2_126_3477_n873,
         DP_OP_424J2_126_3477_n872, DP_OP_424J2_126_3477_n871,
         DP_OP_424J2_126_3477_n870, DP_OP_424J2_126_3477_n869,
         DP_OP_424J2_126_3477_n868, DP_OP_424J2_126_3477_n867,
         DP_OP_424J2_126_3477_n866, DP_OP_424J2_126_3477_n865,
         DP_OP_424J2_126_3477_n864, DP_OP_424J2_126_3477_n863,
         DP_OP_424J2_126_3477_n862, DP_OP_424J2_126_3477_n861,
         DP_OP_424J2_126_3477_n860, DP_OP_424J2_126_3477_n859,
         DP_OP_424J2_126_3477_n858, DP_OP_424J2_126_3477_n857,
         DP_OP_424J2_126_3477_n856, DP_OP_424J2_126_3477_n855,
         DP_OP_424J2_126_3477_n854, DP_OP_424J2_126_3477_n853,
         DP_OP_424J2_126_3477_n852, DP_OP_424J2_126_3477_n851,
         DP_OP_424J2_126_3477_n850, DP_OP_424J2_126_3477_n849,
         DP_OP_424J2_126_3477_n848, DP_OP_424J2_126_3477_n847,
         DP_OP_424J2_126_3477_n846, DP_OP_424J2_126_3477_n845,
         DP_OP_424J2_126_3477_n844, DP_OP_424J2_126_3477_n843,
         DP_OP_424J2_126_3477_n842, DP_OP_424J2_126_3477_n841,
         DP_OP_424J2_126_3477_n840, DP_OP_424J2_126_3477_n839,
         DP_OP_424J2_126_3477_n838, DP_OP_424J2_126_3477_n837,
         DP_OP_424J2_126_3477_n836, DP_OP_424J2_126_3477_n835,
         DP_OP_424J2_126_3477_n834, DP_OP_424J2_126_3477_n833,
         DP_OP_424J2_126_3477_n832, DP_OP_424J2_126_3477_n831,
         DP_OP_424J2_126_3477_n830, DP_OP_424J2_126_3477_n829,
         DP_OP_424J2_126_3477_n828, DP_OP_424J2_126_3477_n827,
         DP_OP_424J2_126_3477_n826, DP_OP_424J2_126_3477_n825,
         DP_OP_424J2_126_3477_n824, DP_OP_424J2_126_3477_n823,
         DP_OP_424J2_126_3477_n822, DP_OP_424J2_126_3477_n821,
         DP_OP_424J2_126_3477_n820, DP_OP_424J2_126_3477_n819,
         DP_OP_424J2_126_3477_n818, DP_OP_424J2_126_3477_n817,
         DP_OP_424J2_126_3477_n816, DP_OP_424J2_126_3477_n815,
         DP_OP_424J2_126_3477_n814, DP_OP_424J2_126_3477_n813,
         DP_OP_424J2_126_3477_n812, DP_OP_424J2_126_3477_n811,
         DP_OP_424J2_126_3477_n810, DP_OP_424J2_126_3477_n809,
         DP_OP_424J2_126_3477_n808, DP_OP_424J2_126_3477_n807,
         DP_OP_424J2_126_3477_n806, DP_OP_424J2_126_3477_n805,
         DP_OP_424J2_126_3477_n804, DP_OP_424J2_126_3477_n803,
         DP_OP_424J2_126_3477_n802, DP_OP_424J2_126_3477_n801,
         DP_OP_424J2_126_3477_n800, DP_OP_424J2_126_3477_n799,
         DP_OP_424J2_126_3477_n798, DP_OP_424J2_126_3477_n797,
         DP_OP_424J2_126_3477_n796, DP_OP_424J2_126_3477_n795,
         DP_OP_424J2_126_3477_n794, DP_OP_424J2_126_3477_n793,
         DP_OP_424J2_126_3477_n792, DP_OP_424J2_126_3477_n791,
         DP_OP_424J2_126_3477_n790, DP_OP_424J2_126_3477_n789,
         DP_OP_424J2_126_3477_n788, DP_OP_424J2_126_3477_n787,
         DP_OP_424J2_126_3477_n786, DP_OP_424J2_126_3477_n785,
         DP_OP_424J2_126_3477_n784, DP_OP_424J2_126_3477_n783,
         DP_OP_424J2_126_3477_n782, DP_OP_424J2_126_3477_n781,
         DP_OP_424J2_126_3477_n780, DP_OP_424J2_126_3477_n779,
         DP_OP_424J2_126_3477_n778, DP_OP_424J2_126_3477_n777,
         DP_OP_424J2_126_3477_n776, DP_OP_424J2_126_3477_n775,
         DP_OP_424J2_126_3477_n774, DP_OP_424J2_126_3477_n773,
         DP_OP_424J2_126_3477_n772, DP_OP_424J2_126_3477_n771,
         DP_OP_424J2_126_3477_n770, DP_OP_424J2_126_3477_n769,
         DP_OP_424J2_126_3477_n768, DP_OP_424J2_126_3477_n767,
         DP_OP_424J2_126_3477_n766, DP_OP_424J2_126_3477_n765,
         DP_OP_424J2_126_3477_n764, DP_OP_424J2_126_3477_n763,
         DP_OP_424J2_126_3477_n762, DP_OP_424J2_126_3477_n761,
         DP_OP_424J2_126_3477_n760, DP_OP_424J2_126_3477_n759,
         DP_OP_424J2_126_3477_n758, DP_OP_424J2_126_3477_n757,
         DP_OP_424J2_126_3477_n756, DP_OP_424J2_126_3477_n755,
         DP_OP_424J2_126_3477_n754, DP_OP_424J2_126_3477_n753,
         DP_OP_424J2_126_3477_n752, DP_OP_424J2_126_3477_n751,
         DP_OP_424J2_126_3477_n750, DP_OP_424J2_126_3477_n749,
         DP_OP_424J2_126_3477_n748, DP_OP_424J2_126_3477_n747,
         DP_OP_424J2_126_3477_n746, DP_OP_424J2_126_3477_n745,
         DP_OP_424J2_126_3477_n744, DP_OP_424J2_126_3477_n743,
         DP_OP_424J2_126_3477_n742, DP_OP_424J2_126_3477_n741,
         DP_OP_424J2_126_3477_n740, DP_OP_424J2_126_3477_n739,
         DP_OP_424J2_126_3477_n738, DP_OP_424J2_126_3477_n737,
         DP_OP_424J2_126_3477_n736, DP_OP_424J2_126_3477_n735,
         DP_OP_424J2_126_3477_n734, DP_OP_424J2_126_3477_n733,
         DP_OP_424J2_126_3477_n732, DP_OP_424J2_126_3477_n731,
         DP_OP_424J2_126_3477_n730, DP_OP_424J2_126_3477_n729,
         DP_OP_424J2_126_3477_n728, DP_OP_424J2_126_3477_n727,
         DP_OP_424J2_126_3477_n726, DP_OP_424J2_126_3477_n725,
         DP_OP_424J2_126_3477_n724, DP_OP_424J2_126_3477_n723,
         DP_OP_424J2_126_3477_n722, DP_OP_424J2_126_3477_n721,
         DP_OP_424J2_126_3477_n720, DP_OP_424J2_126_3477_n719,
         DP_OP_424J2_126_3477_n718, DP_OP_424J2_126_3477_n717,
         DP_OP_424J2_126_3477_n716, DP_OP_424J2_126_3477_n715,
         DP_OP_424J2_126_3477_n714, DP_OP_424J2_126_3477_n713,
         DP_OP_424J2_126_3477_n712, DP_OP_424J2_126_3477_n711,
         DP_OP_424J2_126_3477_n710, DP_OP_424J2_126_3477_n709,
         DP_OP_424J2_126_3477_n708, DP_OP_424J2_126_3477_n707,
         DP_OP_424J2_126_3477_n706, DP_OP_424J2_126_3477_n705,
         DP_OP_424J2_126_3477_n704, DP_OP_424J2_126_3477_n703,
         DP_OP_424J2_126_3477_n702, DP_OP_424J2_126_3477_n701,
         DP_OP_424J2_126_3477_n700, DP_OP_424J2_126_3477_n699,
         DP_OP_424J2_126_3477_n698, DP_OP_424J2_126_3477_n697,
         DP_OP_424J2_126_3477_n696, DP_OP_424J2_126_3477_n695,
         DP_OP_424J2_126_3477_n694, DP_OP_424J2_126_3477_n693,
         DP_OP_424J2_126_3477_n692, DP_OP_424J2_126_3477_n691,
         DP_OP_424J2_126_3477_n690, DP_OP_424J2_126_3477_n689,
         DP_OP_424J2_126_3477_n688, DP_OP_424J2_126_3477_n687,
         DP_OP_424J2_126_3477_n686, DP_OP_424J2_126_3477_n685,
         DP_OP_424J2_126_3477_n684, DP_OP_424J2_126_3477_n683,
         DP_OP_424J2_126_3477_n682, DP_OP_424J2_126_3477_n681,
         DP_OP_424J2_126_3477_n680, DP_OP_424J2_126_3477_n679,
         DP_OP_424J2_126_3477_n678, DP_OP_424J2_126_3477_n677,
         DP_OP_424J2_126_3477_n676, DP_OP_424J2_126_3477_n675,
         DP_OP_424J2_126_3477_n674, DP_OP_424J2_126_3477_n673,
         DP_OP_424J2_126_3477_n672, DP_OP_424J2_126_3477_n671,
         DP_OP_424J2_126_3477_n670, DP_OP_424J2_126_3477_n669,
         DP_OP_424J2_126_3477_n668, DP_OP_424J2_126_3477_n667,
         DP_OP_424J2_126_3477_n666, DP_OP_424J2_126_3477_n665,
         DP_OP_424J2_126_3477_n664, DP_OP_424J2_126_3477_n663,
         DP_OP_424J2_126_3477_n662, DP_OP_424J2_126_3477_n661,
         DP_OP_424J2_126_3477_n660, DP_OP_424J2_126_3477_n659,
         DP_OP_424J2_126_3477_n658, DP_OP_424J2_126_3477_n657,
         DP_OP_424J2_126_3477_n656, DP_OP_424J2_126_3477_n655,
         DP_OP_424J2_126_3477_n654, DP_OP_424J2_126_3477_n653,
         DP_OP_424J2_126_3477_n652, DP_OP_424J2_126_3477_n651,
         DP_OP_424J2_126_3477_n650, DP_OP_424J2_126_3477_n649,
         DP_OP_424J2_126_3477_n648, DP_OP_424J2_126_3477_n647,
         DP_OP_424J2_126_3477_n646, DP_OP_424J2_126_3477_n645,
         DP_OP_424J2_126_3477_n644, DP_OP_424J2_126_3477_n643,
         DP_OP_424J2_126_3477_n642, DP_OP_424J2_126_3477_n641,
         DP_OP_424J2_126_3477_n640, DP_OP_424J2_126_3477_n639,
         DP_OP_424J2_126_3477_n638, DP_OP_424J2_126_3477_n637,
         DP_OP_424J2_126_3477_n636, DP_OP_424J2_126_3477_n635,
         DP_OP_424J2_126_3477_n634, DP_OP_424J2_126_3477_n633,
         DP_OP_424J2_126_3477_n632, DP_OP_424J2_126_3477_n631,
         DP_OP_424J2_126_3477_n630, DP_OP_424J2_126_3477_n629,
         DP_OP_424J2_126_3477_n628, DP_OP_424J2_126_3477_n627,
         DP_OP_424J2_126_3477_n626, DP_OP_424J2_126_3477_n625,
         DP_OP_424J2_126_3477_n624, DP_OP_424J2_126_3477_n623,
         DP_OP_424J2_126_3477_n622, DP_OP_424J2_126_3477_n621,
         DP_OP_424J2_126_3477_n620, DP_OP_424J2_126_3477_n619,
         DP_OP_424J2_126_3477_n618, DP_OP_424J2_126_3477_n617,
         DP_OP_424J2_126_3477_n616, DP_OP_424J2_126_3477_n615,
         DP_OP_424J2_126_3477_n614, DP_OP_424J2_126_3477_n613,
         DP_OP_424J2_126_3477_n612, DP_OP_424J2_126_3477_n611,
         DP_OP_424J2_126_3477_n610, DP_OP_424J2_126_3477_n609,
         DP_OP_424J2_126_3477_n608, DP_OP_424J2_126_3477_n607,
         DP_OP_424J2_126_3477_n606, DP_OP_424J2_126_3477_n605,
         DP_OP_424J2_126_3477_n604, DP_OP_424J2_126_3477_n603,
         DP_OP_424J2_126_3477_n602, DP_OP_424J2_126_3477_n601,
         DP_OP_424J2_126_3477_n600, DP_OP_424J2_126_3477_n599,
         DP_OP_424J2_126_3477_n598, DP_OP_424J2_126_3477_n597,
         DP_OP_424J2_126_3477_n596, DP_OP_424J2_126_3477_n595,
         DP_OP_424J2_126_3477_n594, DP_OP_424J2_126_3477_n593,
         DP_OP_424J2_126_3477_n592, DP_OP_424J2_126_3477_n591,
         DP_OP_424J2_126_3477_n590, DP_OP_424J2_126_3477_n589,
         DP_OP_424J2_126_3477_n588, DP_OP_424J2_126_3477_n587,
         DP_OP_424J2_126_3477_n586, DP_OP_424J2_126_3477_n585,
         DP_OP_424J2_126_3477_n584, DP_OP_424J2_126_3477_n583,
         DP_OP_424J2_126_3477_n582, DP_OP_424J2_126_3477_n581,
         DP_OP_424J2_126_3477_n580, DP_OP_424J2_126_3477_n579,
         DP_OP_424J2_126_3477_n578, DP_OP_424J2_126_3477_n577,
         DP_OP_424J2_126_3477_n576, DP_OP_424J2_126_3477_n575,
         DP_OP_424J2_126_3477_n574, DP_OP_424J2_126_3477_n573,
         DP_OP_424J2_126_3477_n572, DP_OP_424J2_126_3477_n571,
         DP_OP_424J2_126_3477_n570, DP_OP_424J2_126_3477_n569,
         DP_OP_424J2_126_3477_n568, DP_OP_424J2_126_3477_n567,
         DP_OP_424J2_126_3477_n566, DP_OP_424J2_126_3477_n565,
         DP_OP_424J2_126_3477_n564, DP_OP_424J2_126_3477_n563,
         DP_OP_424J2_126_3477_n562, DP_OP_424J2_126_3477_n561,
         DP_OP_424J2_126_3477_n560, DP_OP_424J2_126_3477_n559,
         DP_OP_424J2_126_3477_n558, DP_OP_424J2_126_3477_n557,
         DP_OP_424J2_126_3477_n556, DP_OP_424J2_126_3477_n555,
         DP_OP_424J2_126_3477_n554, DP_OP_424J2_126_3477_n553,
         DP_OP_424J2_126_3477_n552, DP_OP_424J2_126_3477_n551,
         DP_OP_424J2_126_3477_n550, DP_OP_424J2_126_3477_n549,
         DP_OP_424J2_126_3477_n548, DP_OP_424J2_126_3477_n547,
         DP_OP_424J2_126_3477_n546, DP_OP_424J2_126_3477_n545,
         DP_OP_424J2_126_3477_n544, DP_OP_424J2_126_3477_n543,
         DP_OP_424J2_126_3477_n542, DP_OP_424J2_126_3477_n541,
         DP_OP_424J2_126_3477_n540, DP_OP_424J2_126_3477_n539,
         DP_OP_424J2_126_3477_n538, DP_OP_424J2_126_3477_n537,
         DP_OP_424J2_126_3477_n536, DP_OP_424J2_126_3477_n535,
         DP_OP_424J2_126_3477_n534, DP_OP_424J2_126_3477_n533,
         DP_OP_424J2_126_3477_n532, DP_OP_424J2_126_3477_n531,
         DP_OP_424J2_126_3477_n530, DP_OP_424J2_126_3477_n529,
         DP_OP_424J2_126_3477_n528, DP_OP_424J2_126_3477_n527,
         DP_OP_424J2_126_3477_n526, DP_OP_424J2_126_3477_n525,
         DP_OP_424J2_126_3477_n524, DP_OP_424J2_126_3477_n523,
         DP_OP_424J2_126_3477_n522, DP_OP_424J2_126_3477_n521,
         DP_OP_424J2_126_3477_n520, DP_OP_424J2_126_3477_n519,
         DP_OP_424J2_126_3477_n518, DP_OP_424J2_126_3477_n517,
         DP_OP_424J2_126_3477_n516, DP_OP_424J2_126_3477_n515,
         DP_OP_424J2_126_3477_n514, DP_OP_424J2_126_3477_n513,
         DP_OP_424J2_126_3477_n512, DP_OP_424J2_126_3477_n511,
         DP_OP_424J2_126_3477_n510, DP_OP_424J2_126_3477_n509,
         DP_OP_424J2_126_3477_n508, DP_OP_424J2_126_3477_n507,
         DP_OP_424J2_126_3477_n506, DP_OP_424J2_126_3477_n505,
         DP_OP_424J2_126_3477_n504, DP_OP_424J2_126_3477_n503,
         DP_OP_424J2_126_3477_n502, DP_OP_424J2_126_3477_n501,
         DP_OP_424J2_126_3477_n500, DP_OP_424J2_126_3477_n499,
         DP_OP_424J2_126_3477_n498, DP_OP_424J2_126_3477_n497,
         DP_OP_424J2_126_3477_n496, DP_OP_424J2_126_3477_n495,
         DP_OP_424J2_126_3477_n494, DP_OP_424J2_126_3477_n493,
         DP_OP_424J2_126_3477_n492, DP_OP_424J2_126_3477_n491,
         DP_OP_424J2_126_3477_n490, DP_OP_424J2_126_3477_n489,
         DP_OP_424J2_126_3477_n488, DP_OP_424J2_126_3477_n487,
         DP_OP_424J2_126_3477_n486, DP_OP_424J2_126_3477_n485,
         DP_OP_424J2_126_3477_n484, DP_OP_424J2_126_3477_n483,
         DP_OP_424J2_126_3477_n482, DP_OP_424J2_126_3477_n481,
         DP_OP_424J2_126_3477_n480, DP_OP_424J2_126_3477_n479,
         DP_OP_424J2_126_3477_n478, DP_OP_424J2_126_3477_n477,
         DP_OP_424J2_126_3477_n476, DP_OP_424J2_126_3477_n475,
         DP_OP_424J2_126_3477_n474, DP_OP_424J2_126_3477_n473,
         DP_OP_424J2_126_3477_n472, DP_OP_424J2_126_3477_n471,
         DP_OP_424J2_126_3477_n470, DP_OP_424J2_126_3477_n469,
         DP_OP_424J2_126_3477_n468, DP_OP_424J2_126_3477_n467,
         DP_OP_424J2_126_3477_n466, DP_OP_424J2_126_3477_n465,
         DP_OP_424J2_126_3477_n464, DP_OP_424J2_126_3477_n463,
         DP_OP_424J2_126_3477_n462, DP_OP_424J2_126_3477_n461,
         DP_OP_424J2_126_3477_n460, DP_OP_424J2_126_3477_n459,
         DP_OP_424J2_126_3477_n458, DP_OP_424J2_126_3477_n457,
         DP_OP_424J2_126_3477_n456, DP_OP_424J2_126_3477_n455,
         DP_OP_424J2_126_3477_n454, DP_OP_424J2_126_3477_n453,
         DP_OP_424J2_126_3477_n452, DP_OP_424J2_126_3477_n451,
         DP_OP_424J2_126_3477_n450, DP_OP_424J2_126_3477_n449,
         DP_OP_424J2_126_3477_n448, DP_OP_424J2_126_3477_n447,
         DP_OP_424J2_126_3477_n446, DP_OP_424J2_126_3477_n445,
         DP_OP_424J2_126_3477_n444, DP_OP_424J2_126_3477_n443,
         DP_OP_424J2_126_3477_n442, DP_OP_424J2_126_3477_n441,
         DP_OP_424J2_126_3477_n440, DP_OP_424J2_126_3477_n439,
         DP_OP_424J2_126_3477_n438, DP_OP_424J2_126_3477_n437,
         DP_OP_424J2_126_3477_n436, DP_OP_424J2_126_3477_n435,
         DP_OP_424J2_126_3477_n434, DP_OP_424J2_126_3477_n433,
         DP_OP_424J2_126_3477_n432, DP_OP_424J2_126_3477_n431,
         DP_OP_424J2_126_3477_n430, DP_OP_424J2_126_3477_n429,
         DP_OP_424J2_126_3477_n428, DP_OP_424J2_126_3477_n427,
         DP_OP_424J2_126_3477_n426, DP_OP_424J2_126_3477_n425,
         DP_OP_424J2_126_3477_n424, DP_OP_424J2_126_3477_n423,
         DP_OP_424J2_126_3477_n422, DP_OP_424J2_126_3477_n421,
         DP_OP_424J2_126_3477_n420, DP_OP_424J2_126_3477_n419,
         DP_OP_424J2_126_3477_n418, DP_OP_424J2_126_3477_n417,
         DP_OP_424J2_126_3477_n416, DP_OP_424J2_126_3477_n415,
         DP_OP_424J2_126_3477_n414, DP_OP_424J2_126_3477_n413,
         DP_OP_424J2_126_3477_n412, DP_OP_424J2_126_3477_n411,
         DP_OP_424J2_126_3477_n410, DP_OP_424J2_126_3477_n409,
         DP_OP_424J2_126_3477_n408, DP_OP_424J2_126_3477_n407,
         DP_OP_424J2_126_3477_n406, DP_OP_424J2_126_3477_n405,
         DP_OP_424J2_126_3477_n404, DP_OP_424J2_126_3477_n403,
         DP_OP_424J2_126_3477_n402, DP_OP_424J2_126_3477_n401,
         DP_OP_424J2_126_3477_n400, DP_OP_424J2_126_3477_n399,
         DP_OP_424J2_126_3477_n398, DP_OP_424J2_126_3477_n397,
         DP_OP_424J2_126_3477_n396, DP_OP_424J2_126_3477_n395,
         DP_OP_424J2_126_3477_n394, DP_OP_424J2_126_3477_n393,
         DP_OP_424J2_126_3477_n392, DP_OP_424J2_126_3477_n391,
         DP_OP_424J2_126_3477_n390, DP_OP_424J2_126_3477_n389,
         DP_OP_424J2_126_3477_n388, DP_OP_424J2_126_3477_n387,
         DP_OP_424J2_126_3477_n386, DP_OP_424J2_126_3477_n385,
         DP_OP_424J2_126_3477_n384, DP_OP_424J2_126_3477_n383,
         DP_OP_424J2_126_3477_n382, DP_OP_424J2_126_3477_n381,
         DP_OP_424J2_126_3477_n380, DP_OP_424J2_126_3477_n379,
         DP_OP_424J2_126_3477_n378, DP_OP_424J2_126_3477_n377,
         DP_OP_424J2_126_3477_n376, DP_OP_424J2_126_3477_n375,
         DP_OP_424J2_126_3477_n374, DP_OP_424J2_126_3477_n373,
         DP_OP_424J2_126_3477_n372, DP_OP_424J2_126_3477_n371,
         DP_OP_424J2_126_3477_n370, DP_OP_424J2_126_3477_n369,
         DP_OP_424J2_126_3477_n368, DP_OP_424J2_126_3477_n367,
         DP_OP_424J2_126_3477_n366, DP_OP_424J2_126_3477_n365,
         DP_OP_424J2_126_3477_n364, DP_OP_424J2_126_3477_n363,
         DP_OP_424J2_126_3477_n362, DP_OP_424J2_126_3477_n361,
         DP_OP_424J2_126_3477_n360, DP_OP_424J2_126_3477_n359,
         DP_OP_424J2_126_3477_n358, DP_OP_424J2_126_3477_n357,
         DP_OP_424J2_126_3477_n356, DP_OP_424J2_126_3477_n355,
         DP_OP_424J2_126_3477_n354, DP_OP_424J2_126_3477_n353,
         DP_OP_424J2_126_3477_n352, DP_OP_424J2_126_3477_n351,
         DP_OP_424J2_126_3477_n350, DP_OP_424J2_126_3477_n349,
         DP_OP_424J2_126_3477_n348, DP_OP_424J2_126_3477_n347,
         DP_OP_424J2_126_3477_n346, DP_OP_424J2_126_3477_n345,
         DP_OP_424J2_126_3477_n344, DP_OP_424J2_126_3477_n343,
         DP_OP_424J2_126_3477_n342, DP_OP_424J2_126_3477_n341,
         DP_OP_424J2_126_3477_n340, DP_OP_424J2_126_3477_n339,
         DP_OP_424J2_126_3477_n338, DP_OP_424J2_126_3477_n337,
         DP_OP_424J2_126_3477_n336, DP_OP_424J2_126_3477_n335,
         DP_OP_424J2_126_3477_n334, DP_OP_424J2_126_3477_n333,
         DP_OP_424J2_126_3477_n332, DP_OP_424J2_126_3477_n331,
         DP_OP_424J2_126_3477_n330, DP_OP_424J2_126_3477_n329,
         DP_OP_424J2_126_3477_n328, DP_OP_424J2_126_3477_n327,
         DP_OP_424J2_126_3477_n326, DP_OP_424J2_126_3477_n325,
         DP_OP_424J2_126_3477_n324, DP_OP_424J2_126_3477_n323,
         DP_OP_424J2_126_3477_n322, DP_OP_424J2_126_3477_n321,
         DP_OP_424J2_126_3477_n320, DP_OP_424J2_126_3477_n319,
         DP_OP_424J2_126_3477_n318, DP_OP_424J2_126_3477_n317,
         DP_OP_424J2_126_3477_n316, DP_OP_424J2_126_3477_n315,
         DP_OP_424J2_126_3477_n314, DP_OP_424J2_126_3477_n313,
         DP_OP_424J2_126_3477_n312, DP_OP_424J2_126_3477_n311,
         DP_OP_424J2_126_3477_n310, DP_OP_424J2_126_3477_n309,
         DP_OP_424J2_126_3477_n308, DP_OP_424J2_126_3477_n307,
         DP_OP_424J2_126_3477_n306, DP_OP_424J2_126_3477_n305,
         DP_OP_424J2_126_3477_n304, DP_OP_424J2_126_3477_n303,
         DP_OP_424J2_126_3477_n302, DP_OP_424J2_126_3477_n301,
         DP_OP_424J2_126_3477_n300, DP_OP_424J2_126_3477_n299,
         DP_OP_424J2_126_3477_n298, DP_OP_424J2_126_3477_n297,
         DP_OP_424J2_126_3477_n296, DP_OP_424J2_126_3477_n295,
         DP_OP_424J2_126_3477_n294, DP_OP_424J2_126_3477_n293,
         DP_OP_424J2_126_3477_n292, DP_OP_424J2_126_3477_n291,
         DP_OP_424J2_126_3477_n290, DP_OP_424J2_126_3477_n289,
         DP_OP_424J2_126_3477_n288, DP_OP_424J2_126_3477_n287,
         DP_OP_424J2_126_3477_n286, DP_OP_424J2_126_3477_n285,
         DP_OP_424J2_126_3477_n284, DP_OP_424J2_126_3477_n283,
         DP_OP_424J2_126_3477_n282, DP_OP_424J2_126_3477_n281,
         DP_OP_424J2_126_3477_n280, DP_OP_424J2_126_3477_n279,
         DP_OP_424J2_126_3477_n278, DP_OP_424J2_126_3477_n277,
         DP_OP_424J2_126_3477_n276, DP_OP_424J2_126_3477_n275,
         DP_OP_424J2_126_3477_n274, DP_OP_424J2_126_3477_n273,
         DP_OP_424J2_126_3477_n272, DP_OP_424J2_126_3477_n271,
         DP_OP_424J2_126_3477_n270, DP_OP_424J2_126_3477_n269,
         DP_OP_424J2_126_3477_n268, DP_OP_424J2_126_3477_n267,
         DP_OP_424J2_126_3477_n266, DP_OP_424J2_126_3477_n265,
         DP_OP_424J2_126_3477_n264, DP_OP_424J2_126_3477_n263,
         DP_OP_424J2_126_3477_n262, DP_OP_424J2_126_3477_n261,
         DP_OP_424J2_126_3477_n260, DP_OP_424J2_126_3477_n259,
         DP_OP_424J2_126_3477_n258, DP_OP_424J2_126_3477_n257,
         DP_OP_424J2_126_3477_n256, DP_OP_424J2_126_3477_n255,
         DP_OP_424J2_126_3477_n254, DP_OP_424J2_126_3477_n253,
         DP_OP_424J2_126_3477_n252, DP_OP_424J2_126_3477_n251,
         DP_OP_424J2_126_3477_n250, DP_OP_424J2_126_3477_n249,
         DP_OP_424J2_126_3477_n248, DP_OP_424J2_126_3477_n247,
         DP_OP_424J2_126_3477_n246, DP_OP_424J2_126_3477_n245,
         DP_OP_424J2_126_3477_n244, DP_OP_424J2_126_3477_n243,
         DP_OP_424J2_126_3477_n242, DP_OP_424J2_126_3477_n241,
         DP_OP_424J2_126_3477_n240, DP_OP_424J2_126_3477_n239,
         DP_OP_424J2_126_3477_n238, DP_OP_424J2_126_3477_n237,
         DP_OP_424J2_126_3477_n236, DP_OP_424J2_126_3477_n235,
         DP_OP_424J2_126_3477_n234, DP_OP_424J2_126_3477_n233,
         DP_OP_424J2_126_3477_n232, DP_OP_424J2_126_3477_n231,
         DP_OP_424J2_126_3477_n230, DP_OP_424J2_126_3477_n229,
         DP_OP_424J2_126_3477_n228, DP_OP_424J2_126_3477_n227,
         DP_OP_424J2_126_3477_n226, DP_OP_424J2_126_3477_n225,
         DP_OP_424J2_126_3477_n224, DP_OP_424J2_126_3477_n223,
         DP_OP_424J2_126_3477_n222, DP_OP_424J2_126_3477_n221,
         DP_OP_424J2_126_3477_n220, DP_OP_424J2_126_3477_n219,
         DP_OP_424J2_126_3477_n218, DP_OP_424J2_126_3477_n217,
         DP_OP_424J2_126_3477_n216, DP_OP_424J2_126_3477_n215,
         DP_OP_424J2_126_3477_n214, DP_OP_424J2_126_3477_n213,
         DP_OP_424J2_126_3477_n212, DP_OP_424J2_126_3477_n211,
         DP_OP_424J2_126_3477_n210, DP_OP_424J2_126_3477_n209,
         DP_OP_424J2_126_3477_n208, DP_OP_424J2_126_3477_n207,
         DP_OP_424J2_126_3477_n206, DP_OP_424J2_126_3477_n205,
         DP_OP_424J2_126_3477_n204, DP_OP_424J2_126_3477_n203,
         DP_OP_424J2_126_3477_n202, DP_OP_424J2_126_3477_n201,
         DP_OP_424J2_126_3477_n200, DP_OP_424J2_126_3477_n199,
         DP_OP_424J2_126_3477_n198, DP_OP_424J2_126_3477_n197,
         DP_OP_424J2_126_3477_n196, DP_OP_424J2_126_3477_n195,
         DP_OP_424J2_126_3477_n194, DP_OP_424J2_126_3477_n193,
         DP_OP_424J2_126_3477_n192, DP_OP_424J2_126_3477_n191,
         DP_OP_424J2_126_3477_n190, DP_OP_424J2_126_3477_n189,
         DP_OP_424J2_126_3477_n188, DP_OP_424J2_126_3477_n187,
         DP_OP_424J2_126_3477_n186, DP_OP_424J2_126_3477_n185,
         DP_OP_424J2_126_3477_n184, DP_OP_424J2_126_3477_n183,
         DP_OP_424J2_126_3477_n182, DP_OP_424J2_126_3477_n181,
         DP_OP_424J2_126_3477_n180, DP_OP_424J2_126_3477_n179,
         DP_OP_424J2_126_3477_n178, DP_OP_424J2_126_3477_n177,
         DP_OP_424J2_126_3477_n176, DP_OP_424J2_126_3477_n175,
         DP_OP_424J2_126_3477_n174, DP_OP_424J2_126_3477_n173,
         DP_OP_424J2_126_3477_n172, DP_OP_424J2_126_3477_n171,
         DP_OP_424J2_126_3477_n170, DP_OP_424J2_126_3477_n169,
         DP_OP_424J2_126_3477_n168, DP_OP_424J2_126_3477_n167,
         DP_OP_424J2_126_3477_n166, DP_OP_424J2_126_3477_n165,
         DP_OP_424J2_126_3477_n164, DP_OP_424J2_126_3477_n163,
         DP_OP_424J2_126_3477_n162, DP_OP_424J2_126_3477_n161,
         DP_OP_424J2_126_3477_n160, DP_OP_424J2_126_3477_n159,
         DP_OP_424J2_126_3477_n158, DP_OP_424J2_126_3477_n157,
         DP_OP_424J2_126_3477_n156, DP_OP_424J2_126_3477_n155,
         DP_OP_424J2_126_3477_n154, DP_OP_424J2_126_3477_n153,
         DP_OP_424J2_126_3477_n131, DP_OP_424J2_126_3477_n130,
         DP_OP_424J2_126_3477_n129, DP_OP_424J2_126_3477_n128,
         DP_OP_424J2_126_3477_n127, DP_OP_424J2_126_3477_n126,
         DP_OP_424J2_126_3477_n123, DP_OP_424J2_126_3477_n122,
         DP_OP_424J2_126_3477_n121, DP_OP_424J2_126_3477_n120,
         DP_OP_424J2_126_3477_n119, DP_OP_424J2_126_3477_n118,
         DP_OP_424J2_126_3477_n115, DP_OP_424J2_126_3477_n114,
         DP_OP_424J2_126_3477_n113, DP_OP_424J2_126_3477_n112,
         DP_OP_424J2_126_3477_n111, DP_OP_424J2_126_3477_n110,
         DP_OP_424J2_126_3477_n107, DP_OP_424J2_126_3477_n106,
         DP_OP_424J2_126_3477_n105, DP_OP_424J2_126_3477_n104,
         DP_OP_424J2_126_3477_n103, DP_OP_424J2_126_3477_n102,
         DP_OP_424J2_126_3477_n101, DP_OP_424J2_126_3477_n99,
         DP_OP_424J2_126_3477_n98, DP_OP_424J2_126_3477_n95,
         DP_OP_424J2_126_3477_n94, DP_OP_424J2_126_3477_n93,
         DP_OP_424J2_126_3477_n92, DP_OP_424J2_126_3477_n90,
         DP_OP_424J2_126_3477_n88, DP_OP_424J2_126_3477_n87,
         DP_OP_424J2_126_3477_n86, DP_OP_424J2_126_3477_n85,
         DP_OP_424J2_126_3477_n84, DP_OP_424J2_126_3477_n83,
         DP_OP_424J2_126_3477_n82, DP_OP_424J2_126_3477_n80,
         DP_OP_424J2_126_3477_n79, DP_OP_424J2_126_3477_n78,
         DP_OP_424J2_126_3477_n77, DP_OP_424J2_126_3477_n76,
         DP_OP_424J2_126_3477_n75, DP_OP_424J2_126_3477_n74,
         DP_OP_424J2_126_3477_n73, DP_OP_424J2_126_3477_n69,
         DP_OP_424J2_126_3477_n68, DP_OP_424J2_126_3477_n67,
         DP_OP_424J2_126_3477_n66, DP_OP_424J2_126_3477_n65,
         DP_OP_424J2_126_3477_n64, DP_OP_424J2_126_3477_n62,
         DP_OP_424J2_126_3477_n60, DP_OP_424J2_126_3477_n59,
         DP_OP_424J2_126_3477_n57, DP_OP_424J2_126_3477_n56,
         DP_OP_424J2_126_3477_n55, DP_OP_424J2_126_3477_n53,
         DP_OP_424J2_126_3477_n52, DP_OP_424J2_126_3477_n51,
         DP_OP_424J2_126_3477_n50, DP_OP_424J2_126_3477_n46,
         DP_OP_424J2_126_3477_n45, DP_OP_424J2_126_3477_n42,
         DP_OP_424J2_126_3477_n41, DP_OP_424J2_126_3477_n39,
         DP_OP_424J2_126_3477_n38, DP_OP_424J2_126_3477_n37,
         DP_OP_424J2_126_3477_n36, DP_OP_424J2_126_3477_n35,
         DP_OP_424J2_126_3477_n34, DP_OP_424J2_126_3477_n33,
         DP_OP_424J2_126_3477_n32, DP_OP_424J2_126_3477_n31,
         DP_OP_424J2_126_3477_n30, DP_OP_424J2_126_3477_n29,
         DP_OP_424J2_126_3477_n28, DP_OP_424J2_126_3477_n27,
         DP_OP_424J2_126_3477_n26, DP_OP_424J2_126_3477_n25,
         DP_OP_424J2_126_3477_n24, DP_OP_424J2_126_3477_n4,
         DP_OP_424J2_126_3477_n3, DP_OP_424J2_126_3477_n2,
         DP_OP_422J2_124_3477_n2918, DP_OP_422J2_124_3477_n2917,
         DP_OP_422J2_124_3477_n2916, DP_OP_422J2_124_3477_n2913,
         DP_OP_422J2_124_3477_n2912, DP_OP_422J2_124_3477_n2909,
         DP_OP_422J2_124_3477_n2908, DP_OP_422J2_124_3477_n2906,
         DP_OP_422J2_124_3477_n2905, DP_OP_422J2_124_3477_n2904,
         DP_OP_422J2_124_3477_n2903, DP_OP_422J2_124_3477_n2902,
         DP_OP_422J2_124_3477_n2901, DP_OP_422J2_124_3477_n2900,
         DP_OP_422J2_124_3477_n2899, DP_OP_422J2_124_3477_n2898,
         DP_OP_422J2_124_3477_n2897, DP_OP_422J2_124_3477_n2896,
         DP_OP_422J2_124_3477_n2895, DP_OP_422J2_124_3477_n2894,
         DP_OP_422J2_124_3477_n2893, DP_OP_422J2_124_3477_n2892,
         DP_OP_422J2_124_3477_n2891, DP_OP_422J2_124_3477_n2890,
         DP_OP_422J2_124_3477_n2889, DP_OP_422J2_124_3477_n2888,
         DP_OP_422J2_124_3477_n2887, DP_OP_422J2_124_3477_n2886,
         DP_OP_422J2_124_3477_n2885, DP_OP_422J2_124_3477_n2884,
         DP_OP_422J2_124_3477_n2883, DP_OP_422J2_124_3477_n2882,
         DP_OP_422J2_124_3477_n2881, DP_OP_422J2_124_3477_n2880,
         DP_OP_422J2_124_3477_n2879, DP_OP_422J2_124_3477_n2878,
         DP_OP_422J2_124_3477_n2877, DP_OP_422J2_124_3477_n2876,
         DP_OP_422J2_124_3477_n2875, DP_OP_422J2_124_3477_n2873,
         DP_OP_422J2_124_3477_n2872, DP_OP_422J2_124_3477_n2871,
         DP_OP_422J2_124_3477_n2870, DP_OP_422J2_124_3477_n2869,
         DP_OP_422J2_124_3477_n2868, DP_OP_422J2_124_3477_n2865,
         DP_OP_422J2_124_3477_n2864, DP_OP_422J2_124_3477_n2862,
         DP_OP_422J2_124_3477_n2861, DP_OP_422J2_124_3477_n2860,
         DP_OP_422J2_124_3477_n2859, DP_OP_422J2_124_3477_n2858,
         DP_OP_422J2_124_3477_n2857, DP_OP_422J2_124_3477_n2856,
         DP_OP_422J2_124_3477_n2855, DP_OP_422J2_124_3477_n2854,
         DP_OP_422J2_124_3477_n2853, DP_OP_422J2_124_3477_n2852,
         DP_OP_422J2_124_3477_n2851, DP_OP_422J2_124_3477_n2850,
         DP_OP_422J2_124_3477_n2849, DP_OP_422J2_124_3477_n2848,
         DP_OP_422J2_124_3477_n2847, DP_OP_422J2_124_3477_n2846,
         DP_OP_422J2_124_3477_n2845, DP_OP_422J2_124_3477_n2844,
         DP_OP_422J2_124_3477_n2843, DP_OP_422J2_124_3477_n2842,
         DP_OP_422J2_124_3477_n2841, DP_OP_422J2_124_3477_n2840,
         DP_OP_422J2_124_3477_n2839, DP_OP_422J2_124_3477_n2838,
         DP_OP_422J2_124_3477_n2837, DP_OP_422J2_124_3477_n2836,
         DP_OP_422J2_124_3477_n2835, DP_OP_422J2_124_3477_n2834,
         DP_OP_422J2_124_3477_n2833, DP_OP_422J2_124_3477_n2832,
         DP_OP_422J2_124_3477_n2831, DP_OP_422J2_124_3477_n2830,
         DP_OP_422J2_124_3477_n2827, DP_OP_422J2_124_3477_n2825,
         DP_OP_422J2_124_3477_n2820, DP_OP_422J2_124_3477_n2819,
         DP_OP_422J2_124_3477_n2818, DP_OP_422J2_124_3477_n2817,
         DP_OP_422J2_124_3477_n2816, DP_OP_422J2_124_3477_n2815,
         DP_OP_422J2_124_3477_n2814, DP_OP_422J2_124_3477_n2813,
         DP_OP_422J2_124_3477_n2812, DP_OP_422J2_124_3477_n2811,
         DP_OP_422J2_124_3477_n2810, DP_OP_422J2_124_3477_n2809,
         DP_OP_422J2_124_3477_n2808, DP_OP_422J2_124_3477_n2807,
         DP_OP_422J2_124_3477_n2806, DP_OP_422J2_124_3477_n2805,
         DP_OP_422J2_124_3477_n2804, DP_OP_422J2_124_3477_n2803,
         DP_OP_422J2_124_3477_n2802, DP_OP_422J2_124_3477_n2801,
         DP_OP_422J2_124_3477_n2800, DP_OP_422J2_124_3477_n2799,
         DP_OP_422J2_124_3477_n2798, DP_OP_422J2_124_3477_n2797,
         DP_OP_422J2_124_3477_n2796, DP_OP_422J2_124_3477_n2795,
         DP_OP_422J2_124_3477_n2794, DP_OP_422J2_124_3477_n2793,
         DP_OP_422J2_124_3477_n2792, DP_OP_422J2_124_3477_n2791,
         DP_OP_422J2_124_3477_n2790, DP_OP_422J2_124_3477_n2789,
         DP_OP_422J2_124_3477_n2788, DP_OP_422J2_124_3477_n2787,
         DP_OP_422J2_124_3477_n2786, DP_OP_422J2_124_3477_n2785,
         DP_OP_422J2_124_3477_n2784, DP_OP_422J2_124_3477_n2782,
         DP_OP_422J2_124_3477_n2781, DP_OP_422J2_124_3477_n2780,
         DP_OP_422J2_124_3477_n2777, DP_OP_422J2_124_3477_n2776,
         DP_OP_422J2_124_3477_n2774, DP_OP_422J2_124_3477_n2773,
         DP_OP_422J2_124_3477_n2772, DP_OP_422J2_124_3477_n2771,
         DP_OP_422J2_124_3477_n2770, DP_OP_422J2_124_3477_n2769,
         DP_OP_422J2_124_3477_n2768, DP_OP_422J2_124_3477_n2767,
         DP_OP_422J2_124_3477_n2766, DP_OP_422J2_124_3477_n2765,
         DP_OP_422J2_124_3477_n2764, DP_OP_422J2_124_3477_n2763,
         DP_OP_422J2_124_3477_n2762, DP_OP_422J2_124_3477_n2761,
         DP_OP_422J2_124_3477_n2760, DP_OP_422J2_124_3477_n2759,
         DP_OP_422J2_124_3477_n2758, DP_OP_422J2_124_3477_n2757,
         DP_OP_422J2_124_3477_n2756, DP_OP_422J2_124_3477_n2755,
         DP_OP_422J2_124_3477_n2754, DP_OP_422J2_124_3477_n2753,
         DP_OP_422J2_124_3477_n2752, DP_OP_422J2_124_3477_n2751,
         DP_OP_422J2_124_3477_n2750, DP_OP_422J2_124_3477_n2749,
         DP_OP_422J2_124_3477_n2748, DP_OP_422J2_124_3477_n2747,
         DP_OP_422J2_124_3477_n2746, DP_OP_422J2_124_3477_n2745,
         DP_OP_422J2_124_3477_n2744, DP_OP_422J2_124_3477_n2743,
         DP_OP_422J2_124_3477_n2742, DP_OP_422J2_124_3477_n2741,
         DP_OP_422J2_124_3477_n2740, DP_OP_422J2_124_3477_n2739,
         DP_OP_422J2_124_3477_n2736, DP_OP_422J2_124_3477_n2735,
         DP_OP_422J2_124_3477_n2734, DP_OP_422J2_124_3477_n2733,
         DP_OP_422J2_124_3477_n2732, DP_OP_422J2_124_3477_n2731,
         DP_OP_422J2_124_3477_n2730, DP_OP_422J2_124_3477_n2729,
         DP_OP_422J2_124_3477_n2728, DP_OP_422J2_124_3477_n2727,
         DP_OP_422J2_124_3477_n2726, DP_OP_422J2_124_3477_n2725,
         DP_OP_422J2_124_3477_n2724, DP_OP_422J2_124_3477_n2723,
         DP_OP_422J2_124_3477_n2722, DP_OP_422J2_124_3477_n2721,
         DP_OP_422J2_124_3477_n2720, DP_OP_422J2_124_3477_n2719,
         DP_OP_422J2_124_3477_n2718, DP_OP_422J2_124_3477_n2717,
         DP_OP_422J2_124_3477_n2716, DP_OP_422J2_124_3477_n2715,
         DP_OP_422J2_124_3477_n2714, DP_OP_422J2_124_3477_n2713,
         DP_OP_422J2_124_3477_n2712, DP_OP_422J2_124_3477_n2711,
         DP_OP_422J2_124_3477_n2710, DP_OP_422J2_124_3477_n2709,
         DP_OP_422J2_124_3477_n2708, DP_OP_422J2_124_3477_n2707,
         DP_OP_422J2_124_3477_n2706, DP_OP_422J2_124_3477_n2705,
         DP_OP_422J2_124_3477_n2704, DP_OP_422J2_124_3477_n2703,
         DP_OP_422J2_124_3477_n2702, DP_OP_422J2_124_3477_n2701,
         DP_OP_422J2_124_3477_n2700, DP_OP_422J2_124_3477_n2699,
         DP_OP_422J2_124_3477_n2698, DP_OP_422J2_124_3477_n2697,
         DP_OP_422J2_124_3477_n2696, DP_OP_422J2_124_3477_n2695,
         DP_OP_422J2_124_3477_n2694, DP_OP_422J2_124_3477_n2692,
         DP_OP_422J2_124_3477_n2690, DP_OP_422J2_124_3477_n2689,
         DP_OP_422J2_124_3477_n2688, DP_OP_422J2_124_3477_n2687,
         DP_OP_422J2_124_3477_n2686, DP_OP_422J2_124_3477_n2685,
         DP_OP_422J2_124_3477_n2684, DP_OP_422J2_124_3477_n2683,
         DP_OP_422J2_124_3477_n2682, DP_OP_422J2_124_3477_n2681,
         DP_OP_422J2_124_3477_n2680, DP_OP_422J2_124_3477_n2679,
         DP_OP_422J2_124_3477_n2678, DP_OP_422J2_124_3477_n2677,
         DP_OP_422J2_124_3477_n2676, DP_OP_422J2_124_3477_n2675,
         DP_OP_422J2_124_3477_n2674, DP_OP_422J2_124_3477_n2673,
         DP_OP_422J2_124_3477_n2672, DP_OP_422J2_124_3477_n2671,
         DP_OP_422J2_124_3477_n2670, DP_OP_422J2_124_3477_n2669,
         DP_OP_422J2_124_3477_n2668, DP_OP_422J2_124_3477_n2667,
         DP_OP_422J2_124_3477_n2666, DP_OP_422J2_124_3477_n2665,
         DP_OP_422J2_124_3477_n2664, DP_OP_422J2_124_3477_n2663,
         DP_OP_422J2_124_3477_n2662, DP_OP_422J2_124_3477_n2661,
         DP_OP_422J2_124_3477_n2660, DP_OP_422J2_124_3477_n2659,
         DP_OP_422J2_124_3477_n2658, DP_OP_422J2_124_3477_n2657,
         DP_OP_422J2_124_3477_n2656, DP_OP_422J2_124_3477_n2655,
         DP_OP_422J2_124_3477_n2654, DP_OP_422J2_124_3477_n2653,
         DP_OP_422J2_124_3477_n2652, DP_OP_422J2_124_3477_n2651,
         DP_OP_422J2_124_3477_n2650, DP_OP_422J2_124_3477_n2649,
         DP_OP_422J2_124_3477_n2648, DP_OP_422J2_124_3477_n2647,
         DP_OP_422J2_124_3477_n2646, DP_OP_422J2_124_3477_n2645,
         DP_OP_422J2_124_3477_n2644, DP_OP_422J2_124_3477_n2643,
         DP_OP_422J2_124_3477_n2642, DP_OP_422J2_124_3477_n2641,
         DP_OP_422J2_124_3477_n2640, DP_OP_422J2_124_3477_n2639,
         DP_OP_422J2_124_3477_n2638, DP_OP_422J2_124_3477_n2637,
         DP_OP_422J2_124_3477_n2636, DP_OP_422J2_124_3477_n2635,
         DP_OP_422J2_124_3477_n2634, DP_OP_422J2_124_3477_n2633,
         DP_OP_422J2_124_3477_n2632, DP_OP_422J2_124_3477_n2631,
         DP_OP_422J2_124_3477_n2630, DP_OP_422J2_124_3477_n2629,
         DP_OP_422J2_124_3477_n2628, DP_OP_422J2_124_3477_n2627,
         DP_OP_422J2_124_3477_n2626, DP_OP_422J2_124_3477_n2625,
         DP_OP_422J2_124_3477_n2624, DP_OP_422J2_124_3477_n2623,
         DP_OP_422J2_124_3477_n2622, DP_OP_422J2_124_3477_n2621,
         DP_OP_422J2_124_3477_n2620, DP_OP_422J2_124_3477_n2619,
         DP_OP_422J2_124_3477_n2618, DP_OP_422J2_124_3477_n2617,
         DP_OP_422J2_124_3477_n2616, DP_OP_422J2_124_3477_n2615,
         DP_OP_422J2_124_3477_n2614, DP_OP_422J2_124_3477_n2613,
         DP_OP_422J2_124_3477_n2612, DP_OP_422J2_124_3477_n2611,
         DP_OP_422J2_124_3477_n2610, DP_OP_422J2_124_3477_n2609,
         DP_OP_422J2_124_3477_n2608, DP_OP_422J2_124_3477_n2607,
         DP_OP_422J2_124_3477_n2606, DP_OP_422J2_124_3477_n2605,
         DP_OP_422J2_124_3477_n2604, DP_OP_422J2_124_3477_n2603,
         DP_OP_422J2_124_3477_n2602, DP_OP_422J2_124_3477_n2601,
         DP_OP_422J2_124_3477_n2600, DP_OP_422J2_124_3477_n2599,
         DP_OP_422J2_124_3477_n2598, DP_OP_422J2_124_3477_n2597,
         DP_OP_422J2_124_3477_n2596, DP_OP_422J2_124_3477_n2595,
         DP_OP_422J2_124_3477_n2594, DP_OP_422J2_124_3477_n2593,
         DP_OP_422J2_124_3477_n2592, DP_OP_422J2_124_3477_n2591,
         DP_OP_422J2_124_3477_n2590, DP_OP_422J2_124_3477_n2589,
         DP_OP_422J2_124_3477_n2588, DP_OP_422J2_124_3477_n2587,
         DP_OP_422J2_124_3477_n2586, DP_OP_422J2_124_3477_n2585,
         DP_OP_422J2_124_3477_n2584, DP_OP_422J2_124_3477_n2583,
         DP_OP_422J2_124_3477_n2582, DP_OP_422J2_124_3477_n2581,
         DP_OP_422J2_124_3477_n2580, DP_OP_422J2_124_3477_n2579,
         DP_OP_422J2_124_3477_n2578, DP_OP_422J2_124_3477_n2577,
         DP_OP_422J2_124_3477_n2576, DP_OP_422J2_124_3477_n2575,
         DP_OP_422J2_124_3477_n2574, DP_OP_422J2_124_3477_n2573,
         DP_OP_422J2_124_3477_n2572, DP_OP_422J2_124_3477_n2571,
         DP_OP_422J2_124_3477_n2570, DP_OP_422J2_124_3477_n2569,
         DP_OP_422J2_124_3477_n2568, DP_OP_422J2_124_3477_n2567,
         DP_OP_422J2_124_3477_n2566, DP_OP_422J2_124_3477_n2564,
         DP_OP_422J2_124_3477_n2563, DP_OP_422J2_124_3477_n2562,
         DP_OP_422J2_124_3477_n2560, DP_OP_422J2_124_3477_n2559,
         DP_OP_422J2_124_3477_n2558, DP_OP_422J2_124_3477_n2557,
         DP_OP_422J2_124_3477_n2556, DP_OP_422J2_124_3477_n2555,
         DP_OP_422J2_124_3477_n2554, DP_OP_422J2_124_3477_n2553,
         DP_OP_422J2_124_3477_n2552, DP_OP_422J2_124_3477_n2551,
         DP_OP_422J2_124_3477_n2550, DP_OP_422J2_124_3477_n2549,
         DP_OP_422J2_124_3477_n2548, DP_OP_422J2_124_3477_n2547,
         DP_OP_422J2_124_3477_n2546, DP_OP_422J2_124_3477_n2545,
         DP_OP_422J2_124_3477_n2544, DP_OP_422J2_124_3477_n2543,
         DP_OP_422J2_124_3477_n2542, DP_OP_422J2_124_3477_n2541,
         DP_OP_422J2_124_3477_n2540, DP_OP_422J2_124_3477_n2539,
         DP_OP_422J2_124_3477_n2538, DP_OP_422J2_124_3477_n2537,
         DP_OP_422J2_124_3477_n2536, DP_OP_422J2_124_3477_n2535,
         DP_OP_422J2_124_3477_n2534, DP_OP_422J2_124_3477_n2533,
         DP_OP_422J2_124_3477_n2532, DP_OP_422J2_124_3477_n2531,
         DP_OP_422J2_124_3477_n2530, DP_OP_422J2_124_3477_n2529,
         DP_OP_422J2_124_3477_n2528, DP_OP_422J2_124_3477_n2527,
         DP_OP_422J2_124_3477_n2526, DP_OP_422J2_124_3477_n2525,
         DP_OP_422J2_124_3477_n2524, DP_OP_422J2_124_3477_n2523,
         DP_OP_422J2_124_3477_n2522, DP_OP_422J2_124_3477_n2521,
         DP_OP_422J2_124_3477_n2520, DP_OP_422J2_124_3477_n2518,
         DP_OP_422J2_124_3477_n2514, DP_OP_422J2_124_3477_n2513,
         DP_OP_422J2_124_3477_n2512, DP_OP_422J2_124_3477_n2511,
         DP_OP_422J2_124_3477_n2510, DP_OP_422J2_124_3477_n2509,
         DP_OP_422J2_124_3477_n2508, DP_OP_422J2_124_3477_n2507,
         DP_OP_422J2_124_3477_n2506, DP_OP_422J2_124_3477_n2505,
         DP_OP_422J2_124_3477_n2504, DP_OP_422J2_124_3477_n2503,
         DP_OP_422J2_124_3477_n2502, DP_OP_422J2_124_3477_n2501,
         DP_OP_422J2_124_3477_n2500, DP_OP_422J2_124_3477_n2499,
         DP_OP_422J2_124_3477_n2498, DP_OP_422J2_124_3477_n2497,
         DP_OP_422J2_124_3477_n2496, DP_OP_422J2_124_3477_n2495,
         DP_OP_422J2_124_3477_n2494, DP_OP_422J2_124_3477_n2493,
         DP_OP_422J2_124_3477_n2492, DP_OP_422J2_124_3477_n2491,
         DP_OP_422J2_124_3477_n2490, DP_OP_422J2_124_3477_n2489,
         DP_OP_422J2_124_3477_n2488, DP_OP_422J2_124_3477_n2487,
         DP_OP_422J2_124_3477_n2486, DP_OP_422J2_124_3477_n2485,
         DP_OP_422J2_124_3477_n2484, DP_OP_422J2_124_3477_n2483,
         DP_OP_422J2_124_3477_n2482, DP_OP_422J2_124_3477_n2481,
         DP_OP_422J2_124_3477_n2480, DP_OP_422J2_124_3477_n2479,
         DP_OP_422J2_124_3477_n2478, DP_OP_422J2_124_3477_n2477,
         DP_OP_422J2_124_3477_n2476, DP_OP_422J2_124_3477_n2473,
         DP_OP_422J2_124_3477_n2472, DP_OP_422J2_124_3477_n2470,
         DP_OP_422J2_124_3477_n2469, DP_OP_422J2_124_3477_n2468,
         DP_OP_422J2_124_3477_n2467, DP_OP_422J2_124_3477_n2466,
         DP_OP_422J2_124_3477_n2465, DP_OP_422J2_124_3477_n2464,
         DP_OP_422J2_124_3477_n2463, DP_OP_422J2_124_3477_n2462,
         DP_OP_422J2_124_3477_n2461, DP_OP_422J2_124_3477_n2460,
         DP_OP_422J2_124_3477_n2459, DP_OP_422J2_124_3477_n2458,
         DP_OP_422J2_124_3477_n2457, DP_OP_422J2_124_3477_n2456,
         DP_OP_422J2_124_3477_n2455, DP_OP_422J2_124_3477_n2454,
         DP_OP_422J2_124_3477_n2453, DP_OP_422J2_124_3477_n2452,
         DP_OP_422J2_124_3477_n2451, DP_OP_422J2_124_3477_n2450,
         DP_OP_422J2_124_3477_n2449, DP_OP_422J2_124_3477_n2448,
         DP_OP_422J2_124_3477_n2447, DP_OP_422J2_124_3477_n2446,
         DP_OP_422J2_124_3477_n2445, DP_OP_422J2_124_3477_n2444,
         DP_OP_422J2_124_3477_n2443, DP_OP_422J2_124_3477_n2442,
         DP_OP_422J2_124_3477_n2441, DP_OP_422J2_124_3477_n2440,
         DP_OP_422J2_124_3477_n2439, DP_OP_422J2_124_3477_n2438,
         DP_OP_422J2_124_3477_n2437, DP_OP_422J2_124_3477_n2436,
         DP_OP_422J2_124_3477_n2435, DP_OP_422J2_124_3477_n2434,
         DP_OP_422J2_124_3477_n2433, DP_OP_422J2_124_3477_n2432,
         DP_OP_422J2_124_3477_n2430, DP_OP_422J2_124_3477_n2429,
         DP_OP_422J2_124_3477_n2428, DP_OP_422J2_124_3477_n2427,
         DP_OP_422J2_124_3477_n2424, DP_OP_422J2_124_3477_n2423,
         DP_OP_422J2_124_3477_n2422, DP_OP_422J2_124_3477_n2421,
         DP_OP_422J2_124_3477_n2420, DP_OP_422J2_124_3477_n2419,
         DP_OP_422J2_124_3477_n2418, DP_OP_422J2_124_3477_n2417,
         DP_OP_422J2_124_3477_n2416, DP_OP_422J2_124_3477_n2415,
         DP_OP_422J2_124_3477_n2414, DP_OP_422J2_124_3477_n2413,
         DP_OP_422J2_124_3477_n2412, DP_OP_422J2_124_3477_n2411,
         DP_OP_422J2_124_3477_n2410, DP_OP_422J2_124_3477_n2409,
         DP_OP_422J2_124_3477_n2408, DP_OP_422J2_124_3477_n2407,
         DP_OP_422J2_124_3477_n2406, DP_OP_422J2_124_3477_n2405,
         DP_OP_422J2_124_3477_n2404, DP_OP_422J2_124_3477_n2403,
         DP_OP_422J2_124_3477_n2402, DP_OP_422J2_124_3477_n2401,
         DP_OP_422J2_124_3477_n2400, DP_OP_422J2_124_3477_n2399,
         DP_OP_422J2_124_3477_n2398, DP_OP_422J2_124_3477_n2397,
         DP_OP_422J2_124_3477_n2396, DP_OP_422J2_124_3477_n2395,
         DP_OP_422J2_124_3477_n2394, DP_OP_422J2_124_3477_n2393,
         DP_OP_422J2_124_3477_n2392, DP_OP_422J2_124_3477_n2391,
         DP_OP_422J2_124_3477_n2390, DP_OP_422J2_124_3477_n2389,
         DP_OP_422J2_124_3477_n2388, DP_OP_422J2_124_3477_n2387,
         DP_OP_422J2_124_3477_n2386, DP_OP_422J2_124_3477_n2385,
         DP_OP_422J2_124_3477_n2384, DP_OP_422J2_124_3477_n2383,
         DP_OP_422J2_124_3477_n2382, DP_OP_422J2_124_3477_n2381,
         DP_OP_422J2_124_3477_n2380, DP_OP_422J2_124_3477_n2379,
         DP_OP_422J2_124_3477_n2378, DP_OP_422J2_124_3477_n2377,
         DP_OP_422J2_124_3477_n2376, DP_OP_422J2_124_3477_n2375,
         DP_OP_422J2_124_3477_n2374, DP_OP_422J2_124_3477_n2373,
         DP_OP_422J2_124_3477_n2372, DP_OP_422J2_124_3477_n2371,
         DP_OP_422J2_124_3477_n2370, DP_OP_422J2_124_3477_n2369,
         DP_OP_422J2_124_3477_n2368, DP_OP_422J2_124_3477_n2367,
         DP_OP_422J2_124_3477_n2366, DP_OP_422J2_124_3477_n2365,
         DP_OP_422J2_124_3477_n2364, DP_OP_422J2_124_3477_n2363,
         DP_OP_422J2_124_3477_n2362, DP_OP_422J2_124_3477_n2361,
         DP_OP_422J2_124_3477_n2360, DP_OP_422J2_124_3477_n2359,
         DP_OP_422J2_124_3477_n2358, DP_OP_422J2_124_3477_n2357,
         DP_OP_422J2_124_3477_n2356, DP_OP_422J2_124_3477_n2355,
         DP_OP_422J2_124_3477_n2354, DP_OP_422J2_124_3477_n2353,
         DP_OP_422J2_124_3477_n2352, DP_OP_422J2_124_3477_n2351,
         DP_OP_422J2_124_3477_n2350, DP_OP_422J2_124_3477_n2349,
         DP_OP_422J2_124_3477_n2347, DP_OP_422J2_124_3477_n2346,
         DP_OP_422J2_124_3477_n2345, DP_OP_422J2_124_3477_n2344,
         DP_OP_422J2_124_3477_n2343, DP_OP_422J2_124_3477_n2342,
         DP_OP_422J2_124_3477_n2341, DP_OP_422J2_124_3477_n2340,
         DP_OP_422J2_124_3477_n2339, DP_OP_422J2_124_3477_n2338,
         DP_OP_422J2_124_3477_n2336, DP_OP_422J2_124_3477_n2335,
         DP_OP_422J2_124_3477_n2334, DP_OP_422J2_124_3477_n2333,
         DP_OP_422J2_124_3477_n2332, DP_OP_422J2_124_3477_n2331,
         DP_OP_422J2_124_3477_n2330, DP_OP_422J2_124_3477_n2329,
         DP_OP_422J2_124_3477_n2328, DP_OP_422J2_124_3477_n2327,
         DP_OP_422J2_124_3477_n2326, DP_OP_422J2_124_3477_n2325,
         DP_OP_422J2_124_3477_n2324, DP_OP_422J2_124_3477_n2323,
         DP_OP_422J2_124_3477_n2322, DP_OP_422J2_124_3477_n2321,
         DP_OP_422J2_124_3477_n2320, DP_OP_422J2_124_3477_n2319,
         DP_OP_422J2_124_3477_n2318, DP_OP_422J2_124_3477_n2317,
         DP_OP_422J2_124_3477_n2316, DP_OP_422J2_124_3477_n2315,
         DP_OP_422J2_124_3477_n2314, DP_OP_422J2_124_3477_n2313,
         DP_OP_422J2_124_3477_n2312, DP_OP_422J2_124_3477_n2311,
         DP_OP_422J2_124_3477_n2310, DP_OP_422J2_124_3477_n2309,
         DP_OP_422J2_124_3477_n2308, DP_OP_422J2_124_3477_n2307,
         DP_OP_422J2_124_3477_n2306, DP_OP_422J2_124_3477_n2305,
         DP_OP_422J2_124_3477_n2304, DP_OP_422J2_124_3477_n2302,
         DP_OP_422J2_124_3477_n2301, DP_OP_422J2_124_3477_n2299,
         DP_OP_422J2_124_3477_n2298, DP_OP_422J2_124_3477_n2295,
         DP_OP_422J2_124_3477_n2294, DP_OP_422J2_124_3477_n2292,
         DP_OP_422J2_124_3477_n2291, DP_OP_422J2_124_3477_n2290,
         DP_OP_422J2_124_3477_n2289, DP_OP_422J2_124_3477_n2288,
         DP_OP_422J2_124_3477_n2287, DP_OP_422J2_124_3477_n2286,
         DP_OP_422J2_124_3477_n2285, DP_OP_422J2_124_3477_n2284,
         DP_OP_422J2_124_3477_n2283, DP_OP_422J2_124_3477_n2282,
         DP_OP_422J2_124_3477_n2281, DP_OP_422J2_124_3477_n2280,
         DP_OP_422J2_124_3477_n2279, DP_OP_422J2_124_3477_n2278,
         DP_OP_422J2_124_3477_n2277, DP_OP_422J2_124_3477_n2276,
         DP_OP_422J2_124_3477_n2275, DP_OP_422J2_124_3477_n2274,
         DP_OP_422J2_124_3477_n2273, DP_OP_422J2_124_3477_n2272,
         DP_OP_422J2_124_3477_n2271, DP_OP_422J2_124_3477_n2270,
         DP_OP_422J2_124_3477_n2269, DP_OP_422J2_124_3477_n2268,
         DP_OP_422J2_124_3477_n2267, DP_OP_422J2_124_3477_n2266,
         DP_OP_422J2_124_3477_n2265, DP_OP_422J2_124_3477_n2264,
         DP_OP_422J2_124_3477_n2263, DP_OP_422J2_124_3477_n2262,
         DP_OP_422J2_124_3477_n2261, DP_OP_422J2_124_3477_n2260,
         DP_OP_422J2_124_3477_n2259, DP_OP_422J2_124_3477_n2258,
         DP_OP_422J2_124_3477_n2257, DP_OP_422J2_124_3477_n2250,
         DP_OP_422J2_124_3477_n2249, DP_OP_422J2_124_3477_n2248,
         DP_OP_422J2_124_3477_n2247, DP_OP_422J2_124_3477_n2246,
         DP_OP_422J2_124_3477_n2245, DP_OP_422J2_124_3477_n2244,
         DP_OP_422J2_124_3477_n2243, DP_OP_422J2_124_3477_n2242,
         DP_OP_422J2_124_3477_n2241, DP_OP_422J2_124_3477_n2240,
         DP_OP_422J2_124_3477_n2239, DP_OP_422J2_124_3477_n2238,
         DP_OP_422J2_124_3477_n2237, DP_OP_422J2_124_3477_n2236,
         DP_OP_422J2_124_3477_n2235, DP_OP_422J2_124_3477_n2234,
         DP_OP_422J2_124_3477_n2233, DP_OP_422J2_124_3477_n2232,
         DP_OP_422J2_124_3477_n2231, DP_OP_422J2_124_3477_n2230,
         DP_OP_422J2_124_3477_n2229, DP_OP_422J2_124_3477_n2228,
         DP_OP_422J2_124_3477_n2227, DP_OP_422J2_124_3477_n2226,
         DP_OP_422J2_124_3477_n2225, DP_OP_422J2_124_3477_n2224,
         DP_OP_422J2_124_3477_n2223, DP_OP_422J2_124_3477_n2222,
         DP_OP_422J2_124_3477_n2221, DP_OP_422J2_124_3477_n2220,
         DP_OP_422J2_124_3477_n2219, DP_OP_422J2_124_3477_n2218,
         DP_OP_422J2_124_3477_n2217, DP_OP_422J2_124_3477_n2216,
         DP_OP_422J2_124_3477_n2215, DP_OP_422J2_124_3477_n2214,
         DP_OP_422J2_124_3477_n2213, DP_OP_422J2_124_3477_n2211,
         DP_OP_422J2_124_3477_n2210, DP_OP_422J2_124_3477_n2209,
         DP_OP_422J2_124_3477_n2208, DP_OP_422J2_124_3477_n2207,
         DP_OP_422J2_124_3477_n2204, DP_OP_422J2_124_3477_n2203,
         DP_OP_422J2_124_3477_n2202, DP_OP_422J2_124_3477_n2201,
         DP_OP_422J2_124_3477_n2200, DP_OP_422J2_124_3477_n2199,
         DP_OP_422J2_124_3477_n2198, DP_OP_422J2_124_3477_n2197,
         DP_OP_422J2_124_3477_n2196, DP_OP_422J2_124_3477_n2195,
         DP_OP_422J2_124_3477_n2194, DP_OP_422J2_124_3477_n2193,
         DP_OP_422J2_124_3477_n2192, DP_OP_422J2_124_3477_n2191,
         DP_OP_422J2_124_3477_n2190, DP_OP_422J2_124_3477_n2189,
         DP_OP_422J2_124_3477_n2188, DP_OP_422J2_124_3477_n2187,
         DP_OP_422J2_124_3477_n2186, DP_OP_422J2_124_3477_n2185,
         DP_OP_422J2_124_3477_n2184, DP_OP_422J2_124_3477_n2183,
         DP_OP_422J2_124_3477_n2182, DP_OP_422J2_124_3477_n2181,
         DP_OP_422J2_124_3477_n2180, DP_OP_422J2_124_3477_n2179,
         DP_OP_422J2_124_3477_n2178, DP_OP_422J2_124_3477_n2177,
         DP_OP_422J2_124_3477_n2176, DP_OP_422J2_124_3477_n2175,
         DP_OP_422J2_124_3477_n2174, DP_OP_422J2_124_3477_n2173,
         DP_OP_422J2_124_3477_n2171, DP_OP_422J2_124_3477_n2170,
         DP_OP_422J2_124_3477_n2169, DP_OP_422J2_124_3477_n2168,
         DP_OP_422J2_124_3477_n2165, DP_OP_422J2_124_3477_n2164,
         DP_OP_422J2_124_3477_n2163, DP_OP_422J2_124_3477_n2162,
         DP_OP_422J2_124_3477_n2160, DP_OP_422J2_124_3477_n2159,
         DP_OP_422J2_124_3477_n2158, DP_OP_422J2_124_3477_n2157,
         DP_OP_422J2_124_3477_n2156, DP_OP_422J2_124_3477_n2155,
         DP_OP_422J2_124_3477_n2154, DP_OP_422J2_124_3477_n2153,
         DP_OP_422J2_124_3477_n2152, DP_OP_422J2_124_3477_n2151,
         DP_OP_422J2_124_3477_n2150, DP_OP_422J2_124_3477_n2149,
         DP_OP_422J2_124_3477_n2148, DP_OP_422J2_124_3477_n2147,
         DP_OP_422J2_124_3477_n2146, DP_OP_422J2_124_3477_n2145,
         DP_OP_422J2_124_3477_n2144, DP_OP_422J2_124_3477_n2143,
         DP_OP_422J2_124_3477_n2142, DP_OP_422J2_124_3477_n2141,
         DP_OP_422J2_124_3477_n2140, DP_OP_422J2_124_3477_n2139,
         DP_OP_422J2_124_3477_n2138, DP_OP_422J2_124_3477_n2137,
         DP_OP_422J2_124_3477_n2136, DP_OP_422J2_124_3477_n2135,
         DP_OP_422J2_124_3477_n2134, DP_OP_422J2_124_3477_n2133,
         DP_OP_422J2_124_3477_n2132, DP_OP_422J2_124_3477_n2131,
         DP_OP_422J2_124_3477_n2130, DP_OP_422J2_124_3477_n2129,
         DP_OP_422J2_124_3477_n2128, DP_OP_422J2_124_3477_n2127,
         DP_OP_422J2_124_3477_n2125, DP_OP_422J2_124_3477_n2124,
         DP_OP_422J2_124_3477_n2121, DP_OP_422J2_124_3477_n2120,
         DP_OP_422J2_124_3477_n2118, DP_OP_422J2_124_3477_n2117,
         DP_OP_422J2_124_3477_n2116, DP_OP_422J2_124_3477_n2115,
         DP_OP_422J2_124_3477_n2114, DP_OP_422J2_124_3477_n2113,
         DP_OP_422J2_124_3477_n2112, DP_OP_422J2_124_3477_n2111,
         DP_OP_422J2_124_3477_n2110, DP_OP_422J2_124_3477_n2109,
         DP_OP_422J2_124_3477_n2108, DP_OP_422J2_124_3477_n2107,
         DP_OP_422J2_124_3477_n2106, DP_OP_422J2_124_3477_n2105,
         DP_OP_422J2_124_3477_n2104, DP_OP_422J2_124_3477_n2103,
         DP_OP_422J2_124_3477_n2102, DP_OP_422J2_124_3477_n2101,
         DP_OP_422J2_124_3477_n2100, DP_OP_422J2_124_3477_n2099,
         DP_OP_422J2_124_3477_n2098, DP_OP_422J2_124_3477_n2097,
         DP_OP_422J2_124_3477_n2096, DP_OP_422J2_124_3477_n2095,
         DP_OP_422J2_124_3477_n2094, DP_OP_422J2_124_3477_n2093,
         DP_OP_422J2_124_3477_n2092, DP_OP_422J2_124_3477_n2091,
         DP_OP_422J2_124_3477_n2090, DP_OP_422J2_124_3477_n2089,
         DP_OP_422J2_124_3477_n2088, DP_OP_422J2_124_3477_n2087,
         DP_OP_422J2_124_3477_n2086, DP_OP_422J2_124_3477_n2085,
         DP_OP_422J2_124_3477_n2083, DP_OP_422J2_124_3477_n2082,
         DP_OP_422J2_124_3477_n2081, DP_OP_422J2_124_3477_n2078,
         DP_OP_422J2_124_3477_n2076, DP_OP_422J2_124_3477_n2074,
         DP_OP_422J2_124_3477_n2073, DP_OP_422J2_124_3477_n2072,
         DP_OP_422J2_124_3477_n2071, DP_OP_422J2_124_3477_n2070,
         DP_OP_422J2_124_3477_n2069, DP_OP_422J2_124_3477_n2068,
         DP_OP_422J2_124_3477_n2067, DP_OP_422J2_124_3477_n2066,
         DP_OP_422J2_124_3477_n2065, DP_OP_422J2_124_3477_n2064,
         DP_OP_422J2_124_3477_n2063, DP_OP_422J2_124_3477_n2062,
         DP_OP_422J2_124_3477_n2061, DP_OP_422J2_124_3477_n2060,
         DP_OP_422J2_124_3477_n2059, DP_OP_422J2_124_3477_n2058,
         DP_OP_422J2_124_3477_n2057, DP_OP_422J2_124_3477_n2056,
         DP_OP_422J2_124_3477_n2055, DP_OP_422J2_124_3477_n2054,
         DP_OP_422J2_124_3477_n2053, DP_OP_422J2_124_3477_n2052,
         DP_OP_422J2_124_3477_n2051, DP_OP_422J2_124_3477_n2050,
         DP_OP_422J2_124_3477_n2049, DP_OP_422J2_124_3477_n2048,
         DP_OP_422J2_124_3477_n2047, DP_OP_422J2_124_3477_n2046,
         DP_OP_422J2_124_3477_n2045, DP_OP_422J2_124_3477_n2044,
         DP_OP_422J2_124_3477_n2043, DP_OP_422J2_124_3477_n2042,
         DP_OP_422J2_124_3477_n2041, DP_OP_422J2_124_3477_n2040,
         DP_OP_422J2_124_3477_n2039, DP_OP_422J2_124_3477_n2037,
         DP_OP_422J2_124_3477_n2036, DP_OP_422J2_124_3477_n2035,
         DP_OP_422J2_124_3477_n2033, DP_OP_422J2_124_3477_n2032,
         DP_OP_422J2_124_3477_n2031, DP_OP_422J2_124_3477_n2029,
         DP_OP_422J2_124_3477_n2028, DP_OP_422J2_124_3477_n2027,
         DP_OP_422J2_124_3477_n2026, DP_OP_422J2_124_3477_n2025,
         DP_OP_422J2_124_3477_n2024, DP_OP_422J2_124_3477_n2023,
         DP_OP_422J2_124_3477_n2022, DP_OP_422J2_124_3477_n2021,
         DP_OP_422J2_124_3477_n2020, DP_OP_422J2_124_3477_n2019,
         DP_OP_422J2_124_3477_n2018, DP_OP_422J2_124_3477_n2017,
         DP_OP_422J2_124_3477_n2016, DP_OP_422J2_124_3477_n2015,
         DP_OP_422J2_124_3477_n2014, DP_OP_422J2_124_3477_n2013,
         DP_OP_422J2_124_3477_n2012, DP_OP_422J2_124_3477_n2011,
         DP_OP_422J2_124_3477_n2010, DP_OP_422J2_124_3477_n2009,
         DP_OP_422J2_124_3477_n2008, DP_OP_422J2_124_3477_n2007,
         DP_OP_422J2_124_3477_n2006, DP_OP_422J2_124_3477_n2005,
         DP_OP_422J2_124_3477_n2004, DP_OP_422J2_124_3477_n2003,
         DP_OP_422J2_124_3477_n2002, DP_OP_422J2_124_3477_n2001,
         DP_OP_422J2_124_3477_n2000, DP_OP_422J2_124_3477_n1999,
         DP_OP_422J2_124_3477_n1998, DP_OP_422J2_124_3477_n1997,
         DP_OP_422J2_124_3477_n1996, DP_OP_422J2_124_3477_n1995,
         DP_OP_422J2_124_3477_n1994, DP_OP_422J2_124_3477_n1991,
         DP_OP_422J2_124_3477_n1989, DP_OP_422J2_124_3477_n1988,
         DP_OP_422J2_124_3477_n1985, DP_OP_422J2_124_3477_n1984,
         DP_OP_422J2_124_3477_n1983, DP_OP_422J2_124_3477_n1982,
         DP_OP_422J2_124_3477_n1981, DP_OP_422J2_124_3477_n1980,
         DP_OP_422J2_124_3477_n1979, DP_OP_422J2_124_3477_n1978,
         DP_OP_422J2_124_3477_n1977, DP_OP_422J2_124_3477_n1976,
         DP_OP_422J2_124_3477_n1975, DP_OP_422J2_124_3477_n1974,
         DP_OP_422J2_124_3477_n1973, DP_OP_422J2_124_3477_n1972,
         DP_OP_422J2_124_3477_n1971, DP_OP_422J2_124_3477_n1970,
         DP_OP_422J2_124_3477_n1969, DP_OP_422J2_124_3477_n1968,
         DP_OP_422J2_124_3477_n1967, DP_OP_422J2_124_3477_n1966,
         DP_OP_422J2_124_3477_n1965, DP_OP_422J2_124_3477_n1964,
         DP_OP_422J2_124_3477_n1963, DP_OP_422J2_124_3477_n1962,
         DP_OP_422J2_124_3477_n1961, DP_OP_422J2_124_3477_n1960,
         DP_OP_422J2_124_3477_n1959, DP_OP_422J2_124_3477_n1958,
         DP_OP_422J2_124_3477_n1957, DP_OP_422J2_124_3477_n1956,
         DP_OP_422J2_124_3477_n1955, DP_OP_422J2_124_3477_n1954,
         DP_OP_422J2_124_3477_n1952, DP_OP_422J2_124_3477_n1951,
         DP_OP_422J2_124_3477_n1950, DP_OP_422J2_124_3477_n1949,
         DP_OP_422J2_124_3477_n1945, DP_OP_422J2_124_3477_n1943,
         DP_OP_422J2_124_3477_n1941, DP_OP_422J2_124_3477_n1940,
         DP_OP_422J2_124_3477_n1939, DP_OP_422J2_124_3477_n1938,
         DP_OP_422J2_124_3477_n1937, DP_OP_422J2_124_3477_n1936,
         DP_OP_422J2_124_3477_n1935, DP_OP_422J2_124_3477_n1934,
         DP_OP_422J2_124_3477_n1933, DP_OP_422J2_124_3477_n1932,
         DP_OP_422J2_124_3477_n1931, DP_OP_422J2_124_3477_n1930,
         DP_OP_422J2_124_3477_n1929, DP_OP_422J2_124_3477_n1928,
         DP_OP_422J2_124_3477_n1927, DP_OP_422J2_124_3477_n1926,
         DP_OP_422J2_124_3477_n1925, DP_OP_422J2_124_3477_n1924,
         DP_OP_422J2_124_3477_n1923, DP_OP_422J2_124_3477_n1922,
         DP_OP_422J2_124_3477_n1921, DP_OP_422J2_124_3477_n1920,
         DP_OP_422J2_124_3477_n1919, DP_OP_422J2_124_3477_n1918,
         DP_OP_422J2_124_3477_n1917, DP_OP_422J2_124_3477_n1916,
         DP_OP_422J2_124_3477_n1915, DP_OP_422J2_124_3477_n1914,
         DP_OP_422J2_124_3477_n1913, DP_OP_422J2_124_3477_n1912,
         DP_OP_422J2_124_3477_n1911, DP_OP_422J2_124_3477_n1910,
         DP_OP_422J2_124_3477_n1909, DP_OP_422J2_124_3477_n1908,
         DP_OP_422J2_124_3477_n1907, DP_OP_422J2_124_3477_n1906,
         DP_OP_422J2_124_3477_n1905, DP_OP_422J2_124_3477_n1904,
         DP_OP_422J2_124_3477_n1903, DP_OP_422J2_124_3477_n1902,
         DP_OP_422J2_124_3477_n1900, DP_OP_422J2_124_3477_n1899,
         DP_OP_422J2_124_3477_n1898, DP_OP_422J2_124_3477_n1897,
         DP_OP_422J2_124_3477_n1896, DP_OP_422J2_124_3477_n1895,
         DP_OP_422J2_124_3477_n1894, DP_OP_422J2_124_3477_n1893,
         DP_OP_422J2_124_3477_n1892, DP_OP_422J2_124_3477_n1891,
         DP_OP_422J2_124_3477_n1890, DP_OP_422J2_124_3477_n1889,
         DP_OP_422J2_124_3477_n1888, DP_OP_422J2_124_3477_n1887,
         DP_OP_422J2_124_3477_n1886, DP_OP_422J2_124_3477_n1885,
         DP_OP_422J2_124_3477_n1884, DP_OP_422J2_124_3477_n1883,
         DP_OP_422J2_124_3477_n1882, DP_OP_422J2_124_3477_n1881,
         DP_OP_422J2_124_3477_n1880, DP_OP_422J2_124_3477_n1879,
         DP_OP_422J2_124_3477_n1878, DP_OP_422J2_124_3477_n1877,
         DP_OP_422J2_124_3477_n1876, DP_OP_422J2_124_3477_n1875,
         DP_OP_422J2_124_3477_n1874, DP_OP_422J2_124_3477_n1873,
         DP_OP_422J2_124_3477_n1872, DP_OP_422J2_124_3477_n1871,
         DP_OP_422J2_124_3477_n1870, DP_OP_422J2_124_3477_n1869,
         DP_OP_422J2_124_3477_n1868, DP_OP_422J2_124_3477_n1867,
         DP_OP_422J2_124_3477_n1866, DP_OP_422J2_124_3477_n1865,
         DP_OP_422J2_124_3477_n1864, DP_OP_422J2_124_3477_n1863,
         DP_OP_422J2_124_3477_n1862, DP_OP_422J2_124_3477_n1861,
         DP_OP_422J2_124_3477_n1859, DP_OP_422J2_124_3477_n1858,
         DP_OP_422J2_124_3477_n1855, DP_OP_422J2_124_3477_n1854,
         DP_OP_422J2_124_3477_n1853, DP_OP_422J2_124_3477_n1852,
         DP_OP_422J2_124_3477_n1851, DP_OP_422J2_124_3477_n1850,
         DP_OP_422J2_124_3477_n1849, DP_OP_422J2_124_3477_n1848,
         DP_OP_422J2_124_3477_n1847, DP_OP_422J2_124_3477_n1846,
         DP_OP_422J2_124_3477_n1845, DP_OP_422J2_124_3477_n1844,
         DP_OP_422J2_124_3477_n1843, DP_OP_422J2_124_3477_n1842,
         DP_OP_422J2_124_3477_n1841, DP_OP_422J2_124_3477_n1840,
         DP_OP_422J2_124_3477_n1839, DP_OP_422J2_124_3477_n1838,
         DP_OP_422J2_124_3477_n1837, DP_OP_422J2_124_3477_n1836,
         DP_OP_422J2_124_3477_n1835, DP_OP_422J2_124_3477_n1834,
         DP_OP_422J2_124_3477_n1833, DP_OP_422J2_124_3477_n1832,
         DP_OP_422J2_124_3477_n1831, DP_OP_422J2_124_3477_n1830,
         DP_OP_422J2_124_3477_n1829, DP_OP_422J2_124_3477_n1828,
         DP_OP_422J2_124_3477_n1827, DP_OP_422J2_124_3477_n1826,
         DP_OP_422J2_124_3477_n1825, DP_OP_422J2_124_3477_n1824,
         DP_OP_422J2_124_3477_n1823, DP_OP_422J2_124_3477_n1822,
         DP_OP_422J2_124_3477_n1788, DP_OP_422J2_124_3477_n1787,
         DP_OP_422J2_124_3477_n1786, DP_OP_422J2_124_3477_n1785,
         DP_OP_422J2_124_3477_n1784, DP_OP_422J2_124_3477_n1783,
         DP_OP_422J2_124_3477_n1782, DP_OP_422J2_124_3477_n1781,
         DP_OP_422J2_124_3477_n1780, DP_OP_422J2_124_3477_n1779,
         DP_OP_422J2_124_3477_n1778, DP_OP_422J2_124_3477_n1777,
         DP_OP_422J2_124_3477_n1776, DP_OP_422J2_124_3477_n1775,
         DP_OP_422J2_124_3477_n1774, DP_OP_422J2_124_3477_n1773,
         DP_OP_422J2_124_3477_n1772, DP_OP_422J2_124_3477_n1771,
         DP_OP_422J2_124_3477_n1770, DP_OP_422J2_124_3477_n1769,
         DP_OP_422J2_124_3477_n1768, DP_OP_422J2_124_3477_n1767,
         DP_OP_422J2_124_3477_n1766, DP_OP_422J2_124_3477_n1765,
         DP_OP_422J2_124_3477_n1764, DP_OP_422J2_124_3477_n1763,
         DP_OP_422J2_124_3477_n1762, DP_OP_422J2_124_3477_n1761,
         DP_OP_422J2_124_3477_n1760, DP_OP_422J2_124_3477_n1759,
         DP_OP_422J2_124_3477_n1758, DP_OP_422J2_124_3477_n1757,
         DP_OP_422J2_124_3477_n1756, DP_OP_422J2_124_3477_n1755,
         DP_OP_422J2_124_3477_n1754, DP_OP_422J2_124_3477_n1753,
         DP_OP_422J2_124_3477_n1752, DP_OP_422J2_124_3477_n1751,
         DP_OP_422J2_124_3477_n1750, DP_OP_422J2_124_3477_n1749,
         DP_OP_422J2_124_3477_n1748, DP_OP_422J2_124_3477_n1747,
         DP_OP_422J2_124_3477_n1746, DP_OP_422J2_124_3477_n1745,
         DP_OP_422J2_124_3477_n1744, DP_OP_422J2_124_3477_n1743,
         DP_OP_422J2_124_3477_n1742, DP_OP_422J2_124_3477_n1741,
         DP_OP_422J2_124_3477_n1740, DP_OP_422J2_124_3477_n1739,
         DP_OP_422J2_124_3477_n1738, DP_OP_422J2_124_3477_n1737,
         DP_OP_422J2_124_3477_n1736, DP_OP_422J2_124_3477_n1735,
         DP_OP_422J2_124_3477_n1734, DP_OP_422J2_124_3477_n1733,
         DP_OP_422J2_124_3477_n1732, DP_OP_422J2_124_3477_n1731,
         DP_OP_422J2_124_3477_n1730, DP_OP_422J2_124_3477_n1729,
         DP_OP_422J2_124_3477_n1728, DP_OP_422J2_124_3477_n1727,
         DP_OP_422J2_124_3477_n1726, DP_OP_422J2_124_3477_n1725,
         DP_OP_422J2_124_3477_n1724, DP_OP_422J2_124_3477_n1723,
         DP_OP_422J2_124_3477_n1722, DP_OP_422J2_124_3477_n1721,
         DP_OP_422J2_124_3477_n1720, DP_OP_422J2_124_3477_n1719,
         DP_OP_422J2_124_3477_n1718, DP_OP_422J2_124_3477_n1717,
         DP_OP_422J2_124_3477_n1716, DP_OP_422J2_124_3477_n1715,
         DP_OP_422J2_124_3477_n1714, DP_OP_422J2_124_3477_n1713,
         DP_OP_422J2_124_3477_n1712, DP_OP_422J2_124_3477_n1711,
         DP_OP_422J2_124_3477_n1710, DP_OP_422J2_124_3477_n1709,
         DP_OP_422J2_124_3477_n1708, DP_OP_422J2_124_3477_n1707,
         DP_OP_422J2_124_3477_n1706, DP_OP_422J2_124_3477_n1705,
         DP_OP_422J2_124_3477_n1704, DP_OP_422J2_124_3477_n1703,
         DP_OP_422J2_124_3477_n1702, DP_OP_422J2_124_3477_n1701,
         DP_OP_422J2_124_3477_n1700, DP_OP_422J2_124_3477_n1699,
         DP_OP_422J2_124_3477_n1698, DP_OP_422J2_124_3477_n1697,
         DP_OP_422J2_124_3477_n1696, DP_OP_422J2_124_3477_n1695,
         DP_OP_422J2_124_3477_n1694, DP_OP_422J2_124_3477_n1693,
         DP_OP_422J2_124_3477_n1692, DP_OP_422J2_124_3477_n1691,
         DP_OP_422J2_124_3477_n1690, DP_OP_422J2_124_3477_n1689,
         DP_OP_422J2_124_3477_n1688, DP_OP_422J2_124_3477_n1687,
         DP_OP_422J2_124_3477_n1686, DP_OP_422J2_124_3477_n1685,
         DP_OP_422J2_124_3477_n1684, DP_OP_422J2_124_3477_n1683,
         DP_OP_422J2_124_3477_n1682, DP_OP_422J2_124_3477_n1681,
         DP_OP_422J2_124_3477_n1680, DP_OP_422J2_124_3477_n1679,
         DP_OP_422J2_124_3477_n1678, DP_OP_422J2_124_3477_n1677,
         DP_OP_422J2_124_3477_n1676, DP_OP_422J2_124_3477_n1675,
         DP_OP_422J2_124_3477_n1674, DP_OP_422J2_124_3477_n1673,
         DP_OP_422J2_124_3477_n1672, DP_OP_422J2_124_3477_n1671,
         DP_OP_422J2_124_3477_n1670, DP_OP_422J2_124_3477_n1669,
         DP_OP_422J2_124_3477_n1668, DP_OP_422J2_124_3477_n1667,
         DP_OP_422J2_124_3477_n1666, DP_OP_422J2_124_3477_n1665,
         DP_OP_422J2_124_3477_n1664, DP_OP_422J2_124_3477_n1663,
         DP_OP_422J2_124_3477_n1662, DP_OP_422J2_124_3477_n1661,
         DP_OP_422J2_124_3477_n1660, DP_OP_422J2_124_3477_n1659,
         DP_OP_422J2_124_3477_n1658, DP_OP_422J2_124_3477_n1657,
         DP_OP_422J2_124_3477_n1656, DP_OP_422J2_124_3477_n1655,
         DP_OP_422J2_124_3477_n1654, DP_OP_422J2_124_3477_n1653,
         DP_OP_422J2_124_3477_n1652, DP_OP_422J2_124_3477_n1651,
         DP_OP_422J2_124_3477_n1650, DP_OP_422J2_124_3477_n1649,
         DP_OP_422J2_124_3477_n1648, DP_OP_422J2_124_3477_n1647,
         DP_OP_422J2_124_3477_n1646, DP_OP_422J2_124_3477_n1645,
         DP_OP_422J2_124_3477_n1644, DP_OP_422J2_124_3477_n1643,
         DP_OP_422J2_124_3477_n1642, DP_OP_422J2_124_3477_n1641,
         DP_OP_422J2_124_3477_n1640, DP_OP_422J2_124_3477_n1639,
         DP_OP_422J2_124_3477_n1638, DP_OP_422J2_124_3477_n1637,
         DP_OP_422J2_124_3477_n1636, DP_OP_422J2_124_3477_n1635,
         DP_OP_422J2_124_3477_n1634, DP_OP_422J2_124_3477_n1633,
         DP_OP_422J2_124_3477_n1632, DP_OP_422J2_124_3477_n1631,
         DP_OP_422J2_124_3477_n1630, DP_OP_422J2_124_3477_n1629,
         DP_OP_422J2_124_3477_n1628, DP_OP_422J2_124_3477_n1627,
         DP_OP_422J2_124_3477_n1626, DP_OP_422J2_124_3477_n1625,
         DP_OP_422J2_124_3477_n1624, DP_OP_422J2_124_3477_n1623,
         DP_OP_422J2_124_3477_n1622, DP_OP_422J2_124_3477_n1621,
         DP_OP_422J2_124_3477_n1620, DP_OP_422J2_124_3477_n1619,
         DP_OP_422J2_124_3477_n1618, DP_OP_422J2_124_3477_n1617,
         DP_OP_422J2_124_3477_n1616, DP_OP_422J2_124_3477_n1615,
         DP_OP_422J2_124_3477_n1614, DP_OP_422J2_124_3477_n1613,
         DP_OP_422J2_124_3477_n1612, DP_OP_422J2_124_3477_n1611,
         DP_OP_422J2_124_3477_n1610, DP_OP_422J2_124_3477_n1609,
         DP_OP_422J2_124_3477_n1608, DP_OP_422J2_124_3477_n1607,
         DP_OP_422J2_124_3477_n1606, DP_OP_422J2_124_3477_n1605,
         DP_OP_422J2_124_3477_n1604, DP_OP_422J2_124_3477_n1603,
         DP_OP_422J2_124_3477_n1602, DP_OP_422J2_124_3477_n1601,
         DP_OP_422J2_124_3477_n1600, DP_OP_422J2_124_3477_n1599,
         DP_OP_422J2_124_3477_n1598, DP_OP_422J2_124_3477_n1597,
         DP_OP_422J2_124_3477_n1596, DP_OP_422J2_124_3477_n1595,
         DP_OP_422J2_124_3477_n1594, DP_OP_422J2_124_3477_n1593,
         DP_OP_422J2_124_3477_n1592, DP_OP_422J2_124_3477_n1591,
         DP_OP_422J2_124_3477_n1590, DP_OP_422J2_124_3477_n1589,
         DP_OP_422J2_124_3477_n1588, DP_OP_422J2_124_3477_n1587,
         DP_OP_422J2_124_3477_n1586, DP_OP_422J2_124_3477_n1585,
         DP_OP_422J2_124_3477_n1584, DP_OP_422J2_124_3477_n1583,
         DP_OP_422J2_124_3477_n1582, DP_OP_422J2_124_3477_n1581,
         DP_OP_422J2_124_3477_n1580, DP_OP_422J2_124_3477_n1579,
         DP_OP_422J2_124_3477_n1578, DP_OP_422J2_124_3477_n1577,
         DP_OP_422J2_124_3477_n1576, DP_OP_422J2_124_3477_n1575,
         DP_OP_422J2_124_3477_n1574, DP_OP_422J2_124_3477_n1573,
         DP_OP_422J2_124_3477_n1572, DP_OP_422J2_124_3477_n1571,
         DP_OP_422J2_124_3477_n1570, DP_OP_422J2_124_3477_n1569,
         DP_OP_422J2_124_3477_n1568, DP_OP_422J2_124_3477_n1567,
         DP_OP_422J2_124_3477_n1566, DP_OP_422J2_124_3477_n1565,
         DP_OP_422J2_124_3477_n1564, DP_OP_422J2_124_3477_n1563,
         DP_OP_422J2_124_3477_n1562, DP_OP_422J2_124_3477_n1561,
         DP_OP_422J2_124_3477_n1560, DP_OP_422J2_124_3477_n1559,
         DP_OP_422J2_124_3477_n1558, DP_OP_422J2_124_3477_n1557,
         DP_OP_422J2_124_3477_n1556, DP_OP_422J2_124_3477_n1555,
         DP_OP_422J2_124_3477_n1554, DP_OP_422J2_124_3477_n1553,
         DP_OP_422J2_124_3477_n1552, DP_OP_422J2_124_3477_n1551,
         DP_OP_422J2_124_3477_n1550, DP_OP_422J2_124_3477_n1549,
         DP_OP_422J2_124_3477_n1548, DP_OP_422J2_124_3477_n1547,
         DP_OP_422J2_124_3477_n1546, DP_OP_422J2_124_3477_n1545,
         DP_OP_422J2_124_3477_n1544, DP_OP_422J2_124_3477_n1543,
         DP_OP_422J2_124_3477_n1542, DP_OP_422J2_124_3477_n1541,
         DP_OP_422J2_124_3477_n1540, DP_OP_422J2_124_3477_n1539,
         DP_OP_422J2_124_3477_n1538, DP_OP_422J2_124_3477_n1537,
         DP_OP_422J2_124_3477_n1536, DP_OP_422J2_124_3477_n1535,
         DP_OP_422J2_124_3477_n1534, DP_OP_422J2_124_3477_n1533,
         DP_OP_422J2_124_3477_n1532, DP_OP_422J2_124_3477_n1531,
         DP_OP_422J2_124_3477_n1530, DP_OP_422J2_124_3477_n1529,
         DP_OP_422J2_124_3477_n1528, DP_OP_422J2_124_3477_n1527,
         DP_OP_422J2_124_3477_n1526, DP_OP_422J2_124_3477_n1525,
         DP_OP_422J2_124_3477_n1524, DP_OP_422J2_124_3477_n1523,
         DP_OP_422J2_124_3477_n1522, DP_OP_422J2_124_3477_n1521,
         DP_OP_422J2_124_3477_n1520, DP_OP_422J2_124_3477_n1519,
         DP_OP_422J2_124_3477_n1518, DP_OP_422J2_124_3477_n1517,
         DP_OP_422J2_124_3477_n1516, DP_OP_422J2_124_3477_n1515,
         DP_OP_422J2_124_3477_n1514, DP_OP_422J2_124_3477_n1513,
         DP_OP_422J2_124_3477_n1512, DP_OP_422J2_124_3477_n1511,
         DP_OP_422J2_124_3477_n1510, DP_OP_422J2_124_3477_n1509,
         DP_OP_422J2_124_3477_n1508, DP_OP_422J2_124_3477_n1507,
         DP_OP_422J2_124_3477_n1506, DP_OP_422J2_124_3477_n1505,
         DP_OP_422J2_124_3477_n1504, DP_OP_422J2_124_3477_n1503,
         DP_OP_422J2_124_3477_n1502, DP_OP_422J2_124_3477_n1501,
         DP_OP_422J2_124_3477_n1500, DP_OP_422J2_124_3477_n1499,
         DP_OP_422J2_124_3477_n1498, DP_OP_422J2_124_3477_n1497,
         DP_OP_422J2_124_3477_n1496, DP_OP_422J2_124_3477_n1495,
         DP_OP_422J2_124_3477_n1494, DP_OP_422J2_124_3477_n1493,
         DP_OP_422J2_124_3477_n1492, DP_OP_422J2_124_3477_n1491,
         DP_OP_422J2_124_3477_n1490, DP_OP_422J2_124_3477_n1489,
         DP_OP_422J2_124_3477_n1488, DP_OP_422J2_124_3477_n1487,
         DP_OP_422J2_124_3477_n1486, DP_OP_422J2_124_3477_n1485,
         DP_OP_422J2_124_3477_n1484, DP_OP_422J2_124_3477_n1483,
         DP_OP_422J2_124_3477_n1482, DP_OP_422J2_124_3477_n1481,
         DP_OP_422J2_124_3477_n1480, DP_OP_422J2_124_3477_n1479,
         DP_OP_422J2_124_3477_n1478, DP_OP_422J2_124_3477_n1477,
         DP_OP_422J2_124_3477_n1476, DP_OP_422J2_124_3477_n1475,
         DP_OP_422J2_124_3477_n1474, DP_OP_422J2_124_3477_n1473,
         DP_OP_422J2_124_3477_n1472, DP_OP_422J2_124_3477_n1471,
         DP_OP_422J2_124_3477_n1470, DP_OP_422J2_124_3477_n1469,
         DP_OP_422J2_124_3477_n1468, DP_OP_422J2_124_3477_n1467,
         DP_OP_422J2_124_3477_n1466, DP_OP_422J2_124_3477_n1465,
         DP_OP_422J2_124_3477_n1464, DP_OP_422J2_124_3477_n1463,
         DP_OP_422J2_124_3477_n1462, DP_OP_422J2_124_3477_n1461,
         DP_OP_422J2_124_3477_n1460, DP_OP_422J2_124_3477_n1459,
         DP_OP_422J2_124_3477_n1458, DP_OP_422J2_124_3477_n1457,
         DP_OP_422J2_124_3477_n1456, DP_OP_422J2_124_3477_n1455,
         DP_OP_422J2_124_3477_n1454, DP_OP_422J2_124_3477_n1453,
         DP_OP_422J2_124_3477_n1452, DP_OP_422J2_124_3477_n1451,
         DP_OP_422J2_124_3477_n1450, DP_OP_422J2_124_3477_n1449,
         DP_OP_422J2_124_3477_n1448, DP_OP_422J2_124_3477_n1447,
         DP_OP_422J2_124_3477_n1446, DP_OP_422J2_124_3477_n1445,
         DP_OP_422J2_124_3477_n1444, DP_OP_422J2_124_3477_n1443,
         DP_OP_422J2_124_3477_n1442, DP_OP_422J2_124_3477_n1441,
         DP_OP_422J2_124_3477_n1440, DP_OP_422J2_124_3477_n1439,
         DP_OP_422J2_124_3477_n1438, DP_OP_422J2_124_3477_n1437,
         DP_OP_422J2_124_3477_n1436, DP_OP_422J2_124_3477_n1435,
         DP_OP_422J2_124_3477_n1434, DP_OP_422J2_124_3477_n1433,
         DP_OP_422J2_124_3477_n1432, DP_OP_422J2_124_3477_n1431,
         DP_OP_422J2_124_3477_n1430, DP_OP_422J2_124_3477_n1429,
         DP_OP_422J2_124_3477_n1428, DP_OP_422J2_124_3477_n1427,
         DP_OP_422J2_124_3477_n1426, DP_OP_422J2_124_3477_n1425,
         DP_OP_422J2_124_3477_n1424, DP_OP_422J2_124_3477_n1423,
         DP_OP_422J2_124_3477_n1422, DP_OP_422J2_124_3477_n1421,
         DP_OP_422J2_124_3477_n1420, DP_OP_422J2_124_3477_n1419,
         DP_OP_422J2_124_3477_n1418, DP_OP_422J2_124_3477_n1417,
         DP_OP_422J2_124_3477_n1416, DP_OP_422J2_124_3477_n1415,
         DP_OP_422J2_124_3477_n1414, DP_OP_422J2_124_3477_n1413,
         DP_OP_422J2_124_3477_n1412, DP_OP_422J2_124_3477_n1411,
         DP_OP_422J2_124_3477_n1410, DP_OP_422J2_124_3477_n1409,
         DP_OP_422J2_124_3477_n1408, DP_OP_422J2_124_3477_n1407,
         DP_OP_422J2_124_3477_n1406, DP_OP_422J2_124_3477_n1405,
         DP_OP_422J2_124_3477_n1404, DP_OP_422J2_124_3477_n1403,
         DP_OP_422J2_124_3477_n1402, DP_OP_422J2_124_3477_n1401,
         DP_OP_422J2_124_3477_n1400, DP_OP_422J2_124_3477_n1399,
         DP_OP_422J2_124_3477_n1398, DP_OP_422J2_124_3477_n1397,
         DP_OP_422J2_124_3477_n1396, DP_OP_422J2_124_3477_n1395,
         DP_OP_422J2_124_3477_n1394, DP_OP_422J2_124_3477_n1393,
         DP_OP_422J2_124_3477_n1392, DP_OP_422J2_124_3477_n1391,
         DP_OP_422J2_124_3477_n1390, DP_OP_422J2_124_3477_n1389,
         DP_OP_422J2_124_3477_n1388, DP_OP_422J2_124_3477_n1387,
         DP_OP_422J2_124_3477_n1386, DP_OP_422J2_124_3477_n1385,
         DP_OP_422J2_124_3477_n1384, DP_OP_422J2_124_3477_n1383,
         DP_OP_422J2_124_3477_n1382, DP_OP_422J2_124_3477_n1381,
         DP_OP_422J2_124_3477_n1380, DP_OP_422J2_124_3477_n1379,
         DP_OP_422J2_124_3477_n1378, DP_OP_422J2_124_3477_n1377,
         DP_OP_422J2_124_3477_n1376, DP_OP_422J2_124_3477_n1375,
         DP_OP_422J2_124_3477_n1374, DP_OP_422J2_124_3477_n1373,
         DP_OP_422J2_124_3477_n1372, DP_OP_422J2_124_3477_n1371,
         DP_OP_422J2_124_3477_n1370, DP_OP_422J2_124_3477_n1369,
         DP_OP_422J2_124_3477_n1368, DP_OP_422J2_124_3477_n1367,
         DP_OP_422J2_124_3477_n1366, DP_OP_422J2_124_3477_n1365,
         DP_OP_422J2_124_3477_n1364, DP_OP_422J2_124_3477_n1363,
         DP_OP_422J2_124_3477_n1362, DP_OP_422J2_124_3477_n1361,
         DP_OP_422J2_124_3477_n1360, DP_OP_422J2_124_3477_n1359,
         DP_OP_422J2_124_3477_n1358, DP_OP_422J2_124_3477_n1357,
         DP_OP_422J2_124_3477_n1356, DP_OP_422J2_124_3477_n1355,
         DP_OP_422J2_124_3477_n1354, DP_OP_422J2_124_3477_n1353,
         DP_OP_422J2_124_3477_n1352, DP_OP_422J2_124_3477_n1351,
         DP_OP_422J2_124_3477_n1350, DP_OP_422J2_124_3477_n1349,
         DP_OP_422J2_124_3477_n1348, DP_OP_422J2_124_3477_n1347,
         DP_OP_422J2_124_3477_n1346, DP_OP_422J2_124_3477_n1345,
         DP_OP_422J2_124_3477_n1344, DP_OP_422J2_124_3477_n1343,
         DP_OP_422J2_124_3477_n1342, DP_OP_422J2_124_3477_n1341,
         DP_OP_422J2_124_3477_n1340, DP_OP_422J2_124_3477_n1339,
         DP_OP_422J2_124_3477_n1338, DP_OP_422J2_124_3477_n1337,
         DP_OP_422J2_124_3477_n1336, DP_OP_422J2_124_3477_n1335,
         DP_OP_422J2_124_3477_n1334, DP_OP_422J2_124_3477_n1333,
         DP_OP_422J2_124_3477_n1332, DP_OP_422J2_124_3477_n1331,
         DP_OP_422J2_124_3477_n1330, DP_OP_422J2_124_3477_n1329,
         DP_OP_422J2_124_3477_n1328, DP_OP_422J2_124_3477_n1327,
         DP_OP_422J2_124_3477_n1326, DP_OP_422J2_124_3477_n1325,
         DP_OP_422J2_124_3477_n1324, DP_OP_422J2_124_3477_n1323,
         DP_OP_422J2_124_3477_n1322, DP_OP_422J2_124_3477_n1321,
         DP_OP_422J2_124_3477_n1320, DP_OP_422J2_124_3477_n1319,
         DP_OP_422J2_124_3477_n1318, DP_OP_422J2_124_3477_n1317,
         DP_OP_422J2_124_3477_n1316, DP_OP_422J2_124_3477_n1315,
         DP_OP_422J2_124_3477_n1314, DP_OP_422J2_124_3477_n1313,
         DP_OP_422J2_124_3477_n1312, DP_OP_422J2_124_3477_n1311,
         DP_OP_422J2_124_3477_n1310, DP_OP_422J2_124_3477_n1309,
         DP_OP_422J2_124_3477_n1308, DP_OP_422J2_124_3477_n1307,
         DP_OP_422J2_124_3477_n1306, DP_OP_422J2_124_3477_n1305,
         DP_OP_422J2_124_3477_n1304, DP_OP_422J2_124_3477_n1303,
         DP_OP_422J2_124_3477_n1302, DP_OP_422J2_124_3477_n1301,
         DP_OP_422J2_124_3477_n1300, DP_OP_422J2_124_3477_n1299,
         DP_OP_422J2_124_3477_n1298, DP_OP_422J2_124_3477_n1297,
         DP_OP_422J2_124_3477_n1296, DP_OP_422J2_124_3477_n1295,
         DP_OP_422J2_124_3477_n1294, DP_OP_422J2_124_3477_n1293,
         DP_OP_422J2_124_3477_n1292, DP_OP_422J2_124_3477_n1291,
         DP_OP_422J2_124_3477_n1290, DP_OP_422J2_124_3477_n1289,
         DP_OP_422J2_124_3477_n1288, DP_OP_422J2_124_3477_n1287,
         DP_OP_422J2_124_3477_n1286, DP_OP_422J2_124_3477_n1285,
         DP_OP_422J2_124_3477_n1284, DP_OP_422J2_124_3477_n1283,
         DP_OP_422J2_124_3477_n1282, DP_OP_422J2_124_3477_n1281,
         DP_OP_422J2_124_3477_n1280, DP_OP_422J2_124_3477_n1279,
         DP_OP_422J2_124_3477_n1278, DP_OP_422J2_124_3477_n1277,
         DP_OP_422J2_124_3477_n1276, DP_OP_422J2_124_3477_n1275,
         DP_OP_422J2_124_3477_n1274, DP_OP_422J2_124_3477_n1273,
         DP_OP_422J2_124_3477_n1272, DP_OP_422J2_124_3477_n1271,
         DP_OP_422J2_124_3477_n1270, DP_OP_422J2_124_3477_n1269,
         DP_OP_422J2_124_3477_n1268, DP_OP_422J2_124_3477_n1267,
         DP_OP_422J2_124_3477_n1266, DP_OP_422J2_124_3477_n1265,
         DP_OP_422J2_124_3477_n1264, DP_OP_422J2_124_3477_n1263,
         DP_OP_422J2_124_3477_n1262, DP_OP_422J2_124_3477_n1261,
         DP_OP_422J2_124_3477_n1260, DP_OP_422J2_124_3477_n1259,
         DP_OP_422J2_124_3477_n1258, DP_OP_422J2_124_3477_n1257,
         DP_OP_422J2_124_3477_n1256, DP_OP_422J2_124_3477_n1255,
         DP_OP_422J2_124_3477_n1254, DP_OP_422J2_124_3477_n1253,
         DP_OP_422J2_124_3477_n1252, DP_OP_422J2_124_3477_n1251,
         DP_OP_422J2_124_3477_n1250, DP_OP_422J2_124_3477_n1249,
         DP_OP_422J2_124_3477_n1248, DP_OP_422J2_124_3477_n1247,
         DP_OP_422J2_124_3477_n1246, DP_OP_422J2_124_3477_n1245,
         DP_OP_422J2_124_3477_n1244, DP_OP_422J2_124_3477_n1243,
         DP_OP_422J2_124_3477_n1242, DP_OP_422J2_124_3477_n1241,
         DP_OP_422J2_124_3477_n1240, DP_OP_422J2_124_3477_n1239,
         DP_OP_422J2_124_3477_n1238, DP_OP_422J2_124_3477_n1237,
         DP_OP_422J2_124_3477_n1236, DP_OP_422J2_124_3477_n1235,
         DP_OP_422J2_124_3477_n1234, DP_OP_422J2_124_3477_n1233,
         DP_OP_422J2_124_3477_n1232, DP_OP_422J2_124_3477_n1231,
         DP_OP_422J2_124_3477_n1230, DP_OP_422J2_124_3477_n1229,
         DP_OP_422J2_124_3477_n1228, DP_OP_422J2_124_3477_n1227,
         DP_OP_422J2_124_3477_n1226, DP_OP_422J2_124_3477_n1225,
         DP_OP_422J2_124_3477_n1224, DP_OP_422J2_124_3477_n1223,
         DP_OP_422J2_124_3477_n1222, DP_OP_422J2_124_3477_n1221,
         DP_OP_422J2_124_3477_n1220, DP_OP_422J2_124_3477_n1219,
         DP_OP_422J2_124_3477_n1218, DP_OP_422J2_124_3477_n1217,
         DP_OP_422J2_124_3477_n1216, DP_OP_422J2_124_3477_n1215,
         DP_OP_422J2_124_3477_n1214, DP_OP_422J2_124_3477_n1213,
         DP_OP_422J2_124_3477_n1212, DP_OP_422J2_124_3477_n1211,
         DP_OP_422J2_124_3477_n1210, DP_OP_422J2_124_3477_n1209,
         DP_OP_422J2_124_3477_n1208, DP_OP_422J2_124_3477_n1207,
         DP_OP_422J2_124_3477_n1206, DP_OP_422J2_124_3477_n1205,
         DP_OP_422J2_124_3477_n1204, DP_OP_422J2_124_3477_n1203,
         DP_OP_422J2_124_3477_n1202, DP_OP_422J2_124_3477_n1201,
         DP_OP_422J2_124_3477_n1200, DP_OP_422J2_124_3477_n1199,
         DP_OP_422J2_124_3477_n1198, DP_OP_422J2_124_3477_n1197,
         DP_OP_422J2_124_3477_n1196, DP_OP_422J2_124_3477_n1195,
         DP_OP_422J2_124_3477_n1194, DP_OP_422J2_124_3477_n1193,
         DP_OP_422J2_124_3477_n1192, DP_OP_422J2_124_3477_n1191,
         DP_OP_422J2_124_3477_n1190, DP_OP_422J2_124_3477_n1189,
         DP_OP_422J2_124_3477_n1188, DP_OP_422J2_124_3477_n1187,
         DP_OP_422J2_124_3477_n1186, DP_OP_422J2_124_3477_n1185,
         DP_OP_422J2_124_3477_n1184, DP_OP_422J2_124_3477_n1183,
         DP_OP_422J2_124_3477_n1182, DP_OP_422J2_124_3477_n1181,
         DP_OP_422J2_124_3477_n1180, DP_OP_422J2_124_3477_n1179,
         DP_OP_422J2_124_3477_n1178, DP_OP_422J2_124_3477_n1177,
         DP_OP_422J2_124_3477_n1176, DP_OP_422J2_124_3477_n1175,
         DP_OP_422J2_124_3477_n1174, DP_OP_422J2_124_3477_n1173,
         DP_OP_422J2_124_3477_n1172, DP_OP_422J2_124_3477_n1171,
         DP_OP_422J2_124_3477_n1170, DP_OP_422J2_124_3477_n1169,
         DP_OP_422J2_124_3477_n1168, DP_OP_422J2_124_3477_n1167,
         DP_OP_422J2_124_3477_n1166, DP_OP_422J2_124_3477_n1165,
         DP_OP_422J2_124_3477_n1164, DP_OP_422J2_124_3477_n1163,
         DP_OP_422J2_124_3477_n1162, DP_OP_422J2_124_3477_n1161,
         DP_OP_422J2_124_3477_n1160, DP_OP_422J2_124_3477_n1159,
         DP_OP_422J2_124_3477_n1158, DP_OP_422J2_124_3477_n1157,
         DP_OP_422J2_124_3477_n1156, DP_OP_422J2_124_3477_n1155,
         DP_OP_422J2_124_3477_n1154, DP_OP_422J2_124_3477_n1153,
         DP_OP_422J2_124_3477_n1152, DP_OP_422J2_124_3477_n1151,
         DP_OP_422J2_124_3477_n1150, DP_OP_422J2_124_3477_n1149,
         DP_OP_422J2_124_3477_n1148, DP_OP_422J2_124_3477_n1147,
         DP_OP_422J2_124_3477_n1146, DP_OP_422J2_124_3477_n1145,
         DP_OP_422J2_124_3477_n1144, DP_OP_422J2_124_3477_n1143,
         DP_OP_422J2_124_3477_n1142, DP_OP_422J2_124_3477_n1141,
         DP_OP_422J2_124_3477_n1140, DP_OP_422J2_124_3477_n1139,
         DP_OP_422J2_124_3477_n1138, DP_OP_422J2_124_3477_n1137,
         DP_OP_422J2_124_3477_n1136, DP_OP_422J2_124_3477_n1135,
         DP_OP_422J2_124_3477_n1134, DP_OP_422J2_124_3477_n1133,
         DP_OP_422J2_124_3477_n1132, DP_OP_422J2_124_3477_n1131,
         DP_OP_422J2_124_3477_n1130, DP_OP_422J2_124_3477_n1129,
         DP_OP_422J2_124_3477_n1128, DP_OP_422J2_124_3477_n1127,
         DP_OP_422J2_124_3477_n1126, DP_OP_422J2_124_3477_n1125,
         DP_OP_422J2_124_3477_n1124, DP_OP_422J2_124_3477_n1123,
         DP_OP_422J2_124_3477_n1122, DP_OP_422J2_124_3477_n1121,
         DP_OP_422J2_124_3477_n1120, DP_OP_422J2_124_3477_n1119,
         DP_OP_422J2_124_3477_n1118, DP_OP_422J2_124_3477_n1117,
         DP_OP_422J2_124_3477_n1116, DP_OP_422J2_124_3477_n1115,
         DP_OP_422J2_124_3477_n1114, DP_OP_422J2_124_3477_n1113,
         DP_OP_422J2_124_3477_n1112, DP_OP_422J2_124_3477_n1111,
         DP_OP_422J2_124_3477_n1110, DP_OP_422J2_124_3477_n1109,
         DP_OP_422J2_124_3477_n1108, DP_OP_422J2_124_3477_n1107,
         DP_OP_422J2_124_3477_n1106, DP_OP_422J2_124_3477_n1105,
         DP_OP_422J2_124_3477_n1104, DP_OP_422J2_124_3477_n1103,
         DP_OP_422J2_124_3477_n1102, DP_OP_422J2_124_3477_n1101,
         DP_OP_422J2_124_3477_n1100, DP_OP_422J2_124_3477_n1099,
         DP_OP_422J2_124_3477_n1098, DP_OP_422J2_124_3477_n1097,
         DP_OP_422J2_124_3477_n1096, DP_OP_422J2_124_3477_n1095,
         DP_OP_422J2_124_3477_n1094, DP_OP_422J2_124_3477_n1093,
         DP_OP_422J2_124_3477_n1092, DP_OP_422J2_124_3477_n1091,
         DP_OP_422J2_124_3477_n1090, DP_OP_422J2_124_3477_n1089,
         DP_OP_422J2_124_3477_n1088, DP_OP_422J2_124_3477_n1087,
         DP_OP_422J2_124_3477_n1086, DP_OP_422J2_124_3477_n1085,
         DP_OP_422J2_124_3477_n1084, DP_OP_422J2_124_3477_n1083,
         DP_OP_422J2_124_3477_n1082, DP_OP_422J2_124_3477_n1081,
         DP_OP_422J2_124_3477_n1080, DP_OP_422J2_124_3477_n1079,
         DP_OP_422J2_124_3477_n1078, DP_OP_422J2_124_3477_n1077,
         DP_OP_422J2_124_3477_n1076, DP_OP_422J2_124_3477_n1075,
         DP_OP_422J2_124_3477_n1074, DP_OP_422J2_124_3477_n1073,
         DP_OP_422J2_124_3477_n1072, DP_OP_422J2_124_3477_n1071,
         DP_OP_422J2_124_3477_n1070, DP_OP_422J2_124_3477_n1069,
         DP_OP_422J2_124_3477_n1068, DP_OP_422J2_124_3477_n1067,
         DP_OP_422J2_124_3477_n1066, DP_OP_422J2_124_3477_n1065,
         DP_OP_422J2_124_3477_n1064, DP_OP_422J2_124_3477_n1063,
         DP_OP_422J2_124_3477_n1062, DP_OP_422J2_124_3477_n1061,
         DP_OP_422J2_124_3477_n1060, DP_OP_422J2_124_3477_n1059,
         DP_OP_422J2_124_3477_n1058, DP_OP_422J2_124_3477_n1057,
         DP_OP_422J2_124_3477_n1056, DP_OP_422J2_124_3477_n1055,
         DP_OP_422J2_124_3477_n1054, DP_OP_422J2_124_3477_n1053,
         DP_OP_422J2_124_3477_n1052, DP_OP_422J2_124_3477_n1051,
         DP_OP_422J2_124_3477_n1050, DP_OP_422J2_124_3477_n1049,
         DP_OP_422J2_124_3477_n1048, DP_OP_422J2_124_3477_n1047,
         DP_OP_422J2_124_3477_n1046, DP_OP_422J2_124_3477_n1045,
         DP_OP_422J2_124_3477_n1044, DP_OP_422J2_124_3477_n1043,
         DP_OP_422J2_124_3477_n1042, DP_OP_422J2_124_3477_n1041,
         DP_OP_422J2_124_3477_n1040, DP_OP_422J2_124_3477_n1039,
         DP_OP_422J2_124_3477_n1038, DP_OP_422J2_124_3477_n1037,
         DP_OP_422J2_124_3477_n1036, DP_OP_422J2_124_3477_n1035,
         DP_OP_422J2_124_3477_n1034, DP_OP_422J2_124_3477_n1033,
         DP_OP_422J2_124_3477_n1032, DP_OP_422J2_124_3477_n1031,
         DP_OP_422J2_124_3477_n1030, DP_OP_422J2_124_3477_n1029,
         DP_OP_422J2_124_3477_n1028, DP_OP_422J2_124_3477_n1027,
         DP_OP_422J2_124_3477_n1026, DP_OP_422J2_124_3477_n1025,
         DP_OP_422J2_124_3477_n1024, DP_OP_422J2_124_3477_n1023,
         DP_OP_422J2_124_3477_n1022, DP_OP_422J2_124_3477_n1021,
         DP_OP_422J2_124_3477_n1020, DP_OP_422J2_124_3477_n1019,
         DP_OP_422J2_124_3477_n1018, DP_OP_422J2_124_3477_n1017,
         DP_OP_422J2_124_3477_n1016, DP_OP_422J2_124_3477_n1015,
         DP_OP_422J2_124_3477_n1014, DP_OP_422J2_124_3477_n1013,
         DP_OP_422J2_124_3477_n1012, DP_OP_422J2_124_3477_n1011,
         DP_OP_422J2_124_3477_n1010, DP_OP_422J2_124_3477_n1009,
         DP_OP_422J2_124_3477_n1008, DP_OP_422J2_124_3477_n1007,
         DP_OP_422J2_124_3477_n1006, DP_OP_422J2_124_3477_n1005,
         DP_OP_422J2_124_3477_n1004, DP_OP_422J2_124_3477_n1003,
         DP_OP_422J2_124_3477_n1002, DP_OP_422J2_124_3477_n1001,
         DP_OP_422J2_124_3477_n1000, DP_OP_422J2_124_3477_n999,
         DP_OP_422J2_124_3477_n998, DP_OP_422J2_124_3477_n997,
         DP_OP_422J2_124_3477_n996, DP_OP_422J2_124_3477_n995,
         DP_OP_422J2_124_3477_n994, DP_OP_422J2_124_3477_n993,
         DP_OP_422J2_124_3477_n992, DP_OP_422J2_124_3477_n991,
         DP_OP_422J2_124_3477_n990, DP_OP_422J2_124_3477_n989,
         DP_OP_422J2_124_3477_n988, DP_OP_422J2_124_3477_n987,
         DP_OP_422J2_124_3477_n986, DP_OP_422J2_124_3477_n985,
         DP_OP_422J2_124_3477_n984, DP_OP_422J2_124_3477_n983,
         DP_OP_422J2_124_3477_n982, DP_OP_422J2_124_3477_n981,
         DP_OP_422J2_124_3477_n980, DP_OP_422J2_124_3477_n979,
         DP_OP_422J2_124_3477_n978, DP_OP_422J2_124_3477_n977,
         DP_OP_422J2_124_3477_n976, DP_OP_422J2_124_3477_n975,
         DP_OP_422J2_124_3477_n974, DP_OP_422J2_124_3477_n973,
         DP_OP_422J2_124_3477_n972, DP_OP_422J2_124_3477_n971,
         DP_OP_422J2_124_3477_n970, DP_OP_422J2_124_3477_n969,
         DP_OP_422J2_124_3477_n968, DP_OP_422J2_124_3477_n967,
         DP_OP_422J2_124_3477_n966, DP_OP_422J2_124_3477_n965,
         DP_OP_422J2_124_3477_n964, DP_OP_422J2_124_3477_n963,
         DP_OP_422J2_124_3477_n962, DP_OP_422J2_124_3477_n961,
         DP_OP_422J2_124_3477_n960, DP_OP_422J2_124_3477_n959,
         DP_OP_422J2_124_3477_n958, DP_OP_422J2_124_3477_n957,
         DP_OP_422J2_124_3477_n956, DP_OP_422J2_124_3477_n955,
         DP_OP_422J2_124_3477_n954, DP_OP_422J2_124_3477_n953,
         DP_OP_422J2_124_3477_n952, DP_OP_422J2_124_3477_n951,
         DP_OP_422J2_124_3477_n950, DP_OP_422J2_124_3477_n949,
         DP_OP_422J2_124_3477_n948, DP_OP_422J2_124_3477_n947,
         DP_OP_422J2_124_3477_n946, DP_OP_422J2_124_3477_n945,
         DP_OP_422J2_124_3477_n944, DP_OP_422J2_124_3477_n943,
         DP_OP_422J2_124_3477_n942, DP_OP_422J2_124_3477_n941,
         DP_OP_422J2_124_3477_n940, DP_OP_422J2_124_3477_n939,
         DP_OP_422J2_124_3477_n938, DP_OP_422J2_124_3477_n937,
         DP_OP_422J2_124_3477_n936, DP_OP_422J2_124_3477_n935,
         DP_OP_422J2_124_3477_n934, DP_OP_422J2_124_3477_n933,
         DP_OP_422J2_124_3477_n932, DP_OP_422J2_124_3477_n931,
         DP_OP_422J2_124_3477_n930, DP_OP_422J2_124_3477_n929,
         DP_OP_422J2_124_3477_n928, DP_OP_422J2_124_3477_n927,
         DP_OP_422J2_124_3477_n926, DP_OP_422J2_124_3477_n925,
         DP_OP_422J2_124_3477_n924, DP_OP_422J2_124_3477_n923,
         DP_OP_422J2_124_3477_n922, DP_OP_422J2_124_3477_n921,
         DP_OP_422J2_124_3477_n920, DP_OP_422J2_124_3477_n919,
         DP_OP_422J2_124_3477_n918, DP_OP_422J2_124_3477_n917,
         DP_OP_422J2_124_3477_n916, DP_OP_422J2_124_3477_n915,
         DP_OP_422J2_124_3477_n914, DP_OP_422J2_124_3477_n913,
         DP_OP_422J2_124_3477_n912, DP_OP_422J2_124_3477_n911,
         DP_OP_422J2_124_3477_n910, DP_OP_422J2_124_3477_n909,
         DP_OP_422J2_124_3477_n908, DP_OP_422J2_124_3477_n907,
         DP_OP_422J2_124_3477_n906, DP_OP_422J2_124_3477_n905,
         DP_OP_422J2_124_3477_n904, DP_OP_422J2_124_3477_n903,
         DP_OP_422J2_124_3477_n902, DP_OP_422J2_124_3477_n901,
         DP_OP_422J2_124_3477_n900, DP_OP_422J2_124_3477_n899,
         DP_OP_422J2_124_3477_n898, DP_OP_422J2_124_3477_n897,
         DP_OP_422J2_124_3477_n896, DP_OP_422J2_124_3477_n895,
         DP_OP_422J2_124_3477_n894, DP_OP_422J2_124_3477_n893,
         DP_OP_422J2_124_3477_n892, DP_OP_422J2_124_3477_n891,
         DP_OP_422J2_124_3477_n890, DP_OP_422J2_124_3477_n889,
         DP_OP_422J2_124_3477_n888, DP_OP_422J2_124_3477_n887,
         DP_OP_422J2_124_3477_n886, DP_OP_422J2_124_3477_n885,
         DP_OP_422J2_124_3477_n884, DP_OP_422J2_124_3477_n883,
         DP_OP_422J2_124_3477_n882, DP_OP_422J2_124_3477_n881,
         DP_OP_422J2_124_3477_n880, DP_OP_422J2_124_3477_n879,
         DP_OP_422J2_124_3477_n878, DP_OP_422J2_124_3477_n877,
         DP_OP_422J2_124_3477_n876, DP_OP_422J2_124_3477_n875,
         DP_OP_422J2_124_3477_n874, DP_OP_422J2_124_3477_n873,
         DP_OP_422J2_124_3477_n872, DP_OP_422J2_124_3477_n871,
         DP_OP_422J2_124_3477_n870, DP_OP_422J2_124_3477_n869,
         DP_OP_422J2_124_3477_n868, DP_OP_422J2_124_3477_n867,
         DP_OP_422J2_124_3477_n866, DP_OP_422J2_124_3477_n865,
         DP_OP_422J2_124_3477_n864, DP_OP_422J2_124_3477_n863,
         DP_OP_422J2_124_3477_n862, DP_OP_422J2_124_3477_n861,
         DP_OP_422J2_124_3477_n860, DP_OP_422J2_124_3477_n859,
         DP_OP_422J2_124_3477_n858, DP_OP_422J2_124_3477_n857,
         DP_OP_422J2_124_3477_n856, DP_OP_422J2_124_3477_n855,
         DP_OP_422J2_124_3477_n854, DP_OP_422J2_124_3477_n853,
         DP_OP_422J2_124_3477_n852, DP_OP_422J2_124_3477_n851,
         DP_OP_422J2_124_3477_n850, DP_OP_422J2_124_3477_n849,
         DP_OP_422J2_124_3477_n848, DP_OP_422J2_124_3477_n847,
         DP_OP_422J2_124_3477_n846, DP_OP_422J2_124_3477_n845,
         DP_OP_422J2_124_3477_n844, DP_OP_422J2_124_3477_n843,
         DP_OP_422J2_124_3477_n842, DP_OP_422J2_124_3477_n841,
         DP_OP_422J2_124_3477_n840, DP_OP_422J2_124_3477_n839,
         DP_OP_422J2_124_3477_n838, DP_OP_422J2_124_3477_n837,
         DP_OP_422J2_124_3477_n836, DP_OP_422J2_124_3477_n835,
         DP_OP_422J2_124_3477_n834, DP_OP_422J2_124_3477_n833,
         DP_OP_422J2_124_3477_n832, DP_OP_422J2_124_3477_n831,
         DP_OP_422J2_124_3477_n830, DP_OP_422J2_124_3477_n829,
         DP_OP_422J2_124_3477_n828, DP_OP_422J2_124_3477_n827,
         DP_OP_422J2_124_3477_n826, DP_OP_422J2_124_3477_n825,
         DP_OP_422J2_124_3477_n824, DP_OP_422J2_124_3477_n823,
         DP_OP_422J2_124_3477_n822, DP_OP_422J2_124_3477_n821,
         DP_OP_422J2_124_3477_n820, DP_OP_422J2_124_3477_n819,
         DP_OP_422J2_124_3477_n818, DP_OP_422J2_124_3477_n817,
         DP_OP_422J2_124_3477_n816, DP_OP_422J2_124_3477_n815,
         DP_OP_422J2_124_3477_n814, DP_OP_422J2_124_3477_n813,
         DP_OP_422J2_124_3477_n812, DP_OP_422J2_124_3477_n811,
         DP_OP_422J2_124_3477_n810, DP_OP_422J2_124_3477_n809,
         DP_OP_422J2_124_3477_n808, DP_OP_422J2_124_3477_n807,
         DP_OP_422J2_124_3477_n806, DP_OP_422J2_124_3477_n805,
         DP_OP_422J2_124_3477_n804, DP_OP_422J2_124_3477_n803,
         DP_OP_422J2_124_3477_n802, DP_OP_422J2_124_3477_n801,
         DP_OP_422J2_124_3477_n800, DP_OP_422J2_124_3477_n799,
         DP_OP_422J2_124_3477_n798, DP_OP_422J2_124_3477_n797,
         DP_OP_422J2_124_3477_n796, DP_OP_422J2_124_3477_n795,
         DP_OP_422J2_124_3477_n794, DP_OP_422J2_124_3477_n793,
         DP_OP_422J2_124_3477_n792, DP_OP_422J2_124_3477_n791,
         DP_OP_422J2_124_3477_n790, DP_OP_422J2_124_3477_n789,
         DP_OP_422J2_124_3477_n788, DP_OP_422J2_124_3477_n787,
         DP_OP_422J2_124_3477_n786, DP_OP_422J2_124_3477_n785,
         DP_OP_422J2_124_3477_n784, DP_OP_422J2_124_3477_n783,
         DP_OP_422J2_124_3477_n782, DP_OP_422J2_124_3477_n781,
         DP_OP_422J2_124_3477_n780, DP_OP_422J2_124_3477_n779,
         DP_OP_422J2_124_3477_n778, DP_OP_422J2_124_3477_n777,
         DP_OP_422J2_124_3477_n776, DP_OP_422J2_124_3477_n775,
         DP_OP_422J2_124_3477_n774, DP_OP_422J2_124_3477_n773,
         DP_OP_422J2_124_3477_n772, DP_OP_422J2_124_3477_n771,
         DP_OP_422J2_124_3477_n770, DP_OP_422J2_124_3477_n769,
         DP_OP_422J2_124_3477_n768, DP_OP_422J2_124_3477_n767,
         DP_OP_422J2_124_3477_n766, DP_OP_422J2_124_3477_n765,
         DP_OP_422J2_124_3477_n764, DP_OP_422J2_124_3477_n763,
         DP_OP_422J2_124_3477_n762, DP_OP_422J2_124_3477_n761,
         DP_OP_422J2_124_3477_n760, DP_OP_422J2_124_3477_n759,
         DP_OP_422J2_124_3477_n758, DP_OP_422J2_124_3477_n757,
         DP_OP_422J2_124_3477_n756, DP_OP_422J2_124_3477_n755,
         DP_OP_422J2_124_3477_n754, DP_OP_422J2_124_3477_n753,
         DP_OP_422J2_124_3477_n752, DP_OP_422J2_124_3477_n751,
         DP_OP_422J2_124_3477_n750, DP_OP_422J2_124_3477_n749,
         DP_OP_422J2_124_3477_n748, DP_OP_422J2_124_3477_n747,
         DP_OP_422J2_124_3477_n746, DP_OP_422J2_124_3477_n745,
         DP_OP_422J2_124_3477_n744, DP_OP_422J2_124_3477_n743,
         DP_OP_422J2_124_3477_n742, DP_OP_422J2_124_3477_n741,
         DP_OP_422J2_124_3477_n740, DP_OP_422J2_124_3477_n739,
         DP_OP_422J2_124_3477_n738, DP_OP_422J2_124_3477_n737,
         DP_OP_422J2_124_3477_n736, DP_OP_422J2_124_3477_n735,
         DP_OP_422J2_124_3477_n734, DP_OP_422J2_124_3477_n733,
         DP_OP_422J2_124_3477_n732, DP_OP_422J2_124_3477_n731,
         DP_OP_422J2_124_3477_n730, DP_OP_422J2_124_3477_n729,
         DP_OP_422J2_124_3477_n728, DP_OP_422J2_124_3477_n727,
         DP_OP_422J2_124_3477_n726, DP_OP_422J2_124_3477_n725,
         DP_OP_422J2_124_3477_n724, DP_OP_422J2_124_3477_n723,
         DP_OP_422J2_124_3477_n722, DP_OP_422J2_124_3477_n721,
         DP_OP_422J2_124_3477_n720, DP_OP_422J2_124_3477_n719,
         DP_OP_422J2_124_3477_n718, DP_OP_422J2_124_3477_n717,
         DP_OP_422J2_124_3477_n716, DP_OP_422J2_124_3477_n715,
         DP_OP_422J2_124_3477_n714, DP_OP_422J2_124_3477_n713,
         DP_OP_422J2_124_3477_n712, DP_OP_422J2_124_3477_n711,
         DP_OP_422J2_124_3477_n710, DP_OP_422J2_124_3477_n709,
         DP_OP_422J2_124_3477_n708, DP_OP_422J2_124_3477_n707,
         DP_OP_422J2_124_3477_n706, DP_OP_422J2_124_3477_n705,
         DP_OP_422J2_124_3477_n704, DP_OP_422J2_124_3477_n703,
         DP_OP_422J2_124_3477_n702, DP_OP_422J2_124_3477_n701,
         DP_OP_422J2_124_3477_n700, DP_OP_422J2_124_3477_n699,
         DP_OP_422J2_124_3477_n698, DP_OP_422J2_124_3477_n697,
         DP_OP_422J2_124_3477_n696, DP_OP_422J2_124_3477_n695,
         DP_OP_422J2_124_3477_n694, DP_OP_422J2_124_3477_n693,
         DP_OP_422J2_124_3477_n692, DP_OP_422J2_124_3477_n691,
         DP_OP_422J2_124_3477_n690, DP_OP_422J2_124_3477_n689,
         DP_OP_422J2_124_3477_n688, DP_OP_422J2_124_3477_n687,
         DP_OP_422J2_124_3477_n686, DP_OP_422J2_124_3477_n685,
         DP_OP_422J2_124_3477_n684, DP_OP_422J2_124_3477_n683,
         DP_OP_422J2_124_3477_n682, DP_OP_422J2_124_3477_n681,
         DP_OP_422J2_124_3477_n680, DP_OP_422J2_124_3477_n679,
         DP_OP_422J2_124_3477_n678, DP_OP_422J2_124_3477_n677,
         DP_OP_422J2_124_3477_n676, DP_OP_422J2_124_3477_n675,
         DP_OP_422J2_124_3477_n674, DP_OP_422J2_124_3477_n673,
         DP_OP_422J2_124_3477_n672, DP_OP_422J2_124_3477_n671,
         DP_OP_422J2_124_3477_n670, DP_OP_422J2_124_3477_n669,
         DP_OP_422J2_124_3477_n668, DP_OP_422J2_124_3477_n667,
         DP_OP_422J2_124_3477_n666, DP_OP_422J2_124_3477_n665,
         DP_OP_422J2_124_3477_n664, DP_OP_422J2_124_3477_n663,
         DP_OP_422J2_124_3477_n662, DP_OP_422J2_124_3477_n661,
         DP_OP_422J2_124_3477_n660, DP_OP_422J2_124_3477_n659,
         DP_OP_422J2_124_3477_n658, DP_OP_422J2_124_3477_n657,
         DP_OP_422J2_124_3477_n656, DP_OP_422J2_124_3477_n655,
         DP_OP_422J2_124_3477_n654, DP_OP_422J2_124_3477_n653,
         DP_OP_422J2_124_3477_n652, DP_OP_422J2_124_3477_n651,
         DP_OP_422J2_124_3477_n650, DP_OP_422J2_124_3477_n649,
         DP_OP_422J2_124_3477_n648, DP_OP_422J2_124_3477_n647,
         DP_OP_422J2_124_3477_n646, DP_OP_422J2_124_3477_n645,
         DP_OP_422J2_124_3477_n644, DP_OP_422J2_124_3477_n643,
         DP_OP_422J2_124_3477_n642, DP_OP_422J2_124_3477_n641,
         DP_OP_422J2_124_3477_n640, DP_OP_422J2_124_3477_n639,
         DP_OP_422J2_124_3477_n638, DP_OP_422J2_124_3477_n637,
         DP_OP_422J2_124_3477_n636, DP_OP_422J2_124_3477_n635,
         DP_OP_422J2_124_3477_n634, DP_OP_422J2_124_3477_n633,
         DP_OP_422J2_124_3477_n632, DP_OP_422J2_124_3477_n631,
         DP_OP_422J2_124_3477_n630, DP_OP_422J2_124_3477_n629,
         DP_OP_422J2_124_3477_n628, DP_OP_422J2_124_3477_n627,
         DP_OP_422J2_124_3477_n626, DP_OP_422J2_124_3477_n625,
         DP_OP_422J2_124_3477_n624, DP_OP_422J2_124_3477_n623,
         DP_OP_422J2_124_3477_n622, DP_OP_422J2_124_3477_n621,
         DP_OP_422J2_124_3477_n620, DP_OP_422J2_124_3477_n619,
         DP_OP_422J2_124_3477_n618, DP_OP_422J2_124_3477_n617,
         DP_OP_422J2_124_3477_n616, DP_OP_422J2_124_3477_n615,
         DP_OP_422J2_124_3477_n614, DP_OP_422J2_124_3477_n613,
         DP_OP_422J2_124_3477_n612, DP_OP_422J2_124_3477_n611,
         DP_OP_422J2_124_3477_n610, DP_OP_422J2_124_3477_n609,
         DP_OP_422J2_124_3477_n608, DP_OP_422J2_124_3477_n607,
         DP_OP_422J2_124_3477_n606, DP_OP_422J2_124_3477_n605,
         DP_OP_422J2_124_3477_n604, DP_OP_422J2_124_3477_n603,
         DP_OP_422J2_124_3477_n602, DP_OP_422J2_124_3477_n601,
         DP_OP_422J2_124_3477_n600, DP_OP_422J2_124_3477_n599,
         DP_OP_422J2_124_3477_n598, DP_OP_422J2_124_3477_n597,
         DP_OP_422J2_124_3477_n596, DP_OP_422J2_124_3477_n595,
         DP_OP_422J2_124_3477_n594, DP_OP_422J2_124_3477_n593,
         DP_OP_422J2_124_3477_n592, DP_OP_422J2_124_3477_n591,
         DP_OP_422J2_124_3477_n590, DP_OP_422J2_124_3477_n589,
         DP_OP_422J2_124_3477_n588, DP_OP_422J2_124_3477_n587,
         DP_OP_422J2_124_3477_n586, DP_OP_422J2_124_3477_n585,
         DP_OP_422J2_124_3477_n584, DP_OP_422J2_124_3477_n583,
         DP_OP_422J2_124_3477_n582, DP_OP_422J2_124_3477_n581,
         DP_OP_422J2_124_3477_n580, DP_OP_422J2_124_3477_n579,
         DP_OP_422J2_124_3477_n578, DP_OP_422J2_124_3477_n577,
         DP_OP_422J2_124_3477_n576, DP_OP_422J2_124_3477_n575,
         DP_OP_422J2_124_3477_n574, DP_OP_422J2_124_3477_n573,
         DP_OP_422J2_124_3477_n572, DP_OP_422J2_124_3477_n571,
         DP_OP_422J2_124_3477_n570, DP_OP_422J2_124_3477_n569,
         DP_OP_422J2_124_3477_n568, DP_OP_422J2_124_3477_n567,
         DP_OP_422J2_124_3477_n566, DP_OP_422J2_124_3477_n565,
         DP_OP_422J2_124_3477_n564, DP_OP_422J2_124_3477_n563,
         DP_OP_422J2_124_3477_n562, DP_OP_422J2_124_3477_n561,
         DP_OP_422J2_124_3477_n560, DP_OP_422J2_124_3477_n559,
         DP_OP_422J2_124_3477_n558, DP_OP_422J2_124_3477_n557,
         DP_OP_422J2_124_3477_n556, DP_OP_422J2_124_3477_n555,
         DP_OP_422J2_124_3477_n554, DP_OP_422J2_124_3477_n553,
         DP_OP_422J2_124_3477_n552, DP_OP_422J2_124_3477_n551,
         DP_OP_422J2_124_3477_n550, DP_OP_422J2_124_3477_n549,
         DP_OP_422J2_124_3477_n548, DP_OP_422J2_124_3477_n547,
         DP_OP_422J2_124_3477_n546, DP_OP_422J2_124_3477_n545,
         DP_OP_422J2_124_3477_n544, DP_OP_422J2_124_3477_n543,
         DP_OP_422J2_124_3477_n542, DP_OP_422J2_124_3477_n541,
         DP_OP_422J2_124_3477_n540, DP_OP_422J2_124_3477_n539,
         DP_OP_422J2_124_3477_n538, DP_OP_422J2_124_3477_n537,
         DP_OP_422J2_124_3477_n536, DP_OP_422J2_124_3477_n535,
         DP_OP_422J2_124_3477_n534, DP_OP_422J2_124_3477_n533,
         DP_OP_422J2_124_3477_n532, DP_OP_422J2_124_3477_n531,
         DP_OP_422J2_124_3477_n530, DP_OP_422J2_124_3477_n529,
         DP_OP_422J2_124_3477_n528, DP_OP_422J2_124_3477_n527,
         DP_OP_422J2_124_3477_n526, DP_OP_422J2_124_3477_n525,
         DP_OP_422J2_124_3477_n524, DP_OP_422J2_124_3477_n523,
         DP_OP_422J2_124_3477_n522, DP_OP_422J2_124_3477_n521,
         DP_OP_422J2_124_3477_n520, DP_OP_422J2_124_3477_n519,
         DP_OP_422J2_124_3477_n518, DP_OP_422J2_124_3477_n517,
         DP_OP_422J2_124_3477_n516, DP_OP_422J2_124_3477_n515,
         DP_OP_422J2_124_3477_n514, DP_OP_422J2_124_3477_n513,
         DP_OP_422J2_124_3477_n512, DP_OP_422J2_124_3477_n511,
         DP_OP_422J2_124_3477_n510, DP_OP_422J2_124_3477_n509,
         DP_OP_422J2_124_3477_n508, DP_OP_422J2_124_3477_n507,
         DP_OP_422J2_124_3477_n506, DP_OP_422J2_124_3477_n505,
         DP_OP_422J2_124_3477_n504, DP_OP_422J2_124_3477_n503,
         DP_OP_422J2_124_3477_n502, DP_OP_422J2_124_3477_n501,
         DP_OP_422J2_124_3477_n500, DP_OP_422J2_124_3477_n499,
         DP_OP_422J2_124_3477_n498, DP_OP_422J2_124_3477_n497,
         DP_OP_422J2_124_3477_n496, DP_OP_422J2_124_3477_n495,
         DP_OP_422J2_124_3477_n494, DP_OP_422J2_124_3477_n493,
         DP_OP_422J2_124_3477_n492, DP_OP_422J2_124_3477_n491,
         DP_OP_422J2_124_3477_n490, DP_OP_422J2_124_3477_n489,
         DP_OP_422J2_124_3477_n488, DP_OP_422J2_124_3477_n487,
         DP_OP_422J2_124_3477_n486, DP_OP_422J2_124_3477_n485,
         DP_OP_422J2_124_3477_n484, DP_OP_422J2_124_3477_n483,
         DP_OP_422J2_124_3477_n482, DP_OP_422J2_124_3477_n481,
         DP_OP_422J2_124_3477_n480, DP_OP_422J2_124_3477_n479,
         DP_OP_422J2_124_3477_n478, DP_OP_422J2_124_3477_n477,
         DP_OP_422J2_124_3477_n476, DP_OP_422J2_124_3477_n475,
         DP_OP_422J2_124_3477_n474, DP_OP_422J2_124_3477_n473,
         DP_OP_422J2_124_3477_n472, DP_OP_422J2_124_3477_n471,
         DP_OP_422J2_124_3477_n470, DP_OP_422J2_124_3477_n469,
         DP_OP_422J2_124_3477_n468, DP_OP_422J2_124_3477_n467,
         DP_OP_422J2_124_3477_n466, DP_OP_422J2_124_3477_n465,
         DP_OP_422J2_124_3477_n464, DP_OP_422J2_124_3477_n463,
         DP_OP_422J2_124_3477_n462, DP_OP_422J2_124_3477_n461,
         DP_OP_422J2_124_3477_n460, DP_OP_422J2_124_3477_n459,
         DP_OP_422J2_124_3477_n458, DP_OP_422J2_124_3477_n457,
         DP_OP_422J2_124_3477_n456, DP_OP_422J2_124_3477_n455,
         DP_OP_422J2_124_3477_n454, DP_OP_422J2_124_3477_n453,
         DP_OP_422J2_124_3477_n452, DP_OP_422J2_124_3477_n451,
         DP_OP_422J2_124_3477_n450, DP_OP_422J2_124_3477_n449,
         DP_OP_422J2_124_3477_n448, DP_OP_422J2_124_3477_n447,
         DP_OP_422J2_124_3477_n446, DP_OP_422J2_124_3477_n445,
         DP_OP_422J2_124_3477_n444, DP_OP_422J2_124_3477_n443,
         DP_OP_422J2_124_3477_n442, DP_OP_422J2_124_3477_n441,
         DP_OP_422J2_124_3477_n440, DP_OP_422J2_124_3477_n439,
         DP_OP_422J2_124_3477_n438, DP_OP_422J2_124_3477_n437,
         DP_OP_422J2_124_3477_n436, DP_OP_422J2_124_3477_n435,
         DP_OP_422J2_124_3477_n434, DP_OP_422J2_124_3477_n433,
         DP_OP_422J2_124_3477_n432, DP_OP_422J2_124_3477_n431,
         DP_OP_422J2_124_3477_n430, DP_OP_422J2_124_3477_n429,
         DP_OP_422J2_124_3477_n428, DP_OP_422J2_124_3477_n427,
         DP_OP_422J2_124_3477_n426, DP_OP_422J2_124_3477_n425,
         DP_OP_422J2_124_3477_n424, DP_OP_422J2_124_3477_n423,
         DP_OP_422J2_124_3477_n422, DP_OP_422J2_124_3477_n421,
         DP_OP_422J2_124_3477_n420, DP_OP_422J2_124_3477_n419,
         DP_OP_422J2_124_3477_n418, DP_OP_422J2_124_3477_n417,
         DP_OP_422J2_124_3477_n416, DP_OP_422J2_124_3477_n415,
         DP_OP_422J2_124_3477_n414, DP_OP_422J2_124_3477_n413,
         DP_OP_422J2_124_3477_n412, DP_OP_422J2_124_3477_n411,
         DP_OP_422J2_124_3477_n410, DP_OP_422J2_124_3477_n409,
         DP_OP_422J2_124_3477_n408, DP_OP_422J2_124_3477_n407,
         DP_OP_422J2_124_3477_n406, DP_OP_422J2_124_3477_n405,
         DP_OP_422J2_124_3477_n404, DP_OP_422J2_124_3477_n403,
         DP_OP_422J2_124_3477_n402, DP_OP_422J2_124_3477_n401,
         DP_OP_422J2_124_3477_n400, DP_OP_422J2_124_3477_n399,
         DP_OP_422J2_124_3477_n398, DP_OP_422J2_124_3477_n397,
         DP_OP_422J2_124_3477_n396, DP_OP_422J2_124_3477_n395,
         DP_OP_422J2_124_3477_n394, DP_OP_422J2_124_3477_n393,
         DP_OP_422J2_124_3477_n392, DP_OP_422J2_124_3477_n391,
         DP_OP_422J2_124_3477_n390, DP_OP_422J2_124_3477_n389,
         DP_OP_422J2_124_3477_n388, DP_OP_422J2_124_3477_n387,
         DP_OP_422J2_124_3477_n386, DP_OP_422J2_124_3477_n385,
         DP_OP_422J2_124_3477_n384, DP_OP_422J2_124_3477_n383,
         DP_OP_422J2_124_3477_n382, DP_OP_422J2_124_3477_n381,
         DP_OP_422J2_124_3477_n380, DP_OP_422J2_124_3477_n379,
         DP_OP_422J2_124_3477_n378, DP_OP_422J2_124_3477_n377,
         DP_OP_422J2_124_3477_n376, DP_OP_422J2_124_3477_n375,
         DP_OP_422J2_124_3477_n374, DP_OP_422J2_124_3477_n373,
         DP_OP_422J2_124_3477_n372, DP_OP_422J2_124_3477_n371,
         DP_OP_422J2_124_3477_n370, DP_OP_422J2_124_3477_n369,
         DP_OP_422J2_124_3477_n368, DP_OP_422J2_124_3477_n367,
         DP_OP_422J2_124_3477_n366, DP_OP_422J2_124_3477_n365,
         DP_OP_422J2_124_3477_n364, DP_OP_422J2_124_3477_n363,
         DP_OP_422J2_124_3477_n362, DP_OP_422J2_124_3477_n361,
         DP_OP_422J2_124_3477_n360, DP_OP_422J2_124_3477_n359,
         DP_OP_422J2_124_3477_n358, DP_OP_422J2_124_3477_n357,
         DP_OP_422J2_124_3477_n356, DP_OP_422J2_124_3477_n355,
         DP_OP_422J2_124_3477_n354, DP_OP_422J2_124_3477_n353,
         DP_OP_422J2_124_3477_n352, DP_OP_422J2_124_3477_n351,
         DP_OP_422J2_124_3477_n350, DP_OP_422J2_124_3477_n349,
         DP_OP_422J2_124_3477_n348, DP_OP_422J2_124_3477_n347,
         DP_OP_422J2_124_3477_n346, DP_OP_422J2_124_3477_n345,
         DP_OP_422J2_124_3477_n344, DP_OP_422J2_124_3477_n343,
         DP_OP_422J2_124_3477_n342, DP_OP_422J2_124_3477_n341,
         DP_OP_422J2_124_3477_n340, DP_OP_422J2_124_3477_n339,
         DP_OP_422J2_124_3477_n338, DP_OP_422J2_124_3477_n337,
         DP_OP_422J2_124_3477_n336, DP_OP_422J2_124_3477_n335,
         DP_OP_422J2_124_3477_n334, DP_OP_422J2_124_3477_n333,
         DP_OP_422J2_124_3477_n332, DP_OP_422J2_124_3477_n331,
         DP_OP_422J2_124_3477_n330, DP_OP_422J2_124_3477_n329,
         DP_OP_422J2_124_3477_n328, DP_OP_422J2_124_3477_n327,
         DP_OP_422J2_124_3477_n326, DP_OP_422J2_124_3477_n325,
         DP_OP_422J2_124_3477_n324, DP_OP_422J2_124_3477_n323,
         DP_OP_422J2_124_3477_n322, DP_OP_422J2_124_3477_n321,
         DP_OP_422J2_124_3477_n320, DP_OP_422J2_124_3477_n319,
         DP_OP_422J2_124_3477_n318, DP_OP_422J2_124_3477_n317,
         DP_OP_422J2_124_3477_n316, DP_OP_422J2_124_3477_n315,
         DP_OP_422J2_124_3477_n314, DP_OP_422J2_124_3477_n313,
         DP_OP_422J2_124_3477_n312, DP_OP_422J2_124_3477_n311,
         DP_OP_422J2_124_3477_n310, DP_OP_422J2_124_3477_n309,
         DP_OP_422J2_124_3477_n308, DP_OP_422J2_124_3477_n307,
         DP_OP_422J2_124_3477_n306, DP_OP_422J2_124_3477_n305,
         DP_OP_422J2_124_3477_n304, DP_OP_422J2_124_3477_n303,
         DP_OP_422J2_124_3477_n302, DP_OP_422J2_124_3477_n301,
         DP_OP_422J2_124_3477_n300, DP_OP_422J2_124_3477_n299,
         DP_OP_422J2_124_3477_n298, DP_OP_422J2_124_3477_n297,
         DP_OP_422J2_124_3477_n296, DP_OP_422J2_124_3477_n295,
         DP_OP_422J2_124_3477_n294, DP_OP_422J2_124_3477_n293,
         DP_OP_422J2_124_3477_n292, DP_OP_422J2_124_3477_n291,
         DP_OP_422J2_124_3477_n290, DP_OP_422J2_124_3477_n289,
         DP_OP_422J2_124_3477_n288, DP_OP_422J2_124_3477_n287,
         DP_OP_422J2_124_3477_n286, DP_OP_422J2_124_3477_n285,
         DP_OP_422J2_124_3477_n284, DP_OP_422J2_124_3477_n283,
         DP_OP_422J2_124_3477_n282, DP_OP_422J2_124_3477_n281,
         DP_OP_422J2_124_3477_n280, DP_OP_422J2_124_3477_n279,
         DP_OP_422J2_124_3477_n278, DP_OP_422J2_124_3477_n277,
         DP_OP_422J2_124_3477_n276, DP_OP_422J2_124_3477_n275,
         DP_OP_422J2_124_3477_n274, DP_OP_422J2_124_3477_n273,
         DP_OP_422J2_124_3477_n272, DP_OP_422J2_124_3477_n271,
         DP_OP_422J2_124_3477_n270, DP_OP_422J2_124_3477_n269,
         DP_OP_422J2_124_3477_n268, DP_OP_422J2_124_3477_n267,
         DP_OP_422J2_124_3477_n266, DP_OP_422J2_124_3477_n265,
         DP_OP_422J2_124_3477_n264, DP_OP_422J2_124_3477_n263,
         DP_OP_422J2_124_3477_n262, DP_OP_422J2_124_3477_n261,
         DP_OP_422J2_124_3477_n260, DP_OP_422J2_124_3477_n259,
         DP_OP_422J2_124_3477_n258, DP_OP_422J2_124_3477_n257,
         DP_OP_422J2_124_3477_n256, DP_OP_422J2_124_3477_n255,
         DP_OP_422J2_124_3477_n254, DP_OP_422J2_124_3477_n253,
         DP_OP_422J2_124_3477_n252, DP_OP_422J2_124_3477_n251,
         DP_OP_422J2_124_3477_n250, DP_OP_422J2_124_3477_n249,
         DP_OP_422J2_124_3477_n248, DP_OP_422J2_124_3477_n247,
         DP_OP_422J2_124_3477_n246, DP_OP_422J2_124_3477_n245,
         DP_OP_422J2_124_3477_n244, DP_OP_422J2_124_3477_n243,
         DP_OP_422J2_124_3477_n242, DP_OP_422J2_124_3477_n241,
         DP_OP_422J2_124_3477_n240, DP_OP_422J2_124_3477_n239,
         DP_OP_422J2_124_3477_n238, DP_OP_422J2_124_3477_n237,
         DP_OP_422J2_124_3477_n236, DP_OP_422J2_124_3477_n235,
         DP_OP_422J2_124_3477_n234, DP_OP_422J2_124_3477_n233,
         DP_OP_422J2_124_3477_n232, DP_OP_422J2_124_3477_n231,
         DP_OP_422J2_124_3477_n230, DP_OP_422J2_124_3477_n229,
         DP_OP_422J2_124_3477_n228, DP_OP_422J2_124_3477_n227,
         DP_OP_422J2_124_3477_n226, DP_OP_422J2_124_3477_n225,
         DP_OP_422J2_124_3477_n224, DP_OP_422J2_124_3477_n223,
         DP_OP_422J2_124_3477_n222, DP_OP_422J2_124_3477_n221,
         DP_OP_422J2_124_3477_n220, DP_OP_422J2_124_3477_n219,
         DP_OP_422J2_124_3477_n218, DP_OP_422J2_124_3477_n217,
         DP_OP_422J2_124_3477_n216, DP_OP_422J2_124_3477_n215,
         DP_OP_422J2_124_3477_n214, DP_OP_422J2_124_3477_n213,
         DP_OP_422J2_124_3477_n212, DP_OP_422J2_124_3477_n211,
         DP_OP_422J2_124_3477_n210, DP_OP_422J2_124_3477_n209,
         DP_OP_422J2_124_3477_n208, DP_OP_422J2_124_3477_n207,
         DP_OP_422J2_124_3477_n206, DP_OP_422J2_124_3477_n205,
         DP_OP_422J2_124_3477_n204, DP_OP_422J2_124_3477_n203,
         DP_OP_422J2_124_3477_n202, DP_OP_422J2_124_3477_n201,
         DP_OP_422J2_124_3477_n200, DP_OP_422J2_124_3477_n199,
         DP_OP_422J2_124_3477_n198, DP_OP_422J2_124_3477_n197,
         DP_OP_422J2_124_3477_n196, DP_OP_422J2_124_3477_n195,
         DP_OP_422J2_124_3477_n194, DP_OP_422J2_124_3477_n193,
         DP_OP_422J2_124_3477_n192, DP_OP_422J2_124_3477_n191,
         DP_OP_422J2_124_3477_n190, DP_OP_422J2_124_3477_n189,
         DP_OP_422J2_124_3477_n188, DP_OP_422J2_124_3477_n187,
         DP_OP_422J2_124_3477_n186, DP_OP_422J2_124_3477_n185,
         DP_OP_422J2_124_3477_n184, DP_OP_422J2_124_3477_n183,
         DP_OP_422J2_124_3477_n182, DP_OP_422J2_124_3477_n181,
         DP_OP_422J2_124_3477_n180, DP_OP_422J2_124_3477_n179,
         DP_OP_422J2_124_3477_n178, DP_OP_422J2_124_3477_n177,
         DP_OP_422J2_124_3477_n176, DP_OP_422J2_124_3477_n175,
         DP_OP_422J2_124_3477_n174, DP_OP_422J2_124_3477_n173,
         DP_OP_422J2_124_3477_n172, DP_OP_422J2_124_3477_n171,
         DP_OP_422J2_124_3477_n170, DP_OP_422J2_124_3477_n169,
         DP_OP_422J2_124_3477_n168, DP_OP_422J2_124_3477_n167,
         DP_OP_422J2_124_3477_n166, DP_OP_422J2_124_3477_n165,
         DP_OP_422J2_124_3477_n164, DP_OP_422J2_124_3477_n163,
         DP_OP_422J2_124_3477_n162, DP_OP_422J2_124_3477_n161,
         DP_OP_422J2_124_3477_n160, DP_OP_422J2_124_3477_n159,
         DP_OP_422J2_124_3477_n158, DP_OP_422J2_124_3477_n157,
         DP_OP_422J2_124_3477_n156, DP_OP_422J2_124_3477_n155,
         DP_OP_422J2_124_3477_n154, DP_OP_422J2_124_3477_n153,
         DP_OP_422J2_124_3477_n131, DP_OP_422J2_124_3477_n130,
         DP_OP_422J2_124_3477_n129, DP_OP_422J2_124_3477_n128,
         DP_OP_422J2_124_3477_n127, DP_OP_422J2_124_3477_n126,
         DP_OP_422J2_124_3477_n123, DP_OP_422J2_124_3477_n122,
         DP_OP_422J2_124_3477_n121, DP_OP_422J2_124_3477_n120,
         DP_OP_422J2_124_3477_n119, DP_OP_422J2_124_3477_n118,
         DP_OP_422J2_124_3477_n115, DP_OP_422J2_124_3477_n114,
         DP_OP_422J2_124_3477_n113, DP_OP_422J2_124_3477_n112,
         DP_OP_422J2_124_3477_n111, DP_OP_422J2_124_3477_n110,
         DP_OP_422J2_124_3477_n107, DP_OP_422J2_124_3477_n106,
         DP_OP_422J2_124_3477_n105, DP_OP_422J2_124_3477_n104,
         DP_OP_422J2_124_3477_n103, DP_OP_422J2_124_3477_n102,
         DP_OP_422J2_124_3477_n101, DP_OP_422J2_124_3477_n99,
         DP_OP_422J2_124_3477_n98, DP_OP_422J2_124_3477_n95,
         DP_OP_422J2_124_3477_n94, DP_OP_422J2_124_3477_n93,
         DP_OP_422J2_124_3477_n92, DP_OP_422J2_124_3477_n90,
         DP_OP_422J2_124_3477_n88, DP_OP_422J2_124_3477_n87,
         DP_OP_422J2_124_3477_n86, DP_OP_422J2_124_3477_n85,
         DP_OP_422J2_124_3477_n84, DP_OP_422J2_124_3477_n83,
         DP_OP_422J2_124_3477_n82, DP_OP_422J2_124_3477_n80,
         DP_OP_422J2_124_3477_n79, DP_OP_422J2_124_3477_n78,
         DP_OP_422J2_124_3477_n77, DP_OP_422J2_124_3477_n76,
         DP_OP_422J2_124_3477_n75, DP_OP_422J2_124_3477_n74,
         DP_OP_422J2_124_3477_n73, DP_OP_422J2_124_3477_n69,
         DP_OP_422J2_124_3477_n68, DP_OP_422J2_124_3477_n67,
         DP_OP_422J2_124_3477_n66, DP_OP_422J2_124_3477_n65,
         DP_OP_422J2_124_3477_n64, DP_OP_422J2_124_3477_n62,
         DP_OP_422J2_124_3477_n60, DP_OP_422J2_124_3477_n59,
         DP_OP_422J2_124_3477_n57, DP_OP_422J2_124_3477_n56,
         DP_OP_422J2_124_3477_n55, DP_OP_422J2_124_3477_n53,
         DP_OP_422J2_124_3477_n52, DP_OP_422J2_124_3477_n51,
         DP_OP_422J2_124_3477_n50, DP_OP_422J2_124_3477_n46,
         DP_OP_422J2_124_3477_n45, DP_OP_422J2_124_3477_n42,
         DP_OP_422J2_124_3477_n41, DP_OP_422J2_124_3477_n39,
         DP_OP_422J2_124_3477_n38, DP_OP_422J2_124_3477_n37,
         DP_OP_422J2_124_3477_n36, DP_OP_422J2_124_3477_n35,
         DP_OP_422J2_124_3477_n34, DP_OP_422J2_124_3477_n33,
         DP_OP_422J2_124_3477_n32, DP_OP_422J2_124_3477_n31,
         DP_OP_422J2_124_3477_n30, DP_OP_422J2_124_3477_n29,
         DP_OP_422J2_124_3477_n28, DP_OP_422J2_124_3477_n27,
         DP_OP_422J2_124_3477_n26, DP_OP_422J2_124_3477_n25,
         DP_OP_422J2_124_3477_n24, DP_OP_422J2_124_3477_n4,
         DP_OP_422J2_124_3477_n3, DP_OP_422J2_124_3477_n2,
         DP_OP_423J2_125_3477_n2913, DP_OP_423J2_125_3477_n2911,
         DP_OP_423J2_125_3477_n2910, DP_OP_423J2_125_3477_n2909,
         DP_OP_423J2_125_3477_n2908, DP_OP_423J2_125_3477_n2907,
         DP_OP_423J2_125_3477_n2906, DP_OP_423J2_125_3477_n2904,
         DP_OP_423J2_125_3477_n2903, DP_OP_423J2_125_3477_n2902,
         DP_OP_423J2_125_3477_n2901, DP_OP_423J2_125_3477_n2900,
         DP_OP_423J2_125_3477_n2899, DP_OP_423J2_125_3477_n2898,
         DP_OP_423J2_125_3477_n2897, DP_OP_423J2_125_3477_n2896,
         DP_OP_423J2_125_3477_n2895, DP_OP_423J2_125_3477_n2894,
         DP_OP_423J2_125_3477_n2893, DP_OP_423J2_125_3477_n2892,
         DP_OP_423J2_125_3477_n2891, DP_OP_423J2_125_3477_n2890,
         DP_OP_423J2_125_3477_n2889, DP_OP_423J2_125_3477_n2888,
         DP_OP_423J2_125_3477_n2887, DP_OP_423J2_125_3477_n2886,
         DP_OP_423J2_125_3477_n2885, DP_OP_423J2_125_3477_n2884,
         DP_OP_423J2_125_3477_n2883, DP_OP_423J2_125_3477_n2882,
         DP_OP_423J2_125_3477_n2881, DP_OP_423J2_125_3477_n2880,
         DP_OP_423J2_125_3477_n2879, DP_OP_423J2_125_3477_n2878,
         DP_OP_423J2_125_3477_n2877, DP_OP_423J2_125_3477_n2876,
         DP_OP_423J2_125_3477_n2875, DP_OP_423J2_125_3477_n2874,
         DP_OP_423J2_125_3477_n2873, DP_OP_423J2_125_3477_n2872,
         DP_OP_423J2_125_3477_n2871, DP_OP_423J2_125_3477_n2870,
         DP_OP_423J2_125_3477_n2869, DP_OP_423J2_125_3477_n2868,
         DP_OP_423J2_125_3477_n2867, DP_OP_423J2_125_3477_n2866,
         DP_OP_423J2_125_3477_n2865, DP_OP_423J2_125_3477_n2864,
         DP_OP_423J2_125_3477_n2861, DP_OP_423J2_125_3477_n2860,
         DP_OP_423J2_125_3477_n2859, DP_OP_423J2_125_3477_n2857,
         DP_OP_423J2_125_3477_n2856, DP_OP_423J2_125_3477_n2855,
         DP_OP_423J2_125_3477_n2854, DP_OP_423J2_125_3477_n2853,
         DP_OP_423J2_125_3477_n2852, DP_OP_423J2_125_3477_n2851,
         DP_OP_423J2_125_3477_n2850, DP_OP_423J2_125_3477_n2849,
         DP_OP_423J2_125_3477_n2848, DP_OP_423J2_125_3477_n2847,
         DP_OP_423J2_125_3477_n2846, DP_OP_423J2_125_3477_n2845,
         DP_OP_423J2_125_3477_n2844, DP_OP_423J2_125_3477_n2843,
         DP_OP_423J2_125_3477_n2842, DP_OP_423J2_125_3477_n2841,
         DP_OP_423J2_125_3477_n2840, DP_OP_423J2_125_3477_n2839,
         DP_OP_423J2_125_3477_n2838, DP_OP_423J2_125_3477_n2837,
         DP_OP_423J2_125_3477_n2836, DP_OP_423J2_125_3477_n2835,
         DP_OP_423J2_125_3477_n2834, DP_OP_423J2_125_3477_n2833,
         DP_OP_423J2_125_3477_n2832, DP_OP_423J2_125_3477_n2831,
         DP_OP_423J2_125_3477_n2830, DP_OP_423J2_125_3477_n2829,
         DP_OP_423J2_125_3477_n2828, DP_OP_423J2_125_3477_n2827,
         DP_OP_423J2_125_3477_n2826, DP_OP_423J2_125_3477_n2824,
         DP_OP_423J2_125_3477_n2823, DP_OP_423J2_125_3477_n2813,
         DP_OP_423J2_125_3477_n2812, DP_OP_423J2_125_3477_n2811,
         DP_OP_423J2_125_3477_n2810, DP_OP_423J2_125_3477_n2809,
         DP_OP_423J2_125_3477_n2808, DP_OP_423J2_125_3477_n2807,
         DP_OP_423J2_125_3477_n2806, DP_OP_423J2_125_3477_n2805,
         DP_OP_423J2_125_3477_n2804, DP_OP_423J2_125_3477_n2803,
         DP_OP_423J2_125_3477_n2802, DP_OP_423J2_125_3477_n2801,
         DP_OP_423J2_125_3477_n2800, DP_OP_423J2_125_3477_n2799,
         DP_OP_423J2_125_3477_n2798, DP_OP_423J2_125_3477_n2797,
         DP_OP_423J2_125_3477_n2796, DP_OP_423J2_125_3477_n2795,
         DP_OP_423J2_125_3477_n2794, DP_OP_423J2_125_3477_n2793,
         DP_OP_423J2_125_3477_n2792, DP_OP_423J2_125_3477_n2791,
         DP_OP_423J2_125_3477_n2790, DP_OP_423J2_125_3477_n2789,
         DP_OP_423J2_125_3477_n2788, DP_OP_423J2_125_3477_n2787,
         DP_OP_423J2_125_3477_n2786, DP_OP_423J2_125_3477_n2785,
         DP_OP_423J2_125_3477_n2784, DP_OP_423J2_125_3477_n2783,
         DP_OP_423J2_125_3477_n2782, DP_OP_423J2_125_3477_n2781,
         DP_OP_423J2_125_3477_n2779, DP_OP_423J2_125_3477_n2778,
         DP_OP_423J2_125_3477_n2777, DP_OP_423J2_125_3477_n2776,
         DP_OP_423J2_125_3477_n2775, DP_OP_423J2_125_3477_n2772,
         DP_OP_423J2_125_3477_n2770, DP_OP_423J2_125_3477_n2769,
         DP_OP_423J2_125_3477_n2768, DP_OP_423J2_125_3477_n2767,
         DP_OP_423J2_125_3477_n2766, DP_OP_423J2_125_3477_n2765,
         DP_OP_423J2_125_3477_n2764, DP_OP_423J2_125_3477_n2763,
         DP_OP_423J2_125_3477_n2762, DP_OP_423J2_125_3477_n2761,
         DP_OP_423J2_125_3477_n2760, DP_OP_423J2_125_3477_n2759,
         DP_OP_423J2_125_3477_n2758, DP_OP_423J2_125_3477_n2757,
         DP_OP_423J2_125_3477_n2756, DP_OP_423J2_125_3477_n2755,
         DP_OP_423J2_125_3477_n2754, DP_OP_423J2_125_3477_n2753,
         DP_OP_423J2_125_3477_n2752, DP_OP_423J2_125_3477_n2751,
         DP_OP_423J2_125_3477_n2750, DP_OP_423J2_125_3477_n2749,
         DP_OP_423J2_125_3477_n2748, DP_OP_423J2_125_3477_n2747,
         DP_OP_423J2_125_3477_n2746, DP_OP_423J2_125_3477_n2745,
         DP_OP_423J2_125_3477_n2744, DP_OP_423J2_125_3477_n2743,
         DP_OP_423J2_125_3477_n2742, DP_OP_423J2_125_3477_n2741,
         DP_OP_423J2_125_3477_n2740, DP_OP_423J2_125_3477_n2739,
         DP_OP_423J2_125_3477_n2738, DP_OP_423J2_125_3477_n2737,
         DP_OP_423J2_125_3477_n2734, DP_OP_423J2_125_3477_n2733,
         DP_OP_423J2_125_3477_n2732, DP_OP_423J2_125_3477_n2731,
         DP_OP_423J2_125_3477_n2730, DP_OP_423J2_125_3477_n2729,
         DP_OP_423J2_125_3477_n2726, DP_OP_423J2_125_3477_n2725,
         DP_OP_423J2_125_3477_n2724, DP_OP_423J2_125_3477_n2723,
         DP_OP_423J2_125_3477_n2722, DP_OP_423J2_125_3477_n2721,
         DP_OP_423J2_125_3477_n2720, DP_OP_423J2_125_3477_n2719,
         DP_OP_423J2_125_3477_n2718, DP_OP_423J2_125_3477_n2717,
         DP_OP_423J2_125_3477_n2716, DP_OP_423J2_125_3477_n2715,
         DP_OP_423J2_125_3477_n2714, DP_OP_423J2_125_3477_n2713,
         DP_OP_423J2_125_3477_n2712, DP_OP_423J2_125_3477_n2711,
         DP_OP_423J2_125_3477_n2710, DP_OP_423J2_125_3477_n2709,
         DP_OP_423J2_125_3477_n2708, DP_OP_423J2_125_3477_n2707,
         DP_OP_423J2_125_3477_n2706, DP_OP_423J2_125_3477_n2705,
         DP_OP_423J2_125_3477_n2704, DP_OP_423J2_125_3477_n2703,
         DP_OP_423J2_125_3477_n2702, DP_OP_423J2_125_3477_n2701,
         DP_OP_423J2_125_3477_n2700, DP_OP_423J2_125_3477_n2699,
         DP_OP_423J2_125_3477_n2698, DP_OP_423J2_125_3477_n2697,
         DP_OP_423J2_125_3477_n2696, DP_OP_423J2_125_3477_n2695,
         DP_OP_423J2_125_3477_n2693, DP_OP_423J2_125_3477_n2690,
         DP_OP_423J2_125_3477_n2688, DP_OP_423J2_125_3477_n2684,
         DP_OP_423J2_125_3477_n2683, DP_OP_423J2_125_3477_n2682,
         DP_OP_423J2_125_3477_n2681, DP_OP_423J2_125_3477_n2680,
         DP_OP_423J2_125_3477_n2679, DP_OP_423J2_125_3477_n2678,
         DP_OP_423J2_125_3477_n2677, DP_OP_423J2_125_3477_n2676,
         DP_OP_423J2_125_3477_n2675, DP_OP_423J2_125_3477_n2674,
         DP_OP_423J2_125_3477_n2673, DP_OP_423J2_125_3477_n2672,
         DP_OP_423J2_125_3477_n2671, DP_OP_423J2_125_3477_n2670,
         DP_OP_423J2_125_3477_n2669, DP_OP_423J2_125_3477_n2668,
         DP_OP_423J2_125_3477_n2667, DP_OP_423J2_125_3477_n2666,
         DP_OP_423J2_125_3477_n2665, DP_OP_423J2_125_3477_n2664,
         DP_OP_423J2_125_3477_n2663, DP_OP_423J2_125_3477_n2662,
         DP_OP_423J2_125_3477_n2661, DP_OP_423J2_125_3477_n2660,
         DP_OP_423J2_125_3477_n2659, DP_OP_423J2_125_3477_n2658,
         DP_OP_423J2_125_3477_n2657, DP_OP_423J2_125_3477_n2656,
         DP_OP_423J2_125_3477_n2655, DP_OP_423J2_125_3477_n2654,
         DP_OP_423J2_125_3477_n2653, DP_OP_423J2_125_3477_n2651,
         DP_OP_423J2_125_3477_n2649, DP_OP_423J2_125_3477_n2648,
         DP_OP_423J2_125_3477_n2647, DP_OP_423J2_125_3477_n2646,
         DP_OP_423J2_125_3477_n2645, DP_OP_423J2_125_3477_n2643,
         DP_OP_423J2_125_3477_n2642, DP_OP_423J2_125_3477_n2640,
         DP_OP_423J2_125_3477_n2639, DP_OP_423J2_125_3477_n2638,
         DP_OP_423J2_125_3477_n2637, DP_OP_423J2_125_3477_n2636,
         DP_OP_423J2_125_3477_n2635, DP_OP_423J2_125_3477_n2634,
         DP_OP_423J2_125_3477_n2633, DP_OP_423J2_125_3477_n2632,
         DP_OP_423J2_125_3477_n2631, DP_OP_423J2_125_3477_n2630,
         DP_OP_423J2_125_3477_n2629, DP_OP_423J2_125_3477_n2628,
         DP_OP_423J2_125_3477_n2627, DP_OP_423J2_125_3477_n2626,
         DP_OP_423J2_125_3477_n2625, DP_OP_423J2_125_3477_n2624,
         DP_OP_423J2_125_3477_n2623, DP_OP_423J2_125_3477_n2622,
         DP_OP_423J2_125_3477_n2621, DP_OP_423J2_125_3477_n2620,
         DP_OP_423J2_125_3477_n2619, DP_OP_423J2_125_3477_n2618,
         DP_OP_423J2_125_3477_n2617, DP_OP_423J2_125_3477_n2616,
         DP_OP_423J2_125_3477_n2615, DP_OP_423J2_125_3477_n2614,
         DP_OP_423J2_125_3477_n2613, DP_OP_423J2_125_3477_n2612,
         DP_OP_423J2_125_3477_n2611, DP_OP_423J2_125_3477_n2610,
         DP_OP_423J2_125_3477_n2609, DP_OP_423J2_125_3477_n2607,
         DP_OP_423J2_125_3477_n2605, DP_OP_423J2_125_3477_n2604,
         DP_OP_423J2_125_3477_n2603, DP_OP_423J2_125_3477_n2602,
         DP_OP_423J2_125_3477_n2601, DP_OP_423J2_125_3477_n2600,
         DP_OP_423J2_125_3477_n2599, DP_OP_423J2_125_3477_n2596,
         DP_OP_423J2_125_3477_n2595, DP_OP_423J2_125_3477_n2594,
         DP_OP_423J2_125_3477_n2593, DP_OP_423J2_125_3477_n2592,
         DP_OP_423J2_125_3477_n2591, DP_OP_423J2_125_3477_n2590,
         DP_OP_423J2_125_3477_n2589, DP_OP_423J2_125_3477_n2588,
         DP_OP_423J2_125_3477_n2587, DP_OP_423J2_125_3477_n2586,
         DP_OP_423J2_125_3477_n2585, DP_OP_423J2_125_3477_n2584,
         DP_OP_423J2_125_3477_n2583, DP_OP_423J2_125_3477_n2582,
         DP_OP_423J2_125_3477_n2581, DP_OP_423J2_125_3477_n2580,
         DP_OP_423J2_125_3477_n2579, DP_OP_423J2_125_3477_n2578,
         DP_OP_423J2_125_3477_n2577, DP_OP_423J2_125_3477_n2576,
         DP_OP_423J2_125_3477_n2575, DP_OP_423J2_125_3477_n2574,
         DP_OP_423J2_125_3477_n2573, DP_OP_423J2_125_3477_n2572,
         DP_OP_423J2_125_3477_n2571, DP_OP_423J2_125_3477_n2570,
         DP_OP_423J2_125_3477_n2569, DP_OP_423J2_125_3477_n2568,
         DP_OP_423J2_125_3477_n2567, DP_OP_423J2_125_3477_n2566,
         DP_OP_423J2_125_3477_n2565, DP_OP_423J2_125_3477_n2562,
         DP_OP_423J2_125_3477_n2561, DP_OP_423J2_125_3477_n2559,
         DP_OP_423J2_125_3477_n2558, DP_OP_423J2_125_3477_n2554,
         DP_OP_423J2_125_3477_n2553, DP_OP_423J2_125_3477_n2552,
         DP_OP_423J2_125_3477_n2551, DP_OP_423J2_125_3477_n2550,
         DP_OP_423J2_125_3477_n2549, DP_OP_423J2_125_3477_n2548,
         DP_OP_423J2_125_3477_n2547, DP_OP_423J2_125_3477_n2546,
         DP_OP_423J2_125_3477_n2545, DP_OP_423J2_125_3477_n2544,
         DP_OP_423J2_125_3477_n2543, DP_OP_423J2_125_3477_n2542,
         DP_OP_423J2_125_3477_n2541, DP_OP_423J2_125_3477_n2540,
         DP_OP_423J2_125_3477_n2539, DP_OP_423J2_125_3477_n2538,
         DP_OP_423J2_125_3477_n2537, DP_OP_423J2_125_3477_n2536,
         DP_OP_423J2_125_3477_n2535, DP_OP_423J2_125_3477_n2534,
         DP_OP_423J2_125_3477_n2533, DP_OP_423J2_125_3477_n2532,
         DP_OP_423J2_125_3477_n2531, DP_OP_423J2_125_3477_n2530,
         DP_OP_423J2_125_3477_n2529, DP_OP_423J2_125_3477_n2528,
         DP_OP_423J2_125_3477_n2527, DP_OP_423J2_125_3477_n2526,
         DP_OP_423J2_125_3477_n2525, DP_OP_423J2_125_3477_n2524,
         DP_OP_423J2_125_3477_n2523, DP_OP_423J2_125_3477_n2522,
         DP_OP_423J2_125_3477_n2521, DP_OP_423J2_125_3477_n2520,
         DP_OP_423J2_125_3477_n2519, DP_OP_423J2_125_3477_n2517,
         DP_OP_423J2_125_3477_n2516, DP_OP_423J2_125_3477_n2515,
         DP_OP_423J2_125_3477_n2510, DP_OP_423J2_125_3477_n2509,
         DP_OP_423J2_125_3477_n2508, DP_OP_423J2_125_3477_n2507,
         DP_OP_423J2_125_3477_n2506, DP_OP_423J2_125_3477_n2505,
         DP_OP_423J2_125_3477_n2504, DP_OP_423J2_125_3477_n2503,
         DP_OP_423J2_125_3477_n2502, DP_OP_423J2_125_3477_n2501,
         DP_OP_423J2_125_3477_n2500, DP_OP_423J2_125_3477_n2499,
         DP_OP_423J2_125_3477_n2498, DP_OP_423J2_125_3477_n2497,
         DP_OP_423J2_125_3477_n2496, DP_OP_423J2_125_3477_n2495,
         DP_OP_423J2_125_3477_n2494, DP_OP_423J2_125_3477_n2493,
         DP_OP_423J2_125_3477_n2492, DP_OP_423J2_125_3477_n2491,
         DP_OP_423J2_125_3477_n2490, DP_OP_423J2_125_3477_n2489,
         DP_OP_423J2_125_3477_n2488, DP_OP_423J2_125_3477_n2487,
         DP_OP_423J2_125_3477_n2486, DP_OP_423J2_125_3477_n2485,
         DP_OP_423J2_125_3477_n2484, DP_OP_423J2_125_3477_n2483,
         DP_OP_423J2_125_3477_n2482, DP_OP_423J2_125_3477_n2481,
         DP_OP_423J2_125_3477_n2480, DP_OP_423J2_125_3477_n2479,
         DP_OP_423J2_125_3477_n2478, DP_OP_423J2_125_3477_n2477,
         DP_OP_423J2_125_3477_n2476, DP_OP_423J2_125_3477_n2475,
         DP_OP_423J2_125_3477_n2474, DP_OP_423J2_125_3477_n2472,
         DP_OP_423J2_125_3477_n2471, DP_OP_423J2_125_3477_n2470,
         DP_OP_423J2_125_3477_n2469, DP_OP_423J2_125_3477_n2468,
         DP_OP_423J2_125_3477_n2467, DP_OP_423J2_125_3477_n2466,
         DP_OP_423J2_125_3477_n2465, DP_OP_423J2_125_3477_n2464,
         DP_OP_423J2_125_3477_n2463, DP_OP_423J2_125_3477_n2462,
         DP_OP_423J2_125_3477_n2461, DP_OP_423J2_125_3477_n2460,
         DP_OP_423J2_125_3477_n2459, DP_OP_423J2_125_3477_n2458,
         DP_OP_423J2_125_3477_n2457, DP_OP_423J2_125_3477_n2456,
         DP_OP_423J2_125_3477_n2455, DP_OP_423J2_125_3477_n2454,
         DP_OP_423J2_125_3477_n2453, DP_OP_423J2_125_3477_n2452,
         DP_OP_423J2_125_3477_n2451, DP_OP_423J2_125_3477_n2450,
         DP_OP_423J2_125_3477_n2449, DP_OP_423J2_125_3477_n2448,
         DP_OP_423J2_125_3477_n2447, DP_OP_423J2_125_3477_n2446,
         DP_OP_423J2_125_3477_n2445, DP_OP_423J2_125_3477_n2444,
         DP_OP_423J2_125_3477_n2443, DP_OP_423J2_125_3477_n2442,
         DP_OP_423J2_125_3477_n2441, DP_OP_423J2_125_3477_n2440,
         DP_OP_423J2_125_3477_n2439, DP_OP_423J2_125_3477_n2438,
         DP_OP_423J2_125_3477_n2437, DP_OP_423J2_125_3477_n2436,
         DP_OP_423J2_125_3477_n2435, DP_OP_423J2_125_3477_n2434,
         DP_OP_423J2_125_3477_n2433, DP_OP_423J2_125_3477_n2432,
         DP_OP_423J2_125_3477_n2431, DP_OP_423J2_125_3477_n2430,
         DP_OP_423J2_125_3477_n2429, DP_OP_423J2_125_3477_n2428,
         DP_OP_423J2_125_3477_n2425, DP_OP_423J2_125_3477_n2424,
         DP_OP_423J2_125_3477_n2421, DP_OP_423J2_125_3477_n2420,
         DP_OP_423J2_125_3477_n2419, DP_OP_423J2_125_3477_n2418,
         DP_OP_423J2_125_3477_n2417, DP_OP_423J2_125_3477_n2416,
         DP_OP_423J2_125_3477_n2415, DP_OP_423J2_125_3477_n2414,
         DP_OP_423J2_125_3477_n2413, DP_OP_423J2_125_3477_n2412,
         DP_OP_423J2_125_3477_n2411, DP_OP_423J2_125_3477_n2410,
         DP_OP_423J2_125_3477_n2409, DP_OP_423J2_125_3477_n2408,
         DP_OP_423J2_125_3477_n2407, DP_OP_423J2_125_3477_n2406,
         DP_OP_423J2_125_3477_n2405, DP_OP_423J2_125_3477_n2404,
         DP_OP_423J2_125_3477_n2403, DP_OP_423J2_125_3477_n2402,
         DP_OP_423J2_125_3477_n2401, DP_OP_423J2_125_3477_n2400,
         DP_OP_423J2_125_3477_n2399, DP_OP_423J2_125_3477_n2398,
         DP_OP_423J2_125_3477_n2397, DP_OP_423J2_125_3477_n2396,
         DP_OP_423J2_125_3477_n2395, DP_OP_423J2_125_3477_n2394,
         DP_OP_423J2_125_3477_n2393, DP_OP_423J2_125_3477_n2392,
         DP_OP_423J2_125_3477_n2391, DP_OP_423J2_125_3477_n2390,
         DP_OP_423J2_125_3477_n2389, DP_OP_423J2_125_3477_n2388,
         DP_OP_423J2_125_3477_n2387, DP_OP_423J2_125_3477_n2386,
         DP_OP_423J2_125_3477_n2377, DP_OP_423J2_125_3477_n2376,
         DP_OP_423J2_125_3477_n2375, DP_OP_423J2_125_3477_n2374,
         DP_OP_423J2_125_3477_n2373, DP_OP_423J2_125_3477_n2372,
         DP_OP_423J2_125_3477_n2371, DP_OP_423J2_125_3477_n2370,
         DP_OP_423J2_125_3477_n2369, DP_OP_423J2_125_3477_n2368,
         DP_OP_423J2_125_3477_n2367, DP_OP_423J2_125_3477_n2366,
         DP_OP_423J2_125_3477_n2365, DP_OP_423J2_125_3477_n2364,
         DP_OP_423J2_125_3477_n2363, DP_OP_423J2_125_3477_n2362,
         DP_OP_423J2_125_3477_n2361, DP_OP_423J2_125_3477_n2360,
         DP_OP_423J2_125_3477_n2359, DP_OP_423J2_125_3477_n2358,
         DP_OP_423J2_125_3477_n2357, DP_OP_423J2_125_3477_n2356,
         DP_OP_423J2_125_3477_n2355, DP_OP_423J2_125_3477_n2354,
         DP_OP_423J2_125_3477_n2353, DP_OP_423J2_125_3477_n2352,
         DP_OP_423J2_125_3477_n2351, DP_OP_423J2_125_3477_n2350,
         DP_OP_423J2_125_3477_n2349, DP_OP_423J2_125_3477_n2348,
         DP_OP_423J2_125_3477_n2347, DP_OP_423J2_125_3477_n2346,
         DP_OP_423J2_125_3477_n2345, DP_OP_423J2_125_3477_n2344,
         DP_OP_423J2_125_3477_n2343, DP_OP_423J2_125_3477_n2341,
         DP_OP_423J2_125_3477_n2339, DP_OP_423J2_125_3477_n2334,
         DP_OP_423J2_125_3477_n2333, DP_OP_423J2_125_3477_n2332,
         DP_OP_423J2_125_3477_n2331, DP_OP_423J2_125_3477_n2330,
         DP_OP_423J2_125_3477_n2329, DP_OP_423J2_125_3477_n2328,
         DP_OP_423J2_125_3477_n2327, DP_OP_423J2_125_3477_n2326,
         DP_OP_423J2_125_3477_n2325, DP_OP_423J2_125_3477_n2324,
         DP_OP_423J2_125_3477_n2323, DP_OP_423J2_125_3477_n2322,
         DP_OP_423J2_125_3477_n2321, DP_OP_423J2_125_3477_n2320,
         DP_OP_423J2_125_3477_n2319, DP_OP_423J2_125_3477_n2318,
         DP_OP_423J2_125_3477_n2317, DP_OP_423J2_125_3477_n2316,
         DP_OP_423J2_125_3477_n2315, DP_OP_423J2_125_3477_n2314,
         DP_OP_423J2_125_3477_n2313, DP_OP_423J2_125_3477_n2312,
         DP_OP_423J2_125_3477_n2311, DP_OP_423J2_125_3477_n2310,
         DP_OP_423J2_125_3477_n2309, DP_OP_423J2_125_3477_n2308,
         DP_OP_423J2_125_3477_n2307, DP_OP_423J2_125_3477_n2306,
         DP_OP_423J2_125_3477_n2305, DP_OP_423J2_125_3477_n2304,
         DP_OP_423J2_125_3477_n2303, DP_OP_423J2_125_3477_n2302,
         DP_OP_423J2_125_3477_n2301, DP_OP_423J2_125_3477_n2299,
         DP_OP_423J2_125_3477_n2298, DP_OP_423J2_125_3477_n2295,
         DP_OP_423J2_125_3477_n2294, DP_OP_423J2_125_3477_n2291,
         DP_OP_423J2_125_3477_n2288, DP_OP_423J2_125_3477_n2287,
         DP_OP_423J2_125_3477_n2286, DP_OP_423J2_125_3477_n2285,
         DP_OP_423J2_125_3477_n2284, DP_OP_423J2_125_3477_n2283,
         DP_OP_423J2_125_3477_n2282, DP_OP_423J2_125_3477_n2281,
         DP_OP_423J2_125_3477_n2280, DP_OP_423J2_125_3477_n2279,
         DP_OP_423J2_125_3477_n2278, DP_OP_423J2_125_3477_n2277,
         DP_OP_423J2_125_3477_n2276, DP_OP_423J2_125_3477_n2275,
         DP_OP_423J2_125_3477_n2274, DP_OP_423J2_125_3477_n2273,
         DP_OP_423J2_125_3477_n2272, DP_OP_423J2_125_3477_n2271,
         DP_OP_423J2_125_3477_n2270, DP_OP_423J2_125_3477_n2269,
         DP_OP_423J2_125_3477_n2268, DP_OP_423J2_125_3477_n2267,
         DP_OP_423J2_125_3477_n2266, DP_OP_423J2_125_3477_n2265,
         DP_OP_423J2_125_3477_n2264, DP_OP_423J2_125_3477_n2263,
         DP_OP_423J2_125_3477_n2262, DP_OP_423J2_125_3477_n2261,
         DP_OP_423J2_125_3477_n2260, DP_OP_423J2_125_3477_n2259,
         DP_OP_423J2_125_3477_n2258, DP_OP_423J2_125_3477_n2257,
         DP_OP_423J2_125_3477_n2256, DP_OP_423J2_125_3477_n2254,
         DP_OP_423J2_125_3477_n2251, DP_OP_423J2_125_3477_n2247,
         DP_OP_423J2_125_3477_n2244, DP_OP_423J2_125_3477_n2243,
         DP_OP_423J2_125_3477_n2242, DP_OP_423J2_125_3477_n2241,
         DP_OP_423J2_125_3477_n2240, DP_OP_423J2_125_3477_n2239,
         DP_OP_423J2_125_3477_n2238, DP_OP_423J2_125_3477_n2237,
         DP_OP_423J2_125_3477_n2236, DP_OP_423J2_125_3477_n2235,
         DP_OP_423J2_125_3477_n2234, DP_OP_423J2_125_3477_n2233,
         DP_OP_423J2_125_3477_n2232, DP_OP_423J2_125_3477_n2231,
         DP_OP_423J2_125_3477_n2230, DP_OP_423J2_125_3477_n2229,
         DP_OP_423J2_125_3477_n2228, DP_OP_423J2_125_3477_n2227,
         DP_OP_423J2_125_3477_n2226, DP_OP_423J2_125_3477_n2225,
         DP_OP_423J2_125_3477_n2224, DP_OP_423J2_125_3477_n2223,
         DP_OP_423J2_125_3477_n2222, DP_OP_423J2_125_3477_n2221,
         DP_OP_423J2_125_3477_n2220, DP_OP_423J2_125_3477_n2219,
         DP_OP_423J2_125_3477_n2218, DP_OP_423J2_125_3477_n2217,
         DP_OP_423J2_125_3477_n2216, DP_OP_423J2_125_3477_n2215,
         DP_OP_423J2_125_3477_n2214, DP_OP_423J2_125_3477_n2213,
         DP_OP_423J2_125_3477_n2212, DP_OP_423J2_125_3477_n2211,
         DP_OP_423J2_125_3477_n2209, DP_OP_423J2_125_3477_n2205,
         DP_OP_423J2_125_3477_n2204, DP_OP_423J2_125_3477_n2200,
         DP_OP_423J2_125_3477_n2199, DP_OP_423J2_125_3477_n2198,
         DP_OP_423J2_125_3477_n2197, DP_OP_423J2_125_3477_n2196,
         DP_OP_423J2_125_3477_n2195, DP_OP_423J2_125_3477_n2194,
         DP_OP_423J2_125_3477_n2193, DP_OP_423J2_125_3477_n2192,
         DP_OP_423J2_125_3477_n2191, DP_OP_423J2_125_3477_n2190,
         DP_OP_423J2_125_3477_n2189, DP_OP_423J2_125_3477_n2188,
         DP_OP_423J2_125_3477_n2187, DP_OP_423J2_125_3477_n2186,
         DP_OP_423J2_125_3477_n2185, DP_OP_423J2_125_3477_n2184,
         DP_OP_423J2_125_3477_n2183, DP_OP_423J2_125_3477_n2182,
         DP_OP_423J2_125_3477_n2181, DP_OP_423J2_125_3477_n2180,
         DP_OP_423J2_125_3477_n2179, DP_OP_423J2_125_3477_n2178,
         DP_OP_423J2_125_3477_n2177, DP_OP_423J2_125_3477_n2176,
         DP_OP_423J2_125_3477_n2175, DP_OP_423J2_125_3477_n2174,
         DP_OP_423J2_125_3477_n2173, DP_OP_423J2_125_3477_n2172,
         DP_OP_423J2_125_3477_n2171, DP_OP_423J2_125_3477_n2170,
         DP_OP_423J2_125_3477_n2169, DP_OP_423J2_125_3477_n2168,
         DP_OP_423J2_125_3477_n2167, DP_OP_423J2_125_3477_n2165,
         DP_OP_423J2_125_3477_n2164, DP_OP_423J2_125_3477_n2163,
         DP_OP_423J2_125_3477_n2161, DP_OP_423J2_125_3477_n2160,
         DP_OP_423J2_125_3477_n2158, DP_OP_423J2_125_3477_n2157,
         DP_OP_423J2_125_3477_n2156, DP_OP_423J2_125_3477_n2155,
         DP_OP_423J2_125_3477_n2154, DP_OP_423J2_125_3477_n2153,
         DP_OP_423J2_125_3477_n2152, DP_OP_423J2_125_3477_n2151,
         DP_OP_423J2_125_3477_n2150, DP_OP_423J2_125_3477_n2149,
         DP_OP_423J2_125_3477_n2148, DP_OP_423J2_125_3477_n2147,
         DP_OP_423J2_125_3477_n2146, DP_OP_423J2_125_3477_n2145,
         DP_OP_423J2_125_3477_n2144, DP_OP_423J2_125_3477_n2143,
         DP_OP_423J2_125_3477_n2142, DP_OP_423J2_125_3477_n2141,
         DP_OP_423J2_125_3477_n2140, DP_OP_423J2_125_3477_n2139,
         DP_OP_423J2_125_3477_n2138, DP_OP_423J2_125_3477_n2137,
         DP_OP_423J2_125_3477_n2136, DP_OP_423J2_125_3477_n2135,
         DP_OP_423J2_125_3477_n2134, DP_OP_423J2_125_3477_n2133,
         DP_OP_423J2_125_3477_n2132, DP_OP_423J2_125_3477_n2131,
         DP_OP_423J2_125_3477_n2130, DP_OP_423J2_125_3477_n2129,
         DP_OP_423J2_125_3477_n2128, DP_OP_423J2_125_3477_n2127,
         DP_OP_423J2_125_3477_n2126, DP_OP_423J2_125_3477_n2125,
         DP_OP_423J2_125_3477_n2122, DP_OP_423J2_125_3477_n2117,
         DP_OP_423J2_125_3477_n2116, DP_OP_423J2_125_3477_n2115,
         DP_OP_423J2_125_3477_n2114, DP_OP_423J2_125_3477_n2112,
         DP_OP_423J2_125_3477_n2111, DP_OP_423J2_125_3477_n2110,
         DP_OP_423J2_125_3477_n2109, DP_OP_423J2_125_3477_n2108,
         DP_OP_423J2_125_3477_n2107, DP_OP_423J2_125_3477_n2106,
         DP_OP_423J2_125_3477_n2105, DP_OP_423J2_125_3477_n2104,
         DP_OP_423J2_125_3477_n2103, DP_OP_423J2_125_3477_n2102,
         DP_OP_423J2_125_3477_n2101, DP_OP_423J2_125_3477_n2100,
         DP_OP_423J2_125_3477_n2099, DP_OP_423J2_125_3477_n2098,
         DP_OP_423J2_125_3477_n2097, DP_OP_423J2_125_3477_n2096,
         DP_OP_423J2_125_3477_n2095, DP_OP_423J2_125_3477_n2094,
         DP_OP_423J2_125_3477_n2093, DP_OP_423J2_125_3477_n2092,
         DP_OP_423J2_125_3477_n2091, DP_OP_423J2_125_3477_n2090,
         DP_OP_423J2_125_3477_n2089, DP_OP_423J2_125_3477_n2088,
         DP_OP_423J2_125_3477_n2087, DP_OP_423J2_125_3477_n2086,
         DP_OP_423J2_125_3477_n2085, DP_OP_423J2_125_3477_n2084,
         DP_OP_423J2_125_3477_n2083, DP_OP_423J2_125_3477_n2082,
         DP_OP_423J2_125_3477_n2081, DP_OP_423J2_125_3477_n2080,
         DP_OP_423J2_125_3477_n2077, DP_OP_423J2_125_3477_n2076,
         DP_OP_423J2_125_3477_n2074, DP_OP_423J2_125_3477_n2073,
         DP_OP_423J2_125_3477_n2068, DP_OP_423J2_125_3477_n2067,
         DP_OP_423J2_125_3477_n2066, DP_OP_423J2_125_3477_n2065,
         DP_OP_423J2_125_3477_n2064, DP_OP_423J2_125_3477_n2063,
         DP_OP_423J2_125_3477_n2062, DP_OP_423J2_125_3477_n2061,
         DP_OP_423J2_125_3477_n2060, DP_OP_423J2_125_3477_n2059,
         DP_OP_423J2_125_3477_n2058, DP_OP_423J2_125_3477_n2057,
         DP_OP_423J2_125_3477_n2056, DP_OP_423J2_125_3477_n2055,
         DP_OP_423J2_125_3477_n2054, DP_OP_423J2_125_3477_n2053,
         DP_OP_423J2_125_3477_n2052, DP_OP_423J2_125_3477_n2051,
         DP_OP_423J2_125_3477_n2050, DP_OP_423J2_125_3477_n2049,
         DP_OP_423J2_125_3477_n2048, DP_OP_423J2_125_3477_n2047,
         DP_OP_423J2_125_3477_n2046, DP_OP_423J2_125_3477_n2045,
         DP_OP_423J2_125_3477_n2044, DP_OP_423J2_125_3477_n2043,
         DP_OP_423J2_125_3477_n2042, DP_OP_423J2_125_3477_n2041,
         DP_OP_423J2_125_3477_n2040, DP_OP_423J2_125_3477_n2039,
         DP_OP_423J2_125_3477_n2038, DP_OP_423J2_125_3477_n2037,
         DP_OP_423J2_125_3477_n2034, DP_OP_423J2_125_3477_n2033,
         DP_OP_423J2_125_3477_n2032, DP_OP_423J2_125_3477_n2031,
         DP_OP_423J2_125_3477_n2030, DP_OP_423J2_125_3477_n2029,
         DP_OP_423J2_125_3477_n2028, DP_OP_423J2_125_3477_n2024,
         DP_OP_423J2_125_3477_n2023, DP_OP_423J2_125_3477_n2022,
         DP_OP_423J2_125_3477_n2021, DP_OP_423J2_125_3477_n2020,
         DP_OP_423J2_125_3477_n2019, DP_OP_423J2_125_3477_n2018,
         DP_OP_423J2_125_3477_n2017, DP_OP_423J2_125_3477_n2016,
         DP_OP_423J2_125_3477_n2015, DP_OP_423J2_125_3477_n2014,
         DP_OP_423J2_125_3477_n2013, DP_OP_423J2_125_3477_n2012,
         DP_OP_423J2_125_3477_n2011, DP_OP_423J2_125_3477_n2010,
         DP_OP_423J2_125_3477_n2009, DP_OP_423J2_125_3477_n2008,
         DP_OP_423J2_125_3477_n2007, DP_OP_423J2_125_3477_n2006,
         DP_OP_423J2_125_3477_n2005, DP_OP_423J2_125_3477_n2004,
         DP_OP_423J2_125_3477_n2003, DP_OP_423J2_125_3477_n2002,
         DP_OP_423J2_125_3477_n2001, DP_OP_423J2_125_3477_n2000,
         DP_OP_423J2_125_3477_n1999, DP_OP_423J2_125_3477_n1998,
         DP_OP_423J2_125_3477_n1997, DP_OP_423J2_125_3477_n1996,
         DP_OP_423J2_125_3477_n1995, DP_OP_423J2_125_3477_n1994,
         DP_OP_423J2_125_3477_n1993, DP_OP_423J2_125_3477_n1992,
         DP_OP_423J2_125_3477_n1991, DP_OP_423J2_125_3477_n1989,
         DP_OP_423J2_125_3477_n1986, DP_OP_423J2_125_3477_n1985,
         DP_OP_423J2_125_3477_n1983, DP_OP_423J2_125_3477_n1980,
         DP_OP_423J2_125_3477_n1979, DP_OP_423J2_125_3477_n1978,
         DP_OP_423J2_125_3477_n1977, DP_OP_423J2_125_3477_n1976,
         DP_OP_423J2_125_3477_n1975, DP_OP_423J2_125_3477_n1974,
         DP_OP_423J2_125_3477_n1973, DP_OP_423J2_125_3477_n1972,
         DP_OP_423J2_125_3477_n1971, DP_OP_423J2_125_3477_n1970,
         DP_OP_423J2_125_3477_n1969, DP_OP_423J2_125_3477_n1968,
         DP_OP_423J2_125_3477_n1967, DP_OP_423J2_125_3477_n1966,
         DP_OP_423J2_125_3477_n1965, DP_OP_423J2_125_3477_n1964,
         DP_OP_423J2_125_3477_n1963, DP_OP_423J2_125_3477_n1962,
         DP_OP_423J2_125_3477_n1961, DP_OP_423J2_125_3477_n1960,
         DP_OP_423J2_125_3477_n1959, DP_OP_423J2_125_3477_n1958,
         DP_OP_423J2_125_3477_n1957, DP_OP_423J2_125_3477_n1956,
         DP_OP_423J2_125_3477_n1955, DP_OP_423J2_125_3477_n1954,
         DP_OP_423J2_125_3477_n1953, DP_OP_423J2_125_3477_n1952,
         DP_OP_423J2_125_3477_n1951, DP_OP_423J2_125_3477_n1950,
         DP_OP_423J2_125_3477_n1949, DP_OP_423J2_125_3477_n1948,
         DP_OP_423J2_125_3477_n1947, DP_OP_423J2_125_3477_n1943,
         DP_OP_423J2_125_3477_n1939, DP_OP_423J2_125_3477_n1937,
         DP_OP_423J2_125_3477_n1936, DP_OP_423J2_125_3477_n1935,
         DP_OP_423J2_125_3477_n1934, DP_OP_423J2_125_3477_n1933,
         DP_OP_423J2_125_3477_n1932, DP_OP_423J2_125_3477_n1931,
         DP_OP_423J2_125_3477_n1930, DP_OP_423J2_125_3477_n1929,
         DP_OP_423J2_125_3477_n1928, DP_OP_423J2_125_3477_n1927,
         DP_OP_423J2_125_3477_n1926, DP_OP_423J2_125_3477_n1925,
         DP_OP_423J2_125_3477_n1924, DP_OP_423J2_125_3477_n1923,
         DP_OP_423J2_125_3477_n1922, DP_OP_423J2_125_3477_n1921,
         DP_OP_423J2_125_3477_n1920, DP_OP_423J2_125_3477_n1919,
         DP_OP_423J2_125_3477_n1918, DP_OP_423J2_125_3477_n1917,
         DP_OP_423J2_125_3477_n1916, DP_OP_423J2_125_3477_n1915,
         DP_OP_423J2_125_3477_n1914, DP_OP_423J2_125_3477_n1913,
         DP_OP_423J2_125_3477_n1912, DP_OP_423J2_125_3477_n1911,
         DP_OP_423J2_125_3477_n1910, DP_OP_423J2_125_3477_n1909,
         DP_OP_423J2_125_3477_n1908, DP_OP_423J2_125_3477_n1907,
         DP_OP_423J2_125_3477_n1906, DP_OP_423J2_125_3477_n1905,
         DP_OP_423J2_125_3477_n1904, DP_OP_423J2_125_3477_n1901,
         DP_OP_423J2_125_3477_n1899, DP_OP_423J2_125_3477_n1898,
         DP_OP_423J2_125_3477_n1897, DP_OP_423J2_125_3477_n1896,
         DP_OP_423J2_125_3477_n1893, DP_OP_423J2_125_3477_n1892,
         DP_OP_423J2_125_3477_n1891, DP_OP_423J2_125_3477_n1890,
         DP_OP_423J2_125_3477_n1889, DP_OP_423J2_125_3477_n1888,
         DP_OP_423J2_125_3477_n1887, DP_OP_423J2_125_3477_n1886,
         DP_OP_423J2_125_3477_n1885, DP_OP_423J2_125_3477_n1884,
         DP_OP_423J2_125_3477_n1883, DP_OP_423J2_125_3477_n1882,
         DP_OP_423J2_125_3477_n1881, DP_OP_423J2_125_3477_n1880,
         DP_OP_423J2_125_3477_n1879, DP_OP_423J2_125_3477_n1878,
         DP_OP_423J2_125_3477_n1877, DP_OP_423J2_125_3477_n1876,
         DP_OP_423J2_125_3477_n1875, DP_OP_423J2_125_3477_n1874,
         DP_OP_423J2_125_3477_n1873, DP_OP_423J2_125_3477_n1872,
         DP_OP_423J2_125_3477_n1871, DP_OP_423J2_125_3477_n1870,
         DP_OP_423J2_125_3477_n1869, DP_OP_423J2_125_3477_n1868,
         DP_OP_423J2_125_3477_n1867, DP_OP_423J2_125_3477_n1866,
         DP_OP_423J2_125_3477_n1865, DP_OP_423J2_125_3477_n1864,
         DP_OP_423J2_125_3477_n1863, DP_OP_423J2_125_3477_n1862,
         DP_OP_423J2_125_3477_n1861, DP_OP_423J2_125_3477_n1860,
         DP_OP_423J2_125_3477_n1859, DP_OP_423J2_125_3477_n1858,
         DP_OP_423J2_125_3477_n1856, DP_OP_423J2_125_3477_n1853,
         DP_OP_423J2_125_3477_n1852, DP_OP_423J2_125_3477_n1850,
         DP_OP_423J2_125_3477_n1849, DP_OP_423J2_125_3477_n1848,
         DP_OP_423J2_125_3477_n1847, DP_OP_423J2_125_3477_n1846,
         DP_OP_423J2_125_3477_n1845, DP_OP_423J2_125_3477_n1844,
         DP_OP_423J2_125_3477_n1843, DP_OP_423J2_125_3477_n1842,
         DP_OP_423J2_125_3477_n1841, DP_OP_423J2_125_3477_n1840,
         DP_OP_423J2_125_3477_n1839, DP_OP_423J2_125_3477_n1838,
         DP_OP_423J2_125_3477_n1837, DP_OP_423J2_125_3477_n1836,
         DP_OP_423J2_125_3477_n1835, DP_OP_423J2_125_3477_n1834,
         DP_OP_423J2_125_3477_n1833, DP_OP_423J2_125_3477_n1832,
         DP_OP_423J2_125_3477_n1831, DP_OP_423J2_125_3477_n1830,
         DP_OP_423J2_125_3477_n1829, DP_OP_423J2_125_3477_n1828,
         DP_OP_423J2_125_3477_n1827, DP_OP_423J2_125_3477_n1826,
         DP_OP_423J2_125_3477_n1825, DP_OP_423J2_125_3477_n1824,
         DP_OP_423J2_125_3477_n1823, DP_OP_423J2_125_3477_n1822,
         DP_OP_423J2_125_3477_n1821, DP_OP_423J2_125_3477_n1820,
         DP_OP_423J2_125_3477_n1819, DP_OP_423J2_125_3477_n1818,
         DP_OP_423J2_125_3477_n1817, DP_OP_423J2_125_3477_n1783,
         DP_OP_423J2_125_3477_n1782, DP_OP_423J2_125_3477_n1781,
         DP_OP_423J2_125_3477_n1780, DP_OP_423J2_125_3477_n1779,
         DP_OP_423J2_125_3477_n1778, DP_OP_423J2_125_3477_n1777,
         DP_OP_423J2_125_3477_n1776, DP_OP_423J2_125_3477_n1775,
         DP_OP_423J2_125_3477_n1774, DP_OP_423J2_125_3477_n1773,
         DP_OP_423J2_125_3477_n1772, DP_OP_423J2_125_3477_n1771,
         DP_OP_423J2_125_3477_n1770, DP_OP_423J2_125_3477_n1769,
         DP_OP_423J2_125_3477_n1768, DP_OP_423J2_125_3477_n1767,
         DP_OP_423J2_125_3477_n1766, DP_OP_423J2_125_3477_n1765,
         DP_OP_423J2_125_3477_n1764, DP_OP_423J2_125_3477_n1763,
         DP_OP_423J2_125_3477_n1762, DP_OP_423J2_125_3477_n1761,
         DP_OP_423J2_125_3477_n1760, DP_OP_423J2_125_3477_n1759,
         DP_OP_423J2_125_3477_n1758, DP_OP_423J2_125_3477_n1757,
         DP_OP_423J2_125_3477_n1756, DP_OP_423J2_125_3477_n1755,
         DP_OP_423J2_125_3477_n1754, DP_OP_423J2_125_3477_n1753,
         DP_OP_423J2_125_3477_n1752, DP_OP_423J2_125_3477_n1751,
         DP_OP_423J2_125_3477_n1750, DP_OP_423J2_125_3477_n1749,
         DP_OP_423J2_125_3477_n1748, DP_OP_423J2_125_3477_n1747,
         DP_OP_423J2_125_3477_n1746, DP_OP_423J2_125_3477_n1745,
         DP_OP_423J2_125_3477_n1744, DP_OP_423J2_125_3477_n1743,
         DP_OP_423J2_125_3477_n1742, DP_OP_423J2_125_3477_n1741,
         DP_OP_423J2_125_3477_n1740, DP_OP_423J2_125_3477_n1739,
         DP_OP_423J2_125_3477_n1738, DP_OP_423J2_125_3477_n1737,
         DP_OP_423J2_125_3477_n1736, DP_OP_423J2_125_3477_n1735,
         DP_OP_423J2_125_3477_n1734, DP_OP_423J2_125_3477_n1733,
         DP_OP_423J2_125_3477_n1732, DP_OP_423J2_125_3477_n1731,
         DP_OP_423J2_125_3477_n1730, DP_OP_423J2_125_3477_n1729,
         DP_OP_423J2_125_3477_n1728, DP_OP_423J2_125_3477_n1727,
         DP_OP_423J2_125_3477_n1726, DP_OP_423J2_125_3477_n1725,
         DP_OP_423J2_125_3477_n1724, DP_OP_423J2_125_3477_n1723,
         DP_OP_423J2_125_3477_n1722, DP_OP_423J2_125_3477_n1721,
         DP_OP_423J2_125_3477_n1720, DP_OP_423J2_125_3477_n1719,
         DP_OP_423J2_125_3477_n1718, DP_OP_423J2_125_3477_n1717,
         DP_OP_423J2_125_3477_n1716, DP_OP_423J2_125_3477_n1715,
         DP_OP_423J2_125_3477_n1714, DP_OP_423J2_125_3477_n1713,
         DP_OP_423J2_125_3477_n1712, DP_OP_423J2_125_3477_n1711,
         DP_OP_423J2_125_3477_n1710, DP_OP_423J2_125_3477_n1709,
         DP_OP_423J2_125_3477_n1708, DP_OP_423J2_125_3477_n1707,
         DP_OP_423J2_125_3477_n1706, DP_OP_423J2_125_3477_n1705,
         DP_OP_423J2_125_3477_n1704, DP_OP_423J2_125_3477_n1703,
         DP_OP_423J2_125_3477_n1702, DP_OP_423J2_125_3477_n1701,
         DP_OP_423J2_125_3477_n1700, DP_OP_423J2_125_3477_n1699,
         DP_OP_423J2_125_3477_n1698, DP_OP_423J2_125_3477_n1697,
         DP_OP_423J2_125_3477_n1696, DP_OP_423J2_125_3477_n1695,
         DP_OP_423J2_125_3477_n1694, DP_OP_423J2_125_3477_n1693,
         DP_OP_423J2_125_3477_n1692, DP_OP_423J2_125_3477_n1691,
         DP_OP_423J2_125_3477_n1690, DP_OP_423J2_125_3477_n1689,
         DP_OP_423J2_125_3477_n1688, DP_OP_423J2_125_3477_n1687,
         DP_OP_423J2_125_3477_n1686, DP_OP_423J2_125_3477_n1685,
         DP_OP_423J2_125_3477_n1684, DP_OP_423J2_125_3477_n1683,
         DP_OP_423J2_125_3477_n1682, DP_OP_423J2_125_3477_n1681,
         DP_OP_423J2_125_3477_n1680, DP_OP_423J2_125_3477_n1679,
         DP_OP_423J2_125_3477_n1678, DP_OP_423J2_125_3477_n1677,
         DP_OP_423J2_125_3477_n1676, DP_OP_423J2_125_3477_n1675,
         DP_OP_423J2_125_3477_n1674, DP_OP_423J2_125_3477_n1673,
         DP_OP_423J2_125_3477_n1672, DP_OP_423J2_125_3477_n1671,
         DP_OP_423J2_125_3477_n1670, DP_OP_423J2_125_3477_n1669,
         DP_OP_423J2_125_3477_n1668, DP_OP_423J2_125_3477_n1667,
         DP_OP_423J2_125_3477_n1666, DP_OP_423J2_125_3477_n1665,
         DP_OP_423J2_125_3477_n1664, DP_OP_423J2_125_3477_n1663,
         DP_OP_423J2_125_3477_n1662, DP_OP_423J2_125_3477_n1661,
         DP_OP_423J2_125_3477_n1660, DP_OP_423J2_125_3477_n1659,
         DP_OP_423J2_125_3477_n1658, DP_OP_423J2_125_3477_n1657,
         DP_OP_423J2_125_3477_n1656, DP_OP_423J2_125_3477_n1655,
         DP_OP_423J2_125_3477_n1654, DP_OP_423J2_125_3477_n1653,
         DP_OP_423J2_125_3477_n1652, DP_OP_423J2_125_3477_n1651,
         DP_OP_423J2_125_3477_n1650, DP_OP_423J2_125_3477_n1649,
         DP_OP_423J2_125_3477_n1648, DP_OP_423J2_125_3477_n1647,
         DP_OP_423J2_125_3477_n1646, DP_OP_423J2_125_3477_n1645,
         DP_OP_423J2_125_3477_n1644, DP_OP_423J2_125_3477_n1643,
         DP_OP_423J2_125_3477_n1642, DP_OP_423J2_125_3477_n1641,
         DP_OP_423J2_125_3477_n1640, DP_OP_423J2_125_3477_n1639,
         DP_OP_423J2_125_3477_n1638, DP_OP_423J2_125_3477_n1637,
         DP_OP_423J2_125_3477_n1636, DP_OP_423J2_125_3477_n1635,
         DP_OP_423J2_125_3477_n1634, DP_OP_423J2_125_3477_n1633,
         DP_OP_423J2_125_3477_n1632, DP_OP_423J2_125_3477_n1631,
         DP_OP_423J2_125_3477_n1630, DP_OP_423J2_125_3477_n1629,
         DP_OP_423J2_125_3477_n1628, DP_OP_423J2_125_3477_n1627,
         DP_OP_423J2_125_3477_n1626, DP_OP_423J2_125_3477_n1625,
         DP_OP_423J2_125_3477_n1624, DP_OP_423J2_125_3477_n1623,
         DP_OP_423J2_125_3477_n1622, DP_OP_423J2_125_3477_n1621,
         DP_OP_423J2_125_3477_n1620, DP_OP_423J2_125_3477_n1619,
         DP_OP_423J2_125_3477_n1618, DP_OP_423J2_125_3477_n1617,
         DP_OP_423J2_125_3477_n1616, DP_OP_423J2_125_3477_n1615,
         DP_OP_423J2_125_3477_n1614, DP_OP_423J2_125_3477_n1613,
         DP_OP_423J2_125_3477_n1612, DP_OP_423J2_125_3477_n1611,
         DP_OP_423J2_125_3477_n1610, DP_OP_423J2_125_3477_n1609,
         DP_OP_423J2_125_3477_n1608, DP_OP_423J2_125_3477_n1607,
         DP_OP_423J2_125_3477_n1606, DP_OP_423J2_125_3477_n1605,
         DP_OP_423J2_125_3477_n1604, DP_OP_423J2_125_3477_n1603,
         DP_OP_423J2_125_3477_n1602, DP_OP_423J2_125_3477_n1601,
         DP_OP_423J2_125_3477_n1600, DP_OP_423J2_125_3477_n1599,
         DP_OP_423J2_125_3477_n1598, DP_OP_423J2_125_3477_n1597,
         DP_OP_423J2_125_3477_n1596, DP_OP_423J2_125_3477_n1595,
         DP_OP_423J2_125_3477_n1594, DP_OP_423J2_125_3477_n1593,
         DP_OP_423J2_125_3477_n1592, DP_OP_423J2_125_3477_n1591,
         DP_OP_423J2_125_3477_n1590, DP_OP_423J2_125_3477_n1589,
         DP_OP_423J2_125_3477_n1588, DP_OP_423J2_125_3477_n1587,
         DP_OP_423J2_125_3477_n1586, DP_OP_423J2_125_3477_n1585,
         DP_OP_423J2_125_3477_n1584, DP_OP_423J2_125_3477_n1583,
         DP_OP_423J2_125_3477_n1582, DP_OP_423J2_125_3477_n1581,
         DP_OP_423J2_125_3477_n1580, DP_OP_423J2_125_3477_n1579,
         DP_OP_423J2_125_3477_n1578, DP_OP_423J2_125_3477_n1577,
         DP_OP_423J2_125_3477_n1576, DP_OP_423J2_125_3477_n1575,
         DP_OP_423J2_125_3477_n1574, DP_OP_423J2_125_3477_n1573,
         DP_OP_423J2_125_3477_n1572, DP_OP_423J2_125_3477_n1571,
         DP_OP_423J2_125_3477_n1570, DP_OP_423J2_125_3477_n1569,
         DP_OP_423J2_125_3477_n1568, DP_OP_423J2_125_3477_n1567,
         DP_OP_423J2_125_3477_n1566, DP_OP_423J2_125_3477_n1565,
         DP_OP_423J2_125_3477_n1564, DP_OP_423J2_125_3477_n1563,
         DP_OP_423J2_125_3477_n1562, DP_OP_423J2_125_3477_n1561,
         DP_OP_423J2_125_3477_n1560, DP_OP_423J2_125_3477_n1559,
         DP_OP_423J2_125_3477_n1558, DP_OP_423J2_125_3477_n1557,
         DP_OP_423J2_125_3477_n1556, DP_OP_423J2_125_3477_n1555,
         DP_OP_423J2_125_3477_n1554, DP_OP_423J2_125_3477_n1553,
         DP_OP_423J2_125_3477_n1552, DP_OP_423J2_125_3477_n1551,
         DP_OP_423J2_125_3477_n1550, DP_OP_423J2_125_3477_n1549,
         DP_OP_423J2_125_3477_n1548, DP_OP_423J2_125_3477_n1547,
         DP_OP_423J2_125_3477_n1546, DP_OP_423J2_125_3477_n1545,
         DP_OP_423J2_125_3477_n1544, DP_OP_423J2_125_3477_n1543,
         DP_OP_423J2_125_3477_n1542, DP_OP_423J2_125_3477_n1541,
         DP_OP_423J2_125_3477_n1540, DP_OP_423J2_125_3477_n1539,
         DP_OP_423J2_125_3477_n1538, DP_OP_423J2_125_3477_n1537,
         DP_OP_423J2_125_3477_n1536, DP_OP_423J2_125_3477_n1535,
         DP_OP_423J2_125_3477_n1534, DP_OP_423J2_125_3477_n1533,
         DP_OP_423J2_125_3477_n1532, DP_OP_423J2_125_3477_n1531,
         DP_OP_423J2_125_3477_n1530, DP_OP_423J2_125_3477_n1529,
         DP_OP_423J2_125_3477_n1528, DP_OP_423J2_125_3477_n1527,
         DP_OP_423J2_125_3477_n1526, DP_OP_423J2_125_3477_n1525,
         DP_OP_423J2_125_3477_n1524, DP_OP_423J2_125_3477_n1523,
         DP_OP_423J2_125_3477_n1522, DP_OP_423J2_125_3477_n1521,
         DP_OP_423J2_125_3477_n1520, DP_OP_423J2_125_3477_n1519,
         DP_OP_423J2_125_3477_n1518, DP_OP_423J2_125_3477_n1517,
         DP_OP_423J2_125_3477_n1516, DP_OP_423J2_125_3477_n1515,
         DP_OP_423J2_125_3477_n1514, DP_OP_423J2_125_3477_n1513,
         DP_OP_423J2_125_3477_n1512, DP_OP_423J2_125_3477_n1511,
         DP_OP_423J2_125_3477_n1510, DP_OP_423J2_125_3477_n1509,
         DP_OP_423J2_125_3477_n1508, DP_OP_423J2_125_3477_n1507,
         DP_OP_423J2_125_3477_n1506, DP_OP_423J2_125_3477_n1505,
         DP_OP_423J2_125_3477_n1504, DP_OP_423J2_125_3477_n1503,
         DP_OP_423J2_125_3477_n1502, DP_OP_423J2_125_3477_n1501,
         DP_OP_423J2_125_3477_n1500, DP_OP_423J2_125_3477_n1499,
         DP_OP_423J2_125_3477_n1498, DP_OP_423J2_125_3477_n1497,
         DP_OP_423J2_125_3477_n1496, DP_OP_423J2_125_3477_n1495,
         DP_OP_423J2_125_3477_n1494, DP_OP_423J2_125_3477_n1493,
         DP_OP_423J2_125_3477_n1492, DP_OP_423J2_125_3477_n1491,
         DP_OP_423J2_125_3477_n1490, DP_OP_423J2_125_3477_n1489,
         DP_OP_423J2_125_3477_n1488, DP_OP_423J2_125_3477_n1487,
         DP_OP_423J2_125_3477_n1486, DP_OP_423J2_125_3477_n1485,
         DP_OP_423J2_125_3477_n1484, DP_OP_423J2_125_3477_n1483,
         DP_OP_423J2_125_3477_n1482, DP_OP_423J2_125_3477_n1481,
         DP_OP_423J2_125_3477_n1480, DP_OP_423J2_125_3477_n1479,
         DP_OP_423J2_125_3477_n1478, DP_OP_423J2_125_3477_n1477,
         DP_OP_423J2_125_3477_n1476, DP_OP_423J2_125_3477_n1475,
         DP_OP_423J2_125_3477_n1474, DP_OP_423J2_125_3477_n1473,
         DP_OP_423J2_125_3477_n1472, DP_OP_423J2_125_3477_n1471,
         DP_OP_423J2_125_3477_n1470, DP_OP_423J2_125_3477_n1469,
         DP_OP_423J2_125_3477_n1468, DP_OP_423J2_125_3477_n1467,
         DP_OP_423J2_125_3477_n1466, DP_OP_423J2_125_3477_n1465,
         DP_OP_423J2_125_3477_n1464, DP_OP_423J2_125_3477_n1463,
         DP_OP_423J2_125_3477_n1462, DP_OP_423J2_125_3477_n1461,
         DP_OP_423J2_125_3477_n1460, DP_OP_423J2_125_3477_n1459,
         DP_OP_423J2_125_3477_n1458, DP_OP_423J2_125_3477_n1457,
         DP_OP_423J2_125_3477_n1456, DP_OP_423J2_125_3477_n1455,
         DP_OP_423J2_125_3477_n1454, DP_OP_423J2_125_3477_n1453,
         DP_OP_423J2_125_3477_n1452, DP_OP_423J2_125_3477_n1451,
         DP_OP_423J2_125_3477_n1450, DP_OP_423J2_125_3477_n1449,
         DP_OP_423J2_125_3477_n1448, DP_OP_423J2_125_3477_n1447,
         DP_OP_423J2_125_3477_n1446, DP_OP_423J2_125_3477_n1445,
         DP_OP_423J2_125_3477_n1444, DP_OP_423J2_125_3477_n1443,
         DP_OP_423J2_125_3477_n1442, DP_OP_423J2_125_3477_n1441,
         DP_OP_423J2_125_3477_n1440, DP_OP_423J2_125_3477_n1439,
         DP_OP_423J2_125_3477_n1438, DP_OP_423J2_125_3477_n1437,
         DP_OP_423J2_125_3477_n1436, DP_OP_423J2_125_3477_n1435,
         DP_OP_423J2_125_3477_n1434, DP_OP_423J2_125_3477_n1433,
         DP_OP_423J2_125_3477_n1432, DP_OP_423J2_125_3477_n1431,
         DP_OP_423J2_125_3477_n1430, DP_OP_423J2_125_3477_n1429,
         DP_OP_423J2_125_3477_n1428, DP_OP_423J2_125_3477_n1427,
         DP_OP_423J2_125_3477_n1426, DP_OP_423J2_125_3477_n1425,
         DP_OP_423J2_125_3477_n1424, DP_OP_423J2_125_3477_n1423,
         DP_OP_423J2_125_3477_n1422, DP_OP_423J2_125_3477_n1421,
         DP_OP_423J2_125_3477_n1420, DP_OP_423J2_125_3477_n1419,
         DP_OP_423J2_125_3477_n1418, DP_OP_423J2_125_3477_n1417,
         DP_OP_423J2_125_3477_n1416, DP_OP_423J2_125_3477_n1415,
         DP_OP_423J2_125_3477_n1414, DP_OP_423J2_125_3477_n1413,
         DP_OP_423J2_125_3477_n1412, DP_OP_423J2_125_3477_n1411,
         DP_OP_423J2_125_3477_n1410, DP_OP_423J2_125_3477_n1409,
         DP_OP_423J2_125_3477_n1408, DP_OP_423J2_125_3477_n1407,
         DP_OP_423J2_125_3477_n1406, DP_OP_423J2_125_3477_n1405,
         DP_OP_423J2_125_3477_n1404, DP_OP_423J2_125_3477_n1403,
         DP_OP_423J2_125_3477_n1402, DP_OP_423J2_125_3477_n1401,
         DP_OP_423J2_125_3477_n1400, DP_OP_423J2_125_3477_n1399,
         DP_OP_423J2_125_3477_n1398, DP_OP_423J2_125_3477_n1397,
         DP_OP_423J2_125_3477_n1396, DP_OP_423J2_125_3477_n1395,
         DP_OP_423J2_125_3477_n1394, DP_OP_423J2_125_3477_n1393,
         DP_OP_423J2_125_3477_n1392, DP_OP_423J2_125_3477_n1391,
         DP_OP_423J2_125_3477_n1390, DP_OP_423J2_125_3477_n1389,
         DP_OP_423J2_125_3477_n1388, DP_OP_423J2_125_3477_n1387,
         DP_OP_423J2_125_3477_n1386, DP_OP_423J2_125_3477_n1385,
         DP_OP_423J2_125_3477_n1384, DP_OP_423J2_125_3477_n1383,
         DP_OP_423J2_125_3477_n1382, DP_OP_423J2_125_3477_n1381,
         DP_OP_423J2_125_3477_n1380, DP_OP_423J2_125_3477_n1379,
         DP_OP_423J2_125_3477_n1378, DP_OP_423J2_125_3477_n1377,
         DP_OP_423J2_125_3477_n1376, DP_OP_423J2_125_3477_n1375,
         DP_OP_423J2_125_3477_n1374, DP_OP_423J2_125_3477_n1373,
         DP_OP_423J2_125_3477_n1372, DP_OP_423J2_125_3477_n1371,
         DP_OP_423J2_125_3477_n1370, DP_OP_423J2_125_3477_n1369,
         DP_OP_423J2_125_3477_n1368, DP_OP_423J2_125_3477_n1367,
         DP_OP_423J2_125_3477_n1366, DP_OP_423J2_125_3477_n1365,
         DP_OP_423J2_125_3477_n1364, DP_OP_423J2_125_3477_n1363,
         DP_OP_423J2_125_3477_n1362, DP_OP_423J2_125_3477_n1361,
         DP_OP_423J2_125_3477_n1360, DP_OP_423J2_125_3477_n1359,
         DP_OP_423J2_125_3477_n1358, DP_OP_423J2_125_3477_n1357,
         DP_OP_423J2_125_3477_n1356, DP_OP_423J2_125_3477_n1355,
         DP_OP_423J2_125_3477_n1354, DP_OP_423J2_125_3477_n1353,
         DP_OP_423J2_125_3477_n1352, DP_OP_423J2_125_3477_n1351,
         DP_OP_423J2_125_3477_n1350, DP_OP_423J2_125_3477_n1349,
         DP_OP_423J2_125_3477_n1348, DP_OP_423J2_125_3477_n1347,
         DP_OP_423J2_125_3477_n1346, DP_OP_423J2_125_3477_n1345,
         DP_OP_423J2_125_3477_n1344, DP_OP_423J2_125_3477_n1343,
         DP_OP_423J2_125_3477_n1342, DP_OP_423J2_125_3477_n1341,
         DP_OP_423J2_125_3477_n1340, DP_OP_423J2_125_3477_n1339,
         DP_OP_423J2_125_3477_n1338, DP_OP_423J2_125_3477_n1337,
         DP_OP_423J2_125_3477_n1336, DP_OP_423J2_125_3477_n1335,
         DP_OP_423J2_125_3477_n1334, DP_OP_423J2_125_3477_n1333,
         DP_OP_423J2_125_3477_n1332, DP_OP_423J2_125_3477_n1331,
         DP_OP_423J2_125_3477_n1330, DP_OP_423J2_125_3477_n1329,
         DP_OP_423J2_125_3477_n1328, DP_OP_423J2_125_3477_n1327,
         DP_OP_423J2_125_3477_n1326, DP_OP_423J2_125_3477_n1325,
         DP_OP_423J2_125_3477_n1324, DP_OP_423J2_125_3477_n1323,
         DP_OP_423J2_125_3477_n1322, DP_OP_423J2_125_3477_n1321,
         DP_OP_423J2_125_3477_n1320, DP_OP_423J2_125_3477_n1319,
         DP_OP_423J2_125_3477_n1318, DP_OP_423J2_125_3477_n1317,
         DP_OP_423J2_125_3477_n1316, DP_OP_423J2_125_3477_n1315,
         DP_OP_423J2_125_3477_n1314, DP_OP_423J2_125_3477_n1313,
         DP_OP_423J2_125_3477_n1312, DP_OP_423J2_125_3477_n1311,
         DP_OP_423J2_125_3477_n1310, DP_OP_423J2_125_3477_n1309,
         DP_OP_423J2_125_3477_n1308, DP_OP_423J2_125_3477_n1307,
         DP_OP_423J2_125_3477_n1306, DP_OP_423J2_125_3477_n1305,
         DP_OP_423J2_125_3477_n1304, DP_OP_423J2_125_3477_n1303,
         DP_OP_423J2_125_3477_n1302, DP_OP_423J2_125_3477_n1301,
         DP_OP_423J2_125_3477_n1300, DP_OP_423J2_125_3477_n1299,
         DP_OP_423J2_125_3477_n1298, DP_OP_423J2_125_3477_n1297,
         DP_OP_423J2_125_3477_n1296, DP_OP_423J2_125_3477_n1295,
         DP_OP_423J2_125_3477_n1294, DP_OP_423J2_125_3477_n1293,
         DP_OP_423J2_125_3477_n1292, DP_OP_423J2_125_3477_n1291,
         DP_OP_423J2_125_3477_n1290, DP_OP_423J2_125_3477_n1289,
         DP_OP_423J2_125_3477_n1288, DP_OP_423J2_125_3477_n1287,
         DP_OP_423J2_125_3477_n1286, DP_OP_423J2_125_3477_n1285,
         DP_OP_423J2_125_3477_n1284, DP_OP_423J2_125_3477_n1283,
         DP_OP_423J2_125_3477_n1282, DP_OP_423J2_125_3477_n1281,
         DP_OP_423J2_125_3477_n1280, DP_OP_423J2_125_3477_n1279,
         DP_OP_423J2_125_3477_n1278, DP_OP_423J2_125_3477_n1277,
         DP_OP_423J2_125_3477_n1276, DP_OP_423J2_125_3477_n1275,
         DP_OP_423J2_125_3477_n1274, DP_OP_423J2_125_3477_n1273,
         DP_OP_423J2_125_3477_n1272, DP_OP_423J2_125_3477_n1271,
         DP_OP_423J2_125_3477_n1270, DP_OP_423J2_125_3477_n1269,
         DP_OP_423J2_125_3477_n1268, DP_OP_423J2_125_3477_n1267,
         DP_OP_423J2_125_3477_n1266, DP_OP_423J2_125_3477_n1265,
         DP_OP_423J2_125_3477_n1264, DP_OP_423J2_125_3477_n1263,
         DP_OP_423J2_125_3477_n1262, DP_OP_423J2_125_3477_n1261,
         DP_OP_423J2_125_3477_n1260, DP_OP_423J2_125_3477_n1259,
         DP_OP_423J2_125_3477_n1258, DP_OP_423J2_125_3477_n1257,
         DP_OP_423J2_125_3477_n1256, DP_OP_423J2_125_3477_n1255,
         DP_OP_423J2_125_3477_n1254, DP_OP_423J2_125_3477_n1253,
         DP_OP_423J2_125_3477_n1252, DP_OP_423J2_125_3477_n1251,
         DP_OP_423J2_125_3477_n1250, DP_OP_423J2_125_3477_n1249,
         DP_OP_423J2_125_3477_n1248, DP_OP_423J2_125_3477_n1247,
         DP_OP_423J2_125_3477_n1246, DP_OP_423J2_125_3477_n1245,
         DP_OP_423J2_125_3477_n1244, DP_OP_423J2_125_3477_n1243,
         DP_OP_423J2_125_3477_n1242, DP_OP_423J2_125_3477_n1241,
         DP_OP_423J2_125_3477_n1240, DP_OP_423J2_125_3477_n1239,
         DP_OP_423J2_125_3477_n1238, DP_OP_423J2_125_3477_n1237,
         DP_OP_423J2_125_3477_n1236, DP_OP_423J2_125_3477_n1235,
         DP_OP_423J2_125_3477_n1234, DP_OP_423J2_125_3477_n1233,
         DP_OP_423J2_125_3477_n1232, DP_OP_423J2_125_3477_n1231,
         DP_OP_423J2_125_3477_n1230, DP_OP_423J2_125_3477_n1229,
         DP_OP_423J2_125_3477_n1228, DP_OP_423J2_125_3477_n1227,
         DP_OP_423J2_125_3477_n1226, DP_OP_423J2_125_3477_n1225,
         DP_OP_423J2_125_3477_n1224, DP_OP_423J2_125_3477_n1223,
         DP_OP_423J2_125_3477_n1222, DP_OP_423J2_125_3477_n1221,
         DP_OP_423J2_125_3477_n1220, DP_OP_423J2_125_3477_n1219,
         DP_OP_423J2_125_3477_n1218, DP_OP_423J2_125_3477_n1217,
         DP_OP_423J2_125_3477_n1216, DP_OP_423J2_125_3477_n1215,
         DP_OP_423J2_125_3477_n1214, DP_OP_423J2_125_3477_n1213,
         DP_OP_423J2_125_3477_n1212, DP_OP_423J2_125_3477_n1211,
         DP_OP_423J2_125_3477_n1210, DP_OP_423J2_125_3477_n1209,
         DP_OP_423J2_125_3477_n1208, DP_OP_423J2_125_3477_n1207,
         DP_OP_423J2_125_3477_n1206, DP_OP_423J2_125_3477_n1205,
         DP_OP_423J2_125_3477_n1204, DP_OP_423J2_125_3477_n1203,
         DP_OP_423J2_125_3477_n1202, DP_OP_423J2_125_3477_n1201,
         DP_OP_423J2_125_3477_n1200, DP_OP_423J2_125_3477_n1199,
         DP_OP_423J2_125_3477_n1198, DP_OP_423J2_125_3477_n1197,
         DP_OP_423J2_125_3477_n1196, DP_OP_423J2_125_3477_n1195,
         DP_OP_423J2_125_3477_n1194, DP_OP_423J2_125_3477_n1193,
         DP_OP_423J2_125_3477_n1192, DP_OP_423J2_125_3477_n1191,
         DP_OP_423J2_125_3477_n1190, DP_OP_423J2_125_3477_n1189,
         DP_OP_423J2_125_3477_n1188, DP_OP_423J2_125_3477_n1187,
         DP_OP_423J2_125_3477_n1186, DP_OP_423J2_125_3477_n1185,
         DP_OP_423J2_125_3477_n1184, DP_OP_423J2_125_3477_n1183,
         DP_OP_423J2_125_3477_n1182, DP_OP_423J2_125_3477_n1181,
         DP_OP_423J2_125_3477_n1180, DP_OP_423J2_125_3477_n1179,
         DP_OP_423J2_125_3477_n1178, DP_OP_423J2_125_3477_n1177,
         DP_OP_423J2_125_3477_n1176, DP_OP_423J2_125_3477_n1175,
         DP_OP_423J2_125_3477_n1174, DP_OP_423J2_125_3477_n1173,
         DP_OP_423J2_125_3477_n1172, DP_OP_423J2_125_3477_n1171,
         DP_OP_423J2_125_3477_n1170, DP_OP_423J2_125_3477_n1169,
         DP_OP_423J2_125_3477_n1168, DP_OP_423J2_125_3477_n1167,
         DP_OP_423J2_125_3477_n1166, DP_OP_423J2_125_3477_n1165,
         DP_OP_423J2_125_3477_n1164, DP_OP_423J2_125_3477_n1163,
         DP_OP_423J2_125_3477_n1162, DP_OP_423J2_125_3477_n1161,
         DP_OP_423J2_125_3477_n1160, DP_OP_423J2_125_3477_n1159,
         DP_OP_423J2_125_3477_n1158, DP_OP_423J2_125_3477_n1157,
         DP_OP_423J2_125_3477_n1156, DP_OP_423J2_125_3477_n1155,
         DP_OP_423J2_125_3477_n1154, DP_OP_423J2_125_3477_n1153,
         DP_OP_423J2_125_3477_n1152, DP_OP_423J2_125_3477_n1151,
         DP_OP_423J2_125_3477_n1150, DP_OP_423J2_125_3477_n1149,
         DP_OP_423J2_125_3477_n1148, DP_OP_423J2_125_3477_n1147,
         DP_OP_423J2_125_3477_n1146, DP_OP_423J2_125_3477_n1145,
         DP_OP_423J2_125_3477_n1144, DP_OP_423J2_125_3477_n1143,
         DP_OP_423J2_125_3477_n1142, DP_OP_423J2_125_3477_n1141,
         DP_OP_423J2_125_3477_n1140, DP_OP_423J2_125_3477_n1139,
         DP_OP_423J2_125_3477_n1138, DP_OP_423J2_125_3477_n1137,
         DP_OP_423J2_125_3477_n1136, DP_OP_423J2_125_3477_n1135,
         DP_OP_423J2_125_3477_n1134, DP_OP_423J2_125_3477_n1133,
         DP_OP_423J2_125_3477_n1132, DP_OP_423J2_125_3477_n1131,
         DP_OP_423J2_125_3477_n1130, DP_OP_423J2_125_3477_n1129,
         DP_OP_423J2_125_3477_n1128, DP_OP_423J2_125_3477_n1127,
         DP_OP_423J2_125_3477_n1126, DP_OP_423J2_125_3477_n1125,
         DP_OP_423J2_125_3477_n1124, DP_OP_423J2_125_3477_n1123,
         DP_OP_423J2_125_3477_n1122, DP_OP_423J2_125_3477_n1121,
         DP_OP_423J2_125_3477_n1120, DP_OP_423J2_125_3477_n1119,
         DP_OP_423J2_125_3477_n1118, DP_OP_423J2_125_3477_n1117,
         DP_OP_423J2_125_3477_n1116, DP_OP_423J2_125_3477_n1115,
         DP_OP_423J2_125_3477_n1114, DP_OP_423J2_125_3477_n1113,
         DP_OP_423J2_125_3477_n1112, DP_OP_423J2_125_3477_n1111,
         DP_OP_423J2_125_3477_n1110, DP_OP_423J2_125_3477_n1109,
         DP_OP_423J2_125_3477_n1108, DP_OP_423J2_125_3477_n1107,
         DP_OP_423J2_125_3477_n1106, DP_OP_423J2_125_3477_n1105,
         DP_OP_423J2_125_3477_n1104, DP_OP_423J2_125_3477_n1103,
         DP_OP_423J2_125_3477_n1102, DP_OP_423J2_125_3477_n1101,
         DP_OP_423J2_125_3477_n1100, DP_OP_423J2_125_3477_n1099,
         DP_OP_423J2_125_3477_n1098, DP_OP_423J2_125_3477_n1097,
         DP_OP_423J2_125_3477_n1096, DP_OP_423J2_125_3477_n1095,
         DP_OP_423J2_125_3477_n1094, DP_OP_423J2_125_3477_n1093,
         DP_OP_423J2_125_3477_n1092, DP_OP_423J2_125_3477_n1091,
         DP_OP_423J2_125_3477_n1090, DP_OP_423J2_125_3477_n1089,
         DP_OP_423J2_125_3477_n1088, DP_OP_423J2_125_3477_n1087,
         DP_OP_423J2_125_3477_n1086, DP_OP_423J2_125_3477_n1085,
         DP_OP_423J2_125_3477_n1084, DP_OP_423J2_125_3477_n1083,
         DP_OP_423J2_125_3477_n1082, DP_OP_423J2_125_3477_n1081,
         DP_OP_423J2_125_3477_n1080, DP_OP_423J2_125_3477_n1079,
         DP_OP_423J2_125_3477_n1078, DP_OP_423J2_125_3477_n1077,
         DP_OP_423J2_125_3477_n1076, DP_OP_423J2_125_3477_n1075,
         DP_OP_423J2_125_3477_n1074, DP_OP_423J2_125_3477_n1073,
         DP_OP_423J2_125_3477_n1072, DP_OP_423J2_125_3477_n1071,
         DP_OP_423J2_125_3477_n1070, DP_OP_423J2_125_3477_n1069,
         DP_OP_423J2_125_3477_n1068, DP_OP_423J2_125_3477_n1067,
         DP_OP_423J2_125_3477_n1066, DP_OP_423J2_125_3477_n1065,
         DP_OP_423J2_125_3477_n1064, DP_OP_423J2_125_3477_n1063,
         DP_OP_423J2_125_3477_n1062, DP_OP_423J2_125_3477_n1061,
         DP_OP_423J2_125_3477_n1060, DP_OP_423J2_125_3477_n1059,
         DP_OP_423J2_125_3477_n1058, DP_OP_423J2_125_3477_n1057,
         DP_OP_423J2_125_3477_n1056, DP_OP_423J2_125_3477_n1055,
         DP_OP_423J2_125_3477_n1054, DP_OP_423J2_125_3477_n1053,
         DP_OP_423J2_125_3477_n1052, DP_OP_423J2_125_3477_n1051,
         DP_OP_423J2_125_3477_n1050, DP_OP_423J2_125_3477_n1049,
         DP_OP_423J2_125_3477_n1048, DP_OP_423J2_125_3477_n1047,
         DP_OP_423J2_125_3477_n1046, DP_OP_423J2_125_3477_n1045,
         DP_OP_423J2_125_3477_n1044, DP_OP_423J2_125_3477_n1043,
         DP_OP_423J2_125_3477_n1042, DP_OP_423J2_125_3477_n1041,
         DP_OP_423J2_125_3477_n1040, DP_OP_423J2_125_3477_n1039,
         DP_OP_423J2_125_3477_n1038, DP_OP_423J2_125_3477_n1037,
         DP_OP_423J2_125_3477_n1036, DP_OP_423J2_125_3477_n1035,
         DP_OP_423J2_125_3477_n1034, DP_OP_423J2_125_3477_n1033,
         DP_OP_423J2_125_3477_n1032, DP_OP_423J2_125_3477_n1031,
         DP_OP_423J2_125_3477_n1030, DP_OP_423J2_125_3477_n1029,
         DP_OP_423J2_125_3477_n1028, DP_OP_423J2_125_3477_n1027,
         DP_OP_423J2_125_3477_n1026, DP_OP_423J2_125_3477_n1025,
         DP_OP_423J2_125_3477_n1024, DP_OP_423J2_125_3477_n1023,
         DP_OP_423J2_125_3477_n1022, DP_OP_423J2_125_3477_n1021,
         DP_OP_423J2_125_3477_n1020, DP_OP_423J2_125_3477_n1019,
         DP_OP_423J2_125_3477_n1018, DP_OP_423J2_125_3477_n1017,
         DP_OP_423J2_125_3477_n1016, DP_OP_423J2_125_3477_n1015,
         DP_OP_423J2_125_3477_n1014, DP_OP_423J2_125_3477_n1013,
         DP_OP_423J2_125_3477_n1012, DP_OP_423J2_125_3477_n1011,
         DP_OP_423J2_125_3477_n1010, DP_OP_423J2_125_3477_n1009,
         DP_OP_423J2_125_3477_n1008, DP_OP_423J2_125_3477_n1007,
         DP_OP_423J2_125_3477_n1006, DP_OP_423J2_125_3477_n1005,
         DP_OP_423J2_125_3477_n1004, DP_OP_423J2_125_3477_n1003,
         DP_OP_423J2_125_3477_n1002, DP_OP_423J2_125_3477_n1001,
         DP_OP_423J2_125_3477_n1000, DP_OP_423J2_125_3477_n999,
         DP_OP_423J2_125_3477_n998, DP_OP_423J2_125_3477_n997,
         DP_OP_423J2_125_3477_n996, DP_OP_423J2_125_3477_n995,
         DP_OP_423J2_125_3477_n994, DP_OP_423J2_125_3477_n993,
         DP_OP_423J2_125_3477_n992, DP_OP_423J2_125_3477_n991,
         DP_OP_423J2_125_3477_n990, DP_OP_423J2_125_3477_n989,
         DP_OP_423J2_125_3477_n988, DP_OP_423J2_125_3477_n987,
         DP_OP_423J2_125_3477_n986, DP_OP_423J2_125_3477_n985,
         DP_OP_423J2_125_3477_n984, DP_OP_423J2_125_3477_n983,
         DP_OP_423J2_125_3477_n982, DP_OP_423J2_125_3477_n981,
         DP_OP_423J2_125_3477_n980, DP_OP_423J2_125_3477_n979,
         DP_OP_423J2_125_3477_n978, DP_OP_423J2_125_3477_n977,
         DP_OP_423J2_125_3477_n976, DP_OP_423J2_125_3477_n975,
         DP_OP_423J2_125_3477_n974, DP_OP_423J2_125_3477_n973,
         DP_OP_423J2_125_3477_n972, DP_OP_423J2_125_3477_n971,
         DP_OP_423J2_125_3477_n970, DP_OP_423J2_125_3477_n969,
         DP_OP_423J2_125_3477_n968, DP_OP_423J2_125_3477_n967,
         DP_OP_423J2_125_3477_n966, DP_OP_423J2_125_3477_n965,
         DP_OP_423J2_125_3477_n964, DP_OP_423J2_125_3477_n963,
         DP_OP_423J2_125_3477_n962, DP_OP_423J2_125_3477_n961,
         DP_OP_423J2_125_3477_n960, DP_OP_423J2_125_3477_n959,
         DP_OP_423J2_125_3477_n958, DP_OP_423J2_125_3477_n957,
         DP_OP_423J2_125_3477_n956, DP_OP_423J2_125_3477_n955,
         DP_OP_423J2_125_3477_n954, DP_OP_423J2_125_3477_n953,
         DP_OP_423J2_125_3477_n952, DP_OP_423J2_125_3477_n951,
         DP_OP_423J2_125_3477_n950, DP_OP_423J2_125_3477_n949,
         DP_OP_423J2_125_3477_n948, DP_OP_423J2_125_3477_n947,
         DP_OP_423J2_125_3477_n946, DP_OP_423J2_125_3477_n945,
         DP_OP_423J2_125_3477_n944, DP_OP_423J2_125_3477_n943,
         DP_OP_423J2_125_3477_n942, DP_OP_423J2_125_3477_n941,
         DP_OP_423J2_125_3477_n940, DP_OP_423J2_125_3477_n939,
         DP_OP_423J2_125_3477_n938, DP_OP_423J2_125_3477_n937,
         DP_OP_423J2_125_3477_n936, DP_OP_423J2_125_3477_n935,
         DP_OP_423J2_125_3477_n934, DP_OP_423J2_125_3477_n933,
         DP_OP_423J2_125_3477_n932, DP_OP_423J2_125_3477_n931,
         DP_OP_423J2_125_3477_n930, DP_OP_423J2_125_3477_n929,
         DP_OP_423J2_125_3477_n928, DP_OP_423J2_125_3477_n927,
         DP_OP_423J2_125_3477_n926, DP_OP_423J2_125_3477_n925,
         DP_OP_423J2_125_3477_n924, DP_OP_423J2_125_3477_n923,
         DP_OP_423J2_125_3477_n922, DP_OP_423J2_125_3477_n921,
         DP_OP_423J2_125_3477_n920, DP_OP_423J2_125_3477_n919,
         DP_OP_423J2_125_3477_n918, DP_OP_423J2_125_3477_n917,
         DP_OP_423J2_125_3477_n916, DP_OP_423J2_125_3477_n915,
         DP_OP_423J2_125_3477_n914, DP_OP_423J2_125_3477_n913,
         DP_OP_423J2_125_3477_n912, DP_OP_423J2_125_3477_n911,
         DP_OP_423J2_125_3477_n910, DP_OP_423J2_125_3477_n909,
         DP_OP_423J2_125_3477_n908, DP_OP_423J2_125_3477_n907,
         DP_OP_423J2_125_3477_n906, DP_OP_423J2_125_3477_n905,
         DP_OP_423J2_125_3477_n904, DP_OP_423J2_125_3477_n903,
         DP_OP_423J2_125_3477_n902, DP_OP_423J2_125_3477_n901,
         DP_OP_423J2_125_3477_n900, DP_OP_423J2_125_3477_n899,
         DP_OP_423J2_125_3477_n898, DP_OP_423J2_125_3477_n897,
         DP_OP_423J2_125_3477_n896, DP_OP_423J2_125_3477_n895,
         DP_OP_423J2_125_3477_n894, DP_OP_423J2_125_3477_n893,
         DP_OP_423J2_125_3477_n892, DP_OP_423J2_125_3477_n891,
         DP_OP_423J2_125_3477_n890, DP_OP_423J2_125_3477_n889,
         DP_OP_423J2_125_3477_n888, DP_OP_423J2_125_3477_n887,
         DP_OP_423J2_125_3477_n886, DP_OP_423J2_125_3477_n885,
         DP_OP_423J2_125_3477_n884, DP_OP_423J2_125_3477_n883,
         DP_OP_423J2_125_3477_n882, DP_OP_423J2_125_3477_n881,
         DP_OP_423J2_125_3477_n880, DP_OP_423J2_125_3477_n879,
         DP_OP_423J2_125_3477_n878, DP_OP_423J2_125_3477_n877,
         DP_OP_423J2_125_3477_n876, DP_OP_423J2_125_3477_n875,
         DP_OP_423J2_125_3477_n874, DP_OP_423J2_125_3477_n873,
         DP_OP_423J2_125_3477_n872, DP_OP_423J2_125_3477_n871,
         DP_OP_423J2_125_3477_n870, DP_OP_423J2_125_3477_n869,
         DP_OP_423J2_125_3477_n868, DP_OP_423J2_125_3477_n867,
         DP_OP_423J2_125_3477_n866, DP_OP_423J2_125_3477_n865,
         DP_OP_423J2_125_3477_n864, DP_OP_423J2_125_3477_n863,
         DP_OP_423J2_125_3477_n862, DP_OP_423J2_125_3477_n861,
         DP_OP_423J2_125_3477_n860, DP_OP_423J2_125_3477_n859,
         DP_OP_423J2_125_3477_n858, DP_OP_423J2_125_3477_n857,
         DP_OP_423J2_125_3477_n856, DP_OP_423J2_125_3477_n855,
         DP_OP_423J2_125_3477_n854, DP_OP_423J2_125_3477_n853,
         DP_OP_423J2_125_3477_n852, DP_OP_423J2_125_3477_n851,
         DP_OP_423J2_125_3477_n850, DP_OP_423J2_125_3477_n849,
         DP_OP_423J2_125_3477_n848, DP_OP_423J2_125_3477_n847,
         DP_OP_423J2_125_3477_n846, DP_OP_423J2_125_3477_n845,
         DP_OP_423J2_125_3477_n844, DP_OP_423J2_125_3477_n843,
         DP_OP_423J2_125_3477_n842, DP_OP_423J2_125_3477_n841,
         DP_OP_423J2_125_3477_n840, DP_OP_423J2_125_3477_n839,
         DP_OP_423J2_125_3477_n838, DP_OP_423J2_125_3477_n837,
         DP_OP_423J2_125_3477_n836, DP_OP_423J2_125_3477_n835,
         DP_OP_423J2_125_3477_n834, DP_OP_423J2_125_3477_n833,
         DP_OP_423J2_125_3477_n832, DP_OP_423J2_125_3477_n831,
         DP_OP_423J2_125_3477_n830, DP_OP_423J2_125_3477_n829,
         DP_OP_423J2_125_3477_n828, DP_OP_423J2_125_3477_n827,
         DP_OP_423J2_125_3477_n826, DP_OP_423J2_125_3477_n825,
         DP_OP_423J2_125_3477_n824, DP_OP_423J2_125_3477_n823,
         DP_OP_423J2_125_3477_n822, DP_OP_423J2_125_3477_n821,
         DP_OP_423J2_125_3477_n820, DP_OP_423J2_125_3477_n819,
         DP_OP_423J2_125_3477_n818, DP_OP_423J2_125_3477_n817,
         DP_OP_423J2_125_3477_n816, DP_OP_423J2_125_3477_n815,
         DP_OP_423J2_125_3477_n814, DP_OP_423J2_125_3477_n813,
         DP_OP_423J2_125_3477_n812, DP_OP_423J2_125_3477_n811,
         DP_OP_423J2_125_3477_n810, DP_OP_423J2_125_3477_n809,
         DP_OP_423J2_125_3477_n808, DP_OP_423J2_125_3477_n807,
         DP_OP_423J2_125_3477_n806, DP_OP_423J2_125_3477_n805,
         DP_OP_423J2_125_3477_n804, DP_OP_423J2_125_3477_n803,
         DP_OP_423J2_125_3477_n802, DP_OP_423J2_125_3477_n801,
         DP_OP_423J2_125_3477_n800, DP_OP_423J2_125_3477_n799,
         DP_OP_423J2_125_3477_n798, DP_OP_423J2_125_3477_n797,
         DP_OP_423J2_125_3477_n796, DP_OP_423J2_125_3477_n795,
         DP_OP_423J2_125_3477_n794, DP_OP_423J2_125_3477_n793,
         DP_OP_423J2_125_3477_n792, DP_OP_423J2_125_3477_n791,
         DP_OP_423J2_125_3477_n790, DP_OP_423J2_125_3477_n789,
         DP_OP_423J2_125_3477_n788, DP_OP_423J2_125_3477_n787,
         DP_OP_423J2_125_3477_n786, DP_OP_423J2_125_3477_n785,
         DP_OP_423J2_125_3477_n784, DP_OP_423J2_125_3477_n783,
         DP_OP_423J2_125_3477_n782, DP_OP_423J2_125_3477_n781,
         DP_OP_423J2_125_3477_n780, DP_OP_423J2_125_3477_n779,
         DP_OP_423J2_125_3477_n778, DP_OP_423J2_125_3477_n777,
         DP_OP_423J2_125_3477_n776, DP_OP_423J2_125_3477_n775,
         DP_OP_423J2_125_3477_n774, DP_OP_423J2_125_3477_n773,
         DP_OP_423J2_125_3477_n772, DP_OP_423J2_125_3477_n771,
         DP_OP_423J2_125_3477_n770, DP_OP_423J2_125_3477_n769,
         DP_OP_423J2_125_3477_n768, DP_OP_423J2_125_3477_n767,
         DP_OP_423J2_125_3477_n766, DP_OP_423J2_125_3477_n765,
         DP_OP_423J2_125_3477_n764, DP_OP_423J2_125_3477_n763,
         DP_OP_423J2_125_3477_n762, DP_OP_423J2_125_3477_n761,
         DP_OP_423J2_125_3477_n760, DP_OP_423J2_125_3477_n759,
         DP_OP_423J2_125_3477_n758, DP_OP_423J2_125_3477_n757,
         DP_OP_423J2_125_3477_n756, DP_OP_423J2_125_3477_n755,
         DP_OP_423J2_125_3477_n754, DP_OP_423J2_125_3477_n753,
         DP_OP_423J2_125_3477_n752, DP_OP_423J2_125_3477_n751,
         DP_OP_423J2_125_3477_n750, DP_OP_423J2_125_3477_n749,
         DP_OP_423J2_125_3477_n748, DP_OP_423J2_125_3477_n747,
         DP_OP_423J2_125_3477_n746, DP_OP_423J2_125_3477_n745,
         DP_OP_423J2_125_3477_n744, DP_OP_423J2_125_3477_n743,
         DP_OP_423J2_125_3477_n742, DP_OP_423J2_125_3477_n741,
         DP_OP_423J2_125_3477_n740, DP_OP_423J2_125_3477_n739,
         DP_OP_423J2_125_3477_n738, DP_OP_423J2_125_3477_n737,
         DP_OP_423J2_125_3477_n736, DP_OP_423J2_125_3477_n735,
         DP_OP_423J2_125_3477_n734, DP_OP_423J2_125_3477_n733,
         DP_OP_423J2_125_3477_n732, DP_OP_423J2_125_3477_n731,
         DP_OP_423J2_125_3477_n730, DP_OP_423J2_125_3477_n729,
         DP_OP_423J2_125_3477_n728, DP_OP_423J2_125_3477_n727,
         DP_OP_423J2_125_3477_n726, DP_OP_423J2_125_3477_n725,
         DP_OP_423J2_125_3477_n724, DP_OP_423J2_125_3477_n723,
         DP_OP_423J2_125_3477_n722, DP_OP_423J2_125_3477_n721,
         DP_OP_423J2_125_3477_n720, DP_OP_423J2_125_3477_n719,
         DP_OP_423J2_125_3477_n718, DP_OP_423J2_125_3477_n717,
         DP_OP_423J2_125_3477_n716, DP_OP_423J2_125_3477_n715,
         DP_OP_423J2_125_3477_n714, DP_OP_423J2_125_3477_n713,
         DP_OP_423J2_125_3477_n712, DP_OP_423J2_125_3477_n711,
         DP_OP_423J2_125_3477_n710, DP_OP_423J2_125_3477_n709,
         DP_OP_423J2_125_3477_n708, DP_OP_423J2_125_3477_n707,
         DP_OP_423J2_125_3477_n706, DP_OP_423J2_125_3477_n705,
         DP_OP_423J2_125_3477_n704, DP_OP_423J2_125_3477_n703,
         DP_OP_423J2_125_3477_n702, DP_OP_423J2_125_3477_n701,
         DP_OP_423J2_125_3477_n700, DP_OP_423J2_125_3477_n699,
         DP_OP_423J2_125_3477_n698, DP_OP_423J2_125_3477_n697,
         DP_OP_423J2_125_3477_n696, DP_OP_423J2_125_3477_n695,
         DP_OP_423J2_125_3477_n694, DP_OP_423J2_125_3477_n693,
         DP_OP_423J2_125_3477_n692, DP_OP_423J2_125_3477_n691,
         DP_OP_423J2_125_3477_n690, DP_OP_423J2_125_3477_n689,
         DP_OP_423J2_125_3477_n688, DP_OP_423J2_125_3477_n687,
         DP_OP_423J2_125_3477_n686, DP_OP_423J2_125_3477_n685,
         DP_OP_423J2_125_3477_n684, DP_OP_423J2_125_3477_n683,
         DP_OP_423J2_125_3477_n682, DP_OP_423J2_125_3477_n681,
         DP_OP_423J2_125_3477_n680, DP_OP_423J2_125_3477_n679,
         DP_OP_423J2_125_3477_n678, DP_OP_423J2_125_3477_n677,
         DP_OP_423J2_125_3477_n676, DP_OP_423J2_125_3477_n675,
         DP_OP_423J2_125_3477_n674, DP_OP_423J2_125_3477_n673,
         DP_OP_423J2_125_3477_n672, DP_OP_423J2_125_3477_n671,
         DP_OP_423J2_125_3477_n670, DP_OP_423J2_125_3477_n669,
         DP_OP_423J2_125_3477_n668, DP_OP_423J2_125_3477_n667,
         DP_OP_423J2_125_3477_n666, DP_OP_423J2_125_3477_n665,
         DP_OP_423J2_125_3477_n664, DP_OP_423J2_125_3477_n663,
         DP_OP_423J2_125_3477_n662, DP_OP_423J2_125_3477_n661,
         DP_OP_423J2_125_3477_n660, DP_OP_423J2_125_3477_n659,
         DP_OP_423J2_125_3477_n658, DP_OP_423J2_125_3477_n657,
         DP_OP_423J2_125_3477_n656, DP_OP_423J2_125_3477_n655,
         DP_OP_423J2_125_3477_n654, DP_OP_423J2_125_3477_n653,
         DP_OP_423J2_125_3477_n652, DP_OP_423J2_125_3477_n651,
         DP_OP_423J2_125_3477_n650, DP_OP_423J2_125_3477_n649,
         DP_OP_423J2_125_3477_n648, DP_OP_423J2_125_3477_n647,
         DP_OP_423J2_125_3477_n646, DP_OP_423J2_125_3477_n645,
         DP_OP_423J2_125_3477_n644, DP_OP_423J2_125_3477_n643,
         DP_OP_423J2_125_3477_n642, DP_OP_423J2_125_3477_n641,
         DP_OP_423J2_125_3477_n640, DP_OP_423J2_125_3477_n639,
         DP_OP_423J2_125_3477_n638, DP_OP_423J2_125_3477_n637,
         DP_OP_423J2_125_3477_n636, DP_OP_423J2_125_3477_n635,
         DP_OP_423J2_125_3477_n634, DP_OP_423J2_125_3477_n633,
         DP_OP_423J2_125_3477_n632, DP_OP_423J2_125_3477_n631,
         DP_OP_423J2_125_3477_n630, DP_OP_423J2_125_3477_n629,
         DP_OP_423J2_125_3477_n628, DP_OP_423J2_125_3477_n627,
         DP_OP_423J2_125_3477_n626, DP_OP_423J2_125_3477_n625,
         DP_OP_423J2_125_3477_n624, DP_OP_423J2_125_3477_n623,
         DP_OP_423J2_125_3477_n622, DP_OP_423J2_125_3477_n621,
         DP_OP_423J2_125_3477_n620, DP_OP_423J2_125_3477_n619,
         DP_OP_423J2_125_3477_n618, DP_OP_423J2_125_3477_n617,
         DP_OP_423J2_125_3477_n616, DP_OP_423J2_125_3477_n615,
         DP_OP_423J2_125_3477_n614, DP_OP_423J2_125_3477_n613,
         DP_OP_423J2_125_3477_n612, DP_OP_423J2_125_3477_n611,
         DP_OP_423J2_125_3477_n610, DP_OP_423J2_125_3477_n609,
         DP_OP_423J2_125_3477_n608, DP_OP_423J2_125_3477_n607,
         DP_OP_423J2_125_3477_n606, DP_OP_423J2_125_3477_n605,
         DP_OP_423J2_125_3477_n604, DP_OP_423J2_125_3477_n603,
         DP_OP_423J2_125_3477_n602, DP_OP_423J2_125_3477_n601,
         DP_OP_423J2_125_3477_n600, DP_OP_423J2_125_3477_n599,
         DP_OP_423J2_125_3477_n598, DP_OP_423J2_125_3477_n597,
         DP_OP_423J2_125_3477_n596, DP_OP_423J2_125_3477_n595,
         DP_OP_423J2_125_3477_n594, DP_OP_423J2_125_3477_n593,
         DP_OP_423J2_125_3477_n592, DP_OP_423J2_125_3477_n591,
         DP_OP_423J2_125_3477_n590, DP_OP_423J2_125_3477_n589,
         DP_OP_423J2_125_3477_n588, DP_OP_423J2_125_3477_n587,
         DP_OP_423J2_125_3477_n586, DP_OP_423J2_125_3477_n585,
         DP_OP_423J2_125_3477_n584, DP_OP_423J2_125_3477_n583,
         DP_OP_423J2_125_3477_n582, DP_OP_423J2_125_3477_n581,
         DP_OP_423J2_125_3477_n580, DP_OP_423J2_125_3477_n579,
         DP_OP_423J2_125_3477_n578, DP_OP_423J2_125_3477_n577,
         DP_OP_423J2_125_3477_n576, DP_OP_423J2_125_3477_n575,
         DP_OP_423J2_125_3477_n574, DP_OP_423J2_125_3477_n573,
         DP_OP_423J2_125_3477_n572, DP_OP_423J2_125_3477_n571,
         DP_OP_423J2_125_3477_n570, DP_OP_423J2_125_3477_n569,
         DP_OP_423J2_125_3477_n568, DP_OP_423J2_125_3477_n567,
         DP_OP_423J2_125_3477_n566, DP_OP_423J2_125_3477_n565,
         DP_OP_423J2_125_3477_n564, DP_OP_423J2_125_3477_n563,
         DP_OP_423J2_125_3477_n562, DP_OP_423J2_125_3477_n561,
         DP_OP_423J2_125_3477_n560, DP_OP_423J2_125_3477_n559,
         DP_OP_423J2_125_3477_n558, DP_OP_423J2_125_3477_n557,
         DP_OP_423J2_125_3477_n556, DP_OP_423J2_125_3477_n555,
         DP_OP_423J2_125_3477_n554, DP_OP_423J2_125_3477_n553,
         DP_OP_423J2_125_3477_n552, DP_OP_423J2_125_3477_n551,
         DP_OP_423J2_125_3477_n550, DP_OP_423J2_125_3477_n549,
         DP_OP_423J2_125_3477_n548, DP_OP_423J2_125_3477_n547,
         DP_OP_423J2_125_3477_n546, DP_OP_423J2_125_3477_n545,
         DP_OP_423J2_125_3477_n544, DP_OP_423J2_125_3477_n543,
         DP_OP_423J2_125_3477_n542, DP_OP_423J2_125_3477_n541,
         DP_OP_423J2_125_3477_n540, DP_OP_423J2_125_3477_n539,
         DP_OP_423J2_125_3477_n538, DP_OP_423J2_125_3477_n537,
         DP_OP_423J2_125_3477_n536, DP_OP_423J2_125_3477_n535,
         DP_OP_423J2_125_3477_n534, DP_OP_423J2_125_3477_n533,
         DP_OP_423J2_125_3477_n532, DP_OP_423J2_125_3477_n531,
         DP_OP_423J2_125_3477_n530, DP_OP_423J2_125_3477_n529,
         DP_OP_423J2_125_3477_n528, DP_OP_423J2_125_3477_n527,
         DP_OP_423J2_125_3477_n526, DP_OP_423J2_125_3477_n525,
         DP_OP_423J2_125_3477_n524, DP_OP_423J2_125_3477_n523,
         DP_OP_423J2_125_3477_n522, DP_OP_423J2_125_3477_n521,
         DP_OP_423J2_125_3477_n520, DP_OP_423J2_125_3477_n519,
         DP_OP_423J2_125_3477_n518, DP_OP_423J2_125_3477_n517,
         DP_OP_423J2_125_3477_n516, DP_OP_423J2_125_3477_n515,
         DP_OP_423J2_125_3477_n514, DP_OP_423J2_125_3477_n513,
         DP_OP_423J2_125_3477_n512, DP_OP_423J2_125_3477_n511,
         DP_OP_423J2_125_3477_n510, DP_OP_423J2_125_3477_n509,
         DP_OP_423J2_125_3477_n508, DP_OP_423J2_125_3477_n507,
         DP_OP_423J2_125_3477_n506, DP_OP_423J2_125_3477_n505,
         DP_OP_423J2_125_3477_n504, DP_OP_423J2_125_3477_n503,
         DP_OP_423J2_125_3477_n502, DP_OP_423J2_125_3477_n501,
         DP_OP_423J2_125_3477_n500, DP_OP_423J2_125_3477_n499,
         DP_OP_423J2_125_3477_n498, DP_OP_423J2_125_3477_n497,
         DP_OP_423J2_125_3477_n496, DP_OP_423J2_125_3477_n495,
         DP_OP_423J2_125_3477_n494, DP_OP_423J2_125_3477_n493,
         DP_OP_423J2_125_3477_n492, DP_OP_423J2_125_3477_n491,
         DP_OP_423J2_125_3477_n490, DP_OP_423J2_125_3477_n489,
         DP_OP_423J2_125_3477_n488, DP_OP_423J2_125_3477_n487,
         DP_OP_423J2_125_3477_n486, DP_OP_423J2_125_3477_n485,
         DP_OP_423J2_125_3477_n484, DP_OP_423J2_125_3477_n483,
         DP_OP_423J2_125_3477_n482, DP_OP_423J2_125_3477_n481,
         DP_OP_423J2_125_3477_n480, DP_OP_423J2_125_3477_n479,
         DP_OP_423J2_125_3477_n478, DP_OP_423J2_125_3477_n477,
         DP_OP_423J2_125_3477_n476, DP_OP_423J2_125_3477_n475,
         DP_OP_423J2_125_3477_n474, DP_OP_423J2_125_3477_n473,
         DP_OP_423J2_125_3477_n472, DP_OP_423J2_125_3477_n471,
         DP_OP_423J2_125_3477_n470, DP_OP_423J2_125_3477_n469,
         DP_OP_423J2_125_3477_n468, DP_OP_423J2_125_3477_n467,
         DP_OP_423J2_125_3477_n466, DP_OP_423J2_125_3477_n465,
         DP_OP_423J2_125_3477_n464, DP_OP_423J2_125_3477_n463,
         DP_OP_423J2_125_3477_n462, DP_OP_423J2_125_3477_n461,
         DP_OP_423J2_125_3477_n460, DP_OP_423J2_125_3477_n459,
         DP_OP_423J2_125_3477_n458, DP_OP_423J2_125_3477_n457,
         DP_OP_423J2_125_3477_n456, DP_OP_423J2_125_3477_n455,
         DP_OP_423J2_125_3477_n454, DP_OP_423J2_125_3477_n453,
         DP_OP_423J2_125_3477_n452, DP_OP_423J2_125_3477_n451,
         DP_OP_423J2_125_3477_n450, DP_OP_423J2_125_3477_n449,
         DP_OP_423J2_125_3477_n448, DP_OP_423J2_125_3477_n447,
         DP_OP_423J2_125_3477_n446, DP_OP_423J2_125_3477_n445,
         DP_OP_423J2_125_3477_n444, DP_OP_423J2_125_3477_n443,
         DP_OP_423J2_125_3477_n442, DP_OP_423J2_125_3477_n441,
         DP_OP_423J2_125_3477_n440, DP_OP_423J2_125_3477_n439,
         DP_OP_423J2_125_3477_n438, DP_OP_423J2_125_3477_n437,
         DP_OP_423J2_125_3477_n436, DP_OP_423J2_125_3477_n435,
         DP_OP_423J2_125_3477_n434, DP_OP_423J2_125_3477_n433,
         DP_OP_423J2_125_3477_n432, DP_OP_423J2_125_3477_n431,
         DP_OP_423J2_125_3477_n430, DP_OP_423J2_125_3477_n429,
         DP_OP_423J2_125_3477_n428, DP_OP_423J2_125_3477_n427,
         DP_OP_423J2_125_3477_n426, DP_OP_423J2_125_3477_n425,
         DP_OP_423J2_125_3477_n424, DP_OP_423J2_125_3477_n423,
         DP_OP_423J2_125_3477_n422, DP_OP_423J2_125_3477_n421,
         DP_OP_423J2_125_3477_n420, DP_OP_423J2_125_3477_n419,
         DP_OP_423J2_125_3477_n418, DP_OP_423J2_125_3477_n417,
         DP_OP_423J2_125_3477_n416, DP_OP_423J2_125_3477_n415,
         DP_OP_423J2_125_3477_n414, DP_OP_423J2_125_3477_n413,
         DP_OP_423J2_125_3477_n412, DP_OP_423J2_125_3477_n411,
         DP_OP_423J2_125_3477_n410, DP_OP_423J2_125_3477_n409,
         DP_OP_423J2_125_3477_n408, DP_OP_423J2_125_3477_n407,
         DP_OP_423J2_125_3477_n406, DP_OP_423J2_125_3477_n405,
         DP_OP_423J2_125_3477_n404, DP_OP_423J2_125_3477_n403,
         DP_OP_423J2_125_3477_n402, DP_OP_423J2_125_3477_n401,
         DP_OP_423J2_125_3477_n400, DP_OP_423J2_125_3477_n399,
         DP_OP_423J2_125_3477_n398, DP_OP_423J2_125_3477_n397,
         DP_OP_423J2_125_3477_n396, DP_OP_423J2_125_3477_n395,
         DP_OP_423J2_125_3477_n394, DP_OP_423J2_125_3477_n393,
         DP_OP_423J2_125_3477_n392, DP_OP_423J2_125_3477_n391,
         DP_OP_423J2_125_3477_n390, DP_OP_423J2_125_3477_n389,
         DP_OP_423J2_125_3477_n388, DP_OP_423J2_125_3477_n387,
         DP_OP_423J2_125_3477_n386, DP_OP_423J2_125_3477_n385,
         DP_OP_423J2_125_3477_n384, DP_OP_423J2_125_3477_n383,
         DP_OP_423J2_125_3477_n382, DP_OP_423J2_125_3477_n381,
         DP_OP_423J2_125_3477_n380, DP_OP_423J2_125_3477_n379,
         DP_OP_423J2_125_3477_n378, DP_OP_423J2_125_3477_n377,
         DP_OP_423J2_125_3477_n376, DP_OP_423J2_125_3477_n375,
         DP_OP_423J2_125_3477_n374, DP_OP_423J2_125_3477_n373,
         DP_OP_423J2_125_3477_n372, DP_OP_423J2_125_3477_n371,
         DP_OP_423J2_125_3477_n370, DP_OP_423J2_125_3477_n369,
         DP_OP_423J2_125_3477_n368, DP_OP_423J2_125_3477_n367,
         DP_OP_423J2_125_3477_n366, DP_OP_423J2_125_3477_n365,
         DP_OP_423J2_125_3477_n364, DP_OP_423J2_125_3477_n363,
         DP_OP_423J2_125_3477_n362, DP_OP_423J2_125_3477_n361,
         DP_OP_423J2_125_3477_n360, DP_OP_423J2_125_3477_n359,
         DP_OP_423J2_125_3477_n358, DP_OP_423J2_125_3477_n357,
         DP_OP_423J2_125_3477_n356, DP_OP_423J2_125_3477_n355,
         DP_OP_423J2_125_3477_n354, DP_OP_423J2_125_3477_n353,
         DP_OP_423J2_125_3477_n352, DP_OP_423J2_125_3477_n351,
         DP_OP_423J2_125_3477_n350, DP_OP_423J2_125_3477_n349,
         DP_OP_423J2_125_3477_n348, DP_OP_423J2_125_3477_n347,
         DP_OP_423J2_125_3477_n346, DP_OP_423J2_125_3477_n345,
         DP_OP_423J2_125_3477_n344, DP_OP_423J2_125_3477_n343,
         DP_OP_423J2_125_3477_n342, DP_OP_423J2_125_3477_n341,
         DP_OP_423J2_125_3477_n340, DP_OP_423J2_125_3477_n339,
         DP_OP_423J2_125_3477_n338, DP_OP_423J2_125_3477_n337,
         DP_OP_423J2_125_3477_n336, DP_OP_423J2_125_3477_n335,
         DP_OP_423J2_125_3477_n334, DP_OP_423J2_125_3477_n333,
         DP_OP_423J2_125_3477_n332, DP_OP_423J2_125_3477_n331,
         DP_OP_423J2_125_3477_n330, DP_OP_423J2_125_3477_n329,
         DP_OP_423J2_125_3477_n328, DP_OP_423J2_125_3477_n327,
         DP_OP_423J2_125_3477_n326, DP_OP_423J2_125_3477_n325,
         DP_OP_423J2_125_3477_n324, DP_OP_423J2_125_3477_n323,
         DP_OP_423J2_125_3477_n322, DP_OP_423J2_125_3477_n321,
         DP_OP_423J2_125_3477_n320, DP_OP_423J2_125_3477_n319,
         DP_OP_423J2_125_3477_n318, DP_OP_423J2_125_3477_n317,
         DP_OP_423J2_125_3477_n316, DP_OP_423J2_125_3477_n315,
         DP_OP_423J2_125_3477_n314, DP_OP_423J2_125_3477_n313,
         DP_OP_423J2_125_3477_n312, DP_OP_423J2_125_3477_n311,
         DP_OP_423J2_125_3477_n310, DP_OP_423J2_125_3477_n309,
         DP_OP_423J2_125_3477_n308, DP_OP_423J2_125_3477_n307,
         DP_OP_423J2_125_3477_n306, DP_OP_423J2_125_3477_n305,
         DP_OP_423J2_125_3477_n304, DP_OP_423J2_125_3477_n303,
         DP_OP_423J2_125_3477_n302, DP_OP_423J2_125_3477_n301,
         DP_OP_423J2_125_3477_n300, DP_OP_423J2_125_3477_n299,
         DP_OP_423J2_125_3477_n298, DP_OP_423J2_125_3477_n297,
         DP_OP_423J2_125_3477_n296, DP_OP_423J2_125_3477_n295,
         DP_OP_423J2_125_3477_n294, DP_OP_423J2_125_3477_n293,
         DP_OP_423J2_125_3477_n292, DP_OP_423J2_125_3477_n291,
         DP_OP_423J2_125_3477_n290, DP_OP_423J2_125_3477_n289,
         DP_OP_423J2_125_3477_n288, DP_OP_423J2_125_3477_n287,
         DP_OP_423J2_125_3477_n286, DP_OP_423J2_125_3477_n285,
         DP_OP_423J2_125_3477_n284, DP_OP_423J2_125_3477_n283,
         DP_OP_423J2_125_3477_n282, DP_OP_423J2_125_3477_n281,
         DP_OP_423J2_125_3477_n280, DP_OP_423J2_125_3477_n279,
         DP_OP_423J2_125_3477_n278, DP_OP_423J2_125_3477_n277,
         DP_OP_423J2_125_3477_n276, DP_OP_423J2_125_3477_n275,
         DP_OP_423J2_125_3477_n274, DP_OP_423J2_125_3477_n273,
         DP_OP_423J2_125_3477_n272, DP_OP_423J2_125_3477_n271,
         DP_OP_423J2_125_3477_n270, DP_OP_423J2_125_3477_n269,
         DP_OP_423J2_125_3477_n268, DP_OP_423J2_125_3477_n267,
         DP_OP_423J2_125_3477_n266, DP_OP_423J2_125_3477_n265,
         DP_OP_423J2_125_3477_n264, DP_OP_423J2_125_3477_n263,
         DP_OP_423J2_125_3477_n262, DP_OP_423J2_125_3477_n261,
         DP_OP_423J2_125_3477_n260, DP_OP_423J2_125_3477_n259,
         DP_OP_423J2_125_3477_n258, DP_OP_423J2_125_3477_n257,
         DP_OP_423J2_125_3477_n256, DP_OP_423J2_125_3477_n255,
         DP_OP_423J2_125_3477_n254, DP_OP_423J2_125_3477_n253,
         DP_OP_423J2_125_3477_n252, DP_OP_423J2_125_3477_n251,
         DP_OP_423J2_125_3477_n250, DP_OP_423J2_125_3477_n249,
         DP_OP_423J2_125_3477_n248, DP_OP_423J2_125_3477_n247,
         DP_OP_423J2_125_3477_n246, DP_OP_423J2_125_3477_n245,
         DP_OP_423J2_125_3477_n244, DP_OP_423J2_125_3477_n243,
         DP_OP_423J2_125_3477_n242, DP_OP_423J2_125_3477_n241,
         DP_OP_423J2_125_3477_n240, DP_OP_423J2_125_3477_n239,
         DP_OP_423J2_125_3477_n238, DP_OP_423J2_125_3477_n237,
         DP_OP_423J2_125_3477_n236, DP_OP_423J2_125_3477_n235,
         DP_OP_423J2_125_3477_n234, DP_OP_423J2_125_3477_n233,
         DP_OP_423J2_125_3477_n232, DP_OP_423J2_125_3477_n231,
         DP_OP_423J2_125_3477_n230, DP_OP_423J2_125_3477_n229,
         DP_OP_423J2_125_3477_n228, DP_OP_423J2_125_3477_n227,
         DP_OP_423J2_125_3477_n226, DP_OP_423J2_125_3477_n225,
         DP_OP_423J2_125_3477_n224, DP_OP_423J2_125_3477_n223,
         DP_OP_423J2_125_3477_n222, DP_OP_423J2_125_3477_n221,
         DP_OP_423J2_125_3477_n220, DP_OP_423J2_125_3477_n219,
         DP_OP_423J2_125_3477_n218, DP_OP_423J2_125_3477_n217,
         DP_OP_423J2_125_3477_n216, DP_OP_423J2_125_3477_n215,
         DP_OP_423J2_125_3477_n214, DP_OP_423J2_125_3477_n213,
         DP_OP_423J2_125_3477_n212, DP_OP_423J2_125_3477_n211,
         DP_OP_423J2_125_3477_n210, DP_OP_423J2_125_3477_n209,
         DP_OP_423J2_125_3477_n208, DP_OP_423J2_125_3477_n207,
         DP_OP_423J2_125_3477_n206, DP_OP_423J2_125_3477_n205,
         DP_OP_423J2_125_3477_n204, DP_OP_423J2_125_3477_n203,
         DP_OP_423J2_125_3477_n202, DP_OP_423J2_125_3477_n201,
         DP_OP_423J2_125_3477_n200, DP_OP_423J2_125_3477_n199,
         DP_OP_423J2_125_3477_n198, DP_OP_423J2_125_3477_n197,
         DP_OP_423J2_125_3477_n196, DP_OP_423J2_125_3477_n195,
         DP_OP_423J2_125_3477_n194, DP_OP_423J2_125_3477_n193,
         DP_OP_423J2_125_3477_n192, DP_OP_423J2_125_3477_n191,
         DP_OP_423J2_125_3477_n190, DP_OP_423J2_125_3477_n189,
         DP_OP_423J2_125_3477_n188, DP_OP_423J2_125_3477_n187,
         DP_OP_423J2_125_3477_n186, DP_OP_423J2_125_3477_n185,
         DP_OP_423J2_125_3477_n184, DP_OP_423J2_125_3477_n183,
         DP_OP_423J2_125_3477_n182, DP_OP_423J2_125_3477_n181,
         DP_OP_423J2_125_3477_n180, DP_OP_423J2_125_3477_n179,
         DP_OP_423J2_125_3477_n178, DP_OP_423J2_125_3477_n177,
         DP_OP_423J2_125_3477_n176, DP_OP_423J2_125_3477_n175,
         DP_OP_423J2_125_3477_n174, DP_OP_423J2_125_3477_n173,
         DP_OP_423J2_125_3477_n172, DP_OP_423J2_125_3477_n171,
         DP_OP_423J2_125_3477_n170, DP_OP_423J2_125_3477_n169,
         DP_OP_423J2_125_3477_n168, DP_OP_423J2_125_3477_n167,
         DP_OP_423J2_125_3477_n166, DP_OP_423J2_125_3477_n165,
         DP_OP_423J2_125_3477_n164, DP_OP_423J2_125_3477_n163,
         DP_OP_423J2_125_3477_n162, DP_OP_423J2_125_3477_n161,
         DP_OP_423J2_125_3477_n160, DP_OP_423J2_125_3477_n159,
         DP_OP_423J2_125_3477_n158, DP_OP_423J2_125_3477_n157,
         DP_OP_423J2_125_3477_n156, DP_OP_423J2_125_3477_n155,
         DP_OP_423J2_125_3477_n154, DP_OP_423J2_125_3477_n153,
         DP_OP_423J2_125_3477_n152, DP_OP_423J2_125_3477_n151,
         DP_OP_423J2_125_3477_n150, DP_OP_423J2_125_3477_n149,
         DP_OP_423J2_125_3477_n148, DP_OP_423J2_125_3477_n127,
         DP_OP_423J2_125_3477_n126, DP_OP_423J2_125_3477_n125,
         DP_OP_423J2_125_3477_n124, DP_OP_423J2_125_3477_n121,
         DP_OP_423J2_125_3477_n120, DP_OP_423J2_125_3477_n119,
         DP_OP_423J2_125_3477_n118, DP_OP_423J2_125_3477_n117,
         DP_OP_423J2_125_3477_n116, DP_OP_423J2_125_3477_n113,
         DP_OP_423J2_125_3477_n112, DP_OP_423J2_125_3477_n111,
         DP_OP_423J2_125_3477_n110, DP_OP_423J2_125_3477_n109,
         DP_OP_423J2_125_3477_n108, DP_OP_423J2_125_3477_n105,
         DP_OP_423J2_125_3477_n104, DP_OP_423J2_125_3477_n103,
         DP_OP_423J2_125_3477_n102, DP_OP_423J2_125_3477_n101,
         DP_OP_423J2_125_3477_n100, DP_OP_423J2_125_3477_n99,
         DP_OP_423J2_125_3477_n97, DP_OP_423J2_125_3477_n96,
         DP_OP_423J2_125_3477_n93, DP_OP_423J2_125_3477_n92,
         DP_OP_423J2_125_3477_n91, DP_OP_423J2_125_3477_n90,
         DP_OP_423J2_125_3477_n88, DP_OP_423J2_125_3477_n86,
         DP_OP_423J2_125_3477_n85, DP_OP_423J2_125_3477_n84,
         DP_OP_423J2_125_3477_n83, DP_OP_423J2_125_3477_n82,
         DP_OP_423J2_125_3477_n81, DP_OP_423J2_125_3477_n80,
         DP_OP_423J2_125_3477_n78, DP_OP_423J2_125_3477_n77,
         DP_OP_423J2_125_3477_n76, DP_OP_423J2_125_3477_n75,
         DP_OP_423J2_125_3477_n74, DP_OP_423J2_125_3477_n73,
         DP_OP_423J2_125_3477_n72, DP_OP_423J2_125_3477_n71,
         DP_OP_423J2_125_3477_n67, DP_OP_423J2_125_3477_n66,
         DP_OP_423J2_125_3477_n65, DP_OP_423J2_125_3477_n64,
         DP_OP_423J2_125_3477_n63, DP_OP_423J2_125_3477_n62,
         DP_OP_423J2_125_3477_n60, DP_OP_423J2_125_3477_n58,
         DP_OP_423J2_125_3477_n57, DP_OP_423J2_125_3477_n55,
         DP_OP_423J2_125_3477_n54, DP_OP_423J2_125_3477_n53,
         DP_OP_423J2_125_3477_n51, DP_OP_423J2_125_3477_n50,
         DP_OP_423J2_125_3477_n49, DP_OP_423J2_125_3477_n48,
         DP_OP_423J2_125_3477_n44, DP_OP_423J2_125_3477_n43,
         DP_OP_423J2_125_3477_n40, DP_OP_423J2_125_3477_n39,
         DP_OP_423J2_125_3477_n37, DP_OP_423J2_125_3477_n36,
         DP_OP_423J2_125_3477_n35, DP_OP_423J2_125_3477_n34,
         DP_OP_423J2_125_3477_n33, DP_OP_423J2_125_3477_n32,
         DP_OP_423J2_125_3477_n31, DP_OP_423J2_125_3477_n30,
         DP_OP_423J2_125_3477_n29, DP_OP_423J2_125_3477_n28,
         DP_OP_423J2_125_3477_n27, DP_OP_423J2_125_3477_n26,
         DP_OP_423J2_125_3477_n25, DP_OP_423J2_125_3477_n24,
         DP_OP_423J2_125_3477_n23, DP_OP_423J2_125_3477_n22,
         DP_OP_423J2_125_3477_n3, DP_OP_423J2_125_3477_n2, n1, n3, n5010, n6,
         n8, n900, n11, n12, n13, n14, n17, n18, n20, n21, n23, n24, n25, n26,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n701, n71,
         n72, n73, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n901, n91, n92, n93, n94, n95, n96, n97, n99, n101,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n211, n212, n213, n214,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n5001, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687;
  wire   [31:0] conv2_sum_a;
  wire   [31:0] conv2_sum_b;
  wire   [31:0] tmp_big1;
  wire   [31:0] conv2_sum_c;
  wire   [31:0] conv2_sum_d;
  wire   [31:0] tmp_big2;
  wire   [93:0] conv_weight_box;
  wire   [31:0] n_conv2_sum_a;
  wire   [31:0] n_conv2_sum_b;
  wire   [31:0] n_conv2_sum_c;
  wire   [31:0] n_conv2_sum_d;

  DFFSSRX1_HVT conv2_sum_c_reg_31_ ( .D(1'b0), .SETB(n331), .RSTB(
        n_conv2_sum_c[31]), .CLK(clk), .Q(conv2_sum_c[31]), .QN(n314) );
  DFFSSRX1_HVT conv2_sum_c_reg_30_ ( .D(1'b0), .SETB(n347), .RSTB(
        n_conv2_sum_c[30]), .CLK(clk), .Q(conv2_sum_c[30]), .QN(n414) );
  DFFSSRX1_HVT conv2_sum_c_reg_29_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_c[29]), .CLK(clk), .Q(conv2_sum_c[29]), .QN(n424) );
  DFFSSRX1_HVT conv2_sum_c_reg_28_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_c[28]), .CLK(clk), .Q(conv2_sum_c[28]), .QN(n407) );
  DFFSSRX1_HVT conv2_sum_c_reg_27_ ( .D(1'b0), .SETB(n330), .RSTB(
        n_conv2_sum_c[27]), .CLK(clk), .Q(conv2_sum_c[27]), .QN(n378) );
  DFFSSRX1_HVT conv2_sum_c_reg_26_ ( .D(1'b0), .SETB(n347), .RSTB(
        n_conv2_sum_c[26]), .CLK(clk), .Q(conv2_sum_c[26]), .QN(n396) );
  DFFSSRX1_HVT conv2_sum_c_reg_25_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_c[25]), .CLK(clk), .Q(conv2_sum_c[25]), .QN(n425) );
  DFFSSRX1_HVT conv2_sum_c_reg_24_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_c[24]), .CLK(clk), .Q(conv2_sum_c[24]), .QN(n408) );
  DFFSSRX1_HVT conv2_sum_c_reg_23_ ( .D(1'b0), .SETB(n331), .RSTB(
        n_conv2_sum_c[23]), .CLK(clk), .Q(conv2_sum_c[23]), .QN(n383) );
  DFFSSRX1_HVT conv2_sum_c_reg_22_ ( .D(1'b0), .SETB(n347), .RSTB(
        n_conv2_sum_c[22]), .CLK(clk), .Q(conv2_sum_c[22]), .QN(n415) );
  DFFSSRX1_HVT conv2_sum_c_reg_21_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_c[21]), .CLK(clk), .Q(conv2_sum_c[21]), .QN(n426) );
  DFFSSRX1_HVT conv2_sum_c_reg_20_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_c[20]), .CLK(clk), .Q(conv2_sum_c[20]), .QN(n419) );
  DFFSSRX1_HVT conv2_sum_c_reg_19_ ( .D(1'b0), .SETB(n330), .RSTB(
        n_conv2_sum_c[19]), .CLK(clk), .Q(conv2_sum_c[19]), .QN(n379) );
  DFFSSRX1_HVT conv2_sum_c_reg_18_ ( .D(1'b0), .SETB(n347), .RSTB(
        n_conv2_sum_c[18]), .CLK(clk), .Q(conv2_sum_c[18]), .QN(n416) );
  DFFSSRX1_HVT conv2_sum_c_reg_17_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_c[17]), .CLK(clk), .Q(conv2_sum_c[17]), .QN(n427) );
  DFFSSRX1_HVT conv2_sum_c_reg_16_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_c[16]), .CLK(clk), .Q(conv2_sum_c[16]), .QN(n299) );
  DFFSSRX1_HVT conv2_sum_c_reg_15_ ( .D(1'b0), .SETB(n331), .RSTB(
        n_conv2_sum_c[15]), .CLK(clk), .Q(conv2_sum_c[15]), .QN(n374) );
  DFFSSRX1_HVT conv2_sum_c_reg_14_ ( .D(1'b0), .SETB(n347), .RSTB(
        n_conv2_sum_c[14]), .CLK(clk), .Q(conv2_sum_c[14]), .QN(n417) );
  DFFSSRX1_HVT conv2_sum_c_reg_13_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_c[13]), .CLK(clk), .Q(conv2_sum_c[13]), .QN(n401) );
  DFFSSRX1_HVT conv2_sum_c_reg_12_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_c[12]), .CLK(clk), .Q(conv2_sum_c[12]), .QN(n404) );
  DFFSSRX1_HVT conv2_sum_c_reg_11_ ( .D(1'b0), .SETB(n330), .RSTB(
        n_conv2_sum_c[11]), .CLK(clk), .Q(conv2_sum_c[11]), .QN(n370) );
  DFFSSRX1_HVT conv2_sum_c_reg_10_ ( .D(1'b0), .SETB(n347), .RSTB(
        n_conv2_sum_c[10]), .CLK(clk), .Q(conv2_sum_c[10]), .QN(n393) );
  DFFSSRX1_HVT conv2_sum_c_reg_9_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_c[9]), .CLK(clk), .Q(conv2_sum_c[9]), .QN(n402) );
  DFFSSRX1_HVT conv2_sum_c_reg_8_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_c[8]), .CLK(clk), .Q(conv2_sum_c[8]), .QN(n276) );
  DFFSSRX1_HVT conv2_sum_c_reg_7_ ( .D(1'b0), .SETB(n331), .RSTB(
        n_conv2_sum_c[7]), .CLK(clk), .Q(conv2_sum_c[7]), .QN(n375) );
  DFFSSRX1_HVT conv2_sum_c_reg_6_ ( .D(1'b0), .SETB(n347), .RSTB(
        n_conv2_sum_c[6]), .CLK(clk), .Q(conv2_sum_c[6]), .QN(n395) );
  DFFSSRX1_HVT conv2_sum_c_reg_5_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_c[5]), .CLK(clk), .Q(conv2_sum_c[5]), .QN(n367) );
  DFFSSRX1_HVT conv2_sum_c_reg_4_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_c[4]), .CLK(clk), .Q(conv2_sum_c[4]), .QN(n389) );
  DFFSSRX1_HVT conv2_sum_c_reg_3_ ( .D(1'b0), .SETB(n330), .RSTB(
        n_conv2_sum_c[3]), .CLK(clk), .Q(conv2_sum_c[3]), .QN(n371) );
  DFFSSRX1_HVT conv2_sum_c_reg_2_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_c[2]), .CLK(clk), .Q(conv2_sum_c[2]), .QN(n394) );
  DFFSSRX1_HVT conv2_sum_c_reg_1_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_c[1]), .CLK(clk), .Q(conv2_sum_c[1]), .QN(n286) );
  DFFSSRX1_HVT conv2_sum_c_reg_0_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_c[0]), .CLK(clk), .Q(conv2_sum_c[0]), .QN(n278) );
  DFFSSRX1_HVT conv2_sum_d_reg_31_ ( .D(1'b0), .SETB(n331), .RSTB(
        n_conv2_sum_d[31]), .CLK(clk), .Q(conv2_sum_d[31]), .QN(n381) );
  DFFSSRX1_HVT conv2_sum_d_reg_30_ ( .D(1'b0), .SETB(n347), .RSTB(
        n_conv2_sum_d[30]), .CLK(clk), .Q(conv2_sum_d[30]), .QN(n321) );
  DFFSSRX1_HVT conv2_sum_d_reg_29_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_d[29]), .CLK(clk), .Q(conv2_sum_d[29]), .QN(n327) );
  DFFSSRX1_HVT conv2_sum_d_reg_28_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_d[28]), .CLK(clk), .Q(conv2_sum_d[28]), .QN(n325) );
  DFFSSRX1_HVT conv2_sum_d_reg_27_ ( .D(1'b0), .SETB(n330), .RSTB(
        n_conv2_sum_d[27]), .CLK(clk), .Q(conv2_sum_d[27]), .QN(n317) );
  DFFSSRX1_HVT conv2_sum_d_reg_26_ ( .D(1'b0), .SETB(n347), .RSTB(
        n_conv2_sum_d[26]), .CLK(clk), .Q(conv2_sum_d[26]), .QN(n318) );
  DFFSSRX1_HVT conv2_sum_d_reg_25_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_d[25]), .CLK(clk), .Q(conv2_sum_d[25]), .QN(n329) );
  DFFSSRX1_HVT conv2_sum_d_reg_24_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_d[24]), .CLK(clk), .Q(conv2_sum_d[24]), .QN(n322) );
  DFFSSRX1_HVT conv2_sum_d_reg_23_ ( .D(1'b0), .SETB(n331), .RSTB(
        n_conv2_sum_d[23]), .CLK(clk), .Q(conv2_sum_d[23]), .QN(n303) );
  DFFSSRX1_HVT conv2_sum_d_reg_22_ ( .D(1'b0), .SETB(n347), .RSTB(
        n_conv2_sum_d[22]), .CLK(clk), .Q(conv2_sum_d[22]), .QN(n307) );
  DFFSSRX1_HVT conv2_sum_d_reg_21_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_d[21]), .CLK(clk), .Q(conv2_sum_d[21]), .QN(n310) );
  DFFSSRX1_HVT conv2_sum_d_reg_20_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_d[20]), .CLK(clk), .Q(conv2_sum_d[20]), .QN(n309) );
  DFFSSRX1_HVT conv2_sum_d_reg_19_ ( .D(1'b0), .SETB(n330), .RSTB(
        n_conv2_sum_d[19]), .CLK(clk), .Q(conv2_sum_d[19]), .QN(n305) );
  DFFSSRX1_HVT conv2_sum_d_reg_18_ ( .D(1'b0), .SETB(n347), .RSTB(
        n_conv2_sum_d[18]), .CLK(clk), .Q(conv2_sum_d[18]), .QN(n312) );
  DFFSSRX1_HVT conv2_sum_d_reg_17_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_d[17]), .CLK(clk), .Q(conv2_sum_d[17]), .QN(n301) );
  DFFSSRX1_HVT conv2_sum_d_reg_16_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_d[16]), .CLK(clk), .Q(conv2_sum_d[16]), .QN(n398) );
  DFFSSRX1_HVT conv2_sum_d_reg_15_ ( .D(1'b0), .SETB(n331), .RSTB(
        n_conv2_sum_d[15]), .CLK(clk), .Q(conv2_sum_d[15]), .QN(n294) );
  DFFSSRX1_HVT conv2_sum_d_reg_14_ ( .D(1'b0), .SETB(n347), .RSTB(
        n_conv2_sum_d[14]), .CLK(clk), .Q(conv2_sum_d[14]), .QN(n297) );
  DFFSSRX1_HVT conv2_sum_d_reg_13_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_d[13]), .CLK(clk), .Q(conv2_sum_d[13]), .QN(n289) );
  DFFSSRX1_HVT conv2_sum_d_reg_12_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_d[12]), .CLK(clk), .Q(conv2_sum_d[12]), .QN(n287) );
  DFFSSRX1_HVT conv2_sum_d_reg_11_ ( .D(1'b0), .SETB(n330), .RSTB(
        n_conv2_sum_d[11]), .CLK(clk), .Q(conv2_sum_d[11]), .QN(n282) );
  DFFSSRX1_HVT conv2_sum_d_reg_10_ ( .D(1'b0), .SETB(n347), .RSTB(
        n_conv2_sum_d[10]), .CLK(clk), .Q(conv2_sum_d[10]), .QN(n284) );
  DFFSSRX1_HVT conv2_sum_d_reg_9_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_d[9]), .CLK(clk), .Q(conv2_sum_d[9]), .QN(n291) );
  DFFSSRX1_HVT conv2_sum_d_reg_8_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_d[8]), .CLK(clk), .Q(conv2_sum_d[8]), .QN(n387) );
  DFFSSRX1_HVT conv2_sum_d_reg_7_ ( .D(1'b0), .SETB(n331), .RSTB(
        n_conv2_sum_d[7]), .CLK(clk), .Q(conv2_sum_d[7]), .QN(n265) );
  DFFSSRX1_HVT conv2_sum_d_reg_6_ ( .D(1'b0), .SETB(n347), .RSTB(
        n_conv2_sum_d[6]), .CLK(clk), .Q(conv2_sum_d[6]), .QN(n275) );
  DFFSSRX1_HVT conv2_sum_d_reg_5_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_d[5]), .CLK(clk), .Q(conv2_sum_d[5]), .QN(n268) );
  DFFSSRX1_HVT conv2_sum_d_reg_4_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_d[4]), .CLK(clk), .Q(conv2_sum_d[4]), .QN(n272) );
  DFFSSRX1_HVT conv2_sum_d_reg_3_ ( .D(1'b0), .SETB(n330), .RSTB(
        n_conv2_sum_d[3]), .CLK(clk), .Q(conv2_sum_d[3]), .QN(n267) );
  DFFSSRX1_HVT conv2_sum_d_reg_2_ ( .D(1'b0), .SETB(n347), .RSTB(
        n_conv2_sum_d[2]), .CLK(clk), .Q(conv2_sum_d[2]), .QN(n270) );
  DFFSSRX1_HVT conv2_sum_d_reg_1_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_d[1]), .CLK(clk), .Q(conv2_sum_d[1]), .QN(n385) );
  DFFSSRX1_HVT conv2_sum_d_reg_0_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_d[0]), .CLK(clk), .Q(conv2_sum_d[0]), .QN(n280) );
  DFFSSRX1_HVT conv2_sum_a_reg_31_ ( .D(1'b0), .SETB(n331), .RSTB(
        n_conv2_sum_a[31]), .CLK(clk), .Q(conv2_sum_a[31]), .QN(n315) );
  DFFSSRX1_HVT conv2_sum_a_reg_30_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_a[30]), .CLK(clk), .Q(conv2_sum_a[30]), .QN(n409) );
  DFFSSRX1_HVT conv2_sum_a_reg_29_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_a[29]), .CLK(clk), .Q(conv2_sum_a[29]), .QN(n420) );
  DFFSSRX1_HVT conv2_sum_a_reg_28_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_a[28]), .CLK(clk), .Q(conv2_sum_a[28]), .QN(n405) );
  DFFSSRX1_HVT conv2_sum_a_reg_27_ ( .D(1'b0), .SETB(n330), .RSTB(
        n_conv2_sum_a[27]), .CLK(clk), .Q(conv2_sum_a[27]), .QN(n376) );
  DFFSSRX1_HVT conv2_sum_a_reg_26_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_a[26]), .CLK(clk), .Q(conv2_sum_a[26]), .QN(n410) );
  DFFSSRX1_HVT conv2_sum_a_reg_25_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_a[25]), .CLK(clk), .Q(conv2_sum_a[25]), .QN(n421) );
  DFFSSRX1_HVT conv2_sum_a_reg_24_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_a[24]), .CLK(clk), .Q(conv2_sum_a[24]), .QN(n418) );
  DFFSSRX1_HVT conv2_sum_a_reg_23_ ( .D(1'b0), .SETB(n331), .RSTB(
        n_conv2_sum_a[23]), .CLK(clk), .Q(conv2_sum_a[23]), .QN(n382) );
  DFFSSRX1_HVT conv2_sum_a_reg_22_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_a[22]), .CLK(clk), .Q(conv2_sum_a[22]), .QN(n411) );
  DFFSSRX1_HVT conv2_sum_a_reg_21_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_a[21]), .CLK(clk), .Q(conv2_sum_a[21]), .QN(n422) );
  DFFSSRX1_HVT conv2_sum_a_reg_20_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_a[20]), .CLK(clk), .Q(conv2_sum_a[20]), .QN(n406) );
  DFFSSRX1_HVT conv2_sum_a_reg_19_ ( .D(1'b0), .SETB(n330), .RSTB(
        n_conv2_sum_a[19]), .CLK(clk), .Q(conv2_sum_a[19]), .QN(n377) );
  DFFSSRX1_HVT conv2_sum_a_reg_18_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_a[18]), .CLK(clk), .Q(conv2_sum_a[18]), .QN(n412) );
  DFFSSRX1_HVT conv2_sum_a_reg_17_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_a[17]), .CLK(clk), .Q(conv2_sum_a[17]), .QN(n423) );
  DFFSSRX1_HVT conv2_sum_a_reg_16_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_a[16]), .CLK(clk), .Q(conv2_sum_a[16]), .QN(n298) );
  DFFSSRX1_HVT conv2_sum_a_reg_15_ ( .D(1'b0), .SETB(n331), .RSTB(
        n_conv2_sum_a[15]), .CLK(clk), .Q(conv2_sum_a[15]), .QN(n372) );
  DFFSSRX1_HVT conv2_sum_a_reg_14_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_a[14]), .CLK(clk), .Q(conv2_sum_a[14]), .QN(n413) );
  DFFSSRX1_HVT conv2_sum_a_reg_13_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_a[13]), .CLK(clk), .Q(conv2_sum_a[13]), .QN(n399) );
  DFFSSRX1_HVT conv2_sum_a_reg_12_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_a[12]), .CLK(clk), .Q(conv2_sum_a[12]), .QN(n403) );
  DFFSSRX1_HVT conv2_sum_a_reg_11_ ( .D(1'b0), .SETB(n330), .RSTB(
        n_conv2_sum_a[11]), .CLK(clk), .Q(conv2_sum_a[11]), .QN(n368) );
  DFFSSRX1_HVT conv2_sum_a_reg_10_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_a[10]), .CLK(clk), .Q(conv2_sum_a[10]), .QN(n390) );
  DFFSSRX1_HVT conv2_sum_a_reg_9_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_a[9]), .CLK(clk), .Q(conv2_sum_a[9]), .QN(n400) );
  DFFSSRX1_HVT conv2_sum_a_reg_8_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_a[8]), .CLK(clk), .Q(conv2_sum_a[8]), .QN(n277) );
  DFFSSRX1_HVT conv2_sum_a_reg_7_ ( .D(1'b0), .SETB(n331), .RSTB(
        n_conv2_sum_a[7]), .CLK(clk), .Q(conv2_sum_a[7]), .QN(n373) );
  DFFSSRX1_HVT conv2_sum_a_reg_6_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_a[6]), .CLK(clk), .Q(conv2_sum_a[6]), .QN(n392) );
  DFFSSRX1_HVT conv2_sum_a_reg_5_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_a[5]), .CLK(clk), .Q(conv2_sum_a[5]), .QN(n366) );
  DFFSSRX1_HVT conv2_sum_a_reg_4_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_a[4]), .CLK(clk), .Q(conv2_sum_a[4]), .QN(n388) );
  DFFSSRX1_HVT conv2_sum_a_reg_3_ ( .D(1'b0), .SETB(n330), .RSTB(
        n_conv2_sum_a[3]), .CLK(clk), .Q(conv2_sum_a[3]), .QN(n369) );
  DFFSSRX1_HVT conv2_sum_a_reg_2_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_a[2]), .CLK(clk), .Q(conv2_sum_a[2]), .QN(n391) );
  DFFSSRX1_HVT conv2_sum_a_reg_1_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_a[1]), .CLK(clk), .Q(conv2_sum_a[1]), .QN(n285) );
  DFFSSRX1_HVT conv2_sum_a_reg_0_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_a[0]), .CLK(clk), .Q(conv2_sum_a[0]), .QN(n279) );
  DFFSSRX1_HVT conv2_sum_b_reg_31_ ( .D(1'b0), .SETB(n331), .RSTB(
        n_conv2_sum_b[31]), .CLK(clk), .Q(conv2_sum_b[31]), .QN(n380) );
  DFFSSRX1_HVT conv2_sum_b_reg_30_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_b[30]), .CLK(clk), .Q(conv2_sum_b[30]), .QN(n320) );
  DFFSSRX1_HVT conv2_sum_b_reg_29_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_b[29]), .CLK(clk), .Q(conv2_sum_b[29]), .QN(n326) );
  DFFSSRX1_HVT conv2_sum_b_reg_28_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_b[28]), .CLK(clk), .Q(conv2_sum_b[28]), .QN(n323) );
  DFFSSRX1_HVT conv2_sum_b_reg_27_ ( .D(1'b0), .SETB(n330), .RSTB(
        n_conv2_sum_b[27]), .CLK(clk), .Q(conv2_sum_b[27]), .QN(n316) );
  DFFSSRX1_HVT conv2_sum_b_reg_26_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_b[26]), .CLK(clk), .Q(conv2_sum_b[26]), .QN(n319) );
  DFFSSRX1_HVT conv2_sum_b_reg_25_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_b[25]), .CLK(clk), .Q(conv2_sum_b[25]), .QN(n328) );
  DFFSSRX1_HVT conv2_sum_b_reg_24_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_b[24]), .CLK(clk), .Q(conv2_sum_b[24]), .QN(n324) );
  DFFSSRX1_HVT conv2_sum_b_reg_23_ ( .D(1'b0), .SETB(n331), .RSTB(
        n_conv2_sum_b[23]), .CLK(clk), .Q(conv2_sum_b[23]), .QN(n302) );
  DFFSSRX1_HVT conv2_sum_b_reg_22_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_b[22]), .CLK(clk), .Q(conv2_sum_b[22]), .QN(n306) );
  DFFSSRX1_HVT conv2_sum_b_reg_21_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_b[21]), .CLK(clk), .Q(conv2_sum_b[21]), .QN(n311) );
  DFFSSRX1_HVT conv2_sum_b_reg_20_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_b[20]), .CLK(clk), .Q(conv2_sum_b[20]), .QN(n308) );
  DFFSSRX1_HVT conv2_sum_b_reg_19_ ( .D(1'b0), .SETB(n330), .RSTB(
        n_conv2_sum_b[19]), .CLK(clk), .Q(conv2_sum_b[19]), .QN(n304) );
  DFFSSRX1_HVT conv2_sum_b_reg_18_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_b[18]), .CLK(clk), .Q(conv2_sum_b[18]), .QN(n313) );
  DFFSSRX1_HVT conv2_sum_b_reg_17_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_b[17]), .CLK(clk), .Q(conv2_sum_b[17]), .QN(n300) );
  DFFSSRX1_HVT conv2_sum_b_reg_16_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_b[16]), .CLK(clk), .Q(conv2_sum_b[16]), .QN(n397) );
  DFFSSRX1_HVT conv2_sum_b_reg_15_ ( .D(1'b0), .SETB(n331), .RSTB(
        n_conv2_sum_b[15]), .CLK(clk), .Q(conv2_sum_b[15]), .QN(n295) );
  DFFSSRX1_HVT conv2_sum_b_reg_14_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_b[14]), .CLK(clk), .Q(conv2_sum_b[14]), .QN(n296) );
  DFFSSRX1_HVT conv2_sum_b_reg_13_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_b[13]), .CLK(clk), .Q(conv2_sum_b[13]), .QN(n290) );
  DFFSSRX1_HVT conv2_sum_b_reg_12_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_b[12]), .CLK(clk), .Q(conv2_sum_b[12]), .QN(n288) );
  DFFSSRX1_HVT conv2_sum_b_reg_11_ ( .D(1'b0), .SETB(n330), .RSTB(
        n_conv2_sum_b[11]), .CLK(clk), .Q(conv2_sum_b[11]), .QN(n281) );
  DFFSSRX1_HVT conv2_sum_b_reg_10_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_b[10]), .CLK(clk), .Q(conv2_sum_b[10]), .QN(n283) );
  DFFSSRX1_HVT conv2_sum_b_reg_9_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_b[9]), .CLK(clk), .Q(conv2_sum_b[9]), .QN(n292) );
  DFFSSRX1_HVT conv2_sum_b_reg_8_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_b[8]), .CLK(clk), .Q(conv2_sum_b[8]), .QN(n386) );
  DFFSSRX1_HVT conv2_sum_b_reg_7_ ( .D(1'b0), .SETB(n331), .RSTB(
        n_conv2_sum_b[7]), .CLK(clk), .Q(conv2_sum_b[7]), .QN(n264) );
  DFFSSRX1_HVT conv2_sum_b_reg_6_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_b[6]), .CLK(clk), .Q(conv2_sum_b[6]), .QN(n274) );
  DFFSSRX1_HVT conv2_sum_b_reg_5_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_b[5]), .CLK(clk), .Q(conv2_sum_b[5]), .QN(n269) );
  DFFSSRX1_HVT conv2_sum_b_reg_4_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_b[4]), .CLK(clk), .Q(conv2_sum_b[4]), .QN(n273) );
  DFFSSRX1_HVT conv2_sum_b_reg_3_ ( .D(1'b0), .SETB(n330), .RSTB(
        n_conv2_sum_b[3]), .CLK(clk), .Q(conv2_sum_b[3]), .QN(n266) );
  DFFSSRX1_HVT conv2_sum_b_reg_2_ ( .D(1'b0), .SETB(n344), .RSTB(
        n_conv2_sum_b[2]), .CLK(clk), .Q(conv2_sum_b[2]), .QN(n271) );
  DFFSSRX1_HVT conv2_sum_b_reg_1_ ( .D(1'b0), .SETB(n346), .RSTB(
        n_conv2_sum_b[1]), .CLK(clk), .Q(conv2_sum_b[1]), .QN(n384) );
  DFFSSRX1_HVT conv2_sum_b_reg_0_ ( .D(1'b0), .SETB(n345), .RSTB(
        n_conv2_sum_b[0]), .CLK(clk), .Q(conv2_sum_b[0]), .QN(n293) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2130 ( .A1(DP_OP_425J2_127_3477_n2908), 
        .A2(DP_OP_425J2_127_3477_n2918), .Y(DP_OP_425J2_127_3477_n2900) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2129 ( .A1(DP_OP_425J2_127_3477_n2907), .A2(
        DP_OP_425J2_127_3477_n2918), .Y(DP_OP_425J2_127_3477_n2899) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2122 ( .A1(DP_OP_425J2_127_3477_n2908), 
        .A2(DP_OP_425J2_127_3477_n2917), .Y(DP_OP_425J2_127_3477_n2892) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2121 ( .A1(DP_OP_425J2_127_3477_n2907), .A2(
        DP_OP_425J2_127_3477_n2917), .Y(DP_OP_425J2_127_3477_n2891) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2114 ( .A1(DP_OP_425J2_127_3477_n2908), 
        .A2(DP_OP_425J2_127_3477_n2916), .Y(DP_OP_425J2_127_3477_n2884) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2113 ( .A1(DP_OP_425J2_127_3477_n2907), .A2(
        DP_OP_425J2_127_3477_n2916), .Y(DP_OP_425J2_127_3477_n2883) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2112 ( .A1(DP_OP_425J2_127_3477_n2914), .A2(
        DP_OP_425J2_127_3477_n2915), .Y(DP_OP_425J2_127_3477_n2882) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2111 ( .A1(DP_OP_425J2_127_3477_n2913), .A2(
        DP_OP_425J2_127_3477_n2915), .Y(DP_OP_425J2_127_3477_n2881) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2110 ( .A1(DP_OP_425J2_127_3477_n2912), .A2(
        DP_OP_425J2_127_3477_n2915), .Y(DP_OP_425J2_127_3477_n2880) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2109 ( .A1(DP_OP_425J2_127_3477_n2911), .A2(
        DP_OP_425J2_127_3477_n2915), .Y(DP_OP_425J2_127_3477_n2879) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2108 ( .A1(DP_OP_425J2_127_3477_n2910), .A2(
        DP_OP_425J2_127_3477_n2915), .Y(DP_OP_425J2_127_3477_n2878) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2107 ( .A1(DP_OP_425J2_127_3477_n2909), .A2(
        DP_OP_425J2_127_3477_n2915), .Y(DP_OP_425J2_127_3477_n2877) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2106 ( .A1(DP_OP_425J2_127_3477_n2908), .A2(
        DP_OP_425J2_127_3477_n2915), .Y(DP_OP_425J2_127_3477_n2876) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2105 ( .A1(DP_OP_425J2_127_3477_n2907), 
        .A2(DP_OP_425J2_127_3477_n2915), .Y(DP_OP_425J2_127_3477_n2875) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2086 ( .A1(DP_OP_425J2_127_3477_n2864), 
        .A2(DP_OP_425J2_127_3477_n2874), .Y(DP_OP_425J2_127_3477_n2856) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2085 ( .A1(DP_OP_424J2_126_3477_n1854), .A2(
        DP_OP_425J2_127_3477_n2874), .Y(DP_OP_425J2_127_3477_n2855) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2078 ( .A1(DP_OP_425J2_127_3477_n2864), 
        .A2(DP_OP_423J2_125_3477_n2868), .Y(DP_OP_425J2_127_3477_n2848) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2077 ( .A1(DP_OP_424J2_126_3477_n1854), .A2(
        DP_OP_422J2_124_3477_n2873), .Y(DP_OP_425J2_127_3477_n2847) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2070 ( .A1(DP_OP_425J2_127_3477_n2864), 
        .A2(DP_OP_425J2_127_3477_n2872), .Y(DP_OP_425J2_127_3477_n2840) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2069 ( .A1(DP_OP_424J2_126_3477_n1854), .A2(
        DP_OP_425J2_127_3477_n2872), .Y(DP_OP_425J2_127_3477_n2839) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2068 ( .A1(DP_OP_425J2_127_3477_n2870), .A2(
        DP_OP_425J2_127_3477_n2871), .Y(DP_OP_425J2_127_3477_n2838) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2067 ( .A1(DP_OP_425J2_127_3477_n2869), .A2(
        DP_OP_425J2_127_3477_n2871), .Y(DP_OP_425J2_127_3477_n2837) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2066 ( .A1(DP_OP_425J2_127_3477_n2868), .A2(
        DP_OP_425J2_127_3477_n2871), .Y(DP_OP_425J2_127_3477_n2836) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2065 ( .A1(DP_OP_424J2_126_3477_n1858), .A2(
        DP_OP_425J2_127_3477_n2871), .Y(DP_OP_425J2_127_3477_n2835) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2064 ( .A1(DP_OP_424J2_126_3477_n1857), .A2(
        DP_OP_425J2_127_3477_n2871), .Y(DP_OP_425J2_127_3477_n2834) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2063 ( .A1(DP_OP_425J2_127_3477_n2865), .A2(
        DP_OP_425J2_127_3477_n2871), .Y(DP_OP_425J2_127_3477_n2833) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2062 ( .A1(DP_OP_425J2_127_3477_n2864), .A2(
        DP_OP_425J2_127_3477_n2871), .Y(DP_OP_425J2_127_3477_n2832) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2061 ( .A1(DP_OP_424J2_126_3477_n1854), 
        .A2(DP_OP_425J2_127_3477_n2871), .Y(DP_OP_425J2_127_3477_n2831) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2042 ( .A1(DP_OP_425J2_127_3477_n2820), 
        .A2(DP_OP_425J2_127_3477_n2830), .Y(DP_OP_425J2_127_3477_n2812) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2041 ( .A1(DP_OP_424J2_126_3477_n1898), .A2(
        DP_OP_425J2_127_3477_n2830), .Y(DP_OP_425J2_127_3477_n2811) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2034 ( .A1(DP_OP_425J2_127_3477_n2820), 
        .A2(DP_OP_425J2_127_3477_n2829), .Y(DP_OP_425J2_127_3477_n2804) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2033 ( .A1(DP_OP_424J2_126_3477_n1898), .A2(
        DP_OP_425J2_127_3477_n2829), .Y(DP_OP_425J2_127_3477_n2803) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2025 ( .A1(DP_OP_424J2_126_3477_n1898), .A2(
        DP_OP_425J2_127_3477_n2828), .Y(DP_OP_425J2_127_3477_n2795) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2024 ( .A1(DP_OP_425J2_127_3477_n2826), .A2(
        DP_OP_425J2_127_3477_n2827), .Y(DP_OP_425J2_127_3477_n2794) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2023 ( .A1(DP_OP_424J2_126_3477_n1904), .A2(
        DP_OP_425J2_127_3477_n2827), .Y(DP_OP_425J2_127_3477_n2793) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2022 ( .A1(DP_OP_424J2_126_3477_n1903), .A2(
        DP_OP_425J2_127_3477_n2827), .Y(DP_OP_425J2_127_3477_n2792) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2021 ( .A1(DP_OP_425J2_127_3477_n2823), .A2(
        DP_OP_425J2_127_3477_n2827), .Y(DP_OP_425J2_127_3477_n2791) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2020 ( .A1(DP_OP_424J2_126_3477_n1901), .A2(
        DP_OP_425J2_127_3477_n2827), .Y(DP_OP_425J2_127_3477_n2790) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2019 ( .A1(DP_OP_425J2_127_3477_n2821), .A2(
        DP_OP_425J2_127_3477_n2827), .Y(DP_OP_425J2_127_3477_n2789) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2018 ( .A1(DP_OP_425J2_127_3477_n2820), .A2(
        DP_OP_425J2_127_3477_n2827), .Y(DP_OP_425J2_127_3477_n2788) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2017 ( .A1(DP_OP_424J2_126_3477_n1898), 
        .A2(DP_OP_425J2_127_3477_n2827), .Y(DP_OP_425J2_127_3477_n2787) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1998 ( .A1(DP_OP_423J2_125_3477_n1850), 
        .A2(DP_OP_425J2_127_3477_n2786), .Y(DP_OP_425J2_127_3477_n2768) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1997 ( .A1(DP_OP_423J2_125_3477_n1849), .A2(
        DP_OP_425J2_127_3477_n2786), .Y(DP_OP_425J2_127_3477_n2767) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1989 ( .A1(DP_OP_424J2_126_3477_n1942), .A2(
        DP_OP_425J2_127_3477_n2785), .Y(DP_OP_425J2_127_3477_n2759) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1982 ( .A1(DP_OP_423J2_125_3477_n1850), 
        .A2(DP_OP_422J2_124_3477_n2784), .Y(DP_OP_425J2_127_3477_n2752) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1981 ( .A1(DP_OP_423J2_125_3477_n1849), .A2(
        DP_OP_423J2_125_3477_n2779), .Y(DP_OP_425J2_127_3477_n2751) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1980 ( .A1(DP_OP_424J2_126_3477_n1949), .A2(
        DP_OP_425J2_127_3477_n2783), .Y(DP_OP_425J2_127_3477_n2750) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1979 ( .A1(DP_OP_424J2_126_3477_n1948), .A2(
        DP_OP_425J2_127_3477_n2783), .Y(DP_OP_425J2_127_3477_n2749) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1978 ( .A1(DP_OP_425J2_127_3477_n2780), .A2(
        DP_OP_425J2_127_3477_n2783), .Y(DP_OP_425J2_127_3477_n2748) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1977 ( .A1(DP_OP_425J2_127_3477_n2779), .A2(
        DP_OP_425J2_127_3477_n2783), .Y(DP_OP_425J2_127_3477_n2747) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1976 ( .A1(DP_OP_425J2_127_3477_n2778), .A2(
        DP_OP_425J2_127_3477_n2783), .Y(DP_OP_425J2_127_3477_n2746) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1975 ( .A1(DP_OP_425J2_127_3477_n2777), .A2(
        DP_OP_425J2_127_3477_n2783), .Y(DP_OP_425J2_127_3477_n2745) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1974 ( .A1(DP_OP_423J2_125_3477_n1850), .A2(
        DP_OP_425J2_127_3477_n2783), .Y(DP_OP_425J2_127_3477_n2744) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1973 ( .A1(DP_OP_423J2_125_3477_n1849), 
        .A2(DP_OP_425J2_127_3477_n2783), .Y(DP_OP_425J2_127_3477_n2743) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1954 ( .A1(DP_OP_425J2_127_3477_n2732), 
        .A2(DP_OP_423J2_125_3477_n2737), .Y(DP_OP_425J2_127_3477_n2724) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1953 ( .A1(DP_OP_424J2_126_3477_n1986), .A2(
        DP_OP_424J2_126_3477_n2742), .Y(DP_OP_425J2_127_3477_n2723) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1945 ( .A1(DP_OP_423J2_125_3477_n1893), .A2(
        DP_OP_425J2_127_3477_n2741), .Y(DP_OP_425J2_127_3477_n2715) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1937 ( .A1(DP_OP_423J2_125_3477_n1893), .A2(
        DP_OP_425J2_127_3477_n2740), .Y(DP_OP_425J2_127_3477_n2707) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1936 ( .A1(DP_OP_425J2_127_3477_n2738), .A2(
        DP_OP_425J2_127_3477_n2739), .Y(DP_OP_425J2_127_3477_n2706) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1935 ( .A1(DP_OP_423J2_125_3477_n1899), .A2(
        DP_OP_425J2_127_3477_n2739), .Y(DP_OP_425J2_127_3477_n2705) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1934 ( .A1(DP_OP_423J2_125_3477_n1898), .A2(
        DP_OP_425J2_127_3477_n2739), .Y(DP_OP_425J2_127_3477_n2704) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1933 ( .A1(DP_OP_425J2_127_3477_n2735), .A2(
        DP_OP_425J2_127_3477_n2739), .Y(DP_OP_425J2_127_3477_n2703) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1932 ( .A1(DP_OP_425J2_127_3477_n2734), .A2(
        DP_OP_425J2_127_3477_n2739), .Y(DP_OP_425J2_127_3477_n2702) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1931 ( .A1(DP_OP_422J2_124_3477_n2865), .A2(
        DP_OP_425J2_127_3477_n2739), .Y(DP_OP_425J2_127_3477_n2701) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1930 ( .A1(DP_OP_425J2_127_3477_n2732), .A2(
        DP_OP_425J2_127_3477_n2739), .Y(DP_OP_425J2_127_3477_n2700) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1929 ( .A1(DP_OP_424J2_126_3477_n1986), 
        .A2(DP_OP_425J2_127_3477_n2739), .Y(DP_OP_425J2_127_3477_n2699) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1910 ( .A1(DP_OP_425J2_127_3477_n2688), 
        .A2(DP_OP_423J2_125_3477_n2696), .Y(DP_OP_425J2_127_3477_n2680) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1909 ( .A1(DP_OP_423J2_125_3477_n1937), .A2(
        DP_OP_423J2_125_3477_n2696), .Y(DP_OP_425J2_127_3477_n2679) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1901 ( .A1(DP_OP_423J2_125_3477_n1937), .A2(
        DP_OP_423J2_125_3477_n2695), .Y(DP_OP_425J2_127_3477_n2671) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1894 ( .A1(DP_OP_425J2_127_3477_n2688), 
        .A2(DP_OP_425J2_127_3477_n2696), .Y(DP_OP_425J2_127_3477_n2664) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1893 ( .A1(DP_OP_423J2_125_3477_n1937), .A2(
        DP_OP_425J2_127_3477_n2696), .Y(DP_OP_425J2_127_3477_n2663) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1892 ( .A1(DP_OP_425J2_127_3477_n2694), .A2(
        DP_OP_424J2_126_3477_n2695), .Y(DP_OP_425J2_127_3477_n2662) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1891 ( .A1(DP_OP_423J2_125_3477_n1943), .A2(
        DP_OP_423J2_125_3477_n2693), .Y(DP_OP_425J2_127_3477_n2661) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1890 ( .A1(DP_OP_425J2_127_3477_n2692), .A2(
        DP_OP_423J2_125_3477_n2693), .Y(DP_OP_425J2_127_3477_n2660) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1889 ( .A1(DP_OP_425J2_127_3477_n2691), .A2(
        DP_OP_424J2_126_3477_n2695), .Y(DP_OP_425J2_127_3477_n2659) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1888 ( .A1(DP_OP_425J2_127_3477_n2690), .A2(
        DP_OP_423J2_125_3477_n2693), .Y(DP_OP_425J2_127_3477_n2658) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1887 ( .A1(DP_OP_423J2_125_3477_n1939), .A2(
        DP_OP_424J2_126_3477_n2695), .Y(DP_OP_425J2_127_3477_n2657) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1886 ( .A1(DP_OP_425J2_127_3477_n2688), .A2(
        DP_OP_424J2_126_3477_n2695), .Y(DP_OP_425J2_127_3477_n2656) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1885 ( .A1(DP_OP_423J2_125_3477_n1937), 
        .A2(DP_OP_423J2_125_3477_n2693), .Y(DP_OP_425J2_127_3477_n2655) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1866 ( .A1(DP_OP_425J2_127_3477_n2644), 
        .A2(DP_OP_425J2_127_3477_n2654), .Y(DP_OP_425J2_127_3477_n2636) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1865 ( .A1(DP_OP_425J2_127_3477_n2643), .A2(
        DP_OP_425J2_127_3477_n2654), .Y(DP_OP_425J2_127_3477_n2635) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1858 ( .A1(DP_OP_425J2_127_3477_n2644), 
        .A2(DP_OP_424J2_126_3477_n2653), .Y(DP_OP_425J2_127_3477_n2628) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1857 ( .A1(DP_OP_425J2_127_3477_n2643), .A2(
        DP_OP_423J2_125_3477_n2651), .Y(DP_OP_425J2_127_3477_n2627) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1850 ( .A1(DP_OP_425J2_127_3477_n2644), 
        .A2(DP_OP_425J2_127_3477_n2652), .Y(DP_OP_425J2_127_3477_n2620) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1849 ( .A1(DP_OP_425J2_127_3477_n2643), .A2(
        DP_OP_425J2_127_3477_n2652), .Y(DP_OP_425J2_127_3477_n2619) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1848 ( .A1(DP_OP_425J2_127_3477_n2650), .A2(
        DP_OP_422J2_124_3477_n2653), .Y(DP_OP_425J2_127_3477_n2618) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1847 ( .A1(DP_OP_425J2_127_3477_n2649), .A2(
        DP_OP_422J2_124_3477_n2653), .Y(DP_OP_425J2_127_3477_n2617) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1846 ( .A1(DP_OP_423J2_125_3477_n1986), .A2(
        DP_OP_424J2_126_3477_n2651), .Y(DP_OP_425J2_127_3477_n2616) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1845 ( .A1(DP_OP_424J2_126_3477_n2078), .A2(
        DP_OP_423J2_125_3477_n2649), .Y(DP_OP_425J2_127_3477_n2615) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1844 ( .A1(DP_OP_425J2_127_3477_n2646), .A2(
        DP_OP_422J2_124_3477_n2653), .Y(DP_OP_425J2_127_3477_n2614) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1843 ( .A1(DP_OP_423J2_125_3477_n1983), .A2(
        DP_OP_423J2_125_3477_n2649), .Y(DP_OP_425J2_127_3477_n2613) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1842 ( .A1(DP_OP_425J2_127_3477_n2644), .A2(
        DP_OP_423J2_125_3477_n2649), .Y(DP_OP_425J2_127_3477_n2612) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1841 ( .A1(DP_OP_425J2_127_3477_n2643), 
        .A2(DP_OP_422J2_124_3477_n2653), .Y(DP_OP_425J2_127_3477_n2611) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1822 ( .A1(DP_OP_424J2_126_3477_n2119), 
        .A2(DP_OP_425J2_127_3477_n2610), .Y(DP_OP_425J2_127_3477_n2592) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1821 ( .A1(DP_OP_424J2_126_3477_n2118), .A2(
        DP_OP_425J2_127_3477_n2610), .Y(DP_OP_425J2_127_3477_n2591) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1814 ( .A1(DP_OP_424J2_126_3477_n2119), 
        .A2(DP_OP_424J2_126_3477_n2609), .Y(DP_OP_425J2_127_3477_n2584) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1813 ( .A1(DP_OP_422J2_124_3477_n2731), .A2(
        DP_OP_424J2_126_3477_n2609), .Y(DP_OP_425J2_127_3477_n2583) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1806 ( .A1(DP_OP_424J2_126_3477_n2119), 
        .A2(n451), .Y(DP_OP_425J2_127_3477_n2576) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1805 ( .A1(DP_OP_422J2_124_3477_n2731), .A2(
        n451), .Y(DP_OP_425J2_127_3477_n2575) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1804 ( .A1(DP_OP_424J2_126_3477_n2125), .A2(
        DP_OP_424J2_126_3477_n2607), .Y(DP_OP_425J2_127_3477_n2574) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1803 ( .A1(DP_OP_424J2_126_3477_n2124), .A2(
        DP_OP_423J2_125_3477_n2605), .Y(DP_OP_425J2_127_3477_n2573) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1802 ( .A1(DP_OP_423J2_125_3477_n2030), .A2(
        DP_OP_424J2_126_3477_n2607), .Y(DP_OP_425J2_127_3477_n2572) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1801 ( .A1(DP_OP_423J2_125_3477_n2029), .A2(
        DP_OP_424J2_126_3477_n2607), .Y(DP_OP_425J2_127_3477_n2571) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1800 ( .A1(DP_OP_423J2_125_3477_n2028), .A2(
        DP_OP_423J2_125_3477_n2605), .Y(DP_OP_425J2_127_3477_n2570) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1799 ( .A1(DP_OP_424J2_126_3477_n2120), .A2(
        DP_OP_424J2_126_3477_n2607), .Y(DP_OP_425J2_127_3477_n2569) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1798 ( .A1(DP_OP_424J2_126_3477_n2119), .A2(
        DP_OP_422J2_124_3477_n2609), .Y(DP_OP_425J2_127_3477_n2568) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1797 ( .A1(DP_OP_422J2_124_3477_n2731), 
        .A2(DP_OP_423J2_125_3477_n2605), .Y(DP_OP_425J2_127_3477_n2567) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1779 ( .A1(DP_OP_425J2_127_3477_n2557), 
        .A2(DP_OP_425J2_127_3477_n2566), .Y(DP_OP_425J2_127_3477_n2549) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1778 ( .A1(DP_OP_424J2_126_3477_n2163), 
        .A2(DP_OP_425J2_127_3477_n2566), .Y(DP_OP_425J2_127_3477_n2548) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1777 ( .A1(DP_OP_425J2_127_3477_n2555), .A2(
        DP_OP_425J2_127_3477_n2566), .Y(DP_OP_425J2_127_3477_n2547) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1770 ( .A1(DP_OP_422J2_124_3477_n2690), 
        .A2(DP_OP_425J2_127_3477_n2565), .Y(DP_OP_425J2_127_3477_n2540) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1769 ( .A1(DP_OP_425J2_127_3477_n2555), .A2(
        DP_OP_425J2_127_3477_n2565), .Y(DP_OP_425J2_127_3477_n2539) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1762 ( .A1(DP_OP_422J2_124_3477_n2690), 
        .A2(DP_OP_425J2_127_3477_n2564), .Y(DP_OP_425J2_127_3477_n2532) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1761 ( .A1(DP_OP_425J2_127_3477_n2555), .A2(
        DP_OP_425J2_127_3477_n2564), .Y(DP_OP_425J2_127_3477_n2531) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1760 ( .A1(DP_OP_422J2_124_3477_n2696), .A2(
        DP_OP_425J2_127_3477_n2563), .Y(DP_OP_425J2_127_3477_n2530) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1759 ( .A1(DP_OP_422J2_124_3477_n2695), .A2(
        DP_OP_425J2_127_3477_n2563), .Y(DP_OP_425J2_127_3477_n2529) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1758 ( .A1(DP_OP_423J2_125_3477_n2074), .A2(
        DP_OP_425J2_127_3477_n2563), .Y(DP_OP_425J2_127_3477_n2528) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1757 ( .A1(DP_OP_425J2_127_3477_n2559), .A2(
        DP_OP_425J2_127_3477_n2563), .Y(DP_OP_425J2_127_3477_n2527) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1756 ( .A1(DP_OP_425J2_127_3477_n2558), .A2(
        DP_OP_425J2_127_3477_n2563), .Y(DP_OP_425J2_127_3477_n2526) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1755 ( .A1(DP_OP_425J2_127_3477_n2557), .A2(
        DP_OP_425J2_127_3477_n2563), .Y(DP_OP_425J2_127_3477_n2525) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1754 ( .A1(DP_OP_424J2_126_3477_n2163), .A2(
        DP_OP_425J2_127_3477_n2563), .Y(DP_OP_425J2_127_3477_n2524) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1753 ( .A1(DP_OP_425J2_127_3477_n2555), 
        .A2(DP_OP_425J2_127_3477_n2563), .Y(DP_OP_425J2_127_3477_n2523) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1734 ( .A1(DP_OP_422J2_124_3477_n2646), 
        .A2(DP_OP_424J2_126_3477_n2522), .Y(DP_OP_425J2_127_3477_n2504) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1733 ( .A1(DP_OP_425J2_127_3477_n2511), .A2(
        DP_OP_424J2_126_3477_n2522), .Y(DP_OP_425J2_127_3477_n2503) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1726 ( .A1(DP_OP_423J2_125_3477_n2114), 
        .A2(DP_OP_422J2_124_3477_n2523), .Y(DP_OP_425J2_127_3477_n2496) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1725 ( .A1(DP_OP_425J2_127_3477_n2511), .A2(
        DP_OP_422J2_124_3477_n2523), .Y(DP_OP_425J2_127_3477_n2495) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1718 ( .A1(DP_OP_422J2_124_3477_n2646), 
        .A2(n444), .Y(DP_OP_425J2_127_3477_n2488) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1717 ( .A1(DP_OP_425J2_127_3477_n2511), .A2(
        DP_OP_422J2_124_3477_n2522), .Y(DP_OP_425J2_127_3477_n2487) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1716 ( .A1(DP_OP_425J2_127_3477_n2518), .A2(
        DP_OP_425J2_127_3477_n2519), .Y(DP_OP_425J2_127_3477_n2486) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1715 ( .A1(DP_OP_422J2_124_3477_n2651), .A2(
        DP_OP_425J2_127_3477_n2519), .Y(DP_OP_425J2_127_3477_n2485) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1714 ( .A1(DP_OP_424J2_126_3477_n2211), .A2(
        DP_OP_425J2_127_3477_n2519), .Y(DP_OP_425J2_127_3477_n2484) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1713 ( .A1(DP_OP_423J2_125_3477_n2117), .A2(
        DP_OP_425J2_127_3477_n2519), .Y(DP_OP_425J2_127_3477_n2483) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1712 ( .A1(DP_OP_422J2_124_3477_n2648), .A2(
        DP_OP_425J2_127_3477_n2519), .Y(DP_OP_425J2_127_3477_n2482) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1711 ( .A1(DP_OP_423J2_125_3477_n2115), .A2(
        DP_OP_425J2_127_3477_n2519), .Y(DP_OP_425J2_127_3477_n2481) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1710 ( .A1(DP_OP_423J2_125_3477_n2114), .A2(
        DP_OP_425J2_127_3477_n2519), .Y(DP_OP_425J2_127_3477_n2480) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1709 ( .A1(DP_OP_425J2_127_3477_n2511), 
        .A2(DP_OP_425J2_127_3477_n2519), .Y(DP_OP_425J2_127_3477_n2479) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1691 ( .A1(DP_OP_425J2_127_3477_n2469), 
        .A2(DP_OP_423J2_125_3477_n2476), .Y(DP_OP_425J2_127_3477_n2461) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1690 ( .A1(DP_OP_423J2_125_3477_n2158), 
        .A2(DP_OP_424J2_126_3477_n2478), .Y(DP_OP_425J2_127_3477_n2460) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1689 ( .A1(DP_OP_423J2_125_3477_n2157), .A2(
        DP_OP_422J2_124_3477_n2480), .Y(DP_OP_425J2_127_3477_n2459) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1682 ( .A1(DP_OP_423J2_125_3477_n2158), 
        .A2(DP_OP_425J2_127_3477_n2477), .Y(DP_OP_425J2_127_3477_n2452) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1681 ( .A1(DP_OP_423J2_125_3477_n2157), .A2(
        DP_OP_425J2_127_3477_n2477), .Y(DP_OP_425J2_127_3477_n2451) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1674 ( .A1(DP_OP_423J2_125_3477_n2158), 
        .A2(DP_OP_425J2_127_3477_n2476), .Y(DP_OP_425J2_127_3477_n2444) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1673 ( .A1(DP_OP_423J2_125_3477_n2157), .A2(
        DP_OP_425J2_127_3477_n2476), .Y(DP_OP_425J2_127_3477_n2443) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1672 ( .A1(DP_OP_423J2_125_3477_n2164), .A2(
        DP_OP_425J2_127_3477_n2475), .Y(DP_OP_425J2_127_3477_n2442) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1671 ( .A1(DP_OP_423J2_125_3477_n2163), .A2(
        DP_OP_425J2_127_3477_n2475), .Y(DP_OP_425J2_127_3477_n2441) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1670 ( .A1(DP_OP_425J2_127_3477_n2472), .A2(
        DP_OP_425J2_127_3477_n2475), .Y(DP_OP_425J2_127_3477_n2440) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1669 ( .A1(DP_OP_423J2_125_3477_n2161), .A2(
        DP_OP_425J2_127_3477_n2475), .Y(DP_OP_425J2_127_3477_n2439) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1668 ( .A1(DP_OP_423J2_125_3477_n2160), .A2(
        DP_OP_425J2_127_3477_n2475), .Y(DP_OP_425J2_127_3477_n2438) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1667 ( .A1(DP_OP_425J2_127_3477_n2469), .A2(
        DP_OP_425J2_127_3477_n2475), .Y(DP_OP_425J2_127_3477_n2437) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1666 ( .A1(DP_OP_423J2_125_3477_n2158), .A2(
        DP_OP_425J2_127_3477_n2475), .Y(DP_OP_425J2_127_3477_n2436) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1665 ( .A1(DP_OP_423J2_125_3477_n2157), 
        .A2(DP_OP_425J2_127_3477_n2475), .Y(DP_OP_425J2_127_3477_n2435) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1646 ( .A1(DP_OP_425J2_127_3477_n2424), 
        .A2(DP_OP_425J2_127_3477_n2434), .Y(DP_OP_425J2_127_3477_n2416) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1645 ( .A1(DP_OP_425J2_127_3477_n2423), .A2(
        DP_OP_425J2_127_3477_n2434), .Y(DP_OP_425J2_127_3477_n2415) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1638 ( .A1(DP_OP_425J2_127_3477_n2424), 
        .A2(DP_OP_425J2_127_3477_n2433), .Y(DP_OP_425J2_127_3477_n2408) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1637 ( .A1(DP_OP_425J2_127_3477_n2423), .A2(
        DP_OP_425J2_127_3477_n2433), .Y(DP_OP_425J2_127_3477_n2407) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1630 ( .A1(DP_OP_425J2_127_3477_n2424), 
        .A2(DP_OP_423J2_125_3477_n2430), .Y(DP_OP_425J2_127_3477_n2400) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1629 ( .A1(DP_OP_425J2_127_3477_n2423), .A2(
        DP_OP_423J2_125_3477_n2430), .Y(DP_OP_425J2_127_3477_n2399) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1628 ( .A1(DP_OP_425J2_127_3477_n2430), .A2(
        DP_OP_425J2_127_3477_n2431), .Y(DP_OP_425J2_127_3477_n2398) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1627 ( .A1(DP_OP_425J2_127_3477_n2429), .A2(
        DP_OP_425J2_127_3477_n2431), .Y(DP_OP_425J2_127_3477_n2397) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1626 ( .A1(DP_OP_425J2_127_3477_n2428), .A2(
        DP_OP_425J2_127_3477_n2431), .Y(DP_OP_425J2_127_3477_n2396) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1625 ( .A1(DP_OP_425J2_127_3477_n2427), .A2(
        DP_OP_425J2_127_3477_n2431), .Y(DP_OP_425J2_127_3477_n2395) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1624 ( .A1(DP_OP_422J2_124_3477_n2560), .A2(
        DP_OP_425J2_127_3477_n2431), .Y(DP_OP_425J2_127_3477_n2394) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1623 ( .A1(DP_OP_422J2_124_3477_n2559), .A2(
        DP_OP_425J2_127_3477_n2431), .Y(DP_OP_425J2_127_3477_n2393) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1622 ( .A1(DP_OP_425J2_127_3477_n2424), .A2(
        DP_OP_425J2_127_3477_n2431), .Y(DP_OP_425J2_127_3477_n2392) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1621 ( .A1(DP_OP_425J2_127_3477_n2423), 
        .A2(DP_OP_425J2_127_3477_n2431), .Y(DP_OP_425J2_127_3477_n2391) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1601 ( .A1(DP_OP_424J2_126_3477_n2338), .A2(
        DP_OP_424J2_126_3477_n2390), .Y(DP_OP_425J2_127_3477_n2371) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1595 ( .A1(DP_OP_425J2_127_3477_n2381), 
        .A2(DP_OP_424J2_126_3477_n2389), .Y(DP_OP_425J2_127_3477_n2365) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1593 ( .A1(DP_OP_424J2_126_3477_n2338), .A2(
        DP_OP_422J2_124_3477_n2391), .Y(DP_OP_425J2_127_3477_n2363) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1586 ( .A1(DP_OP_422J2_124_3477_n2514), 
        .A2(DP_OP_422J2_124_3477_n2390), .Y(DP_OP_425J2_127_3477_n2356) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1585 ( .A1(DP_OP_422J2_124_3477_n2513), .A2(
        DP_OP_422J2_124_3477_n2390), .Y(DP_OP_425J2_127_3477_n2355) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1584 ( .A1(DP_OP_425J2_127_3477_n2386), .A2(
        DP_OP_425J2_127_3477_n2387), .Y(DP_OP_425J2_127_3477_n1579) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1583 ( .A1(DP_OP_424J2_126_3477_n2344), .A2(
        DP_OP_425J2_127_3477_n2387), .Y(DP_OP_425J2_127_3477_n2354) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1582 ( .A1(DP_OP_425J2_127_3477_n2384), .A2(
        DP_OP_425J2_127_3477_n2387), .Y(DP_OP_425J2_127_3477_n2353) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1581 ( .A1(DP_OP_425J2_127_3477_n2383), .A2(
        DP_OP_425J2_127_3477_n2387), .Y(DP_OP_425J2_127_3477_n2352) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1580 ( .A1(DP_OP_425J2_127_3477_n2382), .A2(
        DP_OP_425J2_127_3477_n2387), .Y(DP_OP_425J2_127_3477_n2351) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1579 ( .A1(DP_OP_425J2_127_3477_n2381), .A2(
        DP_OP_425J2_127_3477_n2387), .Y(DP_OP_425J2_127_3477_n671) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1578 ( .A1(DP_OP_422J2_124_3477_n2514), .A2(
        DP_OP_425J2_127_3477_n2387), .Y(DP_OP_425J2_127_3477_n2350) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1577 ( .A1(DP_OP_424J2_126_3477_n2338), 
        .A2(DP_OP_425J2_127_3477_n2387), .Y(DP_OP_425J2_127_3477_n361) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1559 ( .A1(DP_OP_425J2_127_3477_n2340), 
        .A2(DP_OP_425J2_127_3477_n2349), .Y(DP_OP_425J2_127_3477_n2332) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1558 ( .A1(DP_OP_425J2_127_3477_n2339), 
        .A2(DP_OP_425J2_127_3477_n2349), .Y(DP_OP_425J2_127_3477_n2331) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1557 ( .A1(DP_OP_424J2_126_3477_n2423), .A2(
        DP_OP_425J2_127_3477_n2349), .Y(DP_OP_425J2_127_3477_n2330) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1550 ( .A1(DP_OP_425J2_127_3477_n2339), 
        .A2(DP_OP_425J2_127_3477_n2348), .Y(DP_OP_425J2_127_3477_n2323) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1549 ( .A1(DP_OP_423J2_125_3477_n2509), .A2(
        DP_OP_425J2_127_3477_n2348), .Y(DP_OP_425J2_127_3477_n2322) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1542 ( .A1(DP_OP_425J2_127_3477_n2339), 
        .A2(DP_OP_425J2_127_3477_n2347), .Y(DP_OP_425J2_127_3477_n2315) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1541 ( .A1(DP_OP_423J2_125_3477_n2509), .A2(
        DP_OP_425J2_127_3477_n2347), .Y(DP_OP_425J2_127_3477_n2314) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1540 ( .A1(DP_OP_424J2_126_3477_n2430), .A2(
        DP_OP_425J2_127_3477_n2346), .Y(DP_OP_425J2_127_3477_n2313) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1539 ( .A1(DP_OP_422J2_124_3477_n2211), .A2(
        DP_OP_425J2_127_3477_n2346), .Y(DP_OP_425J2_127_3477_n2312) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1538 ( .A1(DP_OP_422J2_124_3477_n2210), .A2(
        DP_OP_425J2_127_3477_n2346), .Y(DP_OP_425J2_127_3477_n2311) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1537 ( .A1(DP_OP_425J2_127_3477_n2342), .A2(
        DP_OP_425J2_127_3477_n2346), .Y(DP_OP_425J2_127_3477_n2310) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1536 ( .A1(DP_OP_425J2_127_3477_n2341), .A2(
        DP_OP_425J2_127_3477_n2346), .Y(DP_OP_425J2_127_3477_n2309) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1535 ( .A1(DP_OP_425J2_127_3477_n2340), .A2(
        DP_OP_425J2_127_3477_n2346), .Y(DP_OP_425J2_127_3477_n2308) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1534 ( .A1(DP_OP_425J2_127_3477_n2339), .A2(
        DP_OP_425J2_127_3477_n2346), .Y(DP_OP_425J2_127_3477_n2307) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1533 ( .A1(DP_OP_423J2_125_3477_n2509), 
        .A2(DP_OP_425J2_127_3477_n2346), .Y(DP_OP_425J2_127_3477_n2306) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1514 ( .A1(DP_OP_423J2_125_3477_n2554), 
        .A2(DP_OP_425J2_127_3477_n2305), .Y(DP_OP_425J2_127_3477_n2287) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1513 ( .A1(DP_OP_425J2_127_3477_n2294), .A2(
        DP_OP_425J2_127_3477_n2305), .Y(DP_OP_425J2_127_3477_n2286) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1506 ( .A1(DP_OP_423J2_125_3477_n2554), 
        .A2(DP_OP_425J2_127_3477_n2304), .Y(DP_OP_425J2_127_3477_n2279) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1505 ( .A1(DP_OP_425J2_127_3477_n2294), .A2(
        DP_OP_425J2_127_3477_n2304), .Y(DP_OP_425J2_127_3477_n2278) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1498 ( .A1(DP_OP_423J2_125_3477_n2554), 
        .A2(DP_OP_423J2_125_3477_n2298), .Y(DP_OP_425J2_127_3477_n2271) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1497 ( .A1(DP_OP_425J2_127_3477_n2294), .A2(
        DP_OP_422J2_124_3477_n2302), .Y(DP_OP_425J2_127_3477_n2270) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1496 ( .A1(DP_OP_422J2_124_3477_n2168), .A2(
        DP_OP_425J2_127_3477_n2302), .Y(DP_OP_425J2_127_3477_n2269) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1495 ( .A1(DP_OP_425J2_127_3477_n2300), .A2(
        DP_OP_425J2_127_3477_n2302), .Y(DP_OP_425J2_127_3477_n2268) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1494 ( .A1(DP_OP_423J2_125_3477_n2558), .A2(
        DP_OP_425J2_127_3477_n2302), .Y(DP_OP_425J2_127_3477_n2267) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1493 ( .A1(DP_OP_424J2_126_3477_n2471), .A2(
        DP_OP_425J2_127_3477_n2302), .Y(DP_OP_425J2_127_3477_n2266) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1492 ( .A1(DP_OP_425J2_127_3477_n2297), .A2(
        DP_OP_425J2_127_3477_n2302), .Y(DP_OP_425J2_127_3477_n2265) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1491 ( .A1(DP_OP_425J2_127_3477_n2296), .A2(
        DP_OP_425J2_127_3477_n2302), .Y(DP_OP_425J2_127_3477_n2264) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1490 ( .A1(DP_OP_422J2_124_3477_n2162), .A2(
        DP_OP_425J2_127_3477_n2302), .Y(DP_OP_425J2_127_3477_n2263) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1489 ( .A1(DP_OP_425J2_127_3477_n2294), 
        .A2(DP_OP_425J2_127_3477_n2302), .Y(DP_OP_425J2_127_3477_n2262) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1470 ( .A1(DP_OP_424J2_126_3477_n2512), 
        .A2(DP_OP_425J2_127_3477_n2261), .Y(DP_OP_425J2_127_3477_n2243) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1469 ( .A1(DP_OP_425J2_127_3477_n2250), .A2(
        DP_OP_425J2_127_3477_n2261), .Y(DP_OP_425J2_127_3477_n2242) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1462 ( .A1(DP_OP_422J2_124_3477_n2118), 
        .A2(DP_OP_425J2_127_3477_n2260), .Y(DP_OP_425J2_127_3477_n2235) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1461 ( .A1(DP_OP_425J2_127_3477_n2250), .A2(
        DP_OP_425J2_127_3477_n2260), .Y(DP_OP_425J2_127_3477_n2234) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1453 ( .A1(DP_OP_425J2_127_3477_n2250), .A2(
        DP_OP_425J2_127_3477_n2259), .Y(DP_OP_425J2_127_3477_n2226) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1452 ( .A1(DP_OP_423J2_125_3477_n2604), .A2(
        DP_OP_422J2_124_3477_n2257), .Y(DP_OP_425J2_127_3477_n2225) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1451 ( .A1(DP_OP_423J2_125_3477_n2603), .A2(
        n450), .Y(DP_OP_425J2_127_3477_n2224) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1450 ( .A1(DP_OP_425J2_127_3477_n2255), .A2(
        n450), .Y(DP_OP_425J2_127_3477_n2223) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1449 ( .A1(DP_OP_422J2_124_3477_n2121), .A2(
        n450), .Y(DP_OP_425J2_127_3477_n2222) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1448 ( .A1(DP_OP_423J2_125_3477_n2600), .A2(
        DP_OP_424J2_126_3477_n2258), .Y(DP_OP_425J2_127_3477_n2221) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1447 ( .A1(DP_OP_425J2_127_3477_n2252), .A2(
        n450), .Y(DP_OP_425J2_127_3477_n2220) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1446 ( .A1(DP_OP_424J2_126_3477_n2512), .A2(
        n450), .Y(DP_OP_425J2_127_3477_n2219) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1445 ( .A1(DP_OP_425J2_127_3477_n2250), 
        .A2(n450), .Y(DP_OP_425J2_127_3477_n2218) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1426 ( .A1(DP_OP_423J2_125_3477_n2642), 
        .A2(DP_OP_425J2_127_3477_n2217), .Y(DP_OP_425J2_127_3477_n2199) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1425 ( .A1(DP_OP_424J2_126_3477_n2555), .A2(
        DP_OP_425J2_127_3477_n2217), .Y(DP_OP_425J2_127_3477_n2198) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1417 ( .A1(DP_OP_424J2_126_3477_n2555), .A2(
        DP_OP_423J2_125_3477_n2211), .Y(DP_OP_425J2_127_3477_n2190) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1410 ( .A1(DP_OP_423J2_125_3477_n2642), 
        .A2(DP_OP_425J2_127_3477_n2215), .Y(DP_OP_425J2_127_3477_n2183) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1409 ( .A1(DP_OP_422J2_124_3477_n2073), .A2(
        DP_OP_425J2_127_3477_n2215), .Y(DP_OP_425J2_127_3477_n2182) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1408 ( .A1(DP_OP_425J2_127_3477_n2213), .A2(
        DP_OP_425J2_127_3477_n2214), .Y(DP_OP_425J2_127_3477_n2181) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1407 ( .A1(DP_OP_423J2_125_3477_n2647), .A2(
        DP_OP_425J2_127_3477_n2214), .Y(DP_OP_425J2_127_3477_n2180) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1406 ( .A1(DP_OP_422J2_124_3477_n2078), .A2(
        DP_OP_425J2_127_3477_n2214), .Y(DP_OP_425J2_127_3477_n2179) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1405 ( .A1(DP_OP_424J2_126_3477_n2559), .A2(
        DP_OP_425J2_127_3477_n2214), .Y(DP_OP_425J2_127_3477_n2178) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1404 ( .A1(DP_OP_425J2_127_3477_n2209), .A2(
        DP_OP_425J2_127_3477_n2214), .Y(DP_OP_425J2_127_3477_n2177) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1403 ( .A1(DP_OP_424J2_126_3477_n2557), .A2(
        DP_OP_425J2_127_3477_n2214), .Y(DP_OP_425J2_127_3477_n2176) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1402 ( .A1(DP_OP_423J2_125_3477_n2642), .A2(
        DP_OP_425J2_127_3477_n2214), .Y(DP_OP_425J2_127_3477_n2175) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1401 ( .A1(DP_OP_424J2_126_3477_n2555), 
        .A2(DP_OP_425J2_127_3477_n2214), .Y(DP_OP_425J2_127_3477_n2174) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1382 ( .A1(DP_OP_425J2_127_3477_n2163), 
        .A2(DP_OP_425J2_127_3477_n2173), .Y(DP_OP_425J2_127_3477_n2155) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1381 ( .A1(DP_OP_425J2_127_3477_n2162), .A2(
        DP_OP_425J2_127_3477_n2173), .Y(DP_OP_425J2_127_3477_n2154) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1374 ( .A1(DP_OP_425J2_127_3477_n2163), 
        .A2(DP_OP_425J2_127_3477_n2172), .Y(DP_OP_425J2_127_3477_n2147) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1373 ( .A1(DP_OP_425J2_127_3477_n2162), .A2(
        DP_OP_425J2_127_3477_n2172), .Y(DP_OP_425J2_127_3477_n2146) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1366 ( .A1(DP_OP_425J2_127_3477_n2163), 
        .A2(n452), .Y(DP_OP_425J2_127_3477_n2139) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1365 ( .A1(DP_OP_425J2_127_3477_n2162), .A2(
        n452), .Y(DP_OP_425J2_127_3477_n2138) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1364 ( .A1(DP_OP_425J2_127_3477_n2169), .A2(
        DP_OP_423J2_125_3477_n2165), .Y(DP_OP_425J2_127_3477_n2137) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1363 ( .A1(DP_OP_425J2_127_3477_n2168), .A2(
        DP_OP_423J2_125_3477_n2165), .Y(DP_OP_425J2_127_3477_n2136) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1362 ( .A1(DP_OP_423J2_125_3477_n2690), .A2(
        DP_OP_422J2_124_3477_n2169), .Y(DP_OP_425J2_127_3477_n2135) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1361 ( .A1(DP_OP_425J2_127_3477_n2166), .A2(
        DP_OP_424J2_126_3477_n2170), .Y(DP_OP_425J2_127_3477_n2134) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1360 ( .A1(DP_OP_423J2_125_3477_n2688), .A2(
        DP_OP_422J2_124_3477_n2169), .Y(DP_OP_425J2_127_3477_n2133) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1359 ( .A1(DP_OP_425J2_127_3477_n2164), .A2(
        DP_OP_424J2_126_3477_n2170), .Y(DP_OP_425J2_127_3477_n2132) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1358 ( .A1(DP_OP_425J2_127_3477_n2163), .A2(
        DP_OP_422J2_124_3477_n2169), .Y(DP_OP_425J2_127_3477_n2131) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1357 ( .A1(DP_OP_425J2_127_3477_n2162), 
        .A2(DP_OP_423J2_125_3477_n2165), .Y(DP_OP_425J2_127_3477_n2130) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1337 ( .A1(DP_OP_425J2_127_3477_n2118), .A2(
        DP_OP_425J2_127_3477_n2129), .Y(DP_OP_425J2_127_3477_n2110) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1330 ( .A1(DP_OP_425J2_127_3477_n2119), 
        .A2(DP_OP_425J2_127_3477_n2128), .Y(DP_OP_425J2_127_3477_n2103) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1329 ( .A1(DP_OP_425J2_127_3477_n2118), .A2(
        DP_OP_425J2_127_3477_n2128), .Y(DP_OP_425J2_127_3477_n2102) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1322 ( .A1(DP_OP_425J2_127_3477_n2119), 
        .A2(DP_OP_425J2_127_3477_n2127), .Y(DP_OP_425J2_127_3477_n2095) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1321 ( .A1(DP_OP_425J2_127_3477_n2118), .A2(
        DP_OP_425J2_127_3477_n2127), .Y(DP_OP_425J2_127_3477_n2094) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1320 ( .A1(DP_OP_424J2_126_3477_n2650), .A2(
        DP_OP_425J2_127_3477_n2126), .Y(DP_OP_425J2_127_3477_n2093) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1319 ( .A1(DP_OP_424J2_126_3477_n2649), .A2(
        DP_OP_425J2_127_3477_n2126), .Y(DP_OP_425J2_127_3477_n2092) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1318 ( .A1(DP_OP_423J2_125_3477_n2731), .A2(
        DP_OP_425J2_127_3477_n2126), .Y(DP_OP_425J2_127_3477_n2091) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1317 ( .A1(DP_OP_425J2_127_3477_n2122), .A2(
        DP_OP_425J2_127_3477_n2126), .Y(DP_OP_425J2_127_3477_n2090) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1316 ( .A1(DP_OP_422J2_124_3477_n1989), .A2(
        DP_OP_425J2_127_3477_n2126), .Y(DP_OP_425J2_127_3477_n2089) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1315 ( .A1(DP_OP_425J2_127_3477_n2120), .A2(
        DP_OP_425J2_127_3477_n2126), .Y(DP_OP_425J2_127_3477_n2088) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1314 ( .A1(DP_OP_425J2_127_3477_n2119), .A2(
        DP_OP_425J2_127_3477_n2126), .Y(DP_OP_425J2_127_3477_n2087) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1313 ( .A1(DP_OP_425J2_127_3477_n2118), 
        .A2(DP_OP_425J2_127_3477_n2126), .Y(DP_OP_425J2_127_3477_n2086) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1294 ( .A1(DP_OP_425J2_127_3477_n2075), 
        .A2(n441), .Y(DP_OP_425J2_127_3477_n2067) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1293 ( .A1(DP_OP_425J2_127_3477_n2074), .A2(
        n441), .Y(DP_OP_425J2_127_3477_n2066) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1286 ( .A1(DP_OP_425J2_127_3477_n2075), 
        .A2(DP_OP_425J2_127_3477_n2084), .Y(DP_OP_425J2_127_3477_n2059) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1285 ( .A1(DP_OP_425J2_127_3477_n2074), .A2(
        DP_OP_425J2_127_3477_n2084), .Y(DP_OP_425J2_127_3477_n2058) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1277 ( .A1(DP_OP_425J2_127_3477_n2074), .A2(
        DP_OP_425J2_127_3477_n2083), .Y(DP_OP_425J2_127_3477_n2050) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1276 ( .A1(DP_OP_423J2_125_3477_n2777), .A2(
        DP_OP_424J2_126_3477_n2082), .Y(DP_OP_425J2_127_3477_n2049) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1275 ( .A1(DP_OP_423J2_125_3477_n2776), .A2(
        DP_OP_422J2_124_3477_n2081), .Y(DP_OP_425J2_127_3477_n2048) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1274 ( .A1(DP_OP_425J2_127_3477_n2079), .A2(
        DP_OP_424J2_126_3477_n2082), .Y(DP_OP_425J2_127_3477_n2047) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1273 ( .A1(DP_OP_425J2_127_3477_n2078), .A2(
        DP_OP_424J2_126_3477_n2082), .Y(DP_OP_425J2_127_3477_n2046) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1272 ( .A1(DP_OP_425J2_127_3477_n2077), .A2(
        DP_OP_422J2_124_3477_n2081), .Y(DP_OP_425J2_127_3477_n2045) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1271 ( .A1(DP_OP_423J2_125_3477_n2772), .A2(
        DP_OP_424J2_126_3477_n2082), .Y(DP_OP_425J2_127_3477_n2044) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1270 ( .A1(DP_OP_425J2_127_3477_n2075), .A2(
        DP_OP_424J2_126_3477_n2082), .Y(DP_OP_425J2_127_3477_n2043) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1269 ( .A1(DP_OP_425J2_127_3477_n2074), 
        .A2(DP_OP_422J2_124_3477_n2081), .Y(DP_OP_425J2_127_3477_n2042) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1250 ( .A1(DP_OP_422J2_124_3477_n1899), 
        .A2(DP_OP_425J2_127_3477_n2041), .Y(DP_OP_425J2_127_3477_n2023) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1249 ( .A1(DP_OP_424J2_126_3477_n2731), .A2(
        DP_OP_425J2_127_3477_n2041), .Y(DP_OP_425J2_127_3477_n2022) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1242 ( .A1(DP_OP_424J2_126_3477_n2732), 
        .A2(DP_OP_425J2_127_3477_n2040), .Y(DP_OP_425J2_127_3477_n2015) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1241 ( .A1(DP_OP_424J2_126_3477_n2731), .A2(
        DP_OP_425J2_127_3477_n2040), .Y(DP_OP_425J2_127_3477_n2014) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1234 ( .A1(DP_OP_422J2_124_3477_n1899), 
        .A2(DP_OP_425J2_127_3477_n2039), .Y(DP_OP_425J2_127_3477_n2007) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1233 ( .A1(DP_OP_422J2_124_3477_n1898), .A2(
        DP_OP_425J2_127_3477_n2039), .Y(DP_OP_425J2_127_3477_n2006) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1232 ( .A1(DP_OP_422J2_124_3477_n1905), .A2(
        DP_OP_424J2_126_3477_n2038), .Y(DP_OP_425J2_127_3477_n2005) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1231 ( .A1(DP_OP_424J2_126_3477_n2737), .A2(
        DP_OP_424J2_126_3477_n2038), .Y(DP_OP_425J2_127_3477_n2004) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1230 ( .A1(DP_OP_424J2_126_3477_n2736), .A2(
        DP_OP_424J2_126_3477_n2038), .Y(DP_OP_425J2_127_3477_n2003) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1229 ( .A1(DP_OP_422J2_124_3477_n1902), .A2(
        DP_OP_423J2_125_3477_n2033), .Y(DP_OP_425J2_127_3477_n2002) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1228 ( .A1(DP_OP_425J2_127_3477_n2033), .A2(
        DP_OP_423J2_125_3477_n2033), .Y(DP_OP_425J2_127_3477_n2001) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1227 ( .A1(DP_OP_424J2_126_3477_n2733), .A2(
        DP_OP_424J2_126_3477_n2038), .Y(DP_OP_425J2_127_3477_n2000) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1226 ( .A1(DP_OP_424J2_126_3477_n2732), .A2(
        DP_OP_423J2_125_3477_n2033), .Y(DP_OP_425J2_127_3477_n1999) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1225 ( .A1(DP_OP_424J2_126_3477_n2731), 
        .A2(DP_OP_424J2_126_3477_n2038), .Y(DP_OP_425J2_127_3477_n1998) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1206 ( .A1(DP_OP_423J2_125_3477_n2859), 
        .A2(DP_OP_425J2_127_3477_n1997), .Y(DP_OP_425J2_127_3477_n1979) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1205 ( .A1(DP_OP_422J2_124_3477_n1854), .A2(
        DP_OP_425J2_127_3477_n1997), .Y(DP_OP_425J2_127_3477_n1978) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1197 ( .A1(DP_OP_422J2_124_3477_n1854), .A2(
        DP_OP_423J2_125_3477_n1991), .Y(DP_OP_425J2_127_3477_n1970) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1189 ( .A1(DP_OP_422J2_124_3477_n1854), .A2(
        DP_OP_425J2_127_3477_n1995), .Y(DP_OP_425J2_127_3477_n1962) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1188 ( .A1(DP_OP_423J2_125_3477_n2865), .A2(
        DP_OP_424J2_126_3477_n1994), .Y(DP_OP_425J2_127_3477_n1961) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1187 ( .A1(DP_OP_425J2_127_3477_n1992), .A2(
        DP_OP_422J2_124_3477_n1994), .Y(DP_OP_425J2_127_3477_n1960) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1186 ( .A1(DP_OP_425J2_127_3477_n1991), .A2(
        DP_OP_424J2_126_3477_n1994), .Y(DP_OP_425J2_127_3477_n1959) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1185 ( .A1(DP_OP_425J2_127_3477_n1990), .A2(
        DP_OP_422J2_124_3477_n1994), .Y(DP_OP_425J2_127_3477_n1958) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1184 ( .A1(DP_OP_425J2_127_3477_n1989), .A2(
        DP_OP_424J2_126_3477_n1994), .Y(DP_OP_425J2_127_3477_n1957) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1183 ( .A1(DP_OP_423J2_125_3477_n2860), .A2(
        DP_OP_424J2_126_3477_n1994), .Y(DP_OP_425J2_127_3477_n1956) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1182 ( .A1(DP_OP_423J2_125_3477_n2859), .A2(
        DP_OP_424J2_126_3477_n1994), .Y(DP_OP_425J2_127_3477_n1955) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1181 ( .A1(DP_OP_424J2_126_3477_n2775), 
        .A2(DP_OP_422J2_124_3477_n1994), .Y(DP_OP_425J2_127_3477_n1954) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1162 ( .A1(DP_OP_423J2_125_3477_n2903), 
        .A2(DP_OP_425J2_127_3477_n1953), .Y(DP_OP_425J2_127_3477_n1935) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1161 ( .A1(DP_OP_423J2_125_3477_n2902), .A2(
        DP_OP_425J2_127_3477_n1953), .Y(DP_OP_425J2_127_3477_n1934) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1154 ( .A1(DP_OP_423J2_125_3477_n2903), 
        .A2(DP_OP_424J2_126_3477_n1952), .Y(DP_OP_425J2_127_3477_n1927) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1153 ( .A1(DP_OP_423J2_125_3477_n2902), .A2(
        DP_OP_424J2_126_3477_n1952), .Y(DP_OP_425J2_127_3477_n1926) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1146 ( .A1(DP_OP_423J2_125_3477_n2903), 
        .A2(DP_OP_425J2_127_3477_n1951), .Y(DP_OP_425J2_127_3477_n1919) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1145 ( .A1(DP_OP_423J2_125_3477_n2902), .A2(
        DP_OP_425J2_127_3477_n1951), .Y(DP_OP_425J2_127_3477_n1918) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1144 ( .A1(DP_OP_423J2_125_3477_n2909), .A2(
        DP_OP_425J2_127_3477_n1950), .Y(DP_OP_425J2_127_3477_n1917) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1143 ( .A1(DP_OP_423J2_125_3477_n2908), .A2(
        DP_OP_425J2_127_3477_n1950), .Y(DP_OP_425J2_127_3477_n1916) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1142 ( .A1(DP_OP_423J2_125_3477_n2907), .A2(
        DP_OP_425J2_127_3477_n1950), .Y(DP_OP_425J2_127_3477_n1915) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1141 ( .A1(DP_OP_423J2_125_3477_n2906), .A2(
        DP_OP_425J2_127_3477_n1950), .Y(DP_OP_425J2_127_3477_n1914) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1140 ( .A1(DP_OP_425J2_127_3477_n1945), .A2(
        DP_OP_425J2_127_3477_n1950), .Y(DP_OP_425J2_127_3477_n1913) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1139 ( .A1(DP_OP_423J2_125_3477_n2904), .A2(
        DP_OP_425J2_127_3477_n1950), .Y(DP_OP_425J2_127_3477_n1912) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1138 ( .A1(DP_OP_423J2_125_3477_n2903), .A2(
        DP_OP_425J2_127_3477_n1950), .Y(DP_OP_425J2_127_3477_n1911) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1137 ( .A1(DP_OP_423J2_125_3477_n2902), 
        .A2(DP_OP_425J2_127_3477_n1950), .Y(DP_OP_425J2_127_3477_n1910) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1118 ( .A1(DP_OP_424J2_126_3477_n2864), 
        .A2(DP_OP_424J2_126_3477_n1909), .Y(DP_OP_425J2_127_3477_n1891) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1117 ( .A1(DP_OP_424J2_126_3477_n2863), .A2(
        DP_OP_424J2_126_3477_n1909), .Y(DP_OP_425J2_127_3477_n1890) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1110 ( .A1(DP_OP_424J2_126_3477_n2864), 
        .A2(n449), .Y(DP_OP_425J2_127_3477_n1883) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1109 ( .A1(DP_OP_424J2_126_3477_n2863), .A2(
        n449), .Y(DP_OP_425J2_127_3477_n1882) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1102 ( .A1(DP_OP_424J2_126_3477_n2864), 
        .A2(DP_OP_425J2_127_3477_n1907), .Y(DP_OP_425J2_127_3477_n1875) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1101 ( .A1(DP_OP_424J2_126_3477_n2863), .A2(
        DP_OP_425J2_127_3477_n1907), .Y(DP_OP_425J2_127_3477_n1874) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1100 ( .A1(DP_OP_425J2_127_3477_n1905), .A2(
        DP_OP_423J2_125_3477_n1901), .Y(DP_OP_425J2_127_3477_n1873) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1099 ( .A1(DP_OP_424J2_126_3477_n2869), .A2(
        DP_OP_423J2_125_3477_n1901), .Y(DP_OP_425J2_127_3477_n1872) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1098 ( .A1(DP_OP_425J2_127_3477_n1903), .A2(
        DP_OP_423J2_125_3477_n1901), .Y(DP_OP_425J2_127_3477_n1871) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1097 ( .A1(DP_OP_424J2_126_3477_n2867), .A2(
        DP_OP_424J2_126_3477_n1906), .Y(DP_OP_425J2_127_3477_n1870) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1096 ( .A1(DP_OP_425J2_127_3477_n1901), .A2(
        DP_OP_424J2_126_3477_n1906), .Y(DP_OP_425J2_127_3477_n1869) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1095 ( .A1(DP_OP_424J2_126_3477_n2865), .A2(
        DP_OP_423J2_125_3477_n1901), .Y(DP_OP_425J2_127_3477_n1868) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1094 ( .A1(DP_OP_424J2_126_3477_n2864), .A2(
        DP_OP_422J2_124_3477_n1906), .Y(DP_OP_425J2_127_3477_n1867) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1093 ( .A1(DP_OP_424J2_126_3477_n2863), 
        .A2(DP_OP_424J2_126_3477_n1906), .Y(DP_OP_425J2_127_3477_n1866) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1074 ( .A1(DP_OP_425J2_127_3477_n1855), 
        .A2(DP_OP_424J2_126_3477_n1865), .Y(DP_OP_425J2_127_3477_n1847) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1073 ( .A1(DP_OP_425J2_127_3477_n1854), .A2(
        DP_OP_423J2_125_3477_n1860), .Y(DP_OP_425J2_127_3477_n1846) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1066 ( .A1(DP_OP_425J2_127_3477_n1855), 
        .A2(DP_OP_425J2_127_3477_n1864), .Y(DP_OP_425J2_127_3477_n1839) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1065 ( .A1(DP_OP_425J2_127_3477_n1854), .A2(
        DP_OP_425J2_127_3477_n1864), .Y(DP_OP_425J2_127_3477_n1838) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1058 ( .A1(DP_OP_425J2_127_3477_n1855), 
        .A2(DP_OP_425J2_127_3477_n1863), .Y(DP_OP_425J2_127_3477_n1831) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1057 ( .A1(DP_OP_425J2_127_3477_n1854), .A2(
        DP_OP_425J2_127_3477_n1863), .Y(DP_OP_425J2_127_3477_n1830) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1056 ( .A1(DP_OP_425J2_127_3477_n1861), .A2(
        DP_OP_425J2_127_3477_n1862), .Y(DP_OP_425J2_127_3477_n1829) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1055 ( .A1(DP_OP_425J2_127_3477_n1860), .A2(
        DP_OP_425J2_127_3477_n1862), .Y(DP_OP_425J2_127_3477_n1828) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1054 ( .A1(DP_OP_424J2_126_3477_n2912), .A2(
        DP_OP_425J2_127_3477_n1862), .Y(DP_OP_425J2_127_3477_n1827) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1053 ( .A1(DP_OP_425J2_127_3477_n1858), .A2(
        DP_OP_425J2_127_3477_n1862), .Y(DP_OP_425J2_127_3477_n1826) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1052 ( .A1(DP_OP_424J2_126_3477_n2910), .A2(
        DP_OP_425J2_127_3477_n1862), .Y(DP_OP_425J2_127_3477_n1825) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1051 ( .A1(DP_OP_424J2_126_3477_n2909), .A2(
        DP_OP_425J2_127_3477_n1862), .Y(DP_OP_425J2_127_3477_n1824) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1050 ( .A1(DP_OP_425J2_127_3477_n1855), .A2(
        DP_OP_425J2_127_3477_n1862), .Y(DP_OP_425J2_127_3477_n1823) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1049 ( .A1(DP_OP_425J2_127_3477_n1854), 
        .A2(DP_OP_425J2_127_3477_n1862), .Y(DP_OP_425J2_127_3477_n1822) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1001 ( .A1(n297), .A2(
        DP_OP_423J2_125_3477_n2), .Y(DP_OP_425J2_127_3477_n189) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U999 ( .A1(n398), .A2(n341), .Y(
        DP_OP_425J2_127_3477_n181) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U998 ( .A1(n301), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_425J2_127_3477_n179) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U996 ( .A1(n305), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_425J2_127_3477_n175) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U995 ( .A1(n309), .A2(n343), .Y(
        DP_OP_425J2_127_3477_n173) );
  HADDX1_HVT DP_OP_425J2_127_3477_U983 ( .A0(DP_OP_425J2_127_3477_n2117), .B0(
        DP_OP_425J2_127_3477_n2730), .C1(DP_OP_425J2_127_3477_n1771), .SO(
        DP_OP_425J2_127_3477_n1772) );
  FADDX1_HVT DP_OP_425J2_127_3477_U982 ( .A(DP_OP_425J2_127_3477_n2642), .B(
        DP_OP_425J2_127_3477_n1788), .CI(DP_OP_425J2_127_3477_n2293), .CO(
        DP_OP_425J2_127_3477_n1769), .S(DP_OP_425J2_127_3477_n1770) );
  FADDX1_HVT DP_OP_425J2_127_3477_U981 ( .A(DP_OP_425J2_127_3477_n1853), .B(
        DP_OP_425J2_127_3477_n2686), .CI(DP_OP_425J2_127_3477_n2073), .CO(
        DP_OP_425J2_127_3477_n1767), .S(DP_OP_425J2_127_3477_n1768) );
  FADDX1_HVT DP_OP_425J2_127_3477_U980 ( .A(DP_OP_425J2_127_3477_n2205), .B(
        DP_OP_425J2_127_3477_n2029), .CI(DP_OP_425J2_127_3477_n1941), .CO(
        DP_OP_425J2_127_3477_n1765), .S(DP_OP_425J2_127_3477_n1766) );
  FADDX1_HVT DP_OP_425J2_127_3477_U979 ( .A(DP_OP_425J2_127_3477_n2554), .B(
        DP_OP_425J2_127_3477_n1985), .CI(DP_OP_425J2_127_3477_n2510), .CO(
        DP_OP_425J2_127_3477_n1763), .S(DP_OP_425J2_127_3477_n1764) );
  FADDX1_HVT DP_OP_425J2_127_3477_U978 ( .A(DP_OP_425J2_127_3477_n2422), .B(
        DP_OP_425J2_127_3477_n2337), .CI(DP_OP_425J2_127_3477_n1897), .CO(
        DP_OP_425J2_127_3477_n1761), .S(DP_OP_425J2_127_3477_n1762) );
  FADDX1_HVT DP_OP_425J2_127_3477_U977 ( .A(DP_OP_425J2_127_3477_n2598), .B(
        DP_OP_425J2_127_3477_n2466), .CI(DP_OP_425J2_127_3477_n2774), .CO(
        DP_OP_425J2_127_3477_n1759), .S(DP_OP_425J2_127_3477_n1760) );
  FADDX1_HVT DP_OP_425J2_127_3477_U976 ( .A(DP_OP_425J2_127_3477_n2862), .B(
        DP_OP_425J2_127_3477_n2249), .CI(DP_OP_425J2_127_3477_n2906), .CO(
        DP_OP_425J2_127_3477_n1757), .S(DP_OP_425J2_127_3477_n1758) );
  FADDX1_HVT DP_OP_425J2_127_3477_U975 ( .A(DP_OP_425J2_127_3477_n2378), .B(
        DP_OP_425J2_127_3477_n2161), .CI(DP_OP_425J2_127_3477_n2818), .CO(
        DP_OP_425J2_127_3477_n1755), .S(DP_OP_425J2_127_3477_n1756) );
  FADDX1_HVT DP_OP_425J2_127_3477_U974 ( .A(DP_OP_425J2_127_3477_n1772), .B(
        DP_OP_425J2_127_3477_n1762), .CI(DP_OP_425J2_127_3477_n1764), .CO(
        DP_OP_425J2_127_3477_n1753), .S(DP_OP_425J2_127_3477_n1754) );
  FADDX1_HVT DP_OP_425J2_127_3477_U973 ( .A(DP_OP_425J2_127_3477_n1766), .B(
        DP_OP_425J2_127_3477_n1760), .CI(DP_OP_425J2_127_3477_n1758), .CO(
        DP_OP_425J2_127_3477_n1751), .S(DP_OP_425J2_127_3477_n1752) );
  FADDX1_HVT DP_OP_425J2_127_3477_U972 ( .A(DP_OP_425J2_127_3477_n1770), .B(
        DP_OP_425J2_127_3477_n1768), .CI(DP_OP_425J2_127_3477_n1756), .CO(
        DP_OP_425J2_127_3477_n1749), .S(DP_OP_425J2_127_3477_n1750) );
  HADDX1_HVT DP_OP_425J2_127_3477_U971 ( .A0(DP_OP_425J2_127_3477_n2116), .B0(
        DP_OP_425J2_127_3477_n2729), .C1(DP_OP_425J2_127_3477_n1747), .SO(
        DP_OP_425J2_127_3477_n1748) );
  FADDX1_HVT DP_OP_425J2_127_3477_U970 ( .A(DP_OP_425J2_127_3477_n2553), .B(
        DP_OP_425J2_127_3477_n2153), .CI(DP_OP_425J2_127_3477_n2072), .CO(
        DP_OP_425J2_127_3477_n1745), .S(DP_OP_425J2_127_3477_n1746) );
  FADDX1_HVT DP_OP_425J2_127_3477_U969 ( .A(DP_OP_425J2_127_3477_n2597), .B(
        DP_OP_425J2_127_3477_n2414), .CI(DP_OP_425J2_127_3477_n2292), .CO(
        DP_OP_425J2_127_3477_n1743), .S(DP_OP_425J2_127_3477_n1744) );
  FADDX1_HVT DP_OP_425J2_127_3477_U968 ( .A(DP_OP_425J2_127_3477_n2641), .B(
        DP_OP_425J2_127_3477_n1787), .CI(DP_OP_425J2_127_3477_n2285), .CO(
        DP_OP_425J2_127_3477_n1741), .S(DP_OP_425J2_127_3477_n1742) );
  FADDX1_HVT DP_OP_425J2_127_3477_U967 ( .A(DP_OP_425J2_127_3477_n2465), .B(
        DP_OP_425J2_127_3477_n2502), .CI(DP_OP_425J2_127_3477_n2810), .CO(
        DP_OP_425J2_127_3477_n1739), .S(DP_OP_425J2_127_3477_n1740) );
  FADDX1_HVT DP_OP_425J2_127_3477_U966 ( .A(DP_OP_425J2_127_3477_n2336), .B(
        DP_OP_425J2_127_3477_n2065), .CI(DP_OP_425J2_127_3477_n2898), .CO(
        DP_OP_425J2_127_3477_n1737), .S(DP_OP_425J2_127_3477_n1738) );
  FADDX1_HVT DP_OP_425J2_127_3477_U965 ( .A(DP_OP_425J2_127_3477_n2204), .B(
        DP_OP_425J2_127_3477_n2329), .CI(DP_OP_425J2_127_3477_n2854), .CO(
        DP_OP_425J2_127_3477_n1735), .S(DP_OP_425J2_127_3477_n1736) );
  FADDX1_HVT DP_OP_425J2_127_3477_U964 ( .A(DP_OP_425J2_127_3477_n1852), .B(
        DP_OP_425J2_127_3477_n2685), .CI(DP_OP_425J2_127_3477_n2546), .CO(
        DP_OP_425J2_127_3477_n1733), .S(DP_OP_425J2_127_3477_n1734) );
  FADDX1_HVT DP_OP_425J2_127_3477_U963 ( .A(DP_OP_425J2_127_3477_n2421), .B(
        DP_OP_425J2_127_3477_n2028), .CI(DP_OP_425J2_127_3477_n1940), .CO(
        DP_OP_425J2_127_3477_n1731), .S(DP_OP_425J2_127_3477_n1732) );
  FADDX1_HVT DP_OP_425J2_127_3477_U962 ( .A(DP_OP_425J2_127_3477_n1845), .B(
        DP_OP_425J2_127_3477_n1984), .CI(DP_OP_425J2_127_3477_n1896), .CO(
        DP_OP_425J2_127_3477_n1729), .S(DP_OP_425J2_127_3477_n1730) );
  FADDX1_HVT DP_OP_425J2_127_3477_U961 ( .A(DP_OP_425J2_127_3477_n2590), .B(
        DP_OP_425J2_127_3477_n2634), .CI(DP_OP_425J2_127_3477_n2509), .CO(
        DP_OP_425J2_127_3477_n1727), .S(DP_OP_425J2_127_3477_n1728) );
  FADDX1_HVT DP_OP_425J2_127_3477_U960 ( .A(DP_OP_425J2_127_3477_n2861), .B(
        DP_OP_425J2_127_3477_n2773), .CI(DP_OP_425J2_127_3477_n2458), .CO(
        DP_OP_425J2_127_3477_n1725), .S(DP_OP_425J2_127_3477_n1726) );
  FADDX1_HVT DP_OP_425J2_127_3477_U959 ( .A(DP_OP_425J2_127_3477_n2766), .B(
        DP_OP_425J2_127_3477_n1977), .CI(DP_OP_425J2_127_3477_n2370), .CO(
        DP_OP_425J2_127_3477_n1723), .S(DP_OP_425J2_127_3477_n1724) );
  FADDX1_HVT DP_OP_425J2_127_3477_U958 ( .A(DP_OP_425J2_127_3477_n2109), .B(
        DP_OP_425J2_127_3477_n2248), .CI(DP_OP_425J2_127_3477_n2197), .CO(
        DP_OP_425J2_127_3477_n1721), .S(DP_OP_425J2_127_3477_n1722) );
  FADDX1_HVT DP_OP_425J2_127_3477_U957 ( .A(DP_OP_425J2_127_3477_n1889), .B(
        DP_OP_425J2_127_3477_n2678), .CI(DP_OP_425J2_127_3477_n2241), .CO(
        DP_OP_425J2_127_3477_n1719), .S(DP_OP_425J2_127_3477_n1720) );
  FADDX1_HVT DP_OP_425J2_127_3477_U956 ( .A(DP_OP_425J2_127_3477_n2905), .B(
        DP_OP_425J2_127_3477_n1933), .CI(DP_OP_425J2_127_3477_n2817), .CO(
        DP_OP_425J2_127_3477_n1717), .S(DP_OP_425J2_127_3477_n1718) );
  FADDX1_HVT DP_OP_425J2_127_3477_U955 ( .A(DP_OP_425J2_127_3477_n2722), .B(
        DP_OP_425J2_127_3477_n2021), .CI(DP_OP_425J2_127_3477_n2160), .CO(
        DP_OP_425J2_127_3477_n1715), .S(DP_OP_425J2_127_3477_n1716) );
  FADDX1_HVT DP_OP_425J2_127_3477_U954 ( .A(DP_OP_425J2_127_3477_n2377), .B(
        DP_OP_425J2_127_3477_n1771), .CI(DP_OP_425J2_127_3477_n1748), .CO(
        DP_OP_425J2_127_3477_n1713), .S(DP_OP_425J2_127_3477_n1714) );
  FADDX1_HVT DP_OP_425J2_127_3477_U953 ( .A(DP_OP_425J2_127_3477_n1759), .B(
        DP_OP_425J2_127_3477_n1769), .CI(DP_OP_425J2_127_3477_n1757), .CO(
        DP_OP_425J2_127_3477_n1711), .S(DP_OP_425J2_127_3477_n1712) );
  FADDX1_HVT DP_OP_425J2_127_3477_U952 ( .A(DP_OP_425J2_127_3477_n1765), .B(
        DP_OP_425J2_127_3477_n1767), .CI(DP_OP_425J2_127_3477_n1761), .CO(
        DP_OP_425J2_127_3477_n1709), .S(DP_OP_425J2_127_3477_n1710) );
  FADDX1_HVT DP_OP_425J2_127_3477_U951 ( .A(DP_OP_425J2_127_3477_n1763), .B(
        DP_OP_425J2_127_3477_n1755), .CI(DP_OP_425J2_127_3477_n1738), .CO(
        DP_OP_425J2_127_3477_n1707), .S(DP_OP_425J2_127_3477_n1708) );
  FADDX1_HVT DP_OP_425J2_127_3477_U950 ( .A(DP_OP_425J2_127_3477_n1736), .B(
        DP_OP_425J2_127_3477_n1730), .CI(DP_OP_425J2_127_3477_n1726), .CO(
        DP_OP_425J2_127_3477_n1705), .S(DP_OP_425J2_127_3477_n1706) );
  FADDX1_HVT DP_OP_425J2_127_3477_U949 ( .A(DP_OP_425J2_127_3477_n1742), .B(
        DP_OP_425J2_127_3477_n1744), .CI(DP_OP_425J2_127_3477_n1728), .CO(
        DP_OP_425J2_127_3477_n1703), .S(DP_OP_425J2_127_3477_n1704) );
  FADDX1_HVT DP_OP_425J2_127_3477_U948 ( .A(DP_OP_425J2_127_3477_n1740), .B(
        DP_OP_425J2_127_3477_n1746), .CI(DP_OP_425J2_127_3477_n1732), .CO(
        DP_OP_425J2_127_3477_n1701), .S(DP_OP_425J2_127_3477_n1702) );
  FADDX1_HVT DP_OP_425J2_127_3477_U947 ( .A(DP_OP_425J2_127_3477_n1734), .B(
        DP_OP_425J2_127_3477_n1724), .CI(DP_OP_425J2_127_3477_n1722), .CO(
        DP_OP_425J2_127_3477_n1699), .S(DP_OP_425J2_127_3477_n1700) );
  FADDX1_HVT DP_OP_425J2_127_3477_U946 ( .A(DP_OP_425J2_127_3477_n1720), .B(
        DP_OP_425J2_127_3477_n1716), .CI(DP_OP_425J2_127_3477_n1718), .CO(
        DP_OP_425J2_127_3477_n1697), .S(DP_OP_425J2_127_3477_n1698) );
  FADDX1_HVT DP_OP_425J2_127_3477_U945 ( .A(DP_OP_425J2_127_3477_n1714), .B(
        DP_OP_425J2_127_3477_n1753), .CI(DP_OP_425J2_127_3477_n1751), .CO(
        DP_OP_425J2_127_3477_n1695), .S(DP_OP_425J2_127_3477_n1696) );
  FADDX1_HVT DP_OP_425J2_127_3477_U944 ( .A(DP_OP_425J2_127_3477_n1712), .B(
        DP_OP_425J2_127_3477_n1710), .CI(DP_OP_425J2_127_3477_n1749), .CO(
        DP_OP_425J2_127_3477_n1693), .S(DP_OP_425J2_127_3477_n1694) );
  FADDX1_HVT DP_OP_425J2_127_3477_U943 ( .A(DP_OP_425J2_127_3477_n1708), .B(
        DP_OP_425J2_127_3477_n1706), .CI(DP_OP_425J2_127_3477_n1704), .CO(
        DP_OP_425J2_127_3477_n1691), .S(DP_OP_425J2_127_3477_n1692) );
  FADDX1_HVT DP_OP_425J2_127_3477_U942 ( .A(DP_OP_425J2_127_3477_n1702), .B(
        DP_OP_425J2_127_3477_n1700), .CI(DP_OP_425J2_127_3477_n1698), .CO(
        DP_OP_425J2_127_3477_n1689), .S(DP_OP_425J2_127_3477_n1690) );
  FADDX1_HVT DP_OP_425J2_127_3477_U941 ( .A(DP_OP_425J2_127_3477_n1696), .B(
        DP_OP_425J2_127_3477_n1694), .CI(DP_OP_425J2_127_3477_n1692), .CO(
        DP_OP_425J2_127_3477_n1687), .S(DP_OP_425J2_127_3477_n1688) );
  HADDX1_HVT DP_OP_425J2_127_3477_U940 ( .A0(DP_OP_425J2_127_3477_n2115), .B0(
        DP_OP_425J2_127_3477_n2152), .C1(DP_OP_425J2_127_3477_n1685), .SO(
        DP_OP_425J2_127_3477_n1686) );
  FADDX1_HVT DP_OP_425J2_127_3477_U939 ( .A(DP_OP_425J2_127_3477_n2552), .B(
        DP_OP_425J2_127_3477_n2582), .CI(DP_OP_425J2_127_3477_n2145), .CO(
        DP_OP_425J2_127_3477_n1683), .S(DP_OP_425J2_127_3477_n1684) );
  FADDX1_HVT DP_OP_425J2_127_3477_U938 ( .A(DP_OP_425J2_127_3477_n2335), .B(
        DP_OP_425J2_127_3477_n1969), .CI(DP_OP_425J2_127_3477_n2291), .CO(
        DP_OP_425J2_127_3477_n1681), .S(DP_OP_425J2_127_3477_n1682) );
  FADDX1_HVT DP_OP_425J2_127_3477_U937 ( .A(DP_OP_425J2_127_3477_n1851), .B(
        DP_OP_425J2_127_3477_n2538), .CI(DP_OP_425J2_127_3477_n2277), .CO(
        DP_OP_425J2_127_3477_n1679), .S(DP_OP_425J2_127_3477_n1680) );
  FADDX1_HVT DP_OP_425J2_127_3477_U936 ( .A(DP_OP_425J2_127_3477_n2420), .B(
        DP_OP_425J2_127_3477_n2413), .CI(DP_OP_425J2_127_3477_n2071), .CO(
        DP_OP_425J2_127_3477_n1677), .S(DP_OP_425J2_127_3477_n1678) );
  FADDX1_HVT DP_OP_425J2_127_3477_U935 ( .A(DP_OP_425J2_127_3477_n2640), .B(
        DP_OP_425J2_127_3477_n2728), .CI(DP_OP_425J2_127_3477_n2284), .CO(
        DP_OP_425J2_127_3477_n1675), .S(DP_OP_425J2_127_3477_n1676) );
  FADDX1_HVT DP_OP_425J2_127_3477_U934 ( .A(DP_OP_425J2_127_3477_n2464), .B(
        DP_OP_425J2_127_3477_n1786), .CI(DP_OP_425J2_127_3477_n2809), .CO(
        DP_OP_425J2_127_3477_n1673), .S(DP_OP_425J2_127_3477_n1674) );
  FADDX1_HVT DP_OP_425J2_127_3477_U933 ( .A(DP_OP_425J2_127_3477_n2596), .B(
        DP_OP_425J2_127_3477_n2064), .CI(DP_OP_425J2_127_3477_n2057), .CO(
        DP_OP_425J2_127_3477_n1671), .S(DP_OP_425J2_127_3477_n1672) );
  FADDX1_HVT DP_OP_425J2_127_3477_U932 ( .A(DP_OP_425J2_127_3477_n2203), .B(
        DP_OP_425J2_127_3477_n2027), .CI(DP_OP_425J2_127_3477_n2321), .CO(
        DP_OP_425J2_127_3477_n1669), .S(DP_OP_425J2_127_3477_n1670) );
  FADDX1_HVT DP_OP_425J2_127_3477_U931 ( .A(DP_OP_425J2_127_3477_n2890), .B(
        DP_OP_425J2_127_3477_n2684), .CI(DP_OP_425J2_127_3477_n2897), .CO(
        DP_OP_425J2_127_3477_n1667), .S(DP_OP_425J2_127_3477_n1668) );
  FADDX1_HVT DP_OP_425J2_127_3477_U930 ( .A(DP_OP_425J2_127_3477_n2846), .B(
        DP_OP_425J2_127_3477_n2501), .CI(DP_OP_425J2_127_3477_n2853), .CO(
        DP_OP_425J2_127_3477_n1665), .S(DP_OP_425J2_127_3477_n1666) );
  FADDX1_HVT DP_OP_425J2_127_3477_U929 ( .A(DP_OP_425J2_127_3477_n1983), .B(
        DP_OP_425J2_127_3477_n2328), .CI(DP_OP_425J2_127_3477_n2545), .CO(
        DP_OP_425J2_127_3477_n1663), .S(DP_OP_425J2_127_3477_n1664) );
  FADDX1_HVT DP_OP_425J2_127_3477_U928 ( .A(DP_OP_425J2_127_3477_n2589), .B(
        DP_OP_425J2_127_3477_n2758), .CI(DP_OP_425J2_127_3477_n2714), .CO(
        DP_OP_425J2_127_3477_n1661), .S(DP_OP_425J2_127_3477_n1662) );
  FADDX1_HVT DP_OP_425J2_127_3477_U927 ( .A(DP_OP_425J2_127_3477_n1844), .B(
        DP_OP_425J2_127_3477_n2633), .CI(DP_OP_425J2_127_3477_n1939), .CO(
        DP_OP_425J2_127_3477_n1659), .S(DP_OP_425J2_127_3477_n1660) );
  FADDX1_HVT DP_OP_425J2_127_3477_U926 ( .A(DP_OP_425J2_127_3477_n2860), .B(
        DP_OP_425J2_127_3477_n2508), .CI(DP_OP_425J2_127_3477_n2189), .CO(
        DP_OP_425J2_127_3477_n1657), .S(DP_OP_425J2_127_3477_n1658) );
  FADDX1_HVT DP_OP_425J2_127_3477_U925 ( .A(DP_OP_425J2_127_3477_n2772), .B(
        DP_OP_425J2_127_3477_n1895), .CI(DP_OP_425J2_127_3477_n1925), .CO(
        DP_OP_425J2_127_3477_n1655), .S(DP_OP_425J2_127_3477_n1656) );
  FADDX1_HVT DP_OP_425J2_127_3477_U924 ( .A(DP_OP_425J2_127_3477_n2233), .B(
        DP_OP_425J2_127_3477_n2450), .CI(DP_OP_425J2_127_3477_n1881), .CO(
        DP_OP_425J2_127_3477_n1653), .S(DP_OP_425J2_127_3477_n1654) );
  FADDX1_HVT DP_OP_425J2_127_3477_U923 ( .A(DP_OP_425J2_127_3477_n2101), .B(
        DP_OP_425J2_127_3477_n2670), .CI(DP_OP_425J2_127_3477_n2457), .CO(
        DP_OP_425J2_127_3477_n1651), .S(DP_OP_425J2_127_3477_n1652) );
  FADDX1_HVT DP_OP_425J2_127_3477_U922 ( .A(DP_OP_425J2_127_3477_n2765), .B(
        DP_OP_425J2_127_3477_n1837), .CI(DP_OP_425J2_127_3477_n2013), .CO(
        DP_OP_425J2_127_3477_n1649), .S(DP_OP_425J2_127_3477_n1650) );
  FADDX1_HVT DP_OP_425J2_127_3477_U921 ( .A(DP_OP_425J2_127_3477_n1888), .B(
        DP_OP_425J2_127_3477_n2802), .CI(DP_OP_425J2_127_3477_n2240), .CO(
        DP_OP_425J2_127_3477_n1647), .S(DP_OP_425J2_127_3477_n1648) );
  FADDX1_HVT DP_OP_425J2_127_3477_U920 ( .A(DP_OP_425J2_127_3477_n2108), .B(
        DP_OP_425J2_127_3477_n2626), .CI(DP_OP_425J2_127_3477_n2369), .CO(
        DP_OP_425J2_127_3477_n1645), .S(DP_OP_425J2_127_3477_n1646) );
  FADDX1_HVT DP_OP_425J2_127_3477_U919 ( .A(DP_OP_425J2_127_3477_n2494), .B(
        DP_OP_425J2_127_3477_n1976), .CI(DP_OP_425J2_127_3477_n2196), .CO(
        DP_OP_425J2_127_3477_n1643), .S(DP_OP_425J2_127_3477_n1644) );
  FADDX1_HVT DP_OP_425J2_127_3477_U918 ( .A(DP_OP_425J2_127_3477_n2677), .B(
        DP_OP_425J2_127_3477_n2247), .CI(DP_OP_425J2_127_3477_n1932), .CO(
        DP_OP_425J2_127_3477_n1641), .S(DP_OP_425J2_127_3477_n1642) );
  FADDX1_HVT DP_OP_425J2_127_3477_U917 ( .A(DP_OP_425J2_127_3477_n2362), .B(
        DP_OP_425J2_127_3477_n2904), .CI(DP_OP_425J2_127_3477_n2159), .CO(
        DP_OP_425J2_127_3477_n1639), .S(DP_OP_425J2_127_3477_n1640) );
  FADDX1_HVT DP_OP_425J2_127_3477_U916 ( .A(DP_OP_425J2_127_3477_n2376), .B(
        DP_OP_425J2_127_3477_n2406), .CI(DP_OP_425J2_127_3477_n2816), .CO(
        DP_OP_425J2_127_3477_n1637), .S(DP_OP_425J2_127_3477_n1638) );
  FADDX1_HVT DP_OP_425J2_127_3477_U915 ( .A(DP_OP_425J2_127_3477_n2721), .B(
        DP_OP_425J2_127_3477_n2020), .CI(DP_OP_425J2_127_3477_n1747), .CO(
        DP_OP_425J2_127_3477_n1635), .S(DP_OP_425J2_127_3477_n1636) );
  FADDX1_HVT DP_OP_425J2_127_3477_U914 ( .A(DP_OP_425J2_127_3477_n1686), .B(
        DP_OP_425J2_127_3477_n1733), .CI(DP_OP_425J2_127_3477_n1727), .CO(
        DP_OP_425J2_127_3477_n1633), .S(DP_OP_425J2_127_3477_n1634) );
  FADDX1_HVT DP_OP_425J2_127_3477_U913 ( .A(DP_OP_425J2_127_3477_n1745), .B(
        DP_OP_425J2_127_3477_n1729), .CI(DP_OP_425J2_127_3477_n1725), .CO(
        DP_OP_425J2_127_3477_n1631), .S(DP_OP_425J2_127_3477_n1632) );
  FADDX1_HVT DP_OP_425J2_127_3477_U912 ( .A(DP_OP_425J2_127_3477_n1737), .B(
        DP_OP_425J2_127_3477_n1731), .CI(DP_OP_425J2_127_3477_n1735), .CO(
        DP_OP_425J2_127_3477_n1629), .S(DP_OP_425J2_127_3477_n1630) );
  FADDX1_HVT DP_OP_425J2_127_3477_U911 ( .A(DP_OP_425J2_127_3477_n1741), .B(
        DP_OP_425J2_127_3477_n1743), .CI(DP_OP_425J2_127_3477_n1739), .CO(
        DP_OP_425J2_127_3477_n1627), .S(DP_OP_425J2_127_3477_n1628) );
  FADDX1_HVT DP_OP_425J2_127_3477_U910 ( .A(DP_OP_425J2_127_3477_n1723), .B(
        DP_OP_425J2_127_3477_n1719), .CI(DP_OP_425J2_127_3477_n1715), .CO(
        DP_OP_425J2_127_3477_n1625), .S(DP_OP_425J2_127_3477_n1626) );
  FADDX1_HVT DP_OP_425J2_127_3477_U909 ( .A(DP_OP_425J2_127_3477_n1721), .B(
        DP_OP_425J2_127_3477_n1717), .CI(DP_OP_425J2_127_3477_n1668), .CO(
        DP_OP_425J2_127_3477_n1623), .S(DP_OP_425J2_127_3477_n1624) );
  FADDX1_HVT DP_OP_425J2_127_3477_U908 ( .A(DP_OP_425J2_127_3477_n1678), .B(
        DP_OP_425J2_127_3477_n1664), .CI(DP_OP_425J2_127_3477_n1652), .CO(
        DP_OP_425J2_127_3477_n1621), .S(DP_OP_425J2_127_3477_n1622) );
  FADDX1_HVT DP_OP_425J2_127_3477_U907 ( .A(DP_OP_425J2_127_3477_n1676), .B(
        DP_OP_425J2_127_3477_n1662), .CI(DP_OP_425J2_127_3477_n1658), .CO(
        DP_OP_425J2_127_3477_n1619), .S(DP_OP_425J2_127_3477_n1620) );
  FADDX1_HVT DP_OP_425J2_127_3477_U906 ( .A(DP_OP_425J2_127_3477_n1680), .B(
        DP_OP_425J2_127_3477_n1660), .CI(DP_OP_425J2_127_3477_n1654), .CO(
        DP_OP_425J2_127_3477_n1617), .S(DP_OP_425J2_127_3477_n1618) );
  FADDX1_HVT DP_OP_425J2_127_3477_U905 ( .A(DP_OP_425J2_127_3477_n1684), .B(
        DP_OP_425J2_127_3477_n1670), .CI(DP_OP_425J2_127_3477_n1656), .CO(
        DP_OP_425J2_127_3477_n1615), .S(DP_OP_425J2_127_3477_n1616) );
  FADDX1_HVT DP_OP_425J2_127_3477_U904 ( .A(DP_OP_425J2_127_3477_n1672), .B(
        DP_OP_425J2_127_3477_n1682), .CI(DP_OP_425J2_127_3477_n1666), .CO(
        DP_OP_425J2_127_3477_n1613), .S(DP_OP_425J2_127_3477_n1614) );
  FADDX1_HVT DP_OP_425J2_127_3477_U903 ( .A(DP_OP_425J2_127_3477_n1674), .B(
        DP_OP_425J2_127_3477_n1650), .CI(DP_OP_425J2_127_3477_n1646), .CO(
        DP_OP_425J2_127_3477_n1611), .S(DP_OP_425J2_127_3477_n1612) );
  FADDX1_HVT DP_OP_425J2_127_3477_U902 ( .A(DP_OP_425J2_127_3477_n1648), .B(
        DP_OP_425J2_127_3477_n1640), .CI(DP_OP_425J2_127_3477_n1713), .CO(
        DP_OP_425J2_127_3477_n1609), .S(DP_OP_425J2_127_3477_n1610) );
  FADDX1_HVT DP_OP_425J2_127_3477_U901 ( .A(DP_OP_425J2_127_3477_n1644), .B(
        DP_OP_425J2_127_3477_n1642), .CI(DP_OP_425J2_127_3477_n1638), .CO(
        DP_OP_425J2_127_3477_n1607), .S(DP_OP_425J2_127_3477_n1608) );
  FADDX1_HVT DP_OP_425J2_127_3477_U900 ( .A(DP_OP_425J2_127_3477_n1636), .B(
        DP_OP_425J2_127_3477_n1709), .CI(DP_OP_425J2_127_3477_n1711), .CO(
        DP_OP_425J2_127_3477_n1605), .S(DP_OP_425J2_127_3477_n1606) );
  FADDX1_HVT DP_OP_425J2_127_3477_U899 ( .A(DP_OP_425J2_127_3477_n1707), .B(
        DP_OP_425J2_127_3477_n1634), .CI(DP_OP_425J2_127_3477_n1632), .CO(
        DP_OP_425J2_127_3477_n1603), .S(DP_OP_425J2_127_3477_n1604) );
  FADDX1_HVT DP_OP_425J2_127_3477_U898 ( .A(DP_OP_425J2_127_3477_n1630), .B(
        DP_OP_425J2_127_3477_n1705), .CI(DP_OP_425J2_127_3477_n1699), .CO(
        DP_OP_425J2_127_3477_n1601), .S(DP_OP_425J2_127_3477_n1602) );
  FADDX1_HVT DP_OP_425J2_127_3477_U897 ( .A(DP_OP_425J2_127_3477_n1628), .B(
        DP_OP_425J2_127_3477_n1701), .CI(DP_OP_425J2_127_3477_n1703), .CO(
        DP_OP_425J2_127_3477_n1599), .S(DP_OP_425J2_127_3477_n1600) );
  FADDX1_HVT DP_OP_425J2_127_3477_U896 ( .A(DP_OP_425J2_127_3477_n1626), .B(
        DP_OP_425J2_127_3477_n1697), .CI(DP_OP_425J2_127_3477_n1624), .CO(
        DP_OP_425J2_127_3477_n1597), .S(DP_OP_425J2_127_3477_n1598) );
  FADDX1_HVT DP_OP_425J2_127_3477_U895 ( .A(DP_OP_425J2_127_3477_n1622), .B(
        DP_OP_425J2_127_3477_n1614), .CI(DP_OP_425J2_127_3477_n1612), .CO(
        DP_OP_425J2_127_3477_n1595), .S(DP_OP_425J2_127_3477_n1596) );
  FADDX1_HVT DP_OP_425J2_127_3477_U894 ( .A(DP_OP_425J2_127_3477_n1620), .B(
        DP_OP_425J2_127_3477_n1618), .CI(DP_OP_425J2_127_3477_n1616), .CO(
        DP_OP_425J2_127_3477_n1593), .S(DP_OP_425J2_127_3477_n1594) );
  FADDX1_HVT DP_OP_425J2_127_3477_U893 ( .A(DP_OP_425J2_127_3477_n1608), .B(
        DP_OP_425J2_127_3477_n1610), .CI(DP_OP_425J2_127_3477_n1695), .CO(
        DP_OP_425J2_127_3477_n1591), .S(DP_OP_425J2_127_3477_n1592) );
  FADDX1_HVT DP_OP_425J2_127_3477_U892 ( .A(DP_OP_425J2_127_3477_n1606), .B(
        DP_OP_425J2_127_3477_n1693), .CI(DP_OP_425J2_127_3477_n1604), .CO(
        DP_OP_425J2_127_3477_n1589), .S(DP_OP_425J2_127_3477_n1590) );
  FADDX1_HVT DP_OP_425J2_127_3477_U891 ( .A(DP_OP_425J2_127_3477_n1691), .B(
        DP_OP_425J2_127_3477_n1600), .CI(DP_OP_425J2_127_3477_n1689), .CO(
        DP_OP_425J2_127_3477_n1587), .S(DP_OP_425J2_127_3477_n1588) );
  FADDX1_HVT DP_OP_425J2_127_3477_U890 ( .A(DP_OP_425J2_127_3477_n1602), .B(
        DP_OP_425J2_127_3477_n1598), .CI(DP_OP_425J2_127_3477_n1596), .CO(
        DP_OP_425J2_127_3477_n1585), .S(DP_OP_425J2_127_3477_n1586) );
  FADDX1_HVT DP_OP_425J2_127_3477_U889 ( .A(DP_OP_425J2_127_3477_n1594), .B(
        DP_OP_425J2_127_3477_n1592), .CI(DP_OP_425J2_127_3477_n1590), .CO(
        DP_OP_425J2_127_3477_n1583), .S(DP_OP_425J2_127_3477_n1584) );
  FADDX1_HVT DP_OP_425J2_127_3477_U888 ( .A(DP_OP_425J2_127_3477_n1687), .B(
        DP_OP_425J2_127_3477_n1588), .CI(DP_OP_425J2_127_3477_n1586), .CO(
        DP_OP_425J2_127_3477_n1581), .S(DP_OP_425J2_127_3477_n1582) );
  FADDX1_HVT DP_OP_425J2_127_3477_U886 ( .A(DP_OP_425J2_127_3477_n2706), .B(
        DP_OP_425J2_127_3477_n1829), .CI(DP_OP_425J2_127_3477_n2398), .CO(
        DP_OP_425J2_127_3477_n1577), .S(DP_OP_425J2_127_3477_n1578) );
  FADDX1_HVT DP_OP_425J2_127_3477_U885 ( .A(DP_OP_425J2_127_3477_n2005), .B(
        DP_OP_425J2_127_3477_n2181), .CI(DP_OP_425J2_127_3477_n1961), .CO(
        DP_OP_425J2_127_3477_n1575), .S(DP_OP_425J2_127_3477_n1576) );
  FADDX1_HVT DP_OP_425J2_127_3477_U884 ( .A(DP_OP_425J2_127_3477_n2794), .B(
        DP_OP_425J2_127_3477_n2486), .CI(DP_OP_425J2_127_3477_n2750), .CO(
        DP_OP_425J2_127_3477_n1573), .S(DP_OP_425J2_127_3477_n1574) );
  FADDX1_HVT DP_OP_425J2_127_3477_U883 ( .A(DP_OP_425J2_127_3477_n2838), .B(
        DP_OP_425J2_127_3477_n1917), .CI(DP_OP_425J2_127_3477_n2530), .CO(
        DP_OP_425J2_127_3477_n1571), .S(DP_OP_425J2_127_3477_n1572) );
  FADDX1_HVT DP_OP_425J2_127_3477_U882 ( .A(DP_OP_425J2_127_3477_n1873), .B(
        DP_OP_425J2_127_3477_n2442), .CI(DP_OP_425J2_127_3477_n2049), .CO(
        DP_OP_425J2_127_3477_n1569), .S(DP_OP_425J2_127_3477_n1570) );
  FADDX1_HVT DP_OP_425J2_127_3477_U881 ( .A(DP_OP_425J2_127_3477_n2137), .B(
        DP_OP_425J2_127_3477_n2882), .CI(DP_OP_425J2_127_3477_n2574), .CO(
        DP_OP_425J2_127_3477_n1567), .S(DP_OP_425J2_127_3477_n1568) );
  FADDX1_HVT DP_OP_425J2_127_3477_U880 ( .A(DP_OP_425J2_127_3477_n2093), .B(
        DP_OP_425J2_127_3477_n2662), .CI(DP_OP_425J2_127_3477_n2269), .CO(
        DP_OP_425J2_127_3477_n1565), .S(DP_OP_425J2_127_3477_n1566) );
  FADDX1_HVT DP_OP_425J2_127_3477_U879 ( .A(DP_OP_425J2_127_3477_n2618), .B(
        DP_OP_425J2_127_3477_n2313), .CI(DP_OP_425J2_127_3477_n1580), .CO(
        DP_OP_425J2_127_3477_n1563), .S(DP_OP_425J2_127_3477_n1564) );
  FADDX1_HVT DP_OP_425J2_127_3477_U878 ( .A(DP_OP_425J2_127_3477_n2225), .B(
        DP_OP_425J2_127_3477_n2581), .CI(DP_OP_425J2_127_3477_n2283), .CO(
        DP_OP_425J2_127_3477_n1561), .S(DP_OP_425J2_127_3477_n1562) );
  FADDX1_HVT DP_OP_425J2_127_3477_U877 ( .A(DP_OP_425J2_127_3477_n2114), .B(
        DP_OP_425J2_127_3477_n2537), .CI(DP_OP_425J2_127_3477_n2808), .CO(
        DP_OP_425J2_127_3477_n1559), .S(DP_OP_425J2_127_3477_n1560) );
  FADDX1_HVT DP_OP_425J2_127_3477_U876 ( .A(DP_OP_425J2_127_3477_n2551), .B(
        DP_OP_425J2_127_3477_n2412), .CI(DP_OP_425J2_127_3477_n2144), .CO(
        DP_OP_425J2_127_3477_n1557), .S(DP_OP_425J2_127_3477_n1558) );
  FADDX1_HVT DP_OP_425J2_127_3477_U875 ( .A(DP_OP_425J2_127_3477_n2845), .B(
        DP_OP_425J2_127_3477_n1968), .CI(DP_OP_425J2_127_3477_n2070), .CO(
        DP_OP_425J2_127_3477_n1555), .S(DP_OP_425J2_127_3477_n1556) );
  FADDX1_HVT DP_OP_425J2_127_3477_U874 ( .A(DP_OP_425J2_127_3477_n2419), .B(
        DP_OP_425J2_127_3477_n2727), .CI(DP_OP_425J2_127_3477_n2276), .CO(
        DP_OP_425J2_127_3477_n1553), .S(DP_OP_425J2_127_3477_n1554) );
  FADDX1_HVT DP_OP_425J2_127_3477_U873 ( .A(DP_OP_425J2_127_3477_n2595), .B(
        DP_OP_425J2_127_3477_n2151), .CI(DP_OP_425J2_127_3477_n2290), .CO(
        DP_OP_425J2_127_3477_n1551), .S(DP_OP_425J2_127_3477_n1552) );
  FADDX1_HVT DP_OP_425J2_127_3477_U872 ( .A(DP_OP_425J2_127_3477_n1850), .B(
        DP_OP_425J2_127_3477_n1785), .CI(DP_OP_425J2_127_3477_n2056), .CO(
        DP_OP_425J2_127_3477_n1549), .S(DP_OP_425J2_127_3477_n1550) );
  FADDX1_HVT DP_OP_425J2_127_3477_U871 ( .A(DP_OP_425J2_127_3477_n2639), .B(
        DP_OP_425J2_127_3477_n2632), .CI(DP_OP_425J2_127_3477_n2320), .CO(
        DP_OP_425J2_127_3477_n1547), .S(DP_OP_425J2_127_3477_n1548) );
  FADDX1_HVT DP_OP_425J2_127_3477_U870 ( .A(DP_OP_425J2_127_3477_n2463), .B(
        DP_OP_425J2_127_3477_n2063), .CI(DP_OP_425J2_127_3477_n2896), .CO(
        DP_OP_425J2_127_3477_n1545), .S(DP_OP_425J2_127_3477_n1546) );
  FADDX1_HVT DP_OP_425J2_127_3477_U869 ( .A(DP_OP_425J2_127_3477_n2334), .B(
        DP_OP_425J2_127_3477_n2500), .CI(DP_OP_425J2_127_3477_n2852), .CO(
        DP_OP_425J2_127_3477_n1543), .S(DP_OP_425J2_127_3477_n1544) );
  FADDX1_HVT DP_OP_425J2_127_3477_U868 ( .A(DP_OP_425J2_127_3477_n2202), .B(
        DP_OP_425J2_127_3477_n2757), .CI(DP_OP_425J2_127_3477_n2544), .CO(
        DP_OP_425J2_127_3477_n1541), .S(DP_OP_425J2_127_3477_n1542) );
  FADDX1_HVT DP_OP_425J2_127_3477_U867 ( .A(DP_OP_425J2_127_3477_n2889), .B(
        DP_OP_425J2_127_3477_n1843), .CI(DP_OP_425J2_127_3477_n2713), .CO(
        DP_OP_425J2_127_3477_n1539), .S(DP_OP_425J2_127_3477_n1540) );
  FADDX1_HVT DP_OP_425J2_127_3477_U866 ( .A(DP_OP_425J2_127_3477_n2588), .B(
        DP_OP_425J2_127_3477_n2026), .CI(DP_OP_425J2_127_3477_n1938), .CO(
        DP_OP_425J2_127_3477_n1537), .S(DP_OP_425J2_127_3477_n1538) );
  FADDX1_HVT DP_OP_425J2_127_3477_U865 ( .A(DP_OP_425J2_127_3477_n1982), .B(
        DP_OP_425J2_127_3477_n2327), .CI(DP_OP_425J2_127_3477_n2507), .CO(
        DP_OP_425J2_127_3477_n1535), .S(DP_OP_425J2_127_3477_n1536) );
  FADDX1_HVT DP_OP_425J2_127_3477_U864 ( .A(DP_OP_425J2_127_3477_n2683), .B(
        DP_OP_425J2_127_3477_n2100), .CI(DP_OP_425J2_127_3477_n1894), .CO(
        DP_OP_425J2_127_3477_n1533), .S(DP_OP_425J2_127_3477_n1534) );
  FADDX1_HVT DP_OP_425J2_127_3477_U863 ( .A(DP_OP_425J2_127_3477_n2771), .B(
        DP_OP_425J2_127_3477_n2449), .CI(DP_OP_425J2_127_3477_n2188), .CO(
        DP_OP_425J2_127_3477_n1531), .S(DP_OP_425J2_127_3477_n1532) );
  FADDX1_HVT DP_OP_425J2_127_3477_U862 ( .A(DP_OP_425J2_127_3477_n2232), .B(
        DP_OP_425J2_127_3477_n2859), .CI(DP_OP_425J2_127_3477_n1924), .CO(
        DP_OP_425J2_127_3477_n1529), .S(DP_OP_425J2_127_3477_n1530) );
  FADDX1_HVT DP_OP_425J2_127_3477_U861 ( .A(DP_OP_425J2_127_3477_n2669), .B(
        DP_OP_425J2_127_3477_n1836), .CI(DP_OP_425J2_127_3477_n1931), .CO(
        DP_OP_425J2_127_3477_n1527), .S(DP_OP_425J2_127_3477_n1528) );
  FADDX1_HVT DP_OP_425J2_127_3477_U860 ( .A(DP_OP_425J2_127_3477_n2764), .B(
        DP_OP_425J2_127_3477_n1880), .CI(DP_OP_425J2_127_3477_n2368), .CO(
        DP_OP_425J2_127_3477_n1525), .S(DP_OP_425J2_127_3477_n1526) );
  FADDX1_HVT DP_OP_425J2_127_3477_U859 ( .A(DP_OP_425J2_127_3477_n2107), .B(
        DP_OP_425J2_127_3477_n2456), .CI(DP_OP_425J2_127_3477_n2239), .CO(
        DP_OP_425J2_127_3477_n1523), .S(DP_OP_425J2_127_3477_n1524) );
  FADDX1_HVT DP_OP_425J2_127_3477_U858 ( .A(DP_OP_425J2_127_3477_n1887), .B(
        DP_OP_425J2_127_3477_n2625), .CI(DP_OP_425J2_127_3477_n2195), .CO(
        DP_OP_425J2_127_3477_n1521), .S(DP_OP_425J2_127_3477_n1522) );
  FADDX1_HVT DP_OP_425J2_127_3477_U857 ( .A(DP_OP_425J2_127_3477_n2493), .B(
        DP_OP_425J2_127_3477_n2801), .CI(DP_OP_425J2_127_3477_n2012), .CO(
        DP_OP_425J2_127_3477_n1519), .S(DP_OP_425J2_127_3477_n1520) );
  FADDX1_HVT DP_OP_425J2_127_3477_U856 ( .A(DP_OP_425J2_127_3477_n2676), .B(
        DP_OP_425J2_127_3477_n1975), .CI(DP_OP_425J2_127_3477_n2158), .CO(
        DP_OP_425J2_127_3477_n1517), .S(DP_OP_425J2_127_3477_n1518) );
  FADDX1_HVT DP_OP_425J2_127_3477_U855 ( .A(DP_OP_425J2_127_3477_n2361), .B(
        DP_OP_425J2_127_3477_n2246), .CI(DP_OP_425J2_127_3477_n2405), .CO(
        DP_OP_425J2_127_3477_n1515), .S(DP_OP_425J2_127_3477_n1516) );
  FADDX1_HVT DP_OP_425J2_127_3477_U854 ( .A(DP_OP_425J2_127_3477_n2903), .B(
        DP_OP_425J2_127_3477_n2019), .CI(DP_OP_425J2_127_3477_n2815), .CO(
        DP_OP_425J2_127_3477_n1513), .S(DP_OP_425J2_127_3477_n1514) );
  FADDX1_HVT DP_OP_425J2_127_3477_U853 ( .A(DP_OP_425J2_127_3477_n2720), .B(
        DP_OP_425J2_127_3477_n2375), .CI(DP_OP_425J2_127_3477_n1685), .CO(
        DP_OP_425J2_127_3477_n1511), .S(DP_OP_425J2_127_3477_n1512) );
  FADDX1_HVT DP_OP_425J2_127_3477_U852 ( .A(DP_OP_425J2_127_3477_n1683), .B(
        DP_OP_425J2_127_3477_n1659), .CI(DP_OP_425J2_127_3477_n1651), .CO(
        DP_OP_425J2_127_3477_n1509), .S(DP_OP_425J2_127_3477_n1510) );
  FADDX1_HVT DP_OP_425J2_127_3477_U851 ( .A(DP_OP_425J2_127_3477_n1681), .B(
        DP_OP_425J2_127_3477_n1661), .CI(DP_OP_425J2_127_3477_n1653), .CO(
        DP_OP_425J2_127_3477_n1507), .S(DP_OP_425J2_127_3477_n1508) );
  FADDX1_HVT DP_OP_425J2_127_3477_U850 ( .A(DP_OP_425J2_127_3477_n1679), .B(
        DP_OP_425J2_127_3477_n1663), .CI(DP_OP_425J2_127_3477_n1655), .CO(
        DP_OP_425J2_127_3477_n1505), .S(DP_OP_425J2_127_3477_n1506) );
  FADDX1_HVT DP_OP_425J2_127_3477_U849 ( .A(DP_OP_425J2_127_3477_n1677), .B(
        DP_OP_425J2_127_3477_n1675), .CI(DP_OP_425J2_127_3477_n1657), .CO(
        DP_OP_425J2_127_3477_n1503), .S(DP_OP_425J2_127_3477_n1504) );
  FADDX1_HVT DP_OP_425J2_127_3477_U848 ( .A(DP_OP_425J2_127_3477_n1673), .B(
        DP_OP_425J2_127_3477_n1665), .CI(DP_OP_425J2_127_3477_n1667), .CO(
        DP_OP_425J2_127_3477_n1501), .S(DP_OP_425J2_127_3477_n1502) );
  FADDX1_HVT DP_OP_425J2_127_3477_U847 ( .A(DP_OP_425J2_127_3477_n1671), .B(
        DP_OP_425J2_127_3477_n1669), .CI(DP_OP_425J2_127_3477_n1649), .CO(
        DP_OP_425J2_127_3477_n1499), .S(DP_OP_425J2_127_3477_n1500) );
  FADDX1_HVT DP_OP_425J2_127_3477_U846 ( .A(DP_OP_425J2_127_3477_n1647), .B(
        DP_OP_425J2_127_3477_n1568), .CI(DP_OP_425J2_127_3477_n1637), .CO(
        DP_OP_425J2_127_3477_n1497), .S(DP_OP_425J2_127_3477_n1498) );
  FADDX1_HVT DP_OP_425J2_127_3477_U845 ( .A(DP_OP_425J2_127_3477_n1645), .B(
        DP_OP_425J2_127_3477_n1572), .CI(DP_OP_425J2_127_3477_n1564), .CO(
        DP_OP_425J2_127_3477_n1495), .S(DP_OP_425J2_127_3477_n1496) );
  FADDX1_HVT DP_OP_425J2_127_3477_U844 ( .A(DP_OP_425J2_127_3477_n1643), .B(
        DP_OP_425J2_127_3477_n1570), .CI(DP_OP_425J2_127_3477_n1574), .CO(
        DP_OP_425J2_127_3477_n1493), .S(DP_OP_425J2_127_3477_n1494) );
  FADDX1_HVT DP_OP_425J2_127_3477_U843 ( .A(DP_OP_425J2_127_3477_n1641), .B(
        DP_OP_425J2_127_3477_n1578), .CI(DP_OP_425J2_127_3477_n1566), .CO(
        DP_OP_425J2_127_3477_n1491), .S(DP_OP_425J2_127_3477_n1492) );
  FADDX1_HVT DP_OP_425J2_127_3477_U842 ( .A(DP_OP_425J2_127_3477_n1639), .B(
        DP_OP_425J2_127_3477_n1576), .CI(DP_OP_425J2_127_3477_n1635), .CO(
        DP_OP_425J2_127_3477_n1489), .S(DP_OP_425J2_127_3477_n1490) );
  FADDX1_HVT DP_OP_425J2_127_3477_U841 ( .A(DP_OP_425J2_127_3477_n1562), .B(
        DP_OP_425J2_127_3477_n1534), .CI(DP_OP_425J2_127_3477_n1530), .CO(
        DP_OP_425J2_127_3477_n1487), .S(DP_OP_425J2_127_3477_n1488) );
  FADDX1_HVT DP_OP_425J2_127_3477_U840 ( .A(DP_OP_425J2_127_3477_n1560), .B(
        DP_OP_425J2_127_3477_n1538), .CI(DP_OP_425J2_127_3477_n1532), .CO(
        DP_OP_425J2_127_3477_n1485), .S(DP_OP_425J2_127_3477_n1486) );
  FADDX1_HVT DP_OP_425J2_127_3477_U839 ( .A(DP_OP_425J2_127_3477_n1552), .B(
        DP_OP_425J2_127_3477_n1542), .CI(DP_OP_425J2_127_3477_n1536), .CO(
        DP_OP_425J2_127_3477_n1483), .S(DP_OP_425J2_127_3477_n1484) );
  FADDX1_HVT DP_OP_425J2_127_3477_U838 ( .A(DP_OP_425J2_127_3477_n1554), .B(
        DP_OP_425J2_127_3477_n1540), .CI(DP_OP_425J2_127_3477_n1548), .CO(
        DP_OP_425J2_127_3477_n1481), .S(DP_OP_425J2_127_3477_n1482) );
  FADDX1_HVT DP_OP_425J2_127_3477_U837 ( .A(DP_OP_425J2_127_3477_n1546), .B(
        DP_OP_425J2_127_3477_n1544), .CI(DP_OP_425J2_127_3477_n1550), .CO(
        DP_OP_425J2_127_3477_n1479), .S(DP_OP_425J2_127_3477_n1480) );
  FADDX1_HVT DP_OP_425J2_127_3477_U836 ( .A(DP_OP_425J2_127_3477_n1556), .B(
        DP_OP_425J2_127_3477_n1558), .CI(DP_OP_425J2_127_3477_n1528), .CO(
        DP_OP_425J2_127_3477_n1477), .S(DP_OP_425J2_127_3477_n1478) );
  FADDX1_HVT DP_OP_425J2_127_3477_U835 ( .A(DP_OP_425J2_127_3477_n1526), .B(
        DP_OP_425J2_127_3477_n1516), .CI(DP_OP_425J2_127_3477_n1514), .CO(
        DP_OP_425J2_127_3477_n1475), .S(DP_OP_425J2_127_3477_n1476) );
  FADDX1_HVT DP_OP_425J2_127_3477_U834 ( .A(DP_OP_425J2_127_3477_n1522), .B(
        DP_OP_425J2_127_3477_n1524), .CI(DP_OP_425J2_127_3477_n1518), .CO(
        DP_OP_425J2_127_3477_n1473), .S(DP_OP_425J2_127_3477_n1474) );
  FADDX1_HVT DP_OP_425J2_127_3477_U833 ( .A(DP_OP_425J2_127_3477_n1520), .B(
        DP_OP_425J2_127_3477_n1512), .CI(DP_OP_425J2_127_3477_n1633), .CO(
        DP_OP_425J2_127_3477_n1471), .S(DP_OP_425J2_127_3477_n1472) );
  FADDX1_HVT DP_OP_425J2_127_3477_U832 ( .A(DP_OP_425J2_127_3477_n1631), .B(
        DP_OP_425J2_127_3477_n1627), .CI(DP_OP_425J2_127_3477_n1629), .CO(
        DP_OP_425J2_127_3477_n1469), .S(DP_OP_425J2_127_3477_n1470) );
  FADDX1_HVT DP_OP_425J2_127_3477_U831 ( .A(DP_OP_425J2_127_3477_n1625), .B(
        DP_OP_425J2_127_3477_n1623), .CI(DP_OP_425J2_127_3477_n1621), .CO(
        DP_OP_425J2_127_3477_n1467), .S(DP_OP_425J2_127_3477_n1468) );
  FADDX1_HVT DP_OP_425J2_127_3477_U830 ( .A(DP_OP_425J2_127_3477_n1619), .B(
        DP_OP_425J2_127_3477_n1500), .CI(DP_OP_425J2_127_3477_n1611), .CO(
        DP_OP_425J2_127_3477_n1465), .S(DP_OP_425J2_127_3477_n1466) );
  FADDX1_HVT DP_OP_425J2_127_3477_U829 ( .A(DP_OP_425J2_127_3477_n1510), .B(
        DP_OP_425J2_127_3477_n1504), .CI(DP_OP_425J2_127_3477_n1508), .CO(
        DP_OP_425J2_127_3477_n1463), .S(DP_OP_425J2_127_3477_n1464) );
  FADDX1_HVT DP_OP_425J2_127_3477_U828 ( .A(DP_OP_425J2_127_3477_n1617), .B(
        DP_OP_425J2_127_3477_n1615), .CI(DP_OP_425J2_127_3477_n1506), .CO(
        DP_OP_425J2_127_3477_n1461), .S(DP_OP_425J2_127_3477_n1462) );
  FADDX1_HVT DP_OP_425J2_127_3477_U827 ( .A(DP_OP_425J2_127_3477_n1502), .B(
        DP_OP_425J2_127_3477_n1613), .CI(DP_OP_425J2_127_3477_n1496), .CO(
        DP_OP_425J2_127_3477_n1459), .S(DP_OP_425J2_127_3477_n1460) );
  FADDX1_HVT DP_OP_425J2_127_3477_U826 ( .A(DP_OP_425J2_127_3477_n1607), .B(
        DP_OP_425J2_127_3477_n1492), .CI(DP_OP_425J2_127_3477_n1490), .CO(
        DP_OP_425J2_127_3477_n1457), .S(DP_OP_425J2_127_3477_n1458) );
  FADDX1_HVT DP_OP_425J2_127_3477_U825 ( .A(DP_OP_425J2_127_3477_n1494), .B(
        DP_OP_425J2_127_3477_n1609), .CI(DP_OP_425J2_127_3477_n1498), .CO(
        DP_OP_425J2_127_3477_n1455), .S(DP_OP_425J2_127_3477_n1456) );
  FADDX1_HVT DP_OP_425J2_127_3477_U824 ( .A(DP_OP_425J2_127_3477_n1488), .B(
        DP_OP_425J2_127_3477_n1478), .CI(DP_OP_425J2_127_3477_n1605), .CO(
        DP_OP_425J2_127_3477_n1453), .S(DP_OP_425J2_127_3477_n1454) );
  FADDX1_HVT DP_OP_425J2_127_3477_U823 ( .A(DP_OP_425J2_127_3477_n1486), .B(
        DP_OP_425J2_127_3477_n1480), .CI(DP_OP_425J2_127_3477_n1482), .CO(
        DP_OP_425J2_127_3477_n1451), .S(DP_OP_425J2_127_3477_n1452) );
  FADDX1_HVT DP_OP_425J2_127_3477_U822 ( .A(DP_OP_425J2_127_3477_n1484), .B(
        DP_OP_425J2_127_3477_n1476), .CI(DP_OP_425J2_127_3477_n1474), .CO(
        DP_OP_425J2_127_3477_n1449), .S(DP_OP_425J2_127_3477_n1450) );
  FADDX1_HVT DP_OP_425J2_127_3477_U821 ( .A(DP_OP_425J2_127_3477_n1472), .B(
        DP_OP_425J2_127_3477_n1603), .CI(DP_OP_425J2_127_3477_n1599), .CO(
        DP_OP_425J2_127_3477_n1447), .S(DP_OP_425J2_127_3477_n1448) );
  FADDX1_HVT DP_OP_425J2_127_3477_U820 ( .A(DP_OP_425J2_127_3477_n1601), .B(
        DP_OP_425J2_127_3477_n1470), .CI(DP_OP_425J2_127_3477_n1597), .CO(
        DP_OP_425J2_127_3477_n1445), .S(DP_OP_425J2_127_3477_n1446) );
  FADDX1_HVT DP_OP_425J2_127_3477_U819 ( .A(DP_OP_425J2_127_3477_n1468), .B(
        DP_OP_425J2_127_3477_n1593), .CI(DP_OP_425J2_127_3477_n1595), .CO(
        DP_OP_425J2_127_3477_n1443), .S(DP_OP_425J2_127_3477_n1444) );
  FADDX1_HVT DP_OP_425J2_127_3477_U818 ( .A(DP_OP_425J2_127_3477_n1464), .B(
        DP_OP_425J2_127_3477_n1462), .CI(DP_OP_425J2_127_3477_n1460), .CO(
        DP_OP_425J2_127_3477_n1441), .S(DP_OP_425J2_127_3477_n1442) );
  FADDX1_HVT DP_OP_425J2_127_3477_U817 ( .A(DP_OP_425J2_127_3477_n1466), .B(
        DP_OP_425J2_127_3477_n1456), .CI(DP_OP_425J2_127_3477_n1458), .CO(
        DP_OP_425J2_127_3477_n1439), .S(DP_OP_425J2_127_3477_n1440) );
  FADDX1_HVT DP_OP_425J2_127_3477_U816 ( .A(DP_OP_425J2_127_3477_n1591), .B(
        DP_OP_425J2_127_3477_n1454), .CI(DP_OP_425J2_127_3477_n1452), .CO(
        DP_OP_425J2_127_3477_n1437), .S(DP_OP_425J2_127_3477_n1438) );
  FADDX1_HVT DP_OP_425J2_127_3477_U815 ( .A(DP_OP_425J2_127_3477_n1450), .B(
        DP_OP_425J2_127_3477_n1589), .CI(DP_OP_425J2_127_3477_n1448), .CO(
        DP_OP_425J2_127_3477_n1435), .S(DP_OP_425J2_127_3477_n1436) );
  FADDX1_HVT DP_OP_425J2_127_3477_U814 ( .A(DP_OP_425J2_127_3477_n1587), .B(
        DP_OP_425J2_127_3477_n1446), .CI(DP_OP_425J2_127_3477_n1585), .CO(
        DP_OP_425J2_127_3477_n1433), .S(DP_OP_425J2_127_3477_n1434) );
  FADDX1_HVT DP_OP_425J2_127_3477_U813 ( .A(DP_OP_425J2_127_3477_n1444), .B(
        DP_OP_425J2_127_3477_n1442), .CI(DP_OP_425J2_127_3477_n1440), .CO(
        DP_OP_425J2_127_3477_n1431), .S(DP_OP_425J2_127_3477_n1432) );
  FADDX1_HVT DP_OP_425J2_127_3477_U812 ( .A(DP_OP_425J2_127_3477_n1438), .B(
        DP_OP_425J2_127_3477_n1583), .CI(DP_OP_425J2_127_3477_n1436), .CO(
        DP_OP_425J2_127_3477_n1429), .S(DP_OP_425J2_127_3477_n1430) );
  FADDX1_HVT DP_OP_425J2_127_3477_U811 ( .A(DP_OP_425J2_127_3477_n1581), .B(
        DP_OP_425J2_127_3477_n1434), .CI(DP_OP_425J2_127_3477_n1432), .CO(
        DP_OP_425J2_127_3477_n1427), .S(DP_OP_425J2_127_3477_n1428) );
  FADDX1_HVT DP_OP_425J2_127_3477_U810 ( .A(DP_OP_425J2_127_3477_n1579), .B(
        DP_OP_425J2_127_3477_n1828), .CI(DP_OP_425J2_127_3477_n2397), .CO(
        DP_OP_425J2_127_3477_n1425), .S(DP_OP_425J2_127_3477_n1426) );
  FADDX1_HVT DP_OP_425J2_127_3477_U809 ( .A(DP_OP_425J2_127_3477_n2354), .B(
        DP_OP_425J2_127_3477_n1916), .CI(DP_OP_425J2_127_3477_n1960), .CO(
        DP_OP_425J2_127_3477_n1423), .S(DP_OP_425J2_127_3477_n1424) );
  FADDX1_HVT DP_OP_425J2_127_3477_U808 ( .A(DP_OP_425J2_127_3477_n2705), .B(
        DP_OP_425J2_127_3477_n2048), .CI(DP_OP_425J2_127_3477_n2749), .CO(
        DP_OP_425J2_127_3477_n1421), .S(DP_OP_425J2_127_3477_n1422) );
  FADDX1_HVT DP_OP_425J2_127_3477_U807 ( .A(DP_OP_425J2_127_3477_n2004), .B(
        DP_OP_425J2_127_3477_n2485), .CI(DP_OP_425J2_127_3477_n2180), .CO(
        DP_OP_425J2_127_3477_n1419), .S(DP_OP_425J2_127_3477_n1420) );
  FADDX1_HVT DP_OP_425J2_127_3477_U806 ( .A(DP_OP_425J2_127_3477_n2793), .B(
        DP_OP_425J2_127_3477_n2573), .CI(DP_OP_425J2_127_3477_n2529), .CO(
        DP_OP_425J2_127_3477_n1417), .S(DP_OP_425J2_127_3477_n1418) );
  FADDX1_HVT DP_OP_425J2_127_3477_U805 ( .A(DP_OP_425J2_127_3477_n2092), .B(
        DP_OP_425J2_127_3477_n2881), .CI(DP_OP_425J2_127_3477_n2441), .CO(
        DP_OP_425J2_127_3477_n1415), .S(DP_OP_425J2_127_3477_n1416) );
  FADDX1_HVT DP_OP_425J2_127_3477_U804 ( .A(DP_OP_425J2_127_3477_n2136), .B(
        DP_OP_425J2_127_3477_n2837), .CI(DP_OP_425J2_127_3477_n2268), .CO(
        DP_OP_425J2_127_3477_n1413), .S(DP_OP_425J2_127_3477_n1414) );
  FADDX1_HVT DP_OP_425J2_127_3477_U803 ( .A(DP_OP_425J2_127_3477_n2617), .B(
        DP_OP_425J2_127_3477_n1872), .CI(DP_OP_425J2_127_3477_n2661), .CO(
        DP_OP_425J2_127_3477_n1411), .S(DP_OP_425J2_127_3477_n1412) );
  FADDX1_HVT DP_OP_425J2_127_3477_U802 ( .A(DP_OP_425J2_127_3477_n2312), .B(
        DP_OP_425J2_127_3477_n2224), .CI(DP_OP_425J2_127_3477_n2113), .CO(
        DP_OP_425J2_127_3477_n1409), .S(DP_OP_425J2_127_3477_n1410) );
  FADDX1_HVT DP_OP_425J2_127_3477_U801 ( .A(DP_OP_425J2_127_3477_n2462), .B(
        DP_OP_425J2_127_3477_n2580), .CI(DP_OP_425J2_127_3477_n2275), .CO(
        DP_OP_425J2_127_3477_n1407), .S(DP_OP_425J2_127_3477_n1408) );
  FADDX1_HVT DP_OP_425J2_127_3477_U800 ( .A(DP_OP_425J2_127_3477_n1849), .B(
        DP_OP_425J2_127_3477_n2536), .CI(DP_OP_425J2_127_3477_n2143), .CO(
        DP_OP_425J2_127_3477_n1405), .S(DP_OP_425J2_127_3477_n1406) );
  FADDX1_HVT DP_OP_425J2_127_3477_U799 ( .A(DP_OP_425J2_127_3477_n2418), .B(
        DP_OP_425J2_127_3477_n2150), .CI(DP_OP_425J2_127_3477_n2289), .CO(
        DP_OP_425J2_127_3477_n1403), .S(DP_OP_425J2_127_3477_n1404) );
  FADDX1_HVT DP_OP_425J2_127_3477_U798 ( .A(DP_OP_425J2_127_3477_n2550), .B(
        DP_OP_425J2_127_3477_n2726), .CI(DP_OP_425J2_127_3477_n2069), .CO(
        DP_OP_425J2_127_3477_n1401), .S(DP_OP_425J2_127_3477_n1402) );
  FADDX1_HVT DP_OP_425J2_127_3477_U797 ( .A(DP_OP_425J2_127_3477_n2888), .B(
        DP_OP_425J2_127_3477_n2411), .CI(DP_OP_425J2_127_3477_n2807), .CO(
        DP_OP_425J2_127_3477_n1399), .S(DP_OP_425J2_127_3477_n1400) );
  FADDX1_HVT DP_OP_425J2_127_3477_U796 ( .A(DP_OP_425J2_127_3477_n2638), .B(
        DP_OP_425J2_127_3477_n1967), .CI(DP_OP_425J2_127_3477_n2282), .CO(
        DP_OP_425J2_127_3477_n1397), .S(DP_OP_425J2_127_3477_n1398) );
  FADDX1_HVT DP_OP_425J2_127_3477_U795 ( .A(DP_OP_425J2_127_3477_n2844), .B(
        DP_OP_425J2_127_3477_n1784), .CI(DP_OP_425J2_127_3477_n2319), .CO(
        DP_OP_425J2_127_3477_n1395), .S(DP_OP_425J2_127_3477_n1396) );
  FADDX1_HVT DP_OP_425J2_127_3477_U794 ( .A(DP_OP_425J2_127_3477_n2333), .B(
        DP_OP_425J2_127_3477_n2062), .CI(DP_OP_425J2_127_3477_n2055), .CO(
        DP_OP_425J2_127_3477_n1393), .S(DP_OP_425J2_127_3477_n1394) );
  FADDX1_HVT DP_OP_425J2_127_3477_U793 ( .A(DP_OP_425J2_127_3477_n2201), .B(
        DP_OP_425J2_127_3477_n2499), .CI(DP_OP_425J2_127_3477_n2895), .CO(
        DP_OP_425J2_127_3477_n1391), .S(DP_OP_425J2_127_3477_n1392) );
  FADDX1_HVT DP_OP_425J2_127_3477_U792 ( .A(DP_OP_425J2_127_3477_n2594), .B(
        DP_OP_425J2_127_3477_n2631), .CI(DP_OP_425J2_127_3477_n2851), .CO(
        DP_OP_425J2_127_3477_n1389), .S(DP_OP_425J2_127_3477_n1390) );
  FADDX1_HVT DP_OP_425J2_127_3477_U791 ( .A(DP_OP_425J2_127_3477_n2756), .B(
        DP_OP_425J2_127_3477_n2587), .CI(DP_OP_425J2_127_3477_n2543), .CO(
        DP_OP_425J2_127_3477_n1387), .S(DP_OP_425J2_127_3477_n1388) );
  FADDX1_HVT DP_OP_425J2_127_3477_U790 ( .A(DP_OP_425J2_127_3477_n2326), .B(
        DP_OP_425J2_127_3477_n2025), .CI(DP_OP_425J2_127_3477_n2712), .CO(
        DP_OP_425J2_127_3477_n1385), .S(DP_OP_425J2_127_3477_n1386) );
  FADDX1_HVT DP_OP_425J2_127_3477_U789 ( .A(DP_OP_425J2_127_3477_n2682), .B(
        DP_OP_425J2_127_3477_n1842), .CI(DP_OP_425J2_127_3477_n1937), .CO(
        DP_OP_425J2_127_3477_n1383), .S(DP_OP_425J2_127_3477_n1384) );
  FADDX1_HVT DP_OP_425J2_127_3477_U788 ( .A(DP_OP_425J2_127_3477_n1981), .B(
        DP_OP_425J2_127_3477_n2231), .CI(DP_OP_425J2_127_3477_n2448), .CO(
        DP_OP_425J2_127_3477_n1381), .S(DP_OP_425J2_127_3477_n1382) );
  FADDX1_HVT DP_OP_425J2_127_3477_U787 ( .A(DP_OP_425J2_127_3477_n2099), .B(
        DP_OP_425J2_127_3477_n1893), .CI(DP_OP_425J2_127_3477_n1923), .CO(
        DP_OP_425J2_127_3477_n1379), .S(DP_OP_425J2_127_3477_n1380) );
  FADDX1_HVT DP_OP_425J2_127_3477_U786 ( .A(DP_OP_425J2_127_3477_n2858), .B(
        DP_OP_425J2_127_3477_n2506), .CI(DP_OP_425J2_127_3477_n2187), .CO(
        DP_OP_425J2_127_3477_n1377), .S(DP_OP_425J2_127_3477_n1378) );
  FADDX1_HVT DP_OP_425J2_127_3477_U785 ( .A(DP_OP_425J2_127_3477_n2770), .B(
        DP_OP_425J2_127_3477_n2668), .CI(DP_OP_425J2_127_3477_n1879), .CO(
        DP_OP_425J2_127_3477_n1375), .S(DP_OP_425J2_127_3477_n1376) );
  FADDX1_HVT DP_OP_425J2_127_3477_U784 ( .A(DP_OP_425J2_127_3477_n2763), .B(
        DP_OP_425J2_127_3477_n2455), .CI(DP_OP_425J2_127_3477_n2011), .CO(
        DP_OP_425J2_127_3477_n1373), .S(DP_OP_425J2_127_3477_n1374) );
  FADDX1_HVT DP_OP_425J2_127_3477_U783 ( .A(DP_OP_425J2_127_3477_n1886), .B(
        DP_OP_425J2_127_3477_n1835), .CI(DP_OP_425J2_127_3477_n2367), .CO(
        DP_OP_425J2_127_3477_n1371), .S(DP_OP_425J2_127_3477_n1372) );
  FADDX1_HVT DP_OP_425J2_127_3477_U782 ( .A(DP_OP_425J2_127_3477_n2492), .B(
        DP_OP_425J2_127_3477_n2800), .CI(DP_OP_425J2_127_3477_n2194), .CO(
        DP_OP_425J2_127_3477_n1369), .S(DP_OP_425J2_127_3477_n1370) );
  FADDX1_HVT DP_OP_425J2_127_3477_U781 ( .A(DP_OP_425J2_127_3477_n2106), .B(
        DP_OP_425J2_127_3477_n2624), .CI(DP_OP_425J2_127_3477_n2238), .CO(
        DP_OP_425J2_127_3477_n1367), .S(DP_OP_425J2_127_3477_n1368) );
  FADDX1_HVT DP_OP_425J2_127_3477_U780 ( .A(DP_OP_425J2_127_3477_n2675), .B(
        DP_OP_425J2_127_3477_n1974), .CI(DP_OP_425J2_127_3477_n1930), .CO(
        DP_OP_425J2_127_3477_n1365), .S(DP_OP_425J2_127_3477_n1366) );
  FADDX1_HVT DP_OP_425J2_127_3477_U779 ( .A(DP_OP_425J2_127_3477_n2360), .B(
        DP_OP_425J2_127_3477_n2245), .CI(DP_OP_425J2_127_3477_n2157), .CO(
        DP_OP_425J2_127_3477_n1363), .S(DP_OP_425J2_127_3477_n1364) );
  FADDX1_HVT DP_OP_425J2_127_3477_U778 ( .A(DP_OP_425J2_127_3477_n2902), .B(
        DP_OP_425J2_127_3477_n2018), .CI(DP_OP_425J2_127_3477_n2814), .CO(
        DP_OP_425J2_127_3477_n1361), .S(DP_OP_425J2_127_3477_n1362) );
  FADDX1_HVT DP_OP_425J2_127_3477_U777 ( .A(DP_OP_425J2_127_3477_n2719), .B(
        DP_OP_425J2_127_3477_n2374), .CI(DP_OP_425J2_127_3477_n2404), .CO(
        DP_OP_425J2_127_3477_n1359), .S(DP_OP_425J2_127_3477_n1360) );
  FADDX1_HVT DP_OP_425J2_127_3477_U776 ( .A(DP_OP_425J2_127_3477_n1577), .B(
        DP_OP_425J2_127_3477_n1563), .CI(DP_OP_425J2_127_3477_n1565), .CO(
        DP_OP_425J2_127_3477_n1357), .S(DP_OP_425J2_127_3477_n1358) );
  FADDX1_HVT DP_OP_425J2_127_3477_U775 ( .A(DP_OP_425J2_127_3477_n1575), .B(
        DP_OP_425J2_127_3477_n1567), .CI(DP_OP_425J2_127_3477_n1569), .CO(
        DP_OP_425J2_127_3477_n1355), .S(DP_OP_425J2_127_3477_n1356) );
  FADDX1_HVT DP_OP_425J2_127_3477_U774 ( .A(DP_OP_425J2_127_3477_n1573), .B(
        DP_OP_425J2_127_3477_n1571), .CI(DP_OP_425J2_127_3477_n1561), .CO(
        DP_OP_425J2_127_3477_n1353), .S(DP_OP_425J2_127_3477_n1354) );
  FADDX1_HVT DP_OP_425J2_127_3477_U773 ( .A(DP_OP_425J2_127_3477_n1559), .B(
        DP_OP_425J2_127_3477_n1533), .CI(DP_OP_425J2_127_3477_n1529), .CO(
        DP_OP_425J2_127_3477_n1351), .S(DP_OP_425J2_127_3477_n1352) );
  FADDX1_HVT DP_OP_425J2_127_3477_U772 ( .A(DP_OP_425J2_127_3477_n1557), .B(
        DP_OP_425J2_127_3477_n1535), .CI(DP_OP_425J2_127_3477_n1531), .CO(
        DP_OP_425J2_127_3477_n1349), .S(DP_OP_425J2_127_3477_n1350) );
  FADDX1_HVT DP_OP_425J2_127_3477_U771 ( .A(DP_OP_425J2_127_3477_n1555), .B(
        DP_OP_425J2_127_3477_n1539), .CI(DP_OP_425J2_127_3477_n1537), .CO(
        DP_OP_425J2_127_3477_n1347), .S(DP_OP_425J2_127_3477_n1348) );
  FADDX1_HVT DP_OP_425J2_127_3477_U770 ( .A(DP_OP_425J2_127_3477_n1545), .B(
        DP_OP_425J2_127_3477_n1553), .CI(DP_OP_425J2_127_3477_n1541), .CO(
        DP_OP_425J2_127_3477_n1345), .S(DP_OP_425J2_127_3477_n1346) );
  FADDX1_HVT DP_OP_425J2_127_3477_U769 ( .A(DP_OP_425J2_127_3477_n1551), .B(
        DP_OP_425J2_127_3477_n1543), .CI(DP_OP_425J2_127_3477_n1549), .CO(
        DP_OP_425J2_127_3477_n1343), .S(DP_OP_425J2_127_3477_n1344) );
  FADDX1_HVT DP_OP_425J2_127_3477_U768 ( .A(DP_OP_425J2_127_3477_n1547), .B(
        DP_OP_425J2_127_3477_n1527), .CI(DP_OP_425J2_127_3477_n1525), .CO(
        DP_OP_425J2_127_3477_n1341), .S(DP_OP_425J2_127_3477_n1342) );
  FADDX1_HVT DP_OP_425J2_127_3477_U767 ( .A(DP_OP_425J2_127_3477_n1523), .B(
        DP_OP_425J2_127_3477_n1416), .CI(DP_OP_425J2_127_3477_n1513), .CO(
        DP_OP_425J2_127_3477_n1339), .S(DP_OP_425J2_127_3477_n1340) );
  FADDX1_HVT DP_OP_425J2_127_3477_U766 ( .A(DP_OP_425J2_127_3477_n1519), .B(
        DP_OP_425J2_127_3477_n1412), .CI(DP_OP_425J2_127_3477_n1418), .CO(
        DP_OP_425J2_127_3477_n1337), .S(DP_OP_425J2_127_3477_n1338) );
  FADDX1_HVT DP_OP_425J2_127_3477_U765 ( .A(DP_OP_425J2_127_3477_n1521), .B(
        DP_OP_425J2_127_3477_n1420), .CI(DP_OP_425J2_127_3477_n1414), .CO(
        DP_OP_425J2_127_3477_n1335), .S(DP_OP_425J2_127_3477_n1336) );
  FADDX1_HVT DP_OP_425J2_127_3477_U764 ( .A(DP_OP_425J2_127_3477_n1517), .B(
        DP_OP_425J2_127_3477_n1426), .CI(DP_OP_425J2_127_3477_n1422), .CO(
        DP_OP_425J2_127_3477_n1333), .S(DP_OP_425J2_127_3477_n1334) );
  FADDX1_HVT DP_OP_425J2_127_3477_U763 ( .A(DP_OP_425J2_127_3477_n1515), .B(
        DP_OP_425J2_127_3477_n1424), .CI(DP_OP_425J2_127_3477_n1410), .CO(
        DP_OP_425J2_127_3477_n1331), .S(DP_OP_425J2_127_3477_n1332) );
  FADDX1_HVT DP_OP_425J2_127_3477_U762 ( .A(DP_OP_425J2_127_3477_n1511), .B(
        DP_OP_425J2_127_3477_n1384), .CI(DP_OP_425J2_127_3477_n1376), .CO(
        DP_OP_425J2_127_3477_n1329), .S(DP_OP_425J2_127_3477_n1330) );
  FADDX1_HVT DP_OP_425J2_127_3477_U761 ( .A(DP_OP_425J2_127_3477_n1402), .B(
        DP_OP_425J2_127_3477_n1382), .CI(DP_OP_425J2_127_3477_n1378), .CO(
        DP_OP_425J2_127_3477_n1327), .S(DP_OP_425J2_127_3477_n1328) );
  FADDX1_HVT DP_OP_425J2_127_3477_U760 ( .A(DP_OP_425J2_127_3477_n1398), .B(
        DP_OP_425J2_127_3477_n1388), .CI(DP_OP_425J2_127_3477_n1380), .CO(
        DP_OP_425J2_127_3477_n1325), .S(DP_OP_425J2_127_3477_n1326) );
  FADDX1_HVT DP_OP_425J2_127_3477_U759 ( .A(DP_OP_425J2_127_3477_n1396), .B(
        DP_OP_425J2_127_3477_n1392), .CI(DP_OP_425J2_127_3477_n1386), .CO(
        DP_OP_425J2_127_3477_n1323), .S(DP_OP_425J2_127_3477_n1324) );
  FADDX1_HVT DP_OP_425J2_127_3477_U758 ( .A(DP_OP_425J2_127_3477_n1394), .B(
        DP_OP_425J2_127_3477_n1390), .CI(DP_OP_425J2_127_3477_n1408), .CO(
        DP_OP_425J2_127_3477_n1321), .S(DP_OP_425J2_127_3477_n1322) );
  FADDX1_HVT DP_OP_425J2_127_3477_U757 ( .A(DP_OP_425J2_127_3477_n1404), .B(
        DP_OP_425J2_127_3477_n1400), .CI(DP_OP_425J2_127_3477_n1406), .CO(
        DP_OP_425J2_127_3477_n1319), .S(DP_OP_425J2_127_3477_n1320) );
  FADDX1_HVT DP_OP_425J2_127_3477_U756 ( .A(DP_OP_425J2_127_3477_n1374), .B(
        DP_OP_425J2_127_3477_n1364), .CI(DP_OP_425J2_127_3477_n1360), .CO(
        DP_OP_425J2_127_3477_n1317), .S(DP_OP_425J2_127_3477_n1318) );
  FADDX1_HVT DP_OP_425J2_127_3477_U755 ( .A(DP_OP_425J2_127_3477_n1372), .B(
        DP_OP_425J2_127_3477_n1366), .CI(DP_OP_425J2_127_3477_n1362), .CO(
        DP_OP_425J2_127_3477_n1315), .S(DP_OP_425J2_127_3477_n1316) );
  FADDX1_HVT DP_OP_425J2_127_3477_U754 ( .A(DP_OP_425J2_127_3477_n1368), .B(
        DP_OP_425J2_127_3477_n1370), .CI(DP_OP_425J2_127_3477_n1509), .CO(
        DP_OP_425J2_127_3477_n1313), .S(DP_OP_425J2_127_3477_n1314) );
  FADDX1_HVT DP_OP_425J2_127_3477_U753 ( .A(DP_OP_425J2_127_3477_n1507), .B(
        DP_OP_425J2_127_3477_n1505), .CI(DP_OP_425J2_127_3477_n1503), .CO(
        DP_OP_425J2_127_3477_n1311), .S(DP_OP_425J2_127_3477_n1312) );
  FADDX1_HVT DP_OP_425J2_127_3477_U752 ( .A(DP_OP_425J2_127_3477_n1501), .B(
        DP_OP_425J2_127_3477_n1499), .CI(DP_OP_425J2_127_3477_n1493), .CO(
        DP_OP_425J2_127_3477_n1309), .S(DP_OP_425J2_127_3477_n1310) );
  FADDX1_HVT DP_OP_425J2_127_3477_U751 ( .A(DP_OP_425J2_127_3477_n1495), .B(
        DP_OP_425J2_127_3477_n1358), .CI(DP_OP_425J2_127_3477_n1354), .CO(
        DP_OP_425J2_127_3477_n1307), .S(DP_OP_425J2_127_3477_n1308) );
  FADDX1_HVT DP_OP_425J2_127_3477_U750 ( .A(DP_OP_425J2_127_3477_n1497), .B(
        DP_OP_425J2_127_3477_n1489), .CI(DP_OP_425J2_127_3477_n1356), .CO(
        DP_OP_425J2_127_3477_n1305), .S(DP_OP_425J2_127_3477_n1306) );
  FADDX1_HVT DP_OP_425J2_127_3477_U749 ( .A(DP_OP_425J2_127_3477_n1491), .B(
        DP_OP_425J2_127_3477_n1487), .CI(DP_OP_425J2_127_3477_n1485), .CO(
        DP_OP_425J2_127_3477_n1303), .S(DP_OP_425J2_127_3477_n1304) );
  FADDX1_HVT DP_OP_425J2_127_3477_U748 ( .A(DP_OP_425J2_127_3477_n1352), .B(
        DP_OP_425J2_127_3477_n1346), .CI(DP_OP_425J2_127_3477_n1342), .CO(
        DP_OP_425J2_127_3477_n1301), .S(DP_OP_425J2_127_3477_n1302) );
  FADDX1_HVT DP_OP_425J2_127_3477_U747 ( .A(DP_OP_425J2_127_3477_n1483), .B(
        DP_OP_425J2_127_3477_n1344), .CI(DP_OP_425J2_127_3477_n1350), .CO(
        DP_OP_425J2_127_3477_n1299), .S(DP_OP_425J2_127_3477_n1300) );
  FADDX1_HVT DP_OP_425J2_127_3477_U746 ( .A(DP_OP_425J2_127_3477_n1481), .B(
        DP_OP_425J2_127_3477_n1348), .CI(DP_OP_425J2_127_3477_n1477), .CO(
        DP_OP_425J2_127_3477_n1297), .S(DP_OP_425J2_127_3477_n1298) );
  FADDX1_HVT DP_OP_425J2_127_3477_U745 ( .A(DP_OP_425J2_127_3477_n1479), .B(
        DP_OP_425J2_127_3477_n1475), .CI(DP_OP_425J2_127_3477_n1473), .CO(
        DP_OP_425J2_127_3477_n1295), .S(DP_OP_425J2_127_3477_n1296) );
  FADDX1_HVT DP_OP_425J2_127_3477_U744 ( .A(DP_OP_425J2_127_3477_n1336), .B(
        DP_OP_425J2_127_3477_n1332), .CI(DP_OP_425J2_127_3477_n1471), .CO(
        DP_OP_425J2_127_3477_n1293), .S(DP_OP_425J2_127_3477_n1294) );
  FADDX1_HVT DP_OP_425J2_127_3477_U743 ( .A(DP_OP_425J2_127_3477_n1338), .B(
        DP_OP_425J2_127_3477_n1340), .CI(DP_OP_425J2_127_3477_n1334), .CO(
        DP_OP_425J2_127_3477_n1291), .S(DP_OP_425J2_127_3477_n1292) );
  FADDX1_HVT DP_OP_425J2_127_3477_U742 ( .A(DP_OP_425J2_127_3477_n1330), .B(
        DP_OP_425J2_127_3477_n1322), .CI(DP_OP_425J2_127_3477_n1320), .CO(
        DP_OP_425J2_127_3477_n1289), .S(DP_OP_425J2_127_3477_n1290) );
  FADDX1_HVT DP_OP_425J2_127_3477_U741 ( .A(DP_OP_425J2_127_3477_n1326), .B(
        DP_OP_425J2_127_3477_n1328), .CI(DP_OP_425J2_127_3477_n1324), .CO(
        DP_OP_425J2_127_3477_n1287), .S(DP_OP_425J2_127_3477_n1288) );
  FADDX1_HVT DP_OP_425J2_127_3477_U740 ( .A(DP_OP_425J2_127_3477_n1318), .B(
        DP_OP_425J2_127_3477_n1316), .CI(DP_OP_425J2_127_3477_n1469), .CO(
        DP_OP_425J2_127_3477_n1285), .S(DP_OP_425J2_127_3477_n1286) );
  FADDX1_HVT DP_OP_425J2_127_3477_U739 ( .A(DP_OP_425J2_127_3477_n1467), .B(
        DP_OP_425J2_127_3477_n1314), .CI(DP_OP_425J2_127_3477_n1465), .CO(
        DP_OP_425J2_127_3477_n1283), .S(DP_OP_425J2_127_3477_n1284) );
  FADDX1_HVT DP_OP_425J2_127_3477_U738 ( .A(DP_OP_425J2_127_3477_n1463), .B(
        DP_OP_425J2_127_3477_n1312), .CI(DP_OP_425J2_127_3477_n1310), .CO(
        DP_OP_425J2_127_3477_n1281), .S(DP_OP_425J2_127_3477_n1282) );
  FADDX1_HVT DP_OP_425J2_127_3477_U737 ( .A(DP_OP_425J2_127_3477_n1461), .B(
        DP_OP_425J2_127_3477_n1459), .CI(DP_OP_425J2_127_3477_n1457), .CO(
        DP_OP_425J2_127_3477_n1279), .S(DP_OP_425J2_127_3477_n1280) );
  FADDX1_HVT DP_OP_425J2_127_3477_U736 ( .A(DP_OP_425J2_127_3477_n1308), .B(
        DP_OP_425J2_127_3477_n1306), .CI(DP_OP_425J2_127_3477_n1455), .CO(
        DP_OP_425J2_127_3477_n1277), .S(DP_OP_425J2_127_3477_n1278) );
  FADDX1_HVT DP_OP_425J2_127_3477_U735 ( .A(DP_OP_425J2_127_3477_n1304), .B(
        DP_OP_425J2_127_3477_n1453), .CI(DP_OP_425J2_127_3477_n1449), .CO(
        DP_OP_425J2_127_3477_n1275), .S(DP_OP_425J2_127_3477_n1276) );
  FADDX1_HVT DP_OP_425J2_127_3477_U734 ( .A(DP_OP_425J2_127_3477_n1302), .B(
        DP_OP_425J2_127_3477_n1300), .CI(DP_OP_425J2_127_3477_n1296), .CO(
        DP_OP_425J2_127_3477_n1273), .S(DP_OP_425J2_127_3477_n1274) );
  FADDX1_HVT DP_OP_425J2_127_3477_U733 ( .A(DP_OP_425J2_127_3477_n1451), .B(
        DP_OP_425J2_127_3477_n1298), .CI(DP_OP_425J2_127_3477_n1292), .CO(
        DP_OP_425J2_127_3477_n1271), .S(DP_OP_425J2_127_3477_n1272) );
  FADDX1_HVT DP_OP_425J2_127_3477_U732 ( .A(DP_OP_425J2_127_3477_n1294), .B(
        DP_OP_425J2_127_3477_n1290), .CI(DP_OP_425J2_127_3477_n1288), .CO(
        DP_OP_425J2_127_3477_n1269), .S(DP_OP_425J2_127_3477_n1270) );
  FADDX1_HVT DP_OP_425J2_127_3477_U731 ( .A(DP_OP_425J2_127_3477_n1447), .B(
        DP_OP_425J2_127_3477_n1286), .CI(DP_OP_425J2_127_3477_n1445), .CO(
        DP_OP_425J2_127_3477_n1267), .S(DP_OP_425J2_127_3477_n1268) );
  FADDX1_HVT DP_OP_425J2_127_3477_U730 ( .A(DP_OP_425J2_127_3477_n1284), .B(
        DP_OP_425J2_127_3477_n1443), .CI(DP_OP_425J2_127_3477_n1282), .CO(
        DP_OP_425J2_127_3477_n1265), .S(DP_OP_425J2_127_3477_n1266) );
  FADDX1_HVT DP_OP_425J2_127_3477_U729 ( .A(DP_OP_425J2_127_3477_n1441), .B(
        DP_OP_425J2_127_3477_n1280), .CI(DP_OP_425J2_127_3477_n1439), .CO(
        DP_OP_425J2_127_3477_n1263), .S(DP_OP_425J2_127_3477_n1264) );
  FADDX1_HVT DP_OP_425J2_127_3477_U728 ( .A(DP_OP_425J2_127_3477_n1278), .B(
        DP_OP_425J2_127_3477_n1437), .CI(DP_OP_425J2_127_3477_n1276), .CO(
        DP_OP_425J2_127_3477_n1261), .S(DP_OP_425J2_127_3477_n1262) );
  FADDX1_HVT DP_OP_425J2_127_3477_U727 ( .A(DP_OP_425J2_127_3477_n1274), .B(
        DP_OP_425J2_127_3477_n1272), .CI(DP_OP_425J2_127_3477_n1435), .CO(
        DP_OP_425J2_127_3477_n1259), .S(DP_OP_425J2_127_3477_n1260) );
  FADDX1_HVT DP_OP_425J2_127_3477_U726 ( .A(DP_OP_425J2_127_3477_n1270), .B(
        DP_OP_425J2_127_3477_n1268), .CI(DP_OP_425J2_127_3477_n1433), .CO(
        DP_OP_425J2_127_3477_n1257), .S(DP_OP_425J2_127_3477_n1258) );
  FADDX1_HVT DP_OP_425J2_127_3477_U725 ( .A(DP_OP_425J2_127_3477_n1266), .B(
        DP_OP_425J2_127_3477_n1431), .CI(DP_OP_425J2_127_3477_n1264), .CO(
        DP_OP_425J2_127_3477_n1255), .S(DP_OP_425J2_127_3477_n1256) );
  FADDX1_HVT DP_OP_425J2_127_3477_U724 ( .A(DP_OP_425J2_127_3477_n1262), .B(
        DP_OP_425J2_127_3477_n1429), .CI(DP_OP_425J2_127_3477_n1260), .CO(
        DP_OP_425J2_127_3477_n1253), .S(DP_OP_425J2_127_3477_n1254) );
  FADDX1_HVT DP_OP_425J2_127_3477_U723 ( .A(DP_OP_425J2_127_3477_n1258), .B(
        DP_OP_425J2_127_3477_n1427), .CI(DP_OP_425J2_127_3477_n1256), .CO(
        DP_OP_425J2_127_3477_n1251), .S(DP_OP_425J2_127_3477_n1252) );
  HADDX1_HVT DP_OP_425J2_127_3477_U722 ( .A0(DP_OP_425J2_127_3477_n2353), .B0(
        DP_OP_425J2_127_3477_n2440), .C1(DP_OP_425J2_127_3477_n1249), .SO(
        DP_OP_425J2_127_3477_n1250) );
  FADDX1_HVT DP_OP_425J2_127_3477_U721 ( .A(DP_OP_425J2_127_3477_n2704), .B(
        DP_OP_425J2_127_3477_n1827), .CI(DP_OP_425J2_127_3477_n2396), .CO(
        DP_OP_425J2_127_3477_n1247), .S(DP_OP_425J2_127_3477_n1248) );
  FADDX1_HVT DP_OP_425J2_127_3477_U720 ( .A(DP_OP_425J2_127_3477_n2003), .B(
        DP_OP_425J2_127_3477_n2047), .CI(DP_OP_425J2_127_3477_n1959), .CO(
        DP_OP_425J2_127_3477_n1245), .S(DP_OP_425J2_127_3477_n1246) );
  FADDX1_HVT DP_OP_425J2_127_3477_U719 ( .A(DP_OP_425J2_127_3477_n2836), .B(
        DP_OP_425J2_127_3477_n2528), .CI(DP_OP_425J2_127_3477_n2748), .CO(
        DP_OP_425J2_127_3477_n1243), .S(DP_OP_425J2_127_3477_n1244) );
  FADDX1_HVT DP_OP_425J2_127_3477_U718 ( .A(DP_OP_425J2_127_3477_n1871), .B(
        DP_OP_425J2_127_3477_n2484), .CI(DP_OP_425J2_127_3477_n2179), .CO(
        DP_OP_425J2_127_3477_n1241), .S(DP_OP_425J2_127_3477_n1242) );
  FADDX1_HVT DP_OP_425J2_127_3477_U717 ( .A(DP_OP_425J2_127_3477_n2091), .B(
        DP_OP_425J2_127_3477_n2572), .CI(DP_OP_425J2_127_3477_n1915), .CO(
        DP_OP_425J2_127_3477_n1239), .S(DP_OP_425J2_127_3477_n1240) );
  FADDX1_HVT DP_OP_425J2_127_3477_U716 ( .A(DP_OP_425J2_127_3477_n2616), .B(
        DP_OP_425J2_127_3477_n2267), .CI(DP_OP_425J2_127_3477_n2880), .CO(
        DP_OP_425J2_127_3477_n1237), .S(DP_OP_425J2_127_3477_n1238) );
  FADDX1_HVT DP_OP_425J2_127_3477_U715 ( .A(DP_OP_425J2_127_3477_n2135), .B(
        DP_OP_425J2_127_3477_n2311), .CI(DP_OP_425J2_127_3477_n2660), .CO(
        DP_OP_425J2_127_3477_n1235), .S(DP_OP_425J2_127_3477_n1236) );
  FADDX1_HVT DP_OP_425J2_127_3477_U714 ( .A(DP_OP_425J2_127_3477_n2792), .B(
        DP_OP_425J2_127_3477_n2223), .CI(DP_OP_425J2_127_3477_n2112), .CO(
        DP_OP_425J2_127_3477_n1233), .S(DP_OP_425J2_127_3477_n1234) );
  FADDX1_HVT DP_OP_425J2_127_3477_U713 ( .A(DP_OP_425J2_127_3477_n2637), .B(
        DP_OP_425J2_127_3477_n2579), .CI(DP_OP_425J2_127_3477_n2288), .CO(
        DP_OP_425J2_127_3477_n1231), .S(DP_OP_425J2_127_3477_n1232) );
  FADDX1_HVT DP_OP_425J2_127_3477_U712 ( .A(DP_OP_425J2_127_3477_n2417), .B(
        DP_OP_425J2_127_3477_n2725), .CI(DP_OP_425J2_127_3477_n2068), .CO(
        DP_OP_425J2_127_3477_n1229), .S(DP_OP_425J2_127_3477_n1230) );
  FADDX1_HVT DP_OP_425J2_127_3477_U711 ( .A(DP_OP_425J2_127_3477_n2549), .B(
        DP_OP_425J2_127_3477_n1966), .CI(DP_OP_425J2_127_3477_n2274), .CO(
        DP_OP_425J2_127_3477_n1227), .S(DP_OP_425J2_127_3477_n1228) );
  FADDX1_HVT DP_OP_425J2_127_3477_U710 ( .A(DP_OP_425J2_127_3477_n1848), .B(
        DP_OP_425J2_127_3477_n2149), .CI(DP_OP_425J2_127_3477_n2142), .CO(
        DP_OP_425J2_127_3477_n1225), .S(DP_OP_425J2_127_3477_n1226) );
  FADDX1_HVT DP_OP_425J2_127_3477_U709 ( .A(DP_OP_425J2_127_3477_n2332), .B(
        DP_OP_425J2_127_3477_n2410), .CI(DP_OP_425J2_127_3477_n2806), .CO(
        DP_OP_425J2_127_3477_n1223), .S(DP_OP_425J2_127_3477_n1224) );
  FADDX1_HVT DP_OP_425J2_127_3477_U708 ( .A(DP_OP_425J2_127_3477_n2200), .B(
        DP_OP_425J2_127_3477_n2535), .CI(DP_OP_425J2_127_3477_n2281), .CO(
        DP_OP_425J2_127_3477_n1221), .S(DP_OP_425J2_127_3477_n1222) );
  FADDX1_HVT DP_OP_425J2_127_3477_U707 ( .A(DP_OP_425J2_127_3477_n2461), .B(
        DP_OP_425J2_127_3477_n1783), .CI(DP_OP_425J2_127_3477_n2054), .CO(
        DP_OP_425J2_127_3477_n1219), .S(DP_OP_425J2_127_3477_n1220) );
  FADDX1_HVT DP_OP_425J2_127_3477_U706 ( .A(DP_OP_425J2_127_3477_n2887), .B(
        DP_OP_425J2_127_3477_n2061), .CI(DP_OP_425J2_127_3477_n2318), .CO(
        DP_OP_425J2_127_3477_n1217), .S(DP_OP_425J2_127_3477_n1218) );
  FADDX1_HVT DP_OP_425J2_127_3477_U705 ( .A(DP_OP_425J2_127_3477_n2593), .B(
        DP_OP_425J2_127_3477_n2325), .CI(DP_OP_425J2_127_3477_n2894), .CO(
        DP_OP_425J2_127_3477_n1215), .S(DP_OP_425J2_127_3477_n1216) );
  FADDX1_HVT DP_OP_425J2_127_3477_U704 ( .A(DP_OP_425J2_127_3477_n2843), .B(
        DP_OP_425J2_127_3477_n2586), .CI(DP_OP_425J2_127_3477_n2850), .CO(
        DP_OP_425J2_127_3477_n1213), .S(DP_OP_425J2_127_3477_n1214) );
  FADDX1_HVT DP_OP_425J2_127_3477_U703 ( .A(DP_OP_425J2_127_3477_n1980), .B(
        DP_OP_425J2_127_3477_n1841), .CI(DP_OP_425J2_127_3477_n2542), .CO(
        DP_OP_425J2_127_3477_n1211), .S(DP_OP_425J2_127_3477_n1212) );
  FADDX1_HVT DP_OP_425J2_127_3477_U702 ( .A(DP_OP_425J2_127_3477_n2024), .B(
        DP_OP_425J2_127_3477_n2630), .CI(DP_OP_425J2_127_3477_n2711), .CO(
        DP_OP_425J2_127_3477_n1209), .S(DP_OP_425J2_127_3477_n1210) );
  FADDX1_HVT DP_OP_425J2_127_3477_U701 ( .A(DP_OP_425J2_127_3477_n2681), .B(
        DP_OP_425J2_127_3477_n2498), .CI(DP_OP_425J2_127_3477_n1936), .CO(
        DP_OP_425J2_127_3477_n1207), .S(DP_OP_425J2_127_3477_n1208) );
  FADDX1_HVT DP_OP_425J2_127_3477_U700 ( .A(DP_OP_425J2_127_3477_n2755), .B(
        DP_OP_425J2_127_3477_n2857), .CI(DP_OP_425J2_127_3477_n2505), .CO(
        DP_OP_425J2_127_3477_n1205), .S(DP_OP_425J2_127_3477_n1206) );
  FADDX1_HVT DP_OP_425J2_127_3477_U699 ( .A(DP_OP_425J2_127_3477_n2230), .B(
        DP_OP_425J2_127_3477_n2447), .CI(DP_OP_425J2_127_3477_n2186), .CO(
        DP_OP_425J2_127_3477_n1203), .S(DP_OP_425J2_127_3477_n1204) );
  FADDX1_HVT DP_OP_425J2_127_3477_U698 ( .A(DP_OP_425J2_127_3477_n2769), .B(
        DP_OP_425J2_127_3477_n1892), .CI(DP_OP_425J2_127_3477_n1922), .CO(
        DP_OP_425J2_127_3477_n1201), .S(DP_OP_425J2_127_3477_n1202) );
  FADDX1_HVT DP_OP_425J2_127_3477_U697 ( .A(DP_OP_425J2_127_3477_n2098), .B(
        DP_OP_425J2_127_3477_n2667), .CI(DP_OP_425J2_127_3477_n1878), .CO(
        DP_OP_425J2_127_3477_n1199), .S(DP_OP_425J2_127_3477_n1200) );
  FADDX1_HVT DP_OP_425J2_127_3477_U696 ( .A(DP_OP_425J2_127_3477_n2762), .B(
        DP_OP_425J2_127_3477_n2454), .CI(DP_OP_425J2_127_3477_n2010), .CO(
        DP_OP_425J2_127_3477_n1197), .S(DP_OP_425J2_127_3477_n1198) );
  FADDX1_HVT DP_OP_425J2_127_3477_U695 ( .A(DP_OP_425J2_127_3477_n1885), .B(
        DP_OP_425J2_127_3477_n1834), .CI(DP_OP_425J2_127_3477_n2366), .CO(
        DP_OP_425J2_127_3477_n1195), .S(DP_OP_425J2_127_3477_n1196) );
  FADDX1_HVT DP_OP_425J2_127_3477_U694 ( .A(DP_OP_425J2_127_3477_n2491), .B(
        DP_OP_425J2_127_3477_n2799), .CI(DP_OP_425J2_127_3477_n2193), .CO(
        DP_OP_425J2_127_3477_n1193), .S(DP_OP_425J2_127_3477_n1194) );
  FADDX1_HVT DP_OP_425J2_127_3477_U693 ( .A(DP_OP_425J2_127_3477_n2105), .B(
        DP_OP_425J2_127_3477_n2623), .CI(DP_OP_425J2_127_3477_n2237), .CO(
        DP_OP_425J2_127_3477_n1191), .S(DP_OP_425J2_127_3477_n1192) );
  FADDX1_HVT DP_OP_425J2_127_3477_U692 ( .A(DP_OP_425J2_127_3477_n2674), .B(
        DP_OP_425J2_127_3477_n1973), .CI(DP_OP_425J2_127_3477_n1929), .CO(
        DP_OP_425J2_127_3477_n1189), .S(DP_OP_425J2_127_3477_n1190) );
  FADDX1_HVT DP_OP_425J2_127_3477_U691 ( .A(DP_OP_425J2_127_3477_n2359), .B(
        DP_OP_425J2_127_3477_n2244), .CI(DP_OP_425J2_127_3477_n2156), .CO(
        DP_OP_425J2_127_3477_n1187), .S(DP_OP_425J2_127_3477_n1188) );
  FADDX1_HVT DP_OP_425J2_127_3477_U690 ( .A(DP_OP_425J2_127_3477_n2901), .B(
        DP_OP_425J2_127_3477_n2017), .CI(DP_OP_425J2_127_3477_n2813), .CO(
        DP_OP_425J2_127_3477_n1185), .S(DP_OP_425J2_127_3477_n1186) );
  FADDX1_HVT DP_OP_425J2_127_3477_U689 ( .A(DP_OP_425J2_127_3477_n2718), .B(
        DP_OP_425J2_127_3477_n2373), .CI(DP_OP_425J2_127_3477_n2403), .CO(
        DP_OP_425J2_127_3477_n1183), .S(DP_OP_425J2_127_3477_n1184) );
  FADDX1_HVT DP_OP_425J2_127_3477_U688 ( .A(DP_OP_425J2_127_3477_n1250), .B(
        DP_OP_425J2_127_3477_n1425), .CI(DP_OP_425J2_127_3477_n1411), .CO(
        DP_OP_425J2_127_3477_n1181), .S(DP_OP_425J2_127_3477_n1182) );
  FADDX1_HVT DP_OP_425J2_127_3477_U687 ( .A(DP_OP_425J2_127_3477_n1423), .B(
        DP_OP_425J2_127_3477_n1413), .CI(DP_OP_425J2_127_3477_n1409), .CO(
        DP_OP_425J2_127_3477_n1179), .S(DP_OP_425J2_127_3477_n1180) );
  FADDX1_HVT DP_OP_425J2_127_3477_U686 ( .A(DP_OP_425J2_127_3477_n1421), .B(
        DP_OP_425J2_127_3477_n1415), .CI(DP_OP_425J2_127_3477_n1417), .CO(
        DP_OP_425J2_127_3477_n1177), .S(DP_OP_425J2_127_3477_n1178) );
  FADDX1_HVT DP_OP_425J2_127_3477_U685 ( .A(DP_OP_425J2_127_3477_n1419), .B(
        DP_OP_425J2_127_3477_n1407), .CI(DP_OP_425J2_127_3477_n1405), .CO(
        DP_OP_425J2_127_3477_n1175), .S(DP_OP_425J2_127_3477_n1176) );
  FADDX1_HVT DP_OP_425J2_127_3477_U684 ( .A(DP_OP_425J2_127_3477_n1403), .B(
        DP_OP_425J2_127_3477_n1381), .CI(DP_OP_425J2_127_3477_n1375), .CO(
        DP_OP_425J2_127_3477_n1173), .S(DP_OP_425J2_127_3477_n1174) );
  FADDX1_HVT DP_OP_425J2_127_3477_U683 ( .A(DP_OP_425J2_127_3477_n1401), .B(
        DP_OP_425J2_127_3477_n1383), .CI(DP_OP_425J2_127_3477_n1377), .CO(
        DP_OP_425J2_127_3477_n1171), .S(DP_OP_425J2_127_3477_n1172) );
  FADDX1_HVT DP_OP_425J2_127_3477_U682 ( .A(DP_OP_425J2_127_3477_n1399), .B(
        DP_OP_425J2_127_3477_n1385), .CI(DP_OP_425J2_127_3477_n1379), .CO(
        DP_OP_425J2_127_3477_n1169), .S(DP_OP_425J2_127_3477_n1170) );
  FADDX1_HVT DP_OP_425J2_127_3477_U681 ( .A(DP_OP_425J2_127_3477_n1391), .B(
        DP_OP_425J2_127_3477_n1389), .CI(DP_OP_425J2_127_3477_n1387), .CO(
        DP_OP_425J2_127_3477_n1167), .S(DP_OP_425J2_127_3477_n1168) );
  FADDX1_HVT DP_OP_425J2_127_3477_U680 ( .A(DP_OP_425J2_127_3477_n1397), .B(
        DP_OP_425J2_127_3477_n1393), .CI(DP_OP_425J2_127_3477_n1395), .CO(
        DP_OP_425J2_127_3477_n1165), .S(DP_OP_425J2_127_3477_n1166) );
  FADDX1_HVT DP_OP_425J2_127_3477_U679 ( .A(DP_OP_425J2_127_3477_n1373), .B(
        DP_OP_425J2_127_3477_n1244), .CI(DP_OP_425J2_127_3477_n1361), .CO(
        DP_OP_425J2_127_3477_n1163), .S(DP_OP_425J2_127_3477_n1164) );
  FADDX1_HVT DP_OP_425J2_127_3477_U678 ( .A(DP_OP_425J2_127_3477_n1369), .B(
        DP_OP_425J2_127_3477_n1242), .CI(DP_OP_425J2_127_3477_n1359), .CO(
        DP_OP_425J2_127_3477_n1161), .S(DP_OP_425J2_127_3477_n1162) );
  FADDX1_HVT DP_OP_425J2_127_3477_U677 ( .A(DP_OP_425J2_127_3477_n1367), .B(
        DP_OP_425J2_127_3477_n1238), .CI(DP_OP_425J2_127_3477_n1236), .CO(
        DP_OP_425J2_127_3477_n1159), .S(DP_OP_425J2_127_3477_n1160) );
  FADDX1_HVT DP_OP_425J2_127_3477_U676 ( .A(DP_OP_425J2_127_3477_n1371), .B(
        DP_OP_425J2_127_3477_n1246), .CI(DP_OP_425J2_127_3477_n1240), .CO(
        DP_OP_425J2_127_3477_n1157), .S(DP_OP_425J2_127_3477_n1158) );
  FADDX1_HVT DP_OP_425J2_127_3477_U675 ( .A(DP_OP_425J2_127_3477_n1365), .B(
        DP_OP_425J2_127_3477_n1363), .CI(DP_OP_425J2_127_3477_n1248), .CO(
        DP_OP_425J2_127_3477_n1155), .S(DP_OP_425J2_127_3477_n1156) );
  FADDX1_HVT DP_OP_425J2_127_3477_U674 ( .A(DP_OP_425J2_127_3477_n1234), .B(
        DP_OP_425J2_127_3477_n1224), .CI(DP_OP_425J2_127_3477_n1206), .CO(
        DP_OP_425J2_127_3477_n1153), .S(DP_OP_425J2_127_3477_n1154) );
  FADDX1_HVT DP_OP_425J2_127_3477_U673 ( .A(DP_OP_425J2_127_3477_n1226), .B(
        DP_OP_425J2_127_3477_n1208), .CI(DP_OP_425J2_127_3477_n1200), .CO(
        DP_OP_425J2_127_3477_n1151), .S(DP_OP_425J2_127_3477_n1152) );
  FADDX1_HVT DP_OP_425J2_127_3477_U672 ( .A(DP_OP_425J2_127_3477_n1222), .B(
        DP_OP_425J2_127_3477_n1210), .CI(DP_OP_425J2_127_3477_n1204), .CO(
        DP_OP_425J2_127_3477_n1149), .S(DP_OP_425J2_127_3477_n1150) );
  FADDX1_HVT DP_OP_425J2_127_3477_U671 ( .A(DP_OP_425J2_127_3477_n1218), .B(
        DP_OP_425J2_127_3477_n1212), .CI(DP_OP_425J2_127_3477_n1202), .CO(
        DP_OP_425J2_127_3477_n1147), .S(DP_OP_425J2_127_3477_n1148) );
  FADDX1_HVT DP_OP_425J2_127_3477_U670 ( .A(DP_OP_425J2_127_3477_n1220), .B(
        DP_OP_425J2_127_3477_n1232), .CI(DP_OP_425J2_127_3477_n1230), .CO(
        DP_OP_425J2_127_3477_n1145), .S(DP_OP_425J2_127_3477_n1146) );
  FADDX1_HVT DP_OP_425J2_127_3477_U669 ( .A(DP_OP_425J2_127_3477_n1216), .B(
        DP_OP_425J2_127_3477_n1214), .CI(DP_OP_425J2_127_3477_n1228), .CO(
        DP_OP_425J2_127_3477_n1143), .S(DP_OP_425J2_127_3477_n1144) );
  FADDX1_HVT DP_OP_425J2_127_3477_U668 ( .A(DP_OP_425J2_127_3477_n1198), .B(
        DP_OP_425J2_127_3477_n1188), .CI(DP_OP_425J2_127_3477_n1186), .CO(
        DP_OP_425J2_127_3477_n1141), .S(DP_OP_425J2_127_3477_n1142) );
  FADDX1_HVT DP_OP_425J2_127_3477_U667 ( .A(DP_OP_425J2_127_3477_n1194), .B(
        DP_OP_425J2_127_3477_n1190), .CI(DP_OP_425J2_127_3477_n1184), .CO(
        DP_OP_425J2_127_3477_n1139), .S(DP_OP_425J2_127_3477_n1140) );
  FADDX1_HVT DP_OP_425J2_127_3477_U666 ( .A(DP_OP_425J2_127_3477_n1196), .B(
        DP_OP_425J2_127_3477_n1192), .CI(DP_OP_425J2_127_3477_n1357), .CO(
        DP_OP_425J2_127_3477_n1137), .S(DP_OP_425J2_127_3477_n1138) );
  FADDX1_HVT DP_OP_425J2_127_3477_U665 ( .A(DP_OP_425J2_127_3477_n1355), .B(
        DP_OP_425J2_127_3477_n1353), .CI(DP_OP_425J2_127_3477_n1351), .CO(
        DP_OP_425J2_127_3477_n1135), .S(DP_OP_425J2_127_3477_n1136) );
  FADDX1_HVT DP_OP_425J2_127_3477_U664 ( .A(DP_OP_425J2_127_3477_n1349), .B(
        DP_OP_425J2_127_3477_n1343), .CI(DP_OP_425J2_127_3477_n1341), .CO(
        DP_OP_425J2_127_3477_n1133), .S(DP_OP_425J2_127_3477_n1134) );
  FADDX1_HVT DP_OP_425J2_127_3477_U663 ( .A(DP_OP_425J2_127_3477_n1347), .B(
        DP_OP_425J2_127_3477_n1345), .CI(DP_OP_425J2_127_3477_n1182), .CO(
        DP_OP_425J2_127_3477_n1131), .S(DP_OP_425J2_127_3477_n1132) );
  FADDX1_HVT DP_OP_425J2_127_3477_U662 ( .A(DP_OP_425J2_127_3477_n1339), .B(
        DP_OP_425J2_127_3477_n1180), .CI(DP_OP_425J2_127_3477_n1178), .CO(
        DP_OP_425J2_127_3477_n1129), .S(DP_OP_425J2_127_3477_n1130) );
  FADDX1_HVT DP_OP_425J2_127_3477_U661 ( .A(DP_OP_425J2_127_3477_n1337), .B(
        DP_OP_425J2_127_3477_n1333), .CI(DP_OP_425J2_127_3477_n1331), .CO(
        DP_OP_425J2_127_3477_n1127), .S(DP_OP_425J2_127_3477_n1128) );
  FADDX1_HVT DP_OP_425J2_127_3477_U660 ( .A(DP_OP_425J2_127_3477_n1335), .B(
        DP_OP_425J2_127_3477_n1176), .CI(DP_OP_425J2_127_3477_n1329), .CO(
        DP_OP_425J2_127_3477_n1125), .S(DP_OP_425J2_127_3477_n1126) );
  FADDX1_HVT DP_OP_425J2_127_3477_U659 ( .A(DP_OP_425J2_127_3477_n1168), .B(
        DP_OP_425J2_127_3477_n1172), .CI(DP_OP_425J2_127_3477_n1174), .CO(
        DP_OP_425J2_127_3477_n1123), .S(DP_OP_425J2_127_3477_n1124) );
  FADDX1_HVT DP_OP_425J2_127_3477_U658 ( .A(DP_OP_425J2_127_3477_n1327), .B(
        DP_OP_425J2_127_3477_n1170), .CI(DP_OP_425J2_127_3477_n1166), .CO(
        DP_OP_425J2_127_3477_n1121), .S(DP_OP_425J2_127_3477_n1122) );
  FADDX1_HVT DP_OP_425J2_127_3477_U657 ( .A(DP_OP_425J2_127_3477_n1325), .B(
        DP_OP_425J2_127_3477_n1319), .CI(DP_OP_425J2_127_3477_n1321), .CO(
        DP_OP_425J2_127_3477_n1119), .S(DP_OP_425J2_127_3477_n1120) );
  FADDX1_HVT DP_OP_425J2_127_3477_U656 ( .A(DP_OP_425J2_127_3477_n1323), .B(
        DP_OP_425J2_127_3477_n1317), .CI(DP_OP_425J2_127_3477_n1164), .CO(
        DP_OP_425J2_127_3477_n1117), .S(DP_OP_425J2_127_3477_n1118) );
  FADDX1_HVT DP_OP_425J2_127_3477_U655 ( .A(DP_OP_425J2_127_3477_n1315), .B(
        DP_OP_425J2_127_3477_n1162), .CI(DP_OP_425J2_127_3477_n1156), .CO(
        DP_OP_425J2_127_3477_n1115), .S(DP_OP_425J2_127_3477_n1116) );
  FADDX1_HVT DP_OP_425J2_127_3477_U654 ( .A(DP_OP_425J2_127_3477_n1160), .B(
        DP_OP_425J2_127_3477_n1158), .CI(DP_OP_425J2_127_3477_n1154), .CO(
        DP_OP_425J2_127_3477_n1113), .S(DP_OP_425J2_127_3477_n1114) );
  FADDX1_HVT DP_OP_425J2_127_3477_U653 ( .A(DP_OP_425J2_127_3477_n1148), .B(
        DP_OP_425J2_127_3477_n1144), .CI(DP_OP_425J2_127_3477_n1313), .CO(
        DP_OP_425J2_127_3477_n1111), .S(DP_OP_425J2_127_3477_n1112) );
  FADDX1_HVT DP_OP_425J2_127_3477_U652 ( .A(DP_OP_425J2_127_3477_n1150), .B(
        DP_OP_425J2_127_3477_n1146), .CI(DP_OP_425J2_127_3477_n1152), .CO(
        DP_OP_425J2_127_3477_n1109), .S(DP_OP_425J2_127_3477_n1110) );
  FADDX1_HVT DP_OP_425J2_127_3477_U651 ( .A(DP_OP_425J2_127_3477_n1142), .B(
        DP_OP_425J2_127_3477_n1309), .CI(DP_OP_425J2_127_3477_n1138), .CO(
        DP_OP_425J2_127_3477_n1107), .S(DP_OP_425J2_127_3477_n1108) );
  FADDX1_HVT DP_OP_425J2_127_3477_U650 ( .A(DP_OP_425J2_127_3477_n1140), .B(
        DP_OP_425J2_127_3477_n1311), .CI(DP_OP_425J2_127_3477_n1307), .CO(
        DP_OP_425J2_127_3477_n1105), .S(DP_OP_425J2_127_3477_n1106) );
  FADDX1_HVT DP_OP_425J2_127_3477_U649 ( .A(DP_OP_425J2_127_3477_n1305), .B(
        DP_OP_425J2_127_3477_n1136), .CI(DP_OP_425J2_127_3477_n1303), .CO(
        DP_OP_425J2_127_3477_n1103), .S(DP_OP_425J2_127_3477_n1104) );
  FADDX1_HVT DP_OP_425J2_127_3477_U648 ( .A(DP_OP_425J2_127_3477_n1301), .B(
        DP_OP_425J2_127_3477_n1132), .CI(DP_OP_425J2_127_3477_n1295), .CO(
        DP_OP_425J2_127_3477_n1101), .S(DP_OP_425J2_127_3477_n1102) );
  FADDX1_HVT DP_OP_425J2_127_3477_U647 ( .A(DP_OP_425J2_127_3477_n1299), .B(
        DP_OP_425J2_127_3477_n1134), .CI(DP_OP_425J2_127_3477_n1297), .CO(
        DP_OP_425J2_127_3477_n1099), .S(DP_OP_425J2_127_3477_n1100) );
  FADDX1_HVT DP_OP_425J2_127_3477_U646 ( .A(DP_OP_425J2_127_3477_n1293), .B(
        DP_OP_425J2_127_3477_n1128), .CI(DP_OP_425J2_127_3477_n1126), .CO(
        DP_OP_425J2_127_3477_n1097), .S(DP_OP_425J2_127_3477_n1098) );
  FADDX1_HVT DP_OP_425J2_127_3477_U645 ( .A(DP_OP_425J2_127_3477_n1291), .B(
        DP_OP_425J2_127_3477_n1130), .CI(DP_OP_425J2_127_3477_n1289), .CO(
        DP_OP_425J2_127_3477_n1095), .S(DP_OP_425J2_127_3477_n1096) );
  FADDX1_HVT DP_OP_425J2_127_3477_U644 ( .A(DP_OP_425J2_127_3477_n1287), .B(
        DP_OP_425J2_127_3477_n1124), .CI(DP_OP_425J2_127_3477_n1118), .CO(
        DP_OP_425J2_127_3477_n1093), .S(DP_OP_425J2_127_3477_n1094) );
  FADDX1_HVT DP_OP_425J2_127_3477_U643 ( .A(DP_OP_425J2_127_3477_n1120), .B(
        DP_OP_425J2_127_3477_n1122), .CI(DP_OP_425J2_127_3477_n1285), .CO(
        DP_OP_425J2_127_3477_n1091), .S(DP_OP_425J2_127_3477_n1092) );
  FADDX1_HVT DP_OP_425J2_127_3477_U642 ( .A(DP_OP_425J2_127_3477_n1116), .B(
        DP_OP_425J2_127_3477_n1114), .CI(DP_OP_425J2_127_3477_n1110), .CO(
        DP_OP_425J2_127_3477_n1089), .S(DP_OP_425J2_127_3477_n1090) );
  FADDX1_HVT DP_OP_425J2_127_3477_U641 ( .A(DP_OP_425J2_127_3477_n1112), .B(
        DP_OP_425J2_127_3477_n1283), .CI(DP_OP_425J2_127_3477_n1108), .CO(
        DP_OP_425J2_127_3477_n1087), .S(DP_OP_425J2_127_3477_n1088) );
  FADDX1_HVT DP_OP_425J2_127_3477_U640 ( .A(DP_OP_425J2_127_3477_n1281), .B(
        DP_OP_425J2_127_3477_n1279), .CI(DP_OP_425J2_127_3477_n1106), .CO(
        DP_OP_425J2_127_3477_n1085), .S(DP_OP_425J2_127_3477_n1086) );
  FADDX1_HVT DP_OP_425J2_127_3477_U639 ( .A(DP_OP_425J2_127_3477_n1277), .B(
        DP_OP_425J2_127_3477_n1104), .CI(DP_OP_425J2_127_3477_n1275), .CO(
        DP_OP_425J2_127_3477_n1083), .S(DP_OP_425J2_127_3477_n1084) );
  FADDX1_HVT DP_OP_425J2_127_3477_U638 ( .A(DP_OP_425J2_127_3477_n1273), .B(
        DP_OP_425J2_127_3477_n1271), .CI(DP_OP_425J2_127_3477_n1100), .CO(
        DP_OP_425J2_127_3477_n1081), .S(DP_OP_425J2_127_3477_n1082) );
  FADDX1_HVT DP_OP_425J2_127_3477_U637 ( .A(DP_OP_425J2_127_3477_n1102), .B(
        DP_OP_425J2_127_3477_n1098), .CI(DP_OP_425J2_127_3477_n1096), .CO(
        DP_OP_425J2_127_3477_n1079), .S(DP_OP_425J2_127_3477_n1080) );
  FADDX1_HVT DP_OP_425J2_127_3477_U636 ( .A(DP_OP_425J2_127_3477_n1269), .B(
        DP_OP_425J2_127_3477_n1094), .CI(DP_OP_425J2_127_3477_n1092), .CO(
        DP_OP_425J2_127_3477_n1077), .S(DP_OP_425J2_127_3477_n1078) );
  FADDX1_HVT DP_OP_425J2_127_3477_U635 ( .A(DP_OP_425J2_127_3477_n1267), .B(
        DP_OP_425J2_127_3477_n1090), .CI(DP_OP_425J2_127_3477_n1088), .CO(
        DP_OP_425J2_127_3477_n1075), .S(DP_OP_425J2_127_3477_n1076) );
  FADDX1_HVT DP_OP_425J2_127_3477_U634 ( .A(DP_OP_425J2_127_3477_n1265), .B(
        DP_OP_425J2_127_3477_n1263), .CI(DP_OP_425J2_127_3477_n1086), .CO(
        DP_OP_425J2_127_3477_n1073), .S(DP_OP_425J2_127_3477_n1074) );
  FADDX1_HVT DP_OP_425J2_127_3477_U633 ( .A(DP_OP_425J2_127_3477_n1084), .B(
        DP_OP_425J2_127_3477_n1261), .CI(DP_OP_425J2_127_3477_n1082), .CO(
        DP_OP_425J2_127_3477_n1071), .S(DP_OP_425J2_127_3477_n1072) );
  FADDX1_HVT DP_OP_425J2_127_3477_U632 ( .A(DP_OP_425J2_127_3477_n1259), .B(
        DP_OP_425J2_127_3477_n1080), .CI(DP_OP_425J2_127_3477_n1078), .CO(
        DP_OP_425J2_127_3477_n1069), .S(DP_OP_425J2_127_3477_n1070) );
  FADDX1_HVT DP_OP_425J2_127_3477_U631 ( .A(DP_OP_425J2_127_3477_n1257), .B(
        DP_OP_425J2_127_3477_n1076), .CI(DP_OP_425J2_127_3477_n1255), .CO(
        DP_OP_425J2_127_3477_n1067), .S(DP_OP_425J2_127_3477_n1068) );
  FADDX1_HVT DP_OP_425J2_127_3477_U630 ( .A(DP_OP_425J2_127_3477_n1074), .B(
        DP_OP_425J2_127_3477_n1072), .CI(DP_OP_425J2_127_3477_n1253), .CO(
        DP_OP_425J2_127_3477_n1065), .S(DP_OP_425J2_127_3477_n1066) );
  FADDX1_HVT DP_OP_425J2_127_3477_U629 ( .A(DP_OP_425J2_127_3477_n1070), .B(
        DP_OP_425J2_127_3477_n1251), .CI(DP_OP_425J2_127_3477_n1068), .CO(
        DP_OP_425J2_127_3477_n1063), .S(DP_OP_425J2_127_3477_n1064) );
  OR2X1_HVT DP_OP_425J2_127_3477_U628 ( .A1(DP_OP_425J2_127_3477_n2352), .A2(
        DP_OP_425J2_127_3477_n2703), .Y(DP_OP_425J2_127_3477_n1061) );
  FADDX1_HVT DP_OP_425J2_127_3477_U626 ( .A(DP_OP_425J2_127_3477_n2002), .B(
        DP_OP_425J2_127_3477_n1826), .CI(DP_OP_425J2_127_3477_n2395), .CO(
        DP_OP_425J2_127_3477_n1059), .S(DP_OP_425J2_127_3477_n1060) );
  FADDX1_HVT DP_OP_425J2_127_3477_U625 ( .A(DP_OP_425J2_127_3477_n2659), .B(
        DP_OP_425J2_127_3477_n2046), .CI(DP_OP_425J2_127_3477_n2747), .CO(
        DP_OP_425J2_127_3477_n1057), .S(DP_OP_425J2_127_3477_n1058) );
  FADDX1_HVT DP_OP_425J2_127_3477_U624 ( .A(DP_OP_425J2_127_3477_n2310), .B(
        DP_OP_425J2_127_3477_n2527), .CI(DP_OP_425J2_127_3477_n1958), .CO(
        DP_OP_425J2_127_3477_n1055), .S(DP_OP_425J2_127_3477_n1056) );
  FADDX1_HVT DP_OP_425J2_127_3477_U623 ( .A(DP_OP_425J2_127_3477_n2791), .B(
        DP_OP_425J2_127_3477_n2483), .CI(DP_OP_425J2_127_3477_n2178), .CO(
        DP_OP_425J2_127_3477_n1053), .S(DP_OP_425J2_127_3477_n1054) );
  FADDX1_HVT DP_OP_425J2_127_3477_U622 ( .A(DP_OP_425J2_127_3477_n1870), .B(
        DP_OP_425J2_127_3477_n1914), .CI(DP_OP_425J2_127_3477_n2571), .CO(
        DP_OP_425J2_127_3477_n1051), .S(DP_OP_425J2_127_3477_n1052) );
  FADDX1_HVT DP_OP_425J2_127_3477_U621 ( .A(DP_OP_425J2_127_3477_n2090), .B(
        DP_OP_425J2_127_3477_n2879), .CI(DP_OP_425J2_127_3477_n2439), .CO(
        DP_OP_425J2_127_3477_n1049), .S(DP_OP_425J2_127_3477_n1050) );
  FADDX1_HVT DP_OP_425J2_127_3477_U620 ( .A(DP_OP_425J2_127_3477_n2615), .B(
        DP_OP_425J2_127_3477_n2134), .CI(DP_OP_425J2_127_3477_n2266), .CO(
        DP_OP_425J2_127_3477_n1047), .S(DP_OP_425J2_127_3477_n1048) );
  FADDX1_HVT DP_OP_425J2_127_3477_U619 ( .A(DP_OP_425J2_127_3477_n2835), .B(
        DP_OP_425J2_127_3477_n2222), .CI(DP_OP_425J2_127_3477_n2111), .CO(
        DP_OP_425J2_127_3477_n1045), .S(DP_OP_425J2_127_3477_n1046) );
  FADDX1_HVT DP_OP_425J2_127_3477_U618 ( .A(DP_OP_425J2_127_3477_n2636), .B(
        DP_OP_425J2_127_3477_n2578), .CI(DP_OP_425J2_127_3477_n2287), .CO(
        DP_OP_425J2_127_3477_n1043), .S(DP_OP_425J2_127_3477_n1044) );
  FADDX1_HVT DP_OP_425J2_127_3477_U617 ( .A(DP_OP_425J2_127_3477_n2416), .B(
        DP_OP_425J2_127_3477_n2724), .CI(DP_OP_425J2_127_3477_n2067), .CO(
        DP_OP_425J2_127_3477_n1041), .S(DP_OP_425J2_127_3477_n1042) );
  FADDX1_HVT DP_OP_425J2_127_3477_U616 ( .A(DP_OP_425J2_127_3477_n2548), .B(
        DP_OP_425J2_127_3477_n1965), .CI(DP_OP_425J2_127_3477_n2273), .CO(
        DP_OP_425J2_127_3477_n1039), .S(DP_OP_425J2_127_3477_n1040) );
  FADDX1_HVT DP_OP_425J2_127_3477_U615 ( .A(DP_OP_425J2_127_3477_n2331), .B(
        DP_OP_425J2_127_3477_n2534), .CI(DP_OP_425J2_127_3477_n2141), .CO(
        DP_OP_425J2_127_3477_n1037), .S(DP_OP_425J2_127_3477_n1038) );
  FADDX1_HVT DP_OP_425J2_127_3477_U614 ( .A(DP_OP_425J2_127_3477_n2199), .B(
        DP_OP_425J2_127_3477_n2409), .CI(DP_OP_425J2_127_3477_n2805), .CO(
        DP_OP_425J2_127_3477_n1035), .S(DP_OP_425J2_127_3477_n1036) );
  FADDX1_HVT DP_OP_425J2_127_3477_U613 ( .A(DP_OP_425J2_127_3477_n2460), .B(
        DP_OP_425J2_127_3477_n2148), .CI(DP_OP_425J2_127_3477_n2280), .CO(
        DP_OP_425J2_127_3477_n1033), .S(DP_OP_425J2_127_3477_n1034) );
  FADDX1_HVT DP_OP_425J2_127_3477_U612 ( .A(DP_OP_425J2_127_3477_n2592), .B(
        DP_OP_425J2_127_3477_n1782), .CI(DP_OP_425J2_127_3477_n2317), .CO(
        DP_OP_425J2_127_3477_n1031), .S(DP_OP_425J2_127_3477_n1032) );
  FADDX1_HVT DP_OP_425J2_127_3477_U611 ( .A(DP_OP_425J2_127_3477_n1847), .B(
        DP_OP_425J2_127_3477_n2680), .CI(DP_OP_425J2_127_3477_n2053), .CO(
        DP_OP_425J2_127_3477_n1029), .S(DP_OP_425J2_127_3477_n1030) );
  FADDX1_HVT DP_OP_425J2_127_3477_U610 ( .A(DP_OP_425J2_127_3477_n2886), .B(
        DP_OP_425J2_127_3477_n2324), .CI(DP_OP_425J2_127_3477_n2893), .CO(
        DP_OP_425J2_127_3477_n1027), .S(DP_OP_425J2_127_3477_n1028) );
  FADDX1_HVT DP_OP_425J2_127_3477_U609 ( .A(DP_OP_425J2_127_3477_n2842), .B(
        DP_OP_425J2_127_3477_n2585), .CI(DP_OP_425J2_127_3477_n2849), .CO(
        DP_OP_425J2_127_3477_n1025), .S(DP_OP_425J2_127_3477_n1026) );
  FADDX1_HVT DP_OP_425J2_127_3477_U608 ( .A(DP_OP_425J2_127_3477_n2060), .B(
        DP_OP_425J2_127_3477_n2497), .CI(DP_OP_425J2_127_3477_n2541), .CO(
        DP_OP_425J2_127_3477_n1023), .S(DP_OP_425J2_127_3477_n1024) );
  FADDX1_HVT DP_OP_425J2_127_3477_U607 ( .A(DP_OP_425J2_127_3477_n2629), .B(
        DP_OP_425J2_127_3477_n1979), .CI(DP_OP_425J2_127_3477_n2710), .CO(
        DP_OP_425J2_127_3477_n1021), .S(DP_OP_425J2_127_3477_n1022) );
  FADDX1_HVT DP_OP_425J2_127_3477_U606 ( .A(DP_OP_425J2_127_3477_n2023), .B(
        DP_OP_425J2_127_3477_n2754), .CI(DP_OP_425J2_127_3477_n1935), .CO(
        DP_OP_425J2_127_3477_n1019), .S(DP_OP_425J2_127_3477_n1020) );
  FADDX1_HVT DP_OP_425J2_127_3477_U605 ( .A(DP_OP_425J2_127_3477_n1840), .B(
        DP_OP_425J2_127_3477_n2856), .CI(DP_OP_425J2_127_3477_n2504), .CO(
        DP_OP_425J2_127_3477_n1017), .S(DP_OP_425J2_127_3477_n1018) );
  FADDX1_HVT DP_OP_425J2_127_3477_U604 ( .A(DP_OP_425J2_127_3477_n2229), .B(
        DP_OP_425J2_127_3477_n2446), .CI(DP_OP_425J2_127_3477_n2185), .CO(
        DP_OP_425J2_127_3477_n1015), .S(DP_OP_425J2_127_3477_n1016) );
  FADDX1_HVT DP_OP_425J2_127_3477_U603 ( .A(DP_OP_425J2_127_3477_n2768), .B(
        DP_OP_425J2_127_3477_n1891), .CI(DP_OP_425J2_127_3477_n1921), .CO(
        DP_OP_425J2_127_3477_n1013), .S(DP_OP_425J2_127_3477_n1014) );
  FADDX1_HVT DP_OP_425J2_127_3477_U602 ( .A(DP_OP_425J2_127_3477_n2097), .B(
        DP_OP_425J2_127_3477_n2666), .CI(DP_OP_425J2_127_3477_n1877), .CO(
        DP_OP_425J2_127_3477_n1011), .S(DP_OP_425J2_127_3477_n1012) );
  FADDX1_HVT DP_OP_425J2_127_3477_U601 ( .A(DP_OP_425J2_127_3477_n2761), .B(
        DP_OP_425J2_127_3477_n2453), .CI(DP_OP_425J2_127_3477_n2009), .CO(
        DP_OP_425J2_127_3477_n1009), .S(DP_OP_425J2_127_3477_n1010) );
  FADDX1_HVT DP_OP_425J2_127_3477_U600 ( .A(DP_OP_425J2_127_3477_n1884), .B(
        DP_OP_425J2_127_3477_n1833), .CI(DP_OP_425J2_127_3477_n2365), .CO(
        DP_OP_425J2_127_3477_n1007), .S(DP_OP_425J2_127_3477_n1008) );
  FADDX1_HVT DP_OP_425J2_127_3477_U599 ( .A(DP_OP_425J2_127_3477_n2490), .B(
        DP_OP_425J2_127_3477_n2798), .CI(DP_OP_425J2_127_3477_n2192), .CO(
        DP_OP_425J2_127_3477_n1005), .S(DP_OP_425J2_127_3477_n1006) );
  FADDX1_HVT DP_OP_425J2_127_3477_U598 ( .A(DP_OP_425J2_127_3477_n2104), .B(
        DP_OP_425J2_127_3477_n2622), .CI(DP_OP_425J2_127_3477_n2236), .CO(
        DP_OP_425J2_127_3477_n1003), .S(DP_OP_425J2_127_3477_n1004) );
  FADDX1_HVT DP_OP_425J2_127_3477_U597 ( .A(DP_OP_425J2_127_3477_n2673), .B(
        DP_OP_425J2_127_3477_n1972), .CI(DP_OP_425J2_127_3477_n1928), .CO(
        DP_OP_425J2_127_3477_n1001), .S(DP_OP_425J2_127_3477_n1002) );
  FADDX1_HVT DP_OP_425J2_127_3477_U596 ( .A(DP_OP_425J2_127_3477_n2358), .B(
        DP_OP_425J2_127_3477_n2243), .CI(DP_OP_425J2_127_3477_n2155), .CO(
        DP_OP_425J2_127_3477_n999), .S(DP_OP_425J2_127_3477_n1000) );
  FADDX1_HVT DP_OP_425J2_127_3477_U595 ( .A(DP_OP_425J2_127_3477_n2900), .B(
        DP_OP_425J2_127_3477_n2016), .CI(DP_OP_425J2_127_3477_n2812), .CO(
        DP_OP_425J2_127_3477_n997), .S(DP_OP_425J2_127_3477_n998) );
  FADDX1_HVT DP_OP_425J2_127_3477_U594 ( .A(DP_OP_425J2_127_3477_n2372), .B(
        DP_OP_425J2_127_3477_n2402), .CI(DP_OP_425J2_127_3477_n1249), .CO(
        DP_OP_425J2_127_3477_n995), .S(DP_OP_425J2_127_3477_n996) );
  FADDX1_HVT DP_OP_425J2_127_3477_U593 ( .A(DP_OP_425J2_127_3477_n2717), .B(
        DP_OP_425J2_127_3477_n1247), .CI(DP_OP_425J2_127_3477_n1245), .CO(
        DP_OP_425J2_127_3477_n993), .S(DP_OP_425J2_127_3477_n994) );
  FADDX1_HVT DP_OP_425J2_127_3477_U592 ( .A(DP_OP_425J2_127_3477_n1235), .B(
        DP_OP_425J2_127_3477_n1062), .CI(DP_OP_425J2_127_3477_n1233), .CO(
        DP_OP_425J2_127_3477_n991), .S(DP_OP_425J2_127_3477_n992) );
  FADDX1_HVT DP_OP_425J2_127_3477_U591 ( .A(DP_OP_425J2_127_3477_n1243), .B(
        DP_OP_425J2_127_3477_n1237), .CI(DP_OP_425J2_127_3477_n1239), .CO(
        DP_OP_425J2_127_3477_n989), .S(DP_OP_425J2_127_3477_n990) );
  FADDX1_HVT DP_OP_425J2_127_3477_U590 ( .A(DP_OP_425J2_127_3477_n1241), .B(
        DP_OP_425J2_127_3477_n1231), .CI(DP_OP_425J2_127_3477_n1229), .CO(
        DP_OP_425J2_127_3477_n987), .S(DP_OP_425J2_127_3477_n988) );
  FADDX1_HVT DP_OP_425J2_127_3477_U589 ( .A(DP_OP_425J2_127_3477_n1227), .B(
        DP_OP_425J2_127_3477_n1205), .CI(DP_OP_425J2_127_3477_n1199), .CO(
        DP_OP_425J2_127_3477_n985), .S(DP_OP_425J2_127_3477_n986) );
  FADDX1_HVT DP_OP_425J2_127_3477_U588 ( .A(DP_OP_425J2_127_3477_n1225), .B(
        DP_OP_425J2_127_3477_n1207), .CI(DP_OP_425J2_127_3477_n1201), .CO(
        DP_OP_425J2_127_3477_n983), .S(DP_OP_425J2_127_3477_n984) );
  FADDX1_HVT DP_OP_425J2_127_3477_U587 ( .A(DP_OP_425J2_127_3477_n1223), .B(
        DP_OP_425J2_127_3477_n1209), .CI(DP_OP_425J2_127_3477_n1203), .CO(
        DP_OP_425J2_127_3477_n981), .S(DP_OP_425J2_127_3477_n982) );
  FADDX1_HVT DP_OP_425J2_127_3477_U586 ( .A(DP_OP_425J2_127_3477_n1213), .B(
        DP_OP_425J2_127_3477_n1221), .CI(DP_OP_425J2_127_3477_n1211), .CO(
        DP_OP_425J2_127_3477_n979), .S(DP_OP_425J2_127_3477_n980) );
  FADDX1_HVT DP_OP_425J2_127_3477_U585 ( .A(DP_OP_425J2_127_3477_n1217), .B(
        DP_OP_425J2_127_3477_n1215), .CI(DP_OP_425J2_127_3477_n1219), .CO(
        DP_OP_425J2_127_3477_n977), .S(DP_OP_425J2_127_3477_n978) );
  FADDX1_HVT DP_OP_425J2_127_3477_U584 ( .A(DP_OP_425J2_127_3477_n1197), .B(
        DP_OP_425J2_127_3477_n1050), .CI(DP_OP_425J2_127_3477_n1185), .CO(
        DP_OP_425J2_127_3477_n975), .S(DP_OP_425J2_127_3477_n976) );
  FADDX1_HVT DP_OP_425J2_127_3477_U583 ( .A(DP_OP_425J2_127_3477_n1193), .B(
        DP_OP_425J2_127_3477_n1056), .CI(DP_OP_425J2_127_3477_n1183), .CO(
        DP_OP_425J2_127_3477_n973), .S(DP_OP_425J2_127_3477_n974) );
  FADDX1_HVT DP_OP_425J2_127_3477_U582 ( .A(DP_OP_425J2_127_3477_n1195), .B(
        DP_OP_425J2_127_3477_n1052), .CI(DP_OP_425J2_127_3477_n1054), .CO(
        DP_OP_425J2_127_3477_n971), .S(DP_OP_425J2_127_3477_n972) );
  FADDX1_HVT DP_OP_425J2_127_3477_U581 ( .A(DP_OP_425J2_127_3477_n1191), .B(
        DP_OP_425J2_127_3477_n1048), .CI(DP_OP_425J2_127_3477_n1058), .CO(
        DP_OP_425J2_127_3477_n969), .S(DP_OP_425J2_127_3477_n970) );
  FADDX1_HVT DP_OP_425J2_127_3477_U580 ( .A(DP_OP_425J2_127_3477_n1189), .B(
        DP_OP_425J2_127_3477_n1187), .CI(DP_OP_425J2_127_3477_n1060), .CO(
        DP_OP_425J2_127_3477_n967), .S(DP_OP_425J2_127_3477_n968) );
  FADDX1_HVT DP_OP_425J2_127_3477_U579 ( .A(DP_OP_425J2_127_3477_n1046), .B(
        DP_OP_425J2_127_3477_n1038), .CI(DP_OP_425J2_127_3477_n1018), .CO(
        DP_OP_425J2_127_3477_n965), .S(DP_OP_425J2_127_3477_n966) );
  FADDX1_HVT DP_OP_425J2_127_3477_U578 ( .A(DP_OP_425J2_127_3477_n1034), .B(
        DP_OP_425J2_127_3477_n1020), .CI(DP_OP_425J2_127_3477_n1012), .CO(
        DP_OP_425J2_127_3477_n963), .S(DP_OP_425J2_127_3477_n964) );
  FADDX1_HVT DP_OP_425J2_127_3477_U577 ( .A(DP_OP_425J2_127_3477_n1036), .B(
        DP_OP_425J2_127_3477_n1022), .CI(DP_OP_425J2_127_3477_n1016), .CO(
        DP_OP_425J2_127_3477_n961), .S(DP_OP_425J2_127_3477_n962) );
  FADDX1_HVT DP_OP_425J2_127_3477_U576 ( .A(DP_OP_425J2_127_3477_n1030), .B(
        DP_OP_425J2_127_3477_n1024), .CI(DP_OP_425J2_127_3477_n1014), .CO(
        DP_OP_425J2_127_3477_n959), .S(DP_OP_425J2_127_3477_n960) );
  FADDX1_HVT DP_OP_425J2_127_3477_U575 ( .A(DP_OP_425J2_127_3477_n1032), .B(
        DP_OP_425J2_127_3477_n1044), .CI(DP_OP_425J2_127_3477_n1042), .CO(
        DP_OP_425J2_127_3477_n957), .S(DP_OP_425J2_127_3477_n958) );
  FADDX1_HVT DP_OP_425J2_127_3477_U574 ( .A(DP_OP_425J2_127_3477_n1026), .B(
        DP_OP_425J2_127_3477_n1040), .CI(DP_OP_425J2_127_3477_n1028), .CO(
        DP_OP_425J2_127_3477_n955), .S(DP_OP_425J2_127_3477_n956) );
  FADDX1_HVT DP_OP_425J2_127_3477_U573 ( .A(DP_OP_425J2_127_3477_n1010), .B(
        DP_OP_425J2_127_3477_n1000), .CI(DP_OP_425J2_127_3477_n998), .CO(
        DP_OP_425J2_127_3477_n953), .S(DP_OP_425J2_127_3477_n954) );
  FADDX1_HVT DP_OP_425J2_127_3477_U572 ( .A(DP_OP_425J2_127_3477_n1006), .B(
        DP_OP_425J2_127_3477_n1002), .CI(DP_OP_425J2_127_3477_n1181), .CO(
        DP_OP_425J2_127_3477_n951), .S(DP_OP_425J2_127_3477_n952) );
  FADDX1_HVT DP_OP_425J2_127_3477_U571 ( .A(DP_OP_425J2_127_3477_n1004), .B(
        DP_OP_425J2_127_3477_n1008), .CI(DP_OP_425J2_127_3477_n996), .CO(
        DP_OP_425J2_127_3477_n949), .S(DP_OP_425J2_127_3477_n950) );
  FADDX1_HVT DP_OP_425J2_127_3477_U570 ( .A(DP_OP_425J2_127_3477_n1179), .B(
        DP_OP_425J2_127_3477_n1177), .CI(DP_OP_425J2_127_3477_n1175), .CO(
        DP_OP_425J2_127_3477_n947), .S(DP_OP_425J2_127_3477_n948) );
  FADDX1_HVT DP_OP_425J2_127_3477_U569 ( .A(DP_OP_425J2_127_3477_n1173), .B(
        DP_OP_425J2_127_3477_n1165), .CI(DP_OP_425J2_127_3477_n1167), .CO(
        DP_OP_425J2_127_3477_n945), .S(DP_OP_425J2_127_3477_n946) );
  FADDX1_HVT DP_OP_425J2_127_3477_U568 ( .A(DP_OP_425J2_127_3477_n1169), .B(
        DP_OP_425J2_127_3477_n1171), .CI(DP_OP_425J2_127_3477_n994), .CO(
        DP_OP_425J2_127_3477_n943), .S(DP_OP_425J2_127_3477_n944) );
  FADDX1_HVT DP_OP_425J2_127_3477_U567 ( .A(DP_OP_425J2_127_3477_n1163), .B(
        DP_OP_425J2_127_3477_n992), .CI(DP_OP_425J2_127_3477_n990), .CO(
        DP_OP_425J2_127_3477_n941), .S(DP_OP_425J2_127_3477_n942) );
  FADDX1_HVT DP_OP_425J2_127_3477_U566 ( .A(DP_OP_425J2_127_3477_n1157), .B(
        DP_OP_425J2_127_3477_n1159), .CI(DP_OP_425J2_127_3477_n1155), .CO(
        DP_OP_425J2_127_3477_n939), .S(DP_OP_425J2_127_3477_n940) );
  FADDX1_HVT DP_OP_425J2_127_3477_U565 ( .A(DP_OP_425J2_127_3477_n1161), .B(
        DP_OP_425J2_127_3477_n1153), .CI(DP_OP_425J2_127_3477_n988), .CO(
        DP_OP_425J2_127_3477_n937), .S(DP_OP_425J2_127_3477_n938) );
  FADDX1_HVT DP_OP_425J2_127_3477_U564 ( .A(DP_OP_425J2_127_3477_n1151), .B(
        DP_OP_425J2_127_3477_n1149), .CI(DP_OP_425J2_127_3477_n984), .CO(
        DP_OP_425J2_127_3477_n935), .S(DP_OP_425J2_127_3477_n936) );
  FADDX1_HVT DP_OP_425J2_127_3477_U563 ( .A(DP_OP_425J2_127_3477_n980), .B(
        DP_OP_425J2_127_3477_n978), .CI(DP_OP_425J2_127_3477_n986), .CO(
        DP_OP_425J2_127_3477_n933), .S(DP_OP_425J2_127_3477_n934) );
  FADDX1_HVT DP_OP_425J2_127_3477_U562 ( .A(DP_OP_425J2_127_3477_n1147), .B(
        DP_OP_425J2_127_3477_n982), .CI(DP_OP_425J2_127_3477_n1143), .CO(
        DP_OP_425J2_127_3477_n931), .S(DP_OP_425J2_127_3477_n932) );
  FADDX1_HVT DP_OP_425J2_127_3477_U561 ( .A(DP_OP_425J2_127_3477_n1145), .B(
        DP_OP_425J2_127_3477_n1141), .CI(DP_OP_425J2_127_3477_n976), .CO(
        DP_OP_425J2_127_3477_n929), .S(DP_OP_425J2_127_3477_n930) );
  FADDX1_HVT DP_OP_425J2_127_3477_U560 ( .A(DP_OP_425J2_127_3477_n1139), .B(
        DP_OP_425J2_127_3477_n968), .CI(DP_OP_425J2_127_3477_n1137), .CO(
        DP_OP_425J2_127_3477_n927), .S(DP_OP_425J2_127_3477_n928) );
  FADDX1_HVT DP_OP_425J2_127_3477_U559 ( .A(DP_OP_425J2_127_3477_n970), .B(
        DP_OP_425J2_127_3477_n974), .CI(DP_OP_425J2_127_3477_n972), .CO(
        DP_OP_425J2_127_3477_n925), .S(DP_OP_425J2_127_3477_n926) );
  FADDX1_HVT DP_OP_425J2_127_3477_U558 ( .A(DP_OP_425J2_127_3477_n966), .B(
        DP_OP_425J2_127_3477_n962), .CI(DP_OP_425J2_127_3477_n1135), .CO(
        DP_OP_425J2_127_3477_n923), .S(DP_OP_425J2_127_3477_n924) );
  FADDX1_HVT DP_OP_425J2_127_3477_U557 ( .A(DP_OP_425J2_127_3477_n958), .B(
        DP_OP_425J2_127_3477_n964), .CI(DP_OP_425J2_127_3477_n956), .CO(
        DP_OP_425J2_127_3477_n921), .S(DP_OP_425J2_127_3477_n922) );
  FADDX1_HVT DP_OP_425J2_127_3477_U556 ( .A(DP_OP_425J2_127_3477_n960), .B(
        DP_OP_425J2_127_3477_n954), .CI(DP_OP_425J2_127_3477_n950), .CO(
        DP_OP_425J2_127_3477_n919), .S(DP_OP_425J2_127_3477_n920) );
  FADDX1_HVT DP_OP_425J2_127_3477_U555 ( .A(DP_OP_425J2_127_3477_n952), .B(
        DP_OP_425J2_127_3477_n1131), .CI(DP_OP_425J2_127_3477_n1133), .CO(
        DP_OP_425J2_127_3477_n917), .S(DP_OP_425J2_127_3477_n918) );
  FADDX1_HVT DP_OP_425J2_127_3477_U554 ( .A(DP_OP_425J2_127_3477_n1129), .B(
        DP_OP_425J2_127_3477_n948), .CI(DP_OP_425J2_127_3477_n1125), .CO(
        DP_OP_425J2_127_3477_n915), .S(DP_OP_425J2_127_3477_n916) );
  FADDX1_HVT DP_OP_425J2_127_3477_U553 ( .A(DP_OP_425J2_127_3477_n1127), .B(
        DP_OP_425J2_127_3477_n1123), .CI(DP_OP_425J2_127_3477_n1121), .CO(
        DP_OP_425J2_127_3477_n913), .S(DP_OP_425J2_127_3477_n914) );
  FADDX1_HVT DP_OP_425J2_127_3477_U552 ( .A(DP_OP_425J2_127_3477_n1119), .B(
        DP_OP_425J2_127_3477_n944), .CI(DP_OP_425J2_127_3477_n1117), .CO(
        DP_OP_425J2_127_3477_n911), .S(DP_OP_425J2_127_3477_n912) );
  FADDX1_HVT DP_OP_425J2_127_3477_U551 ( .A(DP_OP_425J2_127_3477_n946), .B(
        DP_OP_425J2_127_3477_n942), .CI(DP_OP_425J2_127_3477_n1115), .CO(
        DP_OP_425J2_127_3477_n909), .S(DP_OP_425J2_127_3477_n910) );
  FADDX1_HVT DP_OP_425J2_127_3477_U550 ( .A(DP_OP_425J2_127_3477_n1113), .B(
        DP_OP_425J2_127_3477_n940), .CI(DP_OP_425J2_127_3477_n938), .CO(
        DP_OP_425J2_127_3477_n907), .S(DP_OP_425J2_127_3477_n908) );
  FADDX1_HVT DP_OP_425J2_127_3477_U549 ( .A(DP_OP_425J2_127_3477_n1109), .B(
        DP_OP_425J2_127_3477_n932), .CI(DP_OP_425J2_127_3477_n930), .CO(
        DP_OP_425J2_127_3477_n905), .S(DP_OP_425J2_127_3477_n906) );
  FADDX1_HVT DP_OP_425J2_127_3477_U548 ( .A(DP_OP_425J2_127_3477_n1111), .B(
        DP_OP_425J2_127_3477_n936), .CI(DP_OP_425J2_127_3477_n934), .CO(
        DP_OP_425J2_127_3477_n903), .S(DP_OP_425J2_127_3477_n904) );
  FADDX1_HVT DP_OP_425J2_127_3477_U547 ( .A(DP_OP_425J2_127_3477_n1107), .B(
        DP_OP_425J2_127_3477_n926), .CI(DP_OP_425J2_127_3477_n1105), .CO(
        DP_OP_425J2_127_3477_n901), .S(DP_OP_425J2_127_3477_n902) );
  FADDX1_HVT DP_OP_425J2_127_3477_U546 ( .A(DP_OP_425J2_127_3477_n928), .B(
        DP_OP_425J2_127_3477_n924), .CI(DP_OP_425J2_127_3477_n1103), .CO(
        DP_OP_425J2_127_3477_n899), .S(DP_OP_425J2_127_3477_n900) );
  FADDX1_HVT DP_OP_425J2_127_3477_U545 ( .A(DP_OP_425J2_127_3477_n922), .B(
        DP_OP_425J2_127_3477_n920), .CI(DP_OP_425J2_127_3477_n918), .CO(
        DP_OP_425J2_127_3477_n897), .S(DP_OP_425J2_127_3477_n898) );
  FADDX1_HVT DP_OP_425J2_127_3477_U544 ( .A(DP_OP_425J2_127_3477_n1101), .B(
        DP_OP_425J2_127_3477_n1099), .CI(DP_OP_425J2_127_3477_n1097), .CO(
        DP_OP_425J2_127_3477_n895), .S(DP_OP_425J2_127_3477_n896) );
  FADDX1_HVT DP_OP_425J2_127_3477_U543 ( .A(DP_OP_425J2_127_3477_n916), .B(
        DP_OP_425J2_127_3477_n1095), .CI(DP_OP_425J2_127_3477_n914), .CO(
        DP_OP_425J2_127_3477_n893), .S(DP_OP_425J2_127_3477_n894) );
  FADDX1_HVT DP_OP_425J2_127_3477_U542 ( .A(DP_OP_425J2_127_3477_n1093), .B(
        DP_OP_425J2_127_3477_n1091), .CI(DP_OP_425J2_127_3477_n910), .CO(
        DP_OP_425J2_127_3477_n891), .S(DP_OP_425J2_127_3477_n892) );
  FADDX1_HVT DP_OP_425J2_127_3477_U541 ( .A(DP_OP_425J2_127_3477_n912), .B(
        DP_OP_425J2_127_3477_n908), .CI(DP_OP_425J2_127_3477_n1089), .CO(
        DP_OP_425J2_127_3477_n889), .S(DP_OP_425J2_127_3477_n890) );
  FADDX1_HVT DP_OP_425J2_127_3477_U540 ( .A(DP_OP_425J2_127_3477_n1087), .B(
        DP_OP_425J2_127_3477_n906), .CI(DP_OP_425J2_127_3477_n904), .CO(
        DP_OP_425J2_127_3477_n887), .S(DP_OP_425J2_127_3477_n888) );
  FADDX1_HVT DP_OP_425J2_127_3477_U539 ( .A(DP_OP_425J2_127_3477_n902), .B(
        DP_OP_425J2_127_3477_n1085), .CI(DP_OP_425J2_127_3477_n900), .CO(
        DP_OP_425J2_127_3477_n885), .S(DP_OP_425J2_127_3477_n886) );
  FADDX1_HVT DP_OP_425J2_127_3477_U538 ( .A(DP_OP_425J2_127_3477_n1083), .B(
        DP_OP_425J2_127_3477_n898), .CI(DP_OP_425J2_127_3477_n1081), .CO(
        DP_OP_425J2_127_3477_n883), .S(DP_OP_425J2_127_3477_n884) );
  FADDX1_HVT DP_OP_425J2_127_3477_U537 ( .A(DP_OP_425J2_127_3477_n896), .B(
        DP_OP_425J2_127_3477_n1079), .CI(DP_OP_425J2_127_3477_n894), .CO(
        DP_OP_425J2_127_3477_n881), .S(DP_OP_425J2_127_3477_n882) );
  FADDX1_HVT DP_OP_425J2_127_3477_U536 ( .A(DP_OP_425J2_127_3477_n1077), .B(
        DP_OP_425J2_127_3477_n892), .CI(DP_OP_425J2_127_3477_n890), .CO(
        DP_OP_425J2_127_3477_n879), .S(DP_OP_425J2_127_3477_n880) );
  FADDX1_HVT DP_OP_425J2_127_3477_U535 ( .A(DP_OP_425J2_127_3477_n1075), .B(
        DP_OP_425J2_127_3477_n888), .CI(DP_OP_425J2_127_3477_n1073), .CO(
        DP_OP_425J2_127_3477_n877), .S(DP_OP_425J2_127_3477_n878) );
  FADDX1_HVT DP_OP_425J2_127_3477_U534 ( .A(DP_OP_425J2_127_3477_n886), .B(
        DP_OP_425J2_127_3477_n1071), .CI(DP_OP_425J2_127_3477_n884), .CO(
        DP_OP_425J2_127_3477_n875), .S(DP_OP_425J2_127_3477_n876) );
  FADDX1_HVT DP_OP_425J2_127_3477_U533 ( .A(DP_OP_425J2_127_3477_n882), .B(
        DP_OP_425J2_127_3477_n1069), .CI(DP_OP_425J2_127_3477_n880), .CO(
        DP_OP_425J2_127_3477_n873), .S(DP_OP_425J2_127_3477_n874) );
  FADDX1_HVT DP_OP_425J2_127_3477_U532 ( .A(DP_OP_425J2_127_3477_n1067), .B(
        DP_OP_425J2_127_3477_n878), .CI(DP_OP_425J2_127_3477_n876), .CO(
        DP_OP_425J2_127_3477_n871), .S(DP_OP_425J2_127_3477_n872) );
  FADDX1_HVT DP_OP_425J2_127_3477_U531 ( .A(DP_OP_425J2_127_3477_n1065), .B(
        DP_OP_425J2_127_3477_n874), .CI(DP_OP_425J2_127_3477_n1063), .CO(
        DP_OP_425J2_127_3477_n869), .S(DP_OP_425J2_127_3477_n870) );
  FADDX1_HVT DP_OP_425J2_127_3477_U530 ( .A(DP_OP_425J2_127_3477_n2351), .B(
        DP_OP_425J2_127_3477_n1825), .CI(DP_OP_425J2_127_3477_n1934), .CO(
        DP_OP_425J2_127_3477_n867), .S(DP_OP_425J2_127_3477_n868) );
  FADDX1_HVT DP_OP_425J2_127_3477_U529 ( .A(DP_OP_425J2_127_3477_n2001), .B(
        DP_OP_425J2_127_3477_n2723), .CI(DP_OP_425J2_127_3477_n1890), .CO(
        DP_OP_425J2_127_3477_n865), .S(DP_OP_425J2_127_3477_n866) );
  FADDX1_HVT DP_OP_425J2_127_3477_U528 ( .A(DP_OP_425J2_127_3477_n2702), .B(
        DP_OP_425J2_127_3477_n2526), .CI(DP_OP_425J2_127_3477_n2503), .CO(
        DP_OP_425J2_127_3477_n863), .S(DP_OP_425J2_127_3477_n864) );
  FADDX1_HVT DP_OP_425J2_127_3477_U527 ( .A(DP_OP_425J2_127_3477_n2089), .B(
        DP_OP_425J2_127_3477_n2482), .CI(DP_OP_425J2_127_3477_n2855), .CO(
        DP_OP_425J2_127_3477_n861), .S(DP_OP_425J2_127_3477_n862) );
  FADDX1_HVT DP_OP_425J2_127_3477_U526 ( .A(DP_OP_425J2_127_3477_n1869), .B(
        DP_OP_425J2_127_3477_n2045), .CI(DP_OP_425J2_127_3477_n2767), .CO(
        DP_OP_425J2_127_3477_n859), .S(DP_OP_425J2_127_3477_n860) );
  FADDX1_HVT DP_OP_425J2_127_3477_U525 ( .A(DP_OP_425J2_127_3477_n2658), .B(
        DP_OP_425J2_127_3477_n2438), .CI(DP_OP_425J2_127_3477_n2394), .CO(
        DP_OP_425J2_127_3477_n857), .S(DP_OP_425J2_127_3477_n858) );
  FADDX1_HVT DP_OP_425J2_127_3477_U524 ( .A(DP_OP_425J2_127_3477_n2614), .B(
        DP_OP_425J2_127_3477_n2570), .CI(DP_OP_425J2_127_3477_n2746), .CO(
        DP_OP_425J2_127_3477_n855), .S(DP_OP_425J2_127_3477_n856) );
  FADDX1_HVT DP_OP_425J2_127_3477_U523 ( .A(DP_OP_425J2_127_3477_n2309), .B(
        DP_OP_425J2_127_3477_n2177), .CI(DP_OP_425J2_127_3477_n1957), .CO(
        DP_OP_425J2_127_3477_n853), .S(DP_OP_425J2_127_3477_n854) );
  FADDX1_HVT DP_OP_425J2_127_3477_U522 ( .A(DP_OP_425J2_127_3477_n2834), .B(
        DP_OP_425J2_127_3477_n1978), .CI(DP_OP_425J2_127_3477_n1913), .CO(
        DP_OP_425J2_127_3477_n851), .S(DP_OP_425J2_127_3477_n852) );
  FADDX1_HVT DP_OP_425J2_127_3477_U521 ( .A(DP_OP_425J2_127_3477_n2133), .B(
        DP_OP_425J2_127_3477_n2679), .CI(DP_OP_425J2_127_3477_n2022), .CO(
        DP_OP_425J2_127_3477_n849), .S(DP_OP_425J2_127_3477_n850) );
  FADDX1_HVT DP_OP_425J2_127_3477_U520 ( .A(DP_OP_425J2_127_3477_n2790), .B(
        DP_OP_425J2_127_3477_n2635), .CI(DP_OP_425J2_127_3477_n2330), .CO(
        DP_OP_425J2_127_3477_n847), .S(DP_OP_425J2_127_3477_n848) );
  FADDX1_HVT DP_OP_425J2_127_3477_U519 ( .A(DP_OP_425J2_127_3477_n2265), .B(
        DP_OP_425J2_127_3477_n1846), .CI(DP_OP_425J2_127_3477_n2198), .CO(
        DP_OP_425J2_127_3477_n845), .S(DP_OP_425J2_127_3477_n846) );
  FADDX1_HVT DP_OP_425J2_127_3477_U518 ( .A(DP_OP_425J2_127_3477_n2110), .B(
        DP_OP_425J2_127_3477_n2547), .CI(DP_OP_425J2_127_3477_n2415), .CO(
        DP_OP_425J2_127_3477_n843), .S(DP_OP_425J2_127_3477_n844) );
  FADDX1_HVT DP_OP_425J2_127_3477_U517 ( .A(DP_OP_425J2_127_3477_n2878), .B(
        DP_OP_425J2_127_3477_n2591), .CI(DP_OP_425J2_127_3477_n2459), .CO(
        DP_OP_425J2_127_3477_n841), .S(DP_OP_425J2_127_3477_n842) );
  FADDX1_HVT DP_OP_425J2_127_3477_U516 ( .A(DP_OP_425J2_127_3477_n2066), .B(
        DP_OP_425J2_127_3477_n2577), .CI(DP_OP_425J2_127_3477_n2279), .CO(
        DP_OP_425J2_127_3477_n839), .S(DP_OP_425J2_127_3477_n840) );
  FADDX1_HVT DP_OP_425J2_127_3477_U515 ( .A(DP_OP_425J2_127_3477_n2286), .B(
        DP_OP_425J2_127_3477_n2242), .CI(DP_OP_425J2_127_3477_n2804), .CO(
        DP_OP_425J2_127_3477_n837), .S(DP_OP_425J2_127_3477_n838) );
  FADDX1_HVT DP_OP_425J2_127_3477_U514 ( .A(DP_OP_425J2_127_3477_n2221), .B(
        DP_OP_425J2_127_3477_n2533), .CI(DP_OP_425J2_127_3477_n2316), .CO(
        DP_OP_425J2_127_3477_n835), .S(DP_OP_425J2_127_3477_n836) );
  FADDX1_HVT DP_OP_425J2_127_3477_U513 ( .A(DP_OP_425J2_127_3477_n2841), .B(
        DP_OP_425J2_127_3477_n1964), .CI(DP_OP_425J2_127_3477_n2140), .CO(
        DP_OP_425J2_127_3477_n833), .S(DP_OP_425J2_127_3477_n834) );
  FADDX1_HVT DP_OP_425J2_127_3477_U512 ( .A(DP_OP_425J2_127_3477_n2885), .B(
        DP_OP_425J2_127_3477_n2147), .CI(DP_OP_425J2_127_3477_n2272), .CO(
        DP_OP_425J2_127_3477_n831), .S(DP_OP_425J2_127_3477_n832) );
  FADDX1_HVT DP_OP_425J2_127_3477_U511 ( .A(DP_OP_425J2_127_3477_n2323), .B(
        DP_OP_425J2_127_3477_n2408), .CI(DP_OP_425J2_127_3477_n2052), .CO(
        DP_OP_425J2_127_3477_n829), .S(DP_OP_425J2_127_3477_n830) );
  FADDX1_HVT DP_OP_425J2_127_3477_U510 ( .A(DP_OP_425J2_127_3477_n1839), .B(
        DP_OP_425J2_127_3477_n1781), .CI(DP_OP_425J2_127_3477_n2892), .CO(
        DP_OP_425J2_127_3477_n827), .S(DP_OP_425J2_127_3477_n828) );
  FADDX1_HVT DP_OP_425J2_127_3477_U509 ( .A(DP_OP_425J2_127_3477_n2059), .B(
        DP_OP_425J2_127_3477_n2753), .CI(DP_OP_425J2_127_3477_n2154), .CO(
        DP_OP_425J2_127_3477_n825), .S(DP_OP_425J2_127_3477_n826) );
  FADDX1_HVT DP_OP_425J2_127_3477_U508 ( .A(DP_OP_425J2_127_3477_n2584), .B(
        DP_OP_425J2_127_3477_n2496), .CI(DP_OP_425J2_127_3477_n2848), .CO(
        DP_OP_425J2_127_3477_n823), .S(DP_OP_425J2_127_3477_n824) );
  FADDX1_HVT DP_OP_425J2_127_3477_U507 ( .A(DP_OP_425J2_127_3477_n2628), .B(
        DP_OP_425J2_127_3477_n2228), .CI(DP_OP_425J2_127_3477_n2540), .CO(
        DP_OP_425J2_127_3477_n821), .S(DP_OP_425J2_127_3477_n822) );
  FADDX1_HVT DP_OP_425J2_127_3477_U506 ( .A(DP_OP_425J2_127_3477_n2096), .B(
        DP_OP_425J2_127_3477_n2709), .CI(DP_OP_425J2_127_3477_n2184), .CO(
        DP_OP_425J2_127_3477_n819), .S(DP_OP_425J2_127_3477_n820) );
  FADDX1_HVT DP_OP_425J2_127_3477_U505 ( .A(DP_OP_425J2_127_3477_n2445), .B(
        DP_OP_425J2_127_3477_n2371), .CI(DP_OP_425J2_127_3477_n1920), .CO(
        DP_OP_425J2_127_3477_n817), .S(DP_OP_425J2_127_3477_n818) );
  FADDX1_HVT DP_OP_425J2_127_3477_U504 ( .A(DP_OP_425J2_127_3477_n2899), .B(
        DP_OP_425J2_127_3477_n2760), .CI(DP_OP_425J2_127_3477_n1876), .CO(
        DP_OP_425J2_127_3477_n815), .S(DP_OP_425J2_127_3477_n816) );
  FADDX1_HVT DP_OP_425J2_127_3477_U503 ( .A(DP_OP_425J2_127_3477_n2665), .B(
        DP_OP_425J2_127_3477_n1832), .CI(DP_OP_425J2_127_3477_n1927), .CO(
        DP_OP_425J2_127_3477_n813), .S(DP_OP_425J2_127_3477_n814) );
  FADDX1_HVT DP_OP_425J2_127_3477_U502 ( .A(DP_OP_425J2_127_3477_n2103), .B(
        DP_OP_425J2_127_3477_n2452), .CI(DP_OP_425J2_127_3477_n2235), .CO(
        DP_OP_425J2_127_3477_n811), .S(DP_OP_425J2_127_3477_n812) );
  FADDX1_HVT DP_OP_425J2_127_3477_U501 ( .A(DP_OP_425J2_127_3477_n1883), .B(
        DP_OP_425J2_127_3477_n2811), .CI(DP_OP_425J2_127_3477_n2364), .CO(
        DP_OP_425J2_127_3477_n809), .S(DP_OP_425J2_127_3477_n810) );
  FADDX1_HVT DP_OP_425J2_127_3477_U500 ( .A(DP_OP_425J2_127_3477_n2489), .B(
        DP_OP_425J2_127_3477_n1971), .CI(DP_OP_425J2_127_3477_n2008), .CO(
        DP_OP_425J2_127_3477_n807), .S(DP_OP_425J2_127_3477_n808) );
  FADDX1_HVT DP_OP_425J2_127_3477_U499 ( .A(DP_OP_425J2_127_3477_n2672), .B(
        DP_OP_425J2_127_3477_n2621), .CI(DP_OP_425J2_127_3477_n2191), .CO(
        DP_OP_425J2_127_3477_n805), .S(DP_OP_425J2_127_3477_n806) );
  FADDX1_HVT DP_OP_425J2_127_3477_U498 ( .A(DP_OP_425J2_127_3477_n2357), .B(
        DP_OP_425J2_127_3477_n2797), .CI(DP_OP_425J2_127_3477_n2401), .CO(
        DP_OP_425J2_127_3477_n803), .S(DP_OP_425J2_127_3477_n804) );
  FADDX1_HVT DP_OP_425J2_127_3477_U497 ( .A(DP_OP_425J2_127_3477_n2716), .B(
        DP_OP_425J2_127_3477_n1061), .CI(DP_OP_425J2_127_3477_n2015), .CO(
        DP_OP_425J2_127_3477_n801), .S(DP_OP_425J2_127_3477_n802) );
  FADDX1_HVT DP_OP_425J2_127_3477_U496 ( .A(DP_OP_425J2_127_3477_n1059), .B(
        DP_OP_425J2_127_3477_n1047), .CI(DP_OP_425J2_127_3477_n1045), .CO(
        DP_OP_425J2_127_3477_n799), .S(DP_OP_425J2_127_3477_n800) );
  FADDX1_HVT DP_OP_425J2_127_3477_U495 ( .A(DP_OP_425J2_127_3477_n1057), .B(
        DP_OP_425J2_127_3477_n1049), .CI(DP_OP_425J2_127_3477_n1055), .CO(
        DP_OP_425J2_127_3477_n797), .S(DP_OP_425J2_127_3477_n798) );
  FADDX1_HVT DP_OP_425J2_127_3477_U494 ( .A(DP_OP_425J2_127_3477_n1051), .B(
        DP_OP_425J2_127_3477_n1053), .CI(DP_OP_425J2_127_3477_n1025), .CO(
        DP_OP_425J2_127_3477_n795), .S(DP_OP_425J2_127_3477_n796) );
  FADDX1_HVT DP_OP_425J2_127_3477_U493 ( .A(DP_OP_425J2_127_3477_n1043), .B(
        DP_OP_425J2_127_3477_n1017), .CI(DP_OP_425J2_127_3477_n1011), .CO(
        DP_OP_425J2_127_3477_n793), .S(DP_OP_425J2_127_3477_n794) );
  FADDX1_HVT DP_OP_425J2_127_3477_U492 ( .A(DP_OP_425J2_127_3477_n1041), .B(
        DP_OP_425J2_127_3477_n1019), .CI(DP_OP_425J2_127_3477_n1013), .CO(
        DP_OP_425J2_127_3477_n791), .S(DP_OP_425J2_127_3477_n792) );
  FADDX1_HVT DP_OP_425J2_127_3477_U491 ( .A(DP_OP_425J2_127_3477_n1039), .B(
        DP_OP_425J2_127_3477_n1021), .CI(DP_OP_425J2_127_3477_n1015), .CO(
        DP_OP_425J2_127_3477_n789), .S(DP_OP_425J2_127_3477_n790) );
  FADDX1_HVT DP_OP_425J2_127_3477_U490 ( .A(DP_OP_425J2_127_3477_n1037), .B(
        DP_OP_425J2_127_3477_n1035), .CI(DP_OP_425J2_127_3477_n1023), .CO(
        DP_OP_425J2_127_3477_n787), .S(DP_OP_425J2_127_3477_n788) );
  FADDX1_HVT DP_OP_425J2_127_3477_U489 ( .A(DP_OP_425J2_127_3477_n1031), .B(
        DP_OP_425J2_127_3477_n1033), .CI(DP_OP_425J2_127_3477_n1029), .CO(
        DP_OP_425J2_127_3477_n785), .S(DP_OP_425J2_127_3477_n786) );
  FADDX1_HVT DP_OP_425J2_127_3477_U488 ( .A(DP_OP_425J2_127_3477_n1027), .B(
        DP_OP_425J2_127_3477_n1009), .CI(DP_OP_425J2_127_3477_n1005), .CO(
        DP_OP_425J2_127_3477_n783), .S(DP_OP_425J2_127_3477_n784) );
  FADDX1_HVT DP_OP_425J2_127_3477_U487 ( .A(DP_OP_425J2_127_3477_n1003), .B(
        DP_OP_425J2_127_3477_n844), .CI(DP_OP_425J2_127_3477_n995), .CO(
        DP_OP_425J2_127_3477_n781), .S(DP_OP_425J2_127_3477_n782) );
  FADDX1_HVT DP_OP_425J2_127_3477_U486 ( .A(DP_OP_425J2_127_3477_n1007), .B(
        DP_OP_425J2_127_3477_n846), .CI(DP_OP_425J2_127_3477_n997), .CO(
        DP_OP_425J2_127_3477_n779), .S(DP_OP_425J2_127_3477_n780) );
  FADDX1_HVT DP_OP_425J2_127_3477_U485 ( .A(DP_OP_425J2_127_3477_n1001), .B(
        DP_OP_425J2_127_3477_n848), .CI(DP_OP_425J2_127_3477_n842), .CO(
        DP_OP_425J2_127_3477_n777), .S(DP_OP_425J2_127_3477_n778) );
  FADDX1_HVT DP_OP_425J2_127_3477_U484 ( .A(DP_OP_425J2_127_3477_n999), .B(
        DP_OP_425J2_127_3477_n858), .CI(DP_OP_425J2_127_3477_n856), .CO(
        DP_OP_425J2_127_3477_n775), .S(DP_OP_425J2_127_3477_n776) );
  FADDX1_HVT DP_OP_425J2_127_3477_U483 ( .A(DP_OP_425J2_127_3477_n868), .B(
        DP_OP_425J2_127_3477_n852), .CI(DP_OP_425J2_127_3477_n854), .CO(
        DP_OP_425J2_127_3477_n773), .S(DP_OP_425J2_127_3477_n774) );
  FADDX1_HVT DP_OP_425J2_127_3477_U482 ( .A(DP_OP_425J2_127_3477_n866), .B(
        DP_OP_425J2_127_3477_n850), .CI(DP_OP_425J2_127_3477_n862), .CO(
        DP_OP_425J2_127_3477_n771), .S(DP_OP_425J2_127_3477_n772) );
  FADDX1_HVT DP_OP_425J2_127_3477_U481 ( .A(DP_OP_425J2_127_3477_n864), .B(
        DP_OP_425J2_127_3477_n860), .CI(DP_OP_425J2_127_3477_n840), .CO(
        DP_OP_425J2_127_3477_n769), .S(DP_OP_425J2_127_3477_n770) );
  FADDX1_HVT DP_OP_425J2_127_3477_U480 ( .A(DP_OP_425J2_127_3477_n838), .B(
        DP_OP_425J2_127_3477_n822), .CI(DP_OP_425J2_127_3477_n816), .CO(
        DP_OP_425J2_127_3477_n767), .S(DP_OP_425J2_127_3477_n768) );
  FADDX1_HVT DP_OP_425J2_127_3477_U479 ( .A(DP_OP_425J2_127_3477_n836), .B(
        DP_OP_425J2_127_3477_n826), .CI(DP_OP_425J2_127_3477_n818), .CO(
        DP_OP_425J2_127_3477_n765), .S(DP_OP_425J2_127_3477_n766) );
  FADDX1_HVT DP_OP_425J2_127_3477_U478 ( .A(DP_OP_425J2_127_3477_n832), .B(
        DP_OP_425J2_127_3477_n824), .CI(DP_OP_425J2_127_3477_n820), .CO(
        DP_OP_425J2_127_3477_n763), .S(DP_OP_425J2_127_3477_n764) );
  FADDX1_HVT DP_OP_425J2_127_3477_U477 ( .A(DP_OP_425J2_127_3477_n834), .B(
        DP_OP_425J2_127_3477_n828), .CI(DP_OP_425J2_127_3477_n830), .CO(
        DP_OP_425J2_127_3477_n761), .S(DP_OP_425J2_127_3477_n762) );
  FADDX1_HVT DP_OP_425J2_127_3477_U476 ( .A(DP_OP_425J2_127_3477_n814), .B(
        DP_OP_425J2_127_3477_n804), .CI(DP_OP_425J2_127_3477_n802), .CO(
        DP_OP_425J2_127_3477_n759), .S(DP_OP_425J2_127_3477_n760) );
  FADDX1_HVT DP_OP_425J2_127_3477_U475 ( .A(DP_OP_425J2_127_3477_n810), .B(
        DP_OP_425J2_127_3477_n806), .CI(DP_OP_425J2_127_3477_n993), .CO(
        DP_OP_425J2_127_3477_n757), .S(DP_OP_425J2_127_3477_n758) );
  FADDX1_HVT DP_OP_425J2_127_3477_U474 ( .A(DP_OP_425J2_127_3477_n812), .B(
        DP_OP_425J2_127_3477_n808), .CI(DP_OP_425J2_127_3477_n991), .CO(
        DP_OP_425J2_127_3477_n755), .S(DP_OP_425J2_127_3477_n756) );
  FADDX1_HVT DP_OP_425J2_127_3477_U473 ( .A(DP_OP_425J2_127_3477_n989), .B(
        DP_OP_425J2_127_3477_n987), .CI(DP_OP_425J2_127_3477_n985), .CO(
        DP_OP_425J2_127_3477_n753), .S(DP_OP_425J2_127_3477_n754) );
  FADDX1_HVT DP_OP_425J2_127_3477_U472 ( .A(DP_OP_425J2_127_3477_n983), .B(
        DP_OP_425J2_127_3477_n977), .CI(DP_OP_425J2_127_3477_n979), .CO(
        DP_OP_425J2_127_3477_n751), .S(DP_OP_425J2_127_3477_n752) );
  FADDX1_HVT DP_OP_425J2_127_3477_U471 ( .A(DP_OP_425J2_127_3477_n981), .B(
        DP_OP_425J2_127_3477_n975), .CI(DP_OP_425J2_127_3477_n973), .CO(
        DP_OP_425J2_127_3477_n749), .S(DP_OP_425J2_127_3477_n750) );
  FADDX1_HVT DP_OP_425J2_127_3477_U470 ( .A(DP_OP_425J2_127_3477_n971), .B(
        DP_OP_425J2_127_3477_n798), .CI(DP_OP_425J2_127_3477_n796), .CO(
        DP_OP_425J2_127_3477_n747), .S(DP_OP_425J2_127_3477_n748) );
  FADDX1_HVT DP_OP_425J2_127_3477_U469 ( .A(DP_OP_425J2_127_3477_n969), .B(
        DP_OP_425J2_127_3477_n967), .CI(DP_OP_425J2_127_3477_n800), .CO(
        DP_OP_425J2_127_3477_n745), .S(DP_OP_425J2_127_3477_n746) );
  FADDX1_HVT DP_OP_425J2_127_3477_U468 ( .A(DP_OP_425J2_127_3477_n965), .B(
        DP_OP_425J2_127_3477_n788), .CI(DP_OP_425J2_127_3477_n794), .CO(
        DP_OP_425J2_127_3477_n743), .S(DP_OP_425J2_127_3477_n744) );
  FADDX1_HVT DP_OP_425J2_127_3477_U467 ( .A(DP_OP_425J2_127_3477_n959), .B(
        DP_OP_425J2_127_3477_n792), .CI(DP_OP_425J2_127_3477_n784), .CO(
        DP_OP_425J2_127_3477_n741), .S(DP_OP_425J2_127_3477_n742) );
  FADDX1_HVT DP_OP_425J2_127_3477_U466 ( .A(DP_OP_425J2_127_3477_n963), .B(
        DP_OP_425J2_127_3477_n961), .CI(DP_OP_425J2_127_3477_n790), .CO(
        DP_OP_425J2_127_3477_n739), .S(DP_OP_425J2_127_3477_n740) );
  FADDX1_HVT DP_OP_425J2_127_3477_U465 ( .A(DP_OP_425J2_127_3477_n957), .B(
        DP_OP_425J2_127_3477_n786), .CI(DP_OP_425J2_127_3477_n955), .CO(
        DP_OP_425J2_127_3477_n737), .S(DP_OP_425J2_127_3477_n738) );
  FADDX1_HVT DP_OP_425J2_127_3477_U464 ( .A(DP_OP_425J2_127_3477_n953), .B(
        DP_OP_425J2_127_3477_n772), .CI(DP_OP_425J2_127_3477_n770), .CO(
        DP_OP_425J2_127_3477_n735), .S(DP_OP_425J2_127_3477_n736) );
  FADDX1_HVT DP_OP_425J2_127_3477_U463 ( .A(DP_OP_425J2_127_3477_n951), .B(
        DP_OP_425J2_127_3477_n776), .CI(DP_OP_425J2_127_3477_n774), .CO(
        DP_OP_425J2_127_3477_n733), .S(DP_OP_425J2_127_3477_n734) );
  FADDX1_HVT DP_OP_425J2_127_3477_U462 ( .A(DP_OP_425J2_127_3477_n949), .B(
        DP_OP_425J2_127_3477_n782), .CI(DP_OP_425J2_127_3477_n778), .CO(
        DP_OP_425J2_127_3477_n731), .S(DP_OP_425J2_127_3477_n732) );
  FADDX1_HVT DP_OP_425J2_127_3477_U461 ( .A(DP_OP_425J2_127_3477_n780), .B(
        DP_OP_425J2_127_3477_n768), .CI(DP_OP_425J2_127_3477_n766), .CO(
        DP_OP_425J2_127_3477_n729), .S(DP_OP_425J2_127_3477_n730) );
  FADDX1_HVT DP_OP_425J2_127_3477_U460 ( .A(DP_OP_425J2_127_3477_n762), .B(
        DP_OP_425J2_127_3477_n764), .CI(DP_OP_425J2_127_3477_n947), .CO(
        DP_OP_425J2_127_3477_n727), .S(DP_OP_425J2_127_3477_n728) );
  FADDX1_HVT DP_OP_425J2_127_3477_U459 ( .A(DP_OP_425J2_127_3477_n760), .B(
        DP_OP_425J2_127_3477_n943), .CI(DP_OP_425J2_127_3477_n756), .CO(
        DP_OP_425J2_127_3477_n725), .S(DP_OP_425J2_127_3477_n726) );
  FADDX1_HVT DP_OP_425J2_127_3477_U458 ( .A(DP_OP_425J2_127_3477_n758), .B(
        DP_OP_425J2_127_3477_n945), .CI(DP_OP_425J2_127_3477_n941), .CO(
        DP_OP_425J2_127_3477_n723), .S(DP_OP_425J2_127_3477_n724) );
  FADDX1_HVT DP_OP_425J2_127_3477_U457 ( .A(DP_OP_425J2_127_3477_n939), .B(
        DP_OP_425J2_127_3477_n937), .CI(DP_OP_425J2_127_3477_n754), .CO(
        DP_OP_425J2_127_3477_n721), .S(DP_OP_425J2_127_3477_n722) );
  FADDX1_HVT DP_OP_425J2_127_3477_U456 ( .A(DP_OP_425J2_127_3477_n935), .B(
        DP_OP_425J2_127_3477_n752), .CI(DP_OP_425J2_127_3477_n750), .CO(
        DP_OP_425J2_127_3477_n719), .S(DP_OP_425J2_127_3477_n720) );
  FADDX1_HVT DP_OP_425J2_127_3477_U455 ( .A(DP_OP_425J2_127_3477_n933), .B(
        DP_OP_425J2_127_3477_n931), .CI(DP_OP_425J2_127_3477_n929), .CO(
        DP_OP_425J2_127_3477_n717), .S(DP_OP_425J2_127_3477_n718) );
  FADDX1_HVT DP_OP_425J2_127_3477_U454 ( .A(DP_OP_425J2_127_3477_n927), .B(
        DP_OP_425J2_127_3477_n746), .CI(DP_OP_425J2_127_3477_n748), .CO(
        DP_OP_425J2_127_3477_n715), .S(DP_OP_425J2_127_3477_n716) );
  FADDX1_HVT DP_OP_425J2_127_3477_U453 ( .A(DP_OP_425J2_127_3477_n925), .B(
        DP_OP_425J2_127_3477_n923), .CI(DP_OP_425J2_127_3477_n744), .CO(
        DP_OP_425J2_127_3477_n713), .S(DP_OP_425J2_127_3477_n714) );
  FADDX1_HVT DP_OP_425J2_127_3477_U452 ( .A(DP_OP_425J2_127_3477_n921), .B(
        DP_OP_425J2_127_3477_n742), .CI(DP_OP_425J2_127_3477_n919), .CO(
        DP_OP_425J2_127_3477_n711), .S(DP_OP_425J2_127_3477_n712) );
  FADDX1_HVT DP_OP_425J2_127_3477_U451 ( .A(DP_OP_425J2_127_3477_n740), .B(
        DP_OP_425J2_127_3477_n738), .CI(DP_OP_425J2_127_3477_n736), .CO(
        DP_OP_425J2_127_3477_n709), .S(DP_OP_425J2_127_3477_n710) );
  FADDX1_HVT DP_OP_425J2_127_3477_U450 ( .A(DP_OP_425J2_127_3477_n917), .B(
        DP_OP_425J2_127_3477_n732), .CI(DP_OP_425J2_127_3477_n734), .CO(
        DP_OP_425J2_127_3477_n707), .S(DP_OP_425J2_127_3477_n708) );
  FADDX1_HVT DP_OP_425J2_127_3477_U449 ( .A(DP_OP_425J2_127_3477_n730), .B(
        DP_OP_425J2_127_3477_n915), .CI(DP_OP_425J2_127_3477_n728), .CO(
        DP_OP_425J2_127_3477_n705), .S(DP_OP_425J2_127_3477_n706) );
  FADDX1_HVT DP_OP_425J2_127_3477_U448 ( .A(DP_OP_425J2_127_3477_n913), .B(
        DP_OP_425J2_127_3477_n726), .CI(DP_OP_425J2_127_3477_n724), .CO(
        DP_OP_425J2_127_3477_n703), .S(DP_OP_425J2_127_3477_n704) );
  FADDX1_HVT DP_OP_425J2_127_3477_U447 ( .A(DP_OP_425J2_127_3477_n911), .B(
        DP_OP_425J2_127_3477_n909), .CI(DP_OP_425J2_127_3477_n907), .CO(
        DP_OP_425J2_127_3477_n701), .S(DP_OP_425J2_127_3477_n702) );
  FADDX1_HVT DP_OP_425J2_127_3477_U446 ( .A(DP_OP_425J2_127_3477_n722), .B(
        DP_OP_425J2_127_3477_n905), .CI(DP_OP_425J2_127_3477_n903), .CO(
        DP_OP_425J2_127_3477_n699), .S(DP_OP_425J2_127_3477_n700) );
  FADDX1_HVT DP_OP_425J2_127_3477_U445 ( .A(DP_OP_425J2_127_3477_n720), .B(
        DP_OP_425J2_127_3477_n718), .CI(DP_OP_425J2_127_3477_n901), .CO(
        DP_OP_425J2_127_3477_n697), .S(DP_OP_425J2_127_3477_n698) );
  FADDX1_HVT DP_OP_425J2_127_3477_U444 ( .A(DP_OP_425J2_127_3477_n716), .B(
        DP_OP_425J2_127_3477_n899), .CI(DP_OP_425J2_127_3477_n714), .CO(
        DP_OP_425J2_127_3477_n695), .S(DP_OP_425J2_127_3477_n696) );
  FADDX1_HVT DP_OP_425J2_127_3477_U443 ( .A(DP_OP_425J2_127_3477_n712), .B(
        DP_OP_425J2_127_3477_n710), .CI(DP_OP_425J2_127_3477_n897), .CO(
        DP_OP_425J2_127_3477_n693), .S(DP_OP_425J2_127_3477_n694) );
  FADDX1_HVT DP_OP_425J2_127_3477_U442 ( .A(DP_OP_425J2_127_3477_n708), .B(
        DP_OP_425J2_127_3477_n895), .CI(DP_OP_425J2_127_3477_n706), .CO(
        DP_OP_425J2_127_3477_n691), .S(DP_OP_425J2_127_3477_n692) );
  FADDX1_HVT DP_OP_425J2_127_3477_U441 ( .A(DP_OP_425J2_127_3477_n893), .B(
        DP_OP_425J2_127_3477_n704), .CI(DP_OP_425J2_127_3477_n891), .CO(
        DP_OP_425J2_127_3477_n689), .S(DP_OP_425J2_127_3477_n690) );
  FADDX1_HVT DP_OP_425J2_127_3477_U440 ( .A(DP_OP_425J2_127_3477_n702), .B(
        DP_OP_425J2_127_3477_n889), .CI(DP_OP_425J2_127_3477_n700), .CO(
        DP_OP_425J2_127_3477_n687), .S(DP_OP_425J2_127_3477_n688) );
  FADDX1_HVT DP_OP_425J2_127_3477_U439 ( .A(DP_OP_425J2_127_3477_n887), .B(
        DP_OP_425J2_127_3477_n698), .CI(DP_OP_425J2_127_3477_n885), .CO(
        DP_OP_425J2_127_3477_n685), .S(DP_OP_425J2_127_3477_n686) );
  FADDX1_HVT DP_OP_425J2_127_3477_U438 ( .A(DP_OP_425J2_127_3477_n696), .B(
        DP_OP_425J2_127_3477_n694), .CI(DP_OP_425J2_127_3477_n883), .CO(
        DP_OP_425J2_127_3477_n683), .S(DP_OP_425J2_127_3477_n684) );
  FADDX1_HVT DP_OP_425J2_127_3477_U437 ( .A(DP_OP_425J2_127_3477_n692), .B(
        DP_OP_425J2_127_3477_n881), .CI(DP_OP_425J2_127_3477_n690), .CO(
        DP_OP_425J2_127_3477_n681), .S(DP_OP_425J2_127_3477_n682) );
  FADDX1_HVT DP_OP_425J2_127_3477_U436 ( .A(DP_OP_425J2_127_3477_n879), .B(
        DP_OP_425J2_127_3477_n688), .CI(DP_OP_425J2_127_3477_n877), .CO(
        DP_OP_425J2_127_3477_n679), .S(DP_OP_425J2_127_3477_n680) );
  FADDX1_HVT DP_OP_425J2_127_3477_U435 ( .A(DP_OP_425J2_127_3477_n686), .B(
        DP_OP_425J2_127_3477_n875), .CI(DP_OP_425J2_127_3477_n684), .CO(
        DP_OP_425J2_127_3477_n677), .S(DP_OP_425J2_127_3477_n678) );
  FADDX1_HVT DP_OP_425J2_127_3477_U434 ( .A(DP_OP_425J2_127_3477_n682), .B(
        DP_OP_425J2_127_3477_n873), .CI(DP_OP_425J2_127_3477_n680), .CO(
        DP_OP_425J2_127_3477_n675), .S(DP_OP_425J2_127_3477_n676) );
  FADDX1_HVT DP_OP_425J2_127_3477_U433 ( .A(DP_OP_425J2_127_3477_n871), .B(
        DP_OP_425J2_127_3477_n678), .CI(DP_OP_425J2_127_3477_n676), .CO(
        DP_OP_425J2_127_3477_n673), .S(DP_OP_425J2_127_3477_n674) );
  FADDX1_HVT DP_OP_425J2_127_3477_U431 ( .A(DP_OP_425J2_127_3477_n2000), .B(
        DP_OP_425J2_127_3477_n1824), .CI(DP_OP_425J2_127_3477_n2847), .CO(
        DP_OP_425J2_127_3477_n669), .S(DP_OP_425J2_127_3477_n670) );
  FADDX1_HVT DP_OP_425J2_127_3477_U430 ( .A(DP_OP_425J2_127_3477_n2701), .B(
        DP_OP_425J2_127_3477_n2407), .CI(DP_OP_425J2_127_3477_n2539), .CO(
        DP_OP_425J2_127_3477_n667), .S(DP_OP_425J2_127_3477_n668) );
  FADDX1_HVT DP_OP_425J2_127_3477_U429 ( .A(DP_OP_425J2_127_3477_n2789), .B(
        DP_OP_425J2_127_3477_n2146), .CI(DP_OP_425J2_127_3477_n2393), .CO(
        DP_OP_425J2_127_3477_n665), .S(DP_OP_425J2_127_3477_n666) );
  FADDX1_HVT DP_OP_425J2_127_3477_U428 ( .A(DP_OP_425J2_127_3477_n2613), .B(
        DP_OP_425J2_127_3477_n2437), .CI(DP_OP_425J2_127_3477_n2745), .CO(
        DP_OP_425J2_127_3477_n663), .S(DP_OP_425J2_127_3477_n664) );
  FADDX1_HVT DP_OP_425J2_127_3477_U427 ( .A(DP_OP_425J2_127_3477_n2088), .B(
        DP_OP_425J2_127_3477_n2569), .CI(DP_OP_425J2_127_3477_n1956), .CO(
        DP_OP_425J2_127_3477_n661), .S(DP_OP_425J2_127_3477_n662) );
  FADDX1_HVT DP_OP_425J2_127_3477_U426 ( .A(DP_OP_425J2_127_3477_n2308), .B(
        DP_OP_425J2_127_3477_n2525), .CI(DP_OP_425J2_127_3477_n2481), .CO(
        DP_OP_425J2_127_3477_n659), .S(DP_OP_425J2_127_3477_n660) );
  FADDX1_HVT DP_OP_425J2_127_3477_U425 ( .A(DP_OP_425J2_127_3477_n1868), .B(
        DP_OP_425J2_127_3477_n2176), .CI(DP_OP_425J2_127_3477_n2044), .CO(
        DP_OP_425J2_127_3477_n657), .S(DP_OP_425J2_127_3477_n658) );
  FADDX1_HVT DP_OP_425J2_127_3477_U424 ( .A(DP_OP_425J2_127_3477_n2657), .B(
        DP_OP_425J2_127_3477_n2627), .CI(DP_OP_425J2_127_3477_n1912), .CO(
        DP_OP_425J2_127_3477_n655), .S(DP_OP_425J2_127_3477_n656) );
  FADDX1_HVT DP_OP_425J2_127_3477_U423 ( .A(DP_OP_425J2_127_3477_n2132), .B(
        DP_OP_425J2_127_3477_n1838), .CI(DP_OP_425J2_127_3477_n2058), .CO(
        DP_OP_425J2_127_3477_n653), .S(DP_OP_425J2_127_3477_n654) );
  FADDX1_HVT DP_OP_425J2_127_3477_U422 ( .A(DP_OP_425J2_127_3477_n2833), .B(
        DP_OP_425J2_127_3477_n2322), .CI(DP_OP_425J2_127_3477_n2583), .CO(
        DP_OP_425J2_127_3477_n651), .S(DP_OP_425J2_127_3477_n652) );
  FADDX1_HVT DP_OP_425J2_127_3477_U421 ( .A(DP_OP_425J2_127_3477_n2264), .B(
        DP_OP_425J2_127_3477_n2495), .CI(DP_OP_425J2_127_3477_n2891), .CO(
        DP_OP_425J2_127_3477_n649), .S(DP_OP_425J2_127_3477_n650) );
  FADDX1_HVT DP_OP_425J2_127_3477_U420 ( .A(DP_OP_425J2_127_3477_n2877), .B(
        DP_OP_425J2_127_3477_n2278), .CI(DP_OP_425J2_127_3477_n2803), .CO(
        DP_OP_425J2_127_3477_n647), .S(DP_OP_425J2_127_3477_n648) );
  FADDX1_HVT DP_OP_425J2_127_3477_U419 ( .A(DP_OP_425J2_127_3477_n672), .B(
        DP_OP_425J2_127_3477_n2576), .CI(DP_OP_425J2_127_3477_n2051), .CO(
        DP_OP_425J2_127_3477_n645), .S(DP_OP_425J2_127_3477_n646) );
  FADDX1_HVT DP_OP_425J2_127_3477_U418 ( .A(DP_OP_425J2_127_3477_n2220), .B(
        DP_OP_425J2_127_3477_n1970), .CI(DP_OP_425J2_127_3477_n2315), .CO(
        DP_OP_425J2_127_3477_n643), .S(DP_OP_425J2_127_3477_n644) );
  FADDX1_HVT DP_OP_425J2_127_3477_U417 ( .A(DP_OP_425J2_127_3477_n2840), .B(
        DP_OP_425J2_127_3477_n2451), .CI(DP_OP_425J2_127_3477_n2139), .CO(
        DP_OP_425J2_127_3477_n641), .S(DP_OP_425J2_127_3477_n642) );
  FADDX1_HVT DP_OP_425J2_127_3477_U416 ( .A(DP_OP_425J2_127_3477_n2884), .B(
        DP_OP_425J2_127_3477_n2532), .CI(DP_OP_425J2_127_3477_n2271), .CO(
        DP_OP_425J2_127_3477_n639), .S(DP_OP_425J2_127_3477_n640) );
  FADDX1_HVT DP_OP_425J2_127_3477_U415 ( .A(DP_OP_425J2_127_3477_n2752), .B(
        DP_OP_425J2_127_3477_n1963), .CI(DP_OP_425J2_127_3477_n2234), .CO(
        DP_OP_425J2_127_3477_n637), .S(DP_OP_425J2_127_3477_n638) );
  FADDX1_HVT DP_OP_425J2_127_3477_U414 ( .A(DP_OP_425J2_127_3477_n2759), .B(
        DP_OP_425J2_127_3477_n1780), .CI(DP_OP_425J2_127_3477_n2190), .CO(
        DP_OP_425J2_127_3477_n635), .S(DP_OP_425J2_127_3477_n636) );
  FADDX1_HVT DP_OP_425J2_127_3477_U413 ( .A(DP_OP_425J2_127_3477_n1882), .B(
        DP_OP_425J2_127_3477_n2671), .CI(DP_OP_425J2_127_3477_n2664), .CO(
        DP_OP_425J2_127_3477_n633), .S(DP_OP_425J2_127_3477_n634) );
  FADDX1_HVT DP_OP_425J2_127_3477_U412 ( .A(DP_OP_425J2_127_3477_n2102), .B(
        DP_OP_425J2_127_3477_n2227), .CI(DP_OP_425J2_127_3477_n2363), .CO(
        DP_OP_425J2_127_3477_n631), .S(DP_OP_425J2_127_3477_n632) );
  FADDX1_HVT DP_OP_425J2_127_3477_U411 ( .A(DP_OP_425J2_127_3477_n2095), .B(
        DP_OP_425J2_127_3477_n1926), .CI(DP_OP_425J2_127_3477_n2183), .CO(
        DP_OP_425J2_127_3477_n629), .S(DP_OP_425J2_127_3477_n630) );
  FADDX1_HVT DP_OP_425J2_127_3477_U410 ( .A(DP_OP_425J2_127_3477_n2444), .B(
        DP_OP_425J2_127_3477_n2014), .CI(DP_OP_425J2_127_3477_n1919), .CO(
        DP_OP_425J2_127_3477_n627), .S(DP_OP_425J2_127_3477_n628) );
  FADDX1_HVT DP_OP_425J2_127_3477_U409 ( .A(DP_OP_425J2_127_3477_n2715), .B(
        DP_OP_425J2_127_3477_n2708), .CI(DP_OP_425J2_127_3477_n1875), .CO(
        DP_OP_425J2_127_3477_n625), .S(DP_OP_425J2_127_3477_n626) );
  FADDX1_HVT DP_OP_425J2_127_3477_U408 ( .A(DP_OP_425J2_127_3477_n2488), .B(
        DP_OP_425J2_127_3477_n1831), .CI(DP_OP_425J2_127_3477_n2007), .CO(
        DP_OP_425J2_127_3477_n623), .S(DP_OP_425J2_127_3477_n624) );
  FADDX1_HVT DP_OP_425J2_127_3477_U407 ( .A(DP_OP_425J2_127_3477_n2356), .B(
        DP_OP_425J2_127_3477_n2620), .CI(DP_OP_425J2_127_3477_n2400), .CO(
        DP_OP_425J2_127_3477_n621), .S(DP_OP_425J2_127_3477_n622) );
  FADDX1_HVT DP_OP_425J2_127_3477_U406 ( .A(DP_OP_425J2_127_3477_n2796), .B(
        DP_OP_425J2_127_3477_n867), .CI(DP_OP_425J2_127_3477_n865), .CO(
        DP_OP_425J2_127_3477_n619), .S(DP_OP_425J2_127_3477_n620) );
  FADDX1_HVT DP_OP_425J2_127_3477_U405 ( .A(DP_OP_425J2_127_3477_n863), .B(
        DP_OP_425J2_127_3477_n843), .CI(DP_OP_425J2_127_3477_n841), .CO(
        DP_OP_425J2_127_3477_n617), .S(DP_OP_425J2_127_3477_n618) );
  FADDX1_HVT DP_OP_425J2_127_3477_U404 ( .A(DP_OP_425J2_127_3477_n861), .B(
        DP_OP_425J2_127_3477_n847), .CI(DP_OP_425J2_127_3477_n845), .CO(
        DP_OP_425J2_127_3477_n615), .S(DP_OP_425J2_127_3477_n616) );
  FADDX1_HVT DP_OP_425J2_127_3477_U403 ( .A(DP_OP_425J2_127_3477_n859), .B(
        DP_OP_425J2_127_3477_n849), .CI(DP_OP_425J2_127_3477_n851), .CO(
        DP_OP_425J2_127_3477_n613), .S(DP_OP_425J2_127_3477_n614) );
  FADDX1_HVT DP_OP_425J2_127_3477_U402 ( .A(DP_OP_425J2_127_3477_n857), .B(
        DP_OP_425J2_127_3477_n853), .CI(DP_OP_425J2_127_3477_n855), .CO(
        DP_OP_425J2_127_3477_n611), .S(DP_OP_425J2_127_3477_n612) );
  FADDX1_HVT DP_OP_425J2_127_3477_U401 ( .A(DP_OP_425J2_127_3477_n839), .B(
        DP_OP_425J2_127_3477_n821), .CI(DP_OP_425J2_127_3477_n815), .CO(
        DP_OP_425J2_127_3477_n609), .S(DP_OP_425J2_127_3477_n610) );
  FADDX1_HVT DP_OP_425J2_127_3477_U400 ( .A(DP_OP_425J2_127_3477_n837), .B(
        DP_OP_425J2_127_3477_n823), .CI(DP_OP_425J2_127_3477_n817), .CO(
        DP_OP_425J2_127_3477_n607), .S(DP_OP_425J2_127_3477_n608) );
  FADDX1_HVT DP_OP_425J2_127_3477_U399 ( .A(DP_OP_425J2_127_3477_n835), .B(
        DP_OP_425J2_127_3477_n825), .CI(DP_OP_425J2_127_3477_n819), .CO(
        DP_OP_425J2_127_3477_n605), .S(DP_OP_425J2_127_3477_n606) );
  FADDX1_HVT DP_OP_425J2_127_3477_U398 ( .A(DP_OP_425J2_127_3477_n833), .B(
        DP_OP_425J2_127_3477_n827), .CI(DP_OP_425J2_127_3477_n829), .CO(
        DP_OP_425J2_127_3477_n603), .S(DP_OP_425J2_127_3477_n604) );
  FADDX1_HVT DP_OP_425J2_127_3477_U397 ( .A(DP_OP_425J2_127_3477_n831), .B(
        DP_OP_425J2_127_3477_n813), .CI(DP_OP_425J2_127_3477_n807), .CO(
        DP_OP_425J2_127_3477_n601), .S(DP_OP_425J2_127_3477_n602) );
  FADDX1_HVT DP_OP_425J2_127_3477_U396 ( .A(DP_OP_425J2_127_3477_n811), .B(
        DP_OP_425J2_127_3477_n650), .CI(DP_OP_425J2_127_3477_n648), .CO(
        DP_OP_425J2_127_3477_n599), .S(DP_OP_425J2_127_3477_n600) );
  FADDX1_HVT DP_OP_425J2_127_3477_U395 ( .A(DP_OP_425J2_127_3477_n809), .B(
        DP_OP_425J2_127_3477_n666), .CI(DP_OP_425J2_127_3477_n801), .CO(
        DP_OP_425J2_127_3477_n597), .S(DP_OP_425J2_127_3477_n598) );
  FADDX1_HVT DP_OP_425J2_127_3477_U394 ( .A(DP_OP_425J2_127_3477_n805), .B(
        DP_OP_425J2_127_3477_n654), .CI(DP_OP_425J2_127_3477_n656), .CO(
        DP_OP_425J2_127_3477_n595), .S(DP_OP_425J2_127_3477_n596) );
  FADDX1_HVT DP_OP_425J2_127_3477_U393 ( .A(DP_OP_425J2_127_3477_n803), .B(
        DP_OP_425J2_127_3477_n662), .CI(DP_OP_425J2_127_3477_n658), .CO(
        DP_OP_425J2_127_3477_n593), .S(DP_OP_425J2_127_3477_n594) );
  FADDX1_HVT DP_OP_425J2_127_3477_U392 ( .A(DP_OP_425J2_127_3477_n670), .B(
        DP_OP_425J2_127_3477_n652), .CI(DP_OP_425J2_127_3477_n660), .CO(
        DP_OP_425J2_127_3477_n591), .S(DP_OP_425J2_127_3477_n592) );
  FADDX1_HVT DP_OP_425J2_127_3477_U391 ( .A(DP_OP_425J2_127_3477_n668), .B(
        DP_OP_425J2_127_3477_n664), .CI(DP_OP_425J2_127_3477_n646), .CO(
        DP_OP_425J2_127_3477_n589), .S(DP_OP_425J2_127_3477_n590) );
  FADDX1_HVT DP_OP_425J2_127_3477_U390 ( .A(DP_OP_425J2_127_3477_n644), .B(
        DP_OP_425J2_127_3477_n632), .CI(DP_OP_425J2_127_3477_n626), .CO(
        DP_OP_425J2_127_3477_n587), .S(DP_OP_425J2_127_3477_n588) );
  FADDX1_HVT DP_OP_425J2_127_3477_U389 ( .A(DP_OP_425J2_127_3477_n640), .B(
        DP_OP_425J2_127_3477_n634), .CI(DP_OP_425J2_127_3477_n628), .CO(
        DP_OP_425J2_127_3477_n585), .S(DP_OP_425J2_127_3477_n586) );
  FADDX1_HVT DP_OP_425J2_127_3477_U388 ( .A(DP_OP_425J2_127_3477_n642), .B(
        DP_OP_425J2_127_3477_n636), .CI(DP_OP_425J2_127_3477_n630), .CO(
        DP_OP_425J2_127_3477_n583), .S(DP_OP_425J2_127_3477_n584) );
  FADDX1_HVT DP_OP_425J2_127_3477_U387 ( .A(DP_OP_425J2_127_3477_n638), .B(
        DP_OP_425J2_127_3477_n624), .CI(DP_OP_425J2_127_3477_n622), .CO(
        DP_OP_425J2_127_3477_n581), .S(DP_OP_425J2_127_3477_n582) );
  FADDX1_HVT DP_OP_425J2_127_3477_U386 ( .A(DP_OP_425J2_127_3477_n799), .B(
        DP_OP_425J2_127_3477_n797), .CI(DP_OP_425J2_127_3477_n795), .CO(
        DP_OP_425J2_127_3477_n579), .S(DP_OP_425J2_127_3477_n580) );
  FADDX1_HVT DP_OP_425J2_127_3477_U385 ( .A(DP_OP_425J2_127_3477_n793), .B(
        DP_OP_425J2_127_3477_n785), .CI(DP_OP_425J2_127_3477_n783), .CO(
        DP_OP_425J2_127_3477_n577), .S(DP_OP_425J2_127_3477_n578) );
  FADDX1_HVT DP_OP_425J2_127_3477_U384 ( .A(DP_OP_425J2_127_3477_n791), .B(
        DP_OP_425J2_127_3477_n787), .CI(DP_OP_425J2_127_3477_n789), .CO(
        DP_OP_425J2_127_3477_n575), .S(DP_OP_425J2_127_3477_n576) );
  FADDX1_HVT DP_OP_425J2_127_3477_U383 ( .A(DP_OP_425J2_127_3477_n620), .B(
        DP_OP_425J2_127_3477_n775), .CI(DP_OP_425J2_127_3477_n616), .CO(
        DP_OP_425J2_127_3477_n573), .S(DP_OP_425J2_127_3477_n574) );
  FADDX1_HVT DP_OP_425J2_127_3477_U382 ( .A(DP_OP_425J2_127_3477_n781), .B(
        DP_OP_425J2_127_3477_n614), .CI(DP_OP_425J2_127_3477_n612), .CO(
        DP_OP_425J2_127_3477_n571), .S(DP_OP_425J2_127_3477_n572) );
  FADDX1_HVT DP_OP_425J2_127_3477_U381 ( .A(DP_OP_425J2_127_3477_n779), .B(
        DP_OP_425J2_127_3477_n618), .CI(DP_OP_425J2_127_3477_n769), .CO(
        DP_OP_425J2_127_3477_n569), .S(DP_OP_425J2_127_3477_n570) );
  FADDX1_HVT DP_OP_425J2_127_3477_U380 ( .A(DP_OP_425J2_127_3477_n777), .B(
        DP_OP_425J2_127_3477_n773), .CI(DP_OP_425J2_127_3477_n771), .CO(
        DP_OP_425J2_127_3477_n567), .S(DP_OP_425J2_127_3477_n568) );
  FADDX1_HVT DP_OP_425J2_127_3477_U379 ( .A(DP_OP_425J2_127_3477_n767), .B(
        DP_OP_425J2_127_3477_n761), .CI(DP_OP_425J2_127_3477_n602), .CO(
        DP_OP_425J2_127_3477_n565), .S(DP_OP_425J2_127_3477_n566) );
  FADDX1_HVT DP_OP_425J2_127_3477_U378 ( .A(DP_OP_425J2_127_3477_n608), .B(
        DP_OP_425J2_127_3477_n763), .CI(DP_OP_425J2_127_3477_n604), .CO(
        DP_OP_425J2_127_3477_n563), .S(DP_OP_425J2_127_3477_n564) );
  FADDX1_HVT DP_OP_425J2_127_3477_U377 ( .A(DP_OP_425J2_127_3477_n610), .B(
        DP_OP_425J2_127_3477_n765), .CI(DP_OP_425J2_127_3477_n606), .CO(
        DP_OP_425J2_127_3477_n561), .S(DP_OP_425J2_127_3477_n562) );
  FADDX1_HVT DP_OP_425J2_127_3477_U376 ( .A(DP_OP_425J2_127_3477_n759), .B(
        DP_OP_425J2_127_3477_n594), .CI(DP_OP_425J2_127_3477_n590), .CO(
        DP_OP_425J2_127_3477_n559), .S(DP_OP_425J2_127_3477_n560) );
  FADDX1_HVT DP_OP_425J2_127_3477_U375 ( .A(DP_OP_425J2_127_3477_n757), .B(
        DP_OP_425J2_127_3477_n592), .CI(DP_OP_425J2_127_3477_n755), .CO(
        DP_OP_425J2_127_3477_n557), .S(DP_OP_425J2_127_3477_n558) );
  FADDX1_HVT DP_OP_425J2_127_3477_U374 ( .A(DP_OP_425J2_127_3477_n598), .B(
        DP_OP_425J2_127_3477_n600), .CI(DP_OP_425J2_127_3477_n596), .CO(
        DP_OP_425J2_127_3477_n555), .S(DP_OP_425J2_127_3477_n556) );
  FADDX1_HVT DP_OP_425J2_127_3477_U373 ( .A(DP_OP_425J2_127_3477_n588), .B(
        DP_OP_425J2_127_3477_n753), .CI(DP_OP_425J2_127_3477_n582), .CO(
        DP_OP_425J2_127_3477_n553), .S(DP_OP_425J2_127_3477_n554) );
  FADDX1_HVT DP_OP_425J2_127_3477_U372 ( .A(DP_OP_425J2_127_3477_n584), .B(
        DP_OP_425J2_127_3477_n586), .CI(DP_OP_425J2_127_3477_n751), .CO(
        DP_OP_425J2_127_3477_n551), .S(DP_OP_425J2_127_3477_n552) );
  FADDX1_HVT DP_OP_425J2_127_3477_U371 ( .A(DP_OP_425J2_127_3477_n749), .B(
        DP_OP_425J2_127_3477_n747), .CI(DP_OP_425J2_127_3477_n580), .CO(
        DP_OP_425J2_127_3477_n549), .S(DP_OP_425J2_127_3477_n550) );
  FADDX1_HVT DP_OP_425J2_127_3477_U370 ( .A(DP_OP_425J2_127_3477_n745), .B(
        DP_OP_425J2_127_3477_n743), .CI(DP_OP_425J2_127_3477_n741), .CO(
        DP_OP_425J2_127_3477_n547), .S(DP_OP_425J2_127_3477_n548) );
  FADDX1_HVT DP_OP_425J2_127_3477_U369 ( .A(DP_OP_425J2_127_3477_n739), .B(
        DP_OP_425J2_127_3477_n576), .CI(DP_OP_425J2_127_3477_n578), .CO(
        DP_OP_425J2_127_3477_n545), .S(DP_OP_425J2_127_3477_n546) );
  FADDX1_HVT DP_OP_425J2_127_3477_U368 ( .A(DP_OP_425J2_127_3477_n737), .B(
        DP_OP_425J2_127_3477_n574), .CI(DP_OP_425J2_127_3477_n735), .CO(
        DP_OP_425J2_127_3477_n543), .S(DP_OP_425J2_127_3477_n544) );
  FADDX1_HVT DP_OP_425J2_127_3477_U367 ( .A(DP_OP_425J2_127_3477_n733), .B(
        DP_OP_425J2_127_3477_n568), .CI(DP_OP_425J2_127_3477_n729), .CO(
        DP_OP_425J2_127_3477_n541), .S(DP_OP_425J2_127_3477_n542) );
  FADDX1_HVT DP_OP_425J2_127_3477_U366 ( .A(DP_OP_425J2_127_3477_n572), .B(
        DP_OP_425J2_127_3477_n731), .CI(DP_OP_425J2_127_3477_n570), .CO(
        DP_OP_425J2_127_3477_n539), .S(DP_OP_425J2_127_3477_n540) );
  FADDX1_HVT DP_OP_425J2_127_3477_U365 ( .A(DP_OP_425J2_127_3477_n564), .B(
        DP_OP_425J2_127_3477_n562), .CI(DP_OP_425J2_127_3477_n727), .CO(
        DP_OP_425J2_127_3477_n537), .S(DP_OP_425J2_127_3477_n538) );
  FADDX1_HVT DP_OP_425J2_127_3477_U364 ( .A(DP_OP_425J2_127_3477_n566), .B(
        DP_OP_425J2_127_3477_n725), .CI(DP_OP_425J2_127_3477_n560), .CO(
        DP_OP_425J2_127_3477_n535), .S(DP_OP_425J2_127_3477_n536) );
  FADDX1_HVT DP_OP_425J2_127_3477_U363 ( .A(DP_OP_425J2_127_3477_n723), .B(
        DP_OP_425J2_127_3477_n558), .CI(DP_OP_425J2_127_3477_n556), .CO(
        DP_OP_425J2_127_3477_n533), .S(DP_OP_425J2_127_3477_n534) );
  FADDX1_HVT DP_OP_425J2_127_3477_U362 ( .A(DP_OP_425J2_127_3477_n721), .B(
        DP_OP_425J2_127_3477_n554), .CI(DP_OP_425J2_127_3477_n552), .CO(
        DP_OP_425J2_127_3477_n531), .S(DP_OP_425J2_127_3477_n532) );
  FADDX1_HVT DP_OP_425J2_127_3477_U361 ( .A(DP_OP_425J2_127_3477_n719), .B(
        DP_OP_425J2_127_3477_n717), .CI(DP_OP_425J2_127_3477_n550), .CO(
        DP_OP_425J2_127_3477_n529), .S(DP_OP_425J2_127_3477_n530) );
  FADDX1_HVT DP_OP_425J2_127_3477_U360 ( .A(DP_OP_425J2_127_3477_n715), .B(
        DP_OP_425J2_127_3477_n713), .CI(DP_OP_425J2_127_3477_n548), .CO(
        DP_OP_425J2_127_3477_n527), .S(DP_OP_425J2_127_3477_n528) );
  FADDX1_HVT DP_OP_425J2_127_3477_U359 ( .A(DP_OP_425J2_127_3477_n711), .B(
        DP_OP_425J2_127_3477_n709), .CI(DP_OP_425J2_127_3477_n544), .CO(
        DP_OP_425J2_127_3477_n525), .S(DP_OP_425J2_127_3477_n526) );
  FADDX1_HVT DP_OP_425J2_127_3477_U358 ( .A(DP_OP_425J2_127_3477_n546), .B(
        DP_OP_425J2_127_3477_n707), .CI(DP_OP_425J2_127_3477_n542), .CO(
        DP_OP_425J2_127_3477_n523), .S(DP_OP_425J2_127_3477_n524) );
  FADDX1_HVT DP_OP_425J2_127_3477_U357 ( .A(DP_OP_425J2_127_3477_n540), .B(
        DP_OP_425J2_127_3477_n705), .CI(DP_OP_425J2_127_3477_n538), .CO(
        DP_OP_425J2_127_3477_n521), .S(DP_OP_425J2_127_3477_n522) );
  FADDX1_HVT DP_OP_425J2_127_3477_U356 ( .A(DP_OP_425J2_127_3477_n536), .B(
        DP_OP_425J2_127_3477_n703), .CI(DP_OP_425J2_127_3477_n701), .CO(
        DP_OP_425J2_127_3477_n519), .S(DP_OP_425J2_127_3477_n520) );
  FADDX1_HVT DP_OP_425J2_127_3477_U355 ( .A(DP_OP_425J2_127_3477_n534), .B(
        DP_OP_425J2_127_3477_n532), .CI(DP_OP_425J2_127_3477_n699), .CO(
        DP_OP_425J2_127_3477_n517), .S(DP_OP_425J2_127_3477_n518) );
  FADDX1_HVT DP_OP_425J2_127_3477_U354 ( .A(DP_OP_425J2_127_3477_n697), .B(
        DP_OP_425J2_127_3477_n530), .CI(DP_OP_425J2_127_3477_n695), .CO(
        DP_OP_425J2_127_3477_n515), .S(DP_OP_425J2_127_3477_n516) );
  FADDX1_HVT DP_OP_425J2_127_3477_U353 ( .A(DP_OP_425J2_127_3477_n528), .B(
        DP_OP_425J2_127_3477_n526), .CI(DP_OP_425J2_127_3477_n693), .CO(
        DP_OP_425J2_127_3477_n513), .S(DP_OP_425J2_127_3477_n514) );
  FADDX1_HVT DP_OP_425J2_127_3477_U352 ( .A(DP_OP_425J2_127_3477_n524), .B(
        DP_OP_425J2_127_3477_n691), .CI(DP_OP_425J2_127_3477_n522), .CO(
        DP_OP_425J2_127_3477_n511), .S(DP_OP_425J2_127_3477_n512) );
  FADDX1_HVT DP_OP_425J2_127_3477_U351 ( .A(DP_OP_425J2_127_3477_n689), .B(
        DP_OP_425J2_127_3477_n520), .CI(DP_OP_425J2_127_3477_n687), .CO(
        DP_OP_425J2_127_3477_n509), .S(DP_OP_425J2_127_3477_n510) );
  FADDX1_HVT DP_OP_425J2_127_3477_U350 ( .A(DP_OP_425J2_127_3477_n518), .B(
        DP_OP_425J2_127_3477_n685), .CI(DP_OP_425J2_127_3477_n516), .CO(
        DP_OP_425J2_127_3477_n507), .S(DP_OP_425J2_127_3477_n508) );
  FADDX1_HVT DP_OP_425J2_127_3477_U349 ( .A(DP_OP_425J2_127_3477_n683), .B(
        DP_OP_425J2_127_3477_n514), .CI(DP_OP_425J2_127_3477_n512), .CO(
        DP_OP_425J2_127_3477_n505), .S(DP_OP_425J2_127_3477_n506) );
  FADDX1_HVT DP_OP_425J2_127_3477_U348 ( .A(DP_OP_425J2_127_3477_n681), .B(
        DP_OP_425J2_127_3477_n510), .CI(DP_OP_425J2_127_3477_n679), .CO(
        DP_OP_425J2_127_3477_n503), .S(DP_OP_425J2_127_3477_n504) );
  FADDX1_HVT DP_OP_425J2_127_3477_U347 ( .A(DP_OP_425J2_127_3477_n508), .B(
        DP_OP_425J2_127_3477_n677), .CI(DP_OP_425J2_127_3477_n506), .CO(
        DP_OP_425J2_127_3477_n501), .S(DP_OP_425J2_127_3477_n502) );
  FADDX1_HVT DP_OP_425J2_127_3477_U346 ( .A(DP_OP_425J2_127_3477_n675), .B(
        DP_OP_425J2_127_3477_n504), .CI(DP_OP_425J2_127_3477_n502), .CO(
        DP_OP_425J2_127_3477_n499), .S(DP_OP_425J2_127_3477_n500) );
  FADDX1_HVT DP_OP_425J2_127_3477_U345 ( .A(DP_OP_425J2_127_3477_n671), .B(
        DP_OP_425J2_127_3477_n1823), .CI(DP_OP_425J2_127_3477_n2707), .CO(
        DP_OP_425J2_127_3477_n497), .S(DP_OP_425J2_127_3477_n498) );
  FADDX1_HVT DP_OP_425J2_127_3477_U344 ( .A(DP_OP_425J2_127_3477_n2350), .B(
        DP_OP_425J2_127_3477_n1962), .CI(DP_OP_425J2_127_3477_n2443), .CO(
        DP_OP_425J2_127_3477_n495), .S(DP_OP_425J2_127_3477_n496) );
  FADDX1_HVT DP_OP_425J2_127_3477_U343 ( .A(DP_OP_425J2_127_3477_n1999), .B(
        DP_OP_425J2_127_3477_n2531), .CI(DP_OP_425J2_127_3477_n2226), .CO(
        DP_OP_425J2_127_3477_n493), .S(DP_OP_425J2_127_3477_n494) );
  FADDX1_HVT DP_OP_425J2_127_3477_U342 ( .A(DP_OP_425J2_127_3477_n2700), .B(
        DP_OP_425J2_127_3477_n2480), .CI(DP_OP_425J2_127_3477_n2094), .CO(
        DP_OP_425J2_127_3477_n491), .S(DP_OP_425J2_127_3477_n492) );
  FADDX1_HVT DP_OP_425J2_127_3477_U341 ( .A(DP_OP_425J2_127_3477_n2131), .B(
        DP_OP_425J2_127_3477_n2175), .CI(DP_OP_425J2_127_3477_n2392), .CO(
        DP_OP_425J2_127_3477_n489), .S(DP_OP_425J2_127_3477_n490) );
  FADDX1_HVT DP_OP_425J2_127_3477_U340 ( .A(DP_OP_425J2_127_3477_n2307), .B(
        DP_OP_425J2_127_3477_n2043), .CI(DP_OP_425J2_127_3477_n2744), .CO(
        DP_OP_425J2_127_3477_n487), .S(DP_OP_425J2_127_3477_n488) );
  FADDX1_HVT DP_OP_425J2_127_3477_U339 ( .A(DP_OP_425J2_127_3477_n2788), .B(
        DP_OP_425J2_127_3477_n1911), .CI(DP_OP_425J2_127_3477_n1955), .CO(
        DP_OP_425J2_127_3477_n485), .S(DP_OP_425J2_127_3477_n486) );
  FADDX1_HVT DP_OP_425J2_127_3477_U338 ( .A(DP_OP_425J2_127_3477_n2087), .B(
        DP_OP_425J2_127_3477_n2436), .CI(DP_OP_425J2_127_3477_n2575), .CO(
        DP_OP_425J2_127_3477_n483), .S(DP_OP_425J2_127_3477_n484) );
  FADDX1_HVT DP_OP_425J2_127_3477_U337 ( .A(DP_OP_425J2_127_3477_n2656), .B(
        DP_OP_425J2_127_3477_n2524), .CI(DP_OP_425J2_127_3477_n2568), .CO(
        DP_OP_425J2_127_3477_n481), .S(DP_OP_425J2_127_3477_n482) );
  FADDX1_HVT DP_OP_425J2_127_3477_U336 ( .A(DP_OP_425J2_127_3477_n2612), .B(
        DP_OP_425J2_127_3477_n2839), .CI(DP_OP_425J2_127_3477_n2751), .CO(
        DP_OP_425J2_127_3477_n479), .S(DP_OP_425J2_127_3477_n480) );
  FADDX1_HVT DP_OP_425J2_127_3477_U335 ( .A(DP_OP_425J2_127_3477_n2832), .B(
        DP_OP_425J2_127_3477_n2876), .CI(DP_OP_425J2_127_3477_n2883), .CO(
        DP_OP_425J2_127_3477_n477), .S(DP_OP_425J2_127_3477_n478) );
  FADDX1_HVT DP_OP_425J2_127_3477_U334 ( .A(DP_OP_425J2_127_3477_n1867), .B(
        DP_OP_425J2_127_3477_n2263), .CI(DP_OP_425J2_127_3477_n2050), .CO(
        DP_OP_425J2_127_3477_n475), .S(DP_OP_425J2_127_3477_n476) );
  FADDX1_HVT DP_OP_425J2_127_3477_U333 ( .A(DP_OP_425J2_127_3477_n2314), .B(
        DP_OP_425J2_127_3477_n1779), .CI(DP_OP_425J2_127_3477_n2399), .CO(
        DP_OP_425J2_127_3477_n473), .S(DP_OP_425J2_127_3477_n474) );
  FADDX1_HVT DP_OP_425J2_127_3477_U332 ( .A(DP_OP_425J2_127_3477_n2270), .B(
        DP_OP_425J2_127_3477_n2795), .CI(DP_OP_425J2_127_3477_n2182), .CO(
        DP_OP_425J2_127_3477_n471), .S(DP_OP_425J2_127_3477_n472) );
  FADDX1_HVT DP_OP_425J2_127_3477_U331 ( .A(DP_OP_425J2_127_3477_n2138), .B(
        DP_OP_425J2_127_3477_n2619), .CI(DP_OP_425J2_127_3477_n1918), .CO(
        DP_OP_425J2_127_3477_n469), .S(DP_OP_425J2_127_3477_n470) );
  FADDX1_HVT DP_OP_425J2_127_3477_U330 ( .A(DP_OP_425J2_127_3477_n2219), .B(
        DP_OP_425J2_127_3477_n1830), .CI(DP_OP_425J2_127_3477_n1874), .CO(
        DP_OP_425J2_127_3477_n467), .S(DP_OP_425J2_127_3477_n468) );
  FADDX1_HVT DP_OP_425J2_127_3477_U329 ( .A(DP_OP_425J2_127_3477_n2663), .B(
        DP_OP_425J2_127_3477_n2487), .CI(DP_OP_425J2_127_3477_n2355), .CO(
        DP_OP_425J2_127_3477_n465), .S(DP_OP_425J2_127_3477_n466) );
  FADDX1_HVT DP_OP_425J2_127_3477_U328 ( .A(DP_OP_425J2_127_3477_n2006), .B(
        DP_OP_425J2_127_3477_n669), .CI(DP_OP_425J2_127_3477_n667), .CO(
        DP_OP_425J2_127_3477_n463), .S(DP_OP_425J2_127_3477_n464) );
  FADDX1_HVT DP_OP_425J2_127_3477_U327 ( .A(DP_OP_425J2_127_3477_n665), .B(
        DP_OP_425J2_127_3477_n649), .CI(DP_OP_425J2_127_3477_n647), .CO(
        DP_OP_425J2_127_3477_n461), .S(DP_OP_425J2_127_3477_n462) );
  FADDX1_HVT DP_OP_425J2_127_3477_U326 ( .A(DP_OP_425J2_127_3477_n663), .B(
        DP_OP_425J2_127_3477_n651), .CI(DP_OP_425J2_127_3477_n653), .CO(
        DP_OP_425J2_127_3477_n459), .S(DP_OP_425J2_127_3477_n460) );
  FADDX1_HVT DP_OP_425J2_127_3477_U325 ( .A(DP_OP_425J2_127_3477_n661), .B(
        DP_OP_425J2_127_3477_n655), .CI(DP_OP_425J2_127_3477_n657), .CO(
        DP_OP_425J2_127_3477_n457), .S(DP_OP_425J2_127_3477_n458) );
  FADDX1_HVT DP_OP_425J2_127_3477_U324 ( .A(DP_OP_425J2_127_3477_n659), .B(
        DP_OP_425J2_127_3477_n645), .CI(DP_OP_425J2_127_3477_n643), .CO(
        DP_OP_425J2_127_3477_n455), .S(DP_OP_425J2_127_3477_n456) );
  FADDX1_HVT DP_OP_425J2_127_3477_U323 ( .A(DP_OP_425J2_127_3477_n641), .B(
        DP_OP_425J2_127_3477_n631), .CI(DP_OP_425J2_127_3477_n625), .CO(
        DP_OP_425J2_127_3477_n453), .S(DP_OP_425J2_127_3477_n454) );
  FADDX1_HVT DP_OP_425J2_127_3477_U322 ( .A(DP_OP_425J2_127_3477_n639), .B(
        DP_OP_425J2_127_3477_n633), .CI(DP_OP_425J2_127_3477_n627), .CO(
        DP_OP_425J2_127_3477_n451), .S(DP_OP_425J2_127_3477_n452) );
  FADDX1_HVT DP_OP_425J2_127_3477_U321 ( .A(DP_OP_425J2_127_3477_n637), .B(
        DP_OP_425J2_127_3477_n635), .CI(DP_OP_425J2_127_3477_n629), .CO(
        DP_OP_425J2_127_3477_n449), .S(DP_OP_425J2_127_3477_n450) );
  FADDX1_HVT DP_OP_425J2_127_3477_U320 ( .A(DP_OP_425J2_127_3477_n623), .B(
        DP_OP_425J2_127_3477_n490), .CI(DP_OP_425J2_127_3477_n476), .CO(
        DP_OP_425J2_127_3477_n447), .S(DP_OP_425J2_127_3477_n448) );
  FADDX1_HVT DP_OP_425J2_127_3477_U319 ( .A(DP_OP_425J2_127_3477_n621), .B(
        DP_OP_425J2_127_3477_n488), .CI(DP_OP_425J2_127_3477_n478), .CO(
        DP_OP_425J2_127_3477_n445), .S(DP_OP_425J2_127_3477_n446) );
  FADDX1_HVT DP_OP_425J2_127_3477_U318 ( .A(DP_OP_425J2_127_3477_n496), .B(
        DP_OP_425J2_127_3477_n480), .CI(DP_OP_425J2_127_3477_n486), .CO(
        DP_OP_425J2_127_3477_n443), .S(DP_OP_425J2_127_3477_n444) );
  FADDX1_HVT DP_OP_425J2_127_3477_U317 ( .A(DP_OP_425J2_127_3477_n498), .B(
        DP_OP_425J2_127_3477_n482), .CI(DP_OP_425J2_127_3477_n484), .CO(
        DP_OP_425J2_127_3477_n441), .S(DP_OP_425J2_127_3477_n442) );
  FADDX1_HVT DP_OP_425J2_127_3477_U316 ( .A(DP_OP_425J2_127_3477_n494), .B(
        DP_OP_425J2_127_3477_n492), .CI(DP_OP_425J2_127_3477_n474), .CO(
        DP_OP_425J2_127_3477_n439), .S(DP_OP_425J2_127_3477_n440) );
  FADDX1_HVT DP_OP_425J2_127_3477_U315 ( .A(DP_OP_425J2_127_3477_n472), .B(
        DP_OP_425J2_127_3477_n468), .CI(DP_OP_425J2_127_3477_n466), .CO(
        DP_OP_425J2_127_3477_n437), .S(DP_OP_425J2_127_3477_n438) );
  FADDX1_HVT DP_OP_425J2_127_3477_U314 ( .A(DP_OP_425J2_127_3477_n470), .B(
        DP_OP_425J2_127_3477_n619), .CI(DP_OP_425J2_127_3477_n617), .CO(
        DP_OP_425J2_127_3477_n435), .S(DP_OP_425J2_127_3477_n436) );
  FADDX1_HVT DP_OP_425J2_127_3477_U313 ( .A(DP_OP_425J2_127_3477_n615), .B(
        DP_OP_425J2_127_3477_n611), .CI(DP_OP_425J2_127_3477_n613), .CO(
        DP_OP_425J2_127_3477_n433), .S(DP_OP_425J2_127_3477_n434) );
  FADDX1_HVT DP_OP_425J2_127_3477_U312 ( .A(DP_OP_425J2_127_3477_n609), .B(
        DP_OP_425J2_127_3477_n603), .CI(DP_OP_425J2_127_3477_n601), .CO(
        DP_OP_425J2_127_3477_n431), .S(DP_OP_425J2_127_3477_n432) );
  FADDX1_HVT DP_OP_425J2_127_3477_U311 ( .A(DP_OP_425J2_127_3477_n607), .B(
        DP_OP_425J2_127_3477_n605), .CI(DP_OP_425J2_127_3477_n464), .CO(
        DP_OP_425J2_127_3477_n429), .S(DP_OP_425J2_127_3477_n430) );
  FADDX1_HVT DP_OP_425J2_127_3477_U310 ( .A(DP_OP_425J2_127_3477_n599), .B(
        DP_OP_425J2_127_3477_n458), .CI(DP_OP_425J2_127_3477_n462), .CO(
        DP_OP_425J2_127_3477_n427), .S(DP_OP_425J2_127_3477_n428) );
  FADDX1_HVT DP_OP_425J2_127_3477_U309 ( .A(DP_OP_425J2_127_3477_n597), .B(
        DP_OP_425J2_127_3477_n589), .CI(DP_OP_425J2_127_3477_n460), .CO(
        DP_OP_425J2_127_3477_n425), .S(DP_OP_425J2_127_3477_n426) );
  FADDX1_HVT DP_OP_425J2_127_3477_U308 ( .A(DP_OP_425J2_127_3477_n595), .B(
        DP_OP_425J2_127_3477_n593), .CI(DP_OP_425J2_127_3477_n591), .CO(
        DP_OP_425J2_127_3477_n423), .S(DP_OP_425J2_127_3477_n424) );
  FADDX1_HVT DP_OP_425J2_127_3477_U307 ( .A(DP_OP_425J2_127_3477_n456), .B(
        DP_OP_425J2_127_3477_n587), .CI(DP_OP_425J2_127_3477_n450), .CO(
        DP_OP_425J2_127_3477_n421), .S(DP_OP_425J2_127_3477_n422) );
  FADDX1_HVT DP_OP_425J2_127_3477_U306 ( .A(DP_OP_425J2_127_3477_n585), .B(
        DP_OP_425J2_127_3477_n452), .CI(DP_OP_425J2_127_3477_n581), .CO(
        DP_OP_425J2_127_3477_n419), .S(DP_OP_425J2_127_3477_n420) );
  FADDX1_HVT DP_OP_425J2_127_3477_U305 ( .A(DP_OP_425J2_127_3477_n583), .B(
        DP_OP_425J2_127_3477_n454), .CI(DP_OP_425J2_127_3477_n448), .CO(
        DP_OP_425J2_127_3477_n417), .S(DP_OP_425J2_127_3477_n418) );
  FADDX1_HVT DP_OP_425J2_127_3477_U304 ( .A(DP_OP_425J2_127_3477_n446), .B(
        DP_OP_425J2_127_3477_n444), .CI(DP_OP_425J2_127_3477_n440), .CO(
        DP_OP_425J2_127_3477_n415), .S(DP_OP_425J2_127_3477_n416) );
  FADDX1_HVT DP_OP_425J2_127_3477_U303 ( .A(DP_OP_425J2_127_3477_n442), .B(
        DP_OP_425J2_127_3477_n438), .CI(DP_OP_425J2_127_3477_n579), .CO(
        DP_OP_425J2_127_3477_n413), .S(DP_OP_425J2_127_3477_n414) );
  FADDX1_HVT DP_OP_425J2_127_3477_U302 ( .A(DP_OP_425J2_127_3477_n577), .B(
        DP_OP_425J2_127_3477_n575), .CI(DP_OP_425J2_127_3477_n436), .CO(
        DP_OP_425J2_127_3477_n411), .S(DP_OP_425J2_127_3477_n412) );
  FADDX1_HVT DP_OP_425J2_127_3477_U301 ( .A(DP_OP_425J2_127_3477_n573), .B(
        DP_OP_425J2_127_3477_n567), .CI(DP_OP_425J2_127_3477_n434), .CO(
        DP_OP_425J2_127_3477_n409), .S(DP_OP_425J2_127_3477_n410) );
  FADDX1_HVT DP_OP_425J2_127_3477_U300 ( .A(DP_OP_425J2_127_3477_n571), .B(
        DP_OP_425J2_127_3477_n569), .CI(DP_OP_425J2_127_3477_n565), .CO(
        DP_OP_425J2_127_3477_n407), .S(DP_OP_425J2_127_3477_n408) );
  FADDX1_HVT DP_OP_425J2_127_3477_U299 ( .A(DP_OP_425J2_127_3477_n563), .B(
        DP_OP_425J2_127_3477_n432), .CI(DP_OP_425J2_127_3477_n430), .CO(
        DP_OP_425J2_127_3477_n405), .S(DP_OP_425J2_127_3477_n406) );
  FADDX1_HVT DP_OP_425J2_127_3477_U298 ( .A(DP_OP_425J2_127_3477_n561), .B(
        DP_OP_425J2_127_3477_n559), .CI(DP_OP_425J2_127_3477_n557), .CO(
        DP_OP_425J2_127_3477_n403), .S(DP_OP_425J2_127_3477_n404) );
  FADDX1_HVT DP_OP_425J2_127_3477_U297 ( .A(DP_OP_425J2_127_3477_n555), .B(
        DP_OP_425J2_127_3477_n426), .CI(DP_OP_425J2_127_3477_n424), .CO(
        DP_OP_425J2_127_3477_n401), .S(DP_OP_425J2_127_3477_n402) );
  FADDX1_HVT DP_OP_425J2_127_3477_U296 ( .A(DP_OP_425J2_127_3477_n428), .B(
        DP_OP_425J2_127_3477_n422), .CI(DP_OP_425J2_127_3477_n553), .CO(
        DP_OP_425J2_127_3477_n399), .S(DP_OP_425J2_127_3477_n400) );
  FADDX1_HVT DP_OP_425J2_127_3477_U295 ( .A(DP_OP_425J2_127_3477_n420), .B(
        DP_OP_425J2_127_3477_n551), .CI(DP_OP_425J2_127_3477_n418), .CO(
        DP_OP_425J2_127_3477_n397), .S(DP_OP_425J2_127_3477_n398) );
  FADDX1_HVT DP_OP_425J2_127_3477_U294 ( .A(DP_OP_425J2_127_3477_n416), .B(
        DP_OP_425J2_127_3477_n549), .CI(DP_OP_425J2_127_3477_n414), .CO(
        DP_OP_425J2_127_3477_n395), .S(DP_OP_425J2_127_3477_n396) );
  FADDX1_HVT DP_OP_425J2_127_3477_U293 ( .A(DP_OP_425J2_127_3477_n547), .B(
        DP_OP_425J2_127_3477_n545), .CI(DP_OP_425J2_127_3477_n412), .CO(
        DP_OP_425J2_127_3477_n393), .S(DP_OP_425J2_127_3477_n394) );
  FADDX1_HVT DP_OP_425J2_127_3477_U292 ( .A(DP_OP_425J2_127_3477_n543), .B(
        DP_OP_425J2_127_3477_n410), .CI(DP_OP_425J2_127_3477_n539), .CO(
        DP_OP_425J2_127_3477_n391), .S(DP_OP_425J2_127_3477_n392) );
  FADDX1_HVT DP_OP_425J2_127_3477_U291 ( .A(DP_OP_425J2_127_3477_n541), .B(
        DP_OP_425J2_127_3477_n408), .CI(DP_OP_425J2_127_3477_n537), .CO(
        DP_OP_425J2_127_3477_n389), .S(DP_OP_425J2_127_3477_n390) );
  FADDX1_HVT DP_OP_425J2_127_3477_U290 ( .A(DP_OP_425J2_127_3477_n406), .B(
        DP_OP_425J2_127_3477_n535), .CI(DP_OP_425J2_127_3477_n404), .CO(
        DP_OP_425J2_127_3477_n387), .S(DP_OP_425J2_127_3477_n388) );
  FADDX1_HVT DP_OP_425J2_127_3477_U289 ( .A(DP_OP_425J2_127_3477_n533), .B(
        DP_OP_425J2_127_3477_n402), .CI(DP_OP_425J2_127_3477_n400), .CO(
        DP_OP_425J2_127_3477_n385), .S(DP_OP_425J2_127_3477_n386) );
  FADDX1_HVT DP_OP_425J2_127_3477_U288 ( .A(DP_OP_425J2_127_3477_n531), .B(
        DP_OP_425J2_127_3477_n398), .CI(DP_OP_425J2_127_3477_n529), .CO(
        DP_OP_425J2_127_3477_n383), .S(DP_OP_425J2_127_3477_n384) );
  FADDX1_HVT DP_OP_425J2_127_3477_U287 ( .A(DP_OP_425J2_127_3477_n396), .B(
        DP_OP_425J2_127_3477_n527), .CI(DP_OP_425J2_127_3477_n394), .CO(
        DP_OP_425J2_127_3477_n381), .S(DP_OP_425J2_127_3477_n382) );
  FADDX1_HVT DP_OP_425J2_127_3477_U286 ( .A(DP_OP_425J2_127_3477_n525), .B(
        DP_OP_425J2_127_3477_n523), .CI(DP_OP_425J2_127_3477_n392), .CO(
        DP_OP_425J2_127_3477_n379), .S(DP_OP_425J2_127_3477_n380) );
  FADDX1_HVT DP_OP_425J2_127_3477_U285 ( .A(DP_OP_425J2_127_3477_n390), .B(
        DP_OP_425J2_127_3477_n521), .CI(DP_OP_425J2_127_3477_n388), .CO(
        DP_OP_425J2_127_3477_n377), .S(DP_OP_425J2_127_3477_n378) );
  FADDX1_HVT DP_OP_425J2_127_3477_U284 ( .A(DP_OP_425J2_127_3477_n519), .B(
        DP_OP_425J2_127_3477_n386), .CI(DP_OP_425J2_127_3477_n517), .CO(
        DP_OP_425J2_127_3477_n375), .S(DP_OP_425J2_127_3477_n376) );
  FADDX1_HVT DP_OP_425J2_127_3477_U283 ( .A(DP_OP_425J2_127_3477_n384), .B(
        DP_OP_425J2_127_3477_n515), .CI(DP_OP_425J2_127_3477_n382), .CO(
        DP_OP_425J2_127_3477_n373), .S(DP_OP_425J2_127_3477_n374) );
  FADDX1_HVT DP_OP_425J2_127_3477_U282 ( .A(DP_OP_425J2_127_3477_n513), .B(
        DP_OP_425J2_127_3477_n380), .CI(DP_OP_425J2_127_3477_n511), .CO(
        DP_OP_425J2_127_3477_n371), .S(DP_OP_425J2_127_3477_n372) );
  FADDX1_HVT DP_OP_425J2_127_3477_U281 ( .A(DP_OP_425J2_127_3477_n378), .B(
        DP_OP_425J2_127_3477_n509), .CI(DP_OP_425J2_127_3477_n376), .CO(
        DP_OP_425J2_127_3477_n369), .S(DP_OP_425J2_127_3477_n370) );
  FADDX1_HVT DP_OP_425J2_127_3477_U280 ( .A(DP_OP_425J2_127_3477_n507), .B(
        DP_OP_425J2_127_3477_n374), .CI(DP_OP_425J2_127_3477_n505), .CO(
        DP_OP_425J2_127_3477_n367), .S(DP_OP_425J2_127_3477_n368) );
  FADDX1_HVT DP_OP_425J2_127_3477_U279 ( .A(DP_OP_425J2_127_3477_n372), .B(
        DP_OP_425J2_127_3477_n370), .CI(DP_OP_425J2_127_3477_n503), .CO(
        DP_OP_425J2_127_3477_n365), .S(DP_OP_425J2_127_3477_n366) );
  FADDX1_HVT DP_OP_425J2_127_3477_U278 ( .A(DP_OP_425J2_127_3477_n501), .B(
        DP_OP_425J2_127_3477_n368), .CI(DP_OP_425J2_127_3477_n366), .CO(
        DP_OP_425J2_127_3477_n363), .S(DP_OP_425J2_127_3477_n364) );
  FADDX1_HVT DP_OP_425J2_127_3477_U276 ( .A(DP_OP_425J2_127_3477_n2699), .B(
        DP_OP_425J2_127_3477_n1822), .CI(DP_OP_425J2_127_3477_n2391), .CO(
        DP_OP_425J2_127_3477_n359), .S(DP_OP_425J2_127_3477_n360) );
  FADDX1_HVT DP_OP_425J2_127_3477_U275 ( .A(DP_OP_425J2_127_3477_n1998), .B(
        DP_OP_425J2_127_3477_n1778), .CI(DP_OP_425J2_127_3477_n1954), .CO(
        DP_OP_425J2_127_3477_n357), .S(DP_OP_425J2_127_3477_n358) );
  FADDX1_HVT DP_OP_425J2_127_3477_U274 ( .A(DP_OP_425J2_127_3477_n1866), .B(
        DP_OP_425J2_127_3477_n2567), .CI(DP_OP_425J2_127_3477_n2743), .CO(
        DP_OP_425J2_127_3477_n355), .S(DP_OP_425J2_127_3477_n356) );
  FADDX1_HVT DP_OP_425J2_127_3477_U273 ( .A(DP_OP_425J2_127_3477_n2611), .B(
        DP_OP_425J2_127_3477_n1910), .CI(DP_OP_425J2_127_3477_n2042), .CO(
        DP_OP_425J2_127_3477_n353), .S(DP_OP_425J2_127_3477_n354) );
  FADDX1_HVT DP_OP_425J2_127_3477_U272 ( .A(DP_OP_425J2_127_3477_n2086), .B(
        DP_OP_425J2_127_3477_n2174), .CI(DP_OP_425J2_127_3477_n2435), .CO(
        DP_OP_425J2_127_3477_n351), .S(DP_OP_425J2_127_3477_n352) );
  FADDX1_HVT DP_OP_425J2_127_3477_U271 ( .A(DP_OP_425J2_127_3477_n2130), .B(
        DP_OP_425J2_127_3477_n2479), .CI(DP_OP_425J2_127_3477_n2523), .CO(
        DP_OP_425J2_127_3477_n349), .S(DP_OP_425J2_127_3477_n350) );
  FADDX1_HVT DP_OP_425J2_127_3477_U270 ( .A(DP_OP_425J2_127_3477_n2306), .B(
        DP_OP_425J2_127_3477_n2262), .CI(DP_OP_425J2_127_3477_n2875), .CO(
        DP_OP_425J2_127_3477_n347), .S(DP_OP_425J2_127_3477_n348) );
  FADDX1_HVT DP_OP_425J2_127_3477_U269 ( .A(DP_OP_425J2_127_3477_n2787), .B(
        DP_OP_425J2_127_3477_n2831), .CI(DP_OP_425J2_127_3477_n2655), .CO(
        DP_OP_425J2_127_3477_n345), .S(DP_OP_425J2_127_3477_n346) );
  FADDX1_HVT DP_OP_425J2_127_3477_U268 ( .A(DP_OP_425J2_127_3477_n362), .B(
        DP_OP_425J2_127_3477_n2218), .CI(DP_OP_425J2_127_3477_n497), .CO(
        DP_OP_425J2_127_3477_n343), .S(DP_OP_425J2_127_3477_n344) );
  FADDX1_HVT DP_OP_425J2_127_3477_U267 ( .A(DP_OP_425J2_127_3477_n495), .B(
        DP_OP_425J2_127_3477_n477), .CI(DP_OP_425J2_127_3477_n475), .CO(
        DP_OP_425J2_127_3477_n341), .S(DP_OP_425J2_127_3477_n342) );
  FADDX1_HVT DP_OP_425J2_127_3477_U266 ( .A(DP_OP_425J2_127_3477_n493), .B(
        DP_OP_425J2_127_3477_n479), .CI(DP_OP_425J2_127_3477_n481), .CO(
        DP_OP_425J2_127_3477_n339), .S(DP_OP_425J2_127_3477_n340) );
  FADDX1_HVT DP_OP_425J2_127_3477_U265 ( .A(DP_OP_425J2_127_3477_n491), .B(
        DP_OP_425J2_127_3477_n483), .CI(DP_OP_425J2_127_3477_n485), .CO(
        DP_OP_425J2_127_3477_n337), .S(DP_OP_425J2_127_3477_n338) );
  FADDX1_HVT DP_OP_425J2_127_3477_U264 ( .A(DP_OP_425J2_127_3477_n489), .B(
        DP_OP_425J2_127_3477_n487), .CI(DP_OP_425J2_127_3477_n473), .CO(
        DP_OP_425J2_127_3477_n335), .S(DP_OP_425J2_127_3477_n336) );
  FADDX1_HVT DP_OP_425J2_127_3477_U263 ( .A(DP_OP_425J2_127_3477_n471), .B(
        DP_OP_425J2_127_3477_n467), .CI(DP_OP_425J2_127_3477_n465), .CO(
        DP_OP_425J2_127_3477_n333), .S(DP_OP_425J2_127_3477_n334) );
  FADDX1_HVT DP_OP_425J2_127_3477_U262 ( .A(DP_OP_425J2_127_3477_n469), .B(
        DP_OP_425J2_127_3477_n358), .CI(DP_OP_425J2_127_3477_n360), .CO(
        DP_OP_425J2_127_3477_n331), .S(DP_OP_425J2_127_3477_n332) );
  FADDX1_HVT DP_OP_425J2_127_3477_U261 ( .A(DP_OP_425J2_127_3477_n352), .B(
        DP_OP_425J2_127_3477_n346), .CI(DP_OP_425J2_127_3477_n348), .CO(
        DP_OP_425J2_127_3477_n329), .S(DP_OP_425J2_127_3477_n330) );
  FADDX1_HVT DP_OP_425J2_127_3477_U260 ( .A(DP_OP_425J2_127_3477_n350), .B(
        DP_OP_425J2_127_3477_n356), .CI(DP_OP_425J2_127_3477_n354), .CO(
        DP_OP_425J2_127_3477_n327), .S(DP_OP_425J2_127_3477_n328) );
  FADDX1_HVT DP_OP_425J2_127_3477_U259 ( .A(DP_OP_425J2_127_3477_n463), .B(
        DP_OP_425J2_127_3477_n461), .CI(DP_OP_425J2_127_3477_n457), .CO(
        DP_OP_425J2_127_3477_n325), .S(DP_OP_425J2_127_3477_n326) );
  FADDX1_HVT DP_OP_425J2_127_3477_U258 ( .A(DP_OP_425J2_127_3477_n459), .B(
        DP_OP_425J2_127_3477_n455), .CI(DP_OP_425J2_127_3477_n453), .CO(
        DP_OP_425J2_127_3477_n323), .S(DP_OP_425J2_127_3477_n324) );
  FADDX1_HVT DP_OP_425J2_127_3477_U257 ( .A(DP_OP_425J2_127_3477_n451), .B(
        DP_OP_425J2_127_3477_n449), .CI(DP_OP_425J2_127_3477_n344), .CO(
        DP_OP_425J2_127_3477_n321), .S(DP_OP_425J2_127_3477_n322) );
  FADDX1_HVT DP_OP_425J2_127_3477_U256 ( .A(DP_OP_425J2_127_3477_n447), .B(
        DP_OP_425J2_127_3477_n439), .CI(DP_OP_425J2_127_3477_n336), .CO(
        DP_OP_425J2_127_3477_n319), .S(DP_OP_425J2_127_3477_n320) );
  FADDX1_HVT DP_OP_425J2_127_3477_U255 ( .A(DP_OP_425J2_127_3477_n445), .B(
        DP_OP_425J2_127_3477_n338), .CI(DP_OP_425J2_127_3477_n340), .CO(
        DP_OP_425J2_127_3477_n317), .S(DP_OP_425J2_127_3477_n318) );
  FADDX1_HVT DP_OP_425J2_127_3477_U254 ( .A(DP_OP_425J2_127_3477_n443), .B(
        DP_OP_425J2_127_3477_n441), .CI(DP_OP_425J2_127_3477_n342), .CO(
        DP_OP_425J2_127_3477_n315), .S(DP_OP_425J2_127_3477_n316) );
  FADDX1_HVT DP_OP_425J2_127_3477_U253 ( .A(DP_OP_425J2_127_3477_n437), .B(
        DP_OP_425J2_127_3477_n334), .CI(DP_OP_425J2_127_3477_n435), .CO(
        DP_OP_425J2_127_3477_n313), .S(DP_OP_425J2_127_3477_n314) );
  FADDX1_HVT DP_OP_425J2_127_3477_U252 ( .A(DP_OP_425J2_127_3477_n332), .B(
        DP_OP_425J2_127_3477_n328), .CI(DP_OP_425J2_127_3477_n433), .CO(
        DP_OP_425J2_127_3477_n311), .S(DP_OP_425J2_127_3477_n312) );
  FADDX1_HVT DP_OP_425J2_127_3477_U251 ( .A(DP_OP_425J2_127_3477_n330), .B(
        DP_OP_425J2_127_3477_n431), .CI(DP_OP_425J2_127_3477_n429), .CO(
        DP_OP_425J2_127_3477_n309), .S(DP_OP_425J2_127_3477_n310) );
  FADDX1_HVT DP_OP_425J2_127_3477_U250 ( .A(DP_OP_425J2_127_3477_n326), .B(
        DP_OP_425J2_127_3477_n423), .CI(DP_OP_425J2_127_3477_n324), .CO(
        DP_OP_425J2_127_3477_n307), .S(DP_OP_425J2_127_3477_n308) );
  FADDX1_HVT DP_OP_425J2_127_3477_U249 ( .A(DP_OP_425J2_127_3477_n427), .B(
        DP_OP_425J2_127_3477_n425), .CI(DP_OP_425J2_127_3477_n421), .CO(
        DP_OP_425J2_127_3477_n305), .S(DP_OP_425J2_127_3477_n306) );
  FADDX1_HVT DP_OP_425J2_127_3477_U248 ( .A(DP_OP_425J2_127_3477_n419), .B(
        DP_OP_425J2_127_3477_n322), .CI(DP_OP_425J2_127_3477_n417), .CO(
        DP_OP_425J2_127_3477_n303), .S(DP_OP_425J2_127_3477_n304) );
  FADDX1_HVT DP_OP_425J2_127_3477_U247 ( .A(DP_OP_425J2_127_3477_n320), .B(
        DP_OP_425J2_127_3477_n316), .CI(DP_OP_425J2_127_3477_n413), .CO(
        DP_OP_425J2_127_3477_n301), .S(DP_OP_425J2_127_3477_n302) );
  FADDX1_HVT DP_OP_425J2_127_3477_U246 ( .A(DP_OP_425J2_127_3477_n415), .B(
        DP_OP_425J2_127_3477_n318), .CI(DP_OP_425J2_127_3477_n314), .CO(
        DP_OP_425J2_127_3477_n299), .S(DP_OP_425J2_127_3477_n300) );
  FADDX1_HVT DP_OP_425J2_127_3477_U245 ( .A(DP_OP_425J2_127_3477_n411), .B(
        DP_OP_425J2_127_3477_n312), .CI(DP_OP_425J2_127_3477_n409), .CO(
        DP_OP_425J2_127_3477_n297), .S(DP_OP_425J2_127_3477_n298) );
  FADDX1_HVT DP_OP_425J2_127_3477_U244 ( .A(DP_OP_425J2_127_3477_n407), .B(
        DP_OP_425J2_127_3477_n310), .CI(DP_OP_425J2_127_3477_n405), .CO(
        DP_OP_425J2_127_3477_n295), .S(DP_OP_425J2_127_3477_n296) );
  FADDX1_HVT DP_OP_425J2_127_3477_U243 ( .A(DP_OP_425J2_127_3477_n403), .B(
        DP_OP_425J2_127_3477_n308), .CI(DP_OP_425J2_127_3477_n306), .CO(
        DP_OP_425J2_127_3477_n293), .S(DP_OP_425J2_127_3477_n294) );
  FADDX1_HVT DP_OP_425J2_127_3477_U242 ( .A(DP_OP_425J2_127_3477_n401), .B(
        DP_OP_425J2_127_3477_n399), .CI(DP_OP_425J2_127_3477_n304), .CO(
        DP_OP_425J2_127_3477_n291), .S(DP_OP_425J2_127_3477_n292) );
  FADDX1_HVT DP_OP_425J2_127_3477_U241 ( .A(DP_OP_425J2_127_3477_n397), .B(
        DP_OP_425J2_127_3477_n302), .CI(DP_OP_425J2_127_3477_n395), .CO(
        DP_OP_425J2_127_3477_n289), .S(DP_OP_425J2_127_3477_n290) );
  FADDX1_HVT DP_OP_425J2_127_3477_U240 ( .A(DP_OP_425J2_127_3477_n300), .B(
        DP_OP_425J2_127_3477_n393), .CI(DP_OP_425J2_127_3477_n391), .CO(
        DP_OP_425J2_127_3477_n287), .S(DP_OP_425J2_127_3477_n288) );
  FADDX1_HVT DP_OP_425J2_127_3477_U239 ( .A(DP_OP_425J2_127_3477_n298), .B(
        DP_OP_425J2_127_3477_n389), .CI(DP_OP_425J2_127_3477_n296), .CO(
        DP_OP_425J2_127_3477_n285), .S(DP_OP_425J2_127_3477_n286) );
  FADDX1_HVT DP_OP_425J2_127_3477_U238 ( .A(DP_OP_425J2_127_3477_n387), .B(
        DP_OP_425J2_127_3477_n294), .CI(DP_OP_425J2_127_3477_n385), .CO(
        DP_OP_425J2_127_3477_n283), .S(DP_OP_425J2_127_3477_n284) );
  FADDX1_HVT DP_OP_425J2_127_3477_U237 ( .A(DP_OP_425J2_127_3477_n292), .B(
        DP_OP_425J2_127_3477_n383), .CI(DP_OP_425J2_127_3477_n290), .CO(
        DP_OP_425J2_127_3477_n281), .S(DP_OP_425J2_127_3477_n282) );
  FADDX1_HVT DP_OP_425J2_127_3477_U236 ( .A(DP_OP_425J2_127_3477_n381), .B(
        DP_OP_425J2_127_3477_n288), .CI(DP_OP_425J2_127_3477_n379), .CO(
        DP_OP_425J2_127_3477_n279), .S(DP_OP_425J2_127_3477_n280) );
  FADDX1_HVT DP_OP_425J2_127_3477_U235 ( .A(DP_OP_425J2_127_3477_n286), .B(
        DP_OP_425J2_127_3477_n377), .CI(DP_OP_425J2_127_3477_n284), .CO(
        DP_OP_425J2_127_3477_n277), .S(DP_OP_425J2_127_3477_n278) );
  FADDX1_HVT DP_OP_425J2_127_3477_U234 ( .A(DP_OP_425J2_127_3477_n375), .B(
        DP_OP_425J2_127_3477_n282), .CI(DP_OP_425J2_127_3477_n373), .CO(
        DP_OP_425J2_127_3477_n275), .S(DP_OP_425J2_127_3477_n276) );
  FADDX1_HVT DP_OP_425J2_127_3477_U233 ( .A(DP_OP_425J2_127_3477_n280), .B(
        DP_OP_425J2_127_3477_n371), .CI(DP_OP_425J2_127_3477_n278), .CO(
        DP_OP_425J2_127_3477_n273), .S(DP_OP_425J2_127_3477_n274) );
  FADDX1_HVT DP_OP_425J2_127_3477_U232 ( .A(DP_OP_425J2_127_3477_n369), .B(
        DP_OP_425J2_127_3477_n276), .CI(DP_OP_425J2_127_3477_n367), .CO(
        DP_OP_425J2_127_3477_n271), .S(DP_OP_425J2_127_3477_n272) );
  FADDX1_HVT DP_OP_425J2_127_3477_U231 ( .A(DP_OP_425J2_127_3477_n274), .B(
        DP_OP_425J2_127_3477_n365), .CI(DP_OP_425J2_127_3477_n272), .CO(
        DP_OP_425J2_127_3477_n269), .S(DP_OP_425J2_127_3477_n270) );
  FADDX1_HVT DP_OP_425J2_127_3477_U230 ( .A(DP_OP_425J2_127_3477_n361), .B(
        DP_OP_425J2_127_3477_n1777), .CI(DP_OP_425J2_127_3477_n359), .CO(
        DP_OP_425J2_127_3477_n267), .S(DP_OP_425J2_127_3477_n268) );
  FADDX1_HVT DP_OP_425J2_127_3477_U229 ( .A(DP_OP_425J2_127_3477_n357), .B(
        DP_OP_425J2_127_3477_n345), .CI(DP_OP_425J2_127_3477_n355), .CO(
        DP_OP_425J2_127_3477_n265), .S(DP_OP_425J2_127_3477_n266) );
  FADDX1_HVT DP_OP_425J2_127_3477_U228 ( .A(DP_OP_425J2_127_3477_n353), .B(
        DP_OP_425J2_127_3477_n351), .CI(DP_OP_425J2_127_3477_n349), .CO(
        DP_OP_425J2_127_3477_n263), .S(DP_OP_425J2_127_3477_n264) );
  FADDX1_HVT DP_OP_425J2_127_3477_U227 ( .A(DP_OP_425J2_127_3477_n347), .B(
        DP_OP_425J2_127_3477_n343), .CI(DP_OP_425J2_127_3477_n341), .CO(
        DP_OP_425J2_127_3477_n261), .S(DP_OP_425J2_127_3477_n262) );
  FADDX1_HVT DP_OP_425J2_127_3477_U226 ( .A(DP_OP_425J2_127_3477_n339), .B(
        DP_OP_425J2_127_3477_n337), .CI(DP_OP_425J2_127_3477_n335), .CO(
        DP_OP_425J2_127_3477_n259), .S(DP_OP_425J2_127_3477_n260) );
  FADDX1_HVT DP_OP_425J2_127_3477_U225 ( .A(DP_OP_425J2_127_3477_n333), .B(
        DP_OP_425J2_127_3477_n268), .CI(DP_OP_425J2_127_3477_n331), .CO(
        DP_OP_425J2_127_3477_n257), .S(DP_OP_425J2_127_3477_n258) );
  FADDX1_HVT DP_OP_425J2_127_3477_U224 ( .A(DP_OP_425J2_127_3477_n266), .B(
        DP_OP_425J2_127_3477_n264), .CI(DP_OP_425J2_127_3477_n327), .CO(
        DP_OP_425J2_127_3477_n255), .S(DP_OP_425J2_127_3477_n256) );
  FADDX1_HVT DP_OP_425J2_127_3477_U223 ( .A(DP_OP_425J2_127_3477_n329), .B(
        DP_OP_425J2_127_3477_n325), .CI(DP_OP_425J2_127_3477_n323), .CO(
        DP_OP_425J2_127_3477_n253), .S(DP_OP_425J2_127_3477_n254) );
  FADDX1_HVT DP_OP_425J2_127_3477_U222 ( .A(DP_OP_425J2_127_3477_n321), .B(
        DP_OP_425J2_127_3477_n262), .CI(DP_OP_425J2_127_3477_n319), .CO(
        DP_OP_425J2_127_3477_n251), .S(DP_OP_425J2_127_3477_n252) );
  FADDX1_HVT DP_OP_425J2_127_3477_U221 ( .A(DP_OP_425J2_127_3477_n317), .B(
        DP_OP_425J2_127_3477_n315), .CI(DP_OP_425J2_127_3477_n260), .CO(
        DP_OP_425J2_127_3477_n249), .S(DP_OP_425J2_127_3477_n250) );
  FADDX1_HVT DP_OP_425J2_127_3477_U220 ( .A(DP_OP_425J2_127_3477_n313), .B(
        DP_OP_425J2_127_3477_n258), .CI(DP_OP_425J2_127_3477_n311), .CO(
        DP_OP_425J2_127_3477_n247), .S(DP_OP_425J2_127_3477_n248) );
  FADDX1_HVT DP_OP_425J2_127_3477_U219 ( .A(DP_OP_425J2_127_3477_n256), .B(
        DP_OP_425J2_127_3477_n309), .CI(DP_OP_425J2_127_3477_n254), .CO(
        DP_OP_425J2_127_3477_n245), .S(DP_OP_425J2_127_3477_n246) );
  FADDX1_HVT DP_OP_425J2_127_3477_U218 ( .A(DP_OP_425J2_127_3477_n307), .B(
        DP_OP_425J2_127_3477_n305), .CI(DP_OP_425J2_127_3477_n303), .CO(
        DP_OP_425J2_127_3477_n243), .S(DP_OP_425J2_127_3477_n244) );
  FADDX1_HVT DP_OP_425J2_127_3477_U217 ( .A(DP_OP_425J2_127_3477_n252), .B(
        DP_OP_425J2_127_3477_n301), .CI(DP_OP_425J2_127_3477_n250), .CO(
        DP_OP_425J2_127_3477_n241), .S(DP_OP_425J2_127_3477_n242) );
  FADDX1_HVT DP_OP_425J2_127_3477_U216 ( .A(DP_OP_425J2_127_3477_n299), .B(
        DP_OP_425J2_127_3477_n248), .CI(DP_OP_425J2_127_3477_n297), .CO(
        DP_OP_425J2_127_3477_n239), .S(DP_OP_425J2_127_3477_n240) );
  FADDX1_HVT DP_OP_425J2_127_3477_U215 ( .A(DP_OP_425J2_127_3477_n295), .B(
        DP_OP_425J2_127_3477_n246), .CI(DP_OP_425J2_127_3477_n293), .CO(
        DP_OP_425J2_127_3477_n237), .S(DP_OP_425J2_127_3477_n238) );
  FADDX1_HVT DP_OP_425J2_127_3477_U214 ( .A(DP_OP_425J2_127_3477_n291), .B(
        DP_OP_425J2_127_3477_n244), .CI(DP_OP_425J2_127_3477_n289), .CO(
        DP_OP_425J2_127_3477_n235), .S(DP_OP_425J2_127_3477_n236) );
  FADDX1_HVT DP_OP_425J2_127_3477_U213 ( .A(DP_OP_425J2_127_3477_n242), .B(
        DP_OP_425J2_127_3477_n287), .CI(DP_OP_425J2_127_3477_n240), .CO(
        DP_OP_425J2_127_3477_n233), .S(DP_OP_425J2_127_3477_n234) );
  FADDX1_HVT DP_OP_425J2_127_3477_U212 ( .A(DP_OP_425J2_127_3477_n285), .B(
        DP_OP_425J2_127_3477_n238), .CI(DP_OP_425J2_127_3477_n283), .CO(
        DP_OP_425J2_127_3477_n231), .S(DP_OP_425J2_127_3477_n232) );
  FADDX1_HVT DP_OP_425J2_127_3477_U211 ( .A(DP_OP_425J2_127_3477_n281), .B(
        DP_OP_425J2_127_3477_n236), .CI(DP_OP_425J2_127_3477_n234), .CO(
        DP_OP_425J2_127_3477_n229), .S(DP_OP_425J2_127_3477_n230) );
  FADDX1_HVT DP_OP_425J2_127_3477_U210 ( .A(DP_OP_425J2_127_3477_n279), .B(
        DP_OP_425J2_127_3477_n277), .CI(DP_OP_425J2_127_3477_n232), .CO(
        DP_OP_425J2_127_3477_n227), .S(DP_OP_425J2_127_3477_n228) );
  FADDX1_HVT DP_OP_425J2_127_3477_U209 ( .A(DP_OP_425J2_127_3477_n275), .B(
        DP_OP_425J2_127_3477_n230), .CI(DP_OP_425J2_127_3477_n273), .CO(
        DP_OP_425J2_127_3477_n225), .S(DP_OP_425J2_127_3477_n226) );
  FADDX1_HVT DP_OP_425J2_127_3477_U208 ( .A(DP_OP_425J2_127_3477_n228), .B(
        DP_OP_425J2_127_3477_n271), .CI(DP_OP_425J2_127_3477_n226), .CO(
        DP_OP_425J2_127_3477_n223), .S(DP_OP_425J2_127_3477_n224) );
  FADDX1_HVT DP_OP_425J2_127_3477_U207 ( .A(DP_OP_425J2_127_3477_n1776), .B(
        DP_OP_425J2_127_3477_n267), .CI(DP_OP_425J2_127_3477_n265), .CO(
        DP_OP_425J2_127_3477_n221), .S(DP_OP_425J2_127_3477_n222) );
  FADDX1_HVT DP_OP_425J2_127_3477_U206 ( .A(DP_OP_425J2_127_3477_n263), .B(
        DP_OP_425J2_127_3477_n261), .CI(DP_OP_425J2_127_3477_n259), .CO(
        DP_OP_425J2_127_3477_n219), .S(DP_OP_425J2_127_3477_n220) );
  FADDX1_HVT DP_OP_425J2_127_3477_U205 ( .A(DP_OP_425J2_127_3477_n257), .B(
        DP_OP_425J2_127_3477_n222), .CI(DP_OP_425J2_127_3477_n255), .CO(
        DP_OP_425J2_127_3477_n217), .S(DP_OP_425J2_127_3477_n218) );
  FADDX1_HVT DP_OP_425J2_127_3477_U204 ( .A(DP_OP_425J2_127_3477_n253), .B(
        DP_OP_425J2_127_3477_n251), .CI(DP_OP_425J2_127_3477_n220), .CO(
        DP_OP_425J2_127_3477_n215), .S(DP_OP_425J2_127_3477_n216) );
  FADDX1_HVT DP_OP_425J2_127_3477_U203 ( .A(DP_OP_425J2_127_3477_n249), .B(
        DP_OP_425J2_127_3477_n247), .CI(DP_OP_425J2_127_3477_n218), .CO(
        DP_OP_425J2_127_3477_n213), .S(DP_OP_425J2_127_3477_n214) );
  FADDX1_HVT DP_OP_425J2_127_3477_U202 ( .A(DP_OP_425J2_127_3477_n245), .B(
        DP_OP_425J2_127_3477_n243), .CI(DP_OP_425J2_127_3477_n216), .CO(
        DP_OP_425J2_127_3477_n211), .S(DP_OP_425J2_127_3477_n212) );
  FADDX1_HVT DP_OP_425J2_127_3477_U201 ( .A(DP_OP_425J2_127_3477_n241), .B(
        DP_OP_425J2_127_3477_n214), .CI(DP_OP_425J2_127_3477_n239), .CO(
        DP_OP_425J2_127_3477_n209), .S(DP_OP_425J2_127_3477_n210) );
  FADDX1_HVT DP_OP_425J2_127_3477_U200 ( .A(DP_OP_425J2_127_3477_n237), .B(
        DP_OP_425J2_127_3477_n212), .CI(DP_OP_425J2_127_3477_n235), .CO(
        DP_OP_425J2_127_3477_n207), .S(DP_OP_425J2_127_3477_n208) );
  FADDX1_HVT DP_OP_425J2_127_3477_U199 ( .A(DP_OP_425J2_127_3477_n233), .B(
        DP_OP_425J2_127_3477_n210), .CI(DP_OP_425J2_127_3477_n231), .CO(
        DP_OP_425J2_127_3477_n205), .S(DP_OP_425J2_127_3477_n206) );
  FADDX1_HVT DP_OP_425J2_127_3477_U198 ( .A(DP_OP_425J2_127_3477_n208), .B(
        DP_OP_425J2_127_3477_n229), .CI(DP_OP_425J2_127_3477_n206), .CO(
        DP_OP_425J2_127_3477_n203), .S(DP_OP_425J2_127_3477_n204) );
  FADDX1_HVT DP_OP_425J2_127_3477_U197 ( .A(DP_OP_425J2_127_3477_n227), .B(
        DP_OP_425J2_127_3477_n225), .CI(DP_OP_425J2_127_3477_n204), .CO(
        DP_OP_425J2_127_3477_n201), .S(DP_OP_425J2_127_3477_n202) );
  FADDX1_HVT DP_OP_425J2_127_3477_U196 ( .A(DP_OP_425J2_127_3477_n1775), .B(
        DP_OP_425J2_127_3477_n221), .CI(DP_OP_425J2_127_3477_n219), .CO(
        DP_OP_425J2_127_3477_n199), .S(DP_OP_425J2_127_3477_n200) );
  FADDX1_HVT DP_OP_425J2_127_3477_U195 ( .A(DP_OP_425J2_127_3477_n217), .B(
        DP_OP_425J2_127_3477_n200), .CI(DP_OP_425J2_127_3477_n215), .CO(
        DP_OP_425J2_127_3477_n197), .S(DP_OP_425J2_127_3477_n198) );
  FADDX1_HVT DP_OP_425J2_127_3477_U194 ( .A(DP_OP_425J2_127_3477_n213), .B(
        DP_OP_425J2_127_3477_n211), .CI(DP_OP_425J2_127_3477_n198), .CO(
        DP_OP_425J2_127_3477_n195), .S(DP_OP_425J2_127_3477_n196) );
  FADDX1_HVT DP_OP_425J2_127_3477_U193 ( .A(DP_OP_425J2_127_3477_n209), .B(
        DP_OP_425J2_127_3477_n196), .CI(DP_OP_425J2_127_3477_n207), .CO(
        DP_OP_425J2_127_3477_n193), .S(DP_OP_425J2_127_3477_n194) );
  FADDX1_HVT DP_OP_425J2_127_3477_U192 ( .A(DP_OP_425J2_127_3477_n205), .B(
        DP_OP_425J2_127_3477_n194), .CI(DP_OP_425J2_127_3477_n203), .CO(
        DP_OP_425J2_127_3477_n191), .S(DP_OP_425J2_127_3477_n192) );
  FADDX1_HVT DP_OP_425J2_127_3477_U190 ( .A(DP_OP_425J2_127_3477_n190), .B(
        DP_OP_425J2_127_3477_n199), .CI(DP_OP_425J2_127_3477_n197), .CO(
        DP_OP_425J2_127_3477_n187), .S(DP_OP_425J2_127_3477_n188) );
  FADDX1_HVT DP_OP_425J2_127_3477_U189 ( .A(DP_OP_425J2_127_3477_n188), .B(
        DP_OP_425J2_127_3477_n195), .CI(DP_OP_425J2_127_3477_n193), .CO(
        DP_OP_425J2_127_3477_n185), .S(DP_OP_425J2_127_3477_n186) );
  FADDX1_HVT DP_OP_425J2_127_3477_U188 ( .A(DP_OP_425J2_127_3477_n1774), .B(
        DP_OP_425J2_127_3477_n189), .CI(DP_OP_425J2_127_3477_n187), .CO(
        DP_OP_425J2_127_3477_n183), .S(DP_OP_425J2_127_3477_n184) );
  FADDX1_HVT DP_OP_425J2_127_3477_U171 ( .A(DP_OP_425J2_127_3477_n1754), .B(
        DP_OP_425J2_127_3477_n1752), .CI(DP_OP_425J2_127_3477_n1750), .CO(
        DP_OP_425J2_127_3477_n131), .S(n_conv2_sum_d[0]) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U170 ( .A1(DP_OP_425J2_127_3477_n1688), 
        .A2(DP_OP_425J2_127_3477_n1690), .Y(DP_OP_425J2_127_3477_n130) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U169 ( .A1(DP_OP_425J2_127_3477_n1690), .A2(
        DP_OP_425J2_127_3477_n1688), .Y(DP_OP_425J2_127_3477_n129) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U163 ( .A1(DP_OP_425J2_127_3477_n1582), 
        .A2(DP_OP_425J2_127_3477_n1584), .Y(DP_OP_425J2_127_3477_n127) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U155 ( .A1(DP_OP_425J2_127_3477_n1428), 
        .A2(DP_OP_425J2_127_3477_n1430), .Y(DP_OP_425J2_127_3477_n122) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U154 ( .A1(DP_OP_425J2_127_3477_n1430), .A2(
        DP_OP_425J2_127_3477_n1428), .Y(DP_OP_425J2_127_3477_n121) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U149 ( .A1(DP_OP_425J2_127_3477_n1252), 
        .A2(DP_OP_425J2_127_3477_n1254), .Y(DP_OP_425J2_127_3477_n119) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U141 ( .A1(DP_OP_425J2_127_3477_n1064), 
        .A2(DP_OP_425J2_127_3477_n1066), .Y(DP_OP_425J2_127_3477_n114) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U140 ( .A1(DP_OP_425J2_127_3477_n1066), .A2(
        DP_OP_425J2_127_3477_n1064), .Y(DP_OP_425J2_127_3477_n113) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U135 ( .A1(DP_OP_425J2_127_3477_n870), .A2(
        DP_OP_425J2_127_3477_n872), .Y(DP_OP_425J2_127_3477_n111) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U127 ( .A1(DP_OP_425J2_127_3477_n674), .A2(
        DP_OP_425J2_127_3477_n869), .Y(DP_OP_425J2_127_3477_n106) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U126 ( .A1(DP_OP_425J2_127_3477_n869), .A2(
        DP_OP_425J2_127_3477_n674), .Y(DP_OP_425J2_127_3477_n105) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U120 ( .A1(DP_OP_425J2_127_3477_n500), .A2(
        DP_OP_425J2_127_3477_n673), .Y(DP_OP_425J2_127_3477_n102) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U119 ( .A1(DP_OP_425J2_127_3477_n673), .A2(
        DP_OP_425J2_127_3477_n500), .Y(DP_OP_425J2_127_3477_n101) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U114 ( .A1(DP_OP_425J2_127_3477_n364), .A2(
        DP_OP_425J2_127_3477_n499), .Y(DP_OP_425J2_127_3477_n99) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U113 ( .A1(DP_OP_425J2_127_3477_n499), .A2(
        DP_OP_425J2_127_3477_n364), .Y(DP_OP_425J2_127_3477_n98) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U105 ( .A1(DP_OP_425J2_127_3477_n270), .A2(
        DP_OP_425J2_127_3477_n363), .Y(DP_OP_425J2_127_3477_n93) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U104 ( .A1(DP_OP_425J2_127_3477_n363), .A2(
        DP_OP_425J2_127_3477_n270), .Y(DP_OP_425J2_127_3477_n92) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U97 ( .A1(DP_OP_425J2_127_3477_n224), .A2(
        DP_OP_425J2_127_3477_n269), .Y(DP_OP_425J2_127_3477_n88) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U96 ( .A1(DP_OP_425J2_127_3477_n269), .A2(
        DP_OP_425J2_127_3477_n224), .Y(DP_OP_425J2_127_3477_n87) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U92 ( .A1(DP_OP_425J2_127_3477_n87), .A2(
        DP_OP_425J2_127_3477_n92), .Y(DP_OP_425J2_127_3477_n85) );
  AOI21X1_HVT DP_OP_425J2_127_3477_U91 ( .A1(DP_OP_425J2_127_3477_n94), .A2(
        DP_OP_425J2_127_3477_n85), .A3(DP_OP_425J2_127_3477_n86), .Y(
        DP_OP_425J2_127_3477_n84) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U89 ( .A1(DP_OP_425J2_127_3477_n202), .A2(
        DP_OP_425J2_127_3477_n223), .Y(DP_OP_425J2_127_3477_n83) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U88 ( .A1(DP_OP_425J2_127_3477_n223), .A2(
        DP_OP_425J2_127_3477_n202), .Y(DP_OP_425J2_127_3477_n82) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U83 ( .A1(DP_OP_425J2_127_3477_n201), .A2(
        DP_OP_425J2_127_3477_n192), .Y(DP_OP_425J2_127_3477_n80) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U82 ( .A1(DP_OP_425J2_127_3477_n192), .A2(
        DP_OP_425J2_127_3477_n201), .Y(DP_OP_425J2_127_3477_n79) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U78 ( .A1(DP_OP_425J2_127_3477_n79), .A2(
        DP_OP_425J2_127_3477_n82), .Y(DP_OP_425J2_127_3477_n77) );
  AOI21X1_HVT DP_OP_425J2_127_3477_U77 ( .A1(DP_OP_425J2_127_3477_n86), .A2(
        DP_OP_425J2_127_3477_n77), .A3(DP_OP_425J2_127_3477_n78), .Y(
        DP_OP_425J2_127_3477_n76) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U76 ( .A1(DP_OP_425J2_127_3477_n85), .A2(
        DP_OP_425J2_127_3477_n77), .Y(DP_OP_425J2_127_3477_n75) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U72 ( .A1(DP_OP_425J2_127_3477_n191), .A2(
        DP_OP_425J2_127_3477_n186), .Y(DP_OP_425J2_127_3477_n68) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U71 ( .A1(DP_OP_425J2_127_3477_n186), .A2(
        DP_OP_425J2_127_3477_n191), .Y(DP_OP_425J2_127_3477_n67) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U62 ( .A1(DP_OP_425J2_127_3477_n185), .A2(
        DP_OP_425J2_127_3477_n184), .Y(DP_OP_425J2_127_3477_n65) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U61 ( .A1(DP_OP_425J2_127_3477_n184), .A2(
        DP_OP_425J2_127_3477_n185), .Y(DP_OP_425J2_127_3477_n64) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U54 ( .A1(DP_OP_425J2_127_3477_n183), .A2(
        DP_OP_425J2_127_3477_n182), .Y(DP_OP_425J2_127_3477_n60) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U53 ( .A1(DP_OP_425J2_127_3477_n182), .A2(
        DP_OP_425J2_127_3477_n183), .Y(DP_OP_425J2_127_3477_n59) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U49 ( .A1(DP_OP_425J2_127_3477_n59), .A2(
        DP_OP_425J2_127_3477_n64), .Y(DP_OP_425J2_127_3477_n57) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U47 ( .A1(DP_OP_425J2_127_3477_n69), .A2(
        DP_OP_425J2_127_3477_n57), .Y(DP_OP_425J2_127_3477_n55) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U44 ( .A1(DP_OP_425J2_127_3477_n180), .A2(
        DP_OP_425J2_127_3477_n181), .Y(DP_OP_425J2_127_3477_n53) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U43 ( .A1(DP_OP_425J2_127_3477_n181), .A2(
        DP_OP_425J2_127_3477_n180), .Y(DP_OP_425J2_127_3477_n52) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U39 ( .A1(DP_OP_425J2_127_3477_n52), .A2(
        DP_OP_425J2_127_3477_n55), .Y(DP_OP_425J2_127_3477_n50) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U34 ( .A1(DP_OP_425J2_127_3477_n178), .A2(
        DP_OP_425J2_127_3477_n179), .Y(DP_OP_425J2_127_3477_n46) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U27 ( .A1(DP_OP_425J2_127_3477_n50), .A2(
        DP_OP_425J2_127_3477_n45), .Y(DP_OP_425J2_127_3477_n41) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U24 ( .A1(DP_OP_425J2_127_3477_n176), .A2(
        DP_OP_425J2_127_3477_n177), .Y(DP_OP_425J2_127_3477_n39) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U23 ( .A1(DP_OP_425J2_127_3477_n177), .A2(
        DP_OP_425J2_127_3477_n176), .Y(DP_OP_425J2_127_3477_n38) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U19 ( .A1(DP_OP_425J2_127_3477_n38), .A2(
        DP_OP_425J2_127_3477_n41), .Y(DP_OP_425J2_127_3477_n36) );
  FADDX1_HVT DP_OP_425J2_127_3477_U15 ( .A(DP_OP_425J2_127_3477_n175), .B(
        DP_OP_425J2_127_3477_n174), .CI(DP_OP_425J2_127_3477_n35), .CO(
        DP_OP_425J2_127_3477_n34), .S(n_conv2_sum_d[20]) );
  FADDX1_HVT DP_OP_425J2_127_3477_U14 ( .A(DP_OP_425J2_127_3477_n173), .B(
        DP_OP_425J2_127_3477_n172), .CI(DP_OP_425J2_127_3477_n34), .CO(
        DP_OP_425J2_127_3477_n33), .S(n_conv2_sum_d[21]) );
  FADDX1_HVT DP_OP_425J2_127_3477_U13 ( .A(DP_OP_425J2_127_3477_n171), .B(
        DP_OP_425J2_127_3477_n170), .CI(DP_OP_425J2_127_3477_n33), .CO(
        DP_OP_425J2_127_3477_n32), .S(n_conv2_sum_d[22]) );
  FADDX1_HVT DP_OP_425J2_127_3477_U12 ( .A(DP_OP_425J2_127_3477_n169), .B(
        DP_OP_425J2_127_3477_n168), .CI(DP_OP_425J2_127_3477_n32), .CO(
        DP_OP_425J2_127_3477_n31), .S(n_conv2_sum_d[23]) );
  FADDX1_HVT DP_OP_425J2_127_3477_U11 ( .A(DP_OP_425J2_127_3477_n167), .B(
        DP_OP_425J2_127_3477_n166), .CI(DP_OP_425J2_127_3477_n31), .CO(
        DP_OP_425J2_127_3477_n30), .S(n_conv2_sum_d[24]) );
  FADDX1_HVT DP_OP_425J2_127_3477_U10 ( .A(DP_OP_425J2_127_3477_n165), .B(
        DP_OP_425J2_127_3477_n164), .CI(DP_OP_425J2_127_3477_n30), .CO(
        DP_OP_425J2_127_3477_n29), .S(n_conv2_sum_d[25]) );
  FADDX1_HVT DP_OP_425J2_127_3477_U9 ( .A(DP_OP_425J2_127_3477_n163), .B(
        DP_OP_425J2_127_3477_n162), .CI(DP_OP_425J2_127_3477_n29), .CO(
        DP_OP_425J2_127_3477_n28), .S(n_conv2_sum_d[26]) );
  FADDX1_HVT DP_OP_425J2_127_3477_U8 ( .A(DP_OP_425J2_127_3477_n161), .B(
        DP_OP_425J2_127_3477_n160), .CI(DP_OP_425J2_127_3477_n28), .CO(
        DP_OP_425J2_127_3477_n27), .S(n_conv2_sum_d[27]) );
  FADDX1_HVT DP_OP_425J2_127_3477_U7 ( .A(DP_OP_425J2_127_3477_n159), .B(
        DP_OP_425J2_127_3477_n158), .CI(DP_OP_425J2_127_3477_n27), .CO(
        DP_OP_425J2_127_3477_n26), .S(n_conv2_sum_d[28]) );
  FADDX1_HVT DP_OP_425J2_127_3477_U6 ( .A(DP_OP_425J2_127_3477_n157), .B(
        DP_OP_425J2_127_3477_n156), .CI(DP_OP_425J2_127_3477_n26), .CO(
        DP_OP_425J2_127_3477_n25), .S(n_conv2_sum_d[29]) );
  FADDX1_HVT DP_OP_425J2_127_3477_U5 ( .A(DP_OP_425J2_127_3477_n155), .B(
        DP_OP_425J2_127_3477_n154), .CI(DP_OP_425J2_127_3477_n25), .CO(
        DP_OP_425J2_127_3477_n24), .S(n_conv2_sum_d[30]) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2129 ( .A1(DP_OP_425J2_127_3477_n1854), .A2(
        DP_OP_423J2_125_3477_n2913), .Y(DP_OP_424J2_126_3477_n2899) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2122 ( .A1(DP_OP_425J2_127_3477_n1855), 
        .A2(DP_OP_424J2_126_3477_n2917), .Y(DP_OP_424J2_126_3477_n2892) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2121 ( .A1(DP_OP_425J2_127_3477_n1854), .A2(
        DP_OP_424J2_126_3477_n2917), .Y(DP_OP_424J2_126_3477_n2891) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2114 ( .A1(DP_OP_425J2_127_3477_n1855), 
        .A2(DP_OP_425J2_127_3477_n2916), .Y(DP_OP_424J2_126_3477_n2884) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2113 ( .A1(DP_OP_425J2_127_3477_n1854), .A2(
        DP_OP_425J2_127_3477_n2916), .Y(DP_OP_424J2_126_3477_n2883) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2112 ( .A1(DP_OP_425J2_127_3477_n1861), .A2(
        DP_OP_424J2_126_3477_n2915), .Y(DP_OP_424J2_126_3477_n2882) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2111 ( .A1(DP_OP_425J2_127_3477_n1860), .A2(
        DP_OP_424J2_126_3477_n2915), .Y(DP_OP_424J2_126_3477_n2881) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2110 ( .A1(DP_OP_424J2_126_3477_n2912), .A2(
        DP_OP_424J2_126_3477_n2915), .Y(DP_OP_424J2_126_3477_n2880) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2109 ( .A1(DP_OP_425J2_127_3477_n1858), .A2(
        DP_OP_424J2_126_3477_n2915), .Y(DP_OP_424J2_126_3477_n2879) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2108 ( .A1(DP_OP_424J2_126_3477_n2910), .A2(
        DP_OP_424J2_126_3477_n2915), .Y(DP_OP_424J2_126_3477_n2878) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2107 ( .A1(DP_OP_424J2_126_3477_n2909), .A2(
        DP_OP_424J2_126_3477_n2915), .Y(DP_OP_424J2_126_3477_n2877) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2106 ( .A1(DP_OP_425J2_127_3477_n1855), .A2(
        DP_OP_424J2_126_3477_n2915), .Y(DP_OP_424J2_126_3477_n2876) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2105 ( .A1(DP_OP_425J2_127_3477_n1854), 
        .A2(DP_OP_424J2_126_3477_n2915), .Y(DP_OP_424J2_126_3477_n2875) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2086 ( .A1(DP_OP_424J2_126_3477_n2864), 
        .A2(DP_OP_424J2_126_3477_n2874), .Y(DP_OP_424J2_126_3477_n2856) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2085 ( .A1(DP_OP_424J2_126_3477_n2863), .A2(
        DP_OP_424J2_126_3477_n2874), .Y(DP_OP_424J2_126_3477_n2855) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2078 ( .A1(DP_OP_424J2_126_3477_n2864), 
        .A2(DP_OP_424J2_126_3477_n2873), .Y(DP_OP_424J2_126_3477_n2848) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2077 ( .A1(DP_OP_424J2_126_3477_n2863), .A2(
        DP_OP_424J2_126_3477_n2873), .Y(DP_OP_424J2_126_3477_n2847) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2070 ( .A1(DP_OP_424J2_126_3477_n2864), 
        .A2(DP_OP_425J2_127_3477_n2872), .Y(DP_OP_424J2_126_3477_n2840) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2069 ( .A1(DP_OP_424J2_126_3477_n2863), .A2(
        DP_OP_422J2_124_3477_n2872), .Y(DP_OP_424J2_126_3477_n2839) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2068 ( .A1(DP_OP_425J2_127_3477_n1905), .A2(
        DP_OP_423J2_125_3477_n2866), .Y(DP_OP_424J2_126_3477_n2838) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2067 ( .A1(DP_OP_424J2_126_3477_n2869), .A2(
        DP_OP_423J2_125_3477_n2866), .Y(DP_OP_424J2_126_3477_n2837) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2066 ( .A1(DP_OP_425J2_127_3477_n1903), .A2(
        DP_OP_425J2_127_3477_n2871), .Y(DP_OP_424J2_126_3477_n2836) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2065 ( .A1(DP_OP_424J2_126_3477_n2867), .A2(
        DP_OP_423J2_125_3477_n2866), .Y(DP_OP_424J2_126_3477_n2835) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2064 ( .A1(DP_OP_425J2_127_3477_n1901), .A2(
        DP_OP_423J2_125_3477_n2866), .Y(DP_OP_424J2_126_3477_n2834) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2063 ( .A1(DP_OP_424J2_126_3477_n2865), .A2(
        DP_OP_423J2_125_3477_n2866), .Y(DP_OP_424J2_126_3477_n2833) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2062 ( .A1(DP_OP_424J2_126_3477_n2864), .A2(
        DP_OP_422J2_124_3477_n2871), .Y(DP_OP_424J2_126_3477_n2832) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2061 ( .A1(DP_OP_424J2_126_3477_n2863), 
        .A2(DP_OP_425J2_127_3477_n2871), .Y(DP_OP_424J2_126_3477_n2831) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2042 ( .A1(DP_OP_424J2_126_3477_n2820), 
        .A2(DP_OP_424J2_126_3477_n2830), .Y(DP_OP_424J2_126_3477_n2812) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2041 ( .A1(DP_OP_424J2_126_3477_n2819), .A2(
        DP_OP_424J2_126_3477_n2830), .Y(DP_OP_424J2_126_3477_n2811) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2034 ( .A1(DP_OP_424J2_126_3477_n2820), 
        .A2(DP_OP_424J2_126_3477_n2829), .Y(DP_OP_424J2_126_3477_n2804) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2033 ( .A1(DP_OP_424J2_126_3477_n2819), .A2(
        DP_OP_424J2_126_3477_n2829), .Y(DP_OP_424J2_126_3477_n2803) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2025 ( .A1(DP_OP_424J2_126_3477_n2819), .A2(
        DP_OP_424J2_126_3477_n2828), .Y(DP_OP_424J2_126_3477_n2795) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2024 ( .A1(DP_OP_424J2_126_3477_n2826), .A2(
        DP_OP_424J2_126_3477_n2827), .Y(DP_OP_424J2_126_3477_n2794) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2023 ( .A1(DP_OP_424J2_126_3477_n2825), .A2(
        DP_OP_424J2_126_3477_n2827), .Y(DP_OP_424J2_126_3477_n2793) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2022 ( .A1(DP_OP_424J2_126_3477_n2824), .A2(
        DP_OP_424J2_126_3477_n2827), .Y(DP_OP_424J2_126_3477_n2792) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2021 ( .A1(DP_OP_424J2_126_3477_n2823), .A2(
        DP_OP_424J2_126_3477_n2827), .Y(DP_OP_424J2_126_3477_n2791) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2020 ( .A1(DP_OP_424J2_126_3477_n2822), .A2(
        DP_OP_424J2_126_3477_n2827), .Y(DP_OP_424J2_126_3477_n2790) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2019 ( .A1(DP_OP_424J2_126_3477_n2821), .A2(
        DP_OP_424J2_126_3477_n2827), .Y(DP_OP_424J2_126_3477_n2789) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2018 ( .A1(DP_OP_424J2_126_3477_n2820), .A2(
        DP_OP_424J2_126_3477_n2827), .Y(DP_OP_424J2_126_3477_n2788) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2017 ( .A1(DP_OP_424J2_126_3477_n2819), 
        .A2(DP_OP_424J2_126_3477_n2827), .Y(DP_OP_424J2_126_3477_n2787) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1998 ( .A1(DP_OP_423J2_125_3477_n2859), 
        .A2(DP_OP_422J2_124_3477_n2786), .Y(DP_OP_424J2_126_3477_n2768) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1997 ( .A1(DP_OP_424J2_126_3477_n2775), .A2(
        DP_OP_423J2_125_3477_n2781), .Y(DP_OP_424J2_126_3477_n2767) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1990 ( .A1(DP_OP_423J2_125_3477_n2859), 
        .A2(DP_OP_424J2_126_3477_n2785), .Y(DP_OP_424J2_126_3477_n2760) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1989 ( .A1(DP_OP_424J2_126_3477_n2775), .A2(
        DP_OP_424J2_126_3477_n2785), .Y(DP_OP_424J2_126_3477_n2759) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1982 ( .A1(DP_OP_423J2_125_3477_n2859), 
        .A2(DP_OP_424J2_126_3477_n2784), .Y(DP_OP_424J2_126_3477_n2752) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1981 ( .A1(DP_OP_424J2_126_3477_n2775), .A2(
        DP_OP_424J2_126_3477_n2784), .Y(DP_OP_424J2_126_3477_n2751) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1980 ( .A1(DP_OP_423J2_125_3477_n2865), .A2(
        DP_OP_424J2_126_3477_n2783), .Y(DP_OP_424J2_126_3477_n2750) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1979 ( .A1(DP_OP_423J2_125_3477_n2864), .A2(
        DP_OP_424J2_126_3477_n2783), .Y(DP_OP_424J2_126_3477_n2749) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1978 ( .A1(DP_OP_425J2_127_3477_n1991), .A2(
        DP_OP_424J2_126_3477_n2783), .Y(DP_OP_424J2_126_3477_n2748) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1977 ( .A1(DP_OP_422J2_124_3477_n1858), .A2(
        DP_OP_424J2_126_3477_n2783), .Y(DP_OP_424J2_126_3477_n2747) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1976 ( .A1(DP_OP_425J2_127_3477_n1989), .A2(
        DP_OP_424J2_126_3477_n2783), .Y(DP_OP_424J2_126_3477_n2746) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1975 ( .A1(DP_OP_424J2_126_3477_n2777), .A2(
        DP_OP_424J2_126_3477_n2783), .Y(DP_OP_424J2_126_3477_n2745) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1974 ( .A1(DP_OP_423J2_125_3477_n2859), .A2(
        DP_OP_424J2_126_3477_n2783), .Y(DP_OP_424J2_126_3477_n2744) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1973 ( .A1(DP_OP_424J2_126_3477_n2775), 
        .A2(DP_OP_424J2_126_3477_n2783), .Y(DP_OP_424J2_126_3477_n2743) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1954 ( .A1(DP_OP_424J2_126_3477_n2732), 
        .A2(DP_OP_424J2_126_3477_n2742), .Y(DP_OP_424J2_126_3477_n2724) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1953 ( .A1(DP_OP_424J2_126_3477_n2731), .A2(
        DP_OP_424J2_126_3477_n2742), .Y(DP_OP_424J2_126_3477_n2723) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1945 ( .A1(DP_OP_424J2_126_3477_n2731), .A2(
        DP_OP_424J2_126_3477_n2741), .Y(DP_OP_424J2_126_3477_n2715) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1938 ( .A1(DP_OP_424J2_126_3477_n2732), 
        .A2(DP_OP_424J2_126_3477_n2740), .Y(DP_OP_424J2_126_3477_n2708) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1937 ( .A1(DP_OP_424J2_126_3477_n2731), .A2(
        DP_OP_424J2_126_3477_n2740), .Y(DP_OP_424J2_126_3477_n2707) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1936 ( .A1(DP_OP_424J2_126_3477_n2738), .A2(
        DP_OP_423J2_125_3477_n2734), .Y(DP_OP_424J2_126_3477_n2706) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1935 ( .A1(DP_OP_424J2_126_3477_n2737), .A2(
        DP_OP_425J2_127_3477_n2739), .Y(DP_OP_424J2_126_3477_n2705) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1934 ( .A1(DP_OP_424J2_126_3477_n2736), .A2(
        DP_OP_423J2_125_3477_n2734), .Y(DP_OP_424J2_126_3477_n2704) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1933 ( .A1(DP_OP_424J2_126_3477_n2735), .A2(
        DP_OP_425J2_127_3477_n2739), .Y(DP_OP_424J2_126_3477_n2703) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1932 ( .A1(DP_OP_424J2_126_3477_n2734), .A2(
        DP_OP_423J2_125_3477_n2734), .Y(DP_OP_424J2_126_3477_n2702) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1931 ( .A1(DP_OP_424J2_126_3477_n2733), .A2(
        DP_OP_423J2_125_3477_n2734), .Y(DP_OP_424J2_126_3477_n2701) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1930 ( .A1(DP_OP_424J2_126_3477_n2732), .A2(
        DP_OP_425J2_127_3477_n2739), .Y(DP_OP_424J2_126_3477_n2700) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1929 ( .A1(DP_OP_424J2_126_3477_n2731), 
        .A2(DP_OP_423J2_125_3477_n2734), .Y(DP_OP_424J2_126_3477_n2699) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1910 ( .A1(DP_OP_422J2_124_3477_n1943), 
        .A2(DP_OP_424J2_126_3477_n2698), .Y(DP_OP_424J2_126_3477_n2680) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1909 ( .A1(DP_OP_423J2_125_3477_n2770), .A2(
        DP_OP_424J2_126_3477_n2698), .Y(DP_OP_424J2_126_3477_n2679) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1902 ( .A1(DP_OP_422J2_124_3477_n1943), 
        .A2(DP_OP_424J2_126_3477_n2697), .Y(DP_OP_424J2_126_3477_n2672) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1901 ( .A1(DP_OP_425J2_127_3477_n2074), .A2(
        DP_OP_424J2_126_3477_n2697), .Y(DP_OP_424J2_126_3477_n2671) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1893 ( .A1(DP_OP_423J2_125_3477_n2770), .A2(
        DP_OP_424J2_126_3477_n2696), .Y(DP_OP_424J2_126_3477_n2663) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1892 ( .A1(DP_OP_423J2_125_3477_n2777), .A2(
        DP_OP_424J2_126_3477_n2695), .Y(DP_OP_424J2_126_3477_n2662) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1891 ( .A1(DP_OP_424J2_126_3477_n2693), .A2(
        DP_OP_424J2_126_3477_n2695), .Y(DP_OP_424J2_126_3477_n2661) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1890 ( .A1(DP_OP_423J2_125_3477_n2775), .A2(
        DP_OP_424J2_126_3477_n2695), .Y(DP_OP_424J2_126_3477_n2660) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1889 ( .A1(DP_OP_424J2_126_3477_n2691), .A2(
        DP_OP_424J2_126_3477_n2695), .Y(DP_OP_424J2_126_3477_n2659) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1888 ( .A1(DP_OP_422J2_124_3477_n1945), .A2(
        DP_OP_424J2_126_3477_n2695), .Y(DP_OP_424J2_126_3477_n2658) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1887 ( .A1(DP_OP_424J2_126_3477_n2689), .A2(
        DP_OP_424J2_126_3477_n2695), .Y(DP_OP_424J2_126_3477_n2657) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1886 ( .A1(DP_OP_422J2_124_3477_n1943), .A2(
        DP_OP_424J2_126_3477_n2695), .Y(DP_OP_424J2_126_3477_n2656) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1885 ( .A1(DP_OP_425J2_127_3477_n2074), 
        .A2(DP_OP_424J2_126_3477_n2695), .Y(DP_OP_424J2_126_3477_n2655) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1866 ( .A1(DP_OP_424J2_126_3477_n2644), 
        .A2(DP_OP_424J2_126_3477_n2654), .Y(DP_OP_424J2_126_3477_n2636) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1865 ( .A1(DP_OP_425J2_127_3477_n2118), .A2(
        DP_OP_424J2_126_3477_n2654), .Y(DP_OP_424J2_126_3477_n2635) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1858 ( .A1(DP_OP_424J2_126_3477_n2644), 
        .A2(DP_OP_424J2_126_3477_n2653), .Y(DP_OP_424J2_126_3477_n2628) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1857 ( .A1(DP_OP_423J2_125_3477_n2726), .A2(
        DP_OP_424J2_126_3477_n2653), .Y(DP_OP_424J2_126_3477_n2627) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1850 ( .A1(DP_OP_424J2_126_3477_n2644), 
        .A2(DP_OP_424J2_126_3477_n2652), .Y(DP_OP_424J2_126_3477_n2620) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1849 ( .A1(DP_OP_425J2_127_3477_n2118), .A2(
        DP_OP_424J2_126_3477_n2652), .Y(DP_OP_424J2_126_3477_n2619) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1848 ( .A1(DP_OP_424J2_126_3477_n2650), .A2(
        DP_OP_424J2_126_3477_n2651), .Y(DP_OP_424J2_126_3477_n2618) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1847 ( .A1(DP_OP_424J2_126_3477_n2649), .A2(
        DP_OP_424J2_126_3477_n2651), .Y(DP_OP_424J2_126_3477_n2617) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1846 ( .A1(DP_OP_422J2_124_3477_n1991), .A2(
        DP_OP_424J2_126_3477_n2651), .Y(DP_OP_424J2_126_3477_n2616) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1845 ( .A1(DP_OP_425J2_127_3477_n2122), .A2(
        DP_OP_424J2_126_3477_n2651), .Y(DP_OP_424J2_126_3477_n2615) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1844 ( .A1(DP_OP_422J2_124_3477_n1989), .A2(
        DP_OP_424J2_126_3477_n2651), .Y(DP_OP_424J2_126_3477_n2614) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1843 ( .A1(DP_OP_422J2_124_3477_n1988), .A2(
        DP_OP_424J2_126_3477_n2651), .Y(DP_OP_424J2_126_3477_n2613) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1842 ( .A1(DP_OP_424J2_126_3477_n2644), .A2(
        DP_OP_424J2_126_3477_n2651), .Y(DP_OP_424J2_126_3477_n2612) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1841 ( .A1(DP_OP_423J2_125_3477_n2726), 
        .A2(DP_OP_424J2_126_3477_n2651), .Y(DP_OP_424J2_126_3477_n2611) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1822 ( .A1(DP_OP_424J2_126_3477_n2600), 
        .A2(DP_OP_424J2_126_3477_n2610), .Y(DP_OP_424J2_126_3477_n2592) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1821 ( .A1(DP_OP_422J2_124_3477_n2029), .A2(
        DP_OP_424J2_126_3477_n2610), .Y(DP_OP_424J2_126_3477_n2591) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1814 ( .A1(DP_OP_424J2_126_3477_n2600), 
        .A2(DP_OP_424J2_126_3477_n2609), .Y(DP_OP_424J2_126_3477_n2584) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1813 ( .A1(DP_OP_422J2_124_3477_n2029), .A2(
        DP_OP_424J2_126_3477_n2609), .Y(DP_OP_424J2_126_3477_n2583) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1806 ( .A1(DP_OP_424J2_126_3477_n2600), 
        .A2(DP_OP_424J2_126_3477_n2608), .Y(DP_OP_424J2_126_3477_n2576) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1805 ( .A1(DP_OP_422J2_124_3477_n2029), .A2(
        DP_OP_424J2_126_3477_n2608), .Y(DP_OP_424J2_126_3477_n2575) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1804 ( .A1(DP_OP_422J2_124_3477_n2036), .A2(
        DP_OP_424J2_126_3477_n2607), .Y(DP_OP_424J2_126_3477_n2574) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1803 ( .A1(DP_OP_422J2_124_3477_n2035), .A2(
        DP_OP_424J2_126_3477_n2607), .Y(DP_OP_424J2_126_3477_n2573) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1802 ( .A1(DP_OP_424J2_126_3477_n2604), .A2(
        DP_OP_424J2_126_3477_n2607), .Y(DP_OP_424J2_126_3477_n2572) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1801 ( .A1(DP_OP_422J2_124_3477_n2033), .A2(
        DP_OP_424J2_126_3477_n2607), .Y(DP_OP_424J2_126_3477_n2571) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1800 ( .A1(DP_OP_422J2_124_3477_n2032), .A2(
        DP_OP_424J2_126_3477_n2607), .Y(DP_OP_424J2_126_3477_n2570) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1799 ( .A1(DP_OP_422J2_124_3477_n2031), .A2(
        DP_OP_424J2_126_3477_n2607), .Y(DP_OP_424J2_126_3477_n2569) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1798 ( .A1(DP_OP_424J2_126_3477_n2600), .A2(
        DP_OP_424J2_126_3477_n2607), .Y(DP_OP_424J2_126_3477_n2568) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1797 ( .A1(DP_OP_422J2_124_3477_n2029), 
        .A2(DP_OP_424J2_126_3477_n2607), .Y(DP_OP_424J2_126_3477_n2567) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1778 ( .A1(DP_OP_423J2_125_3477_n2642), 
        .A2(DP_OP_424J2_126_3477_n2566), .Y(DP_OP_424J2_126_3477_n2548) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1777 ( .A1(DP_OP_424J2_126_3477_n2555), .A2(
        DP_OP_424J2_126_3477_n2566), .Y(DP_OP_424J2_126_3477_n2547) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1769 ( .A1(DP_OP_424J2_126_3477_n2555), .A2(
        DP_OP_424J2_126_3477_n2565), .Y(DP_OP_424J2_126_3477_n2539) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1762 ( .A1(DP_OP_422J2_124_3477_n2074), 
        .A2(DP_OP_422J2_124_3477_n2566), .Y(DP_OP_424J2_126_3477_n2532) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1761 ( .A1(DP_OP_424J2_126_3477_n2555), .A2(
        DP_OP_425J2_127_3477_n2564), .Y(DP_OP_424J2_126_3477_n2531) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1760 ( .A1(DP_OP_423J2_125_3477_n2648), .A2(
        DP_OP_424J2_126_3477_n2563), .Y(DP_OP_424J2_126_3477_n2530) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1759 ( .A1(DP_OP_424J2_126_3477_n2561), .A2(
        DP_OP_424J2_126_3477_n2563), .Y(DP_OP_424J2_126_3477_n2529) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1758 ( .A1(DP_OP_422J2_124_3477_n2078), .A2(
        DP_OP_424J2_126_3477_n2563), .Y(DP_OP_424J2_126_3477_n2528) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1757 ( .A1(DP_OP_424J2_126_3477_n2559), .A2(
        DP_OP_424J2_126_3477_n2563), .Y(DP_OP_424J2_126_3477_n2527) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1756 ( .A1(DP_OP_422J2_124_3477_n2076), .A2(
        DP_OP_424J2_126_3477_n2563), .Y(DP_OP_424J2_126_3477_n2526) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1755 ( .A1(DP_OP_424J2_126_3477_n2557), .A2(
        DP_OP_424J2_126_3477_n2563), .Y(DP_OP_424J2_126_3477_n2525) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1754 ( .A1(DP_OP_422J2_124_3477_n2074), .A2(
        DP_OP_424J2_126_3477_n2563), .Y(DP_OP_424J2_126_3477_n2524) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1753 ( .A1(DP_OP_424J2_126_3477_n2555), 
        .A2(DP_OP_424J2_126_3477_n2563), .Y(DP_OP_424J2_126_3477_n2523) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1734 ( .A1(DP_OP_424J2_126_3477_n2512), 
        .A2(DP_OP_424J2_126_3477_n2522), .Y(DP_OP_424J2_126_3477_n2504) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1733 ( .A1(DP_OP_425J2_127_3477_n2250), .A2(
        DP_OP_424J2_126_3477_n2522), .Y(DP_OP_424J2_126_3477_n2503) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1725 ( .A1(DP_OP_425J2_127_3477_n2250), .A2(
        DP_OP_424J2_126_3477_n2521), .Y(DP_OP_424J2_126_3477_n2495) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1718 ( .A1(DP_OP_424J2_126_3477_n2512), 
        .A2(DP_OP_424J2_126_3477_n2520), .Y(DP_OP_424J2_126_3477_n2488) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1717 ( .A1(DP_OP_425J2_127_3477_n2250), .A2(
        DP_OP_424J2_126_3477_n2520), .Y(DP_OP_424J2_126_3477_n2487) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1716 ( .A1(DP_OP_423J2_125_3477_n2604), .A2(
        DP_OP_425J2_127_3477_n2519), .Y(DP_OP_424J2_126_3477_n2486) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1715 ( .A1(DP_OP_424J2_126_3477_n2517), .A2(
        DP_OP_425J2_127_3477_n2519), .Y(DP_OP_424J2_126_3477_n2485) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1714 ( .A1(DP_OP_425J2_127_3477_n2255), .A2(
        DP_OP_425J2_127_3477_n2519), .Y(DP_OP_424J2_126_3477_n2484) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1713 ( .A1(DP_OP_422J2_124_3477_n2121), .A2(
        DP_OP_423J2_125_3477_n2517), .Y(DP_OP_424J2_126_3477_n2483) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1712 ( .A1(DP_OP_423J2_125_3477_n2600), .A2(
        DP_OP_423J2_125_3477_n2517), .Y(DP_OP_424J2_126_3477_n2482) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1711 ( .A1(DP_OP_425J2_127_3477_n2252), .A2(
        DP_OP_425J2_127_3477_n2519), .Y(DP_OP_424J2_126_3477_n2481) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1710 ( .A1(DP_OP_424J2_126_3477_n2512), .A2(
        DP_OP_423J2_125_3477_n2517), .Y(DP_OP_424J2_126_3477_n2480) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1709 ( .A1(DP_OP_422J2_124_3477_n2117), 
        .A2(DP_OP_425J2_127_3477_n2519), .Y(DP_OP_424J2_126_3477_n2479) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1690 ( .A1(DP_OP_423J2_125_3477_n2554), 
        .A2(DP_OP_424J2_126_3477_n2478), .Y(DP_OP_424J2_126_3477_n2460) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1689 ( .A1(DP_OP_425J2_127_3477_n2294), .A2(
        DP_OP_424J2_126_3477_n2478), .Y(DP_OP_424J2_126_3477_n2459) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1682 ( .A1(DP_OP_423J2_125_3477_n2554), 
        .A2(DP_OP_423J2_125_3477_n2475), .Y(DP_OP_424J2_126_3477_n2452) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1681 ( .A1(DP_OP_423J2_125_3477_n2553), .A2(
        DP_OP_423J2_125_3477_n2475), .Y(DP_OP_424J2_126_3477_n2451) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1674 ( .A1(DP_OP_423J2_125_3477_n2554), 
        .A2(DP_OP_422J2_124_3477_n2478), .Y(DP_OP_424J2_126_3477_n2444) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1673 ( .A1(DP_OP_425J2_127_3477_n2294), .A2(
        DP_OP_425J2_127_3477_n2476), .Y(DP_OP_424J2_126_3477_n2443) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1672 ( .A1(DP_OP_424J2_126_3477_n2474), .A2(
        DP_OP_424J2_126_3477_n2475), .Y(DP_OP_424J2_126_3477_n2442) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1671 ( .A1(DP_OP_423J2_125_3477_n2559), .A2(
        DP_OP_424J2_126_3477_n2475), .Y(DP_OP_424J2_126_3477_n2441) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1670 ( .A1(DP_OP_424J2_126_3477_n2472), .A2(
        DP_OP_424J2_126_3477_n2475), .Y(DP_OP_424J2_126_3477_n2440) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1669 ( .A1(DP_OP_424J2_126_3477_n2471), .A2(
        DP_OP_424J2_126_3477_n2475), .Y(DP_OP_424J2_126_3477_n2439) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1668 ( .A1(DP_OP_422J2_124_3477_n2164), .A2(
        DP_OP_424J2_126_3477_n2475), .Y(DP_OP_424J2_126_3477_n2438) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1667 ( .A1(DP_OP_425J2_127_3477_n2296), .A2(
        DP_OP_424J2_126_3477_n2475), .Y(DP_OP_424J2_126_3477_n2437) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1666 ( .A1(DP_OP_423J2_125_3477_n2554), .A2(
        DP_OP_424J2_126_3477_n2475), .Y(DP_OP_424J2_126_3477_n2436) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1665 ( .A1(DP_OP_423J2_125_3477_n2553), 
        .A2(DP_OP_424J2_126_3477_n2475), .Y(DP_OP_424J2_126_3477_n2435) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1646 ( .A1(DP_OP_425J2_127_3477_n2339), 
        .A2(DP_OP_423J2_125_3477_n2432), .Y(DP_OP_424J2_126_3477_n2416) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1645 ( .A1(DP_OP_424J2_126_3477_n2423), .A2(
        DP_OP_425J2_127_3477_n2434), .Y(DP_OP_424J2_126_3477_n2415) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1638 ( .A1(DP_OP_423J2_125_3477_n2510), 
        .A2(DP_OP_425J2_127_3477_n2433), .Y(DP_OP_424J2_126_3477_n2408) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1637 ( .A1(DP_OP_424J2_126_3477_n2423), .A2(
        DP_OP_425J2_127_3477_n2433), .Y(DP_OP_424J2_126_3477_n2407) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1630 ( .A1(DP_OP_423J2_125_3477_n2510), 
        .A2(DP_OP_424J2_126_3477_n2432), .Y(DP_OP_424J2_126_3477_n2400) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1629 ( .A1(DP_OP_424J2_126_3477_n2423), .A2(
        DP_OP_424J2_126_3477_n2432), .Y(DP_OP_424J2_126_3477_n2399) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1628 ( .A1(DP_OP_424J2_126_3477_n2430), .A2(
        DP_OP_423J2_125_3477_n2429), .Y(DP_OP_424J2_126_3477_n2398) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1627 ( .A1(DP_OP_422J2_124_3477_n2211), .A2(
        DP_OP_425J2_127_3477_n2431), .Y(DP_OP_424J2_126_3477_n2397) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1626 ( .A1(DP_OP_424J2_126_3477_n2428), .A2(
        DP_OP_425J2_127_3477_n2431), .Y(DP_OP_424J2_126_3477_n2396) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1625 ( .A1(DP_OP_425J2_127_3477_n2342), .A2(
        DP_OP_423J2_125_3477_n2429), .Y(DP_OP_424J2_126_3477_n2395) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1624 ( .A1(DP_OP_425J2_127_3477_n2341), .A2(
        DP_OP_423J2_125_3477_n2429), .Y(DP_OP_424J2_126_3477_n2394) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1623 ( .A1(DP_OP_425J2_127_3477_n2340), .A2(
        DP_OP_423J2_125_3477_n2429), .Y(DP_OP_424J2_126_3477_n2393) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1622 ( .A1(DP_OP_425J2_127_3477_n2339), .A2(
        DP_OP_425J2_127_3477_n2431), .Y(DP_OP_424J2_126_3477_n2392) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1621 ( .A1(DP_OP_424J2_126_3477_n2423), 
        .A2(DP_OP_423J2_125_3477_n2429), .Y(DP_OP_424J2_126_3477_n2391) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1601 ( .A1(DP_OP_422J2_124_3477_n2249), .A2(
        DP_OP_424J2_126_3477_n2390), .Y(DP_OP_424J2_126_3477_n2371) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1594 ( .A1(DP_OP_422J2_124_3477_n2250), 
        .A2(DP_OP_424J2_126_3477_n2389), .Y(DP_OP_424J2_126_3477_n2364) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1593 ( .A1(DP_OP_422J2_124_3477_n2249), .A2(
        DP_OP_424J2_126_3477_n2389), .Y(DP_OP_424J2_126_3477_n2363) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1586 ( .A1(DP_OP_422J2_124_3477_n2250), 
        .A2(DP_OP_424J2_126_3477_n2388), .Y(DP_OP_424J2_126_3477_n2356) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1585 ( .A1(DP_OP_422J2_124_3477_n2249), .A2(
        DP_OP_424J2_126_3477_n2388), .Y(DP_OP_424J2_126_3477_n2355) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1584 ( .A1(DP_OP_424J2_126_3477_n2386), .A2(
        DP_OP_424J2_126_3477_n2387), .Y(DP_OP_424J2_126_3477_n1579) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1583 ( .A1(DP_OP_424J2_126_3477_n2385), .A2(
        DP_OP_424J2_126_3477_n2387), .Y(DP_OP_424J2_126_3477_n2354) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1582 ( .A1(DP_OP_424J2_126_3477_n2384), .A2(
        DP_OP_424J2_126_3477_n2387), .Y(DP_OP_424J2_126_3477_n2353) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1581 ( .A1(DP_OP_424J2_126_3477_n2383), .A2(
        DP_OP_424J2_126_3477_n2387), .Y(DP_OP_424J2_126_3477_n2352) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1580 ( .A1(DP_OP_424J2_126_3477_n2382), .A2(
        DP_OP_424J2_126_3477_n2387), .Y(DP_OP_424J2_126_3477_n2351) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1579 ( .A1(DP_OP_424J2_126_3477_n2381), .A2(
        DP_OP_424J2_126_3477_n2387), .Y(DP_OP_424J2_126_3477_n671) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1578 ( .A1(DP_OP_422J2_124_3477_n2250), .A2(
        DP_OP_424J2_126_3477_n2387), .Y(DP_OP_424J2_126_3477_n2350) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1577 ( .A1(DP_OP_422J2_124_3477_n2249), 
        .A2(DP_OP_424J2_126_3477_n2387), .Y(DP_OP_424J2_126_3477_n361) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1558 ( .A1(DP_OP_424J2_126_3477_n2339), 
        .A2(DP_OP_424J2_126_3477_n2349), .Y(DP_OP_424J2_126_3477_n2331) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1557 ( .A1(DP_OP_424J2_126_3477_n2338), .A2(
        DP_OP_424J2_126_3477_n2349), .Y(DP_OP_424J2_126_3477_n2330) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1550 ( .A1(DP_OP_424J2_126_3477_n2339), 
        .A2(DP_OP_423J2_125_3477_n2343), .Y(DP_OP_424J2_126_3477_n2323) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1549 ( .A1(DP_OP_424J2_126_3477_n2338), .A2(
        DP_OP_422J2_124_3477_n2347), .Y(DP_OP_424J2_126_3477_n2322) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1542 ( .A1(DP_OP_424J2_126_3477_n2339), 
        .A2(DP_OP_425J2_127_3477_n2347), .Y(DP_OP_424J2_126_3477_n2315) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1541 ( .A1(DP_OP_424J2_126_3477_n2338), .A2(
        n448), .Y(DP_OP_424J2_126_3477_n2314) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1540 ( .A1(DP_OP_422J2_124_3477_n2520), .A2(
        DP_OP_425J2_127_3477_n2346), .Y(DP_OP_424J2_126_3477_n2313) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1539 ( .A1(DP_OP_424J2_126_3477_n2344), .A2(
        DP_OP_425J2_127_3477_n2346), .Y(DP_OP_424J2_126_3477_n2312) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1538 ( .A1(DP_OP_425J2_127_3477_n2384), .A2(
        DP_OP_422J2_124_3477_n2345), .Y(DP_OP_424J2_126_3477_n2311) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1537 ( .A1(DP_OP_424J2_126_3477_n2342), .A2(
        DP_OP_422J2_124_3477_n2345), .Y(DP_OP_424J2_126_3477_n2310) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1536 ( .A1(DP_OP_424J2_126_3477_n2341), .A2(
        DP_OP_425J2_127_3477_n2346), .Y(DP_OP_424J2_126_3477_n2309) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1535 ( .A1(DP_OP_423J2_125_3477_n2247), .A2(
        DP_OP_422J2_124_3477_n2345), .Y(DP_OP_424J2_126_3477_n2308) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1534 ( .A1(DP_OP_424J2_126_3477_n2339), .A2(
        DP_OP_425J2_127_3477_n2346), .Y(DP_OP_424J2_126_3477_n2307) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1533 ( .A1(DP_OP_424J2_126_3477_n2338), 
        .A2(DP_OP_425J2_127_3477_n2346), .Y(DP_OP_424J2_126_3477_n2306) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1514 ( .A1(DP_OP_425J2_127_3477_n2424), 
        .A2(n446), .Y(DP_OP_424J2_126_3477_n2287) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1513 ( .A1(DP_OP_425J2_127_3477_n2423), .A2(
        n446), .Y(DP_OP_424J2_126_3477_n2286) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1506 ( .A1(DP_OP_425J2_127_3477_n2424), 
        .A2(DP_OP_424J2_126_3477_n2304), .Y(DP_OP_424J2_126_3477_n2279) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1505 ( .A1(DP_OP_425J2_127_3477_n2423), .A2(
        DP_OP_424J2_126_3477_n2304), .Y(DP_OP_424J2_126_3477_n2278) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1498 ( .A1(DP_OP_425J2_127_3477_n2424), 
        .A2(n445), .Y(DP_OP_424J2_126_3477_n2271) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1497 ( .A1(DP_OP_425J2_127_3477_n2423), .A2(
        n445), .Y(DP_OP_424J2_126_3477_n2270) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1496 ( .A1(DP_OP_425J2_127_3477_n2430), .A2(
        DP_OP_424J2_126_3477_n2302), .Y(DP_OP_424J2_126_3477_n2269) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1495 ( .A1(DP_OP_425J2_127_3477_n2429), .A2(
        DP_OP_424J2_126_3477_n2302), .Y(DP_OP_424J2_126_3477_n2268) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1494 ( .A1(DP_OP_425J2_127_3477_n2428), .A2(
        DP_OP_424J2_126_3477_n2302), .Y(DP_OP_424J2_126_3477_n2267) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1493 ( .A1(DP_OP_423J2_125_3477_n2205), .A2(
        DP_OP_424J2_126_3477_n2302), .Y(DP_OP_424J2_126_3477_n2266) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1492 ( .A1(DP_OP_423J2_125_3477_n2204), .A2(
        DP_OP_424J2_126_3477_n2302), .Y(DP_OP_424J2_126_3477_n2265) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1491 ( .A1(DP_OP_424J2_126_3477_n2296), .A2(
        DP_OP_424J2_126_3477_n2302), .Y(DP_OP_424J2_126_3477_n2264) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1490 ( .A1(DP_OP_422J2_124_3477_n2558), .A2(
        DP_OP_424J2_126_3477_n2302), .Y(DP_OP_424J2_126_3477_n2263) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1489 ( .A1(DP_OP_425J2_127_3477_n2423), 
        .A2(DP_OP_424J2_126_3477_n2302), .Y(DP_OP_424J2_126_3477_n2262) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1471 ( .A1(DP_OP_422J2_124_3477_n2603), 
        .A2(DP_OP_423J2_125_3477_n2256), .Y(DP_OP_424J2_126_3477_n2244) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1470 ( .A1(DP_OP_422J2_124_3477_n2602), 
        .A2(DP_OP_425J2_127_3477_n2261), .Y(DP_OP_424J2_126_3477_n2243) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1469 ( .A1(DP_OP_422J2_124_3477_n2601), .A2(
        DP_OP_425J2_127_3477_n2261), .Y(DP_OP_424J2_126_3477_n2242) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1461 ( .A1(DP_OP_422J2_124_3477_n2601), .A2(
        DP_OP_424J2_126_3477_n2260), .Y(DP_OP_424J2_126_3477_n2234) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1454 ( .A1(DP_OP_422J2_124_3477_n2602), 
        .A2(DP_OP_422J2_124_3477_n2258), .Y(DP_OP_424J2_126_3477_n2227) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1453 ( .A1(DP_OP_422J2_124_3477_n2601), .A2(
        DP_OP_422J2_124_3477_n2258), .Y(DP_OP_424J2_126_3477_n2226) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1452 ( .A1(DP_OP_422J2_124_3477_n2608), .A2(
        DP_OP_424J2_126_3477_n2258), .Y(DP_OP_424J2_126_3477_n2225) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1451 ( .A1(DP_OP_422J2_124_3477_n2607), .A2(
        DP_OP_424J2_126_3477_n2258), .Y(DP_OP_424J2_126_3477_n2224) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1450 ( .A1(DP_OP_422J2_124_3477_n2606), .A2(
        DP_OP_424J2_126_3477_n2258), .Y(DP_OP_424J2_126_3477_n2223) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1449 ( .A1(DP_OP_422J2_124_3477_n2605), .A2(
        DP_OP_424J2_126_3477_n2258), .Y(DP_OP_424J2_126_3477_n2222) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1448 ( .A1(DP_OP_422J2_124_3477_n2604), .A2(
        DP_OP_424J2_126_3477_n2258), .Y(DP_OP_424J2_126_3477_n2221) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1447 ( .A1(DP_OP_422J2_124_3477_n2603), .A2(
        DP_OP_424J2_126_3477_n2258), .Y(DP_OP_424J2_126_3477_n2220) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1446 ( .A1(DP_OP_422J2_124_3477_n2602), .A2(
        DP_OP_424J2_126_3477_n2258), .Y(DP_OP_424J2_126_3477_n2219) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1445 ( .A1(DP_OP_422J2_124_3477_n2601), 
        .A2(DP_OP_424J2_126_3477_n2258), .Y(DP_OP_424J2_126_3477_n2218) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1426 ( .A1(DP_OP_422J2_124_3477_n2646), 
        .A2(DP_OP_425J2_127_3477_n2217), .Y(DP_OP_424J2_126_3477_n2199) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1425 ( .A1(DP_OP_425J2_127_3477_n2511), .A2(
        DP_OP_423J2_125_3477_n2212), .Y(DP_OP_424J2_126_3477_n2198) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1417 ( .A1(DP_OP_425J2_127_3477_n2511), .A2(
        DP_OP_424J2_126_3477_n2216), .Y(DP_OP_424J2_126_3477_n2190) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1410 ( .A1(DP_OP_422J2_124_3477_n2646), 
        .A2(n443), .Y(DP_OP_424J2_126_3477_n2183) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1409 ( .A1(DP_OP_425J2_127_3477_n2511), .A2(
        n443), .Y(DP_OP_424J2_126_3477_n2182) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1408 ( .A1(DP_OP_422J2_124_3477_n2652), .A2(
        DP_OP_423J2_125_3477_n2209), .Y(DP_OP_424J2_126_3477_n2181) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1407 ( .A1(DP_OP_424J2_126_3477_n2212), .A2(
        DP_OP_425J2_127_3477_n2214), .Y(DP_OP_424J2_126_3477_n2180) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1406 ( .A1(DP_OP_424J2_126_3477_n2211), .A2(
        DP_OP_423J2_125_3477_n2209), .Y(DP_OP_424J2_126_3477_n2179) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1405 ( .A1(DP_OP_422J2_124_3477_n2649), .A2(
        DP_OP_425J2_127_3477_n2214), .Y(DP_OP_424J2_126_3477_n2178) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1404 ( .A1(DP_OP_422J2_124_3477_n2648), .A2(
        DP_OP_423J2_125_3477_n2209), .Y(DP_OP_424J2_126_3477_n2177) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1403 ( .A1(DP_OP_423J2_125_3477_n2115), .A2(
        DP_OP_425J2_127_3477_n2214), .Y(DP_OP_424J2_126_3477_n2176) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1402 ( .A1(DP_OP_423J2_125_3477_n2114), .A2(
        DP_OP_425J2_127_3477_n2214), .Y(DP_OP_424J2_126_3477_n2175) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1401 ( .A1(DP_OP_422J2_124_3477_n2645), 
        .A2(DP_OP_423J2_125_3477_n2209), .Y(DP_OP_424J2_126_3477_n2174) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1382 ( .A1(DP_OP_424J2_126_3477_n2163), 
        .A2(DP_OP_424J2_126_3477_n2173), .Y(DP_OP_424J2_126_3477_n2155) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1381 ( .A1(DP_OP_422J2_124_3477_n2689), .A2(
        DP_OP_424J2_126_3477_n2173), .Y(DP_OP_424J2_126_3477_n2154) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1374 ( .A1(DP_OP_424J2_126_3477_n2163), 
        .A2(DP_OP_422J2_124_3477_n2171), .Y(DP_OP_424J2_126_3477_n2147) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1373 ( .A1(DP_OP_422J2_124_3477_n2689), .A2(
        DP_OP_425J2_127_3477_n2172), .Y(DP_OP_424J2_126_3477_n2146) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1366 ( .A1(DP_OP_424J2_126_3477_n2163), 
        .A2(DP_OP_424J2_126_3477_n2171), .Y(DP_OP_424J2_126_3477_n2139) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1365 ( .A1(DP_OP_425J2_127_3477_n2555), .A2(
        DP_OP_424J2_126_3477_n2171), .Y(DP_OP_424J2_126_3477_n2138) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1364 ( .A1(DP_OP_423J2_125_3477_n2076), .A2(
        DP_OP_424J2_126_3477_n2170), .Y(DP_OP_424J2_126_3477_n2137) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1363 ( .A1(DP_OP_424J2_126_3477_n2168), .A2(
        DP_OP_424J2_126_3477_n2170), .Y(DP_OP_424J2_126_3477_n2136) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1362 ( .A1(DP_OP_423J2_125_3477_n2074), .A2(
        DP_OP_424J2_126_3477_n2170), .Y(DP_OP_424J2_126_3477_n2135) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1361 ( .A1(DP_OP_423J2_125_3477_n2073), .A2(
        DP_OP_424J2_126_3477_n2170), .Y(DP_OP_424J2_126_3477_n2134) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1360 ( .A1(DP_OP_422J2_124_3477_n2692), .A2(
        DP_OP_424J2_126_3477_n2170), .Y(DP_OP_424J2_126_3477_n2133) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1359 ( .A1(DP_OP_424J2_126_3477_n2164), .A2(
        DP_OP_424J2_126_3477_n2170), .Y(DP_OP_424J2_126_3477_n2132) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1358 ( .A1(DP_OP_424J2_126_3477_n2163), .A2(
        DP_OP_424J2_126_3477_n2170), .Y(DP_OP_424J2_126_3477_n2131) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1357 ( .A1(DP_OP_422J2_124_3477_n2689), 
        .A2(DP_OP_424J2_126_3477_n2170), .Y(DP_OP_424J2_126_3477_n2130) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1338 ( .A1(DP_OP_424J2_126_3477_n2119), 
        .A2(DP_OP_424J2_126_3477_n2129), .Y(DP_OP_424J2_126_3477_n2111) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1337 ( .A1(DP_OP_424J2_126_3477_n2118), .A2(
        DP_OP_424J2_126_3477_n2129), .Y(DP_OP_424J2_126_3477_n2110) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1329 ( .A1(DP_OP_424J2_126_3477_n2118), .A2(
        n440), .Y(DP_OP_424J2_126_3477_n2102) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1322 ( .A1(DP_OP_424J2_126_3477_n2119), 
        .A2(DP_OP_424J2_126_3477_n2127), .Y(DP_OP_424J2_126_3477_n2095) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1321 ( .A1(DP_OP_424J2_126_3477_n2118), .A2(
        DP_OP_424J2_126_3477_n2127), .Y(DP_OP_424J2_126_3477_n2094) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1320 ( .A1(DP_OP_424J2_126_3477_n2125), .A2(
        DP_OP_424J2_126_3477_n2126), .Y(DP_OP_424J2_126_3477_n2093) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1319 ( .A1(DP_OP_424J2_126_3477_n2124), .A2(
        DP_OP_424J2_126_3477_n2126), .Y(DP_OP_424J2_126_3477_n2092) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1318 ( .A1(DP_OP_422J2_124_3477_n2736), .A2(
        DP_OP_424J2_126_3477_n2126), .Y(DP_OP_424J2_126_3477_n2091) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1317 ( .A1(DP_OP_423J2_125_3477_n2029), .A2(
        DP_OP_424J2_126_3477_n2126), .Y(DP_OP_424J2_126_3477_n2090) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1316 ( .A1(DP_OP_423J2_125_3477_n2028), .A2(
        DP_OP_424J2_126_3477_n2126), .Y(DP_OP_424J2_126_3477_n2089) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1315 ( .A1(DP_OP_424J2_126_3477_n2120), .A2(
        DP_OP_424J2_126_3477_n2126), .Y(DP_OP_424J2_126_3477_n2088) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1314 ( .A1(DP_OP_424J2_126_3477_n2119), .A2(
        DP_OP_424J2_126_3477_n2126), .Y(DP_OP_424J2_126_3477_n2087) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1313 ( .A1(DP_OP_424J2_126_3477_n2118), 
        .A2(DP_OP_424J2_126_3477_n2126), .Y(DP_OP_424J2_126_3477_n2086) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1294 ( .A1(DP_OP_422J2_124_3477_n2776), 
        .A2(DP_OP_424J2_126_3477_n2085), .Y(DP_OP_424J2_126_3477_n2067) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1293 ( .A1(DP_OP_424J2_126_3477_n2074), .A2(
        DP_OP_424J2_126_3477_n2085), .Y(DP_OP_424J2_126_3477_n2066) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1286 ( .A1(DP_OP_425J2_127_3477_n2644), 
        .A2(DP_OP_424J2_126_3477_n2084), .Y(DP_OP_424J2_126_3477_n2059) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1285 ( .A1(DP_OP_424J2_126_3477_n2074), .A2(
        DP_OP_424J2_126_3477_n2084), .Y(DP_OP_424J2_126_3477_n2058) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1278 ( .A1(DP_OP_425J2_127_3477_n2644), 
        .A2(n447), .Y(DP_OP_424J2_126_3477_n2051) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1277 ( .A1(DP_OP_424J2_126_3477_n2074), .A2(
        n447), .Y(DP_OP_424J2_126_3477_n2050) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1276 ( .A1(DP_OP_425J2_127_3477_n2650), .A2(
        DP_OP_424J2_126_3477_n2082), .Y(DP_OP_424J2_126_3477_n2049) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1275 ( .A1(DP_OP_425J2_127_3477_n2649), .A2(
        DP_OP_424J2_126_3477_n2082), .Y(DP_OP_424J2_126_3477_n2048) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1274 ( .A1(DP_OP_423J2_125_3477_n1986), .A2(
        DP_OP_424J2_126_3477_n2082), .Y(DP_OP_424J2_126_3477_n2047) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1273 ( .A1(DP_OP_424J2_126_3477_n2078), .A2(
        DP_OP_424J2_126_3477_n2082), .Y(DP_OP_424J2_126_3477_n2046) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1272 ( .A1(DP_OP_424J2_126_3477_n2077), .A2(
        DP_OP_424J2_126_3477_n2082), .Y(DP_OP_424J2_126_3477_n2045) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1271 ( .A1(DP_OP_422J2_124_3477_n2777), .A2(
        DP_OP_424J2_126_3477_n2082), .Y(DP_OP_424J2_126_3477_n2044) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1270 ( .A1(DP_OP_422J2_124_3477_n2776), .A2(
        DP_OP_424J2_126_3477_n2082), .Y(DP_OP_424J2_126_3477_n2043) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1269 ( .A1(DP_OP_424J2_126_3477_n2074), 
        .A2(DP_OP_424J2_126_3477_n2082), .Y(DP_OP_424J2_126_3477_n2042) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1250 ( .A1(DP_OP_422J2_124_3477_n2820), 
        .A2(DP_OP_424J2_126_3477_n2041), .Y(DP_OP_424J2_126_3477_n2023) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1249 ( .A1(DP_OP_422J2_124_3477_n2819), .A2(
        DP_OP_424J2_126_3477_n2041), .Y(DP_OP_424J2_126_3477_n2022) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1242 ( .A1(DP_OP_422J2_124_3477_n2820), 
        .A2(DP_OP_424J2_126_3477_n2040), .Y(DP_OP_424J2_126_3477_n2015) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1241 ( .A1(DP_OP_422J2_124_3477_n2819), .A2(
        DP_OP_424J2_126_3477_n2040), .Y(DP_OP_424J2_126_3477_n2014) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1234 ( .A1(DP_OP_422J2_124_3477_n2820), 
        .A2(DP_OP_424J2_126_3477_n2039), .Y(DP_OP_424J2_126_3477_n2007) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1233 ( .A1(DP_OP_422J2_124_3477_n2819), .A2(
        DP_OP_424J2_126_3477_n2039), .Y(DP_OP_424J2_126_3477_n2006) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1232 ( .A1(DP_OP_424J2_126_3477_n2037), .A2(
        DP_OP_424J2_126_3477_n2038), .Y(DP_OP_424J2_126_3477_n2005) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1231 ( .A1(DP_OP_422J2_124_3477_n2825), .A2(
        DP_OP_424J2_126_3477_n2038), .Y(DP_OP_424J2_126_3477_n2004) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1230 ( .A1(DP_OP_424J2_126_3477_n2035), .A2(
        DP_OP_424J2_126_3477_n2038), .Y(DP_OP_424J2_126_3477_n2003) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1229 ( .A1(DP_OP_424J2_126_3477_n2034), .A2(
        DP_OP_424J2_126_3477_n2038), .Y(DP_OP_424J2_126_3477_n2002) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1228 ( .A1(DP_OP_424J2_126_3477_n2033), .A2(
        DP_OP_424J2_126_3477_n2038), .Y(DP_OP_424J2_126_3477_n2001) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1227 ( .A1(DP_OP_424J2_126_3477_n2032), .A2(
        DP_OP_424J2_126_3477_n2038), .Y(DP_OP_424J2_126_3477_n2000) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1226 ( .A1(DP_OP_422J2_124_3477_n2820), .A2(
        DP_OP_424J2_126_3477_n2038), .Y(DP_OP_424J2_126_3477_n1999) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1225 ( .A1(DP_OP_422J2_124_3477_n2819), 
        .A2(DP_OP_424J2_126_3477_n2038), .Y(DP_OP_424J2_126_3477_n1998) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1206 ( .A1(DP_OP_425J2_127_3477_n2732), 
        .A2(DP_OP_423J2_125_3477_n1992), .Y(DP_OP_424J2_126_3477_n1979) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1205 ( .A1(DP_OP_424J2_126_3477_n1986), .A2(
        DP_OP_423J2_125_3477_n1992), .Y(DP_OP_424J2_126_3477_n1978) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1197 ( .A1(DP_OP_424J2_126_3477_n1986), .A2(
        DP_OP_424J2_126_3477_n1996), .Y(DP_OP_424J2_126_3477_n1970) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1190 ( .A1(DP_OP_425J2_127_3477_n2732), 
        .A2(DP_OP_424J2_126_3477_n1995), .Y(DP_OP_424J2_126_3477_n1963) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1189 ( .A1(DP_OP_424J2_126_3477_n1986), .A2(
        DP_OP_424J2_126_3477_n1995), .Y(DP_OP_424J2_126_3477_n1962) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1188 ( .A1(DP_OP_425J2_127_3477_n2738), .A2(
        DP_OP_424J2_126_3477_n1994), .Y(DP_OP_424J2_126_3477_n1961) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1187 ( .A1(DP_OP_423J2_125_3477_n1899), .A2(
        DP_OP_424J2_126_3477_n1994), .Y(DP_OP_424J2_126_3477_n1960) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1186 ( .A1(DP_OP_423J2_125_3477_n1898), .A2(
        DP_OP_424J2_126_3477_n1994), .Y(DP_OP_424J2_126_3477_n1959) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1185 ( .A1(DP_OP_423J2_125_3477_n1897), .A2(
        DP_OP_424J2_126_3477_n1994), .Y(DP_OP_424J2_126_3477_n1958) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1184 ( .A1(DP_OP_423J2_125_3477_n1896), .A2(
        DP_OP_424J2_126_3477_n1994), .Y(DP_OP_424J2_126_3477_n1957) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1183 ( .A1(DP_OP_424J2_126_3477_n1988), .A2(
        DP_OP_424J2_126_3477_n1994), .Y(DP_OP_424J2_126_3477_n1956) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1182 ( .A1(DP_OP_425J2_127_3477_n2732), .A2(
        DP_OP_424J2_126_3477_n1994), .Y(DP_OP_424J2_126_3477_n1955) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1181 ( .A1(DP_OP_424J2_126_3477_n1986), 
        .A2(DP_OP_424J2_126_3477_n1994), .Y(DP_OP_424J2_126_3477_n1954) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1162 ( .A1(DP_OP_423J2_125_3477_n1850), 
        .A2(DP_OP_424J2_126_3477_n1953), .Y(DP_OP_424J2_126_3477_n1935) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1161 ( .A1(DP_OP_424J2_126_3477_n1942), .A2(
        DP_OP_424J2_126_3477_n1953), .Y(DP_OP_424J2_126_3477_n1934) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1154 ( .A1(DP_OP_423J2_125_3477_n1850), 
        .A2(DP_OP_424J2_126_3477_n1952), .Y(DP_OP_424J2_126_3477_n1927) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1153 ( .A1(DP_OP_424J2_126_3477_n1942), .A2(
        DP_OP_424J2_126_3477_n1952), .Y(DP_OP_424J2_126_3477_n1926) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1145 ( .A1(DP_OP_424J2_126_3477_n1942), .A2(
        DP_OP_425J2_127_3477_n1951), .Y(DP_OP_424J2_126_3477_n1918) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1144 ( .A1(DP_OP_424J2_126_3477_n1949), .A2(
        DP_OP_424J2_126_3477_n1950), .Y(DP_OP_424J2_126_3477_n1917) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1143 ( .A1(DP_OP_424J2_126_3477_n1948), .A2(
        DP_OP_424J2_126_3477_n1950), .Y(DP_OP_424J2_126_3477_n1916) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1142 ( .A1(DP_OP_422J2_124_3477_n2912), .A2(
        DP_OP_424J2_126_3477_n1950), .Y(DP_OP_424J2_126_3477_n1915) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1141 ( .A1(DP_OP_425J2_127_3477_n2779), .A2(
        DP_OP_424J2_126_3477_n1950), .Y(DP_OP_424J2_126_3477_n1914) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1140 ( .A1(DP_OP_425J2_127_3477_n2778), .A2(
        DP_OP_424J2_126_3477_n1950), .Y(DP_OP_424J2_126_3477_n1913) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1139 ( .A1(DP_OP_425J2_127_3477_n2777), .A2(
        DP_OP_424J2_126_3477_n1950), .Y(DP_OP_424J2_126_3477_n1912) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1138 ( .A1(DP_OP_423J2_125_3477_n1850), .A2(
        DP_OP_424J2_126_3477_n1950), .Y(DP_OP_424J2_126_3477_n1911) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1137 ( .A1(DP_OP_424J2_126_3477_n1942), 
        .A2(DP_OP_424J2_126_3477_n1950), .Y(DP_OP_424J2_126_3477_n1910) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1118 ( .A1(DP_OP_425J2_127_3477_n2820), 
        .A2(DP_OP_424J2_126_3477_n1909), .Y(DP_OP_424J2_126_3477_n1891) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1117 ( .A1(DP_OP_424J2_126_3477_n1898), .A2(
        DP_OP_424J2_126_3477_n1909), .Y(DP_OP_424J2_126_3477_n1890) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1110 ( .A1(DP_OP_425J2_127_3477_n2820), 
        .A2(DP_OP_424J2_126_3477_n1908), .Y(DP_OP_424J2_126_3477_n1883) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1109 ( .A1(DP_OP_424J2_126_3477_n1898), .A2(
        DP_OP_424J2_126_3477_n1908), .Y(DP_OP_424J2_126_3477_n1882) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1102 ( .A1(DP_OP_425J2_127_3477_n2820), 
        .A2(DP_OP_424J2_126_3477_n1907), .Y(DP_OP_424J2_126_3477_n1875) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1101 ( .A1(DP_OP_424J2_126_3477_n1898), .A2(
        DP_OP_424J2_126_3477_n1907), .Y(DP_OP_424J2_126_3477_n1874) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1100 ( .A1(DP_OP_425J2_127_3477_n2826), .A2(
        DP_OP_424J2_126_3477_n1906), .Y(DP_OP_424J2_126_3477_n1873) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1099 ( .A1(DP_OP_424J2_126_3477_n1904), .A2(
        DP_OP_424J2_126_3477_n1906), .Y(DP_OP_424J2_126_3477_n1872) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1098 ( .A1(DP_OP_424J2_126_3477_n1903), .A2(
        DP_OP_424J2_126_3477_n1906), .Y(DP_OP_424J2_126_3477_n1871) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1097 ( .A1(DP_OP_425J2_127_3477_n2823), .A2(
        DP_OP_424J2_126_3477_n1906), .Y(DP_OP_424J2_126_3477_n1870) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1096 ( .A1(DP_OP_424J2_126_3477_n1901), .A2(
        DP_OP_424J2_126_3477_n1906), .Y(DP_OP_424J2_126_3477_n1869) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1095 ( .A1(DP_OP_425J2_127_3477_n2821), .A2(
        DP_OP_424J2_126_3477_n1906), .Y(DP_OP_424J2_126_3477_n1868) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1094 ( .A1(DP_OP_425J2_127_3477_n2820), .A2(
        DP_OP_424J2_126_3477_n1906), .Y(DP_OP_424J2_126_3477_n1867) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1093 ( .A1(DP_OP_424J2_126_3477_n1898), 
        .A2(DP_OP_424J2_126_3477_n1906), .Y(DP_OP_424J2_126_3477_n1866) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1074 ( .A1(DP_OP_425J2_127_3477_n2864), 
        .A2(DP_OP_424J2_126_3477_n1865), .Y(DP_OP_424J2_126_3477_n1847) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1073 ( .A1(DP_OP_424J2_126_3477_n1854), .A2(
        DP_OP_424J2_126_3477_n1865), .Y(DP_OP_424J2_126_3477_n1846) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1066 ( .A1(DP_OP_425J2_127_3477_n2864), 
        .A2(DP_OP_425J2_127_3477_n1864), .Y(DP_OP_424J2_126_3477_n1839) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1065 ( .A1(DP_OP_424J2_126_3477_n1854), .A2(
        DP_OP_423J2_125_3477_n1859), .Y(DP_OP_424J2_126_3477_n1838) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1058 ( .A1(DP_OP_425J2_127_3477_n2864), 
        .A2(DP_OP_425J2_127_3477_n1863), .Y(DP_OP_424J2_126_3477_n1831) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1057 ( .A1(DP_OP_424J2_126_3477_n1854), .A2(
        DP_OP_425J2_127_3477_n1863), .Y(DP_OP_424J2_126_3477_n1830) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1056 ( .A1(DP_OP_425J2_127_3477_n2870), .A2(
        DP_OP_424J2_126_3477_n1862), .Y(DP_OP_424J2_126_3477_n1829) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1055 ( .A1(DP_OP_425J2_127_3477_n2869), .A2(
        DP_OP_424J2_126_3477_n1862), .Y(DP_OP_424J2_126_3477_n1828) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1054 ( .A1(DP_OP_425J2_127_3477_n2868), .A2(
        DP_OP_424J2_126_3477_n1862), .Y(DP_OP_424J2_126_3477_n1827) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1053 ( .A1(DP_OP_424J2_126_3477_n1858), .A2(
        DP_OP_424J2_126_3477_n1862), .Y(DP_OP_424J2_126_3477_n1826) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1052 ( .A1(DP_OP_424J2_126_3477_n1857), .A2(
        DP_OP_424J2_126_3477_n1862), .Y(DP_OP_424J2_126_3477_n1825) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1051 ( .A1(DP_OP_425J2_127_3477_n2865), .A2(
        DP_OP_424J2_126_3477_n1862), .Y(DP_OP_424J2_126_3477_n1824) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1050 ( .A1(DP_OP_425J2_127_3477_n2864), .A2(
        DP_OP_424J2_126_3477_n1862), .Y(DP_OP_424J2_126_3477_n1823) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1049 ( .A1(DP_OP_424J2_126_3477_n1854), 
        .A2(DP_OP_424J2_126_3477_n1862), .Y(DP_OP_424J2_126_3477_n1822) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1001 ( .A1(n417), .A2(
        DP_OP_425J2_127_3477_n2), .Y(DP_OP_424J2_126_3477_n189) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U999 ( .A1(n299), .A2(n338), .Y(
        DP_OP_424J2_126_3477_n181) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U998 ( .A1(n427), .A2(
        DP_OP_423J2_125_3477_n2), .Y(DP_OP_424J2_126_3477_n179) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U997 ( .A1(n416), .A2(
        DP_OP_424J2_126_3477_n2), .Y(DP_OP_424J2_126_3477_n177) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U996 ( .A1(n379), .A2(n342), .Y(
        DP_OP_424J2_126_3477_n175) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U995 ( .A1(n419), .A2(n340), .Y(
        DP_OP_424J2_126_3477_n173) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U994 ( .A1(n426), .A2(n341), .Y(
        DP_OP_424J2_126_3477_n171) );
  HADDX1_HVT DP_OP_424J2_126_3477_U983 ( .A0(DP_OP_424J2_126_3477_n2642), .B0(
        DP_OP_424J2_126_3477_n2730), .C1(DP_OP_424J2_126_3477_n1771), .SO(
        DP_OP_424J2_126_3477_n1772) );
  FADDX1_HVT DP_OP_424J2_126_3477_U982 ( .A(DP_OP_424J2_126_3477_n2598), .B(
        DP_OP_424J2_126_3477_n1788), .CI(DP_OP_424J2_126_3477_n2293), .CO(
        DP_OP_424J2_126_3477_n1769), .S(DP_OP_424J2_126_3477_n1770) );
  FADDX1_HVT DP_OP_424J2_126_3477_U981 ( .A(DP_OP_424J2_126_3477_n1853), .B(
        DP_OP_424J2_126_3477_n2029), .CI(DP_OP_424J2_126_3477_n2073), .CO(
        DP_OP_424J2_126_3477_n1767), .S(DP_OP_424J2_126_3477_n1768) );
  FADDX1_HVT DP_OP_424J2_126_3477_U980 ( .A(DP_OP_424J2_126_3477_n2205), .B(
        DP_OP_424J2_126_3477_n1985), .CI(DP_OP_424J2_126_3477_n2510), .CO(
        DP_OP_424J2_126_3477_n1765), .S(DP_OP_424J2_126_3477_n1766) );
  FADDX1_HVT DP_OP_424J2_126_3477_U979 ( .A(DP_OP_424J2_126_3477_n2554), .B(
        DP_OP_424J2_126_3477_n2686), .CI(DP_OP_424J2_126_3477_n2774), .CO(
        DP_OP_424J2_126_3477_n1763), .S(DP_OP_424J2_126_3477_n1764) );
  FADDX1_HVT DP_OP_424J2_126_3477_U978 ( .A(DP_OP_424J2_126_3477_n2422), .B(
        DP_OP_424J2_126_3477_n2337), .CI(DP_OP_424J2_126_3477_n2862), .CO(
        DP_OP_424J2_126_3477_n1761), .S(DP_OP_424J2_126_3477_n1762) );
  FADDX1_HVT DP_OP_424J2_126_3477_U977 ( .A(DP_OP_424J2_126_3477_n2466), .B(
        DP_OP_424J2_126_3477_n2117), .CI(DP_OP_424J2_126_3477_n1897), .CO(
        DP_OP_424J2_126_3477_n1759), .S(DP_OP_424J2_126_3477_n1760) );
  FADDX1_HVT DP_OP_424J2_126_3477_U976 ( .A(DP_OP_424J2_126_3477_n1941), .B(
        DP_OP_424J2_126_3477_n2249), .CI(DP_OP_424J2_126_3477_n2906), .CO(
        DP_OP_424J2_126_3477_n1757), .S(DP_OP_424J2_126_3477_n1758) );
  FADDX1_HVT DP_OP_424J2_126_3477_U975 ( .A(DP_OP_424J2_126_3477_n2161), .B(
        DP_OP_424J2_126_3477_n2378), .CI(DP_OP_424J2_126_3477_n2818), .CO(
        DP_OP_424J2_126_3477_n1755), .S(DP_OP_424J2_126_3477_n1756) );
  FADDX1_HVT DP_OP_424J2_126_3477_U974 ( .A(DP_OP_424J2_126_3477_n1772), .B(
        DP_OP_424J2_126_3477_n1762), .CI(DP_OP_424J2_126_3477_n1764), .CO(
        DP_OP_424J2_126_3477_n1753), .S(DP_OP_424J2_126_3477_n1754) );
  FADDX1_HVT DP_OP_424J2_126_3477_U973 ( .A(DP_OP_424J2_126_3477_n1766), .B(
        DP_OP_424J2_126_3477_n1760), .CI(DP_OP_424J2_126_3477_n1768), .CO(
        DP_OP_424J2_126_3477_n1751), .S(DP_OP_424J2_126_3477_n1752) );
  FADDX1_HVT DP_OP_424J2_126_3477_U972 ( .A(DP_OP_424J2_126_3477_n1770), .B(
        DP_OP_424J2_126_3477_n1758), .CI(DP_OP_424J2_126_3477_n1756), .CO(
        DP_OP_424J2_126_3477_n1749), .S(DP_OP_424J2_126_3477_n1750) );
  HADDX1_HVT DP_OP_424J2_126_3477_U971 ( .A0(DP_OP_424J2_126_3477_n2553), .B0(
        DP_OP_424J2_126_3477_n2414), .C1(DP_OP_424J2_126_3477_n1747), .SO(
        DP_OP_424J2_126_3477_n1748) );
  FADDX1_HVT DP_OP_424J2_126_3477_U970 ( .A(DP_OP_424J2_126_3477_n1852), .B(
        DP_OP_424J2_126_3477_n2729), .CI(DP_OP_424J2_126_3477_n2072), .CO(
        DP_OP_424J2_126_3477_n1745), .S(DP_OP_424J2_126_3477_n1746) );
  FADDX1_HVT DP_OP_424J2_126_3477_U969 ( .A(DP_OP_424J2_126_3477_n2336), .B(
        DP_OP_424J2_126_3477_n2153), .CI(DP_OP_424J2_126_3477_n2292), .CO(
        DP_OP_424J2_126_3477_n1743), .S(DP_OP_424J2_126_3477_n1744) );
  FADDX1_HVT DP_OP_424J2_126_3477_U968 ( .A(DP_OP_424J2_126_3477_n2116), .B(
        DP_OP_424J2_126_3477_n1787), .CI(DP_OP_424J2_126_3477_n2509), .CO(
        DP_OP_424J2_126_3477_n1741), .S(DP_OP_424J2_126_3477_n1742) );
  FADDX1_HVT DP_OP_424J2_126_3477_U967 ( .A(DP_OP_424J2_126_3477_n2204), .B(
        DP_OP_424J2_126_3477_n2065), .CI(DP_OP_424J2_126_3477_n2773), .CO(
        DP_OP_424J2_126_3477_n1739), .S(DP_OP_424J2_126_3477_n1740) );
  FADDX1_HVT DP_OP_424J2_126_3477_U966 ( .A(DP_OP_424J2_126_3477_n2465), .B(
        DP_OP_424J2_126_3477_n1984), .CI(DP_OP_424J2_126_3477_n1896), .CO(
        DP_OP_424J2_126_3477_n1737), .S(DP_OP_424J2_126_3477_n1738) );
  FADDX1_HVT DP_OP_424J2_126_3477_U965 ( .A(DP_OP_424J2_126_3477_n2641), .B(
        DP_OP_424J2_126_3477_n2028), .CI(DP_OP_424J2_126_3477_n2861), .CO(
        DP_OP_424J2_126_3477_n1735), .S(DP_OP_424J2_126_3477_n1736) );
  FADDX1_HVT DP_OP_424J2_126_3477_U964 ( .A(DP_OP_424J2_126_3477_n2597), .B(
        DP_OP_424J2_126_3477_n2590), .CI(DP_OP_424J2_126_3477_n2329), .CO(
        DP_OP_424J2_126_3477_n1733), .S(DP_OP_424J2_126_3477_n1734) );
  FADDX1_HVT DP_OP_424J2_126_3477_U963 ( .A(DP_OP_424J2_126_3477_n2421), .B(
        DP_OP_424J2_126_3477_n2634), .CI(DP_OP_424J2_126_3477_n2685), .CO(
        DP_OP_424J2_126_3477_n1731), .S(DP_OP_424J2_126_3477_n1732) );
  FADDX1_HVT DP_OP_424J2_126_3477_U962 ( .A(DP_OP_424J2_126_3477_n1845), .B(
        DP_OP_424J2_126_3477_n2502), .CI(DP_OP_424J2_126_3477_n1940), .CO(
        DP_OP_424J2_126_3477_n1729), .S(DP_OP_424J2_126_3477_n1730) );
  FADDX1_HVT DP_OP_424J2_126_3477_U961 ( .A(DP_OP_424J2_126_3477_n2546), .B(
        DP_OP_424J2_126_3477_n2766), .CI(DP_OP_424J2_126_3477_n2370), .CO(
        DP_OP_424J2_126_3477_n1727), .S(DP_OP_424J2_126_3477_n1728) );
  FADDX1_HVT DP_OP_424J2_126_3477_U960 ( .A(DP_OP_424J2_126_3477_n2854), .B(
        DP_OP_424J2_126_3477_n2458), .CI(DP_OP_424J2_126_3477_n2241), .CO(
        DP_OP_424J2_126_3477_n1725), .S(DP_OP_424J2_126_3477_n1726) );
  FADDX1_HVT DP_OP_424J2_126_3477_U959 ( .A(DP_OP_424J2_126_3477_n2109), .B(
        DP_OP_424J2_126_3477_n2810), .CI(DP_OP_424J2_126_3477_n2197), .CO(
        DP_OP_424J2_126_3477_n1723), .S(DP_OP_424J2_126_3477_n1724) );
  FADDX1_HVT DP_OP_424J2_126_3477_U958 ( .A(DP_OP_424J2_126_3477_n1889), .B(
        DP_OP_424J2_126_3477_n2285), .CI(DP_OP_424J2_126_3477_n1933), .CO(
        DP_OP_424J2_126_3477_n1721), .S(DP_OP_424J2_126_3477_n1722) );
  FADDX1_HVT DP_OP_424J2_126_3477_U957 ( .A(DP_OP_424J2_126_3477_n2678), .B(
        DP_OP_424J2_126_3477_n2898), .CI(DP_OP_424J2_126_3477_n2377), .CO(
        DP_OP_424J2_126_3477_n1719), .S(DP_OP_424J2_126_3477_n1720) );
  FADDX1_HVT DP_OP_424J2_126_3477_U956 ( .A(DP_OP_424J2_126_3477_n2248), .B(
        DP_OP_424J2_126_3477_n1977), .CI(DP_OP_424J2_126_3477_n2905), .CO(
        DP_OP_424J2_126_3477_n1717), .S(DP_OP_424J2_126_3477_n1718) );
  FADDX1_HVT DP_OP_424J2_126_3477_U955 ( .A(DP_OP_424J2_126_3477_n2160), .B(
        DP_OP_424J2_126_3477_n2722), .CI(DP_OP_424J2_126_3477_n2817), .CO(
        DP_OP_424J2_126_3477_n1715), .S(DP_OP_424J2_126_3477_n1716) );
  FADDX1_HVT DP_OP_424J2_126_3477_U954 ( .A(DP_OP_424J2_126_3477_n2021), .B(
        DP_OP_424J2_126_3477_n1771), .CI(DP_OP_424J2_126_3477_n1748), .CO(
        DP_OP_424J2_126_3477_n1713), .S(DP_OP_424J2_126_3477_n1714) );
  FADDX1_HVT DP_OP_424J2_126_3477_U953 ( .A(DP_OP_424J2_126_3477_n1759), .B(
        DP_OP_424J2_126_3477_n1769), .CI(DP_OP_424J2_126_3477_n1767), .CO(
        DP_OP_424J2_126_3477_n1711), .S(DP_OP_424J2_126_3477_n1712) );
  FADDX1_HVT DP_OP_424J2_126_3477_U952 ( .A(DP_OP_424J2_126_3477_n1763), .B(
        DP_OP_424J2_126_3477_n1765), .CI(DP_OP_424J2_126_3477_n1761), .CO(
        DP_OP_424J2_126_3477_n1709), .S(DP_OP_424J2_126_3477_n1710) );
  FADDX1_HVT DP_OP_424J2_126_3477_U951 ( .A(DP_OP_424J2_126_3477_n1757), .B(
        DP_OP_424J2_126_3477_n1755), .CI(DP_OP_424J2_126_3477_n1738), .CO(
        DP_OP_424J2_126_3477_n1707), .S(DP_OP_424J2_126_3477_n1708) );
  FADDX1_HVT DP_OP_424J2_126_3477_U950 ( .A(DP_OP_424J2_126_3477_n1736), .B(
        DP_OP_424J2_126_3477_n1742), .CI(DP_OP_424J2_126_3477_n1730), .CO(
        DP_OP_424J2_126_3477_n1705), .S(DP_OP_424J2_126_3477_n1706) );
  FADDX1_HVT DP_OP_424J2_126_3477_U949 ( .A(DP_OP_424J2_126_3477_n1740), .B(
        DP_OP_424J2_126_3477_n1746), .CI(DP_OP_424J2_126_3477_n1734), .CO(
        DP_OP_424J2_126_3477_n1703), .S(DP_OP_424J2_126_3477_n1704) );
  FADDX1_HVT DP_OP_424J2_126_3477_U948 ( .A(DP_OP_424J2_126_3477_n1732), .B(
        DP_OP_424J2_126_3477_n1744), .CI(DP_OP_424J2_126_3477_n1728), .CO(
        DP_OP_424J2_126_3477_n1701), .S(DP_OP_424J2_126_3477_n1702) );
  FADDX1_HVT DP_OP_424J2_126_3477_U947 ( .A(DP_OP_424J2_126_3477_n1726), .B(
        DP_OP_424J2_126_3477_n1718), .CI(DP_OP_424J2_126_3477_n1716), .CO(
        DP_OP_424J2_126_3477_n1699), .S(DP_OP_424J2_126_3477_n1700) );
  FADDX1_HVT DP_OP_424J2_126_3477_U946 ( .A(DP_OP_424J2_126_3477_n1722), .B(
        DP_OP_424J2_126_3477_n1724), .CI(DP_OP_424J2_126_3477_n1720), .CO(
        DP_OP_424J2_126_3477_n1697), .S(DP_OP_424J2_126_3477_n1698) );
  FADDX1_HVT DP_OP_424J2_126_3477_U945 ( .A(DP_OP_424J2_126_3477_n1714), .B(
        DP_OP_424J2_126_3477_n1753), .CI(DP_OP_424J2_126_3477_n1751), .CO(
        DP_OP_424J2_126_3477_n1695), .S(DP_OP_424J2_126_3477_n1696) );
  FADDX1_HVT DP_OP_424J2_126_3477_U944 ( .A(DP_OP_424J2_126_3477_n1712), .B(
        DP_OP_424J2_126_3477_n1710), .CI(DP_OP_424J2_126_3477_n1749), .CO(
        DP_OP_424J2_126_3477_n1693), .S(DP_OP_424J2_126_3477_n1694) );
  FADDX1_HVT DP_OP_424J2_126_3477_U943 ( .A(DP_OP_424J2_126_3477_n1708), .B(
        DP_OP_424J2_126_3477_n1706), .CI(DP_OP_424J2_126_3477_n1704), .CO(
        DP_OP_424J2_126_3477_n1691), .S(DP_OP_424J2_126_3477_n1692) );
  FADDX1_HVT DP_OP_424J2_126_3477_U942 ( .A(DP_OP_424J2_126_3477_n1702), .B(
        DP_OP_424J2_126_3477_n1700), .CI(DP_OP_424J2_126_3477_n1698), .CO(
        DP_OP_424J2_126_3477_n1689), .S(DP_OP_424J2_126_3477_n1690) );
  FADDX1_HVT DP_OP_424J2_126_3477_U941 ( .A(DP_OP_424J2_126_3477_n1696), .B(
        DP_OP_424J2_126_3477_n1694), .CI(DP_OP_424J2_126_3477_n1692), .CO(
        DP_OP_424J2_126_3477_n1687), .S(DP_OP_424J2_126_3477_n1688) );
  HADDX1_HVT DP_OP_424J2_126_3477_U940 ( .A0(DP_OP_424J2_126_3477_n2464), .B0(
        DP_OP_424J2_126_3477_n2152), .C1(DP_OP_424J2_126_3477_n1685), .SO(
        DP_OP_424J2_126_3477_n1686) );
  FADDX1_HVT DP_OP_424J2_126_3477_U939 ( .A(DP_OP_424J2_126_3477_n2846), .B(
        DP_OP_424J2_126_3477_n2413), .CI(DP_OP_424J2_126_3477_n2071), .CO(
        DP_OP_424J2_126_3477_n1683), .S(DP_OP_424J2_126_3477_n1684) );
  FADDX1_HVT DP_OP_424J2_126_3477_U938 ( .A(DP_OP_424J2_126_3477_n2890), .B(
        DP_OP_424J2_126_3477_n2538), .CI(DP_OP_424J2_126_3477_n2277), .CO(
        DP_OP_424J2_126_3477_n1681), .S(DP_OP_424J2_126_3477_n1682) );
  FADDX1_HVT DP_OP_424J2_126_3477_U937 ( .A(DP_OP_424J2_126_3477_n2596), .B(
        DP_OP_424J2_126_3477_n2728), .CI(DP_OP_424J2_126_3477_n2291), .CO(
        DP_OP_424J2_126_3477_n1679), .S(DP_OP_424J2_126_3477_n1680) );
  FADDX1_HVT DP_OP_424J2_126_3477_U936 ( .A(DP_OP_424J2_126_3477_n2640), .B(
        DP_OP_424J2_126_3477_n1969), .CI(DP_OP_424J2_126_3477_n2145), .CO(
        DP_OP_424J2_126_3477_n1677), .S(DP_OP_424J2_126_3477_n1678) );
  FADDX1_HVT DP_OP_424J2_126_3477_U935 ( .A(DP_OP_424J2_126_3477_n2420), .B(
        DP_OP_424J2_126_3477_n1786), .CI(DP_OP_424J2_126_3477_n2508), .CO(
        DP_OP_424J2_126_3477_n1675), .S(DP_OP_424J2_126_3477_n1676) );
  FADDX1_HVT DP_OP_424J2_126_3477_U934 ( .A(DP_OP_424J2_126_3477_n2203), .B(
        DP_OP_424J2_126_3477_n2633), .CI(DP_OP_424J2_126_3477_n2860), .CO(
        DP_OP_424J2_126_3477_n1673), .S(DP_OP_424J2_126_3477_n1674) );
  FADDX1_HVT DP_OP_424J2_126_3477_U933 ( .A(DP_OP_424J2_126_3477_n1851), .B(
        DP_OP_424J2_126_3477_n2758), .CI(DP_OP_424J2_126_3477_n2772), .CO(
        DP_OP_424J2_126_3477_n1671), .S(DP_OP_424J2_126_3477_n1672) );
  FADDX1_HVT DP_OP_424J2_126_3477_U932 ( .A(DP_OP_424J2_126_3477_n2335), .B(
        DP_OP_424J2_126_3477_n2328), .CI(DP_OP_424J2_126_3477_n2101), .CO(
        DP_OP_424J2_126_3477_n1669), .S(DP_OP_424J2_126_3477_n1670) );
  FADDX1_HVT DP_OP_424J2_126_3477_U931 ( .A(DP_OP_424J2_126_3477_n2115), .B(
        DP_OP_424J2_126_3477_n1983), .CI(DP_OP_424J2_126_3477_n1895), .CO(
        DP_OP_424J2_126_3477_n1667), .S(DP_OP_424J2_126_3477_n1668) );
  FADDX1_HVT DP_OP_424J2_126_3477_U930 ( .A(DP_OP_424J2_126_3477_n2552), .B(
        DP_OP_424J2_126_3477_n2684), .CI(DP_OP_424J2_126_3477_n2450), .CO(
        DP_OP_424J2_126_3477_n1665), .S(DP_OP_424J2_126_3477_n1666) );
  FADDX1_HVT DP_OP_424J2_126_3477_U929 ( .A(DP_OP_424J2_126_3477_n2501), .B(
        DP_OP_424J2_126_3477_n2589), .CI(DP_OP_424J2_126_3477_n2233), .CO(
        DP_OP_424J2_126_3477_n1663), .S(DP_OP_424J2_126_3477_n1664) );
  FADDX1_HVT DP_OP_424J2_126_3477_U928 ( .A(DP_OP_424J2_126_3477_n2064), .B(
        DP_OP_424J2_126_3477_n1844), .CI(DP_OP_424J2_126_3477_n2582), .CO(
        DP_OP_424J2_126_3477_n1661), .S(DP_OP_424J2_126_3477_n1662) );
  FADDX1_HVT DP_OP_424J2_126_3477_U927 ( .A(DP_OP_424J2_126_3477_n2027), .B(
        DP_OP_424J2_126_3477_n1939), .CI(DP_OP_424J2_126_3477_n2714), .CO(
        DP_OP_424J2_126_3477_n1659), .S(DP_OP_424J2_126_3477_n1660) );
  FADDX1_HVT DP_OP_424J2_126_3477_U926 ( .A(DP_OP_424J2_126_3477_n2545), .B(
        DP_OP_424J2_126_3477_n2765), .CI(DP_OP_424J2_126_3477_n2013), .CO(
        DP_OP_424J2_126_3477_n1657), .S(DP_OP_424J2_126_3477_n1658) );
  FADDX1_HVT DP_OP_424J2_126_3477_U925 ( .A(DP_OP_424J2_126_3477_n2853), .B(
        DP_OP_424J2_126_3477_n2457), .CI(DP_OP_424J2_126_3477_n2240), .CO(
        DP_OP_424J2_126_3477_n1655), .S(DP_OP_424J2_126_3477_n1656) );
  FADDX1_HVT DP_OP_424J2_126_3477_U924 ( .A(DP_OP_424J2_126_3477_n2108), .B(
        DP_OP_424J2_126_3477_n2284), .CI(DP_OP_424J2_126_3477_n2369), .CO(
        DP_OP_424J2_126_3477_n1653), .S(DP_OP_424J2_126_3477_n1654) );
  FADDX1_HVT DP_OP_424J2_126_3477_U923 ( .A(DP_OP_424J2_126_3477_n1888), .B(
        DP_OP_424J2_126_3477_n2809), .CI(DP_OP_424J2_126_3477_n2196), .CO(
        DP_OP_424J2_126_3477_n1651), .S(DP_OP_424J2_126_3477_n1652) );
  FADDX1_HVT DP_OP_424J2_126_3477_U922 ( .A(DP_OP_424J2_126_3477_n2494), .B(
        DP_OP_424J2_126_3477_n2670), .CI(DP_OP_424J2_126_3477_n1932), .CO(
        DP_OP_424J2_126_3477_n1649), .S(DP_OP_424J2_126_3477_n1650) );
  FADDX1_HVT DP_OP_424J2_126_3477_U921 ( .A(DP_OP_424J2_126_3477_n2362), .B(
        DP_OP_424J2_126_3477_n2897), .CI(DP_OP_424J2_126_3477_n2904), .CO(
        DP_OP_424J2_126_3477_n1647), .S(DP_OP_424J2_126_3477_n1648) );
  FADDX1_HVT DP_OP_424J2_126_3477_U920 ( .A(DP_OP_424J2_126_3477_n2677), .B(
        DP_OP_424J2_126_3477_n2247), .CI(DP_OP_424J2_126_3477_n2376), .CO(
        DP_OP_424J2_126_3477_n1645), .S(DP_OP_424J2_126_3477_n1646) );
  FADDX1_HVT DP_OP_424J2_126_3477_U919 ( .A(DP_OP_424J2_126_3477_n2057), .B(
        DP_OP_424J2_126_3477_n2321), .CI(DP_OP_424J2_126_3477_n2721), .CO(
        DP_OP_424J2_126_3477_n1643), .S(DP_OP_424J2_126_3477_n1644) );
  FADDX1_HVT DP_OP_424J2_126_3477_U918 ( .A(DP_OP_424J2_126_3477_n2802), .B(
        DP_OP_424J2_126_3477_n2159), .CI(DP_OP_424J2_126_3477_n2816), .CO(
        DP_OP_424J2_126_3477_n1641), .S(DP_OP_424J2_126_3477_n1642) );
  FADDX1_HVT DP_OP_424J2_126_3477_U917 ( .A(DP_OP_424J2_126_3477_n2626), .B(
        DP_OP_424J2_126_3477_n2406), .CI(DP_OP_424J2_126_3477_n2020), .CO(
        DP_OP_424J2_126_3477_n1639), .S(DP_OP_424J2_126_3477_n1640) );
  FADDX1_HVT DP_OP_424J2_126_3477_U916 ( .A(DP_OP_424J2_126_3477_n1976), .B(
        DP_OP_424J2_126_3477_n2189), .CI(DP_OP_424J2_126_3477_n1925), .CO(
        DP_OP_424J2_126_3477_n1637), .S(DP_OP_424J2_126_3477_n1638) );
  FADDX1_HVT DP_OP_424J2_126_3477_U915 ( .A(DP_OP_424J2_126_3477_n1881), .B(
        DP_OP_424J2_126_3477_n1837), .CI(DP_OP_424J2_126_3477_n1747), .CO(
        DP_OP_424J2_126_3477_n1635), .S(DP_OP_424J2_126_3477_n1636) );
  FADDX1_HVT DP_OP_424J2_126_3477_U914 ( .A(DP_OP_424J2_126_3477_n1686), .B(
        DP_OP_424J2_126_3477_n1745), .CI(DP_OP_424J2_126_3477_n1729), .CO(
        DP_OP_424J2_126_3477_n1633), .S(DP_OP_424J2_126_3477_n1634) );
  FADDX1_HVT DP_OP_424J2_126_3477_U913 ( .A(DP_OP_424J2_126_3477_n1743), .B(
        DP_OP_424J2_126_3477_n1731), .CI(DP_OP_424J2_126_3477_n1741), .CO(
        DP_OP_424J2_126_3477_n1631), .S(DP_OP_424J2_126_3477_n1632) );
  FADDX1_HVT DP_OP_424J2_126_3477_U912 ( .A(DP_OP_424J2_126_3477_n1733), .B(
        DP_OP_424J2_126_3477_n1735), .CI(DP_OP_424J2_126_3477_n1737), .CO(
        DP_OP_424J2_126_3477_n1629), .S(DP_OP_424J2_126_3477_n1630) );
  FADDX1_HVT DP_OP_424J2_126_3477_U911 ( .A(DP_OP_424J2_126_3477_n1739), .B(
        DP_OP_424J2_126_3477_n1727), .CI(DP_OP_424J2_126_3477_n1725), .CO(
        DP_OP_424J2_126_3477_n1627), .S(DP_OP_424J2_126_3477_n1628) );
  FADDX1_HVT DP_OP_424J2_126_3477_U910 ( .A(DP_OP_424J2_126_3477_n1723), .B(
        DP_OP_424J2_126_3477_n1717), .CI(DP_OP_424J2_126_3477_n1715), .CO(
        DP_OP_424J2_126_3477_n1625), .S(DP_OP_424J2_126_3477_n1626) );
  FADDX1_HVT DP_OP_424J2_126_3477_U909 ( .A(DP_OP_424J2_126_3477_n1721), .B(
        DP_OP_424J2_126_3477_n1719), .CI(DP_OP_424J2_126_3477_n1668), .CO(
        DP_OP_424J2_126_3477_n1623), .S(DP_OP_424J2_126_3477_n1624) );
  FADDX1_HVT DP_OP_424J2_126_3477_U908 ( .A(DP_OP_424J2_126_3477_n1678), .B(
        DP_OP_424J2_126_3477_n1664), .CI(DP_OP_424J2_126_3477_n1660), .CO(
        DP_OP_424J2_126_3477_n1621), .S(DP_OP_424J2_126_3477_n1622) );
  FADDX1_HVT DP_OP_424J2_126_3477_U907 ( .A(DP_OP_424J2_126_3477_n1676), .B(
        DP_OP_424J2_126_3477_n1670), .CI(DP_OP_424J2_126_3477_n1662), .CO(
        DP_OP_424J2_126_3477_n1619), .S(DP_OP_424J2_126_3477_n1620) );
  FADDX1_HVT DP_OP_424J2_126_3477_U906 ( .A(DP_OP_424J2_126_3477_n1684), .B(
        DP_OP_424J2_126_3477_n1666), .CI(DP_OP_424J2_126_3477_n1672), .CO(
        DP_OP_424J2_126_3477_n1617), .S(DP_OP_424J2_126_3477_n1618) );
  FADDX1_HVT DP_OP_424J2_126_3477_U905 ( .A(DP_OP_424J2_126_3477_n1682), .B(
        DP_OP_424J2_126_3477_n1674), .CI(DP_OP_424J2_126_3477_n1680), .CO(
        DP_OP_424J2_126_3477_n1615), .S(DP_OP_424J2_126_3477_n1616) );
  FADDX1_HVT DP_OP_424J2_126_3477_U904 ( .A(DP_OP_424J2_126_3477_n1658), .B(
        DP_OP_424J2_126_3477_n1644), .CI(DP_OP_424J2_126_3477_n1713), .CO(
        DP_OP_424J2_126_3477_n1613), .S(DP_OP_424J2_126_3477_n1614) );
  FADDX1_HVT DP_OP_424J2_126_3477_U903 ( .A(DP_OP_424J2_126_3477_n1656), .B(
        DP_OP_424J2_126_3477_n1646), .CI(DP_OP_424J2_126_3477_n1642), .CO(
        DP_OP_424J2_126_3477_n1611), .S(DP_OP_424J2_126_3477_n1612) );
  FADDX1_HVT DP_OP_424J2_126_3477_U902 ( .A(DP_OP_424J2_126_3477_n1652), .B(
        DP_OP_424J2_126_3477_n1648), .CI(DP_OP_424J2_126_3477_n1640), .CO(
        DP_OP_424J2_126_3477_n1609), .S(DP_OP_424J2_126_3477_n1610) );
  FADDX1_HVT DP_OP_424J2_126_3477_U901 ( .A(DP_OP_424J2_126_3477_n1654), .B(
        DP_OP_424J2_126_3477_n1650), .CI(DP_OP_424J2_126_3477_n1638), .CO(
        DP_OP_424J2_126_3477_n1607), .S(DP_OP_424J2_126_3477_n1608) );
  FADDX1_HVT DP_OP_424J2_126_3477_U900 ( .A(DP_OP_424J2_126_3477_n1636), .B(
        DP_OP_424J2_126_3477_n1711), .CI(DP_OP_424J2_126_3477_n1709), .CO(
        DP_OP_424J2_126_3477_n1605), .S(DP_OP_424J2_126_3477_n1606) );
  FADDX1_HVT DP_OP_424J2_126_3477_U899 ( .A(DP_OP_424J2_126_3477_n1707), .B(
        DP_OP_424J2_126_3477_n1634), .CI(DP_OP_424J2_126_3477_n1632), .CO(
        DP_OP_424J2_126_3477_n1603), .S(DP_OP_424J2_126_3477_n1604) );
  FADDX1_HVT DP_OP_424J2_126_3477_U898 ( .A(DP_OP_424J2_126_3477_n1705), .B(
        DP_OP_424J2_126_3477_n1630), .CI(DP_OP_424J2_126_3477_n1628), .CO(
        DP_OP_424J2_126_3477_n1601), .S(DP_OP_424J2_126_3477_n1602) );
  FADDX1_HVT DP_OP_424J2_126_3477_U897 ( .A(DP_OP_424J2_126_3477_n1703), .B(
        DP_OP_424J2_126_3477_n1701), .CI(DP_OP_424J2_126_3477_n1699), .CO(
        DP_OP_424J2_126_3477_n1599), .S(DP_OP_424J2_126_3477_n1600) );
  FADDX1_HVT DP_OP_424J2_126_3477_U896 ( .A(DP_OP_424J2_126_3477_n1697), .B(
        DP_OP_424J2_126_3477_n1626), .CI(DP_OP_424J2_126_3477_n1624), .CO(
        DP_OP_424J2_126_3477_n1597), .S(DP_OP_424J2_126_3477_n1598) );
  FADDX1_HVT DP_OP_424J2_126_3477_U895 ( .A(DP_OP_424J2_126_3477_n1622), .B(
        DP_OP_424J2_126_3477_n1616), .CI(DP_OP_424J2_126_3477_n1618), .CO(
        DP_OP_424J2_126_3477_n1595), .S(DP_OP_424J2_126_3477_n1596) );
  FADDX1_HVT DP_OP_424J2_126_3477_U894 ( .A(DP_OP_424J2_126_3477_n1620), .B(
        DP_OP_424J2_126_3477_n1614), .CI(DP_OP_424J2_126_3477_n1612), .CO(
        DP_OP_424J2_126_3477_n1593), .S(DP_OP_424J2_126_3477_n1594) );
  FADDX1_HVT DP_OP_424J2_126_3477_U893 ( .A(DP_OP_424J2_126_3477_n1608), .B(
        DP_OP_424J2_126_3477_n1610), .CI(DP_OP_424J2_126_3477_n1695), .CO(
        DP_OP_424J2_126_3477_n1591), .S(DP_OP_424J2_126_3477_n1592) );
  FADDX1_HVT DP_OP_424J2_126_3477_U892 ( .A(DP_OP_424J2_126_3477_n1606), .B(
        DP_OP_424J2_126_3477_n1693), .CI(DP_OP_424J2_126_3477_n1604), .CO(
        DP_OP_424J2_126_3477_n1589), .S(DP_OP_424J2_126_3477_n1590) );
  FADDX1_HVT DP_OP_424J2_126_3477_U891 ( .A(DP_OP_424J2_126_3477_n1691), .B(
        DP_OP_424J2_126_3477_n1602), .CI(DP_OP_424J2_126_3477_n1600), .CO(
        DP_OP_424J2_126_3477_n1587), .S(DP_OP_424J2_126_3477_n1588) );
  FADDX1_HVT DP_OP_424J2_126_3477_U890 ( .A(DP_OP_424J2_126_3477_n1689), .B(
        DP_OP_424J2_126_3477_n1598), .CI(DP_OP_424J2_126_3477_n1596), .CO(
        DP_OP_424J2_126_3477_n1585), .S(DP_OP_424J2_126_3477_n1586) );
  FADDX1_HVT DP_OP_424J2_126_3477_U889 ( .A(DP_OP_424J2_126_3477_n1594), .B(
        DP_OP_424J2_126_3477_n1592), .CI(DP_OP_424J2_126_3477_n1590), .CO(
        DP_OP_424J2_126_3477_n1583), .S(DP_OP_424J2_126_3477_n1584) );
  FADDX1_HVT DP_OP_424J2_126_3477_U888 ( .A(DP_OP_424J2_126_3477_n1687), .B(
        DP_OP_424J2_126_3477_n1588), .CI(DP_OP_424J2_126_3477_n1586), .CO(
        DP_OP_424J2_126_3477_n1581), .S(DP_OP_424J2_126_3477_n1582) );
  FADDX1_HVT DP_OP_424J2_126_3477_U886 ( .A(DP_OP_424J2_126_3477_n2005), .B(
        DP_OP_424J2_126_3477_n1829), .CI(DP_OP_424J2_126_3477_n2398), .CO(
        DP_OP_424J2_126_3477_n1577), .S(DP_OP_424J2_126_3477_n1578) );
  FADDX1_HVT DP_OP_424J2_126_3477_U885 ( .A(DP_OP_424J2_126_3477_n2706), .B(
        DP_OP_424J2_126_3477_n1917), .CI(DP_OP_424J2_126_3477_n1961), .CO(
        DP_OP_424J2_126_3477_n1575), .S(DP_OP_424J2_126_3477_n1576) );
  FADDX1_HVT DP_OP_424J2_126_3477_U884 ( .A(DP_OP_424J2_126_3477_n2618), .B(
        DP_OP_424J2_126_3477_n2442), .CI(DP_OP_424J2_126_3477_n2750), .CO(
        DP_OP_424J2_126_3477_n1573), .S(DP_OP_424J2_126_3477_n1574) );
  FADDX1_HVT DP_OP_424J2_126_3477_U883 ( .A(DP_OP_424J2_126_3477_n1873), .B(
        DP_OP_424J2_126_3477_n2574), .CI(DP_OP_424J2_126_3477_n2530), .CO(
        DP_OP_424J2_126_3477_n1571), .S(DP_OP_424J2_126_3477_n1572) );
  FADDX1_HVT DP_OP_424J2_126_3477_U882 ( .A(DP_OP_424J2_126_3477_n2662), .B(
        DP_OP_424J2_126_3477_n2049), .CI(DP_OP_424J2_126_3477_n2486), .CO(
        DP_OP_424J2_126_3477_n1569), .S(DP_OP_424J2_126_3477_n1570) );
  FADDX1_HVT DP_OP_424J2_126_3477_U881 ( .A(DP_OP_424J2_126_3477_n2093), .B(
        DP_OP_424J2_126_3477_n2882), .CI(DP_OP_424J2_126_3477_n2181), .CO(
        DP_OP_424J2_126_3477_n1567), .S(DP_OP_424J2_126_3477_n1568) );
  FADDX1_HVT DP_OP_424J2_126_3477_U880 ( .A(DP_OP_424J2_126_3477_n2838), .B(
        DP_OP_424J2_126_3477_n2794), .CI(DP_OP_424J2_126_3477_n2269), .CO(
        DP_OP_424J2_126_3477_n1565), .S(DP_OP_424J2_126_3477_n1566) );
  FADDX1_HVT DP_OP_424J2_126_3477_U879 ( .A(DP_OP_424J2_126_3477_n2137), .B(
        DP_OP_424J2_126_3477_n2313), .CI(DP_OP_424J2_126_3477_n1580), .CO(
        DP_OP_424J2_126_3477_n1563), .S(DP_OP_424J2_126_3477_n1564) );
  FADDX1_HVT DP_OP_424J2_126_3477_U878 ( .A(DP_OP_424J2_126_3477_n2225), .B(
        DP_OP_424J2_126_3477_n2151), .CI(DP_OP_424J2_126_3477_n2276), .CO(
        DP_OP_424J2_126_3477_n1561), .S(DP_OP_424J2_126_3477_n1562) );
  FADDX1_HVT DP_OP_424J2_126_3477_U877 ( .A(DP_OP_424J2_126_3477_n2114), .B(
        DP_OP_424J2_126_3477_n2412), .CI(DP_OP_424J2_126_3477_n2144), .CO(
        DP_OP_424J2_126_3477_n1559), .S(DP_OP_424J2_126_3477_n1560) );
  FADDX1_HVT DP_OP_424J2_126_3477_U876 ( .A(DP_OP_424J2_126_3477_n2334), .B(
        DP_OP_424J2_126_3477_n2727), .CI(DP_OP_424J2_126_3477_n2070), .CO(
        DP_OP_424J2_126_3477_n1557), .S(DP_OP_424J2_126_3477_n1558) );
  FADDX1_HVT DP_OP_424J2_126_3477_U875 ( .A(DP_OP_424J2_126_3477_n2595), .B(
        DP_OP_424J2_126_3477_n1968), .CI(DP_OP_424J2_126_3477_n2290), .CO(
        DP_OP_424J2_126_3477_n1555), .S(DP_OP_424J2_126_3477_n1556) );
  FADDX1_HVT DP_OP_424J2_126_3477_U874 ( .A(DP_OP_424J2_126_3477_n2202), .B(
        DP_OP_424J2_126_3477_n2537), .CI(DP_OP_424J2_126_3477_n2507), .CO(
        DP_OP_424J2_126_3477_n1553), .S(DP_OP_424J2_126_3477_n1554) );
  FADDX1_HVT DP_OP_424J2_126_3477_U873 ( .A(DP_OP_424J2_126_3477_n2463), .B(
        DP_OP_424J2_126_3477_n1785), .CI(DP_OP_424J2_126_3477_n2100), .CO(
        DP_OP_424J2_126_3477_n1551), .S(DP_OP_424J2_126_3477_n1552) );
  FADDX1_HVT DP_OP_424J2_126_3477_U872 ( .A(DP_OP_424J2_126_3477_n2845), .B(
        DP_OP_424J2_126_3477_n2588), .CI(DP_OP_424J2_126_3477_n2771), .CO(
        DP_OP_424J2_126_3477_n1549), .S(DP_OP_424J2_126_3477_n1550) );
  FADDX1_HVT DP_OP_424J2_126_3477_U871 ( .A(DP_OP_424J2_126_3477_n2889), .B(
        DP_OP_424J2_126_3477_n1843), .CI(DP_OP_424J2_126_3477_n2232), .CO(
        DP_OP_424J2_126_3477_n1547), .S(DP_OP_424J2_126_3477_n1548) );
  FADDX1_HVT DP_OP_424J2_126_3477_U870 ( .A(DP_OP_424J2_126_3477_n2419), .B(
        DP_OP_424J2_126_3477_n2327), .CI(DP_OP_424J2_126_3477_n2859), .CO(
        DP_OP_424J2_126_3477_n1545), .S(DP_OP_424J2_126_3477_n1546) );
  FADDX1_HVT DP_OP_424J2_126_3477_U869 ( .A(DP_OP_424J2_126_3477_n2639), .B(
        DP_OP_424J2_126_3477_n2500), .CI(DP_OP_424J2_126_3477_n2449), .CO(
        DP_OP_424J2_126_3477_n1543), .S(DP_OP_424J2_126_3477_n1544) );
  FADDX1_HVT DP_OP_424J2_126_3477_U868 ( .A(DP_OP_424J2_126_3477_n2551), .B(
        DP_OP_424J2_126_3477_n2757), .CI(DP_OP_424J2_126_3477_n1894), .CO(
        DP_OP_424J2_126_3477_n1541), .S(DP_OP_424J2_126_3477_n1542) );
  FADDX1_HVT DP_OP_424J2_126_3477_U867 ( .A(DP_OP_424J2_126_3477_n1850), .B(
        DP_OP_424J2_126_3477_n2683), .CI(DP_OP_424J2_126_3477_n2581), .CO(
        DP_OP_424J2_126_3477_n1539), .S(DP_OP_424J2_126_3477_n1540) );
  FADDX1_HVT DP_OP_424J2_126_3477_U866 ( .A(DP_OP_424J2_126_3477_n2632), .B(
        DP_OP_424J2_126_3477_n2026), .CI(DP_OP_424J2_126_3477_n1982), .CO(
        DP_OP_424J2_126_3477_n1537), .S(DP_OP_424J2_126_3477_n1538) );
  FADDX1_HVT DP_OP_424J2_126_3477_U865 ( .A(DP_OP_424J2_126_3477_n2063), .B(
        DP_OP_424J2_126_3477_n1938), .CI(DP_OP_424J2_126_3477_n2544), .CO(
        DP_OP_424J2_126_3477_n1535), .S(DP_OP_424J2_126_3477_n1536) );
  FADDX1_HVT DP_OP_424J2_126_3477_U864 ( .A(DP_OP_424J2_126_3477_n2713), .B(
        DP_OP_424J2_126_3477_n2764), .CI(DP_OP_424J2_126_3477_n2368), .CO(
        DP_OP_424J2_126_3477_n1533), .S(DP_OP_424J2_126_3477_n1534) );
  FADDX1_HVT DP_OP_424J2_126_3477_U863 ( .A(DP_OP_424J2_126_3477_n2852), .B(
        DP_OP_424J2_126_3477_n2456), .CI(DP_OP_424J2_126_3477_n2239), .CO(
        DP_OP_424J2_126_3477_n1531), .S(DP_OP_424J2_126_3477_n1532) );
  FADDX1_HVT DP_OP_424J2_126_3477_U862 ( .A(DP_OP_424J2_126_3477_n1887), .B(
        DP_OP_424J2_126_3477_n2283), .CI(DP_OP_424J2_126_3477_n2195), .CO(
        DP_OP_424J2_126_3477_n1529), .S(DP_OP_424J2_126_3477_n1530) );
  FADDX1_HVT DP_OP_424J2_126_3477_U861 ( .A(DP_OP_424J2_126_3477_n2107), .B(
        DP_OP_424J2_126_3477_n2808), .CI(DP_OP_424J2_126_3477_n2012), .CO(
        DP_OP_424J2_126_3477_n1527), .S(DP_OP_424J2_126_3477_n1528) );
  FADDX1_HVT DP_OP_424J2_126_3477_U860 ( .A(DP_OP_424J2_126_3477_n2493), .B(
        DP_OP_424J2_126_3477_n2669), .CI(DP_OP_424J2_126_3477_n1931), .CO(
        DP_OP_424J2_126_3477_n1525), .S(DP_OP_424J2_126_3477_n1526) );
  FADDX1_HVT DP_OP_424J2_126_3477_U859 ( .A(DP_OP_424J2_126_3477_n2361), .B(
        DP_OP_424J2_126_3477_n2896), .CI(DP_OP_424J2_126_3477_n2375), .CO(
        DP_OP_424J2_126_3477_n1523), .S(DP_OP_424J2_126_3477_n1524) );
  FADDX1_HVT DP_OP_424J2_126_3477_U858 ( .A(DP_OP_424J2_126_3477_n2676), .B(
        DP_OP_424J2_126_3477_n2246), .CI(DP_OP_424J2_126_3477_n2720), .CO(
        DP_OP_424J2_126_3477_n1521), .S(DP_OP_424J2_126_3477_n1522) );
  FADDX1_HVT DP_OP_424J2_126_3477_U857 ( .A(DP_OP_424J2_126_3477_n2320), .B(
        DP_OP_424J2_126_3477_n2056), .CI(DP_OP_424J2_126_3477_n2903), .CO(
        DP_OP_424J2_126_3477_n1519), .S(DP_OP_424J2_126_3477_n1520) );
  FADDX1_HVT DP_OP_424J2_126_3477_U856 ( .A(DP_OP_424J2_126_3477_n2625), .B(
        DP_OP_424J2_126_3477_n2019), .CI(DP_OP_424J2_126_3477_n2815), .CO(
        DP_OP_424J2_126_3477_n1517), .S(DP_OP_424J2_126_3477_n1518) );
  FADDX1_HVT DP_OP_424J2_126_3477_U855 ( .A(DP_OP_424J2_126_3477_n2801), .B(
        DP_OP_424J2_126_3477_n2158), .CI(DP_OP_424J2_126_3477_n2405), .CO(
        DP_OP_424J2_126_3477_n1515), .S(DP_OP_424J2_126_3477_n1516) );
  FADDX1_HVT DP_OP_424J2_126_3477_U854 ( .A(DP_OP_424J2_126_3477_n1975), .B(
        DP_OP_424J2_126_3477_n1924), .CI(DP_OP_424J2_126_3477_n2188), .CO(
        DP_OP_424J2_126_3477_n1513), .S(DP_OP_424J2_126_3477_n1514) );
  FADDX1_HVT DP_OP_424J2_126_3477_U853 ( .A(DP_OP_424J2_126_3477_n1880), .B(
        DP_OP_424J2_126_3477_n1836), .CI(DP_OP_424J2_126_3477_n1685), .CO(
        DP_OP_424J2_126_3477_n1511), .S(DP_OP_424J2_126_3477_n1512) );
  FADDX1_HVT DP_OP_424J2_126_3477_U852 ( .A(DP_OP_424J2_126_3477_n1683), .B(
        DP_OP_424J2_126_3477_n1661), .CI(DP_OP_424J2_126_3477_n1659), .CO(
        DP_OP_424J2_126_3477_n1509), .S(DP_OP_424J2_126_3477_n1510) );
  FADDX1_HVT DP_OP_424J2_126_3477_U851 ( .A(DP_OP_424J2_126_3477_n1673), .B(
        DP_OP_424J2_126_3477_n1665), .CI(DP_OP_424J2_126_3477_n1663), .CO(
        DP_OP_424J2_126_3477_n1507), .S(DP_OP_424J2_126_3477_n1508) );
  FADDX1_HVT DP_OP_424J2_126_3477_U850 ( .A(DP_OP_424J2_126_3477_n1681), .B(
        DP_OP_424J2_126_3477_n1667), .CI(DP_OP_424J2_126_3477_n1669), .CO(
        DP_OP_424J2_126_3477_n1505), .S(DP_OP_424J2_126_3477_n1506) );
  FADDX1_HVT DP_OP_424J2_126_3477_U849 ( .A(DP_OP_424J2_126_3477_n1679), .B(
        DP_OP_424J2_126_3477_n1671), .CI(DP_OP_424J2_126_3477_n1675), .CO(
        DP_OP_424J2_126_3477_n1503), .S(DP_OP_424J2_126_3477_n1504) );
  FADDX1_HVT DP_OP_424J2_126_3477_U848 ( .A(DP_OP_424J2_126_3477_n1677), .B(
        DP_OP_424J2_126_3477_n1657), .CI(DP_OP_424J2_126_3477_n1655), .CO(
        DP_OP_424J2_126_3477_n1501), .S(DP_OP_424J2_126_3477_n1502) );
  FADDX1_HVT DP_OP_424J2_126_3477_U847 ( .A(DP_OP_424J2_126_3477_n1653), .B(
        DP_OP_424J2_126_3477_n1574), .CI(DP_OP_424J2_126_3477_n1637), .CO(
        DP_OP_424J2_126_3477_n1499), .S(DP_OP_424J2_126_3477_n1500) );
  FADDX1_HVT DP_OP_424J2_126_3477_U846 ( .A(DP_OP_424J2_126_3477_n1649), .B(
        DP_OP_424J2_126_3477_n1572), .CI(DP_OP_424J2_126_3477_n1641), .CO(
        DP_OP_424J2_126_3477_n1497), .S(DP_OP_424J2_126_3477_n1498) );
  FADDX1_HVT DP_OP_424J2_126_3477_U845 ( .A(DP_OP_424J2_126_3477_n1651), .B(
        DP_OP_424J2_126_3477_n1566), .CI(DP_OP_424J2_126_3477_n1639), .CO(
        DP_OP_424J2_126_3477_n1495), .S(DP_OP_424J2_126_3477_n1496) );
  FADDX1_HVT DP_OP_424J2_126_3477_U844 ( .A(DP_OP_424J2_126_3477_n1647), .B(
        DP_OP_424J2_126_3477_n1568), .CI(DP_OP_424J2_126_3477_n1564), .CO(
        DP_OP_424J2_126_3477_n1493), .S(DP_OP_424J2_126_3477_n1494) );
  FADDX1_HVT DP_OP_424J2_126_3477_U843 ( .A(DP_OP_424J2_126_3477_n1645), .B(
        DP_OP_424J2_126_3477_n1578), .CI(DP_OP_424J2_126_3477_n1570), .CO(
        DP_OP_424J2_126_3477_n1491), .S(DP_OP_424J2_126_3477_n1492) );
  FADDX1_HVT DP_OP_424J2_126_3477_U842 ( .A(DP_OP_424J2_126_3477_n1643), .B(
        DP_OP_424J2_126_3477_n1576), .CI(DP_OP_424J2_126_3477_n1635), .CO(
        DP_OP_424J2_126_3477_n1489), .S(DP_OP_424J2_126_3477_n1490) );
  FADDX1_HVT DP_OP_424J2_126_3477_U841 ( .A(DP_OP_424J2_126_3477_n1562), .B(
        DP_OP_424J2_126_3477_n1538), .CI(DP_OP_424J2_126_3477_n1536), .CO(
        DP_OP_424J2_126_3477_n1487), .S(DP_OP_424J2_126_3477_n1488) );
  FADDX1_HVT DP_OP_424J2_126_3477_U840 ( .A(DP_OP_424J2_126_3477_n1558), .B(
        DP_OP_424J2_126_3477_n1560), .CI(DP_OP_424J2_126_3477_n1540), .CO(
        DP_OP_424J2_126_3477_n1485), .S(DP_OP_424J2_126_3477_n1486) );
  FADDX1_HVT DP_OP_424J2_126_3477_U839 ( .A(DP_OP_424J2_126_3477_n1552), .B(
        DP_OP_424J2_126_3477_n1546), .CI(DP_OP_424J2_126_3477_n1544), .CO(
        DP_OP_424J2_126_3477_n1483), .S(DP_OP_424J2_126_3477_n1484) );
  FADDX1_HVT DP_OP_424J2_126_3477_U838 ( .A(DP_OP_424J2_126_3477_n1548), .B(
        DP_OP_424J2_126_3477_n1542), .CI(DP_OP_424J2_126_3477_n1556), .CO(
        DP_OP_424J2_126_3477_n1481), .S(DP_OP_424J2_126_3477_n1482) );
  FADDX1_HVT DP_OP_424J2_126_3477_U837 ( .A(DP_OP_424J2_126_3477_n1550), .B(
        DP_OP_424J2_126_3477_n1554), .CI(DP_OP_424J2_126_3477_n1534), .CO(
        DP_OP_424J2_126_3477_n1479), .S(DP_OP_424J2_126_3477_n1480) );
  FADDX1_HVT DP_OP_424J2_126_3477_U836 ( .A(DP_OP_424J2_126_3477_n1532), .B(
        DP_OP_424J2_126_3477_n1520), .CI(DP_OP_424J2_126_3477_n1516), .CO(
        DP_OP_424J2_126_3477_n1477), .S(DP_OP_424J2_126_3477_n1478) );
  FADDX1_HVT DP_OP_424J2_126_3477_U835 ( .A(DP_OP_424J2_126_3477_n1528), .B(
        DP_OP_424J2_126_3477_n1522), .CI(DP_OP_424J2_126_3477_n1514), .CO(
        DP_OP_424J2_126_3477_n1475), .S(DP_OP_424J2_126_3477_n1476) );
  FADDX1_HVT DP_OP_424J2_126_3477_U834 ( .A(DP_OP_424J2_126_3477_n1526), .B(
        DP_OP_424J2_126_3477_n1524), .CI(DP_OP_424J2_126_3477_n1518), .CO(
        DP_OP_424J2_126_3477_n1473), .S(DP_OP_424J2_126_3477_n1474) );
  FADDX1_HVT DP_OP_424J2_126_3477_U833 ( .A(DP_OP_424J2_126_3477_n1530), .B(
        DP_OP_424J2_126_3477_n1512), .CI(DP_OP_424J2_126_3477_n1633), .CO(
        DP_OP_424J2_126_3477_n1471), .S(DP_OP_424J2_126_3477_n1472) );
  FADDX1_HVT DP_OP_424J2_126_3477_U832 ( .A(DP_OP_424J2_126_3477_n1631), .B(
        DP_OP_424J2_126_3477_n1629), .CI(DP_OP_424J2_126_3477_n1627), .CO(
        DP_OP_424J2_126_3477_n1469), .S(DP_OP_424J2_126_3477_n1470) );
  FADDX1_HVT DP_OP_424J2_126_3477_U831 ( .A(DP_OP_424J2_126_3477_n1625), .B(
        DP_OP_424J2_126_3477_n1623), .CI(DP_OP_424J2_126_3477_n1508), .CO(
        DP_OP_424J2_126_3477_n1467), .S(DP_OP_424J2_126_3477_n1468) );
  FADDX1_HVT DP_OP_424J2_126_3477_U830 ( .A(DP_OP_424J2_126_3477_n1621), .B(
        DP_OP_424J2_126_3477_n1510), .CI(DP_OP_424J2_126_3477_n1502), .CO(
        DP_OP_424J2_126_3477_n1465), .S(DP_OP_424J2_126_3477_n1466) );
  FADDX1_HVT DP_OP_424J2_126_3477_U829 ( .A(DP_OP_424J2_126_3477_n1619), .B(
        DP_OP_424J2_126_3477_n1506), .CI(DP_OP_424J2_126_3477_n1504), .CO(
        DP_OP_424J2_126_3477_n1463), .S(DP_OP_424J2_126_3477_n1464) );
  FADDX1_HVT DP_OP_424J2_126_3477_U828 ( .A(DP_OP_424J2_126_3477_n1617), .B(
        DP_OP_424J2_126_3477_n1615), .CI(DP_OP_424J2_126_3477_n1613), .CO(
        DP_OP_424J2_126_3477_n1461), .S(DP_OP_424J2_126_3477_n1462) );
  FADDX1_HVT DP_OP_424J2_126_3477_U827 ( .A(DP_OP_424J2_126_3477_n1611), .B(
        DP_OP_424J2_126_3477_n1492), .CI(DP_OP_424J2_126_3477_n1490), .CO(
        DP_OP_424J2_126_3477_n1459), .S(DP_OP_424J2_126_3477_n1460) );
  FADDX1_HVT DP_OP_424J2_126_3477_U826 ( .A(DP_OP_424J2_126_3477_n1496), .B(
        DP_OP_424J2_126_3477_n1498), .CI(DP_OP_424J2_126_3477_n1494), .CO(
        DP_OP_424J2_126_3477_n1457), .S(DP_OP_424J2_126_3477_n1458) );
  FADDX1_HVT DP_OP_424J2_126_3477_U825 ( .A(DP_OP_424J2_126_3477_n1609), .B(
        DP_OP_424J2_126_3477_n1607), .CI(DP_OP_424J2_126_3477_n1500), .CO(
        DP_OP_424J2_126_3477_n1455), .S(DP_OP_424J2_126_3477_n1456) );
  FADDX1_HVT DP_OP_424J2_126_3477_U824 ( .A(DP_OP_424J2_126_3477_n1488), .B(
        DP_OP_424J2_126_3477_n1480), .CI(DP_OP_424J2_126_3477_n1605), .CO(
        DP_OP_424J2_126_3477_n1453), .S(DP_OP_424J2_126_3477_n1454) );
  FADDX1_HVT DP_OP_424J2_126_3477_U823 ( .A(DP_OP_424J2_126_3477_n1486), .B(
        DP_OP_424J2_126_3477_n1484), .CI(DP_OP_424J2_126_3477_n1482), .CO(
        DP_OP_424J2_126_3477_n1451), .S(DP_OP_424J2_126_3477_n1452) );
  FADDX1_HVT DP_OP_424J2_126_3477_U822 ( .A(DP_OP_424J2_126_3477_n1478), .B(
        DP_OP_424J2_126_3477_n1474), .CI(DP_OP_424J2_126_3477_n1476), .CO(
        DP_OP_424J2_126_3477_n1449), .S(DP_OP_424J2_126_3477_n1450) );
  FADDX1_HVT DP_OP_424J2_126_3477_U821 ( .A(DP_OP_424J2_126_3477_n1472), .B(
        DP_OP_424J2_126_3477_n1603), .CI(DP_OP_424J2_126_3477_n1601), .CO(
        DP_OP_424J2_126_3477_n1447), .S(DP_OP_424J2_126_3477_n1448) );
  FADDX1_HVT DP_OP_424J2_126_3477_U820 ( .A(DP_OP_424J2_126_3477_n1599), .B(
        DP_OP_424J2_126_3477_n1470), .CI(DP_OP_424J2_126_3477_n1597), .CO(
        DP_OP_424J2_126_3477_n1445), .S(DP_OP_424J2_126_3477_n1446) );
  FADDX1_HVT DP_OP_424J2_126_3477_U819 ( .A(DP_OP_424J2_126_3477_n1468), .B(
        DP_OP_424J2_126_3477_n1595), .CI(DP_OP_424J2_126_3477_n1464), .CO(
        DP_OP_424J2_126_3477_n1443), .S(DP_OP_424J2_126_3477_n1444) );
  FADDX1_HVT DP_OP_424J2_126_3477_U818 ( .A(DP_OP_424J2_126_3477_n1466), .B(
        DP_OP_424J2_126_3477_n1462), .CI(DP_OP_424J2_126_3477_n1593), .CO(
        DP_OP_424J2_126_3477_n1441), .S(DP_OP_424J2_126_3477_n1442) );
  FADDX1_HVT DP_OP_424J2_126_3477_U817 ( .A(DP_OP_424J2_126_3477_n1460), .B(
        DP_OP_424J2_126_3477_n1458), .CI(DP_OP_424J2_126_3477_n1591), .CO(
        DP_OP_424J2_126_3477_n1439), .S(DP_OP_424J2_126_3477_n1440) );
  FADDX1_HVT DP_OP_424J2_126_3477_U816 ( .A(DP_OP_424J2_126_3477_n1456), .B(
        DP_OP_424J2_126_3477_n1454), .CI(DP_OP_424J2_126_3477_n1452), .CO(
        DP_OP_424J2_126_3477_n1437), .S(DP_OP_424J2_126_3477_n1438) );
  FADDX1_HVT DP_OP_424J2_126_3477_U815 ( .A(DP_OP_424J2_126_3477_n1450), .B(
        DP_OP_424J2_126_3477_n1589), .CI(DP_OP_424J2_126_3477_n1448), .CO(
        DP_OP_424J2_126_3477_n1435), .S(DP_OP_424J2_126_3477_n1436) );
  FADDX1_HVT DP_OP_424J2_126_3477_U814 ( .A(DP_OP_424J2_126_3477_n1587), .B(
        DP_OP_424J2_126_3477_n1446), .CI(DP_OP_424J2_126_3477_n1585), .CO(
        DP_OP_424J2_126_3477_n1433), .S(DP_OP_424J2_126_3477_n1434) );
  FADDX1_HVT DP_OP_424J2_126_3477_U813 ( .A(DP_OP_424J2_126_3477_n1444), .B(
        DP_OP_424J2_126_3477_n1442), .CI(DP_OP_424J2_126_3477_n1440), .CO(
        DP_OP_424J2_126_3477_n1431), .S(DP_OP_424J2_126_3477_n1432) );
  FADDX1_HVT DP_OP_424J2_126_3477_U812 ( .A(DP_OP_424J2_126_3477_n1438), .B(
        DP_OP_424J2_126_3477_n1583), .CI(DP_OP_424J2_126_3477_n1436), .CO(
        DP_OP_424J2_126_3477_n1429), .S(DP_OP_424J2_126_3477_n1430) );
  FADDX1_HVT DP_OP_424J2_126_3477_U811 ( .A(DP_OP_424J2_126_3477_n1581), .B(
        DP_OP_424J2_126_3477_n1434), .CI(DP_OP_424J2_126_3477_n1432), .CO(
        DP_OP_424J2_126_3477_n1427), .S(DP_OP_424J2_126_3477_n1428) );
  FADDX1_HVT DP_OP_424J2_126_3477_U810 ( .A(DP_OP_424J2_126_3477_n1579), .B(
        DP_OP_424J2_126_3477_n1828), .CI(DP_OP_424J2_126_3477_n2397), .CO(
        DP_OP_424J2_126_3477_n1425), .S(DP_OP_424J2_126_3477_n1426) );
  FADDX1_HVT DP_OP_424J2_126_3477_U809 ( .A(DP_OP_424J2_126_3477_n2354), .B(
        DP_OP_424J2_126_3477_n1916), .CI(DP_OP_424J2_126_3477_n1960), .CO(
        DP_OP_424J2_126_3477_n1423), .S(DP_OP_424J2_126_3477_n1424) );
  FADDX1_HVT DP_OP_424J2_126_3477_U808 ( .A(DP_OP_424J2_126_3477_n2705), .B(
        DP_OP_424J2_126_3477_n2573), .CI(DP_OP_424J2_126_3477_n2749), .CO(
        DP_OP_424J2_126_3477_n1421), .S(DP_OP_424J2_126_3477_n1422) );
  FADDX1_HVT DP_OP_424J2_126_3477_U807 ( .A(DP_OP_424J2_126_3477_n2004), .B(
        DP_OP_424J2_126_3477_n2485), .CI(DP_OP_424J2_126_3477_n2180), .CO(
        DP_OP_424J2_126_3477_n1419), .S(DP_OP_424J2_126_3477_n1420) );
  FADDX1_HVT DP_OP_424J2_126_3477_U806 ( .A(DP_OP_424J2_126_3477_n2661), .B(
        DP_OP_424J2_126_3477_n2048), .CI(DP_OP_424J2_126_3477_n2441), .CO(
        DP_OP_424J2_126_3477_n1417), .S(DP_OP_424J2_126_3477_n1418) );
  FADDX1_HVT DP_OP_424J2_126_3477_U805 ( .A(DP_OP_424J2_126_3477_n2312), .B(
        DP_OP_424J2_126_3477_n2881), .CI(DP_OP_424J2_126_3477_n2529), .CO(
        DP_OP_424J2_126_3477_n1415), .S(DP_OP_424J2_126_3477_n1416) );
  FADDX1_HVT DP_OP_424J2_126_3477_U804 ( .A(DP_OP_424J2_126_3477_n2837), .B(
        DP_OP_424J2_126_3477_n2136), .CI(DP_OP_424J2_126_3477_n2268), .CO(
        DP_OP_424J2_126_3477_n1413), .S(DP_OP_424J2_126_3477_n1414) );
  FADDX1_HVT DP_OP_424J2_126_3477_U803 ( .A(DP_OP_424J2_126_3477_n2617), .B(
        DP_OP_424J2_126_3477_n1872), .CI(DP_OP_424J2_126_3477_n2793), .CO(
        DP_OP_424J2_126_3477_n1411), .S(DP_OP_424J2_126_3477_n1412) );
  FADDX1_HVT DP_OP_424J2_126_3477_U802 ( .A(DP_OP_424J2_126_3477_n2092), .B(
        DP_OP_424J2_126_3477_n2224), .CI(DP_OP_424J2_126_3477_n1849), .CO(
        DP_OP_424J2_126_3477_n1409), .S(DP_OP_424J2_126_3477_n1410) );
  FADDX1_HVT DP_OP_424J2_126_3477_U801 ( .A(DP_OP_424J2_126_3477_n2462), .B(
        DP_OP_424J2_126_3477_n1967), .CI(DP_OP_424J2_126_3477_n2275), .CO(
        DP_OP_424J2_126_3477_n1407), .S(DP_OP_424J2_126_3477_n1408) );
  FADDX1_HVT DP_OP_424J2_126_3477_U800 ( .A(DP_OP_424J2_126_3477_n2594), .B(
        DP_OP_424J2_126_3477_n2726), .CI(DP_OP_424J2_126_3477_n2143), .CO(
        DP_OP_424J2_126_3477_n1405), .S(DP_OP_424J2_126_3477_n1406) );
  FADDX1_HVT DP_OP_424J2_126_3477_U799 ( .A(DP_OP_424J2_126_3477_n2201), .B(
        DP_OP_424J2_126_3477_n2536), .CI(DP_OP_424J2_126_3477_n2289), .CO(
        DP_OP_424J2_126_3477_n1403), .S(DP_OP_424J2_126_3477_n1404) );
  FADDX1_HVT DP_OP_424J2_126_3477_U798 ( .A(DP_OP_424J2_126_3477_n2333), .B(
        DP_OP_424J2_126_3477_n2411), .CI(DP_OP_424J2_126_3477_n2069), .CO(
        DP_OP_424J2_126_3477_n1401), .S(DP_OP_424J2_126_3477_n1402) );
  FADDX1_HVT DP_OP_424J2_126_3477_U797 ( .A(DP_OP_424J2_126_3477_n2888), .B(
        DP_OP_424J2_126_3477_n2150), .CI(DP_OP_424J2_126_3477_n2506), .CO(
        DP_OP_424J2_126_3477_n1399), .S(DP_OP_424J2_126_3477_n1400) );
  FADDX1_HVT DP_OP_424J2_126_3477_U796 ( .A(DP_OP_424J2_126_3477_n2550), .B(
        DP_OP_424J2_126_3477_n1784), .CI(DP_OP_424J2_126_3477_n2231), .CO(
        DP_OP_424J2_126_3477_n1397), .S(DP_OP_424J2_126_3477_n1398) );
  FADDX1_HVT DP_OP_424J2_126_3477_U795 ( .A(DP_OP_424J2_126_3477_n2418), .B(
        DP_OP_424J2_126_3477_n2062), .CI(DP_OP_424J2_126_3477_n2770), .CO(
        DP_OP_424J2_126_3477_n1395), .S(DP_OP_424J2_126_3477_n1396) );
  FADDX1_HVT DP_OP_424J2_126_3477_U794 ( .A(DP_OP_424J2_126_3477_n2638), .B(
        DP_OP_424J2_126_3477_n2587), .CI(DP_OP_424J2_126_3477_n2099), .CO(
        DP_OP_424J2_126_3477_n1393), .S(DP_OP_424J2_126_3477_n1394) );
  FADDX1_HVT DP_OP_424J2_126_3477_U793 ( .A(DP_OP_424J2_126_3477_n2844), .B(
        DP_OP_424J2_126_3477_n1981), .CI(DP_OP_424J2_126_3477_n1893), .CO(
        DP_OP_424J2_126_3477_n1391), .S(DP_OP_424J2_126_3477_n1392) );
  FADDX1_HVT DP_OP_424J2_126_3477_U792 ( .A(DP_OP_424J2_126_3477_n2113), .B(
        DP_OP_424J2_126_3477_n2326), .CI(DP_OP_424J2_126_3477_n2858), .CO(
        DP_OP_424J2_126_3477_n1389), .S(DP_OP_424J2_126_3477_n1390) );
  FADDX1_HVT DP_OP_424J2_126_3477_U791 ( .A(DP_OP_424J2_126_3477_n1842), .B(
        DP_OP_424J2_126_3477_n2025), .CI(DP_OP_424J2_126_3477_n2448), .CO(
        DP_OP_424J2_126_3477_n1387), .S(DP_OP_424J2_126_3477_n1388) );
  FADDX1_HVT DP_OP_424J2_126_3477_U790 ( .A(DP_OP_424J2_126_3477_n2682), .B(
        DP_OP_424J2_126_3477_n2631), .CI(DP_OP_424J2_126_3477_n2580), .CO(
        DP_OP_424J2_126_3477_n1385), .S(DP_OP_424J2_126_3477_n1386) );
  FADDX1_HVT DP_OP_424J2_126_3477_U789 ( .A(DP_OP_424J2_126_3477_n2756), .B(
        DP_OP_424J2_126_3477_n2499), .CI(DP_OP_424J2_126_3477_n1937), .CO(
        DP_OP_424J2_126_3477_n1383), .S(DP_OP_424J2_126_3477_n1384) );
  FADDX1_HVT DP_OP_424J2_126_3477_U788 ( .A(DP_OP_424J2_126_3477_n2543), .B(
        DP_OP_424J2_126_3477_n2763), .CI(DP_OP_424J2_126_3477_n2238), .CO(
        DP_OP_424J2_126_3477_n1381), .S(DP_OP_424J2_126_3477_n1382) );
  FADDX1_HVT DP_OP_424J2_126_3477_U787 ( .A(DP_OP_424J2_126_3477_n2712), .B(
        DP_OP_424J2_126_3477_n2455), .CI(DP_OP_424J2_126_3477_n2194), .CO(
        DP_OP_424J2_126_3477_n1379), .S(DP_OP_424J2_126_3477_n1380) );
  FADDX1_HVT DP_OP_424J2_126_3477_U786 ( .A(DP_OP_424J2_126_3477_n2851), .B(
        DP_OP_424J2_126_3477_n2807), .CI(DP_OP_424J2_126_3477_n2011), .CO(
        DP_OP_424J2_126_3477_n1377), .S(DP_OP_424J2_126_3477_n1378) );
  FADDX1_HVT DP_OP_424J2_126_3477_U785 ( .A(DP_OP_424J2_126_3477_n1886), .B(
        DP_OP_424J2_126_3477_n2282), .CI(DP_OP_424J2_126_3477_n2367), .CO(
        DP_OP_424J2_126_3477_n1375), .S(DP_OP_424J2_126_3477_n1376) );
  FADDX1_HVT DP_OP_424J2_126_3477_U784 ( .A(DP_OP_424J2_126_3477_n2106), .B(
        DP_OP_424J2_126_3477_n2668), .CI(DP_OP_424J2_126_3477_n1930), .CO(
        DP_OP_424J2_126_3477_n1373), .S(DP_OP_424J2_126_3477_n1374) );
  FADDX1_HVT DP_OP_424J2_126_3477_U783 ( .A(DP_OP_424J2_126_3477_n2492), .B(
        DP_OP_424J2_126_3477_n2895), .CI(DP_OP_424J2_126_3477_n2902), .CO(
        DP_OP_424J2_126_3477_n1371), .S(DP_OP_424J2_126_3477_n1372) );
  FADDX1_HVT DP_OP_424J2_126_3477_U782 ( .A(DP_OP_424J2_126_3477_n2360), .B(
        DP_OP_424J2_126_3477_n2245), .CI(DP_OP_424J2_126_3477_n2719), .CO(
        DP_OP_424J2_126_3477_n1369), .S(DP_OP_424J2_126_3477_n1370) );
  FADDX1_HVT DP_OP_424J2_126_3477_U781 ( .A(DP_OP_424J2_126_3477_n2675), .B(
        DP_OP_424J2_126_3477_n2055), .CI(DP_OP_424J2_126_3477_n2374), .CO(
        DP_OP_424J2_126_3477_n1367), .S(DP_OP_424J2_126_3477_n1368) );
  FADDX1_HVT DP_OP_424J2_126_3477_U780 ( .A(DP_OP_424J2_126_3477_n2319), .B(
        DP_OP_424J2_126_3477_n2624), .CI(DP_OP_424J2_126_3477_n2018), .CO(
        DP_OP_424J2_126_3477_n1365), .S(DP_OP_424J2_126_3477_n1366) );
  FADDX1_HVT DP_OP_424J2_126_3477_U779 ( .A(DP_OP_424J2_126_3477_n1974), .B(
        DP_OP_424J2_126_3477_n2157), .CI(DP_OP_424J2_126_3477_n2814), .CO(
        DP_OP_424J2_126_3477_n1363), .S(DP_OP_424J2_126_3477_n1364) );
  FADDX1_HVT DP_OP_424J2_126_3477_U778 ( .A(DP_OP_424J2_126_3477_n2800), .B(
        DP_OP_424J2_126_3477_n1923), .CI(DP_OP_424J2_126_3477_n2404), .CO(
        DP_OP_424J2_126_3477_n1361), .S(DP_OP_424J2_126_3477_n1362) );
  FADDX1_HVT DP_OP_424J2_126_3477_U777 ( .A(DP_OP_424J2_126_3477_n1879), .B(
        DP_OP_424J2_126_3477_n1835), .CI(DP_OP_424J2_126_3477_n2187), .CO(
        DP_OP_424J2_126_3477_n1359), .S(DP_OP_424J2_126_3477_n1360) );
  FADDX1_HVT DP_OP_424J2_126_3477_U776 ( .A(DP_OP_424J2_126_3477_n1577), .B(
        DP_OP_424J2_126_3477_n1563), .CI(DP_OP_424J2_126_3477_n1565), .CO(
        DP_OP_424J2_126_3477_n1357), .S(DP_OP_424J2_126_3477_n1358) );
  FADDX1_HVT DP_OP_424J2_126_3477_U775 ( .A(DP_OP_424J2_126_3477_n1575), .B(
        DP_OP_424J2_126_3477_n1567), .CI(DP_OP_424J2_126_3477_n1569), .CO(
        DP_OP_424J2_126_3477_n1355), .S(DP_OP_424J2_126_3477_n1356) );
  FADDX1_HVT DP_OP_424J2_126_3477_U774 ( .A(DP_OP_424J2_126_3477_n1573), .B(
        DP_OP_424J2_126_3477_n1571), .CI(DP_OP_424J2_126_3477_n1561), .CO(
        DP_OP_424J2_126_3477_n1353), .S(DP_OP_424J2_126_3477_n1354) );
  FADDX1_HVT DP_OP_424J2_126_3477_U773 ( .A(DP_OP_424J2_126_3477_n1559), .B(
        DP_OP_424J2_126_3477_n1537), .CI(DP_OP_424J2_126_3477_n1535), .CO(
        DP_OP_424J2_126_3477_n1351), .S(DP_OP_424J2_126_3477_n1352) );
  FADDX1_HVT DP_OP_424J2_126_3477_U772 ( .A(DP_OP_424J2_126_3477_n1539), .B(
        DP_OP_424J2_126_3477_n1541), .CI(DP_OP_424J2_126_3477_n1543), .CO(
        DP_OP_424J2_126_3477_n1349), .S(DP_OP_424J2_126_3477_n1350) );
  FADDX1_HVT DP_OP_424J2_126_3477_U771 ( .A(DP_OP_424J2_126_3477_n1557), .B(
        DP_OP_424J2_126_3477_n1545), .CI(DP_OP_424J2_126_3477_n1547), .CO(
        DP_OP_424J2_126_3477_n1347), .S(DP_OP_424J2_126_3477_n1348) );
  FADDX1_HVT DP_OP_424J2_126_3477_U770 ( .A(DP_OP_424J2_126_3477_n1555), .B(
        DP_OP_424J2_126_3477_n1549), .CI(DP_OP_424J2_126_3477_n1551), .CO(
        DP_OP_424J2_126_3477_n1345), .S(DP_OP_424J2_126_3477_n1346) );
  FADDX1_HVT DP_OP_424J2_126_3477_U769 ( .A(DP_OP_424J2_126_3477_n1553), .B(
        DP_OP_424J2_126_3477_n1533), .CI(DP_OP_424J2_126_3477_n1531), .CO(
        DP_OP_424J2_126_3477_n1343), .S(DP_OP_424J2_126_3477_n1344) );
  FADDX1_HVT DP_OP_424J2_126_3477_U768 ( .A(DP_OP_424J2_126_3477_n1527), .B(
        DP_OP_424J2_126_3477_n1414), .CI(DP_OP_424J2_126_3477_n1515), .CO(
        DP_OP_424J2_126_3477_n1341), .S(DP_OP_424J2_126_3477_n1342) );
  FADDX1_HVT DP_OP_424J2_126_3477_U767 ( .A(DP_OP_424J2_126_3477_n1529), .B(
        DP_OP_424J2_126_3477_n1412), .CI(DP_OP_424J2_126_3477_n1513), .CO(
        DP_OP_424J2_126_3477_n1339), .S(DP_OP_424J2_126_3477_n1340) );
  FADDX1_HVT DP_OP_424J2_126_3477_U766 ( .A(DP_OP_424J2_126_3477_n1525), .B(
        DP_OP_424J2_126_3477_n1418), .CI(DP_OP_424J2_126_3477_n1517), .CO(
        DP_OP_424J2_126_3477_n1337), .S(DP_OP_424J2_126_3477_n1338) );
  FADDX1_HVT DP_OP_424J2_126_3477_U765 ( .A(DP_OP_424J2_126_3477_n1523), .B(
        DP_OP_424J2_126_3477_n1420), .CI(DP_OP_424J2_126_3477_n1416), .CO(
        DP_OP_424J2_126_3477_n1335), .S(DP_OP_424J2_126_3477_n1336) );
  FADDX1_HVT DP_OP_424J2_126_3477_U764 ( .A(DP_OP_424J2_126_3477_n1521), .B(
        DP_OP_424J2_126_3477_n1426), .CI(DP_OP_424J2_126_3477_n1422), .CO(
        DP_OP_424J2_126_3477_n1333), .S(DP_OP_424J2_126_3477_n1334) );
  FADDX1_HVT DP_OP_424J2_126_3477_U763 ( .A(DP_OP_424J2_126_3477_n1519), .B(
        DP_OP_424J2_126_3477_n1424), .CI(DP_OP_424J2_126_3477_n1410), .CO(
        DP_OP_424J2_126_3477_n1331), .S(DP_OP_424J2_126_3477_n1332) );
  FADDX1_HVT DP_OP_424J2_126_3477_U762 ( .A(DP_OP_424J2_126_3477_n1511), .B(
        DP_OP_424J2_126_3477_n1388), .CI(DP_OP_424J2_126_3477_n1384), .CO(
        DP_OP_424J2_126_3477_n1329), .S(DP_OP_424J2_126_3477_n1330) );
  FADDX1_HVT DP_OP_424J2_126_3477_U761 ( .A(DP_OP_424J2_126_3477_n1402), .B(
        DP_OP_424J2_126_3477_n1398), .CI(DP_OP_424J2_126_3477_n1386), .CO(
        DP_OP_424J2_126_3477_n1327), .S(DP_OP_424J2_126_3477_n1328) );
  FADDX1_HVT DP_OP_424J2_126_3477_U760 ( .A(DP_OP_424J2_126_3477_n1400), .B(
        DP_OP_424J2_126_3477_n1390), .CI(DP_OP_424J2_126_3477_n1394), .CO(
        DP_OP_424J2_126_3477_n1325), .S(DP_OP_424J2_126_3477_n1326) );
  FADDX1_HVT DP_OP_424J2_126_3477_U759 ( .A(DP_OP_424J2_126_3477_n1396), .B(
        DP_OP_424J2_126_3477_n1408), .CI(DP_OP_424J2_126_3477_n1404), .CO(
        DP_OP_424J2_126_3477_n1323), .S(DP_OP_424J2_126_3477_n1324) );
  FADDX1_HVT DP_OP_424J2_126_3477_U758 ( .A(DP_OP_424J2_126_3477_n1406), .B(
        DP_OP_424J2_126_3477_n1392), .CI(DP_OP_424J2_126_3477_n1382), .CO(
        DP_OP_424J2_126_3477_n1321), .S(DP_OP_424J2_126_3477_n1322) );
  FADDX1_HVT DP_OP_424J2_126_3477_U757 ( .A(DP_OP_424J2_126_3477_n1380), .B(
        DP_OP_424J2_126_3477_n1366), .CI(DP_OP_424J2_126_3477_n1360), .CO(
        DP_OP_424J2_126_3477_n1319), .S(DP_OP_424J2_126_3477_n1320) );
  FADDX1_HVT DP_OP_424J2_126_3477_U756 ( .A(DP_OP_424J2_126_3477_n1378), .B(
        DP_OP_424J2_126_3477_n1368), .CI(DP_OP_424J2_126_3477_n1364), .CO(
        DP_OP_424J2_126_3477_n1317), .S(DP_OP_424J2_126_3477_n1318) );
  FADDX1_HVT DP_OP_424J2_126_3477_U755 ( .A(DP_OP_424J2_126_3477_n1376), .B(
        DP_OP_424J2_126_3477_n1370), .CI(DP_OP_424J2_126_3477_n1362), .CO(
        DP_OP_424J2_126_3477_n1315), .S(DP_OP_424J2_126_3477_n1316) );
  FADDX1_HVT DP_OP_424J2_126_3477_U754 ( .A(DP_OP_424J2_126_3477_n1372), .B(
        DP_OP_424J2_126_3477_n1374), .CI(DP_OP_424J2_126_3477_n1509), .CO(
        DP_OP_424J2_126_3477_n1313), .S(DP_OP_424J2_126_3477_n1314) );
  FADDX1_HVT DP_OP_424J2_126_3477_U753 ( .A(DP_OP_424J2_126_3477_n1507), .B(
        DP_OP_424J2_126_3477_n1505), .CI(DP_OP_424J2_126_3477_n1501), .CO(
        DP_OP_424J2_126_3477_n1311), .S(DP_OP_424J2_126_3477_n1312) );
  FADDX1_HVT DP_OP_424J2_126_3477_U752 ( .A(DP_OP_424J2_126_3477_n1503), .B(
        DP_OP_424J2_126_3477_n1499), .CI(DP_OP_424J2_126_3477_n1497), .CO(
        DP_OP_424J2_126_3477_n1309), .S(DP_OP_424J2_126_3477_n1310) );
  FADDX1_HVT DP_OP_424J2_126_3477_U751 ( .A(DP_OP_424J2_126_3477_n1495), .B(
        DP_OP_424J2_126_3477_n1356), .CI(DP_OP_424J2_126_3477_n1354), .CO(
        DP_OP_424J2_126_3477_n1307), .S(DP_OP_424J2_126_3477_n1308) );
  FADDX1_HVT DP_OP_424J2_126_3477_U750 ( .A(DP_OP_424J2_126_3477_n1493), .B(
        DP_OP_424J2_126_3477_n1489), .CI(DP_OP_424J2_126_3477_n1358), .CO(
        DP_OP_424J2_126_3477_n1305), .S(DP_OP_424J2_126_3477_n1306) );
  FADDX1_HVT DP_OP_424J2_126_3477_U749 ( .A(DP_OP_424J2_126_3477_n1491), .B(
        DP_OP_424J2_126_3477_n1487), .CI(DP_OP_424J2_126_3477_n1485), .CO(
        DP_OP_424J2_126_3477_n1303), .S(DP_OP_424J2_126_3477_n1304) );
  FADDX1_HVT DP_OP_424J2_126_3477_U748 ( .A(DP_OP_424J2_126_3477_n1483), .B(
        DP_OP_424J2_126_3477_n1350), .CI(DP_OP_424J2_126_3477_n1344), .CO(
        DP_OP_424J2_126_3477_n1301), .S(DP_OP_424J2_126_3477_n1302) );
  FADDX1_HVT DP_OP_424J2_126_3477_U747 ( .A(DP_OP_424J2_126_3477_n1481), .B(
        DP_OP_424J2_126_3477_n1352), .CI(DP_OP_424J2_126_3477_n1348), .CO(
        DP_OP_424J2_126_3477_n1299), .S(DP_OP_424J2_126_3477_n1300) );
  FADDX1_HVT DP_OP_424J2_126_3477_U746 ( .A(DP_OP_424J2_126_3477_n1479), .B(
        DP_OP_424J2_126_3477_n1346), .CI(DP_OP_424J2_126_3477_n1477), .CO(
        DP_OP_424J2_126_3477_n1297), .S(DP_OP_424J2_126_3477_n1298) );
  FADDX1_HVT DP_OP_424J2_126_3477_U745 ( .A(DP_OP_424J2_126_3477_n1475), .B(
        DP_OP_424J2_126_3477_n1332), .CI(DP_OP_424J2_126_3477_n1471), .CO(
        DP_OP_424J2_126_3477_n1295), .S(DP_OP_424J2_126_3477_n1296) );
  FADDX1_HVT DP_OP_424J2_126_3477_U744 ( .A(DP_OP_424J2_126_3477_n1338), .B(
        DP_OP_424J2_126_3477_n1336), .CI(DP_OP_424J2_126_3477_n1334), .CO(
        DP_OP_424J2_126_3477_n1293), .S(DP_OP_424J2_126_3477_n1294) );
  FADDX1_HVT DP_OP_424J2_126_3477_U743 ( .A(DP_OP_424J2_126_3477_n1473), .B(
        DP_OP_424J2_126_3477_n1342), .CI(DP_OP_424J2_126_3477_n1340), .CO(
        DP_OP_424J2_126_3477_n1291), .S(DP_OP_424J2_126_3477_n1292) );
  FADDX1_HVT DP_OP_424J2_126_3477_U742 ( .A(DP_OP_424J2_126_3477_n1330), .B(
        DP_OP_424J2_126_3477_n1328), .CI(DP_OP_424J2_126_3477_n1322), .CO(
        DP_OP_424J2_126_3477_n1289), .S(DP_OP_424J2_126_3477_n1290) );
  FADDX1_HVT DP_OP_424J2_126_3477_U741 ( .A(DP_OP_424J2_126_3477_n1324), .B(
        DP_OP_424J2_126_3477_n1326), .CI(DP_OP_424J2_126_3477_n1320), .CO(
        DP_OP_424J2_126_3477_n1287), .S(DP_OP_424J2_126_3477_n1288) );
  FADDX1_HVT DP_OP_424J2_126_3477_U740 ( .A(DP_OP_424J2_126_3477_n1318), .B(
        DP_OP_424J2_126_3477_n1316), .CI(DP_OP_424J2_126_3477_n1469), .CO(
        DP_OP_424J2_126_3477_n1285), .S(DP_OP_424J2_126_3477_n1286) );
  FADDX1_HVT DP_OP_424J2_126_3477_U739 ( .A(DP_OP_424J2_126_3477_n1467), .B(
        DP_OP_424J2_126_3477_n1314), .CI(DP_OP_424J2_126_3477_n1465), .CO(
        DP_OP_424J2_126_3477_n1283), .S(DP_OP_424J2_126_3477_n1284) );
  FADDX1_HVT DP_OP_424J2_126_3477_U738 ( .A(DP_OP_424J2_126_3477_n1463), .B(
        DP_OP_424J2_126_3477_n1312), .CI(DP_OP_424J2_126_3477_n1310), .CO(
        DP_OP_424J2_126_3477_n1281), .S(DP_OP_424J2_126_3477_n1282) );
  FADDX1_HVT DP_OP_424J2_126_3477_U737 ( .A(DP_OP_424J2_126_3477_n1461), .B(
        DP_OP_424J2_126_3477_n1459), .CI(DP_OP_424J2_126_3477_n1457), .CO(
        DP_OP_424J2_126_3477_n1279), .S(DP_OP_424J2_126_3477_n1280) );
  FADDX1_HVT DP_OP_424J2_126_3477_U736 ( .A(DP_OP_424J2_126_3477_n1455), .B(
        DP_OP_424J2_126_3477_n1308), .CI(DP_OP_424J2_126_3477_n1306), .CO(
        DP_OP_424J2_126_3477_n1277), .S(DP_OP_424J2_126_3477_n1278) );
  FADDX1_HVT DP_OP_424J2_126_3477_U735 ( .A(DP_OP_424J2_126_3477_n1304), .B(
        DP_OP_424J2_126_3477_n1453), .CI(DP_OP_424J2_126_3477_n1298), .CO(
        DP_OP_424J2_126_3477_n1275), .S(DP_OP_424J2_126_3477_n1276) );
  FADDX1_HVT DP_OP_424J2_126_3477_U734 ( .A(DP_OP_424J2_126_3477_n1451), .B(
        DP_OP_424J2_126_3477_n1302), .CI(DP_OP_424J2_126_3477_n1300), .CO(
        DP_OP_424J2_126_3477_n1273), .S(DP_OP_424J2_126_3477_n1274) );
  FADDX1_HVT DP_OP_424J2_126_3477_U733 ( .A(DP_OP_424J2_126_3477_n1449), .B(
        DP_OP_424J2_126_3477_n1294), .CI(DP_OP_424J2_126_3477_n1296), .CO(
        DP_OP_424J2_126_3477_n1271), .S(DP_OP_424J2_126_3477_n1272) );
  FADDX1_HVT DP_OP_424J2_126_3477_U732 ( .A(DP_OP_424J2_126_3477_n1292), .B(
        DP_OP_424J2_126_3477_n1290), .CI(DP_OP_424J2_126_3477_n1447), .CO(
        DP_OP_424J2_126_3477_n1269), .S(DP_OP_424J2_126_3477_n1270) );
  FADDX1_HVT DP_OP_424J2_126_3477_U731 ( .A(DP_OP_424J2_126_3477_n1288), .B(
        DP_OP_424J2_126_3477_n1286), .CI(DP_OP_424J2_126_3477_n1445), .CO(
        DP_OP_424J2_126_3477_n1267), .S(DP_OP_424J2_126_3477_n1268) );
  FADDX1_HVT DP_OP_424J2_126_3477_U730 ( .A(DP_OP_424J2_126_3477_n1284), .B(
        DP_OP_424J2_126_3477_n1443), .CI(DP_OP_424J2_126_3477_n1282), .CO(
        DP_OP_424J2_126_3477_n1265), .S(DP_OP_424J2_126_3477_n1266) );
  FADDX1_HVT DP_OP_424J2_126_3477_U729 ( .A(DP_OP_424J2_126_3477_n1441), .B(
        DP_OP_424J2_126_3477_n1280), .CI(DP_OP_424J2_126_3477_n1439), .CO(
        DP_OP_424J2_126_3477_n1263), .S(DP_OP_424J2_126_3477_n1264) );
  FADDX1_HVT DP_OP_424J2_126_3477_U728 ( .A(DP_OP_424J2_126_3477_n1278), .B(
        DP_OP_424J2_126_3477_n1437), .CI(DP_OP_424J2_126_3477_n1276), .CO(
        DP_OP_424J2_126_3477_n1261), .S(DP_OP_424J2_126_3477_n1262) );
  FADDX1_HVT DP_OP_424J2_126_3477_U727 ( .A(DP_OP_424J2_126_3477_n1274), .B(
        DP_OP_424J2_126_3477_n1272), .CI(DP_OP_424J2_126_3477_n1435), .CO(
        DP_OP_424J2_126_3477_n1259), .S(DP_OP_424J2_126_3477_n1260) );
  FADDX1_HVT DP_OP_424J2_126_3477_U726 ( .A(DP_OP_424J2_126_3477_n1270), .B(
        DP_OP_424J2_126_3477_n1268), .CI(DP_OP_424J2_126_3477_n1433), .CO(
        DP_OP_424J2_126_3477_n1257), .S(DP_OP_424J2_126_3477_n1258) );
  FADDX1_HVT DP_OP_424J2_126_3477_U725 ( .A(DP_OP_424J2_126_3477_n1266), .B(
        DP_OP_424J2_126_3477_n1431), .CI(DP_OP_424J2_126_3477_n1264), .CO(
        DP_OP_424J2_126_3477_n1255), .S(DP_OP_424J2_126_3477_n1256) );
  FADDX1_HVT DP_OP_424J2_126_3477_U724 ( .A(DP_OP_424J2_126_3477_n1262), .B(
        DP_OP_424J2_126_3477_n1429), .CI(DP_OP_424J2_126_3477_n1260), .CO(
        DP_OP_424J2_126_3477_n1253), .S(DP_OP_424J2_126_3477_n1254) );
  FADDX1_HVT DP_OP_424J2_126_3477_U723 ( .A(DP_OP_424J2_126_3477_n1258), .B(
        DP_OP_424J2_126_3477_n1427), .CI(DP_OP_424J2_126_3477_n1256), .CO(
        DP_OP_424J2_126_3477_n1251), .S(DP_OP_424J2_126_3477_n1252) );
  HADDX1_HVT DP_OP_424J2_126_3477_U722 ( .A0(DP_OP_424J2_126_3477_n2353), .B0(
        DP_OP_424J2_126_3477_n2440), .C1(DP_OP_424J2_126_3477_n1249), .SO(
        DP_OP_424J2_126_3477_n1250) );
  FADDX1_HVT DP_OP_424J2_126_3477_U721 ( .A(DP_OP_424J2_126_3477_n2003), .B(
        DP_OP_424J2_126_3477_n1827), .CI(DP_OP_424J2_126_3477_n2396), .CO(
        DP_OP_424J2_126_3477_n1247), .S(DP_OP_424J2_126_3477_n1248) );
  FADDX1_HVT DP_OP_424J2_126_3477_U720 ( .A(DP_OP_424J2_126_3477_n2704), .B(
        DP_OP_424J2_126_3477_n2047), .CI(DP_OP_424J2_126_3477_n1959), .CO(
        DP_OP_424J2_126_3477_n1245), .S(DP_OP_424J2_126_3477_n1246) );
  FADDX1_HVT DP_OP_424J2_126_3477_U719 ( .A(DP_OP_424J2_126_3477_n2836), .B(
        DP_OP_424J2_126_3477_n2179), .CI(DP_OP_424J2_126_3477_n2748), .CO(
        DP_OP_424J2_126_3477_n1243), .S(DP_OP_424J2_126_3477_n1244) );
  FADDX1_HVT DP_OP_424J2_126_3477_U718 ( .A(DP_OP_424J2_126_3477_n2311), .B(
        DP_OP_424J2_126_3477_n2484), .CI(DP_OP_424J2_126_3477_n1915), .CO(
        DP_OP_424J2_126_3477_n1241), .S(DP_OP_424J2_126_3477_n1242) );
  FADDX1_HVT DP_OP_424J2_126_3477_U717 ( .A(DP_OP_424J2_126_3477_n2091), .B(
        DP_OP_424J2_126_3477_n2528), .CI(DP_OP_424J2_126_3477_n2572), .CO(
        DP_OP_424J2_126_3477_n1239), .S(DP_OP_424J2_126_3477_n1240) );
  FADDX1_HVT DP_OP_424J2_126_3477_U716 ( .A(DP_OP_424J2_126_3477_n2135), .B(
        DP_OP_424J2_126_3477_n2267), .CI(DP_OP_424J2_126_3477_n2880), .CO(
        DP_OP_424J2_126_3477_n1237), .S(DP_OP_424J2_126_3477_n1238) );
  FADDX1_HVT DP_OP_424J2_126_3477_U715 ( .A(DP_OP_424J2_126_3477_n1871), .B(
        DP_OP_424J2_126_3477_n2792), .CI(DP_OP_424J2_126_3477_n2616), .CO(
        DP_OP_424J2_126_3477_n1235), .S(DP_OP_424J2_126_3477_n1236) );
  FADDX1_HVT DP_OP_424J2_126_3477_U714 ( .A(DP_OP_424J2_126_3477_n2660), .B(
        DP_OP_424J2_126_3477_n2223), .CI(DP_OP_424J2_126_3477_n2637), .CO(
        DP_OP_424J2_126_3477_n1233), .S(DP_OP_424J2_126_3477_n1234) );
  FADDX1_HVT DP_OP_424J2_126_3477_U713 ( .A(DP_OP_424J2_126_3477_n2461), .B(
        DP_OP_424J2_126_3477_n2535), .CI(DP_OP_424J2_126_3477_n2288), .CO(
        DP_OP_424J2_126_3477_n1231), .S(DP_OP_424J2_126_3477_n1232) );
  FADDX1_HVT DP_OP_424J2_126_3477_U712 ( .A(DP_OP_424J2_126_3477_n2593), .B(
        DP_OP_424J2_126_3477_n1966), .CI(DP_OP_424J2_126_3477_n2274), .CO(
        DP_OP_424J2_126_3477_n1229), .S(DP_OP_424J2_126_3477_n1230) );
  FADDX1_HVT DP_OP_424J2_126_3477_U711 ( .A(DP_OP_424J2_126_3477_n2332), .B(
        DP_OP_424J2_126_3477_n2410), .CI(DP_OP_424J2_126_3477_n2142), .CO(
        DP_OP_424J2_126_3477_n1227), .S(DP_OP_424J2_126_3477_n1228) );
  FADDX1_HVT DP_OP_424J2_126_3477_U710 ( .A(DP_OP_424J2_126_3477_n1848), .B(
        DP_OP_424J2_126_3477_n2725), .CI(DP_OP_424J2_126_3477_n2068), .CO(
        DP_OP_424J2_126_3477_n1225), .S(DP_OP_424J2_126_3477_n1226) );
  FADDX1_HVT DP_OP_424J2_126_3477_U709 ( .A(DP_OP_424J2_126_3477_n2112), .B(
        DP_OP_424J2_126_3477_n2149), .CI(DP_OP_424J2_126_3477_n2505), .CO(
        DP_OP_424J2_126_3477_n1223), .S(DP_OP_424J2_126_3477_n1224) );
  FADDX1_HVT DP_OP_424J2_126_3477_U708 ( .A(DP_OP_424J2_126_3477_n2549), .B(
        DP_OP_424J2_126_3477_n1783), .CI(DP_OP_424J2_126_3477_n1892), .CO(
        DP_OP_424J2_126_3477_n1221), .S(DP_OP_424J2_126_3477_n1222) );
  FADDX1_HVT DP_OP_424J2_126_3477_U707 ( .A(DP_OP_424J2_126_3477_n2417), .B(
        DP_OP_424J2_126_3477_n1841), .CI(DP_OP_424J2_126_3477_n2447), .CO(
        DP_OP_424J2_126_3477_n1219), .S(DP_OP_424J2_126_3477_n1220) );
  FADDX1_HVT DP_OP_424J2_126_3477_U706 ( .A(DP_OP_424J2_126_3477_n2200), .B(
        DP_OP_424J2_126_3477_n2755), .CI(DP_OP_424J2_126_3477_n2230), .CO(
        DP_OP_424J2_126_3477_n1217), .S(DP_OP_424J2_126_3477_n1218) );
  FADDX1_HVT DP_OP_424J2_126_3477_U705 ( .A(DP_OP_424J2_126_3477_n2887), .B(
        DP_OP_424J2_126_3477_n2498), .CI(DP_OP_424J2_126_3477_n2769), .CO(
        DP_OP_424J2_126_3477_n1215), .S(DP_OP_424J2_126_3477_n1216) );
  FADDX1_HVT DP_OP_424J2_126_3477_U704 ( .A(DP_OP_424J2_126_3477_n2843), .B(
        DP_OP_424J2_126_3477_n2061), .CI(DP_OP_424J2_126_3477_n2098), .CO(
        DP_OP_424J2_126_3477_n1213), .S(DP_OP_424J2_126_3477_n1214) );
  FADDX1_HVT DP_OP_424J2_126_3477_U703 ( .A(DP_OP_424J2_126_3477_n2024), .B(
        DP_OP_424J2_126_3477_n1980), .CI(DP_OP_424J2_126_3477_n2857), .CO(
        DP_OP_424J2_126_3477_n1211), .S(DP_OP_424J2_126_3477_n1212) );
  FADDX1_HVT DP_OP_424J2_126_3477_U702 ( .A(DP_OP_424J2_126_3477_n2325), .B(
        DP_OP_424J2_126_3477_n2630), .CI(DP_OP_424J2_126_3477_n2579), .CO(
        DP_OP_424J2_126_3477_n1209), .S(DP_OP_424J2_126_3477_n1210) );
  FADDX1_HVT DP_OP_424J2_126_3477_U701 ( .A(DP_OP_424J2_126_3477_n2681), .B(
        DP_OP_424J2_126_3477_n2586), .CI(DP_OP_424J2_126_3477_n1936), .CO(
        DP_OP_424J2_126_3477_n1207), .S(DP_OP_424J2_126_3477_n1208) );
  FADDX1_HVT DP_OP_424J2_126_3477_U700 ( .A(DP_OP_424J2_126_3477_n2711), .B(
        DP_OP_424J2_126_3477_n2762), .CI(DP_OP_424J2_126_3477_n2366), .CO(
        DP_OP_424J2_126_3477_n1205), .S(DP_OP_424J2_126_3477_n1206) );
  FADDX1_HVT DP_OP_424J2_126_3477_U699 ( .A(DP_OP_424J2_126_3477_n2542), .B(
        DP_OP_424J2_126_3477_n2454), .CI(DP_OP_424J2_126_3477_n2237), .CO(
        DP_OP_424J2_126_3477_n1203), .S(DP_OP_424J2_126_3477_n1204) );
  FADDX1_HVT DP_OP_424J2_126_3477_U698 ( .A(DP_OP_424J2_126_3477_n2850), .B(
        DP_OP_424J2_126_3477_n2806), .CI(DP_OP_424J2_126_3477_n2010), .CO(
        DP_OP_424J2_126_3477_n1201), .S(DP_OP_424J2_126_3477_n1202) );
  FADDX1_HVT DP_OP_424J2_126_3477_U697 ( .A(DP_OP_424J2_126_3477_n1885), .B(
        DP_OP_424J2_126_3477_n2281), .CI(DP_OP_424J2_126_3477_n2193), .CO(
        DP_OP_424J2_126_3477_n1199), .S(DP_OP_424J2_126_3477_n1200) );
  FADDX1_HVT DP_OP_424J2_126_3477_U696 ( .A(DP_OP_424J2_126_3477_n2105), .B(
        DP_OP_424J2_126_3477_n2667), .CI(DP_OP_424J2_126_3477_n1929), .CO(
        DP_OP_424J2_126_3477_n1197), .S(DP_OP_424J2_126_3477_n1198) );
  FADDX1_HVT DP_OP_424J2_126_3477_U695 ( .A(DP_OP_424J2_126_3477_n2491), .B(
        DP_OP_424J2_126_3477_n2894), .CI(DP_OP_424J2_126_3477_n2901), .CO(
        DP_OP_424J2_126_3477_n1195), .S(DP_OP_424J2_126_3477_n1196) );
  FADDX1_HVT DP_OP_424J2_126_3477_U694 ( .A(DP_OP_424J2_126_3477_n2359), .B(
        DP_OP_424J2_126_3477_n2244), .CI(DP_OP_424J2_126_3477_n2718), .CO(
        DP_OP_424J2_126_3477_n1193), .S(DP_OP_424J2_126_3477_n1194) );
  FADDX1_HVT DP_OP_424J2_126_3477_U693 ( .A(DP_OP_424J2_126_3477_n2674), .B(
        DP_OP_424J2_126_3477_n2318), .CI(DP_OP_424J2_126_3477_n2373), .CO(
        DP_OP_424J2_126_3477_n1191), .S(DP_OP_424J2_126_3477_n1192) );
  FADDX1_HVT DP_OP_424J2_126_3477_U692 ( .A(DP_OP_424J2_126_3477_n2054), .B(
        DP_OP_424J2_126_3477_n2623), .CI(DP_OP_424J2_126_3477_n2017), .CO(
        DP_OP_424J2_126_3477_n1189), .S(DP_OP_424J2_126_3477_n1190) );
  FADDX1_HVT DP_OP_424J2_126_3477_U691 ( .A(DP_OP_424J2_126_3477_n2799), .B(
        DP_OP_424J2_126_3477_n2403), .CI(DP_OP_424J2_126_3477_n2813), .CO(
        DP_OP_424J2_126_3477_n1187), .S(DP_OP_424J2_126_3477_n1188) );
  FADDX1_HVT DP_OP_424J2_126_3477_U690 ( .A(DP_OP_424J2_126_3477_n1973), .B(
        DP_OP_424J2_126_3477_n1922), .CI(DP_OP_424J2_126_3477_n2156), .CO(
        DP_OP_424J2_126_3477_n1185), .S(DP_OP_424J2_126_3477_n1186) );
  FADDX1_HVT DP_OP_424J2_126_3477_U689 ( .A(DP_OP_424J2_126_3477_n1878), .B(
        DP_OP_424J2_126_3477_n1834), .CI(DP_OP_424J2_126_3477_n2186), .CO(
        DP_OP_424J2_126_3477_n1183), .S(DP_OP_424J2_126_3477_n1184) );
  FADDX1_HVT DP_OP_424J2_126_3477_U688 ( .A(DP_OP_424J2_126_3477_n1250), .B(
        DP_OP_424J2_126_3477_n1425), .CI(DP_OP_424J2_126_3477_n1411), .CO(
        DP_OP_424J2_126_3477_n1181), .S(DP_OP_424J2_126_3477_n1182) );
  FADDX1_HVT DP_OP_424J2_126_3477_U687 ( .A(DP_OP_424J2_126_3477_n1423), .B(
        DP_OP_424J2_126_3477_n1413), .CI(DP_OP_424J2_126_3477_n1409), .CO(
        DP_OP_424J2_126_3477_n1179), .S(DP_OP_424J2_126_3477_n1180) );
  FADDX1_HVT DP_OP_424J2_126_3477_U686 ( .A(DP_OP_424J2_126_3477_n1421), .B(
        DP_OP_424J2_126_3477_n1415), .CI(DP_OP_424J2_126_3477_n1417), .CO(
        DP_OP_424J2_126_3477_n1177), .S(DP_OP_424J2_126_3477_n1178) );
  FADDX1_HVT DP_OP_424J2_126_3477_U685 ( .A(DP_OP_424J2_126_3477_n1419), .B(
        DP_OP_424J2_126_3477_n1407), .CI(DP_OP_424J2_126_3477_n1405), .CO(
        DP_OP_424J2_126_3477_n1175), .S(DP_OP_424J2_126_3477_n1176) );
  FADDX1_HVT DP_OP_424J2_126_3477_U684 ( .A(DP_OP_424J2_126_3477_n1403), .B(
        DP_OP_424J2_126_3477_n1383), .CI(DP_OP_424J2_126_3477_n1385), .CO(
        DP_OP_424J2_126_3477_n1173), .S(DP_OP_424J2_126_3477_n1174) );
  FADDX1_HVT DP_OP_424J2_126_3477_U683 ( .A(DP_OP_424J2_126_3477_n1401), .B(
        DP_OP_424J2_126_3477_n1399), .CI(DP_OP_424J2_126_3477_n1387), .CO(
        DP_OP_424J2_126_3477_n1171), .S(DP_OP_424J2_126_3477_n1172) );
  FADDX1_HVT DP_OP_424J2_126_3477_U682 ( .A(DP_OP_424J2_126_3477_n1397), .B(
        DP_OP_424J2_126_3477_n1389), .CI(DP_OP_424J2_126_3477_n1391), .CO(
        DP_OP_424J2_126_3477_n1169), .S(DP_OP_424J2_126_3477_n1170) );
  FADDX1_HVT DP_OP_424J2_126_3477_U681 ( .A(DP_OP_424J2_126_3477_n1395), .B(
        DP_OP_424J2_126_3477_n1393), .CI(DP_OP_424J2_126_3477_n1381), .CO(
        DP_OP_424J2_126_3477_n1167), .S(DP_OP_424J2_126_3477_n1168) );
  FADDX1_HVT DP_OP_424J2_126_3477_U680 ( .A(DP_OP_424J2_126_3477_n1379), .B(
        DP_OP_424J2_126_3477_n1365), .CI(DP_OP_424J2_126_3477_n1359), .CO(
        DP_OP_424J2_126_3477_n1165), .S(DP_OP_424J2_126_3477_n1166) );
  FADDX1_HVT DP_OP_424J2_126_3477_U679 ( .A(DP_OP_424J2_126_3477_n1377), .B(
        DP_OP_424J2_126_3477_n1248), .CI(DP_OP_424J2_126_3477_n1361), .CO(
        DP_OP_424J2_126_3477_n1163), .S(DP_OP_424J2_126_3477_n1164) );
  FADDX1_HVT DP_OP_424J2_126_3477_U678 ( .A(DP_OP_424J2_126_3477_n1373), .B(
        DP_OP_424J2_126_3477_n1242), .CI(DP_OP_424J2_126_3477_n1363), .CO(
        DP_OP_424J2_126_3477_n1161), .S(DP_OP_424J2_126_3477_n1162) );
  FADDX1_HVT DP_OP_424J2_126_3477_U677 ( .A(DP_OP_424J2_126_3477_n1371), .B(
        DP_OP_424J2_126_3477_n1238), .CI(DP_OP_424J2_126_3477_n1240), .CO(
        DP_OP_424J2_126_3477_n1159), .S(DP_OP_424J2_126_3477_n1160) );
  FADDX1_HVT DP_OP_424J2_126_3477_U676 ( .A(DP_OP_424J2_126_3477_n1375), .B(
        DP_OP_424J2_126_3477_n1236), .CI(DP_OP_424J2_126_3477_n1244), .CO(
        DP_OP_424J2_126_3477_n1157), .S(DP_OP_424J2_126_3477_n1158) );
  FADDX1_HVT DP_OP_424J2_126_3477_U675 ( .A(DP_OP_424J2_126_3477_n1369), .B(
        DP_OP_424J2_126_3477_n1367), .CI(DP_OP_424J2_126_3477_n1246), .CO(
        DP_OP_424J2_126_3477_n1155), .S(DP_OP_424J2_126_3477_n1156) );
  FADDX1_HVT DP_OP_424J2_126_3477_U674 ( .A(DP_OP_424J2_126_3477_n1234), .B(
        DP_OP_424J2_126_3477_n1224), .CI(DP_OP_424J2_126_3477_n1208), .CO(
        DP_OP_424J2_126_3477_n1153), .S(DP_OP_424J2_126_3477_n1154) );
  FADDX1_HVT DP_OP_424J2_126_3477_U673 ( .A(DP_OP_424J2_126_3477_n1226), .B(
        DP_OP_424J2_126_3477_n1212), .CI(DP_OP_424J2_126_3477_n1210), .CO(
        DP_OP_424J2_126_3477_n1151), .S(DP_OP_424J2_126_3477_n1152) );
  FADDX1_HVT DP_OP_424J2_126_3477_U672 ( .A(DP_OP_424J2_126_3477_n1222), .B(
        DP_OP_424J2_126_3477_n1216), .CI(DP_OP_424J2_126_3477_n1218), .CO(
        DP_OP_424J2_126_3477_n1149), .S(DP_OP_424J2_126_3477_n1150) );
  FADDX1_HVT DP_OP_424J2_126_3477_U671 ( .A(DP_OP_424J2_126_3477_n1214), .B(
        DP_OP_424J2_126_3477_n1232), .CI(DP_OP_424J2_126_3477_n1228), .CO(
        DP_OP_424J2_126_3477_n1147), .S(DP_OP_424J2_126_3477_n1148) );
  FADDX1_HVT DP_OP_424J2_126_3477_U670 ( .A(DP_OP_424J2_126_3477_n1230), .B(
        DP_OP_424J2_126_3477_n1220), .CI(DP_OP_424J2_126_3477_n1206), .CO(
        DP_OP_424J2_126_3477_n1145), .S(DP_OP_424J2_126_3477_n1146) );
  FADDX1_HVT DP_OP_424J2_126_3477_U669 ( .A(DP_OP_424J2_126_3477_n1204), .B(
        DP_OP_424J2_126_3477_n1190), .CI(DP_OP_424J2_126_3477_n1184), .CO(
        DP_OP_424J2_126_3477_n1143), .S(DP_OP_424J2_126_3477_n1144) );
  FADDX1_HVT DP_OP_424J2_126_3477_U668 ( .A(DP_OP_424J2_126_3477_n1202), .B(
        DP_OP_424J2_126_3477_n1192), .CI(DP_OP_424J2_126_3477_n1186), .CO(
        DP_OP_424J2_126_3477_n1141), .S(DP_OP_424J2_126_3477_n1142) );
  FADDX1_HVT DP_OP_424J2_126_3477_U667 ( .A(DP_OP_424J2_126_3477_n1198), .B(
        DP_OP_424J2_126_3477_n1194), .CI(DP_OP_424J2_126_3477_n1188), .CO(
        DP_OP_424J2_126_3477_n1139), .S(DP_OP_424J2_126_3477_n1140) );
  FADDX1_HVT DP_OP_424J2_126_3477_U666 ( .A(DP_OP_424J2_126_3477_n1200), .B(
        DP_OP_424J2_126_3477_n1196), .CI(DP_OP_424J2_126_3477_n1357), .CO(
        DP_OP_424J2_126_3477_n1137), .S(DP_OP_424J2_126_3477_n1138) );
  FADDX1_HVT DP_OP_424J2_126_3477_U665 ( .A(DP_OP_424J2_126_3477_n1355), .B(
        DP_OP_424J2_126_3477_n1353), .CI(DP_OP_424J2_126_3477_n1351), .CO(
        DP_OP_424J2_126_3477_n1135), .S(DP_OP_424J2_126_3477_n1136) );
  FADDX1_HVT DP_OP_424J2_126_3477_U664 ( .A(DP_OP_424J2_126_3477_n1349), .B(
        DP_OP_424J2_126_3477_n1345), .CI(DP_OP_424J2_126_3477_n1343), .CO(
        DP_OP_424J2_126_3477_n1133), .S(DP_OP_424J2_126_3477_n1134) );
  FADDX1_HVT DP_OP_424J2_126_3477_U663 ( .A(DP_OP_424J2_126_3477_n1347), .B(
        DP_OP_424J2_126_3477_n1182), .CI(DP_OP_424J2_126_3477_n1341), .CO(
        DP_OP_424J2_126_3477_n1131), .S(DP_OP_424J2_126_3477_n1132) );
  FADDX1_HVT DP_OP_424J2_126_3477_U662 ( .A(DP_OP_424J2_126_3477_n1339), .B(
        DP_OP_424J2_126_3477_n1180), .CI(DP_OP_424J2_126_3477_n1178), .CO(
        DP_OP_424J2_126_3477_n1129), .S(DP_OP_424J2_126_3477_n1130) );
  FADDX1_HVT DP_OP_424J2_126_3477_U661 ( .A(DP_OP_424J2_126_3477_n1337), .B(
        DP_OP_424J2_126_3477_n1333), .CI(DP_OP_424J2_126_3477_n1331), .CO(
        DP_OP_424J2_126_3477_n1127), .S(DP_OP_424J2_126_3477_n1128) );
  FADDX1_HVT DP_OP_424J2_126_3477_U660 ( .A(DP_OP_424J2_126_3477_n1335), .B(
        DP_OP_424J2_126_3477_n1176), .CI(DP_OP_424J2_126_3477_n1329), .CO(
        DP_OP_424J2_126_3477_n1125), .S(DP_OP_424J2_126_3477_n1126) );
  FADDX1_HVT DP_OP_424J2_126_3477_U659 ( .A(DP_OP_424J2_126_3477_n1323), .B(
        DP_OP_424J2_126_3477_n1170), .CI(DP_OP_424J2_126_3477_n1168), .CO(
        DP_OP_424J2_126_3477_n1123), .S(DP_OP_424J2_126_3477_n1124) );
  FADDX1_HVT DP_OP_424J2_126_3477_U658 ( .A(DP_OP_424J2_126_3477_n1327), .B(
        DP_OP_424J2_126_3477_n1325), .CI(DP_OP_424J2_126_3477_n1321), .CO(
        DP_OP_424J2_126_3477_n1121), .S(DP_OP_424J2_126_3477_n1122) );
  FADDX1_HVT DP_OP_424J2_126_3477_U657 ( .A(DP_OP_424J2_126_3477_n1174), .B(
        DP_OP_424J2_126_3477_n1172), .CI(DP_OP_424J2_126_3477_n1319), .CO(
        DP_OP_424J2_126_3477_n1119), .S(DP_OP_424J2_126_3477_n1120) );
  FADDX1_HVT DP_OP_424J2_126_3477_U656 ( .A(DP_OP_424J2_126_3477_n1166), .B(
        DP_OP_424J2_126_3477_n1160), .CI(DP_OP_424J2_126_3477_n1156), .CO(
        DP_OP_424J2_126_3477_n1117), .S(DP_OP_424J2_126_3477_n1118) );
  FADDX1_HVT DP_OP_424J2_126_3477_U655 ( .A(DP_OP_424J2_126_3477_n1317), .B(
        DP_OP_424J2_126_3477_n1158), .CI(DP_OP_424J2_126_3477_n1315), .CO(
        DP_OP_424J2_126_3477_n1115), .S(DP_OP_424J2_126_3477_n1116) );
  FADDX1_HVT DP_OP_424J2_126_3477_U654 ( .A(DP_OP_424J2_126_3477_n1164), .B(
        DP_OP_424J2_126_3477_n1162), .CI(DP_OP_424J2_126_3477_n1154), .CO(
        DP_OP_424J2_126_3477_n1113), .S(DP_OP_424J2_126_3477_n1114) );
  FADDX1_HVT DP_OP_424J2_126_3477_U653 ( .A(DP_OP_424J2_126_3477_n1148), .B(
        DP_OP_424J2_126_3477_n1313), .CI(DP_OP_424J2_126_3477_n1146), .CO(
        DP_OP_424J2_126_3477_n1111), .S(DP_OP_424J2_126_3477_n1112) );
  FADDX1_HVT DP_OP_424J2_126_3477_U652 ( .A(DP_OP_424J2_126_3477_n1152), .B(
        DP_OP_424J2_126_3477_n1150), .CI(DP_OP_424J2_126_3477_n1144), .CO(
        DP_OP_424J2_126_3477_n1109), .S(DP_OP_424J2_126_3477_n1110) );
  FADDX1_HVT DP_OP_424J2_126_3477_U651 ( .A(DP_OP_424J2_126_3477_n1142), .B(
        DP_OP_424J2_126_3477_n1311), .CI(DP_OP_424J2_126_3477_n1309), .CO(
        DP_OP_424J2_126_3477_n1107), .S(DP_OP_424J2_126_3477_n1108) );
  FADDX1_HVT DP_OP_424J2_126_3477_U650 ( .A(DP_OP_424J2_126_3477_n1140), .B(
        DP_OP_424J2_126_3477_n1138), .CI(DP_OP_424J2_126_3477_n1307), .CO(
        DP_OP_424J2_126_3477_n1105), .S(DP_OP_424J2_126_3477_n1106) );
  FADDX1_HVT DP_OP_424J2_126_3477_U649 ( .A(DP_OP_424J2_126_3477_n1305), .B(
        DP_OP_424J2_126_3477_n1136), .CI(DP_OP_424J2_126_3477_n1303), .CO(
        DP_OP_424J2_126_3477_n1103), .S(DP_OP_424J2_126_3477_n1104) );
  FADDX1_HVT DP_OP_424J2_126_3477_U648 ( .A(DP_OP_424J2_126_3477_n1301), .B(
        DP_OP_424J2_126_3477_n1134), .CI(DP_OP_424J2_126_3477_n1132), .CO(
        DP_OP_424J2_126_3477_n1101), .S(DP_OP_424J2_126_3477_n1102) );
  FADDX1_HVT DP_OP_424J2_126_3477_U647 ( .A(DP_OP_424J2_126_3477_n1299), .B(
        DP_OP_424J2_126_3477_n1297), .CI(DP_OP_424J2_126_3477_n1295), .CO(
        DP_OP_424J2_126_3477_n1099), .S(DP_OP_424J2_126_3477_n1100) );
  FADDX1_HVT DP_OP_424J2_126_3477_U646 ( .A(DP_OP_424J2_126_3477_n1293), .B(
        DP_OP_424J2_126_3477_n1128), .CI(DP_OP_424J2_126_3477_n1126), .CO(
        DP_OP_424J2_126_3477_n1097), .S(DP_OP_424J2_126_3477_n1098) );
  FADDX1_HVT DP_OP_424J2_126_3477_U645 ( .A(DP_OP_424J2_126_3477_n1291), .B(
        DP_OP_424J2_126_3477_n1130), .CI(DP_OP_424J2_126_3477_n1289), .CO(
        DP_OP_424J2_126_3477_n1095), .S(DP_OP_424J2_126_3477_n1096) );
  FADDX1_HVT DP_OP_424J2_126_3477_U644 ( .A(DP_OP_424J2_126_3477_n1287), .B(
        DP_OP_424J2_126_3477_n1124), .CI(DP_OP_424J2_126_3477_n1120), .CO(
        DP_OP_424J2_126_3477_n1093), .S(DP_OP_424J2_126_3477_n1094) );
  FADDX1_HVT DP_OP_424J2_126_3477_U643 ( .A(DP_OP_424J2_126_3477_n1122), .B(
        DP_OP_424J2_126_3477_n1118), .CI(DP_OP_424J2_126_3477_n1285), .CO(
        DP_OP_424J2_126_3477_n1091), .S(DP_OP_424J2_126_3477_n1092) );
  FADDX1_HVT DP_OP_424J2_126_3477_U642 ( .A(DP_OP_424J2_126_3477_n1116), .B(
        DP_OP_424J2_126_3477_n1114), .CI(DP_OP_424J2_126_3477_n1112), .CO(
        DP_OP_424J2_126_3477_n1089), .S(DP_OP_424J2_126_3477_n1090) );
  FADDX1_HVT DP_OP_424J2_126_3477_U641 ( .A(DP_OP_424J2_126_3477_n1283), .B(
        DP_OP_424J2_126_3477_n1110), .CI(DP_OP_424J2_126_3477_n1108), .CO(
        DP_OP_424J2_126_3477_n1087), .S(DP_OP_424J2_126_3477_n1088) );
  FADDX1_HVT DP_OP_424J2_126_3477_U640 ( .A(DP_OP_424J2_126_3477_n1281), .B(
        DP_OP_424J2_126_3477_n1106), .CI(DP_OP_424J2_126_3477_n1279), .CO(
        DP_OP_424J2_126_3477_n1085), .S(DP_OP_424J2_126_3477_n1086) );
  FADDX1_HVT DP_OP_424J2_126_3477_U639 ( .A(DP_OP_424J2_126_3477_n1277), .B(
        DP_OP_424J2_126_3477_n1104), .CI(DP_OP_424J2_126_3477_n1275), .CO(
        DP_OP_424J2_126_3477_n1083), .S(DP_OP_424J2_126_3477_n1084) );
  FADDX1_HVT DP_OP_424J2_126_3477_U638 ( .A(DP_OP_424J2_126_3477_n1273), .B(
        DP_OP_424J2_126_3477_n1102), .CI(DP_OP_424J2_126_3477_n1100), .CO(
        DP_OP_424J2_126_3477_n1081), .S(DP_OP_424J2_126_3477_n1082) );
  FADDX1_HVT DP_OP_424J2_126_3477_U637 ( .A(DP_OP_424J2_126_3477_n1271), .B(
        DP_OP_424J2_126_3477_n1098), .CI(DP_OP_424J2_126_3477_n1269), .CO(
        DP_OP_424J2_126_3477_n1079), .S(DP_OP_424J2_126_3477_n1080) );
  FADDX1_HVT DP_OP_424J2_126_3477_U636 ( .A(DP_OP_424J2_126_3477_n1096), .B(
        DP_OP_424J2_126_3477_n1094), .CI(DP_OP_424J2_126_3477_n1267), .CO(
        DP_OP_424J2_126_3477_n1077), .S(DP_OP_424J2_126_3477_n1078) );
  FADDX1_HVT DP_OP_424J2_126_3477_U635 ( .A(DP_OP_424J2_126_3477_n1092), .B(
        DP_OP_424J2_126_3477_n1090), .CI(DP_OP_424J2_126_3477_n1088), .CO(
        DP_OP_424J2_126_3477_n1075), .S(DP_OP_424J2_126_3477_n1076) );
  FADDX1_HVT DP_OP_424J2_126_3477_U634 ( .A(DP_OP_424J2_126_3477_n1265), .B(
        DP_OP_424J2_126_3477_n1086), .CI(DP_OP_424J2_126_3477_n1263), .CO(
        DP_OP_424J2_126_3477_n1073), .S(DP_OP_424J2_126_3477_n1074) );
  FADDX1_HVT DP_OP_424J2_126_3477_U633 ( .A(DP_OP_424J2_126_3477_n1084), .B(
        DP_OP_424J2_126_3477_n1261), .CI(DP_OP_424J2_126_3477_n1082), .CO(
        DP_OP_424J2_126_3477_n1071), .S(DP_OP_424J2_126_3477_n1072) );
  FADDX1_HVT DP_OP_424J2_126_3477_U632 ( .A(DP_OP_424J2_126_3477_n1259), .B(
        DP_OP_424J2_126_3477_n1080), .CI(DP_OP_424J2_126_3477_n1078), .CO(
        DP_OP_424J2_126_3477_n1069), .S(DP_OP_424J2_126_3477_n1070) );
  FADDX1_HVT DP_OP_424J2_126_3477_U631 ( .A(DP_OP_424J2_126_3477_n1257), .B(
        DP_OP_424J2_126_3477_n1076), .CI(DP_OP_424J2_126_3477_n1255), .CO(
        DP_OP_424J2_126_3477_n1067), .S(DP_OP_424J2_126_3477_n1068) );
  FADDX1_HVT DP_OP_424J2_126_3477_U630 ( .A(DP_OP_424J2_126_3477_n1074), .B(
        DP_OP_424J2_126_3477_n1072), .CI(DP_OP_424J2_126_3477_n1253), .CO(
        DP_OP_424J2_126_3477_n1065), .S(DP_OP_424J2_126_3477_n1066) );
  FADDX1_HVT DP_OP_424J2_126_3477_U629 ( .A(DP_OP_424J2_126_3477_n1070), .B(
        DP_OP_424J2_126_3477_n1251), .CI(DP_OP_424J2_126_3477_n1068), .CO(
        DP_OP_424J2_126_3477_n1063), .S(DP_OP_424J2_126_3477_n1064) );
  OR2X1_HVT DP_OP_424J2_126_3477_U628 ( .A1(DP_OP_424J2_126_3477_n2352), .A2(
        DP_OP_424J2_126_3477_n2002), .Y(DP_OP_424J2_126_3477_n1061) );
  FADDX1_HVT DP_OP_424J2_126_3477_U626 ( .A(DP_OP_424J2_126_3477_n2703), .B(
        DP_OP_424J2_126_3477_n1826), .CI(DP_OP_424J2_126_3477_n2395), .CO(
        DP_OP_424J2_126_3477_n1059), .S(DP_OP_424J2_126_3477_n1060) );
  FADDX1_HVT DP_OP_424J2_126_3477_U625 ( .A(DP_OP_424J2_126_3477_n2659), .B(
        DP_OP_424J2_126_3477_n2439), .CI(DP_OP_424J2_126_3477_n2747), .CO(
        DP_OP_424J2_126_3477_n1057), .S(DP_OP_424J2_126_3477_n1058) );
  FADDX1_HVT DP_OP_424J2_126_3477_U624 ( .A(DP_OP_424J2_126_3477_n2090), .B(
        DP_OP_424J2_126_3477_n2046), .CI(DP_OP_424J2_126_3477_n1958), .CO(
        DP_OP_424J2_126_3477_n1055), .S(DP_OP_424J2_126_3477_n1056) );
  FADDX1_HVT DP_OP_424J2_126_3477_U623 ( .A(DP_OP_424J2_126_3477_n2134), .B(
        DP_OP_424J2_126_3477_n2483), .CI(DP_OP_424J2_126_3477_n2178), .CO(
        DP_OP_424J2_126_3477_n1053), .S(DP_OP_424J2_126_3477_n1054) );
  FADDX1_HVT DP_OP_424J2_126_3477_U622 ( .A(DP_OP_424J2_126_3477_n1870), .B(
        DP_OP_424J2_126_3477_n2527), .CI(DP_OP_424J2_126_3477_n2571), .CO(
        DP_OP_424J2_126_3477_n1051), .S(DP_OP_424J2_126_3477_n1052) );
  FADDX1_HVT DP_OP_424J2_126_3477_U621 ( .A(DP_OP_424J2_126_3477_n2791), .B(
        DP_OP_424J2_126_3477_n2879), .CI(DP_OP_424J2_126_3477_n1914), .CO(
        DP_OP_424J2_126_3477_n1049), .S(DP_OP_424J2_126_3477_n1050) );
  FADDX1_HVT DP_OP_424J2_126_3477_U620 ( .A(DP_OP_424J2_126_3477_n2615), .B(
        DP_OP_424J2_126_3477_n2310), .CI(DP_OP_424J2_126_3477_n2266), .CO(
        DP_OP_424J2_126_3477_n1047), .S(DP_OP_424J2_126_3477_n1048) );
  FADDX1_HVT DP_OP_424J2_126_3477_U619 ( .A(DP_OP_424J2_126_3477_n2835), .B(
        DP_OP_424J2_126_3477_n2222), .CI(DP_OP_424J2_126_3477_n2636), .CO(
        DP_OP_424J2_126_3477_n1045), .S(DP_OP_424J2_126_3477_n1046) );
  FADDX1_HVT DP_OP_424J2_126_3477_U618 ( .A(DP_OP_424J2_126_3477_n2460), .B(
        DP_OP_424J2_126_3477_n2534), .CI(DP_OP_424J2_126_3477_n2287), .CO(
        DP_OP_424J2_126_3477_n1043), .S(DP_OP_424J2_126_3477_n1044) );
  FADDX1_HVT DP_OP_424J2_126_3477_U617 ( .A(DP_OP_424J2_126_3477_n2592), .B(
        DP_OP_424J2_126_3477_n1965), .CI(DP_OP_424J2_126_3477_n2273), .CO(
        DP_OP_424J2_126_3477_n1041), .S(DP_OP_424J2_126_3477_n1042) );
  FADDX1_HVT DP_OP_424J2_126_3477_U616 ( .A(DP_OP_424J2_126_3477_n2331), .B(
        DP_OP_424J2_126_3477_n2409), .CI(DP_OP_424J2_126_3477_n2141), .CO(
        DP_OP_424J2_126_3477_n1039), .S(DP_OP_424J2_126_3477_n1040) );
  FADDX1_HVT DP_OP_424J2_126_3477_U615 ( .A(DP_OP_424J2_126_3477_n2111), .B(
        DP_OP_424J2_126_3477_n2724), .CI(DP_OP_424J2_126_3477_n2067), .CO(
        DP_OP_424J2_126_3477_n1037), .S(DP_OP_424J2_126_3477_n1038) );
  FADDX1_HVT DP_OP_424J2_126_3477_U614 ( .A(DP_OP_424J2_126_3477_n2199), .B(
        DP_OP_424J2_126_3477_n2148), .CI(DP_OP_424J2_126_3477_n2504), .CO(
        DP_OP_424J2_126_3477_n1035), .S(DP_OP_424J2_126_3477_n1036) );
  FADDX1_HVT DP_OP_424J2_126_3477_U613 ( .A(DP_OP_424J2_126_3477_n2416), .B(
        DP_OP_424J2_126_3477_n1782), .CI(DP_OP_424J2_126_3477_n2856), .CO(
        DP_OP_424J2_126_3477_n1033), .S(DP_OP_424J2_126_3477_n1034) );
  FADDX1_HVT DP_OP_424J2_126_3477_U612 ( .A(DP_OP_424J2_126_3477_n2548), .B(
        DP_OP_424J2_126_3477_n2324), .CI(DP_OP_424J2_126_3477_n1891), .CO(
        DP_OP_424J2_126_3477_n1031), .S(DP_OP_424J2_126_3477_n1032) );
  FADDX1_HVT DP_OP_424J2_126_3477_U611 ( .A(DP_OP_424J2_126_3477_n1847), .B(
        DP_OP_424J2_126_3477_n1840), .CI(DP_OP_424J2_126_3477_n2229), .CO(
        DP_OP_424J2_126_3477_n1029), .S(DP_OP_424J2_126_3477_n1030) );
  FADDX1_HVT DP_OP_424J2_126_3477_U610 ( .A(DP_OP_424J2_126_3477_n2842), .B(
        DP_OP_424J2_126_3477_n2629), .CI(DP_OP_424J2_126_3477_n2446), .CO(
        DP_OP_424J2_126_3477_n1027), .S(DP_OP_424J2_126_3477_n1028) );
  FADDX1_HVT DP_OP_424J2_126_3477_U609 ( .A(DP_OP_424J2_126_3477_n2886), .B(
        DP_OP_424J2_126_3477_n2585), .CI(DP_OP_424J2_126_3477_n2097), .CO(
        DP_OP_424J2_126_3477_n1025), .S(DP_OP_424J2_126_3477_n1026) );
  FADDX1_HVT DP_OP_424J2_126_3477_U608 ( .A(DP_OP_424J2_126_3477_n2754), .B(
        DP_OP_424J2_126_3477_n2023), .CI(DP_OP_424J2_126_3477_n2768), .CO(
        DP_OP_424J2_126_3477_n1023), .S(DP_OP_424J2_126_3477_n1024) );
  FADDX1_HVT DP_OP_424J2_126_3477_U607 ( .A(DP_OP_424J2_126_3477_n2060), .B(
        DP_OP_424J2_126_3477_n2497), .CI(DP_OP_424J2_126_3477_n2578), .CO(
        DP_OP_424J2_126_3477_n1021), .S(DP_OP_424J2_126_3477_n1022) );
  FADDX1_HVT DP_OP_424J2_126_3477_U606 ( .A(DP_OP_424J2_126_3477_n2680), .B(
        DP_OP_424J2_126_3477_n1979), .CI(DP_OP_424J2_126_3477_n1935), .CO(
        DP_OP_424J2_126_3477_n1019), .S(DP_OP_424J2_126_3477_n1020) );
  FADDX1_HVT DP_OP_424J2_126_3477_U605 ( .A(DP_OP_424J2_126_3477_n2710), .B(
        DP_OP_424J2_126_3477_n2761), .CI(DP_OP_424J2_126_3477_n2365), .CO(
        DP_OP_424J2_126_3477_n1017), .S(DP_OP_424J2_126_3477_n1018) );
  FADDX1_HVT DP_OP_424J2_126_3477_U604 ( .A(DP_OP_424J2_126_3477_n2541), .B(
        DP_OP_424J2_126_3477_n2453), .CI(DP_OP_424J2_126_3477_n2236), .CO(
        DP_OP_424J2_126_3477_n1015), .S(DP_OP_424J2_126_3477_n1016) );
  FADDX1_HVT DP_OP_424J2_126_3477_U603 ( .A(DP_OP_424J2_126_3477_n2849), .B(
        DP_OP_424J2_126_3477_n2805), .CI(DP_OP_424J2_126_3477_n2009), .CO(
        DP_OP_424J2_126_3477_n1013), .S(DP_OP_424J2_126_3477_n1014) );
  FADDX1_HVT DP_OP_424J2_126_3477_U602 ( .A(DP_OP_424J2_126_3477_n1884), .B(
        DP_OP_424J2_126_3477_n2280), .CI(DP_OP_424J2_126_3477_n2192), .CO(
        DP_OP_424J2_126_3477_n1011), .S(DP_OP_424J2_126_3477_n1012) );
  FADDX1_HVT DP_OP_424J2_126_3477_U601 ( .A(DP_OP_424J2_126_3477_n2104), .B(
        DP_OP_424J2_126_3477_n2666), .CI(DP_OP_424J2_126_3477_n1928), .CO(
        DP_OP_424J2_126_3477_n1009), .S(DP_OP_424J2_126_3477_n1010) );
  FADDX1_HVT DP_OP_424J2_126_3477_U600 ( .A(DP_OP_424J2_126_3477_n2490), .B(
        DP_OP_424J2_126_3477_n2893), .CI(DP_OP_424J2_126_3477_n2900), .CO(
        DP_OP_424J2_126_3477_n1007), .S(DP_OP_424J2_126_3477_n1008) );
  FADDX1_HVT DP_OP_424J2_126_3477_U599 ( .A(DP_OP_424J2_126_3477_n2358), .B(
        DP_OP_424J2_126_3477_n2243), .CI(DP_OP_424J2_126_3477_n2717), .CO(
        DP_OP_424J2_126_3477_n1005), .S(DP_OP_424J2_126_3477_n1006) );
  FADDX1_HVT DP_OP_424J2_126_3477_U598 ( .A(DP_OP_424J2_126_3477_n2673), .B(
        DP_OP_424J2_126_3477_n2317), .CI(DP_OP_424J2_126_3477_n2372), .CO(
        DP_OP_424J2_126_3477_n1003), .S(DP_OP_424J2_126_3477_n1004) );
  FADDX1_HVT DP_OP_424J2_126_3477_U597 ( .A(DP_OP_424J2_126_3477_n2053), .B(
        DP_OP_424J2_126_3477_n2622), .CI(DP_OP_424J2_126_3477_n2016), .CO(
        DP_OP_424J2_126_3477_n1001), .S(DP_OP_424J2_126_3477_n1002) );
  FADDX1_HVT DP_OP_424J2_126_3477_U596 ( .A(DP_OP_424J2_126_3477_n2798), .B(
        DP_OP_424J2_126_3477_n2402), .CI(DP_OP_424J2_126_3477_n1249), .CO(
        DP_OP_424J2_126_3477_n999), .S(DP_OP_424J2_126_3477_n1000) );
  FADDX1_HVT DP_OP_424J2_126_3477_U595 ( .A(DP_OP_424J2_126_3477_n1972), .B(
        DP_OP_424J2_126_3477_n2155), .CI(DP_OP_424J2_126_3477_n2812), .CO(
        DP_OP_424J2_126_3477_n997), .S(DP_OP_424J2_126_3477_n998) );
  FADDX1_HVT DP_OP_424J2_126_3477_U594 ( .A(DP_OP_424J2_126_3477_n1877), .B(
        DP_OP_424J2_126_3477_n1921), .CI(DP_OP_424J2_126_3477_n2185), .CO(
        DP_OP_424J2_126_3477_n995), .S(DP_OP_424J2_126_3477_n996) );
  FADDX1_HVT DP_OP_424J2_126_3477_U593 ( .A(DP_OP_424J2_126_3477_n1833), .B(
        DP_OP_424J2_126_3477_n1247), .CI(DP_OP_424J2_126_3477_n1245), .CO(
        DP_OP_424J2_126_3477_n993), .S(DP_OP_424J2_126_3477_n994) );
  FADDX1_HVT DP_OP_424J2_126_3477_U592 ( .A(DP_OP_424J2_126_3477_n1243), .B(
        DP_OP_424J2_126_3477_n1062), .CI(DP_OP_424J2_126_3477_n1233), .CO(
        DP_OP_424J2_126_3477_n991), .S(DP_OP_424J2_126_3477_n992) );
  FADDX1_HVT DP_OP_424J2_126_3477_U591 ( .A(DP_OP_424J2_126_3477_n1241), .B(
        DP_OP_424J2_126_3477_n1235), .CI(DP_OP_424J2_126_3477_n1237), .CO(
        DP_OP_424J2_126_3477_n989), .S(DP_OP_424J2_126_3477_n990) );
  FADDX1_HVT DP_OP_424J2_126_3477_U590 ( .A(DP_OP_424J2_126_3477_n1239), .B(
        DP_OP_424J2_126_3477_n1231), .CI(DP_OP_424J2_126_3477_n1229), .CO(
        DP_OP_424J2_126_3477_n987), .S(DP_OP_424J2_126_3477_n988) );
  FADDX1_HVT DP_OP_424J2_126_3477_U589 ( .A(DP_OP_424J2_126_3477_n1227), .B(
        DP_OP_424J2_126_3477_n1207), .CI(DP_OP_424J2_126_3477_n1209), .CO(
        DP_OP_424J2_126_3477_n985), .S(DP_OP_424J2_126_3477_n986) );
  FADDX1_HVT DP_OP_424J2_126_3477_U588 ( .A(DP_OP_424J2_126_3477_n1225), .B(
        DP_OP_424J2_126_3477_n1213), .CI(DP_OP_424J2_126_3477_n1211), .CO(
        DP_OP_424J2_126_3477_n983), .S(DP_OP_424J2_126_3477_n984) );
  FADDX1_HVT DP_OP_424J2_126_3477_U587 ( .A(DP_OP_424J2_126_3477_n1217), .B(
        DP_OP_424J2_126_3477_n1215), .CI(DP_OP_424J2_126_3477_n1223), .CO(
        DP_OP_424J2_126_3477_n981), .S(DP_OP_424J2_126_3477_n982) );
  FADDX1_HVT DP_OP_424J2_126_3477_U586 ( .A(DP_OP_424J2_126_3477_n1219), .B(
        DP_OP_424J2_126_3477_n1221), .CI(DP_OP_424J2_126_3477_n1203), .CO(
        DP_OP_424J2_126_3477_n979), .S(DP_OP_424J2_126_3477_n980) );
  FADDX1_HVT DP_OP_424J2_126_3477_U585 ( .A(DP_OP_424J2_126_3477_n1205), .B(
        DP_OP_424J2_126_3477_n1189), .CI(DP_OP_424J2_126_3477_n1183), .CO(
        DP_OP_424J2_126_3477_n977), .S(DP_OP_424J2_126_3477_n978) );
  FADDX1_HVT DP_OP_424J2_126_3477_U584 ( .A(DP_OP_424J2_126_3477_n1201), .B(
        DP_OP_424J2_126_3477_n1060), .CI(DP_OP_424J2_126_3477_n1187), .CO(
        DP_OP_424J2_126_3477_n975), .S(DP_OP_424J2_126_3477_n976) );
  FADDX1_HVT DP_OP_424J2_126_3477_U583 ( .A(DP_OP_424J2_126_3477_n1197), .B(
        DP_OP_424J2_126_3477_n1054), .CI(DP_OP_424J2_126_3477_n1185), .CO(
        DP_OP_424J2_126_3477_n973), .S(DP_OP_424J2_126_3477_n974) );
  FADDX1_HVT DP_OP_424J2_126_3477_U582 ( .A(DP_OP_424J2_126_3477_n1199), .B(
        DP_OP_424J2_126_3477_n1050), .CI(DP_OP_424J2_126_3477_n1052), .CO(
        DP_OP_424J2_126_3477_n971), .S(DP_OP_424J2_126_3477_n972) );
  FADDX1_HVT DP_OP_424J2_126_3477_U581 ( .A(DP_OP_424J2_126_3477_n1195), .B(
        DP_OP_424J2_126_3477_n1048), .CI(DP_OP_424J2_126_3477_n1058), .CO(
        DP_OP_424J2_126_3477_n969), .S(DP_OP_424J2_126_3477_n970) );
  FADDX1_HVT DP_OP_424J2_126_3477_U580 ( .A(DP_OP_424J2_126_3477_n1193), .B(
        DP_OP_424J2_126_3477_n1191), .CI(DP_OP_424J2_126_3477_n1056), .CO(
        DP_OP_424J2_126_3477_n967), .S(DP_OP_424J2_126_3477_n968) );
  FADDX1_HVT DP_OP_424J2_126_3477_U579 ( .A(DP_OP_424J2_126_3477_n1046), .B(
        DP_OP_424J2_126_3477_n1038), .CI(DP_OP_424J2_126_3477_n1020), .CO(
        DP_OP_424J2_126_3477_n965), .S(DP_OP_424J2_126_3477_n966) );
  FADDX1_HVT DP_OP_424J2_126_3477_U578 ( .A(DP_OP_424J2_126_3477_n1034), .B(
        DP_OP_424J2_126_3477_n1024), .CI(DP_OP_424J2_126_3477_n1022), .CO(
        DP_OP_424J2_126_3477_n963), .S(DP_OP_424J2_126_3477_n964) );
  FADDX1_HVT DP_OP_424J2_126_3477_U577 ( .A(DP_OP_424J2_126_3477_n1036), .B(
        DP_OP_424J2_126_3477_n1028), .CI(DP_OP_424J2_126_3477_n1030), .CO(
        DP_OP_424J2_126_3477_n961), .S(DP_OP_424J2_126_3477_n962) );
  FADDX1_HVT DP_OP_424J2_126_3477_U576 ( .A(DP_OP_424J2_126_3477_n1026), .B(
        DP_OP_424J2_126_3477_n1044), .CI(DP_OP_424J2_126_3477_n1042), .CO(
        DP_OP_424J2_126_3477_n959), .S(DP_OP_424J2_126_3477_n960) );
  FADDX1_HVT DP_OP_424J2_126_3477_U575 ( .A(DP_OP_424J2_126_3477_n1040), .B(
        DP_OP_424J2_126_3477_n1032), .CI(DP_OP_424J2_126_3477_n1018), .CO(
        DP_OP_424J2_126_3477_n957), .S(DP_OP_424J2_126_3477_n958) );
  FADDX1_HVT DP_OP_424J2_126_3477_U574 ( .A(DP_OP_424J2_126_3477_n1016), .B(
        DP_OP_424J2_126_3477_n1002), .CI(DP_OP_424J2_126_3477_n996), .CO(
        DP_OP_424J2_126_3477_n955), .S(DP_OP_424J2_126_3477_n956) );
  FADDX1_HVT DP_OP_424J2_126_3477_U573 ( .A(DP_OP_424J2_126_3477_n1014), .B(
        DP_OP_424J2_126_3477_n1004), .CI(DP_OP_424J2_126_3477_n998), .CO(
        DP_OP_424J2_126_3477_n953), .S(DP_OP_424J2_126_3477_n954) );
  FADDX1_HVT DP_OP_424J2_126_3477_U572 ( .A(DP_OP_424J2_126_3477_n1010), .B(
        DP_OP_424J2_126_3477_n1006), .CI(DP_OP_424J2_126_3477_n1181), .CO(
        DP_OP_424J2_126_3477_n951), .S(DP_OP_424J2_126_3477_n952) );
  FADDX1_HVT DP_OP_424J2_126_3477_U571 ( .A(DP_OP_424J2_126_3477_n1008), .B(
        DP_OP_424J2_126_3477_n1012), .CI(DP_OP_424J2_126_3477_n1000), .CO(
        DP_OP_424J2_126_3477_n949), .S(DP_OP_424J2_126_3477_n950) );
  FADDX1_HVT DP_OP_424J2_126_3477_U570 ( .A(DP_OP_424J2_126_3477_n1179), .B(
        DP_OP_424J2_126_3477_n1177), .CI(DP_OP_424J2_126_3477_n1175), .CO(
        DP_OP_424J2_126_3477_n947), .S(DP_OP_424J2_126_3477_n948) );
  FADDX1_HVT DP_OP_424J2_126_3477_U569 ( .A(DP_OP_424J2_126_3477_n1173), .B(
        DP_OP_424J2_126_3477_n1167), .CI(DP_OP_424J2_126_3477_n1169), .CO(
        DP_OP_424J2_126_3477_n945), .S(DP_OP_424J2_126_3477_n946) );
  FADDX1_HVT DP_OP_424J2_126_3477_U568 ( .A(DP_OP_424J2_126_3477_n1171), .B(
        DP_OP_424J2_126_3477_n1165), .CI(DP_OP_424J2_126_3477_n994), .CO(
        DP_OP_424J2_126_3477_n943), .S(DP_OP_424J2_126_3477_n944) );
  FADDX1_HVT DP_OP_424J2_126_3477_U567 ( .A(DP_OP_424J2_126_3477_n1163), .B(
        DP_OP_424J2_126_3477_n1155), .CI(DP_OP_424J2_126_3477_n992), .CO(
        DP_OP_424J2_126_3477_n941), .S(DP_OP_424J2_126_3477_n942) );
  FADDX1_HVT DP_OP_424J2_126_3477_U566 ( .A(DP_OP_424J2_126_3477_n1161), .B(
        DP_OP_424J2_126_3477_n1157), .CI(DP_OP_424J2_126_3477_n990), .CO(
        DP_OP_424J2_126_3477_n939), .S(DP_OP_424J2_126_3477_n940) );
  FADDX1_HVT DP_OP_424J2_126_3477_U565 ( .A(DP_OP_424J2_126_3477_n1159), .B(
        DP_OP_424J2_126_3477_n1153), .CI(DP_OP_424J2_126_3477_n988), .CO(
        DP_OP_424J2_126_3477_n937), .S(DP_OP_424J2_126_3477_n938) );
  FADDX1_HVT DP_OP_424J2_126_3477_U564 ( .A(DP_OP_424J2_126_3477_n1151), .B(
        DP_OP_424J2_126_3477_n984), .CI(DP_OP_424J2_126_3477_n980), .CO(
        DP_OP_424J2_126_3477_n935), .S(DP_OP_424J2_126_3477_n936) );
  FADDX1_HVT DP_OP_424J2_126_3477_U563 ( .A(DP_OP_424J2_126_3477_n1145), .B(
        DP_OP_424J2_126_3477_n982), .CI(DP_OP_424J2_126_3477_n986), .CO(
        DP_OP_424J2_126_3477_n933), .S(DP_OP_424J2_126_3477_n934) );
  FADDX1_HVT DP_OP_424J2_126_3477_U562 ( .A(DP_OP_424J2_126_3477_n1149), .B(
        DP_OP_424J2_126_3477_n1147), .CI(DP_OP_424J2_126_3477_n1143), .CO(
        DP_OP_424J2_126_3477_n931), .S(DP_OP_424J2_126_3477_n932) );
  FADDX1_HVT DP_OP_424J2_126_3477_U561 ( .A(DP_OP_424J2_126_3477_n978), .B(
        DP_OP_424J2_126_3477_n968), .CI(DP_OP_424J2_126_3477_n1137), .CO(
        DP_OP_424J2_126_3477_n929), .S(DP_OP_424J2_126_3477_n930) );
  FADDX1_HVT DP_OP_424J2_126_3477_U560 ( .A(DP_OP_424J2_126_3477_n1141), .B(
        DP_OP_424J2_126_3477_n972), .CI(DP_OP_424J2_126_3477_n974), .CO(
        DP_OP_424J2_126_3477_n927), .S(DP_OP_424J2_126_3477_n928) );
  FADDX1_HVT DP_OP_424J2_126_3477_U559 ( .A(DP_OP_424J2_126_3477_n976), .B(
        DP_OP_424J2_126_3477_n970), .CI(DP_OP_424J2_126_3477_n1139), .CO(
        DP_OP_424J2_126_3477_n925), .S(DP_OP_424J2_126_3477_n926) );
  FADDX1_HVT DP_OP_424J2_126_3477_U558 ( .A(DP_OP_424J2_126_3477_n966), .B(
        DP_OP_424J2_126_3477_n960), .CI(DP_OP_424J2_126_3477_n958), .CO(
        DP_OP_424J2_126_3477_n923), .S(DP_OP_424J2_126_3477_n924) );
  FADDX1_HVT DP_OP_424J2_126_3477_U557 ( .A(DP_OP_424J2_126_3477_n962), .B(
        DP_OP_424J2_126_3477_n964), .CI(DP_OP_424J2_126_3477_n1135), .CO(
        DP_OP_424J2_126_3477_n921), .S(DP_OP_424J2_126_3477_n922) );
  FADDX1_HVT DP_OP_424J2_126_3477_U556 ( .A(DP_OP_424J2_126_3477_n956), .B(
        DP_OP_424J2_126_3477_n1133), .CI(DP_OP_424J2_126_3477_n1131), .CO(
        DP_OP_424J2_126_3477_n919), .S(DP_OP_424J2_126_3477_n920) );
  FADDX1_HVT DP_OP_424J2_126_3477_U555 ( .A(DP_OP_424J2_126_3477_n954), .B(
        DP_OP_424J2_126_3477_n952), .CI(DP_OP_424J2_126_3477_n950), .CO(
        DP_OP_424J2_126_3477_n917), .S(DP_OP_424J2_126_3477_n918) );
  FADDX1_HVT DP_OP_424J2_126_3477_U554 ( .A(DP_OP_424J2_126_3477_n1129), .B(
        DP_OP_424J2_126_3477_n948), .CI(DP_OP_424J2_126_3477_n1125), .CO(
        DP_OP_424J2_126_3477_n915), .S(DP_OP_424J2_126_3477_n916) );
  FADDX1_HVT DP_OP_424J2_126_3477_U553 ( .A(DP_OP_424J2_126_3477_n1127), .B(
        DP_OP_424J2_126_3477_n1123), .CI(DP_OP_424J2_126_3477_n1121), .CO(
        DP_OP_424J2_126_3477_n913), .S(DP_OP_424J2_126_3477_n914) );
  FADDX1_HVT DP_OP_424J2_126_3477_U552 ( .A(DP_OP_424J2_126_3477_n1119), .B(
        DP_OP_424J2_126_3477_n946), .CI(DP_OP_424J2_126_3477_n944), .CO(
        DP_OP_424J2_126_3477_n911), .S(DP_OP_424J2_126_3477_n912) );
  FADDX1_HVT DP_OP_424J2_126_3477_U551 ( .A(DP_OP_424J2_126_3477_n1117), .B(
        DP_OP_424J2_126_3477_n940), .CI(DP_OP_424J2_126_3477_n938), .CO(
        DP_OP_424J2_126_3477_n909), .S(DP_OP_424J2_126_3477_n910) );
  FADDX1_HVT DP_OP_424J2_126_3477_U550 ( .A(DP_OP_424J2_126_3477_n1115), .B(
        DP_OP_424J2_126_3477_n942), .CI(DP_OP_424J2_126_3477_n1113), .CO(
        DP_OP_424J2_126_3477_n907), .S(DP_OP_424J2_126_3477_n908) );
  FADDX1_HVT DP_OP_424J2_126_3477_U549 ( .A(DP_OP_424J2_126_3477_n1109), .B(
        DP_OP_424J2_126_3477_n936), .CI(DP_OP_424J2_126_3477_n932), .CO(
        DP_OP_424J2_126_3477_n905), .S(DP_OP_424J2_126_3477_n906) );
  FADDX1_HVT DP_OP_424J2_126_3477_U548 ( .A(DP_OP_424J2_126_3477_n1111), .B(
        DP_OP_424J2_126_3477_n934), .CI(DP_OP_424J2_126_3477_n930), .CO(
        DP_OP_424J2_126_3477_n903), .S(DP_OP_424J2_126_3477_n904) );
  FADDX1_HVT DP_OP_424J2_126_3477_U547 ( .A(DP_OP_424J2_126_3477_n1107), .B(
        DP_OP_424J2_126_3477_n926), .CI(DP_OP_424J2_126_3477_n1105), .CO(
        DP_OP_424J2_126_3477_n901), .S(DP_OP_424J2_126_3477_n902) );
  FADDX1_HVT DP_OP_424J2_126_3477_U546 ( .A(DP_OP_424J2_126_3477_n928), .B(
        DP_OP_424J2_126_3477_n924), .CI(DP_OP_424J2_126_3477_n1103), .CO(
        DP_OP_424J2_126_3477_n899), .S(DP_OP_424J2_126_3477_n900) );
  FADDX1_HVT DP_OP_424J2_126_3477_U545 ( .A(DP_OP_424J2_126_3477_n922), .B(
        DP_OP_424J2_126_3477_n920), .CI(DP_OP_424J2_126_3477_n918), .CO(
        DP_OP_424J2_126_3477_n897), .S(DP_OP_424J2_126_3477_n898) );
  FADDX1_HVT DP_OP_424J2_126_3477_U544 ( .A(DP_OP_424J2_126_3477_n1101), .B(
        DP_OP_424J2_126_3477_n1099), .CI(DP_OP_424J2_126_3477_n1097), .CO(
        DP_OP_424J2_126_3477_n895), .S(DP_OP_424J2_126_3477_n896) );
  FADDX1_HVT DP_OP_424J2_126_3477_U543 ( .A(DP_OP_424J2_126_3477_n916), .B(
        DP_OP_424J2_126_3477_n1095), .CI(DP_OP_424J2_126_3477_n914), .CO(
        DP_OP_424J2_126_3477_n893), .S(DP_OP_424J2_126_3477_n894) );
  FADDX1_HVT DP_OP_424J2_126_3477_U542 ( .A(DP_OP_424J2_126_3477_n1093), .B(
        DP_OP_424J2_126_3477_n912), .CI(DP_OP_424J2_126_3477_n1091), .CO(
        DP_OP_424J2_126_3477_n891), .S(DP_OP_424J2_126_3477_n892) );
  FADDX1_HVT DP_OP_424J2_126_3477_U541 ( .A(DP_OP_424J2_126_3477_n910), .B(
        DP_OP_424J2_126_3477_n908), .CI(DP_OP_424J2_126_3477_n1089), .CO(
        DP_OP_424J2_126_3477_n889), .S(DP_OP_424J2_126_3477_n890) );
  FADDX1_HVT DP_OP_424J2_126_3477_U540 ( .A(DP_OP_424J2_126_3477_n906), .B(
        DP_OP_424J2_126_3477_n1087), .CI(DP_OP_424J2_126_3477_n904), .CO(
        DP_OP_424J2_126_3477_n887), .S(DP_OP_424J2_126_3477_n888) );
  FADDX1_HVT DP_OP_424J2_126_3477_U539 ( .A(DP_OP_424J2_126_3477_n902), .B(
        DP_OP_424J2_126_3477_n1085), .CI(DP_OP_424J2_126_3477_n900), .CO(
        DP_OP_424J2_126_3477_n885), .S(DP_OP_424J2_126_3477_n886) );
  FADDX1_HVT DP_OP_424J2_126_3477_U538 ( .A(DP_OP_424J2_126_3477_n1083), .B(
        DP_OP_424J2_126_3477_n898), .CI(DP_OP_424J2_126_3477_n1081), .CO(
        DP_OP_424J2_126_3477_n883), .S(DP_OP_424J2_126_3477_n884) );
  FADDX1_HVT DP_OP_424J2_126_3477_U537 ( .A(DP_OP_424J2_126_3477_n896), .B(
        DP_OP_424J2_126_3477_n1079), .CI(DP_OP_424J2_126_3477_n894), .CO(
        DP_OP_424J2_126_3477_n881), .S(DP_OP_424J2_126_3477_n882) );
  FADDX1_HVT DP_OP_424J2_126_3477_U536 ( .A(DP_OP_424J2_126_3477_n1077), .B(
        DP_OP_424J2_126_3477_n892), .CI(DP_OP_424J2_126_3477_n890), .CO(
        DP_OP_424J2_126_3477_n879), .S(DP_OP_424J2_126_3477_n880) );
  FADDX1_HVT DP_OP_424J2_126_3477_U535 ( .A(DP_OP_424J2_126_3477_n1075), .B(
        DP_OP_424J2_126_3477_n888), .CI(DP_OP_424J2_126_3477_n1073), .CO(
        DP_OP_424J2_126_3477_n877), .S(DP_OP_424J2_126_3477_n878) );
  FADDX1_HVT DP_OP_424J2_126_3477_U534 ( .A(DP_OP_424J2_126_3477_n886), .B(
        DP_OP_424J2_126_3477_n1071), .CI(DP_OP_424J2_126_3477_n884), .CO(
        DP_OP_424J2_126_3477_n875), .S(DP_OP_424J2_126_3477_n876) );
  FADDX1_HVT DP_OP_424J2_126_3477_U533 ( .A(DP_OP_424J2_126_3477_n882), .B(
        DP_OP_424J2_126_3477_n1069), .CI(DP_OP_424J2_126_3477_n880), .CO(
        DP_OP_424J2_126_3477_n873), .S(DP_OP_424J2_126_3477_n874) );
  FADDX1_HVT DP_OP_424J2_126_3477_U532 ( .A(DP_OP_424J2_126_3477_n1067), .B(
        DP_OP_424J2_126_3477_n878), .CI(DP_OP_424J2_126_3477_n876), .CO(
        DP_OP_424J2_126_3477_n871), .S(DP_OP_424J2_126_3477_n872) );
  FADDX1_HVT DP_OP_424J2_126_3477_U531 ( .A(DP_OP_424J2_126_3477_n1065), .B(
        DP_OP_424J2_126_3477_n874), .CI(DP_OP_424J2_126_3477_n1063), .CO(
        DP_OP_424J2_126_3477_n869), .S(DP_OP_424J2_126_3477_n870) );
  FADDX1_HVT DP_OP_424J2_126_3477_U530 ( .A(DP_OP_424J2_126_3477_n2351), .B(
        DP_OP_424J2_126_3477_n2723), .CI(DP_OP_424J2_126_3477_n2394), .CO(
        DP_OP_424J2_126_3477_n867), .S(DP_OP_424J2_126_3477_n868) );
  FADDX1_HVT DP_OP_424J2_126_3477_U529 ( .A(DP_OP_424J2_126_3477_n2001), .B(
        DP_OP_424J2_126_3477_n1825), .CI(DP_OP_424J2_126_3477_n2503), .CO(
        DP_OP_424J2_126_3477_n865), .S(DP_OP_424J2_126_3477_n866) );
  FADDX1_HVT DP_OP_424J2_126_3477_U528 ( .A(DP_OP_424J2_126_3477_n2702), .B(
        DP_OP_424J2_126_3477_n1913), .CI(DP_OP_424J2_126_3477_n1890), .CO(
        DP_OP_424J2_126_3477_n863), .S(DP_OP_424J2_126_3477_n864) );
  FADDX1_HVT DP_OP_424J2_126_3477_U527 ( .A(DP_OP_424J2_126_3477_n2089), .B(
        DP_OP_424J2_126_3477_n2526), .CI(DP_OP_424J2_126_3477_n2855), .CO(
        DP_OP_424J2_126_3477_n861), .S(DP_OP_424J2_126_3477_n862) );
  FADDX1_HVT DP_OP_424J2_126_3477_U526 ( .A(DP_OP_424J2_126_3477_n1869), .B(
        DP_OP_424J2_126_3477_n2045), .CI(DP_OP_424J2_126_3477_n2767), .CO(
        DP_OP_424J2_126_3477_n859), .S(DP_OP_424J2_126_3477_n860) );
  FADDX1_HVT DP_OP_424J2_126_3477_U525 ( .A(DP_OP_424J2_126_3477_n2658), .B(
        DP_OP_424J2_126_3477_n2177), .CI(DP_OP_424J2_126_3477_n2746), .CO(
        DP_OP_424J2_126_3477_n857), .S(DP_OP_424J2_126_3477_n858) );
  FADDX1_HVT DP_OP_424J2_126_3477_U524 ( .A(DP_OP_424J2_126_3477_n2834), .B(
        DP_OP_424J2_126_3477_n2482), .CI(DP_OP_424J2_126_3477_n1957), .CO(
        DP_OP_424J2_126_3477_n855), .S(DP_OP_424J2_126_3477_n856) );
  FADDX1_HVT DP_OP_424J2_126_3477_U523 ( .A(DP_OP_424J2_126_3477_n2133), .B(
        DP_OP_424J2_126_3477_n2438), .CI(DP_OP_424J2_126_3477_n2570), .CO(
        DP_OP_424J2_126_3477_n853), .S(DP_OP_424J2_126_3477_n854) );
  FADDX1_HVT DP_OP_424J2_126_3477_U522 ( .A(DP_OP_424J2_126_3477_n2790), .B(
        DP_OP_424J2_126_3477_n1978), .CI(DP_OP_424J2_126_3477_n2878), .CO(
        DP_OP_424J2_126_3477_n851), .S(DP_OP_424J2_126_3477_n852) );
  FADDX1_HVT DP_OP_424J2_126_3477_U521 ( .A(DP_OP_424J2_126_3477_n2309), .B(
        DP_OP_424J2_126_3477_n2679), .CI(DP_OP_424J2_126_3477_n2022), .CO(
        DP_OP_424J2_126_3477_n849), .S(DP_OP_424J2_126_3477_n850) );
  FADDX1_HVT DP_OP_424J2_126_3477_U520 ( .A(DP_OP_424J2_126_3477_n2614), .B(
        DP_OP_424J2_126_3477_n2110), .CI(DP_OP_424J2_126_3477_n2330), .CO(
        DP_OP_424J2_126_3477_n847), .S(DP_OP_424J2_126_3477_n848) );
  FADDX1_HVT DP_OP_424J2_126_3477_U519 ( .A(DP_OP_424J2_126_3477_n2265), .B(
        DP_OP_424J2_126_3477_n1846), .CI(DP_OP_424J2_126_3477_n2635), .CO(
        DP_OP_424J2_126_3477_n845), .S(DP_OP_424J2_126_3477_n846) );
  FADDX1_HVT DP_OP_424J2_126_3477_U518 ( .A(DP_OP_424J2_126_3477_n2459), .B(
        DP_OP_424J2_126_3477_n2547), .CI(DP_OP_424J2_126_3477_n2286), .CO(
        DP_OP_424J2_126_3477_n843), .S(DP_OP_424J2_126_3477_n844) );
  FADDX1_HVT DP_OP_424J2_126_3477_U517 ( .A(DP_OP_424J2_126_3477_n2198), .B(
        DP_OP_424J2_126_3477_n2591), .CI(DP_OP_424J2_126_3477_n2066), .CO(
        DP_OP_424J2_126_3477_n841), .S(DP_OP_424J2_126_3477_n842) );
  FADDX1_HVT DP_OP_424J2_126_3477_U516 ( .A(DP_OP_424J2_126_3477_n2415), .B(
        DP_OP_424J2_126_3477_n2221), .CI(DP_OP_424J2_126_3477_n2841), .CO(
        DP_OP_424J2_126_3477_n839), .S(DP_OP_424J2_126_3477_n840) );
  FADDX1_HVT DP_OP_424J2_126_3477_U515 ( .A(DP_OP_424J2_126_3477_n2885), .B(
        DP_OP_424J2_126_3477_n2242), .CI(DP_OP_424J2_126_3477_n2140), .CO(
        DP_OP_424J2_126_3477_n837), .S(DP_OP_424J2_126_3477_n838) );
  FADDX1_HVT DP_OP_424J2_126_3477_U514 ( .A(DP_OP_424J2_126_3477_n1934), .B(
        DP_OP_424J2_126_3477_n1964), .CI(DP_OP_424J2_126_3477_n2272), .CO(
        DP_OP_424J2_126_3477_n835), .S(DP_OP_424J2_126_3477_n836) );
  FADDX1_HVT DP_OP_424J2_126_3477_U513 ( .A(DP_OP_424J2_126_3477_n2059), .B(
        DP_OP_424J2_126_3477_n2408), .CI(DP_OP_424J2_126_3477_n2899), .CO(
        DP_OP_424J2_126_3477_n833), .S(DP_OP_424J2_126_3477_n834) );
  FADDX1_HVT DP_OP_424J2_126_3477_U512 ( .A(DP_OP_424J2_126_3477_n2628), .B(
        DP_OP_424J2_126_3477_n2533), .CI(DP_OP_424J2_126_3477_n2371), .CO(
        DP_OP_424J2_126_3477_n831), .S(DP_OP_424J2_126_3477_n832) );
  FADDX1_HVT DP_OP_424J2_126_3477_U511 ( .A(DP_OP_424J2_126_3477_n1839), .B(
        DP_OP_424J2_126_3477_n2147), .CI(DP_OP_424J2_126_3477_n2154), .CO(
        DP_OP_424J2_126_3477_n829), .S(DP_OP_424J2_126_3477_n830) );
  FADDX1_HVT DP_OP_424J2_126_3477_U510 ( .A(DP_OP_424J2_126_3477_n2323), .B(
        DP_OP_424J2_126_3477_n1781), .CI(DP_OP_424J2_126_3477_n2228), .CO(
        DP_OP_424J2_126_3477_n827), .S(DP_OP_424J2_126_3477_n828) );
  FADDX1_HVT DP_OP_424J2_126_3477_U509 ( .A(DP_OP_424J2_126_3477_n2753), .B(
        DP_OP_424J2_126_3477_n2496), .CI(DP_OP_424J2_126_3477_n2096), .CO(
        DP_OP_424J2_126_3477_n825), .S(DP_OP_424J2_126_3477_n826) );
  FADDX1_HVT DP_OP_424J2_126_3477_U508 ( .A(DP_OP_424J2_126_3477_n2584), .B(
        DP_OP_424J2_126_3477_n2577), .CI(DP_OP_424J2_126_3477_n2445), .CO(
        DP_OP_424J2_126_3477_n823), .S(DP_OP_424J2_126_3477_n824) );
  FADDX1_HVT DP_OP_424J2_126_3477_U507 ( .A(DP_OP_424J2_126_3477_n2540), .B(
        DP_OP_424J2_126_3477_n2760), .CI(DP_OP_424J2_126_3477_n2364), .CO(
        DP_OP_424J2_126_3477_n821), .S(DP_OP_424J2_126_3477_n822) );
  FADDX1_HVT DP_OP_424J2_126_3477_U506 ( .A(DP_OP_424J2_126_3477_n2709), .B(
        DP_OP_424J2_126_3477_n2452), .CI(DP_OP_424J2_126_3477_n2008), .CO(
        DP_OP_424J2_126_3477_n819), .S(DP_OP_424J2_126_3477_n820) );
  FADDX1_HVT DP_OP_424J2_126_3477_U505 ( .A(DP_OP_424J2_126_3477_n2848), .B(
        DP_OP_424J2_126_3477_n2811), .CI(DP_OP_424J2_126_3477_n2191), .CO(
        DP_OP_424J2_126_3477_n817), .S(DP_OP_424J2_126_3477_n818) );
  FADDX1_HVT DP_OP_424J2_126_3477_U504 ( .A(DP_OP_424J2_126_3477_n2489), .B(
        DP_OP_424J2_126_3477_n2279), .CI(DP_OP_424J2_126_3477_n2235), .CO(
        DP_OP_424J2_126_3477_n815), .S(DP_OP_424J2_126_3477_n816) );
  FADDX1_HVT DP_OP_424J2_126_3477_U503 ( .A(DP_OP_424J2_126_3477_n1883), .B(
        DP_OP_424J2_126_3477_n2804), .CI(DP_OP_424J2_126_3477_n1061), .CO(
        DP_OP_424J2_126_3477_n813), .S(DP_OP_424J2_126_3477_n814) );
  FADDX1_HVT DP_OP_424J2_126_3477_U502 ( .A(DP_OP_424J2_126_3477_n2103), .B(
        DP_OP_424J2_126_3477_n2665), .CI(DP_OP_424J2_126_3477_n1927), .CO(
        DP_OP_424J2_126_3477_n811), .S(DP_OP_424J2_126_3477_n812) );
  FADDX1_HVT DP_OP_424J2_126_3477_U501 ( .A(DP_OP_424J2_126_3477_n2357), .B(
        DP_OP_424J2_126_3477_n2892), .CI(DP_OP_424J2_126_3477_n2716), .CO(
        DP_OP_424J2_126_3477_n809), .S(DP_OP_424J2_126_3477_n810) );
  FADDX1_HVT DP_OP_424J2_126_3477_U500 ( .A(DP_OP_424J2_126_3477_n2672), .B(
        DP_OP_424J2_126_3477_n2052), .CI(DP_OP_424J2_126_3477_n2015), .CO(
        DP_OP_424J2_126_3477_n807), .S(DP_OP_424J2_126_3477_n808) );
  FADDX1_HVT DP_OP_424J2_126_3477_U499 ( .A(DP_OP_424J2_126_3477_n2316), .B(
        DP_OP_424J2_126_3477_n2797), .CI(DP_OP_424J2_126_3477_n2401), .CO(
        DP_OP_424J2_126_3477_n805), .S(DP_OP_424J2_126_3477_n806) );
  FADDX1_HVT DP_OP_424J2_126_3477_U498 ( .A(DP_OP_424J2_126_3477_n2621), .B(
        DP_OP_424J2_126_3477_n1920), .CI(DP_OP_424J2_126_3477_n2184), .CO(
        DP_OP_424J2_126_3477_n803), .S(DP_OP_424J2_126_3477_n804) );
  FADDX1_HVT DP_OP_424J2_126_3477_U497 ( .A(DP_OP_424J2_126_3477_n1971), .B(
        DP_OP_424J2_126_3477_n1876), .CI(DP_OP_424J2_126_3477_n1832), .CO(
        DP_OP_424J2_126_3477_n801), .S(DP_OP_424J2_126_3477_n802) );
  FADDX1_HVT DP_OP_424J2_126_3477_U496 ( .A(DP_OP_424J2_126_3477_n1059), .B(
        DP_OP_424J2_126_3477_n1057), .CI(DP_OP_424J2_126_3477_n1045), .CO(
        DP_OP_424J2_126_3477_n799), .S(DP_OP_424J2_126_3477_n800) );
  FADDX1_HVT DP_OP_424J2_126_3477_U495 ( .A(DP_OP_424J2_126_3477_n1047), .B(
        DP_OP_424J2_126_3477_n1055), .CI(DP_OP_424J2_126_3477_n1053), .CO(
        DP_OP_424J2_126_3477_n797), .S(DP_OP_424J2_126_3477_n798) );
  FADDX1_HVT DP_OP_424J2_126_3477_U494 ( .A(DP_OP_424J2_126_3477_n1051), .B(
        DP_OP_424J2_126_3477_n1049), .CI(DP_OP_424J2_126_3477_n1043), .CO(
        DP_OP_424J2_126_3477_n795), .S(DP_OP_424J2_126_3477_n796) );
  FADDX1_HVT DP_OP_424J2_126_3477_U493 ( .A(DP_OP_424J2_126_3477_n1041), .B(
        DP_OP_424J2_126_3477_n1019), .CI(DP_OP_424J2_126_3477_n1021), .CO(
        DP_OP_424J2_126_3477_n793), .S(DP_OP_424J2_126_3477_n794) );
  FADDX1_HVT DP_OP_424J2_126_3477_U492 ( .A(DP_OP_424J2_126_3477_n1039), .B(
        DP_OP_424J2_126_3477_n1025), .CI(DP_OP_424J2_126_3477_n1023), .CO(
        DP_OP_424J2_126_3477_n791), .S(DP_OP_424J2_126_3477_n792) );
  FADDX1_HVT DP_OP_424J2_126_3477_U491 ( .A(DP_OP_424J2_126_3477_n1037), .B(
        DP_OP_424J2_126_3477_n1027), .CI(DP_OP_424J2_126_3477_n1029), .CO(
        DP_OP_424J2_126_3477_n789), .S(DP_OP_424J2_126_3477_n790) );
  FADDX1_HVT DP_OP_424J2_126_3477_U490 ( .A(DP_OP_424J2_126_3477_n1035), .B(
        DP_OP_424J2_126_3477_n1033), .CI(DP_OP_424J2_126_3477_n1031), .CO(
        DP_OP_424J2_126_3477_n787), .S(DP_OP_424J2_126_3477_n788) );
  FADDX1_HVT DP_OP_424J2_126_3477_U489 ( .A(DP_OP_424J2_126_3477_n1015), .B(
        DP_OP_424J2_126_3477_n868), .CI(DP_OP_424J2_126_3477_n995), .CO(
        DP_OP_424J2_126_3477_n785), .S(DP_OP_424J2_126_3477_n786) );
  FADDX1_HVT DP_OP_424J2_126_3477_U488 ( .A(DP_OP_424J2_126_3477_n1017), .B(
        DP_OP_424J2_126_3477_n1001), .CI(DP_OP_424J2_126_3477_n997), .CO(
        DP_OP_424J2_126_3477_n783), .S(DP_OP_424J2_126_3477_n784) );
  FADDX1_HVT DP_OP_424J2_126_3477_U487 ( .A(DP_OP_424J2_126_3477_n1013), .B(
        DP_OP_424J2_126_3477_n866), .CI(DP_OP_424J2_126_3477_n999), .CO(
        DP_OP_424J2_126_3477_n781), .S(DP_OP_424J2_126_3477_n782) );
  FADDX1_HVT DP_OP_424J2_126_3477_U486 ( .A(DP_OP_424J2_126_3477_n1011), .B(
        DP_OP_424J2_126_3477_n846), .CI(DP_OP_424J2_126_3477_n844), .CO(
        DP_OP_424J2_126_3477_n779), .S(DP_OP_424J2_126_3477_n780) );
  FADDX1_HVT DP_OP_424J2_126_3477_U485 ( .A(DP_OP_424J2_126_3477_n1007), .B(
        DP_OP_424J2_126_3477_n860), .CI(DP_OP_424J2_126_3477_n842), .CO(
        DP_OP_424J2_126_3477_n777), .S(DP_OP_424J2_126_3477_n778) );
  FADDX1_HVT DP_OP_424J2_126_3477_U484 ( .A(DP_OP_424J2_126_3477_n1009), .B(
        DP_OP_424J2_126_3477_n858), .CI(DP_OP_424J2_126_3477_n850), .CO(
        DP_OP_424J2_126_3477_n775), .S(DP_OP_424J2_126_3477_n776) );
  FADDX1_HVT DP_OP_424J2_126_3477_U483 ( .A(DP_OP_424J2_126_3477_n1005), .B(
        DP_OP_424J2_126_3477_n852), .CI(DP_OP_424J2_126_3477_n848), .CO(
        DP_OP_424J2_126_3477_n773), .S(DP_OP_424J2_126_3477_n774) );
  FADDX1_HVT DP_OP_424J2_126_3477_U482 ( .A(DP_OP_424J2_126_3477_n1003), .B(
        DP_OP_424J2_126_3477_n854), .CI(DP_OP_424J2_126_3477_n862), .CO(
        DP_OP_424J2_126_3477_n771), .S(DP_OP_424J2_126_3477_n772) );
  FADDX1_HVT DP_OP_424J2_126_3477_U481 ( .A(DP_OP_424J2_126_3477_n864), .B(
        DP_OP_424J2_126_3477_n856), .CI(DP_OP_424J2_126_3477_n840), .CO(
        DP_OP_424J2_126_3477_n769), .S(DP_OP_424J2_126_3477_n770) );
  FADDX1_HVT DP_OP_424J2_126_3477_U480 ( .A(DP_OP_424J2_126_3477_n838), .B(
        DP_OP_424J2_126_3477_n826), .CI(DP_OP_424J2_126_3477_n824), .CO(
        DP_OP_424J2_126_3477_n767), .S(DP_OP_424J2_126_3477_n768) );
  FADDX1_HVT DP_OP_424J2_126_3477_U479 ( .A(DP_OP_424J2_126_3477_n836), .B(
        DP_OP_424J2_126_3477_n832), .CI(DP_OP_424J2_126_3477_n834), .CO(
        DP_OP_424J2_126_3477_n765), .S(DP_OP_424J2_126_3477_n766) );
  FADDX1_HVT DP_OP_424J2_126_3477_U478 ( .A(DP_OP_424J2_126_3477_n828), .B(
        DP_OP_424J2_126_3477_n830), .CI(DP_OP_424J2_126_3477_n820), .CO(
        DP_OP_424J2_126_3477_n763), .S(DP_OP_424J2_126_3477_n764) );
  FADDX1_HVT DP_OP_424J2_126_3477_U477 ( .A(DP_OP_424J2_126_3477_n822), .B(
        DP_OP_424J2_126_3477_n806), .CI(DP_OP_424J2_126_3477_n802), .CO(
        DP_OP_424J2_126_3477_n761), .S(DP_OP_424J2_126_3477_n762) );
  FADDX1_HVT DP_OP_424J2_126_3477_U476 ( .A(DP_OP_424J2_126_3477_n818), .B(
        DP_OP_424J2_126_3477_n808), .CI(DP_OP_424J2_126_3477_n804), .CO(
        DP_OP_424J2_126_3477_n759), .S(DP_OP_424J2_126_3477_n760) );
  FADDX1_HVT DP_OP_424J2_126_3477_U475 ( .A(DP_OP_424J2_126_3477_n812), .B(
        DP_OP_424J2_126_3477_n816), .CI(DP_OP_424J2_126_3477_n810), .CO(
        DP_OP_424J2_126_3477_n757), .S(DP_OP_424J2_126_3477_n758) );
  FADDX1_HVT DP_OP_424J2_126_3477_U474 ( .A(DP_OP_424J2_126_3477_n814), .B(
        DP_OP_424J2_126_3477_n993), .CI(DP_OP_424J2_126_3477_n991), .CO(
        DP_OP_424J2_126_3477_n755), .S(DP_OP_424J2_126_3477_n756) );
  FADDX1_HVT DP_OP_424J2_126_3477_U473 ( .A(DP_OP_424J2_126_3477_n989), .B(
        DP_OP_424J2_126_3477_n987), .CI(DP_OP_424J2_126_3477_n985), .CO(
        DP_OP_424J2_126_3477_n753), .S(DP_OP_424J2_126_3477_n754) );
  FADDX1_HVT DP_OP_424J2_126_3477_U472 ( .A(DP_OP_424J2_126_3477_n983), .B(
        DP_OP_424J2_126_3477_n979), .CI(DP_OP_424J2_126_3477_n981), .CO(
        DP_OP_424J2_126_3477_n751), .S(DP_OP_424J2_126_3477_n752) );
  FADDX1_HVT DP_OP_424J2_126_3477_U471 ( .A(DP_OP_424J2_126_3477_n977), .B(
        DP_OP_424J2_126_3477_n967), .CI(DP_OP_424J2_126_3477_n796), .CO(
        DP_OP_424J2_126_3477_n749), .S(DP_OP_424J2_126_3477_n750) );
  FADDX1_HVT DP_OP_424J2_126_3477_U470 ( .A(DP_OP_424J2_126_3477_n975), .B(
        DP_OP_424J2_126_3477_n800), .CI(DP_OP_424J2_126_3477_n798), .CO(
        DP_OP_424J2_126_3477_n747), .S(DP_OP_424J2_126_3477_n748) );
  FADDX1_HVT DP_OP_424J2_126_3477_U469 ( .A(DP_OP_424J2_126_3477_n973), .B(
        DP_OP_424J2_126_3477_n969), .CI(DP_OP_424J2_126_3477_n971), .CO(
        DP_OP_424J2_126_3477_n745), .S(DP_OP_424J2_126_3477_n746) );
  FADDX1_HVT DP_OP_424J2_126_3477_U468 ( .A(DP_OP_424J2_126_3477_n965), .B(
        DP_OP_424J2_126_3477_n788), .CI(DP_OP_424J2_126_3477_n792), .CO(
        DP_OP_424J2_126_3477_n743), .S(DP_OP_424J2_126_3477_n744) );
  FADDX1_HVT DP_OP_424J2_126_3477_U467 ( .A(DP_OP_424J2_126_3477_n959), .B(
        DP_OP_424J2_126_3477_n790), .CI(DP_OP_424J2_126_3477_n794), .CO(
        DP_OP_424J2_126_3477_n741), .S(DP_OP_424J2_126_3477_n742) );
  FADDX1_HVT DP_OP_424J2_126_3477_U466 ( .A(DP_OP_424J2_126_3477_n963), .B(
        DP_OP_424J2_126_3477_n957), .CI(DP_OP_424J2_126_3477_n961), .CO(
        DP_OP_424J2_126_3477_n739), .S(DP_OP_424J2_126_3477_n740) );
  FADDX1_HVT DP_OP_424J2_126_3477_U465 ( .A(DP_OP_424J2_126_3477_n955), .B(
        DP_OP_424J2_126_3477_n772), .CI(DP_OP_424J2_126_3477_n770), .CO(
        DP_OP_424J2_126_3477_n737), .S(DP_OP_424J2_126_3477_n738) );
  FADDX1_HVT DP_OP_424J2_126_3477_U464 ( .A(DP_OP_424J2_126_3477_n784), .B(
        DP_OP_424J2_126_3477_n949), .CI(DP_OP_424J2_126_3477_n774), .CO(
        DP_OP_424J2_126_3477_n735), .S(DP_OP_424J2_126_3477_n736) );
  FADDX1_HVT DP_OP_424J2_126_3477_U463 ( .A(DP_OP_424J2_126_3477_n786), .B(
        DP_OP_424J2_126_3477_n780), .CI(DP_OP_424J2_126_3477_n776), .CO(
        DP_OP_424J2_126_3477_n733), .S(DP_OP_424J2_126_3477_n734) );
  FADDX1_HVT DP_OP_424J2_126_3477_U462 ( .A(DP_OP_424J2_126_3477_n953), .B(
        DP_OP_424J2_126_3477_n778), .CI(DP_OP_424J2_126_3477_n951), .CO(
        DP_OP_424J2_126_3477_n731), .S(DP_OP_424J2_126_3477_n732) );
  FADDX1_HVT DP_OP_424J2_126_3477_U461 ( .A(DP_OP_424J2_126_3477_n782), .B(
        DP_OP_424J2_126_3477_n768), .CI(DP_OP_424J2_126_3477_n766), .CO(
        DP_OP_424J2_126_3477_n729), .S(DP_OP_424J2_126_3477_n730) );
  FADDX1_HVT DP_OP_424J2_126_3477_U460 ( .A(DP_OP_424J2_126_3477_n947), .B(
        DP_OP_424J2_126_3477_n764), .CI(DP_OP_424J2_126_3477_n762), .CO(
        DP_OP_424J2_126_3477_n727), .S(DP_OP_424J2_126_3477_n728) );
  FADDX1_HVT DP_OP_424J2_126_3477_U459 ( .A(DP_OP_424J2_126_3477_n760), .B(
        DP_OP_424J2_126_3477_n945), .CI(DP_OP_424J2_126_3477_n756), .CO(
        DP_OP_424J2_126_3477_n725), .S(DP_OP_424J2_126_3477_n726) );
  FADDX1_HVT DP_OP_424J2_126_3477_U458 ( .A(DP_OP_424J2_126_3477_n758), .B(
        DP_OP_424J2_126_3477_n943), .CI(DP_OP_424J2_126_3477_n941), .CO(
        DP_OP_424J2_126_3477_n723), .S(DP_OP_424J2_126_3477_n724) );
  FADDX1_HVT DP_OP_424J2_126_3477_U457 ( .A(DP_OP_424J2_126_3477_n939), .B(
        DP_OP_424J2_126_3477_n937), .CI(DP_OP_424J2_126_3477_n754), .CO(
        DP_OP_424J2_126_3477_n721), .S(DP_OP_424J2_126_3477_n722) );
  FADDX1_HVT DP_OP_424J2_126_3477_U456 ( .A(DP_OP_424J2_126_3477_n935), .B(
        DP_OP_424J2_126_3477_n752), .CI(DP_OP_424J2_126_3477_n931), .CO(
        DP_OP_424J2_126_3477_n719), .S(DP_OP_424J2_126_3477_n720) );
  FADDX1_HVT DP_OP_424J2_126_3477_U455 ( .A(DP_OP_424J2_126_3477_n933), .B(
        DP_OP_424J2_126_3477_n929), .CI(DP_OP_424J2_126_3477_n750), .CO(
        DP_OP_424J2_126_3477_n717), .S(DP_OP_424J2_126_3477_n718) );
  FADDX1_HVT DP_OP_424J2_126_3477_U454 ( .A(DP_OP_424J2_126_3477_n927), .B(
        DP_OP_424J2_126_3477_n748), .CI(DP_OP_424J2_126_3477_n746), .CO(
        DP_OP_424J2_126_3477_n715), .S(DP_OP_424J2_126_3477_n716) );
  FADDX1_HVT DP_OP_424J2_126_3477_U453 ( .A(DP_OP_424J2_126_3477_n925), .B(
        DP_OP_424J2_126_3477_n923), .CI(DP_OP_424J2_126_3477_n744), .CO(
        DP_OP_424J2_126_3477_n713), .S(DP_OP_424J2_126_3477_n714) );
  FADDX1_HVT DP_OP_424J2_126_3477_U452 ( .A(DP_OP_424J2_126_3477_n921), .B(
        DP_OP_424J2_126_3477_n740), .CI(DP_OP_424J2_126_3477_n742), .CO(
        DP_OP_424J2_126_3477_n711), .S(DP_OP_424J2_126_3477_n712) );
  FADDX1_HVT DP_OP_424J2_126_3477_U451 ( .A(DP_OP_424J2_126_3477_n919), .B(
        DP_OP_424J2_126_3477_n917), .CI(DP_OP_424J2_126_3477_n732), .CO(
        DP_OP_424J2_126_3477_n709), .S(DP_OP_424J2_126_3477_n710) );
  FADDX1_HVT DP_OP_424J2_126_3477_U450 ( .A(DP_OP_424J2_126_3477_n736), .B(
        DP_OP_424J2_126_3477_n734), .CI(DP_OP_424J2_126_3477_n738), .CO(
        DP_OP_424J2_126_3477_n707), .S(DP_OP_424J2_126_3477_n708) );
  FADDX1_HVT DP_OP_424J2_126_3477_U449 ( .A(DP_OP_424J2_126_3477_n730), .B(
        DP_OP_424J2_126_3477_n915), .CI(DP_OP_424J2_126_3477_n728), .CO(
        DP_OP_424J2_126_3477_n705), .S(DP_OP_424J2_126_3477_n706) );
  FADDX1_HVT DP_OP_424J2_126_3477_U448 ( .A(DP_OP_424J2_126_3477_n913), .B(
        DP_OP_424J2_126_3477_n726), .CI(DP_OP_424J2_126_3477_n724), .CO(
        DP_OP_424J2_126_3477_n703), .S(DP_OP_424J2_126_3477_n704) );
  FADDX1_HVT DP_OP_424J2_126_3477_U447 ( .A(DP_OP_424J2_126_3477_n911), .B(
        DP_OP_424J2_126_3477_n909), .CI(DP_OP_424J2_126_3477_n907), .CO(
        DP_OP_424J2_126_3477_n701), .S(DP_OP_424J2_126_3477_n702) );
  FADDX1_HVT DP_OP_424J2_126_3477_U446 ( .A(DP_OP_424J2_126_3477_n722), .B(
        DP_OP_424J2_126_3477_n905), .CI(DP_OP_424J2_126_3477_n903), .CO(
        DP_OP_424J2_126_3477_n699), .S(DP_OP_424J2_126_3477_n700) );
  FADDX1_HVT DP_OP_424J2_126_3477_U445 ( .A(DP_OP_424J2_126_3477_n720), .B(
        DP_OP_424J2_126_3477_n718), .CI(DP_OP_424J2_126_3477_n901), .CO(
        DP_OP_424J2_126_3477_n697), .S(DP_OP_424J2_126_3477_n698) );
  FADDX1_HVT DP_OP_424J2_126_3477_U444 ( .A(DP_OP_424J2_126_3477_n716), .B(
        DP_OP_424J2_126_3477_n899), .CI(DP_OP_424J2_126_3477_n714), .CO(
        DP_OP_424J2_126_3477_n695), .S(DP_OP_424J2_126_3477_n696) );
  FADDX1_HVT DP_OP_424J2_126_3477_U443 ( .A(DP_OP_424J2_126_3477_n712), .B(
        DP_OP_424J2_126_3477_n897), .CI(DP_OP_424J2_126_3477_n710), .CO(
        DP_OP_424J2_126_3477_n693), .S(DP_OP_424J2_126_3477_n694) );
  FADDX1_HVT DP_OP_424J2_126_3477_U442 ( .A(DP_OP_424J2_126_3477_n708), .B(
        DP_OP_424J2_126_3477_n895), .CI(DP_OP_424J2_126_3477_n706), .CO(
        DP_OP_424J2_126_3477_n691), .S(DP_OP_424J2_126_3477_n692) );
  FADDX1_HVT DP_OP_424J2_126_3477_U441 ( .A(DP_OP_424J2_126_3477_n893), .B(
        DP_OP_424J2_126_3477_n704), .CI(DP_OP_424J2_126_3477_n891), .CO(
        DP_OP_424J2_126_3477_n689), .S(DP_OP_424J2_126_3477_n690) );
  FADDX1_HVT DP_OP_424J2_126_3477_U440 ( .A(DP_OP_424J2_126_3477_n702), .B(
        DP_OP_424J2_126_3477_n889), .CI(DP_OP_424J2_126_3477_n700), .CO(
        DP_OP_424J2_126_3477_n687), .S(DP_OP_424J2_126_3477_n688) );
  FADDX1_HVT DP_OP_424J2_126_3477_U439 ( .A(DP_OP_424J2_126_3477_n887), .B(
        DP_OP_424J2_126_3477_n698), .CI(DP_OP_424J2_126_3477_n885), .CO(
        DP_OP_424J2_126_3477_n685), .S(DP_OP_424J2_126_3477_n686) );
  FADDX1_HVT DP_OP_424J2_126_3477_U438 ( .A(DP_OP_424J2_126_3477_n696), .B(
        DP_OP_424J2_126_3477_n883), .CI(DP_OP_424J2_126_3477_n694), .CO(
        DP_OP_424J2_126_3477_n683), .S(DP_OP_424J2_126_3477_n684) );
  FADDX1_HVT DP_OP_424J2_126_3477_U437 ( .A(DP_OP_424J2_126_3477_n692), .B(
        DP_OP_424J2_126_3477_n881), .CI(DP_OP_424J2_126_3477_n690), .CO(
        DP_OP_424J2_126_3477_n681), .S(DP_OP_424J2_126_3477_n682) );
  FADDX1_HVT DP_OP_424J2_126_3477_U436 ( .A(DP_OP_424J2_126_3477_n879), .B(
        DP_OP_424J2_126_3477_n688), .CI(DP_OP_424J2_126_3477_n877), .CO(
        DP_OP_424J2_126_3477_n679), .S(DP_OP_424J2_126_3477_n680) );
  FADDX1_HVT DP_OP_424J2_126_3477_U435 ( .A(DP_OP_424J2_126_3477_n686), .B(
        DP_OP_424J2_126_3477_n875), .CI(DP_OP_424J2_126_3477_n684), .CO(
        DP_OP_424J2_126_3477_n677), .S(DP_OP_424J2_126_3477_n678) );
  FADDX1_HVT DP_OP_424J2_126_3477_U434 ( .A(DP_OP_424J2_126_3477_n682), .B(
        DP_OP_424J2_126_3477_n873), .CI(DP_OP_424J2_126_3477_n680), .CO(
        DP_OP_424J2_126_3477_n675), .S(DP_OP_424J2_126_3477_n676) );
  FADDX1_HVT DP_OP_424J2_126_3477_U433 ( .A(DP_OP_424J2_126_3477_n871), .B(
        DP_OP_424J2_126_3477_n678), .CI(DP_OP_424J2_126_3477_n676), .CO(
        DP_OP_424J2_126_3477_n673), .S(DP_OP_424J2_126_3477_n674) );
  FADDX1_HVT DP_OP_424J2_126_3477_U431 ( .A(DP_OP_424J2_126_3477_n2000), .B(
        DP_OP_424J2_126_3477_n2146), .CI(DP_OP_424J2_126_3477_n2393), .CO(
        DP_OP_424J2_126_3477_n669), .S(DP_OP_424J2_126_3477_n670) );
  FADDX1_HVT DP_OP_424J2_126_3477_U430 ( .A(DP_OP_424J2_126_3477_n2701), .B(
        DP_OP_424J2_126_3477_n2407), .CI(DP_OP_424J2_126_3477_n1956), .CO(
        DP_OP_424J2_126_3477_n667), .S(DP_OP_424J2_126_3477_n668) );
  FADDX1_HVT DP_OP_424J2_126_3477_U429 ( .A(DP_OP_424J2_126_3477_n2308), .B(
        DP_OP_424J2_126_3477_n1824), .CI(DP_OP_424J2_126_3477_n2745), .CO(
        DP_OP_424J2_126_3477_n665), .S(DP_OP_424J2_126_3477_n666) );
  FADDX1_HVT DP_OP_424J2_126_3477_U428 ( .A(DP_OP_424J2_126_3477_n2132), .B(
        DP_OP_424J2_126_3477_n2437), .CI(DP_OP_424J2_126_3477_n2481), .CO(
        DP_OP_424J2_126_3477_n663), .S(DP_OP_424J2_126_3477_n664) );
  FADDX1_HVT DP_OP_424J2_126_3477_U427 ( .A(DP_OP_424J2_126_3477_n1868), .B(
        DP_OP_424J2_126_3477_n1912), .CI(DP_OP_424J2_126_3477_n2044), .CO(
        DP_OP_424J2_126_3477_n661), .S(DP_OP_424J2_126_3477_n662) );
  FADDX1_HVT DP_OP_424J2_126_3477_U426 ( .A(DP_OP_424J2_126_3477_n2088), .B(
        DP_OP_424J2_126_3477_n2176), .CI(DP_OP_424J2_126_3477_n2569), .CO(
        DP_OP_424J2_126_3477_n659), .S(DP_OP_424J2_126_3477_n660) );
  FADDX1_HVT DP_OP_424J2_126_3477_U425 ( .A(DP_OP_424J2_126_3477_n2789), .B(
        DP_OP_424J2_126_3477_n2877), .CI(DP_OP_424J2_126_3477_n2525), .CO(
        DP_OP_424J2_126_3477_n657), .S(DP_OP_424J2_126_3477_n658) );
  FADDX1_HVT DP_OP_424J2_126_3477_U424 ( .A(DP_OP_424J2_126_3477_n2613), .B(
        DP_OP_424J2_126_3477_n2495), .CI(DP_OP_424J2_126_3477_n2322), .CO(
        DP_OP_424J2_126_3477_n655), .S(DP_OP_424J2_126_3477_n656) );
  FADDX1_HVT DP_OP_424J2_126_3477_U423 ( .A(DP_OP_424J2_126_3477_n2833), .B(
        DP_OP_424J2_126_3477_n2583), .CI(DP_OP_424J2_126_3477_n2627), .CO(
        DP_OP_424J2_126_3477_n653), .S(DP_OP_424J2_126_3477_n654) );
  FADDX1_HVT DP_OP_424J2_126_3477_U422 ( .A(DP_OP_424J2_126_3477_n2657), .B(
        DP_OP_424J2_126_3477_n2058), .CI(DP_OP_424J2_126_3477_n1838), .CO(
        DP_OP_424J2_126_3477_n651), .S(DP_OP_424J2_126_3477_n652) );
  FADDX1_HVT DP_OP_424J2_126_3477_U421 ( .A(DP_OP_424J2_126_3477_n2264), .B(
        DP_OP_424J2_126_3477_n672), .CI(DP_OP_424J2_126_3477_n2220), .CO(
        DP_OP_424J2_126_3477_n649), .S(DP_OP_424J2_126_3477_n650) );
  FADDX1_HVT DP_OP_424J2_126_3477_U420 ( .A(DP_OP_424J2_126_3477_n2840), .B(
        DP_OP_424J2_126_3477_n2451), .CI(DP_OP_424J2_126_3477_n2139), .CO(
        DP_OP_424J2_126_3477_n647), .S(DP_OP_424J2_126_3477_n648) );
  FADDX1_HVT DP_OP_424J2_126_3477_U419 ( .A(DP_OP_424J2_126_3477_n2884), .B(
        DP_OP_424J2_126_3477_n2803), .CI(DP_OP_424J2_126_3477_n2271), .CO(
        DP_OP_424J2_126_3477_n645), .S(DP_OP_424J2_126_3477_n646) );
  FADDX1_HVT DP_OP_424J2_126_3477_U418 ( .A(DP_OP_424J2_126_3477_n2752), .B(
        DP_OP_424J2_126_3477_n2759), .CI(DP_OP_424J2_126_3477_n2363), .CO(
        DP_OP_424J2_126_3477_n643), .S(DP_OP_424J2_126_3477_n644) );
  FADDX1_HVT DP_OP_424J2_126_3477_U417 ( .A(DP_OP_424J2_126_3477_n2539), .B(
        DP_OP_424J2_126_3477_n2278), .CI(DP_OP_424J2_126_3477_n2190), .CO(
        DP_OP_424J2_126_3477_n641), .S(DP_OP_424J2_126_3477_n642) );
  FADDX1_HVT DP_OP_424J2_126_3477_U416 ( .A(DP_OP_424J2_126_3477_n2847), .B(
        DP_OP_424J2_126_3477_n2891), .CI(DP_OP_424J2_126_3477_n2234), .CO(
        DP_OP_424J2_126_3477_n639), .S(DP_OP_424J2_126_3477_n640) );
  FADDX1_HVT DP_OP_424J2_126_3477_U415 ( .A(DP_OP_424J2_126_3477_n1780), .B(
        DP_OP_424J2_126_3477_n2532), .CI(DP_OP_424J2_126_3477_n2708), .CO(
        DP_OP_424J2_126_3477_n637), .S(DP_OP_424J2_126_3477_n638) );
  FADDX1_HVT DP_OP_424J2_126_3477_U414 ( .A(DP_OP_424J2_126_3477_n2102), .B(
        DP_OP_424J2_126_3477_n1963), .CI(DP_OP_424J2_126_3477_n1926), .CO(
        DP_OP_424J2_126_3477_n635), .S(DP_OP_424J2_126_3477_n636) );
  FADDX1_HVT DP_OP_424J2_126_3477_U413 ( .A(DP_OP_424J2_126_3477_n1882), .B(
        DP_OP_424J2_126_3477_n2671), .CI(DP_OP_424J2_126_3477_n2715), .CO(
        DP_OP_424J2_126_3477_n633), .S(DP_OP_424J2_126_3477_n634) );
  FADDX1_HVT DP_OP_424J2_126_3477_U412 ( .A(DP_OP_424J2_126_3477_n2576), .B(
        DP_OP_424J2_126_3477_n2014), .CI(DP_OP_424J2_126_3477_n2664), .CO(
        DP_OP_424J2_126_3477_n631), .S(DP_OP_424J2_126_3477_n632) );
  FADDX1_HVT DP_OP_424J2_126_3477_U411 ( .A(DP_OP_424J2_126_3477_n1970), .B(
        DP_OP_424J2_126_3477_n2095), .CI(DP_OP_424J2_126_3477_n2315), .CO(
        DP_OP_424J2_126_3477_n629), .S(DP_OP_424J2_126_3477_n630) );
  FADDX1_HVT DP_OP_424J2_126_3477_U410 ( .A(DP_OP_424J2_126_3477_n2227), .B(
        DP_OP_424J2_126_3477_n2444), .CI(DP_OP_424J2_126_3477_n2051), .CO(
        DP_OP_424J2_126_3477_n627), .S(DP_OP_424J2_126_3477_n628) );
  FADDX1_HVT DP_OP_424J2_126_3477_U409 ( .A(DP_OP_424J2_126_3477_n2488), .B(
        DP_OP_424J2_126_3477_n2356), .CI(DP_OP_424J2_126_3477_n2007), .CO(
        DP_OP_424J2_126_3477_n625), .S(DP_OP_424J2_126_3477_n626) );
  FADDX1_HVT DP_OP_424J2_126_3477_U408 ( .A(DP_OP_424J2_126_3477_n2796), .B(
        DP_OP_424J2_126_3477_n1919), .CI(DP_OP_424J2_126_3477_n2400), .CO(
        DP_OP_424J2_126_3477_n623), .S(DP_OP_424J2_126_3477_n624) );
  FADDX1_HVT DP_OP_424J2_126_3477_U407 ( .A(DP_OP_424J2_126_3477_n2620), .B(
        DP_OP_424J2_126_3477_n1831), .CI(DP_OP_424J2_126_3477_n2183), .CO(
        DP_OP_424J2_126_3477_n621), .S(DP_OP_424J2_126_3477_n622) );
  FADDX1_HVT DP_OP_424J2_126_3477_U406 ( .A(DP_OP_424J2_126_3477_n1875), .B(
        DP_OP_424J2_126_3477_n867), .CI(DP_OP_424J2_126_3477_n865), .CO(
        DP_OP_424J2_126_3477_n619), .S(DP_OP_424J2_126_3477_n620) );
  FADDX1_HVT DP_OP_424J2_126_3477_U405 ( .A(DP_OP_424J2_126_3477_n863), .B(
        DP_OP_424J2_126_3477_n841), .CI(DP_OP_424J2_126_3477_n839), .CO(
        DP_OP_424J2_126_3477_n617), .S(DP_OP_424J2_126_3477_n618) );
  FADDX1_HVT DP_OP_424J2_126_3477_U404 ( .A(DP_OP_424J2_126_3477_n861), .B(
        DP_OP_424J2_126_3477_n845), .CI(DP_OP_424J2_126_3477_n843), .CO(
        DP_OP_424J2_126_3477_n615), .S(DP_OP_424J2_126_3477_n616) );
  FADDX1_HVT DP_OP_424J2_126_3477_U403 ( .A(DP_OP_424J2_126_3477_n859), .B(
        DP_OP_424J2_126_3477_n847), .CI(DP_OP_424J2_126_3477_n849), .CO(
        DP_OP_424J2_126_3477_n613), .S(DP_OP_424J2_126_3477_n614) );
  FADDX1_HVT DP_OP_424J2_126_3477_U402 ( .A(DP_OP_424J2_126_3477_n857), .B(
        DP_OP_424J2_126_3477_n851), .CI(DP_OP_424J2_126_3477_n853), .CO(
        DP_OP_424J2_126_3477_n611), .S(DP_OP_424J2_126_3477_n612) );
  FADDX1_HVT DP_OP_424J2_126_3477_U401 ( .A(DP_OP_424J2_126_3477_n855), .B(
        DP_OP_424J2_126_3477_n837), .CI(DP_OP_424J2_126_3477_n835), .CO(
        DP_OP_424J2_126_3477_n609), .S(DP_OP_424J2_126_3477_n610) );
  FADDX1_HVT DP_OP_424J2_126_3477_U400 ( .A(DP_OP_424J2_126_3477_n833), .B(
        DP_OP_424J2_126_3477_n825), .CI(DP_OP_424J2_126_3477_n823), .CO(
        DP_OP_424J2_126_3477_n607), .S(DP_OP_424J2_126_3477_n608) );
  FADDX1_HVT DP_OP_424J2_126_3477_U399 ( .A(DP_OP_424J2_126_3477_n831), .B(
        DP_OP_424J2_126_3477_n827), .CI(DP_OP_424J2_126_3477_n829), .CO(
        DP_OP_424J2_126_3477_n605), .S(DP_OP_424J2_126_3477_n606) );
  FADDX1_HVT DP_OP_424J2_126_3477_U398 ( .A(DP_OP_424J2_126_3477_n821), .B(
        DP_OP_424J2_126_3477_n805), .CI(DP_OP_424J2_126_3477_n801), .CO(
        DP_OP_424J2_126_3477_n603), .S(DP_OP_424J2_126_3477_n604) );
  FADDX1_HVT DP_OP_424J2_126_3477_U397 ( .A(DP_OP_424J2_126_3477_n819), .B(
        DP_OP_424J2_126_3477_n807), .CI(DP_OP_424J2_126_3477_n803), .CO(
        DP_OP_424J2_126_3477_n601), .S(DP_OP_424J2_126_3477_n602) );
  FADDX1_HVT DP_OP_424J2_126_3477_U396 ( .A(DP_OP_424J2_126_3477_n817), .B(
        DP_OP_424J2_126_3477_n670), .CI(DP_OP_424J2_126_3477_n654), .CO(
        DP_OP_424J2_126_3477_n599), .S(DP_OP_424J2_126_3477_n600) );
  FADDX1_HVT DP_OP_424J2_126_3477_U395 ( .A(DP_OP_424J2_126_3477_n815), .B(
        DP_OP_424J2_126_3477_n652), .CI(DP_OP_424J2_126_3477_n662), .CO(
        DP_OP_424J2_126_3477_n597), .S(DP_OP_424J2_126_3477_n598) );
  FADDX1_HVT DP_OP_424J2_126_3477_U394 ( .A(DP_OP_424J2_126_3477_n813), .B(
        DP_OP_424J2_126_3477_n658), .CI(DP_OP_424J2_126_3477_n660), .CO(
        DP_OP_424J2_126_3477_n595), .S(DP_OP_424J2_126_3477_n596) );
  FADDX1_HVT DP_OP_424J2_126_3477_U393 ( .A(DP_OP_424J2_126_3477_n811), .B(
        DP_OP_424J2_126_3477_n664), .CI(DP_OP_424J2_126_3477_n666), .CO(
        DP_OP_424J2_126_3477_n593), .S(DP_OP_424J2_126_3477_n594) );
  FADDX1_HVT DP_OP_424J2_126_3477_U392 ( .A(DP_OP_424J2_126_3477_n809), .B(
        DP_OP_424J2_126_3477_n668), .CI(DP_OP_424J2_126_3477_n656), .CO(
        DP_OP_424J2_126_3477_n591), .S(DP_OP_424J2_126_3477_n592) );
  FADDX1_HVT DP_OP_424J2_126_3477_U391 ( .A(DP_OP_424J2_126_3477_n650), .B(
        DP_OP_424J2_126_3477_n648), .CI(DP_OP_424J2_126_3477_n630), .CO(
        DP_OP_424J2_126_3477_n589), .S(DP_OP_424J2_126_3477_n590) );
  FADDX1_HVT DP_OP_424J2_126_3477_U390 ( .A(DP_OP_424J2_126_3477_n646), .B(
        DP_OP_424J2_126_3477_n634), .CI(DP_OP_424J2_126_3477_n628), .CO(
        DP_OP_424J2_126_3477_n587), .S(DP_OP_424J2_126_3477_n588) );
  FADDX1_HVT DP_OP_424J2_126_3477_U389 ( .A(DP_OP_424J2_126_3477_n644), .B(
        DP_OP_424J2_126_3477_n636), .CI(DP_OP_424J2_126_3477_n632), .CO(
        DP_OP_424J2_126_3477_n585), .S(DP_OP_424J2_126_3477_n586) );
  FADDX1_HVT DP_OP_424J2_126_3477_U388 ( .A(DP_OP_424J2_126_3477_n642), .B(
        DP_OP_424J2_126_3477_n640), .CI(DP_OP_424J2_126_3477_n638), .CO(
        DP_OP_424J2_126_3477_n583), .S(DP_OP_424J2_126_3477_n584) );
  FADDX1_HVT DP_OP_424J2_126_3477_U387 ( .A(DP_OP_424J2_126_3477_n626), .B(
        DP_OP_424J2_126_3477_n622), .CI(DP_OP_424J2_126_3477_n624), .CO(
        DP_OP_424J2_126_3477_n581), .S(DP_OP_424J2_126_3477_n582) );
  FADDX1_HVT DP_OP_424J2_126_3477_U386 ( .A(DP_OP_424J2_126_3477_n799), .B(
        DP_OP_424J2_126_3477_n795), .CI(DP_OP_424J2_126_3477_n797), .CO(
        DP_OP_424J2_126_3477_n579), .S(DP_OP_424J2_126_3477_n580) );
  FADDX1_HVT DP_OP_424J2_126_3477_U385 ( .A(DP_OP_424J2_126_3477_n793), .B(
        DP_OP_424J2_126_3477_n787), .CI(DP_OP_424J2_126_3477_n789), .CO(
        DP_OP_424J2_126_3477_n577), .S(DP_OP_424J2_126_3477_n578) );
  FADDX1_HVT DP_OP_424J2_126_3477_U384 ( .A(DP_OP_424J2_126_3477_n791), .B(
        DP_OP_424J2_126_3477_n620), .CI(DP_OP_424J2_126_3477_n785), .CO(
        DP_OP_424J2_126_3477_n575), .S(DP_OP_424J2_126_3477_n576) );
  FADDX1_HVT DP_OP_424J2_126_3477_U383 ( .A(DP_OP_424J2_126_3477_n783), .B(
        DP_OP_424J2_126_3477_n771), .CI(DP_OP_424J2_126_3477_n612), .CO(
        DP_OP_424J2_126_3477_n573), .S(DP_OP_424J2_126_3477_n574) );
  FADDX1_HVT DP_OP_424J2_126_3477_U382 ( .A(DP_OP_424J2_126_3477_n781), .B(
        DP_OP_424J2_126_3477_n618), .CI(DP_OP_424J2_126_3477_n616), .CO(
        DP_OP_424J2_126_3477_n571), .S(DP_OP_424J2_126_3477_n572) );
  FADDX1_HVT DP_OP_424J2_126_3477_U381 ( .A(DP_OP_424J2_126_3477_n779), .B(
        DP_OP_424J2_126_3477_n769), .CI(DP_OP_424J2_126_3477_n614), .CO(
        DP_OP_424J2_126_3477_n569), .S(DP_OP_424J2_126_3477_n570) );
  FADDX1_HVT DP_OP_424J2_126_3477_U380 ( .A(DP_OP_424J2_126_3477_n777), .B(
        DP_OP_424J2_126_3477_n775), .CI(DP_OP_424J2_126_3477_n773), .CO(
        DP_OP_424J2_126_3477_n567), .S(DP_OP_424J2_126_3477_n568) );
  FADDX1_HVT DP_OP_424J2_126_3477_U379 ( .A(DP_OP_424J2_126_3477_n610), .B(
        DP_OP_424J2_126_3477_n767), .CI(DP_OP_424J2_126_3477_n606), .CO(
        DP_OP_424J2_126_3477_n565), .S(DP_OP_424J2_126_3477_n566) );
  FADDX1_HVT DP_OP_424J2_126_3477_U378 ( .A(DP_OP_424J2_126_3477_n765), .B(
        DP_OP_424J2_126_3477_n608), .CI(DP_OP_424J2_126_3477_n763), .CO(
        DP_OP_424J2_126_3477_n563), .S(DP_OP_424J2_126_3477_n564) );
  FADDX1_HVT DP_OP_424J2_126_3477_U377 ( .A(DP_OP_424J2_126_3477_n761), .B(
        DP_OP_424J2_126_3477_n592), .CI(DP_OP_424J2_126_3477_n755), .CO(
        DP_OP_424J2_126_3477_n561), .S(DP_OP_424J2_126_3477_n562) );
  FADDX1_HVT DP_OP_424J2_126_3477_U376 ( .A(DP_OP_424J2_126_3477_n602), .B(
        DP_OP_424J2_126_3477_n757), .CI(DP_OP_424J2_126_3477_n598), .CO(
        DP_OP_424J2_126_3477_n559), .S(DP_OP_424J2_126_3477_n560) );
  FADDX1_HVT DP_OP_424J2_126_3477_U375 ( .A(DP_OP_424J2_126_3477_n604), .B(
        DP_OP_424J2_126_3477_n594), .CI(DP_OP_424J2_126_3477_n596), .CO(
        DP_OP_424J2_126_3477_n557), .S(DP_OP_424J2_126_3477_n558) );
  FADDX1_HVT DP_OP_424J2_126_3477_U374 ( .A(DP_OP_424J2_126_3477_n759), .B(
        DP_OP_424J2_126_3477_n600), .CI(DP_OP_424J2_126_3477_n590), .CO(
        DP_OP_424J2_126_3477_n555), .S(DP_OP_424J2_126_3477_n556) );
  FADDX1_HVT DP_OP_424J2_126_3477_U373 ( .A(DP_OP_424J2_126_3477_n588), .B(
        DP_OP_424J2_126_3477_n584), .CI(DP_OP_424J2_126_3477_n753), .CO(
        DP_OP_424J2_126_3477_n553), .S(DP_OP_424J2_126_3477_n554) );
  FADDX1_HVT DP_OP_424J2_126_3477_U372 ( .A(DP_OP_424J2_126_3477_n586), .B(
        DP_OP_424J2_126_3477_n751), .CI(DP_OP_424J2_126_3477_n582), .CO(
        DP_OP_424J2_126_3477_n551), .S(DP_OP_424J2_126_3477_n552) );
  FADDX1_HVT DP_OP_424J2_126_3477_U371 ( .A(DP_OP_424J2_126_3477_n749), .B(
        DP_OP_424J2_126_3477_n745), .CI(DP_OP_424J2_126_3477_n580), .CO(
        DP_OP_424J2_126_3477_n549), .S(DP_OP_424J2_126_3477_n550) );
  FADDX1_HVT DP_OP_424J2_126_3477_U370 ( .A(DP_OP_424J2_126_3477_n747), .B(
        DP_OP_424J2_126_3477_n743), .CI(DP_OP_424J2_126_3477_n739), .CO(
        DP_OP_424J2_126_3477_n547), .S(DP_OP_424J2_126_3477_n548) );
  FADDX1_HVT DP_OP_424J2_126_3477_U369 ( .A(DP_OP_424J2_126_3477_n741), .B(
        DP_OP_424J2_126_3477_n578), .CI(DP_OP_424J2_126_3477_n576), .CO(
        DP_OP_424J2_126_3477_n545), .S(DP_OP_424J2_126_3477_n546) );
  FADDX1_HVT DP_OP_424J2_126_3477_U368 ( .A(DP_OP_424J2_126_3477_n737), .B(
        DP_OP_424J2_126_3477_n570), .CI(DP_OP_424J2_126_3477_n568), .CO(
        DP_OP_424J2_126_3477_n543), .S(DP_OP_424J2_126_3477_n544) );
  FADDX1_HVT DP_OP_424J2_126_3477_U367 ( .A(DP_OP_424J2_126_3477_n735), .B(
        DP_OP_424J2_126_3477_n572), .CI(DP_OP_424J2_126_3477_n731), .CO(
        DP_OP_424J2_126_3477_n541), .S(DP_OP_424J2_126_3477_n542) );
  FADDX1_HVT DP_OP_424J2_126_3477_U366 ( .A(DP_OP_424J2_126_3477_n733), .B(
        DP_OP_424J2_126_3477_n574), .CI(DP_OP_424J2_126_3477_n729), .CO(
        DP_OP_424J2_126_3477_n539), .S(DP_OP_424J2_126_3477_n540) );
  FADDX1_HVT DP_OP_424J2_126_3477_U365 ( .A(DP_OP_424J2_126_3477_n566), .B(
        DP_OP_424J2_126_3477_n564), .CI(DP_OP_424J2_126_3477_n727), .CO(
        DP_OP_424J2_126_3477_n537), .S(DP_OP_424J2_126_3477_n538) );
  FADDX1_HVT DP_OP_424J2_126_3477_U364 ( .A(DP_OP_424J2_126_3477_n560), .B(
        DP_OP_424J2_126_3477_n556), .CI(DP_OP_424J2_126_3477_n723), .CO(
        DP_OP_424J2_126_3477_n535), .S(DP_OP_424J2_126_3477_n536) );
  FADDX1_HVT DP_OP_424J2_126_3477_U363 ( .A(DP_OP_424J2_126_3477_n558), .B(
        DP_OP_424J2_126_3477_n562), .CI(DP_OP_424J2_126_3477_n725), .CO(
        DP_OP_424J2_126_3477_n533), .S(DP_OP_424J2_126_3477_n534) );
  FADDX1_HVT DP_OP_424J2_126_3477_U362 ( .A(DP_OP_424J2_126_3477_n721), .B(
        DP_OP_424J2_126_3477_n554), .CI(DP_OP_424J2_126_3477_n552), .CO(
        DP_OP_424J2_126_3477_n531), .S(DP_OP_424J2_126_3477_n532) );
  FADDX1_HVT DP_OP_424J2_126_3477_U361 ( .A(DP_OP_424J2_126_3477_n719), .B(
        DP_OP_424J2_126_3477_n717), .CI(DP_OP_424J2_126_3477_n550), .CO(
        DP_OP_424J2_126_3477_n529), .S(DP_OP_424J2_126_3477_n530) );
  FADDX1_HVT DP_OP_424J2_126_3477_U360 ( .A(DP_OP_424J2_126_3477_n715), .B(
        DP_OP_424J2_126_3477_n713), .CI(DP_OP_424J2_126_3477_n548), .CO(
        DP_OP_424J2_126_3477_n527), .S(DP_OP_424J2_126_3477_n528) );
  FADDX1_HVT DP_OP_424J2_126_3477_U359 ( .A(DP_OP_424J2_126_3477_n711), .B(
        DP_OP_424J2_126_3477_n546), .CI(DP_OP_424J2_126_3477_n709), .CO(
        DP_OP_424J2_126_3477_n525), .S(DP_OP_424J2_126_3477_n526) );
  FADDX1_HVT DP_OP_424J2_126_3477_U358 ( .A(DP_OP_424J2_126_3477_n544), .B(
        DP_OP_424J2_126_3477_n542), .CI(DP_OP_424J2_126_3477_n540), .CO(
        DP_OP_424J2_126_3477_n523), .S(DP_OP_424J2_126_3477_n524) );
  FADDX1_HVT DP_OP_424J2_126_3477_U357 ( .A(DP_OP_424J2_126_3477_n707), .B(
        DP_OP_424J2_126_3477_n705), .CI(DP_OP_424J2_126_3477_n538), .CO(
        DP_OP_424J2_126_3477_n521), .S(DP_OP_424J2_126_3477_n522) );
  FADDX1_HVT DP_OP_424J2_126_3477_U356 ( .A(DP_OP_424J2_126_3477_n703), .B(
        DP_OP_424J2_126_3477_n534), .CI(DP_OP_424J2_126_3477_n536), .CO(
        DP_OP_424J2_126_3477_n519), .S(DP_OP_424J2_126_3477_n520) );
  FADDX1_HVT DP_OP_424J2_126_3477_U355 ( .A(DP_OP_424J2_126_3477_n701), .B(
        DP_OP_424J2_126_3477_n532), .CI(DP_OP_424J2_126_3477_n699), .CO(
        DP_OP_424J2_126_3477_n517), .S(DP_OP_424J2_126_3477_n518) );
  FADDX1_HVT DP_OP_424J2_126_3477_U354 ( .A(DP_OP_424J2_126_3477_n697), .B(
        DP_OP_424J2_126_3477_n530), .CI(DP_OP_424J2_126_3477_n695), .CO(
        DP_OP_424J2_126_3477_n515), .S(DP_OP_424J2_126_3477_n516) );
  FADDX1_HVT DP_OP_424J2_126_3477_U353 ( .A(DP_OP_424J2_126_3477_n528), .B(
        DP_OP_424J2_126_3477_n693), .CI(DP_OP_424J2_126_3477_n526), .CO(
        DP_OP_424J2_126_3477_n513), .S(DP_OP_424J2_126_3477_n514) );
  FADDX1_HVT DP_OP_424J2_126_3477_U352 ( .A(DP_OP_424J2_126_3477_n524), .B(
        DP_OP_424J2_126_3477_n691), .CI(DP_OP_424J2_126_3477_n522), .CO(
        DP_OP_424J2_126_3477_n511), .S(DP_OP_424J2_126_3477_n512) );
  FADDX1_HVT DP_OP_424J2_126_3477_U351 ( .A(DP_OP_424J2_126_3477_n689), .B(
        DP_OP_424J2_126_3477_n520), .CI(DP_OP_424J2_126_3477_n687), .CO(
        DP_OP_424J2_126_3477_n509), .S(DP_OP_424J2_126_3477_n510) );
  FADDX1_HVT DP_OP_424J2_126_3477_U350 ( .A(DP_OP_424J2_126_3477_n518), .B(
        DP_OP_424J2_126_3477_n685), .CI(DP_OP_424J2_126_3477_n516), .CO(
        DP_OP_424J2_126_3477_n507), .S(DP_OP_424J2_126_3477_n508) );
  FADDX1_HVT DP_OP_424J2_126_3477_U349 ( .A(DP_OP_424J2_126_3477_n683), .B(
        DP_OP_424J2_126_3477_n514), .CI(DP_OP_424J2_126_3477_n512), .CO(
        DP_OP_424J2_126_3477_n505), .S(DP_OP_424J2_126_3477_n506) );
  FADDX1_HVT DP_OP_424J2_126_3477_U348 ( .A(DP_OP_424J2_126_3477_n681), .B(
        DP_OP_424J2_126_3477_n510), .CI(DP_OP_424J2_126_3477_n679), .CO(
        DP_OP_424J2_126_3477_n503), .S(DP_OP_424J2_126_3477_n504) );
  FADDX1_HVT DP_OP_424J2_126_3477_U347 ( .A(DP_OP_424J2_126_3477_n508), .B(
        DP_OP_424J2_126_3477_n677), .CI(DP_OP_424J2_126_3477_n506), .CO(
        DP_OP_424J2_126_3477_n501), .S(DP_OP_424J2_126_3477_n502) );
  FADDX1_HVT DP_OP_424J2_126_3477_U346 ( .A(DP_OP_424J2_126_3477_n675), .B(
        DP_OP_424J2_126_3477_n504), .CI(DP_OP_424J2_126_3477_n502), .CO(
        DP_OP_424J2_126_3477_n499), .S(DP_OP_424J2_126_3477_n500) );
  FADDX1_HVT DP_OP_424J2_126_3477_U345 ( .A(DP_OP_424J2_126_3477_n671), .B(
        DP_OP_424J2_126_3477_n2531), .CI(DP_OP_424J2_126_3477_n2392), .CO(
        DP_OP_424J2_126_3477_n497), .S(DP_OP_424J2_126_3477_n498) );
  FADDX1_HVT DP_OP_424J2_126_3477_U344 ( .A(DP_OP_424J2_126_3477_n2350), .B(
        DP_OP_424J2_126_3477_n1962), .CI(DP_OP_424J2_126_3477_n2443), .CO(
        DP_OP_424J2_126_3477_n495), .S(DP_OP_424J2_126_3477_n496) );
  FADDX1_HVT DP_OP_424J2_126_3477_U343 ( .A(DP_OP_424J2_126_3477_n1999), .B(
        DP_OP_424J2_126_3477_n1823), .CI(DP_OP_424J2_126_3477_n2094), .CO(
        DP_OP_424J2_126_3477_n493), .S(DP_OP_424J2_126_3477_n494) );
  FADDX1_HVT DP_OP_424J2_126_3477_U342 ( .A(DP_OP_424J2_126_3477_n2700), .B(
        DP_OP_424J2_126_3477_n2043), .CI(DP_OP_424J2_126_3477_n2226), .CO(
        DP_OP_424J2_126_3477_n491), .S(DP_OP_424J2_126_3477_n492) );
  FADDX1_HVT DP_OP_424J2_126_3477_U341 ( .A(DP_OP_424J2_126_3477_n1867), .B(
        DP_OP_424J2_126_3477_n2175), .CI(DP_OP_424J2_126_3477_n2575), .CO(
        DP_OP_424J2_126_3477_n489), .S(DP_OP_424J2_126_3477_n490) );
  FADDX1_HVT DP_OP_424J2_126_3477_U340 ( .A(DP_OP_424J2_126_3477_n2087), .B(
        DP_OP_424J2_126_3477_n2524), .CI(DP_OP_424J2_126_3477_n2744), .CO(
        DP_OP_424J2_126_3477_n487), .S(DP_OP_424J2_126_3477_n488) );
  FADDX1_HVT DP_OP_424J2_126_3477_U339 ( .A(DP_OP_424J2_126_3477_n2788), .B(
        DP_OP_424J2_126_3477_n2568), .CI(DP_OP_424J2_126_3477_n1955), .CO(
        DP_OP_424J2_126_3477_n485), .S(DP_OP_424J2_126_3477_n486) );
  FADDX1_HVT DP_OP_424J2_126_3477_U338 ( .A(DP_OP_424J2_126_3477_n2656), .B(
        DP_OP_424J2_126_3477_n2480), .CI(DP_OP_424J2_126_3477_n1911), .CO(
        DP_OP_424J2_126_3477_n483), .S(DP_OP_424J2_126_3477_n484) );
  FADDX1_HVT DP_OP_424J2_126_3477_U337 ( .A(DP_OP_424J2_126_3477_n2307), .B(
        DP_OP_424J2_126_3477_n2876), .CI(DP_OP_424J2_126_3477_n2436), .CO(
        DP_OP_424J2_126_3477_n481), .S(DP_OP_424J2_126_3477_n482) );
  FADDX1_HVT DP_OP_424J2_126_3477_U336 ( .A(DP_OP_424J2_126_3477_n2832), .B(
        DP_OP_424J2_126_3477_n2883), .CI(DP_OP_424J2_126_3477_n2751), .CO(
        DP_OP_424J2_126_3477_n479), .S(DP_OP_424J2_126_3477_n480) );
  FADDX1_HVT DP_OP_424J2_126_3477_U335 ( .A(DP_OP_424J2_126_3477_n2612), .B(
        DP_OP_424J2_126_3477_n2263), .CI(DP_OP_424J2_126_3477_n2839), .CO(
        DP_OP_424J2_126_3477_n477), .S(DP_OP_424J2_126_3477_n478) );
  FADDX1_HVT DP_OP_424J2_126_3477_U334 ( .A(DP_OP_424J2_126_3477_n2131), .B(
        DP_OP_424J2_126_3477_n2138), .CI(DP_OP_424J2_126_3477_n2270), .CO(
        DP_OP_424J2_126_3477_n475), .S(DP_OP_424J2_126_3477_n476) );
  FADDX1_HVT DP_OP_424J2_126_3477_U333 ( .A(DP_OP_424J2_126_3477_n2219), .B(
        DP_OP_424J2_126_3477_n2663), .CI(DP_OP_424J2_126_3477_n2399), .CO(
        DP_OP_424J2_126_3477_n473), .S(DP_OP_424J2_126_3477_n474) );
  FADDX1_HVT DP_OP_424J2_126_3477_U332 ( .A(DP_OP_424J2_126_3477_n2707), .B(
        DP_OP_424J2_126_3477_n2050), .CI(DP_OP_424J2_126_3477_n2006), .CO(
        DP_OP_424J2_126_3477_n471), .S(DP_OP_424J2_126_3477_n472) );
  FADDX1_HVT DP_OP_424J2_126_3477_U331 ( .A(DP_OP_424J2_126_3477_n1779), .B(
        DP_OP_424J2_126_3477_n2314), .CI(DP_OP_424J2_126_3477_n1918), .CO(
        DP_OP_424J2_126_3477_n469), .S(DP_OP_424J2_126_3477_n470) );
  FADDX1_HVT DP_OP_424J2_126_3477_U330 ( .A(DP_OP_424J2_126_3477_n2487), .B(
        DP_OP_424J2_126_3477_n2355), .CI(DP_OP_424J2_126_3477_n2182), .CO(
        DP_OP_424J2_126_3477_n467), .S(DP_OP_424J2_126_3477_n468) );
  FADDX1_HVT DP_OP_424J2_126_3477_U329 ( .A(DP_OP_424J2_126_3477_n2795), .B(
        DP_OP_424J2_126_3477_n1874), .CI(DP_OP_424J2_126_3477_n1830), .CO(
        DP_OP_424J2_126_3477_n465), .S(DP_OP_424J2_126_3477_n466) );
  FADDX1_HVT DP_OP_424J2_126_3477_U328 ( .A(DP_OP_424J2_126_3477_n2619), .B(
        DP_OP_424J2_126_3477_n669), .CI(DP_OP_424J2_126_3477_n667), .CO(
        DP_OP_424J2_126_3477_n463), .S(DP_OP_424J2_126_3477_n464) );
  FADDX1_HVT DP_OP_424J2_126_3477_U327 ( .A(DP_OP_424J2_126_3477_n665), .B(
        DP_OP_424J2_126_3477_n651), .CI(DP_OP_424J2_126_3477_n649), .CO(
        DP_OP_424J2_126_3477_n461), .S(DP_OP_424J2_126_3477_n462) );
  FADDX1_HVT DP_OP_424J2_126_3477_U326 ( .A(DP_OP_424J2_126_3477_n663), .B(
        DP_OP_424J2_126_3477_n653), .CI(DP_OP_424J2_126_3477_n655), .CO(
        DP_OP_424J2_126_3477_n459), .S(DP_OP_424J2_126_3477_n460) );
  FADDX1_HVT DP_OP_424J2_126_3477_U325 ( .A(DP_OP_424J2_126_3477_n661), .B(
        DP_OP_424J2_126_3477_n657), .CI(DP_OP_424J2_126_3477_n659), .CO(
        DP_OP_424J2_126_3477_n457), .S(DP_OP_424J2_126_3477_n458) );
  FADDX1_HVT DP_OP_424J2_126_3477_U324 ( .A(DP_OP_424J2_126_3477_n647), .B(
        DP_OP_424J2_126_3477_n633), .CI(DP_OP_424J2_126_3477_n627), .CO(
        DP_OP_424J2_126_3477_n455), .S(DP_OP_424J2_126_3477_n456) );
  FADDX1_HVT DP_OP_424J2_126_3477_U323 ( .A(DP_OP_424J2_126_3477_n645), .B(
        DP_OP_424J2_126_3477_n635), .CI(DP_OP_424J2_126_3477_n629), .CO(
        DP_OP_424J2_126_3477_n453), .S(DP_OP_424J2_126_3477_n454) );
  FADDX1_HVT DP_OP_424J2_126_3477_U322 ( .A(DP_OP_424J2_126_3477_n643), .B(
        DP_OP_424J2_126_3477_n637), .CI(DP_OP_424J2_126_3477_n631), .CO(
        DP_OP_424J2_126_3477_n451), .S(DP_OP_424J2_126_3477_n452) );
  FADDX1_HVT DP_OP_424J2_126_3477_U321 ( .A(DP_OP_424J2_126_3477_n641), .B(
        DP_OP_424J2_126_3477_n639), .CI(DP_OP_424J2_126_3477_n625), .CO(
        DP_OP_424J2_126_3477_n449), .S(DP_OP_424J2_126_3477_n450) );
  FADDX1_HVT DP_OP_424J2_126_3477_U320 ( .A(DP_OP_424J2_126_3477_n498), .B(
        DP_OP_424J2_126_3477_n621), .CI(DP_OP_424J2_126_3477_n476), .CO(
        DP_OP_424J2_126_3477_n447), .S(DP_OP_424J2_126_3477_n448) );
  FADDX1_HVT DP_OP_424J2_126_3477_U319 ( .A(DP_OP_424J2_126_3477_n496), .B(
        DP_OP_424J2_126_3477_n488), .CI(DP_OP_424J2_126_3477_n623), .CO(
        DP_OP_424J2_126_3477_n445), .S(DP_OP_424J2_126_3477_n446) );
  FADDX1_HVT DP_OP_424J2_126_3477_U318 ( .A(DP_OP_424J2_126_3477_n492), .B(
        DP_OP_424J2_126_3477_n478), .CI(DP_OP_424J2_126_3477_n486), .CO(
        DP_OP_424J2_126_3477_n443), .S(DP_OP_424J2_126_3477_n444) );
  FADDX1_HVT DP_OP_424J2_126_3477_U317 ( .A(DP_OP_424J2_126_3477_n494), .B(
        DP_OP_424J2_126_3477_n490), .CI(DP_OP_424J2_126_3477_n482), .CO(
        DP_OP_424J2_126_3477_n441), .S(DP_OP_424J2_126_3477_n442) );
  FADDX1_HVT DP_OP_424J2_126_3477_U316 ( .A(DP_OP_424J2_126_3477_n484), .B(
        DP_OP_424J2_126_3477_n480), .CI(DP_OP_424J2_126_3477_n474), .CO(
        DP_OP_424J2_126_3477_n439), .S(DP_OP_424J2_126_3477_n440) );
  FADDX1_HVT DP_OP_424J2_126_3477_U315 ( .A(DP_OP_424J2_126_3477_n472), .B(
        DP_OP_424J2_126_3477_n468), .CI(DP_OP_424J2_126_3477_n466), .CO(
        DP_OP_424J2_126_3477_n437), .S(DP_OP_424J2_126_3477_n438) );
  FADDX1_HVT DP_OP_424J2_126_3477_U314 ( .A(DP_OP_424J2_126_3477_n470), .B(
        DP_OP_424J2_126_3477_n619), .CI(DP_OP_424J2_126_3477_n617), .CO(
        DP_OP_424J2_126_3477_n435), .S(DP_OP_424J2_126_3477_n436) );
  FADDX1_HVT DP_OP_424J2_126_3477_U313 ( .A(DP_OP_424J2_126_3477_n615), .B(
        DP_OP_424J2_126_3477_n611), .CI(DP_OP_424J2_126_3477_n609), .CO(
        DP_OP_424J2_126_3477_n433), .S(DP_OP_424J2_126_3477_n434) );
  FADDX1_HVT DP_OP_424J2_126_3477_U312 ( .A(DP_OP_424J2_126_3477_n613), .B(
        DP_OP_424J2_126_3477_n607), .CI(DP_OP_424J2_126_3477_n605), .CO(
        DP_OP_424J2_126_3477_n431), .S(DP_OP_424J2_126_3477_n432) );
  FADDX1_HVT DP_OP_424J2_126_3477_U311 ( .A(DP_OP_424J2_126_3477_n603), .B(
        DP_OP_424J2_126_3477_n591), .CI(DP_OP_424J2_126_3477_n458), .CO(
        DP_OP_424J2_126_3477_n429), .S(DP_OP_424J2_126_3477_n430) );
  FADDX1_HVT DP_OP_424J2_126_3477_U310 ( .A(DP_OP_424J2_126_3477_n601), .B(
        DP_OP_424J2_126_3477_n595), .CI(DP_OP_424J2_126_3477_n462), .CO(
        DP_OP_424J2_126_3477_n427), .S(DP_OP_424J2_126_3477_n428) );
  FADDX1_HVT DP_OP_424J2_126_3477_U309 ( .A(DP_OP_424J2_126_3477_n464), .B(
        DP_OP_424J2_126_3477_n593), .CI(DP_OP_424J2_126_3477_n460), .CO(
        DP_OP_424J2_126_3477_n425), .S(DP_OP_424J2_126_3477_n426) );
  FADDX1_HVT DP_OP_424J2_126_3477_U308 ( .A(DP_OP_424J2_126_3477_n599), .B(
        DP_OP_424J2_126_3477_n597), .CI(DP_OP_424J2_126_3477_n589), .CO(
        DP_OP_424J2_126_3477_n423), .S(DP_OP_424J2_126_3477_n424) );
  FADDX1_HVT DP_OP_424J2_126_3477_U307 ( .A(DP_OP_424J2_126_3477_n454), .B(
        DP_OP_424J2_126_3477_n583), .CI(DP_OP_424J2_126_3477_n450), .CO(
        DP_OP_424J2_126_3477_n421), .S(DP_OP_424J2_126_3477_n422) );
  FADDX1_HVT DP_OP_424J2_126_3477_U306 ( .A(DP_OP_424J2_126_3477_n587), .B(
        DP_OP_424J2_126_3477_n452), .CI(DP_OP_424J2_126_3477_n585), .CO(
        DP_OP_424J2_126_3477_n419), .S(DP_OP_424J2_126_3477_n420) );
  FADDX1_HVT DP_OP_424J2_126_3477_U305 ( .A(DP_OP_424J2_126_3477_n456), .B(
        DP_OP_424J2_126_3477_n581), .CI(DP_OP_424J2_126_3477_n448), .CO(
        DP_OP_424J2_126_3477_n417), .S(DP_OP_424J2_126_3477_n418) );
  FADDX1_HVT DP_OP_424J2_126_3477_U304 ( .A(DP_OP_424J2_126_3477_n446), .B(
        DP_OP_424J2_126_3477_n444), .CI(DP_OP_424J2_126_3477_n440), .CO(
        DP_OP_424J2_126_3477_n415), .S(DP_OP_424J2_126_3477_n416) );
  FADDX1_HVT DP_OP_424J2_126_3477_U303 ( .A(DP_OP_424J2_126_3477_n442), .B(
        DP_OP_424J2_126_3477_n438), .CI(DP_OP_424J2_126_3477_n579), .CO(
        DP_OP_424J2_126_3477_n413), .S(DP_OP_424J2_126_3477_n414) );
  FADDX1_HVT DP_OP_424J2_126_3477_U302 ( .A(DP_OP_424J2_126_3477_n577), .B(
        DP_OP_424J2_126_3477_n575), .CI(DP_OP_424J2_126_3477_n436), .CO(
        DP_OP_424J2_126_3477_n411), .S(DP_OP_424J2_126_3477_n412) );
  FADDX1_HVT DP_OP_424J2_126_3477_U301 ( .A(DP_OP_424J2_126_3477_n573), .B(
        DP_OP_424J2_126_3477_n567), .CI(DP_OP_424J2_126_3477_n434), .CO(
        DP_OP_424J2_126_3477_n409), .S(DP_OP_424J2_126_3477_n410) );
  FADDX1_HVT DP_OP_424J2_126_3477_U300 ( .A(DP_OP_424J2_126_3477_n571), .B(
        DP_OP_424J2_126_3477_n569), .CI(DP_OP_424J2_126_3477_n565), .CO(
        DP_OP_424J2_126_3477_n407), .S(DP_OP_424J2_126_3477_n408) );
  FADDX1_HVT DP_OP_424J2_126_3477_U299 ( .A(DP_OP_424J2_126_3477_n432), .B(
        DP_OP_424J2_126_3477_n563), .CI(DP_OP_424J2_126_3477_n561), .CO(
        DP_OP_424J2_126_3477_n405), .S(DP_OP_424J2_126_3477_n406) );
  FADDX1_HVT DP_OP_424J2_126_3477_U298 ( .A(DP_OP_424J2_126_3477_n557), .B(
        DP_OP_424J2_126_3477_n555), .CI(DP_OP_424J2_126_3477_n424), .CO(
        DP_OP_424J2_126_3477_n403), .S(DP_OP_424J2_126_3477_n404) );
  FADDX1_HVT DP_OP_424J2_126_3477_U297 ( .A(DP_OP_424J2_126_3477_n559), .B(
        DP_OP_424J2_126_3477_n428), .CI(DP_OP_424J2_126_3477_n426), .CO(
        DP_OP_424J2_126_3477_n401), .S(DP_OP_424J2_126_3477_n402) );
  FADDX1_HVT DP_OP_424J2_126_3477_U296 ( .A(DP_OP_424J2_126_3477_n430), .B(
        DP_OP_424J2_126_3477_n553), .CI(DP_OP_424J2_126_3477_n422), .CO(
        DP_OP_424J2_126_3477_n399), .S(DP_OP_424J2_126_3477_n400) );
  FADDX1_HVT DP_OP_424J2_126_3477_U295 ( .A(DP_OP_424J2_126_3477_n420), .B(
        DP_OP_424J2_126_3477_n551), .CI(DP_OP_424J2_126_3477_n418), .CO(
        DP_OP_424J2_126_3477_n397), .S(DP_OP_424J2_126_3477_n398) );
  FADDX1_HVT DP_OP_424J2_126_3477_U294 ( .A(DP_OP_424J2_126_3477_n416), .B(
        DP_OP_424J2_126_3477_n414), .CI(DP_OP_424J2_126_3477_n549), .CO(
        DP_OP_424J2_126_3477_n395), .S(DP_OP_424J2_126_3477_n396) );
  FADDX1_HVT DP_OP_424J2_126_3477_U293 ( .A(DP_OP_424J2_126_3477_n547), .B(
        DP_OP_424J2_126_3477_n545), .CI(DP_OP_424J2_126_3477_n412), .CO(
        DP_OP_424J2_126_3477_n393), .S(DP_OP_424J2_126_3477_n394) );
  FADDX1_HVT DP_OP_424J2_126_3477_U292 ( .A(DP_OP_424J2_126_3477_n543), .B(
        DP_OP_424J2_126_3477_n410), .CI(DP_OP_424J2_126_3477_n408), .CO(
        DP_OP_424J2_126_3477_n391), .S(DP_OP_424J2_126_3477_n392) );
  FADDX1_HVT DP_OP_424J2_126_3477_U291 ( .A(DP_OP_424J2_126_3477_n541), .B(
        DP_OP_424J2_126_3477_n539), .CI(DP_OP_424J2_126_3477_n537), .CO(
        DP_OP_424J2_126_3477_n389), .S(DP_OP_424J2_126_3477_n390) );
  FADDX1_HVT DP_OP_424J2_126_3477_U290 ( .A(DP_OP_424J2_126_3477_n406), .B(
        DP_OP_424J2_126_3477_n535), .CI(DP_OP_424J2_126_3477_n533), .CO(
        DP_OP_424J2_126_3477_n387), .S(DP_OP_424J2_126_3477_n388) );
  FADDX1_HVT DP_OP_424J2_126_3477_U289 ( .A(DP_OP_424J2_126_3477_n404), .B(
        DP_OP_424J2_126_3477_n402), .CI(DP_OP_424J2_126_3477_n400), .CO(
        DP_OP_424J2_126_3477_n385), .S(DP_OP_424J2_126_3477_n386) );
  FADDX1_HVT DP_OP_424J2_126_3477_U288 ( .A(DP_OP_424J2_126_3477_n531), .B(
        DP_OP_424J2_126_3477_n398), .CI(DP_OP_424J2_126_3477_n529), .CO(
        DP_OP_424J2_126_3477_n383), .S(DP_OP_424J2_126_3477_n384) );
  FADDX1_HVT DP_OP_424J2_126_3477_U287 ( .A(DP_OP_424J2_126_3477_n396), .B(
        DP_OP_424J2_126_3477_n527), .CI(DP_OP_424J2_126_3477_n394), .CO(
        DP_OP_424J2_126_3477_n381), .S(DP_OP_424J2_126_3477_n382) );
  FADDX1_HVT DP_OP_424J2_126_3477_U286 ( .A(DP_OP_424J2_126_3477_n525), .B(
        DP_OP_424J2_126_3477_n523), .CI(DP_OP_424J2_126_3477_n392), .CO(
        DP_OP_424J2_126_3477_n379), .S(DP_OP_424J2_126_3477_n380) );
  FADDX1_HVT DP_OP_424J2_126_3477_U285 ( .A(DP_OP_424J2_126_3477_n390), .B(
        DP_OP_424J2_126_3477_n521), .CI(DP_OP_424J2_126_3477_n519), .CO(
        DP_OP_424J2_126_3477_n377), .S(DP_OP_424J2_126_3477_n378) );
  FADDX1_HVT DP_OP_424J2_126_3477_U284 ( .A(DP_OP_424J2_126_3477_n388), .B(
        DP_OP_424J2_126_3477_n386), .CI(DP_OP_424J2_126_3477_n517), .CO(
        DP_OP_424J2_126_3477_n375), .S(DP_OP_424J2_126_3477_n376) );
  FADDX1_HVT DP_OP_424J2_126_3477_U283 ( .A(DP_OP_424J2_126_3477_n384), .B(
        DP_OP_424J2_126_3477_n515), .CI(DP_OP_424J2_126_3477_n382), .CO(
        DP_OP_424J2_126_3477_n373), .S(DP_OP_424J2_126_3477_n374) );
  FADDX1_HVT DP_OP_424J2_126_3477_U282 ( .A(DP_OP_424J2_126_3477_n513), .B(
        DP_OP_424J2_126_3477_n380), .CI(DP_OP_424J2_126_3477_n511), .CO(
        DP_OP_424J2_126_3477_n371), .S(DP_OP_424J2_126_3477_n372) );
  FADDX1_HVT DP_OP_424J2_126_3477_U281 ( .A(DP_OP_424J2_126_3477_n378), .B(
        DP_OP_424J2_126_3477_n509), .CI(DP_OP_424J2_126_3477_n376), .CO(
        DP_OP_424J2_126_3477_n369), .S(DP_OP_424J2_126_3477_n370) );
  FADDX1_HVT DP_OP_424J2_126_3477_U280 ( .A(DP_OP_424J2_126_3477_n507), .B(
        DP_OP_424J2_126_3477_n374), .CI(DP_OP_424J2_126_3477_n505), .CO(
        DP_OP_424J2_126_3477_n367), .S(DP_OP_424J2_126_3477_n368) );
  FADDX1_HVT DP_OP_424J2_126_3477_U279 ( .A(DP_OP_424J2_126_3477_n372), .B(
        DP_OP_424J2_126_3477_n370), .CI(DP_OP_424J2_126_3477_n503), .CO(
        DP_OP_424J2_126_3477_n365), .S(DP_OP_424J2_126_3477_n366) );
  FADDX1_HVT DP_OP_424J2_126_3477_U278 ( .A(DP_OP_424J2_126_3477_n501), .B(
        DP_OP_424J2_126_3477_n368), .CI(DP_OP_424J2_126_3477_n366), .CO(
        DP_OP_424J2_126_3477_n363), .S(DP_OP_424J2_126_3477_n364) );
  FADDX1_HVT DP_OP_424J2_126_3477_U276 ( .A(DP_OP_424J2_126_3477_n2699), .B(
        DP_OP_424J2_126_3477_n1822), .CI(DP_OP_424J2_126_3477_n2391), .CO(
        DP_OP_424J2_126_3477_n359), .S(DP_OP_424J2_126_3477_n360) );
  FADDX1_HVT DP_OP_424J2_126_3477_U275 ( .A(DP_OP_424J2_126_3477_n1998), .B(
        DP_OP_424J2_126_3477_n1778), .CI(DP_OP_424J2_126_3477_n1954), .CO(
        DP_OP_424J2_126_3477_n357), .S(DP_OP_424J2_126_3477_n358) );
  FADDX1_HVT DP_OP_424J2_126_3477_U274 ( .A(DP_OP_424J2_126_3477_n1866), .B(
        DP_OP_424J2_126_3477_n2567), .CI(DP_OP_424J2_126_3477_n2743), .CO(
        DP_OP_424J2_126_3477_n355), .S(DP_OP_424J2_126_3477_n356) );
  FADDX1_HVT DP_OP_424J2_126_3477_U273 ( .A(DP_OP_424J2_126_3477_n2611), .B(
        DP_OP_424J2_126_3477_n1910), .CI(DP_OP_424J2_126_3477_n2042), .CO(
        DP_OP_424J2_126_3477_n353), .S(DP_OP_424J2_126_3477_n354) );
  FADDX1_HVT DP_OP_424J2_126_3477_U272 ( .A(DP_OP_424J2_126_3477_n2086), .B(
        DP_OP_424J2_126_3477_n2174), .CI(DP_OP_424J2_126_3477_n2435), .CO(
        DP_OP_424J2_126_3477_n351), .S(DP_OP_424J2_126_3477_n352) );
  FADDX1_HVT DP_OP_424J2_126_3477_U271 ( .A(DP_OP_424J2_126_3477_n2130), .B(
        DP_OP_424J2_126_3477_n2479), .CI(DP_OP_424J2_126_3477_n2523), .CO(
        DP_OP_424J2_126_3477_n349), .S(DP_OP_424J2_126_3477_n350) );
  FADDX1_HVT DP_OP_424J2_126_3477_U270 ( .A(DP_OP_424J2_126_3477_n2306), .B(
        DP_OP_424J2_126_3477_n2262), .CI(DP_OP_424J2_126_3477_n2875), .CO(
        DP_OP_424J2_126_3477_n347), .S(DP_OP_424J2_126_3477_n348) );
  FADDX1_HVT DP_OP_424J2_126_3477_U269 ( .A(DP_OP_424J2_126_3477_n2787), .B(
        DP_OP_424J2_126_3477_n2655), .CI(DP_OP_424J2_126_3477_n2831), .CO(
        DP_OP_424J2_126_3477_n345), .S(DP_OP_424J2_126_3477_n346) );
  FADDX1_HVT DP_OP_424J2_126_3477_U268 ( .A(DP_OP_424J2_126_3477_n362), .B(
        DP_OP_424J2_126_3477_n2218), .CI(DP_OP_424J2_126_3477_n497), .CO(
        DP_OP_424J2_126_3477_n343), .S(DP_OP_424J2_126_3477_n344) );
  FADDX1_HVT DP_OP_424J2_126_3477_U267 ( .A(DP_OP_424J2_126_3477_n495), .B(
        DP_OP_424J2_126_3477_n477), .CI(DP_OP_424J2_126_3477_n475), .CO(
        DP_OP_424J2_126_3477_n341), .S(DP_OP_424J2_126_3477_n342) );
  FADDX1_HVT DP_OP_424J2_126_3477_U266 ( .A(DP_OP_424J2_126_3477_n493), .B(
        DP_OP_424J2_126_3477_n479), .CI(DP_OP_424J2_126_3477_n481), .CO(
        DP_OP_424J2_126_3477_n339), .S(DP_OP_424J2_126_3477_n340) );
  FADDX1_HVT DP_OP_424J2_126_3477_U265 ( .A(DP_OP_424J2_126_3477_n491), .B(
        DP_OP_424J2_126_3477_n483), .CI(DP_OP_424J2_126_3477_n485), .CO(
        DP_OP_424J2_126_3477_n337), .S(DP_OP_424J2_126_3477_n338) );
  FADDX1_HVT DP_OP_424J2_126_3477_U264 ( .A(DP_OP_424J2_126_3477_n489), .B(
        DP_OP_424J2_126_3477_n487), .CI(DP_OP_424J2_126_3477_n473), .CO(
        DP_OP_424J2_126_3477_n335), .S(DP_OP_424J2_126_3477_n336) );
  FADDX1_HVT DP_OP_424J2_126_3477_U263 ( .A(DP_OP_424J2_126_3477_n471), .B(
        DP_OP_424J2_126_3477_n467), .CI(DP_OP_424J2_126_3477_n465), .CO(
        DP_OP_424J2_126_3477_n333), .S(DP_OP_424J2_126_3477_n334) );
  FADDX1_HVT DP_OP_424J2_126_3477_U262 ( .A(DP_OP_424J2_126_3477_n469), .B(
        DP_OP_424J2_126_3477_n360), .CI(DP_OP_424J2_126_3477_n358), .CO(
        DP_OP_424J2_126_3477_n331), .S(DP_OP_424J2_126_3477_n332) );
  FADDX1_HVT DP_OP_424J2_126_3477_U261 ( .A(DP_OP_424J2_126_3477_n352), .B(
        DP_OP_424J2_126_3477_n346), .CI(DP_OP_424J2_126_3477_n348), .CO(
        DP_OP_424J2_126_3477_n329), .S(DP_OP_424J2_126_3477_n330) );
  FADDX1_HVT DP_OP_424J2_126_3477_U260 ( .A(DP_OP_424J2_126_3477_n350), .B(
        DP_OP_424J2_126_3477_n356), .CI(DP_OP_424J2_126_3477_n354), .CO(
        DP_OP_424J2_126_3477_n327), .S(DP_OP_424J2_126_3477_n328) );
  FADDX1_HVT DP_OP_424J2_126_3477_U259 ( .A(DP_OP_424J2_126_3477_n463), .B(
        DP_OP_424J2_126_3477_n461), .CI(DP_OP_424J2_126_3477_n457), .CO(
        DP_OP_424J2_126_3477_n325), .S(DP_OP_424J2_126_3477_n326) );
  FADDX1_HVT DP_OP_424J2_126_3477_U258 ( .A(DP_OP_424J2_126_3477_n459), .B(
        DP_OP_424J2_126_3477_n455), .CI(DP_OP_424J2_126_3477_n453), .CO(
        DP_OP_424J2_126_3477_n323), .S(DP_OP_424J2_126_3477_n324) );
  FADDX1_HVT DP_OP_424J2_126_3477_U257 ( .A(DP_OP_424J2_126_3477_n451), .B(
        DP_OP_424J2_126_3477_n449), .CI(DP_OP_424J2_126_3477_n344), .CO(
        DP_OP_424J2_126_3477_n321), .S(DP_OP_424J2_126_3477_n322) );
  FADDX1_HVT DP_OP_424J2_126_3477_U256 ( .A(DP_OP_424J2_126_3477_n447), .B(
        DP_OP_424J2_126_3477_n439), .CI(DP_OP_424J2_126_3477_n336), .CO(
        DP_OP_424J2_126_3477_n319), .S(DP_OP_424J2_126_3477_n320) );
  FADDX1_HVT DP_OP_424J2_126_3477_U255 ( .A(DP_OP_424J2_126_3477_n445), .B(
        DP_OP_424J2_126_3477_n338), .CI(DP_OP_424J2_126_3477_n441), .CO(
        DP_OP_424J2_126_3477_n317), .S(DP_OP_424J2_126_3477_n318) );
  FADDX1_HVT DP_OP_424J2_126_3477_U254 ( .A(DP_OP_424J2_126_3477_n342), .B(
        DP_OP_424J2_126_3477_n340), .CI(DP_OP_424J2_126_3477_n443), .CO(
        DP_OP_424J2_126_3477_n315), .S(DP_OP_424J2_126_3477_n316) );
  FADDX1_HVT DP_OP_424J2_126_3477_U253 ( .A(DP_OP_424J2_126_3477_n437), .B(
        DP_OP_424J2_126_3477_n334), .CI(DP_OP_424J2_126_3477_n435), .CO(
        DP_OP_424J2_126_3477_n313), .S(DP_OP_424J2_126_3477_n314) );
  FADDX1_HVT DP_OP_424J2_126_3477_U252 ( .A(DP_OP_424J2_126_3477_n332), .B(
        DP_OP_424J2_126_3477_n328), .CI(DP_OP_424J2_126_3477_n433), .CO(
        DP_OP_424J2_126_3477_n311), .S(DP_OP_424J2_126_3477_n312) );
  FADDX1_HVT DP_OP_424J2_126_3477_U251 ( .A(DP_OP_424J2_126_3477_n330), .B(
        DP_OP_424J2_126_3477_n431), .CI(DP_OP_424J2_126_3477_n429), .CO(
        DP_OP_424J2_126_3477_n309), .S(DP_OP_424J2_126_3477_n310) );
  FADDX1_HVT DP_OP_424J2_126_3477_U250 ( .A(DP_OP_424J2_126_3477_n427), .B(
        DP_OP_424J2_126_3477_n423), .CI(DP_OP_424J2_126_3477_n326), .CO(
        DP_OP_424J2_126_3477_n307), .S(DP_OP_424J2_126_3477_n308) );
  FADDX1_HVT DP_OP_424J2_126_3477_U249 ( .A(DP_OP_424J2_126_3477_n425), .B(
        DP_OP_424J2_126_3477_n324), .CI(DP_OP_424J2_126_3477_n421), .CO(
        DP_OP_424J2_126_3477_n305), .S(DP_OP_424J2_126_3477_n306) );
  FADDX1_HVT DP_OP_424J2_126_3477_U248 ( .A(DP_OP_424J2_126_3477_n419), .B(
        DP_OP_424J2_126_3477_n322), .CI(DP_OP_424J2_126_3477_n417), .CO(
        DP_OP_424J2_126_3477_n303), .S(DP_OP_424J2_126_3477_n304) );
  FADDX1_HVT DP_OP_424J2_126_3477_U247 ( .A(DP_OP_424J2_126_3477_n415), .B(
        DP_OP_424J2_126_3477_n318), .CI(DP_OP_424J2_126_3477_n413), .CO(
        DP_OP_424J2_126_3477_n301), .S(DP_OP_424J2_126_3477_n302) );
  FADDX1_HVT DP_OP_424J2_126_3477_U246 ( .A(DP_OP_424J2_126_3477_n320), .B(
        DP_OP_424J2_126_3477_n316), .CI(DP_OP_424J2_126_3477_n314), .CO(
        DP_OP_424J2_126_3477_n299), .S(DP_OP_424J2_126_3477_n300) );
  FADDX1_HVT DP_OP_424J2_126_3477_U245 ( .A(DP_OP_424J2_126_3477_n411), .B(
        DP_OP_424J2_126_3477_n312), .CI(DP_OP_424J2_126_3477_n409), .CO(
        DP_OP_424J2_126_3477_n297), .S(DP_OP_424J2_126_3477_n298) );
  FADDX1_HVT DP_OP_424J2_126_3477_U244 ( .A(DP_OP_424J2_126_3477_n407), .B(
        DP_OP_424J2_126_3477_n405), .CI(DP_OP_424J2_126_3477_n310), .CO(
        DP_OP_424J2_126_3477_n295), .S(DP_OP_424J2_126_3477_n296) );
  FADDX1_HVT DP_OP_424J2_126_3477_U243 ( .A(DP_OP_424J2_126_3477_n403), .B(
        DP_OP_424J2_126_3477_n308), .CI(DP_OP_424J2_126_3477_n306), .CO(
        DP_OP_424J2_126_3477_n293), .S(DP_OP_424J2_126_3477_n294) );
  FADDX1_HVT DP_OP_424J2_126_3477_U242 ( .A(DP_OP_424J2_126_3477_n401), .B(
        DP_OP_424J2_126_3477_n399), .CI(DP_OP_424J2_126_3477_n304), .CO(
        DP_OP_424J2_126_3477_n291), .S(DP_OP_424J2_126_3477_n292) );
  FADDX1_HVT DP_OP_424J2_126_3477_U241 ( .A(DP_OP_424J2_126_3477_n397), .B(
        DP_OP_424J2_126_3477_n302), .CI(DP_OP_424J2_126_3477_n395), .CO(
        DP_OP_424J2_126_3477_n289), .S(DP_OP_424J2_126_3477_n290) );
  FADDX1_HVT DP_OP_424J2_126_3477_U240 ( .A(DP_OP_424J2_126_3477_n300), .B(
        DP_OP_424J2_126_3477_n393), .CI(DP_OP_424J2_126_3477_n298), .CO(
        DP_OP_424J2_126_3477_n287), .S(DP_OP_424J2_126_3477_n288) );
  FADDX1_HVT DP_OP_424J2_126_3477_U239 ( .A(DP_OP_424J2_126_3477_n391), .B(
        DP_OP_424J2_126_3477_n389), .CI(DP_OP_424J2_126_3477_n296), .CO(
        DP_OP_424J2_126_3477_n285), .S(DP_OP_424J2_126_3477_n286) );
  FADDX1_HVT DP_OP_424J2_126_3477_U238 ( .A(DP_OP_424J2_126_3477_n387), .B(
        DP_OP_424J2_126_3477_n294), .CI(DP_OP_424J2_126_3477_n385), .CO(
        DP_OP_424J2_126_3477_n283), .S(DP_OP_424J2_126_3477_n284) );
  FADDX1_HVT DP_OP_424J2_126_3477_U237 ( .A(DP_OP_424J2_126_3477_n292), .B(
        DP_OP_424J2_126_3477_n383), .CI(DP_OP_424J2_126_3477_n290), .CO(
        DP_OP_424J2_126_3477_n281), .S(DP_OP_424J2_126_3477_n282) );
  FADDX1_HVT DP_OP_424J2_126_3477_U236 ( .A(DP_OP_424J2_126_3477_n381), .B(
        DP_OP_424J2_126_3477_n288), .CI(DP_OP_424J2_126_3477_n379), .CO(
        DP_OP_424J2_126_3477_n279), .S(DP_OP_424J2_126_3477_n280) );
  FADDX1_HVT DP_OP_424J2_126_3477_U235 ( .A(DP_OP_424J2_126_3477_n286), .B(
        DP_OP_424J2_126_3477_n377), .CI(DP_OP_424J2_126_3477_n284), .CO(
        DP_OP_424J2_126_3477_n277), .S(DP_OP_424J2_126_3477_n278) );
  FADDX1_HVT DP_OP_424J2_126_3477_U234 ( .A(DP_OP_424J2_126_3477_n375), .B(
        DP_OP_424J2_126_3477_n282), .CI(DP_OP_424J2_126_3477_n373), .CO(
        DP_OP_424J2_126_3477_n275), .S(DP_OP_424J2_126_3477_n276) );
  FADDX1_HVT DP_OP_424J2_126_3477_U233 ( .A(DP_OP_424J2_126_3477_n280), .B(
        DP_OP_424J2_126_3477_n371), .CI(DP_OP_424J2_126_3477_n278), .CO(
        DP_OP_424J2_126_3477_n273), .S(DP_OP_424J2_126_3477_n274) );
  FADDX1_HVT DP_OP_424J2_126_3477_U232 ( .A(DP_OP_424J2_126_3477_n369), .B(
        DP_OP_424J2_126_3477_n276), .CI(DP_OP_424J2_126_3477_n367), .CO(
        DP_OP_424J2_126_3477_n271), .S(DP_OP_424J2_126_3477_n272) );
  FADDX1_HVT DP_OP_424J2_126_3477_U231 ( .A(DP_OP_424J2_126_3477_n274), .B(
        DP_OP_424J2_126_3477_n365), .CI(DP_OP_424J2_126_3477_n272), .CO(
        DP_OP_424J2_126_3477_n269), .S(DP_OP_424J2_126_3477_n270) );
  FADDX1_HVT DP_OP_424J2_126_3477_U230 ( .A(DP_OP_424J2_126_3477_n361), .B(
        DP_OP_424J2_126_3477_n1777), .CI(DP_OP_424J2_126_3477_n359), .CO(
        DP_OP_424J2_126_3477_n267), .S(DP_OP_424J2_126_3477_n268) );
  FADDX1_HVT DP_OP_424J2_126_3477_U229 ( .A(DP_OP_424J2_126_3477_n357), .B(
        DP_OP_424J2_126_3477_n345), .CI(DP_OP_424J2_126_3477_n355), .CO(
        DP_OP_424J2_126_3477_n265), .S(DP_OP_424J2_126_3477_n266) );
  FADDX1_HVT DP_OP_424J2_126_3477_U228 ( .A(DP_OP_424J2_126_3477_n353), .B(
        DP_OP_424J2_126_3477_n351), .CI(DP_OP_424J2_126_3477_n349), .CO(
        DP_OP_424J2_126_3477_n263), .S(DP_OP_424J2_126_3477_n264) );
  FADDX1_HVT DP_OP_424J2_126_3477_U227 ( .A(DP_OP_424J2_126_3477_n347), .B(
        DP_OP_424J2_126_3477_n343), .CI(DP_OP_424J2_126_3477_n341), .CO(
        DP_OP_424J2_126_3477_n261), .S(DP_OP_424J2_126_3477_n262) );
  FADDX1_HVT DP_OP_424J2_126_3477_U226 ( .A(DP_OP_424J2_126_3477_n339), .B(
        DP_OP_424J2_126_3477_n337), .CI(DP_OP_424J2_126_3477_n335), .CO(
        DP_OP_424J2_126_3477_n259), .S(DP_OP_424J2_126_3477_n260) );
  FADDX1_HVT DP_OP_424J2_126_3477_U225 ( .A(DP_OP_424J2_126_3477_n333), .B(
        DP_OP_424J2_126_3477_n268), .CI(DP_OP_424J2_126_3477_n331), .CO(
        DP_OP_424J2_126_3477_n257), .S(DP_OP_424J2_126_3477_n258) );
  FADDX1_HVT DP_OP_424J2_126_3477_U224 ( .A(DP_OP_424J2_126_3477_n266), .B(
        DP_OP_424J2_126_3477_n327), .CI(DP_OP_424J2_126_3477_n264), .CO(
        DP_OP_424J2_126_3477_n255), .S(DP_OP_424J2_126_3477_n256) );
  FADDX1_HVT DP_OP_424J2_126_3477_U223 ( .A(DP_OP_424J2_126_3477_n329), .B(
        DP_OP_424J2_126_3477_n325), .CI(DP_OP_424J2_126_3477_n323), .CO(
        DP_OP_424J2_126_3477_n253), .S(DP_OP_424J2_126_3477_n254) );
  FADDX1_HVT DP_OP_424J2_126_3477_U222 ( .A(DP_OP_424J2_126_3477_n321), .B(
        DP_OP_424J2_126_3477_n262), .CI(DP_OP_424J2_126_3477_n319), .CO(
        DP_OP_424J2_126_3477_n251), .S(DP_OP_424J2_126_3477_n252) );
  FADDX1_HVT DP_OP_424J2_126_3477_U221 ( .A(DP_OP_424J2_126_3477_n317), .B(
        DP_OP_424J2_126_3477_n315), .CI(DP_OP_424J2_126_3477_n260), .CO(
        DP_OP_424J2_126_3477_n249), .S(DP_OP_424J2_126_3477_n250) );
  FADDX1_HVT DP_OP_424J2_126_3477_U220 ( .A(DP_OP_424J2_126_3477_n313), .B(
        DP_OP_424J2_126_3477_n258), .CI(DP_OP_424J2_126_3477_n311), .CO(
        DP_OP_424J2_126_3477_n247), .S(DP_OP_424J2_126_3477_n248) );
  FADDX1_HVT DP_OP_424J2_126_3477_U219 ( .A(DP_OP_424J2_126_3477_n256), .B(
        DP_OP_424J2_126_3477_n309), .CI(DP_OP_424J2_126_3477_n307), .CO(
        DP_OP_424J2_126_3477_n245), .S(DP_OP_424J2_126_3477_n246) );
  FADDX1_HVT DP_OP_424J2_126_3477_U218 ( .A(DP_OP_424J2_126_3477_n254), .B(
        DP_OP_424J2_126_3477_n305), .CI(DP_OP_424J2_126_3477_n303), .CO(
        DP_OP_424J2_126_3477_n243), .S(DP_OP_424J2_126_3477_n244) );
  FADDX1_HVT DP_OP_424J2_126_3477_U217 ( .A(DP_OP_424J2_126_3477_n252), .B(
        DP_OP_424J2_126_3477_n301), .CI(DP_OP_424J2_126_3477_n250), .CO(
        DP_OP_424J2_126_3477_n241), .S(DP_OP_424J2_126_3477_n242) );
  FADDX1_HVT DP_OP_424J2_126_3477_U216 ( .A(DP_OP_424J2_126_3477_n299), .B(
        DP_OP_424J2_126_3477_n248), .CI(DP_OP_424J2_126_3477_n297), .CO(
        DP_OP_424J2_126_3477_n239), .S(DP_OP_424J2_126_3477_n240) );
  FADDX1_HVT DP_OP_424J2_126_3477_U215 ( .A(DP_OP_424J2_126_3477_n295), .B(
        DP_OP_424J2_126_3477_n246), .CI(DP_OP_424J2_126_3477_n293), .CO(
        DP_OP_424J2_126_3477_n237), .S(DP_OP_424J2_126_3477_n238) );
  FADDX1_HVT DP_OP_424J2_126_3477_U214 ( .A(DP_OP_424J2_126_3477_n291), .B(
        DP_OP_424J2_126_3477_n244), .CI(DP_OP_424J2_126_3477_n289), .CO(
        DP_OP_424J2_126_3477_n235), .S(DP_OP_424J2_126_3477_n236) );
  FADDX1_HVT DP_OP_424J2_126_3477_U213 ( .A(DP_OP_424J2_126_3477_n242), .B(
        DP_OP_424J2_126_3477_n287), .CI(DP_OP_424J2_126_3477_n240), .CO(
        DP_OP_424J2_126_3477_n233), .S(DP_OP_424J2_126_3477_n234) );
  FADDX1_HVT DP_OP_424J2_126_3477_U212 ( .A(DP_OP_424J2_126_3477_n285), .B(
        DP_OP_424J2_126_3477_n238), .CI(DP_OP_424J2_126_3477_n283), .CO(
        DP_OP_424J2_126_3477_n231), .S(DP_OP_424J2_126_3477_n232) );
  FADDX1_HVT DP_OP_424J2_126_3477_U211 ( .A(DP_OP_424J2_126_3477_n281), .B(
        DP_OP_424J2_126_3477_n236), .CI(DP_OP_424J2_126_3477_n234), .CO(
        DP_OP_424J2_126_3477_n229), .S(DP_OP_424J2_126_3477_n230) );
  FADDX1_HVT DP_OP_424J2_126_3477_U210 ( .A(DP_OP_424J2_126_3477_n279), .B(
        DP_OP_424J2_126_3477_n277), .CI(DP_OP_424J2_126_3477_n232), .CO(
        DP_OP_424J2_126_3477_n227), .S(DP_OP_424J2_126_3477_n228) );
  FADDX1_HVT DP_OP_424J2_126_3477_U209 ( .A(DP_OP_424J2_126_3477_n275), .B(
        DP_OP_424J2_126_3477_n230), .CI(DP_OP_424J2_126_3477_n273), .CO(
        DP_OP_424J2_126_3477_n225), .S(DP_OP_424J2_126_3477_n226) );
  FADDX1_HVT DP_OP_424J2_126_3477_U208 ( .A(DP_OP_424J2_126_3477_n228), .B(
        DP_OP_424J2_126_3477_n271), .CI(DP_OP_424J2_126_3477_n226), .CO(
        DP_OP_424J2_126_3477_n223), .S(DP_OP_424J2_126_3477_n224) );
  FADDX1_HVT DP_OP_424J2_126_3477_U207 ( .A(DP_OP_424J2_126_3477_n1776), .B(
        DP_OP_424J2_126_3477_n267), .CI(DP_OP_424J2_126_3477_n265), .CO(
        DP_OP_424J2_126_3477_n221), .S(DP_OP_424J2_126_3477_n222) );
  FADDX1_HVT DP_OP_424J2_126_3477_U206 ( .A(DP_OP_424J2_126_3477_n263), .B(
        DP_OP_424J2_126_3477_n261), .CI(DP_OP_424J2_126_3477_n259), .CO(
        DP_OP_424J2_126_3477_n219), .S(DP_OP_424J2_126_3477_n220) );
  FADDX1_HVT DP_OP_424J2_126_3477_U205 ( .A(DP_OP_424J2_126_3477_n257), .B(
        DP_OP_424J2_126_3477_n222), .CI(DP_OP_424J2_126_3477_n255), .CO(
        DP_OP_424J2_126_3477_n217), .S(DP_OP_424J2_126_3477_n218) );
  FADDX1_HVT DP_OP_424J2_126_3477_U204 ( .A(DP_OP_424J2_126_3477_n253), .B(
        DP_OP_424J2_126_3477_n251), .CI(DP_OP_424J2_126_3477_n220), .CO(
        DP_OP_424J2_126_3477_n215), .S(DP_OP_424J2_126_3477_n216) );
  FADDX1_HVT DP_OP_424J2_126_3477_U203 ( .A(DP_OP_424J2_126_3477_n249), .B(
        DP_OP_424J2_126_3477_n247), .CI(DP_OP_424J2_126_3477_n218), .CO(
        DP_OP_424J2_126_3477_n213), .S(DP_OP_424J2_126_3477_n214) );
  FADDX1_HVT DP_OP_424J2_126_3477_U202 ( .A(DP_OP_424J2_126_3477_n245), .B(
        DP_OP_424J2_126_3477_n243), .CI(DP_OP_424J2_126_3477_n216), .CO(
        DP_OP_424J2_126_3477_n211), .S(DP_OP_424J2_126_3477_n212) );
  FADDX1_HVT DP_OP_424J2_126_3477_U201 ( .A(DP_OP_424J2_126_3477_n241), .B(
        DP_OP_424J2_126_3477_n214), .CI(DP_OP_424J2_126_3477_n239), .CO(
        DP_OP_424J2_126_3477_n209), .S(DP_OP_424J2_126_3477_n210) );
  FADDX1_HVT DP_OP_424J2_126_3477_U200 ( .A(DP_OP_424J2_126_3477_n237), .B(
        DP_OP_424J2_126_3477_n212), .CI(DP_OP_424J2_126_3477_n235), .CO(
        DP_OP_424J2_126_3477_n207), .S(DP_OP_424J2_126_3477_n208) );
  FADDX1_HVT DP_OP_424J2_126_3477_U199 ( .A(DP_OP_424J2_126_3477_n233), .B(
        DP_OP_424J2_126_3477_n210), .CI(DP_OP_424J2_126_3477_n231), .CO(
        DP_OP_424J2_126_3477_n205), .S(DP_OP_424J2_126_3477_n206) );
  FADDX1_HVT DP_OP_424J2_126_3477_U198 ( .A(DP_OP_424J2_126_3477_n208), .B(
        DP_OP_424J2_126_3477_n229), .CI(DP_OP_424J2_126_3477_n206), .CO(
        DP_OP_424J2_126_3477_n203), .S(DP_OP_424J2_126_3477_n204) );
  FADDX1_HVT DP_OP_424J2_126_3477_U197 ( .A(DP_OP_424J2_126_3477_n227), .B(
        DP_OP_424J2_126_3477_n225), .CI(DP_OP_424J2_126_3477_n204), .CO(
        DP_OP_424J2_126_3477_n201), .S(DP_OP_424J2_126_3477_n202) );
  FADDX1_HVT DP_OP_424J2_126_3477_U196 ( .A(DP_OP_424J2_126_3477_n1775), .B(
        DP_OP_424J2_126_3477_n221), .CI(DP_OP_424J2_126_3477_n219), .CO(
        DP_OP_424J2_126_3477_n199), .S(DP_OP_424J2_126_3477_n200) );
  FADDX1_HVT DP_OP_424J2_126_3477_U195 ( .A(DP_OP_424J2_126_3477_n217), .B(
        DP_OP_424J2_126_3477_n200), .CI(DP_OP_424J2_126_3477_n215), .CO(
        DP_OP_424J2_126_3477_n197), .S(DP_OP_424J2_126_3477_n198) );
  FADDX1_HVT DP_OP_424J2_126_3477_U194 ( .A(DP_OP_424J2_126_3477_n213), .B(
        DP_OP_424J2_126_3477_n211), .CI(DP_OP_424J2_126_3477_n198), .CO(
        DP_OP_424J2_126_3477_n195), .S(DP_OP_424J2_126_3477_n196) );
  FADDX1_HVT DP_OP_424J2_126_3477_U193 ( .A(DP_OP_424J2_126_3477_n209), .B(
        DP_OP_424J2_126_3477_n196), .CI(DP_OP_424J2_126_3477_n207), .CO(
        DP_OP_424J2_126_3477_n193), .S(DP_OP_424J2_126_3477_n194) );
  FADDX1_HVT DP_OP_424J2_126_3477_U192 ( .A(DP_OP_424J2_126_3477_n205), .B(
        DP_OP_424J2_126_3477_n194), .CI(DP_OP_424J2_126_3477_n203), .CO(
        DP_OP_424J2_126_3477_n191), .S(DP_OP_424J2_126_3477_n192) );
  FADDX1_HVT DP_OP_424J2_126_3477_U190 ( .A(DP_OP_424J2_126_3477_n190), .B(
        DP_OP_424J2_126_3477_n199), .CI(DP_OP_424J2_126_3477_n197), .CO(
        DP_OP_424J2_126_3477_n187), .S(DP_OP_424J2_126_3477_n188) );
  FADDX1_HVT DP_OP_424J2_126_3477_U189 ( .A(DP_OP_424J2_126_3477_n188), .B(
        DP_OP_424J2_126_3477_n195), .CI(DP_OP_424J2_126_3477_n193), .CO(
        DP_OP_424J2_126_3477_n185), .S(DP_OP_424J2_126_3477_n186) );
  FADDX1_HVT DP_OP_424J2_126_3477_U188 ( .A(DP_OP_424J2_126_3477_n1774), .B(
        DP_OP_424J2_126_3477_n189), .CI(DP_OP_424J2_126_3477_n187), .CO(
        DP_OP_424J2_126_3477_n183), .S(DP_OP_424J2_126_3477_n184) );
  FADDX1_HVT DP_OP_424J2_126_3477_U171 ( .A(DP_OP_424J2_126_3477_n1754), .B(
        DP_OP_424J2_126_3477_n1752), .CI(DP_OP_424J2_126_3477_n1750), .CO(
        DP_OP_424J2_126_3477_n131), .S(n_conv2_sum_c[0]) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U170 ( .A1(DP_OP_424J2_126_3477_n1688), 
        .A2(DP_OP_424J2_126_3477_n1690), .Y(DP_OP_424J2_126_3477_n130) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U169 ( .A1(DP_OP_424J2_126_3477_n1690), .A2(
        DP_OP_424J2_126_3477_n1688), .Y(DP_OP_424J2_126_3477_n129) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U163 ( .A1(DP_OP_424J2_126_3477_n1582), 
        .A2(DP_OP_424J2_126_3477_n1584), .Y(DP_OP_424J2_126_3477_n127) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U155 ( .A1(DP_OP_424J2_126_3477_n1428), 
        .A2(DP_OP_424J2_126_3477_n1430), .Y(DP_OP_424J2_126_3477_n122) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U154 ( .A1(DP_OP_424J2_126_3477_n1430), .A2(
        DP_OP_424J2_126_3477_n1428), .Y(DP_OP_424J2_126_3477_n121) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U149 ( .A1(DP_OP_424J2_126_3477_n1252), 
        .A2(DP_OP_424J2_126_3477_n1254), .Y(DP_OP_424J2_126_3477_n119) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U141 ( .A1(DP_OP_424J2_126_3477_n1064), 
        .A2(DP_OP_424J2_126_3477_n1066), .Y(DP_OP_424J2_126_3477_n114) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U140 ( .A1(DP_OP_424J2_126_3477_n1066), .A2(
        DP_OP_424J2_126_3477_n1064), .Y(DP_OP_424J2_126_3477_n113) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U135 ( .A1(DP_OP_424J2_126_3477_n870), .A2(
        DP_OP_424J2_126_3477_n872), .Y(DP_OP_424J2_126_3477_n111) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U127 ( .A1(DP_OP_424J2_126_3477_n674), .A2(
        DP_OP_424J2_126_3477_n869), .Y(DP_OP_424J2_126_3477_n106) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U126 ( .A1(DP_OP_424J2_126_3477_n869), .A2(
        DP_OP_424J2_126_3477_n674), .Y(DP_OP_424J2_126_3477_n105) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U120 ( .A1(DP_OP_424J2_126_3477_n500), .A2(
        DP_OP_424J2_126_3477_n673), .Y(DP_OP_424J2_126_3477_n102) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U119 ( .A1(DP_OP_424J2_126_3477_n673), .A2(
        DP_OP_424J2_126_3477_n500), .Y(DP_OP_424J2_126_3477_n101) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U114 ( .A1(DP_OP_424J2_126_3477_n364), .A2(
        DP_OP_424J2_126_3477_n499), .Y(DP_OP_424J2_126_3477_n99) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U113 ( .A1(DP_OP_424J2_126_3477_n499), .A2(
        DP_OP_424J2_126_3477_n364), .Y(DP_OP_424J2_126_3477_n98) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U105 ( .A1(DP_OP_424J2_126_3477_n270), .A2(
        DP_OP_424J2_126_3477_n363), .Y(DP_OP_424J2_126_3477_n93) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U104 ( .A1(DP_OP_424J2_126_3477_n363), .A2(
        DP_OP_424J2_126_3477_n270), .Y(DP_OP_424J2_126_3477_n92) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U97 ( .A1(DP_OP_424J2_126_3477_n224), .A2(
        DP_OP_424J2_126_3477_n269), .Y(DP_OP_424J2_126_3477_n88) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U96 ( .A1(DP_OP_424J2_126_3477_n269), .A2(
        DP_OP_424J2_126_3477_n224), .Y(DP_OP_424J2_126_3477_n87) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U92 ( .A1(DP_OP_424J2_126_3477_n87), .A2(
        DP_OP_424J2_126_3477_n92), .Y(DP_OP_424J2_126_3477_n85) );
  AOI21X1_HVT DP_OP_424J2_126_3477_U91 ( .A1(DP_OP_424J2_126_3477_n94), .A2(
        DP_OP_424J2_126_3477_n85), .A3(DP_OP_424J2_126_3477_n86), .Y(
        DP_OP_424J2_126_3477_n84) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U89 ( .A1(DP_OP_424J2_126_3477_n202), .A2(
        DP_OP_424J2_126_3477_n223), .Y(DP_OP_424J2_126_3477_n83) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U88 ( .A1(DP_OP_424J2_126_3477_n223), .A2(
        DP_OP_424J2_126_3477_n202), .Y(DP_OP_424J2_126_3477_n82) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U83 ( .A1(DP_OP_424J2_126_3477_n201), .A2(
        DP_OP_424J2_126_3477_n192), .Y(DP_OP_424J2_126_3477_n80) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U82 ( .A1(DP_OP_424J2_126_3477_n192), .A2(
        DP_OP_424J2_126_3477_n201), .Y(DP_OP_424J2_126_3477_n79) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U78 ( .A1(DP_OP_424J2_126_3477_n79), .A2(
        DP_OP_424J2_126_3477_n82), .Y(DP_OP_424J2_126_3477_n77) );
  AOI21X1_HVT DP_OP_424J2_126_3477_U77 ( .A1(DP_OP_424J2_126_3477_n86), .A2(
        DP_OP_424J2_126_3477_n77), .A3(DP_OP_424J2_126_3477_n78), .Y(
        DP_OP_424J2_126_3477_n76) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U76 ( .A1(DP_OP_424J2_126_3477_n85), .A2(
        DP_OP_424J2_126_3477_n77), .Y(DP_OP_424J2_126_3477_n75) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U72 ( .A1(DP_OP_424J2_126_3477_n191), .A2(
        DP_OP_424J2_126_3477_n186), .Y(DP_OP_424J2_126_3477_n68) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U62 ( .A1(DP_OP_424J2_126_3477_n185), .A2(
        DP_OP_424J2_126_3477_n184), .Y(DP_OP_424J2_126_3477_n65) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U61 ( .A1(DP_OP_424J2_126_3477_n184), .A2(
        DP_OP_424J2_126_3477_n185), .Y(DP_OP_424J2_126_3477_n64) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U54 ( .A1(DP_OP_424J2_126_3477_n183), .A2(
        DP_OP_424J2_126_3477_n182), .Y(DP_OP_424J2_126_3477_n60) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U53 ( .A1(DP_OP_424J2_126_3477_n182), .A2(
        DP_OP_424J2_126_3477_n183), .Y(DP_OP_424J2_126_3477_n59) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U49 ( .A1(DP_OP_424J2_126_3477_n59), .A2(
        DP_OP_424J2_126_3477_n64), .Y(DP_OP_424J2_126_3477_n57) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U47 ( .A1(DP_OP_424J2_126_3477_n69), .A2(
        DP_OP_424J2_126_3477_n57), .Y(DP_OP_424J2_126_3477_n55) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U44 ( .A1(DP_OP_424J2_126_3477_n180), .A2(
        DP_OP_424J2_126_3477_n181), .Y(DP_OP_424J2_126_3477_n53) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U43 ( .A1(DP_OP_424J2_126_3477_n181), .A2(
        DP_OP_424J2_126_3477_n180), .Y(DP_OP_424J2_126_3477_n52) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U39 ( .A1(DP_OP_424J2_126_3477_n52), .A2(
        DP_OP_424J2_126_3477_n55), .Y(DP_OP_424J2_126_3477_n50) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U34 ( .A1(DP_OP_424J2_126_3477_n178), .A2(
        DP_OP_424J2_126_3477_n179), .Y(DP_OP_424J2_126_3477_n46) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U27 ( .A1(DP_OP_424J2_126_3477_n50), .A2(
        DP_OP_424J2_126_3477_n45), .Y(DP_OP_424J2_126_3477_n41) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U24 ( .A1(DP_OP_424J2_126_3477_n176), .A2(
        DP_OP_424J2_126_3477_n177), .Y(DP_OP_424J2_126_3477_n39) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U23 ( .A1(DP_OP_424J2_126_3477_n177), .A2(
        DP_OP_424J2_126_3477_n176), .Y(DP_OP_424J2_126_3477_n38) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U19 ( .A1(DP_OP_424J2_126_3477_n38), .A2(
        DP_OP_424J2_126_3477_n41), .Y(DP_OP_424J2_126_3477_n36) );
  FADDX1_HVT DP_OP_424J2_126_3477_U15 ( .A(DP_OP_424J2_126_3477_n175), .B(
        DP_OP_424J2_126_3477_n174), .CI(DP_OP_424J2_126_3477_n35), .CO(
        DP_OP_424J2_126_3477_n34), .S(n_conv2_sum_c[20]) );
  FADDX1_HVT DP_OP_424J2_126_3477_U14 ( .A(DP_OP_424J2_126_3477_n173), .B(
        DP_OP_424J2_126_3477_n172), .CI(DP_OP_424J2_126_3477_n34), .CO(
        DP_OP_424J2_126_3477_n33), .S(n_conv2_sum_c[21]) );
  FADDX1_HVT DP_OP_424J2_126_3477_U13 ( .A(DP_OP_424J2_126_3477_n171), .B(
        DP_OP_424J2_126_3477_n170), .CI(DP_OP_424J2_126_3477_n33), .CO(
        DP_OP_424J2_126_3477_n32), .S(n_conv2_sum_c[22]) );
  FADDX1_HVT DP_OP_424J2_126_3477_U12 ( .A(DP_OP_424J2_126_3477_n169), .B(
        DP_OP_424J2_126_3477_n168), .CI(DP_OP_424J2_126_3477_n32), .CO(
        DP_OP_424J2_126_3477_n31), .S(n_conv2_sum_c[23]) );
  FADDX1_HVT DP_OP_424J2_126_3477_U11 ( .A(DP_OP_424J2_126_3477_n167), .B(
        DP_OP_424J2_126_3477_n166), .CI(DP_OP_424J2_126_3477_n31), .CO(
        DP_OP_424J2_126_3477_n30), .S(n_conv2_sum_c[24]) );
  FADDX1_HVT DP_OP_424J2_126_3477_U10 ( .A(DP_OP_424J2_126_3477_n165), .B(
        DP_OP_424J2_126_3477_n164), .CI(DP_OP_424J2_126_3477_n30), .CO(
        DP_OP_424J2_126_3477_n29), .S(n_conv2_sum_c[25]) );
  FADDX1_HVT DP_OP_424J2_126_3477_U9 ( .A(DP_OP_424J2_126_3477_n163), .B(
        DP_OP_424J2_126_3477_n162), .CI(DP_OP_424J2_126_3477_n29), .CO(
        DP_OP_424J2_126_3477_n28), .S(n_conv2_sum_c[26]) );
  FADDX1_HVT DP_OP_424J2_126_3477_U8 ( .A(DP_OP_424J2_126_3477_n161), .B(
        DP_OP_424J2_126_3477_n160), .CI(DP_OP_424J2_126_3477_n28), .CO(
        DP_OP_424J2_126_3477_n27), .S(n_conv2_sum_c[27]) );
  FADDX1_HVT DP_OP_424J2_126_3477_U7 ( .A(DP_OP_424J2_126_3477_n159), .B(
        DP_OP_424J2_126_3477_n158), .CI(DP_OP_424J2_126_3477_n27), .CO(
        DP_OP_424J2_126_3477_n26), .S(n_conv2_sum_c[28]) );
  FADDX1_HVT DP_OP_424J2_126_3477_U6 ( .A(DP_OP_424J2_126_3477_n157), .B(
        DP_OP_424J2_126_3477_n156), .CI(DP_OP_424J2_126_3477_n26), .CO(
        DP_OP_424J2_126_3477_n25), .S(n_conv2_sum_c[29]) );
  FADDX1_HVT DP_OP_424J2_126_3477_U5 ( .A(DP_OP_424J2_126_3477_n155), .B(
        DP_OP_424J2_126_3477_n154), .CI(DP_OP_424J2_126_3477_n25), .CO(
        DP_OP_424J2_126_3477_n24), .S(n_conv2_sum_c[30]) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2129 ( .A1(DP_OP_424J2_126_3477_n1942), .A2(
        DP_OP_422J2_124_3477_n2918), .Y(DP_OP_422J2_124_3477_n2899) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2122 ( .A1(DP_OP_422J2_124_3477_n2908), 
        .A2(DP_OP_422J2_124_3477_n2917), .Y(DP_OP_422J2_124_3477_n2892) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2121 ( .A1(DP_OP_423J2_125_3477_n1849), .A2(
        DP_OP_422J2_124_3477_n2917), .Y(DP_OP_422J2_124_3477_n2891) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2114 ( .A1(DP_OP_422J2_124_3477_n2908), 
        .A2(DP_OP_422J2_124_3477_n2916), .Y(DP_OP_422J2_124_3477_n2884) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2113 ( .A1(DP_OP_424J2_126_3477_n1942), .A2(
        DP_OP_422J2_124_3477_n2916), .Y(DP_OP_422J2_124_3477_n2883) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2112 ( .A1(DP_OP_423J2_125_3477_n1856), .A2(
        DP_OP_424J2_126_3477_n2915), .Y(DP_OP_422J2_124_3477_n2882) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2111 ( .A1(DP_OP_422J2_124_3477_n2913), .A2(
        DP_OP_423J2_125_3477_n2910), .Y(DP_OP_422J2_124_3477_n2881) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2110 ( .A1(DP_OP_422J2_124_3477_n2912), .A2(
        DP_OP_423J2_125_3477_n2910), .Y(DP_OP_422J2_124_3477_n2880) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2109 ( .A1(DP_OP_423J2_125_3477_n1853), .A2(
        DP_OP_424J2_126_3477_n2915), .Y(DP_OP_422J2_124_3477_n2879) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2108 ( .A1(DP_OP_425J2_127_3477_n2778), .A2(
        DP_OP_424J2_126_3477_n2915), .Y(DP_OP_422J2_124_3477_n2878) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2107 ( .A1(DP_OP_422J2_124_3477_n2909), .A2(
        DP_OP_423J2_125_3477_n2910), .Y(DP_OP_422J2_124_3477_n2877) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2106 ( .A1(DP_OP_422J2_124_3477_n2908), .A2(
        DP_OP_423J2_125_3477_n2910), .Y(DP_OP_422J2_124_3477_n2876) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2105 ( .A1(DP_OP_423J2_125_3477_n1849), 
        .A2(DP_OP_424J2_126_3477_n2915), .Y(DP_OP_422J2_124_3477_n2875) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2086 ( .A1(DP_OP_422J2_124_3477_n2864), 
        .A2(DP_OP_425J2_127_3477_n2874), .Y(DP_OP_422J2_124_3477_n2856) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2085 ( .A1(DP_OP_423J2_125_3477_n1893), .A2(
        DP_OP_424J2_126_3477_n2874), .Y(DP_OP_422J2_124_3477_n2855) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2078 ( .A1(DP_OP_422J2_124_3477_n2864), 
        .A2(DP_OP_422J2_124_3477_n2873), .Y(DP_OP_422J2_124_3477_n2848) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2077 ( .A1(DP_OP_424J2_126_3477_n1986), .A2(
        DP_OP_422J2_124_3477_n2873), .Y(DP_OP_422J2_124_3477_n2847) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2070 ( .A1(DP_OP_422J2_124_3477_n2864), 
        .A2(DP_OP_422J2_124_3477_n2872), .Y(DP_OP_422J2_124_3477_n2840) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2069 ( .A1(DP_OP_424J2_126_3477_n1986), .A2(
        DP_OP_422J2_124_3477_n2872), .Y(DP_OP_422J2_124_3477_n2839) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2068 ( .A1(DP_OP_422J2_124_3477_n2870), .A2(
        DP_OP_422J2_124_3477_n2871), .Y(DP_OP_422J2_124_3477_n2838) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2067 ( .A1(DP_OP_422J2_124_3477_n2869), .A2(
        DP_OP_422J2_124_3477_n2871), .Y(DP_OP_422J2_124_3477_n2837) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2066 ( .A1(DP_OP_422J2_124_3477_n2868), .A2(
        DP_OP_422J2_124_3477_n2871), .Y(DP_OP_422J2_124_3477_n2836) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2065 ( .A1(DP_OP_423J2_125_3477_n1897), .A2(
        DP_OP_422J2_124_3477_n2871), .Y(DP_OP_422J2_124_3477_n2835) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2064 ( .A1(DP_OP_423J2_125_3477_n1896), .A2(
        DP_OP_422J2_124_3477_n2871), .Y(DP_OP_422J2_124_3477_n2834) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2063 ( .A1(DP_OP_422J2_124_3477_n2865), .A2(
        DP_OP_422J2_124_3477_n2871), .Y(DP_OP_422J2_124_3477_n2833) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2062 ( .A1(DP_OP_422J2_124_3477_n2864), .A2(
        DP_OP_422J2_124_3477_n2871), .Y(DP_OP_422J2_124_3477_n2832) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2061 ( .A1(DP_OP_423J2_125_3477_n1893), 
        .A2(DP_OP_422J2_124_3477_n2871), .Y(DP_OP_422J2_124_3477_n2831) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2041 ( .A1(DP_OP_422J2_124_3477_n2819), .A2(
        DP_OP_422J2_124_3477_n2830), .Y(DP_OP_422J2_124_3477_n2811) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2034 ( .A1(DP_OP_422J2_124_3477_n2820), 
        .A2(DP_OP_423J2_125_3477_n2824), .Y(DP_OP_422J2_124_3477_n2804) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2033 ( .A1(DP_OP_422J2_124_3477_n2819), .A2(
        DP_OP_424J2_126_3477_n2829), .Y(DP_OP_422J2_124_3477_n2803) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2026 ( .A1(DP_OP_422J2_124_3477_n2820), 
        .A2(DP_OP_424J2_126_3477_n2828), .Y(DP_OP_422J2_124_3477_n2796) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2025 ( .A1(DP_OP_422J2_124_3477_n2819), .A2(
        DP_OP_425J2_127_3477_n2828), .Y(DP_OP_422J2_124_3477_n2795) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2024 ( .A1(DP_OP_424J2_126_3477_n2037), .A2(
        DP_OP_422J2_124_3477_n2827), .Y(DP_OP_422J2_124_3477_n2794) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2023 ( .A1(DP_OP_422J2_124_3477_n2825), .A2(
        DP_OP_422J2_124_3477_n2827), .Y(DP_OP_422J2_124_3477_n2793) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2022 ( .A1(DP_OP_424J2_126_3477_n2035), .A2(
        DP_OP_422J2_124_3477_n2827), .Y(DP_OP_422J2_124_3477_n2792) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2021 ( .A1(DP_OP_424J2_126_3477_n2034), .A2(
        DP_OP_422J2_124_3477_n2827), .Y(DP_OP_422J2_124_3477_n2791) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2020 ( .A1(DP_OP_424J2_126_3477_n2033), .A2(
        DP_OP_422J2_124_3477_n2827), .Y(DP_OP_422J2_124_3477_n2790) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2019 ( .A1(DP_OP_424J2_126_3477_n2032), .A2(
        DP_OP_422J2_124_3477_n2827), .Y(DP_OP_422J2_124_3477_n2789) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2018 ( .A1(DP_OP_422J2_124_3477_n2820), .A2(
        DP_OP_422J2_124_3477_n2827), .Y(DP_OP_422J2_124_3477_n2788) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2017 ( .A1(DP_OP_422J2_124_3477_n2819), 
        .A2(DP_OP_422J2_124_3477_n2827), .Y(DP_OP_422J2_124_3477_n2787) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1998 ( .A1(DP_OP_422J2_124_3477_n2776), 
        .A2(DP_OP_422J2_124_3477_n2786), .Y(DP_OP_422J2_124_3477_n2768) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1997 ( .A1(DP_OP_425J2_127_3477_n2643), .A2(
        DP_OP_422J2_124_3477_n2786), .Y(DP_OP_422J2_124_3477_n2767) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1990 ( .A1(DP_OP_422J2_124_3477_n2776), 
        .A2(DP_OP_422J2_124_3477_n2785), .Y(DP_OP_422J2_124_3477_n2760) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1989 ( .A1(DP_OP_425J2_127_3477_n2643), .A2(
        DP_OP_422J2_124_3477_n2785), .Y(DP_OP_422J2_124_3477_n2759) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1982 ( .A1(DP_OP_422J2_124_3477_n2776), 
        .A2(DP_OP_422J2_124_3477_n2784), .Y(DP_OP_422J2_124_3477_n2752) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1981 ( .A1(DP_OP_425J2_127_3477_n2643), .A2(
        DP_OP_422J2_124_3477_n2784), .Y(DP_OP_422J2_124_3477_n2751) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1980 ( .A1(DP_OP_422J2_124_3477_n2782), .A2(
        DP_OP_424J2_126_3477_n2783), .Y(DP_OP_422J2_124_3477_n2750) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1979 ( .A1(DP_OP_422J2_124_3477_n2781), .A2(
        DP_OP_423J2_125_3477_n2778), .Y(DP_OP_422J2_124_3477_n2749) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1978 ( .A1(DP_OP_422J2_124_3477_n2780), .A2(
        DP_OP_423J2_125_3477_n2778), .Y(DP_OP_422J2_124_3477_n2748) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1977 ( .A1(DP_OP_423J2_125_3477_n1985), .A2(
        DP_OP_424J2_126_3477_n2783), .Y(DP_OP_422J2_124_3477_n2747) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1976 ( .A1(DP_OP_424J2_126_3477_n2077), .A2(
        DP_OP_424J2_126_3477_n2783), .Y(DP_OP_422J2_124_3477_n2746) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1975 ( .A1(DP_OP_422J2_124_3477_n2777), .A2(
        DP_OP_424J2_126_3477_n2783), .Y(DP_OP_422J2_124_3477_n2745) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1974 ( .A1(DP_OP_422J2_124_3477_n2776), .A2(
        DP_OP_424J2_126_3477_n2783), .Y(DP_OP_422J2_124_3477_n2744) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1973 ( .A1(DP_OP_424J2_126_3477_n2074), 
        .A2(DP_OP_423J2_125_3477_n2778), .Y(DP_OP_422J2_124_3477_n2743) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1955 ( .A1(DP_OP_422J2_124_3477_n2733), 
        .A2(DP_OP_422J2_124_3477_n2742), .Y(DP_OP_422J2_124_3477_n2725) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1954 ( .A1(DP_OP_422J2_124_3477_n2732), 
        .A2(DP_OP_422J2_124_3477_n2742), .Y(DP_OP_422J2_124_3477_n2724) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1953 ( .A1(DP_OP_422J2_124_3477_n2731), .A2(
        DP_OP_422J2_124_3477_n2742), .Y(DP_OP_422J2_124_3477_n2723) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1945 ( .A1(DP_OP_422J2_124_3477_n2731), .A2(
        DP_OP_422J2_124_3477_n2741), .Y(DP_OP_422J2_124_3477_n2715) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1938 ( .A1(DP_OP_422J2_124_3477_n2732), 
        .A2(DP_OP_422J2_124_3477_n2740), .Y(DP_OP_422J2_124_3477_n2708) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1937 ( .A1(DP_OP_422J2_124_3477_n2731), .A2(
        DP_OP_422J2_124_3477_n2740), .Y(DP_OP_422J2_124_3477_n2707) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1936 ( .A1(DP_OP_424J2_126_3477_n2125), .A2(
        DP_OP_422J2_124_3477_n2739), .Y(DP_OP_422J2_124_3477_n2706) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1935 ( .A1(DP_OP_424J2_126_3477_n2124), .A2(
        DP_OP_422J2_124_3477_n2739), .Y(DP_OP_422J2_124_3477_n2705) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1934 ( .A1(DP_OP_422J2_124_3477_n2736), .A2(
        DP_OP_422J2_124_3477_n2739), .Y(DP_OP_422J2_124_3477_n2704) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1933 ( .A1(DP_OP_422J2_124_3477_n2735), .A2(
        DP_OP_422J2_124_3477_n2739), .Y(DP_OP_422J2_124_3477_n2703) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1932 ( .A1(DP_OP_422J2_124_3477_n2734), .A2(
        DP_OP_422J2_124_3477_n2739), .Y(DP_OP_422J2_124_3477_n2702) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1931 ( .A1(DP_OP_422J2_124_3477_n2733), .A2(
        DP_OP_422J2_124_3477_n2739), .Y(DP_OP_422J2_124_3477_n671) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1930 ( .A1(DP_OP_422J2_124_3477_n2732), .A2(
        DP_OP_422J2_124_3477_n2739), .Y(DP_OP_422J2_124_3477_n2701) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1929 ( .A1(DP_OP_422J2_124_3477_n2731), 
        .A2(DP_OP_422J2_124_3477_n2739), .Y(DP_OP_422J2_124_3477_n361) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1910 ( .A1(DP_OP_422J2_124_3477_n2690), 
        .A2(DP_OP_422J2_124_3477_n2700), .Y(DP_OP_422J2_124_3477_n2682) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1909 ( .A1(DP_OP_422J2_124_3477_n2689), .A2(
        DP_OP_422J2_124_3477_n2700), .Y(DP_OP_422J2_124_3477_n2681) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1902 ( .A1(DP_OP_422J2_124_3477_n2690), 
        .A2(DP_OP_422J2_124_3477_n2699), .Y(DP_OP_422J2_124_3477_n2674) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1901 ( .A1(DP_OP_422J2_124_3477_n2689), .A2(
        DP_OP_422J2_124_3477_n2699), .Y(DP_OP_422J2_124_3477_n2673) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1894 ( .A1(DP_OP_422J2_124_3477_n2690), 
        .A2(DP_OP_422J2_124_3477_n2698), .Y(DP_OP_422J2_124_3477_n2666) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1893 ( .A1(DP_OP_422J2_124_3477_n2689), .A2(
        DP_OP_422J2_124_3477_n2698), .Y(DP_OP_422J2_124_3477_n2665) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1892 ( .A1(DP_OP_422J2_124_3477_n2696), .A2(
        DP_OP_422J2_124_3477_n2697), .Y(DP_OP_422J2_124_3477_n2664) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1891 ( .A1(DP_OP_422J2_124_3477_n2695), .A2(
        DP_OP_422J2_124_3477_n2697), .Y(DP_OP_422J2_124_3477_n2663) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1890 ( .A1(DP_OP_422J2_124_3477_n2694), .A2(
        DP_OP_422J2_124_3477_n2697), .Y(DP_OP_422J2_124_3477_n2662) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1889 ( .A1(DP_OP_425J2_127_3477_n2559), .A2(
        DP_OP_422J2_124_3477_n2697), .Y(DP_OP_422J2_124_3477_n2661) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1888 ( .A1(DP_OP_422J2_124_3477_n2692), .A2(
        DP_OP_422J2_124_3477_n2697), .Y(DP_OP_422J2_124_3477_n2660) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1887 ( .A1(DP_OP_425J2_127_3477_n2557), .A2(
        DP_OP_422J2_124_3477_n2697), .Y(DP_OP_422J2_124_3477_n2659) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1886 ( .A1(DP_OP_422J2_124_3477_n2690), .A2(
        DP_OP_422J2_124_3477_n2697), .Y(DP_OP_422J2_124_3477_n2658) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1885 ( .A1(DP_OP_422J2_124_3477_n2689), 
        .A2(DP_OP_422J2_124_3477_n2697), .Y(DP_OP_422J2_124_3477_n2657) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1866 ( .A1(DP_OP_422J2_124_3477_n2646), 
        .A2(DP_OP_422J2_124_3477_n2656), .Y(DP_OP_422J2_124_3477_n2638) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1865 ( .A1(DP_OP_422J2_124_3477_n2645), .A2(
        DP_OP_422J2_124_3477_n2656), .Y(DP_OP_422J2_124_3477_n2637) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1858 ( .A1(DP_OP_422J2_124_3477_n2646), 
        .A2(DP_OP_422J2_124_3477_n2655), .Y(DP_OP_422J2_124_3477_n2630) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1857 ( .A1(DP_OP_422J2_124_3477_n2645), .A2(
        DP_OP_422J2_124_3477_n2655), .Y(DP_OP_422J2_124_3477_n2629) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1850 ( .A1(DP_OP_422J2_124_3477_n2646), 
        .A2(DP_OP_422J2_124_3477_n2654), .Y(DP_OP_422J2_124_3477_n2622) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1849 ( .A1(DP_OP_422J2_124_3477_n2645), .A2(
        DP_OP_422J2_124_3477_n2654), .Y(DP_OP_422J2_124_3477_n2621) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1848 ( .A1(DP_OP_422J2_124_3477_n2652), .A2(
        DP_OP_422J2_124_3477_n2653), .Y(DP_OP_422J2_124_3477_n2620) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1847 ( .A1(DP_OP_422J2_124_3477_n2651), .A2(
        DP_OP_422J2_124_3477_n2653), .Y(DP_OP_422J2_124_3477_n2619) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1846 ( .A1(DP_OP_422J2_124_3477_n2650), .A2(
        DP_OP_422J2_124_3477_n2653), .Y(DP_OP_422J2_124_3477_n2618) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1845 ( .A1(DP_OP_422J2_124_3477_n2649), .A2(
        DP_OP_422J2_124_3477_n2653), .Y(DP_OP_422J2_124_3477_n2617) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1844 ( .A1(DP_OP_422J2_124_3477_n2648), .A2(
        DP_OP_422J2_124_3477_n2653), .Y(DP_OP_422J2_124_3477_n2616) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1843 ( .A1(DP_OP_422J2_124_3477_n2647), .A2(
        DP_OP_422J2_124_3477_n2653), .Y(DP_OP_422J2_124_3477_n2615) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1842 ( .A1(DP_OP_422J2_124_3477_n2646), .A2(
        DP_OP_422J2_124_3477_n2653), .Y(DP_OP_422J2_124_3477_n2614) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1841 ( .A1(DP_OP_422J2_124_3477_n2645), 
        .A2(DP_OP_422J2_124_3477_n2653), .Y(DP_OP_422J2_124_3477_n2613) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1822 ( .A1(DP_OP_422J2_124_3477_n2602), 
        .A2(DP_OP_422J2_124_3477_n2612), .Y(DP_OP_422J2_124_3477_n2594) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1821 ( .A1(DP_OP_422J2_124_3477_n2601), .A2(
        DP_OP_422J2_124_3477_n2612), .Y(DP_OP_422J2_124_3477_n2593) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1814 ( .A1(DP_OP_422J2_124_3477_n2602), 
        .A2(DP_OP_422J2_124_3477_n2611), .Y(DP_OP_422J2_124_3477_n2586) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1813 ( .A1(DP_OP_422J2_124_3477_n2601), .A2(
        DP_OP_422J2_124_3477_n2611), .Y(DP_OP_422J2_124_3477_n2585) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1806 ( .A1(DP_OP_422J2_124_3477_n2602), 
        .A2(DP_OP_422J2_124_3477_n2610), .Y(DP_OP_422J2_124_3477_n2578) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1805 ( .A1(DP_OP_422J2_124_3477_n2601), .A2(
        DP_OP_422J2_124_3477_n2610), .Y(DP_OP_422J2_124_3477_n2577) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1804 ( .A1(DP_OP_422J2_124_3477_n2608), .A2(
        DP_OP_422J2_124_3477_n2609), .Y(DP_OP_422J2_124_3477_n2576) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1803 ( .A1(DP_OP_422J2_124_3477_n2607), .A2(
        DP_OP_422J2_124_3477_n2609), .Y(DP_OP_422J2_124_3477_n2575) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1802 ( .A1(DP_OP_422J2_124_3477_n2606), .A2(
        DP_OP_422J2_124_3477_n2609), .Y(DP_OP_422J2_124_3477_n2574) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1801 ( .A1(DP_OP_422J2_124_3477_n2605), .A2(
        DP_OP_422J2_124_3477_n2609), .Y(DP_OP_422J2_124_3477_n2573) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1800 ( .A1(DP_OP_422J2_124_3477_n2604), .A2(
        DP_OP_422J2_124_3477_n2609), .Y(DP_OP_422J2_124_3477_n2572) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1799 ( .A1(DP_OP_422J2_124_3477_n2603), .A2(
        DP_OP_422J2_124_3477_n2609), .Y(DP_OP_422J2_124_3477_n2571) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1798 ( .A1(DP_OP_422J2_124_3477_n2602), .A2(
        DP_OP_422J2_124_3477_n2609), .Y(DP_OP_422J2_124_3477_n2570) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1797 ( .A1(DP_OP_422J2_124_3477_n2601), 
        .A2(DP_OP_422J2_124_3477_n2609), .Y(DP_OP_422J2_124_3477_n2569) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1778 ( .A1(DP_OP_422J2_124_3477_n2558), 
        .A2(DP_OP_422J2_124_3477_n2568), .Y(DP_OP_422J2_124_3477_n2550) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1777 ( .A1(DP_OP_422J2_124_3477_n2557), .A2(
        DP_OP_422J2_124_3477_n2568), .Y(DP_OP_422J2_124_3477_n2549) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1769 ( .A1(DP_OP_422J2_124_3477_n2557), .A2(
        DP_OP_422J2_124_3477_n2567), .Y(DP_OP_422J2_124_3477_n2541) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1761 ( .A1(DP_OP_422J2_124_3477_n2557), .A2(
        DP_OP_422J2_124_3477_n2566), .Y(DP_OP_422J2_124_3477_n2533) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1760 ( .A1(DP_OP_422J2_124_3477_n2564), .A2(
        DP_OP_424J2_126_3477_n2563), .Y(DP_OP_422J2_124_3477_n2532) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1759 ( .A1(DP_OP_422J2_124_3477_n2563), .A2(
        DP_OP_423J2_125_3477_n2561), .Y(DP_OP_422J2_124_3477_n2531) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1758 ( .A1(DP_OP_422J2_124_3477_n2562), .A2(
        DP_OP_424J2_126_3477_n2563), .Y(DP_OP_422J2_124_3477_n2530) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1757 ( .A1(DP_OP_423J2_125_3477_n2205), .A2(
        DP_OP_424J2_126_3477_n2563), .Y(DP_OP_422J2_124_3477_n2529) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1756 ( .A1(DP_OP_422J2_124_3477_n2560), .A2(
        DP_OP_424J2_126_3477_n2563), .Y(DP_OP_422J2_124_3477_n2528) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1755 ( .A1(DP_OP_422J2_124_3477_n2559), .A2(
        DP_OP_424J2_126_3477_n2563), .Y(DP_OP_422J2_124_3477_n2527) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1754 ( .A1(DP_OP_422J2_124_3477_n2558), .A2(
        DP_OP_423J2_125_3477_n2561), .Y(DP_OP_422J2_124_3477_n2526) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1753 ( .A1(DP_OP_422J2_124_3477_n2557), 
        .A2(DP_OP_423J2_125_3477_n2561), .Y(DP_OP_422J2_124_3477_n2525) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1734 ( .A1(DP_OP_422J2_124_3477_n2514), 
        .A2(DP_OP_422J2_124_3477_n2524), .Y(DP_OP_422J2_124_3477_n2506) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1733 ( .A1(DP_OP_422J2_124_3477_n2513), .A2(
        DP_OP_422J2_124_3477_n2524), .Y(DP_OP_422J2_124_3477_n2505) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1725 ( .A1(DP_OP_422J2_124_3477_n2513), .A2(
        DP_OP_422J2_124_3477_n2523), .Y(DP_OP_422J2_124_3477_n2497) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1718 ( .A1(DP_OP_422J2_124_3477_n2514), 
        .A2(DP_OP_422J2_124_3477_n2522), .Y(DP_OP_422J2_124_3477_n2490) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1717 ( .A1(DP_OP_422J2_124_3477_n2513), .A2(
        DP_OP_422J2_124_3477_n2522), .Y(DP_OP_422J2_124_3477_n2489) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1716 ( .A1(DP_OP_422J2_124_3477_n2520), .A2(
        DP_OP_422J2_124_3477_n2521), .Y(DP_OP_422J2_124_3477_n2488) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1715 ( .A1(DP_OP_424J2_126_3477_n2344), .A2(
        DP_OP_422J2_124_3477_n2521), .Y(DP_OP_422J2_124_3477_n2487) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1714 ( .A1(DP_OP_422J2_124_3477_n2518), .A2(
        DP_OP_422J2_124_3477_n2521), .Y(DP_OP_422J2_124_3477_n2486) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1713 ( .A1(DP_OP_424J2_126_3477_n2342), .A2(
        DP_OP_422J2_124_3477_n2521), .Y(DP_OP_422J2_124_3477_n2485) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1712 ( .A1(DP_OP_424J2_126_3477_n2341), .A2(
        DP_OP_422J2_124_3477_n2521), .Y(DP_OP_422J2_124_3477_n2484) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1711 ( .A1(DP_OP_423J2_125_3477_n2247), .A2(
        DP_OP_422J2_124_3477_n2521), .Y(DP_OP_422J2_124_3477_n2483) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1710 ( .A1(DP_OP_422J2_124_3477_n2514), .A2(
        DP_OP_422J2_124_3477_n2521), .Y(DP_OP_422J2_124_3477_n2482) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1709 ( .A1(DP_OP_422J2_124_3477_n2513), 
        .A2(DP_OP_422J2_124_3477_n2521), .Y(DP_OP_422J2_124_3477_n2481) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1690 ( .A1(DP_OP_422J2_124_3477_n2470), 
        .A2(DP_OP_422J2_124_3477_n2480), .Y(DP_OP_422J2_124_3477_n2462) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1689 ( .A1(DP_OP_422J2_124_3477_n2469), .A2(
        DP_OP_422J2_124_3477_n2480), .Y(DP_OP_422J2_124_3477_n2461) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1682 ( .A1(DP_OP_422J2_124_3477_n2470), 
        .A2(DP_OP_422J2_124_3477_n2479), .Y(DP_OP_422J2_124_3477_n2454) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1681 ( .A1(DP_OP_422J2_124_3477_n2469), .A2(
        DP_OP_422J2_124_3477_n2479), .Y(DP_OP_422J2_124_3477_n2453) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1674 ( .A1(DP_OP_422J2_124_3477_n2470), 
        .A2(DP_OP_422J2_124_3477_n2478), .Y(DP_OP_422J2_124_3477_n2446) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1673 ( .A1(DP_OP_422J2_124_3477_n2469), .A2(
        DP_OP_422J2_124_3477_n2478), .Y(DP_OP_422J2_124_3477_n2445) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1672 ( .A1(DP_OP_422J2_124_3477_n2476), .A2(
        DP_OP_422J2_124_3477_n2477), .Y(DP_OP_422J2_124_3477_n2444) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1671 ( .A1(DP_OP_423J2_125_3477_n2295), .A2(
        DP_OP_422J2_124_3477_n2477), .Y(DP_OP_422J2_124_3477_n2443) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1670 ( .A1(DP_OP_423J2_125_3477_n2294), .A2(
        DP_OP_422J2_124_3477_n2477), .Y(DP_OP_422J2_124_3477_n2442) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1669 ( .A1(DP_OP_422J2_124_3477_n2473), .A2(
        DP_OP_422J2_124_3477_n2477), .Y(DP_OP_422J2_124_3477_n2441) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1668 ( .A1(DP_OP_422J2_124_3477_n2472), .A2(
        DP_OP_422J2_124_3477_n2477), .Y(DP_OP_422J2_124_3477_n2440) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1667 ( .A1(DP_OP_423J2_125_3477_n2291), .A2(
        DP_OP_422J2_124_3477_n2477), .Y(DP_OP_422J2_124_3477_n2439) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1666 ( .A1(DP_OP_422J2_124_3477_n2470), .A2(
        DP_OP_422J2_124_3477_n2477), .Y(DP_OP_422J2_124_3477_n2438) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1665 ( .A1(DP_OP_422J2_124_3477_n2469), 
        .A2(DP_OP_422J2_124_3477_n2477), .Y(DP_OP_422J2_124_3477_n2437) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1646 ( .A1(DP_OP_423J2_125_3477_n2334), 
        .A2(DP_OP_422J2_124_3477_n2436), .Y(DP_OP_422J2_124_3477_n2418) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1645 ( .A1(DP_OP_423J2_125_3477_n2333), .A2(
        DP_OP_422J2_124_3477_n2436), .Y(DP_OP_422J2_124_3477_n2417) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1638 ( .A1(DP_OP_423J2_125_3477_n2334), 
        .A2(DP_OP_422J2_124_3477_n2435), .Y(DP_OP_422J2_124_3477_n2410) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1637 ( .A1(DP_OP_423J2_125_3477_n2333), .A2(
        DP_OP_422J2_124_3477_n2435), .Y(DP_OP_422J2_124_3477_n2409) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1630 ( .A1(DP_OP_423J2_125_3477_n2334), 
        .A2(DP_OP_422J2_124_3477_n2434), .Y(DP_OP_422J2_124_3477_n2402) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1629 ( .A1(DP_OP_423J2_125_3477_n2333), .A2(
        DP_OP_422J2_124_3477_n2434), .Y(DP_OP_422J2_124_3477_n2401) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1628 ( .A1(DP_OP_422J2_124_3477_n2432), .A2(
        DP_OP_422J2_124_3477_n2433), .Y(DP_OP_422J2_124_3477_n2400) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1627 ( .A1(DP_OP_423J2_125_3477_n2339), .A2(
        DP_OP_422J2_124_3477_n2433), .Y(DP_OP_422J2_124_3477_n2399) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1626 ( .A1(DP_OP_422J2_124_3477_n2430), .A2(
        DP_OP_422J2_124_3477_n2433), .Y(DP_OP_422J2_124_3477_n2398) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1625 ( .A1(DP_OP_422J2_124_3477_n2429), .A2(
        DP_OP_422J2_124_3477_n2433), .Y(DP_OP_422J2_124_3477_n2397) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1624 ( .A1(DP_OP_422J2_124_3477_n2428), .A2(
        DP_OP_422J2_124_3477_n2433), .Y(DP_OP_422J2_124_3477_n2396) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1623 ( .A1(DP_OP_422J2_124_3477_n2427), .A2(
        DP_OP_422J2_124_3477_n2433), .Y(DP_OP_422J2_124_3477_n2395) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1622 ( .A1(DP_OP_423J2_125_3477_n2334), .A2(
        DP_OP_422J2_124_3477_n2433), .Y(DP_OP_422J2_124_3477_n2394) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1621 ( .A1(DP_OP_423J2_125_3477_n2333), 
        .A2(DP_OP_422J2_124_3477_n2433), .Y(DP_OP_422J2_124_3477_n2393) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1601 ( .A1(DP_OP_422J2_124_3477_n2381), .A2(
        DP_OP_422J2_124_3477_n2392), .Y(DP_OP_422J2_124_3477_n2373) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1594 ( .A1(DP_OP_422J2_124_3477_n2382), 
        .A2(DP_OP_422J2_124_3477_n2391), .Y(DP_OP_422J2_124_3477_n2366) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1593 ( .A1(DP_OP_422J2_124_3477_n2381), .A2(
        DP_OP_422J2_124_3477_n2391), .Y(DP_OP_422J2_124_3477_n2365) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1586 ( .A1(DP_OP_422J2_124_3477_n2382), 
        .A2(DP_OP_422J2_124_3477_n2390), .Y(DP_OP_422J2_124_3477_n2358) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1585 ( .A1(DP_OP_422J2_124_3477_n2381), .A2(
        DP_OP_422J2_124_3477_n2390), .Y(DP_OP_422J2_124_3477_n2357) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1584 ( .A1(DP_OP_422J2_124_3477_n2388), .A2(
        DP_OP_422J2_124_3477_n2389), .Y(DP_OP_422J2_124_3477_n2356) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1583 ( .A1(DP_OP_422J2_124_3477_n2387), .A2(
        DP_OP_422J2_124_3477_n2389), .Y(DP_OP_422J2_124_3477_n2355) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1582 ( .A1(DP_OP_422J2_124_3477_n2386), .A2(
        DP_OP_422J2_124_3477_n2389), .Y(DP_OP_422J2_124_3477_n2354) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1581 ( .A1(DP_OP_422J2_124_3477_n2385), .A2(
        DP_OP_422J2_124_3477_n2389), .Y(DP_OP_422J2_124_3477_n2353) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1580 ( .A1(DP_OP_422J2_124_3477_n2384), .A2(
        DP_OP_422J2_124_3477_n2389), .Y(DP_OP_422J2_124_3477_n2352) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1579 ( .A1(DP_OP_422J2_124_3477_n2383), .A2(
        DP_OP_422J2_124_3477_n2389), .Y(DP_OP_422J2_124_3477_n2351) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1578 ( .A1(DP_OP_422J2_124_3477_n2382), .A2(
        DP_OP_422J2_124_3477_n2389), .Y(DP_OP_422J2_124_3477_n2350) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1577 ( .A1(DP_OP_422J2_124_3477_n2381), 
        .A2(DP_OP_422J2_124_3477_n2389), .Y(DP_OP_422J2_124_3477_n2349) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1559 ( .A1(DP_OP_422J2_124_3477_n2339), 
        .A2(DP_OP_423J2_125_3477_n2344), .Y(DP_OP_422J2_124_3477_n2331) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1558 ( .A1(DP_OP_422J2_124_3477_n2338), 
        .A2(DP_OP_425J2_127_3477_n2349), .Y(DP_OP_422J2_124_3477_n2330) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1557 ( .A1(DP_OP_423J2_125_3477_n2377), .A2(
        DP_OP_423J2_125_3477_n2344), .Y(DP_OP_422J2_124_3477_n2329) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1550 ( .A1(DP_OP_422J2_124_3477_n2338), 
        .A2(DP_OP_422J2_124_3477_n2347), .Y(DP_OP_422J2_124_3477_n2322) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1549 ( .A1(DP_OP_423J2_125_3477_n2377), .A2(
        DP_OP_422J2_124_3477_n2347), .Y(DP_OP_422J2_124_3477_n2321) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1542 ( .A1(DP_OP_422J2_124_3477_n2338), 
        .A2(DP_OP_422J2_124_3477_n2346), .Y(DP_OP_422J2_124_3477_n2314) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1541 ( .A1(DP_OP_423J2_125_3477_n2377), .A2(
        DP_OP_422J2_124_3477_n2346), .Y(DP_OP_422J2_124_3477_n2313) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1540 ( .A1(DP_OP_422J2_124_3477_n2344), .A2(
        DP_OP_422J2_124_3477_n2345), .Y(DP_OP_422J2_124_3477_n2312) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1539 ( .A1(DP_OP_422J2_124_3477_n2343), .A2(
        DP_OP_422J2_124_3477_n2345), .Y(DP_OP_422J2_124_3477_n2311) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1538 ( .A1(DP_OP_422J2_124_3477_n2342), .A2(
        DP_OP_422J2_124_3477_n2345), .Y(DP_OP_422J2_124_3477_n2310) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1537 ( .A1(DP_OP_422J2_124_3477_n2341), .A2(
        DP_OP_422J2_124_3477_n2345), .Y(DP_OP_422J2_124_3477_n2309) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1536 ( .A1(DP_OP_422J2_124_3477_n2340), .A2(
        DP_OP_422J2_124_3477_n2345), .Y(DP_OP_422J2_124_3477_n2308) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1535 ( .A1(DP_OP_422J2_124_3477_n2339), .A2(
        DP_OP_422J2_124_3477_n2345), .Y(DP_OP_422J2_124_3477_n2307) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1534 ( .A1(DP_OP_422J2_124_3477_n2338), .A2(
        DP_OP_422J2_124_3477_n2345), .Y(DP_OP_422J2_124_3477_n2306) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1533 ( .A1(DP_OP_423J2_125_3477_n2377), 
        .A2(DP_OP_422J2_124_3477_n2345), .Y(DP_OP_422J2_124_3477_n2305) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1514 ( .A1(DP_OP_422J2_124_3477_n2294), 
        .A2(DP_OP_422J2_124_3477_n2304), .Y(DP_OP_422J2_124_3477_n2286) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1513 ( .A1(DP_OP_423J2_125_3477_n2421), .A2(
        DP_OP_422J2_124_3477_n2304), .Y(DP_OP_422J2_124_3477_n2285) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1506 ( .A1(DP_OP_422J2_124_3477_n2294), 
        .A2(DP_OP_423J2_125_3477_n2299), .Y(DP_OP_422J2_124_3477_n2278) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1505 ( .A1(DP_OP_423J2_125_3477_n2421), .A2(
        DP_OP_425J2_127_3477_n2304), .Y(DP_OP_422J2_124_3477_n2277) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1498 ( .A1(DP_OP_422J2_124_3477_n2294), 
        .A2(DP_OP_422J2_124_3477_n2302), .Y(DP_OP_422J2_124_3477_n2270) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1497 ( .A1(DP_OP_423J2_125_3477_n2421), .A2(
        DP_OP_422J2_124_3477_n2302), .Y(DP_OP_422J2_124_3477_n2269) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1496 ( .A1(DP_OP_423J2_125_3477_n2428), .A2(
        DP_OP_422J2_124_3477_n2301), .Y(DP_OP_422J2_124_3477_n2268) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1495 ( .A1(DP_OP_422J2_124_3477_n2299), .A2(
        DP_OP_422J2_124_3477_n2301), .Y(DP_OP_422J2_124_3477_n2267) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1494 ( .A1(DP_OP_422J2_124_3477_n2298), .A2(
        DP_OP_422J2_124_3477_n2301), .Y(DP_OP_422J2_124_3477_n2266) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1493 ( .A1(DP_OP_423J2_125_3477_n2425), .A2(
        DP_OP_422J2_124_3477_n2301), .Y(DP_OP_422J2_124_3477_n2265) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1492 ( .A1(DP_OP_423J2_125_3477_n2424), .A2(
        DP_OP_422J2_124_3477_n2301), .Y(DP_OP_422J2_124_3477_n2264) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1491 ( .A1(DP_OP_422J2_124_3477_n2295), .A2(
        DP_OP_422J2_124_3477_n2301), .Y(DP_OP_422J2_124_3477_n2263) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1490 ( .A1(DP_OP_422J2_124_3477_n2294), .A2(
        DP_OP_422J2_124_3477_n2301), .Y(DP_OP_422J2_124_3477_n2262) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1489 ( .A1(DP_OP_423J2_125_3477_n2421), 
        .A2(DP_OP_422J2_124_3477_n2301), .Y(DP_OP_422J2_124_3477_n2261) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1471 ( .A1(DP_OP_424J2_126_3477_n2381), 
        .A2(DP_OP_422J2_124_3477_n2260), .Y(DP_OP_422J2_124_3477_n2243) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1470 ( .A1(DP_OP_422J2_124_3477_n2250), 
        .A2(DP_OP_422J2_124_3477_n2260), .Y(DP_OP_422J2_124_3477_n2242) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1469 ( .A1(DP_OP_422J2_124_3477_n2249), .A2(
        DP_OP_422J2_124_3477_n2260), .Y(DP_OP_422J2_124_3477_n2241) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1462 ( .A1(DP_OP_422J2_124_3477_n2250), 
        .A2(DP_OP_422J2_124_3477_n2259), .Y(DP_OP_422J2_124_3477_n2234) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1461 ( .A1(DP_OP_422J2_124_3477_n2249), .A2(
        DP_OP_422J2_124_3477_n2259), .Y(DP_OP_422J2_124_3477_n2233) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1454 ( .A1(DP_OP_422J2_124_3477_n2250), 
        .A2(DP_OP_422J2_124_3477_n2258), .Y(DP_OP_422J2_124_3477_n2226) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1453 ( .A1(DP_OP_422J2_124_3477_n2249), .A2(
        DP_OP_422J2_124_3477_n2258), .Y(DP_OP_422J2_124_3477_n2225) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1452 ( .A1(DP_OP_424J2_126_3477_n2386), .A2(
        DP_OP_422J2_124_3477_n2257), .Y(DP_OP_422J2_124_3477_n2224) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1451 ( .A1(DP_OP_424J2_126_3477_n2385), .A2(
        DP_OP_422J2_124_3477_n2257), .Y(DP_OP_422J2_124_3477_n2223) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1450 ( .A1(DP_OP_424J2_126_3477_n2384), .A2(
        DP_OP_422J2_124_3477_n2257), .Y(DP_OP_422J2_124_3477_n2222) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1449 ( .A1(DP_OP_424J2_126_3477_n2383), .A2(
        DP_OP_422J2_124_3477_n2257), .Y(DP_OP_422J2_124_3477_n2221) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1448 ( .A1(DP_OP_424J2_126_3477_n2382), .A2(
        DP_OP_422J2_124_3477_n2257), .Y(DP_OP_422J2_124_3477_n2220) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1447 ( .A1(DP_OP_424J2_126_3477_n2381), .A2(
        DP_OP_422J2_124_3477_n2257), .Y(DP_OP_422J2_124_3477_n2219) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1446 ( .A1(DP_OP_422J2_124_3477_n2250), .A2(
        DP_OP_422J2_124_3477_n2257), .Y(DP_OP_422J2_124_3477_n2218) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1445 ( .A1(DP_OP_422J2_124_3477_n2249), 
        .A2(DP_OP_422J2_124_3477_n2257), .Y(DP_OP_422J2_124_3477_n2217) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1426 ( .A1(DP_OP_423J2_125_3477_n2510), 
        .A2(DP_OP_422J2_124_3477_n2216), .Y(DP_OP_422J2_124_3477_n2198) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1425 ( .A1(DP_OP_424J2_126_3477_n2423), .A2(
        DP_OP_422J2_124_3477_n2216), .Y(DP_OP_422J2_124_3477_n2197) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1418 ( .A1(DP_OP_423J2_125_3477_n2510), 
        .A2(DP_OP_422J2_124_3477_n2215), .Y(DP_OP_422J2_124_3477_n2190) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1417 ( .A1(DP_OP_423J2_125_3477_n2509), .A2(
        DP_OP_422J2_124_3477_n2215), .Y(DP_OP_422J2_124_3477_n2189) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1410 ( .A1(DP_OP_425J2_127_3477_n2339), 
        .A2(DP_OP_422J2_124_3477_n2214), .Y(DP_OP_422J2_124_3477_n2182) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1409 ( .A1(DP_OP_424J2_126_3477_n2423), .A2(
        DP_OP_422J2_124_3477_n2214), .Y(DP_OP_422J2_124_3477_n2181) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1408 ( .A1(DP_OP_424J2_126_3477_n2430), .A2(
        DP_OP_422J2_124_3477_n2213), .Y(DP_OP_422J2_124_3477_n2180) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1407 ( .A1(DP_OP_422J2_124_3477_n2211), .A2(
        DP_OP_422J2_124_3477_n2213), .Y(DP_OP_422J2_124_3477_n2179) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1406 ( .A1(DP_OP_422J2_124_3477_n2210), .A2(
        DP_OP_422J2_124_3477_n2213), .Y(DP_OP_422J2_124_3477_n2178) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1405 ( .A1(DP_OP_422J2_124_3477_n2209), .A2(
        DP_OP_422J2_124_3477_n2213), .Y(DP_OP_422J2_124_3477_n2177) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1404 ( .A1(DP_OP_422J2_124_3477_n2208), .A2(
        DP_OP_422J2_124_3477_n2213), .Y(DP_OP_422J2_124_3477_n2176) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1403 ( .A1(DP_OP_422J2_124_3477_n2207), .A2(
        DP_OP_422J2_124_3477_n2213), .Y(DP_OP_422J2_124_3477_n2175) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1402 ( .A1(DP_OP_423J2_125_3477_n2510), .A2(
        DP_OP_422J2_124_3477_n2213), .Y(DP_OP_422J2_124_3477_n2174) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1401 ( .A1(DP_OP_424J2_126_3477_n2423), 
        .A2(DP_OP_422J2_124_3477_n2213), .Y(DP_OP_422J2_124_3477_n2173) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1382 ( .A1(DP_OP_422J2_124_3477_n2162), 
        .A2(DP_OP_424J2_126_3477_n2173), .Y(DP_OP_422J2_124_3477_n2154) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1381 ( .A1(DP_OP_423J2_125_3477_n2553), .A2(
        DP_OP_424J2_126_3477_n2173), .Y(DP_OP_422J2_124_3477_n2153) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1374 ( .A1(DP_OP_422J2_124_3477_n2162), 
        .A2(DP_OP_422J2_124_3477_n2171), .Y(DP_OP_422J2_124_3477_n2146) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1373 ( .A1(DP_OP_423J2_125_3477_n2553), .A2(
        DP_OP_422J2_124_3477_n2171), .Y(DP_OP_422J2_124_3477_n2145) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1366 ( .A1(DP_OP_422J2_124_3477_n2162), 
        .A2(DP_OP_422J2_124_3477_n2170), .Y(DP_OP_422J2_124_3477_n2138) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1365 ( .A1(DP_OP_423J2_125_3477_n2553), .A2(
        DP_OP_422J2_124_3477_n2170), .Y(DP_OP_422J2_124_3477_n2137) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1364 ( .A1(DP_OP_422J2_124_3477_n2168), .A2(
        DP_OP_422J2_124_3477_n2169), .Y(DP_OP_422J2_124_3477_n2136) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1363 ( .A1(DP_OP_425J2_127_3477_n2300), .A2(
        DP_OP_422J2_124_3477_n2169), .Y(DP_OP_422J2_124_3477_n2135) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1362 ( .A1(DP_OP_423J2_125_3477_n2558), .A2(
        DP_OP_422J2_124_3477_n2169), .Y(DP_OP_422J2_124_3477_n2134) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1361 ( .A1(DP_OP_422J2_124_3477_n2165), .A2(
        DP_OP_422J2_124_3477_n2169), .Y(DP_OP_422J2_124_3477_n2133) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1360 ( .A1(DP_OP_422J2_124_3477_n2164), .A2(
        DP_OP_422J2_124_3477_n2169), .Y(DP_OP_422J2_124_3477_n2132) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1359 ( .A1(DP_OP_422J2_124_3477_n2163), .A2(
        DP_OP_422J2_124_3477_n2169), .Y(DP_OP_422J2_124_3477_n2131) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1358 ( .A1(DP_OP_422J2_124_3477_n2162), .A2(
        DP_OP_422J2_124_3477_n2169), .Y(DP_OP_422J2_124_3477_n2130) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1357 ( .A1(DP_OP_425J2_127_3477_n2294), 
        .A2(DP_OP_422J2_124_3477_n2169), .Y(DP_OP_422J2_124_3477_n2129) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1338 ( .A1(DP_OP_422J2_124_3477_n2118), 
        .A2(DP_OP_422J2_124_3477_n2128), .Y(DP_OP_422J2_124_3477_n2110) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1337 ( .A1(DP_OP_422J2_124_3477_n2117), .A2(
        DP_OP_422J2_124_3477_n2128), .Y(DP_OP_422J2_124_3477_n2109) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1330 ( .A1(DP_OP_422J2_124_3477_n2118), 
        .A2(DP_OP_422J2_124_3477_n2127), .Y(DP_OP_422J2_124_3477_n2102) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1329 ( .A1(DP_OP_422J2_124_3477_n2117), .A2(
        DP_OP_422J2_124_3477_n2127), .Y(DP_OP_422J2_124_3477_n2101) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1321 ( .A1(DP_OP_422J2_124_3477_n2117), .A2(
        DP_OP_424J2_126_3477_n2127), .Y(DP_OP_422J2_124_3477_n2093) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1320 ( .A1(DP_OP_422J2_124_3477_n2124), .A2(
        DP_OP_422J2_124_3477_n2125), .Y(DP_OP_422J2_124_3477_n2092) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1319 ( .A1(DP_OP_423J2_125_3477_n2603), .A2(
        DP_OP_422J2_124_3477_n2125), .Y(DP_OP_422J2_124_3477_n2091) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1318 ( .A1(DP_OP_423J2_125_3477_n2602), .A2(
        DP_OP_422J2_124_3477_n2125), .Y(DP_OP_422J2_124_3477_n2090) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1317 ( .A1(DP_OP_422J2_124_3477_n2121), .A2(
        DP_OP_422J2_124_3477_n2125), .Y(DP_OP_422J2_124_3477_n2089) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1316 ( .A1(DP_OP_422J2_124_3477_n2120), .A2(
        DP_OP_422J2_124_3477_n2125), .Y(DP_OP_422J2_124_3477_n2088) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1315 ( .A1(DP_OP_425J2_127_3477_n2252), .A2(
        DP_OP_422J2_124_3477_n2125), .Y(DP_OP_422J2_124_3477_n2087) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1314 ( .A1(DP_OP_422J2_124_3477_n2118), .A2(
        DP_OP_422J2_124_3477_n2125), .Y(DP_OP_422J2_124_3477_n2086) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1313 ( .A1(DP_OP_422J2_124_3477_n2117), 
        .A2(DP_OP_422J2_124_3477_n2125), .Y(DP_OP_422J2_124_3477_n2085) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1294 ( .A1(DP_OP_422J2_124_3477_n2074), 
        .A2(DP_OP_424J2_126_3477_n2085), .Y(DP_OP_422J2_124_3477_n2066) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1293 ( .A1(DP_OP_422J2_124_3477_n2073), .A2(
        n441), .Y(DP_OP_422J2_124_3477_n2065) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1286 ( .A1(DP_OP_422J2_124_3477_n2074), 
        .A2(DP_OP_422J2_124_3477_n2083), .Y(DP_OP_422J2_124_3477_n2058) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1285 ( .A1(DP_OP_422J2_124_3477_n2073), .A2(
        DP_OP_422J2_124_3477_n2083), .Y(DP_OP_422J2_124_3477_n2057) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1278 ( .A1(DP_OP_422J2_124_3477_n2074), 
        .A2(DP_OP_422J2_124_3477_n2082), .Y(DP_OP_422J2_124_3477_n2050) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1277 ( .A1(DP_OP_422J2_124_3477_n2073), .A2(
        DP_OP_422J2_124_3477_n2082), .Y(DP_OP_422J2_124_3477_n2049) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1276 ( .A1(DP_OP_425J2_127_3477_n2213), .A2(
        DP_OP_422J2_124_3477_n2081), .Y(DP_OP_422J2_124_3477_n2048) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1275 ( .A1(DP_OP_423J2_125_3477_n2647), .A2(
        DP_OP_422J2_124_3477_n2081), .Y(DP_OP_422J2_124_3477_n2047) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1274 ( .A1(DP_OP_422J2_124_3477_n2078), .A2(
        DP_OP_422J2_124_3477_n2081), .Y(DP_OP_422J2_124_3477_n2046) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1273 ( .A1(DP_OP_423J2_125_3477_n2645), .A2(
        DP_OP_422J2_124_3477_n2081), .Y(DP_OP_422J2_124_3477_n2045) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1272 ( .A1(DP_OP_422J2_124_3477_n2076), .A2(
        DP_OP_422J2_124_3477_n2081), .Y(DP_OP_422J2_124_3477_n2044) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1271 ( .A1(DP_OP_423J2_125_3477_n2643), .A2(
        DP_OP_422J2_124_3477_n2081), .Y(DP_OP_422J2_124_3477_n2043) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1270 ( .A1(DP_OP_422J2_124_3477_n2074), .A2(
        DP_OP_422J2_124_3477_n2081), .Y(DP_OP_422J2_124_3477_n2042) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1269 ( .A1(DP_OP_422J2_124_3477_n2073), 
        .A2(DP_OP_422J2_124_3477_n2081), .Y(DP_OP_422J2_124_3477_n2041) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1250 ( .A1(DP_OP_424J2_126_3477_n2600), 
        .A2(DP_OP_422J2_124_3477_n2040), .Y(DP_OP_422J2_124_3477_n2022) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1249 ( .A1(DP_OP_422J2_124_3477_n2029), .A2(
        DP_OP_422J2_124_3477_n2040), .Y(DP_OP_422J2_124_3477_n2021) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1242 ( .A1(DP_OP_424J2_126_3477_n2600), 
        .A2(DP_OP_422J2_124_3477_n2039), .Y(DP_OP_422J2_124_3477_n2014) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1241 ( .A1(DP_OP_422J2_124_3477_n2029), .A2(
        DP_OP_422J2_124_3477_n2039), .Y(DP_OP_422J2_124_3477_n2013) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1234 ( .A1(DP_OP_424J2_126_3477_n2600), 
        .A2(DP_OP_423J2_125_3477_n2034), .Y(DP_OP_422J2_124_3477_n2006) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1233 ( .A1(DP_OP_422J2_124_3477_n2029), .A2(
        DP_OP_425J2_127_3477_n2039), .Y(DP_OP_422J2_124_3477_n2005) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1232 ( .A1(DP_OP_422J2_124_3477_n2036), .A2(
        DP_OP_422J2_124_3477_n2037), .Y(DP_OP_422J2_124_3477_n1579) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1231 ( .A1(DP_OP_422J2_124_3477_n2035), .A2(
        DP_OP_422J2_124_3477_n2037), .Y(DP_OP_422J2_124_3477_n2004) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1230 ( .A1(DP_OP_424J2_126_3477_n2604), .A2(
        DP_OP_422J2_124_3477_n2037), .Y(DP_OP_422J2_124_3477_n2003) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1229 ( .A1(DP_OP_422J2_124_3477_n2033), .A2(
        DP_OP_422J2_124_3477_n2037), .Y(DP_OP_422J2_124_3477_n2002) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1228 ( .A1(DP_OP_422J2_124_3477_n2032), .A2(
        DP_OP_422J2_124_3477_n2037), .Y(DP_OP_422J2_124_3477_n2001) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1227 ( .A1(DP_OP_422J2_124_3477_n2031), .A2(
        DP_OP_422J2_124_3477_n2037), .Y(DP_OP_422J2_124_3477_n2000) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1226 ( .A1(DP_OP_424J2_126_3477_n2600), .A2(
        DP_OP_422J2_124_3477_n2037), .Y(DP_OP_422J2_124_3477_n1999) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1225 ( .A1(DP_OP_422J2_124_3477_n2029), 
        .A2(DP_OP_422J2_124_3477_n2037), .Y(DP_OP_422J2_124_3477_n1998) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1207 ( .A1(DP_OP_422J2_124_3477_n1988), 
        .A2(DP_OP_422J2_124_3477_n1997), .Y(DP_OP_422J2_124_3477_n1980) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1206 ( .A1(DP_OP_425J2_127_3477_n2119), 
        .A2(DP_OP_422J2_124_3477_n1997), .Y(DP_OP_422J2_124_3477_n1979) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1205 ( .A1(DP_OP_425J2_127_3477_n2118), .A2(
        DP_OP_422J2_124_3477_n1997), .Y(DP_OP_422J2_124_3477_n1978) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1197 ( .A1(DP_OP_423J2_125_3477_n2726), .A2(
        DP_OP_422J2_124_3477_n1996), .Y(DP_OP_422J2_124_3477_n1970) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1190 ( .A1(DP_OP_425J2_127_3477_n2119), 
        .A2(DP_OP_422J2_124_3477_n1995), .Y(DP_OP_422J2_124_3477_n1963) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1189 ( .A1(DP_OP_423J2_125_3477_n2726), .A2(
        DP_OP_422J2_124_3477_n1995), .Y(DP_OP_422J2_124_3477_n1962) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1188 ( .A1(DP_OP_423J2_125_3477_n2733), .A2(
        DP_OP_422J2_124_3477_n1994), .Y(DP_OP_422J2_124_3477_n1961) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1187 ( .A1(DP_OP_424J2_126_3477_n2649), .A2(
        DP_OP_422J2_124_3477_n1994), .Y(DP_OP_422J2_124_3477_n1960) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1186 ( .A1(DP_OP_422J2_124_3477_n1991), .A2(
        DP_OP_422J2_124_3477_n1994), .Y(DP_OP_422J2_124_3477_n1959) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1185 ( .A1(DP_OP_423J2_125_3477_n2730), .A2(
        DP_OP_422J2_124_3477_n1994), .Y(DP_OP_422J2_124_3477_n1958) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1184 ( .A1(DP_OP_422J2_124_3477_n1989), .A2(
        DP_OP_422J2_124_3477_n1994), .Y(DP_OP_422J2_124_3477_n1957) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1183 ( .A1(DP_OP_422J2_124_3477_n1988), .A2(
        DP_OP_422J2_124_3477_n1994), .Y(DP_OP_422J2_124_3477_n1956) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1182 ( .A1(DP_OP_425J2_127_3477_n2119), .A2(
        DP_OP_422J2_124_3477_n1994), .Y(DP_OP_422J2_124_3477_n1955) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1181 ( .A1(DP_OP_425J2_127_3477_n2118), 
        .A2(DP_OP_422J2_124_3477_n1994), .Y(DP_OP_422J2_124_3477_n1954) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1162 ( .A1(DP_OP_422J2_124_3477_n1943), 
        .A2(DP_OP_425J2_127_3477_n1953), .Y(DP_OP_422J2_124_3477_n1935) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1161 ( .A1(DP_OP_423J2_125_3477_n2770), .A2(
        DP_OP_423J2_125_3477_n1948), .Y(DP_OP_422J2_124_3477_n1934) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1153 ( .A1(DP_OP_423J2_125_3477_n2770), .A2(
        DP_OP_422J2_124_3477_n1952), .Y(DP_OP_422J2_124_3477_n1926) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1146 ( .A1(DP_OP_422J2_124_3477_n1943), 
        .A2(DP_OP_422J2_124_3477_n1951), .Y(DP_OP_422J2_124_3477_n1919) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1145 ( .A1(DP_OP_423J2_125_3477_n2770), .A2(
        DP_OP_422J2_124_3477_n1951), .Y(DP_OP_422J2_124_3477_n1918) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1144 ( .A1(DP_OP_422J2_124_3477_n1949), .A2(
        DP_OP_422J2_124_3477_n1950), .Y(DP_OP_422J2_124_3477_n1917) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1143 ( .A1(DP_OP_424J2_126_3477_n2693), .A2(
        DP_OP_422J2_124_3477_n1950), .Y(DP_OP_422J2_124_3477_n1916) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1142 ( .A1(DP_OP_423J2_125_3477_n2775), .A2(
        DP_OP_422J2_124_3477_n1950), .Y(DP_OP_422J2_124_3477_n1915) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1141 ( .A1(DP_OP_424J2_126_3477_n2691), .A2(
        DP_OP_422J2_124_3477_n1950), .Y(DP_OP_422J2_124_3477_n1914) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1140 ( .A1(DP_OP_422J2_124_3477_n1945), .A2(
        DP_OP_422J2_124_3477_n1950), .Y(DP_OP_422J2_124_3477_n1913) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1139 ( .A1(DP_OP_424J2_126_3477_n2689), .A2(
        DP_OP_422J2_124_3477_n1950), .Y(DP_OP_422J2_124_3477_n1912) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1138 ( .A1(DP_OP_422J2_124_3477_n1943), .A2(
        DP_OP_422J2_124_3477_n1950), .Y(DP_OP_422J2_124_3477_n1911) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1137 ( .A1(DP_OP_423J2_125_3477_n2770), 
        .A2(DP_OP_422J2_124_3477_n1950), .Y(DP_OP_422J2_124_3477_n1910) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1118 ( .A1(DP_OP_422J2_124_3477_n1899), 
        .A2(DP_OP_422J2_124_3477_n1909), .Y(DP_OP_422J2_124_3477_n1891) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1117 ( .A1(DP_OP_422J2_124_3477_n1898), .A2(
        DP_OP_422J2_124_3477_n1909), .Y(DP_OP_422J2_124_3477_n1890) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1110 ( .A1(DP_OP_422J2_124_3477_n1899), 
        .A2(DP_OP_422J2_124_3477_n1908), .Y(DP_OP_422J2_124_3477_n1883) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1109 ( .A1(DP_OP_422J2_124_3477_n1898), .A2(
        DP_OP_422J2_124_3477_n1908), .Y(DP_OP_422J2_124_3477_n1882) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1102 ( .A1(DP_OP_422J2_124_3477_n1899), 
        .A2(DP_OP_422J2_124_3477_n1907), .Y(DP_OP_422J2_124_3477_n1875) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1101 ( .A1(DP_OP_422J2_124_3477_n1898), .A2(
        DP_OP_422J2_124_3477_n1907), .Y(DP_OP_422J2_124_3477_n1874) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1100 ( .A1(DP_OP_422J2_124_3477_n1905), .A2(
        DP_OP_422J2_124_3477_n1906), .Y(DP_OP_422J2_124_3477_n1873) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1099 ( .A1(DP_OP_422J2_124_3477_n1904), .A2(
        DP_OP_422J2_124_3477_n1906), .Y(DP_OP_422J2_124_3477_n1872) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1098 ( .A1(DP_OP_422J2_124_3477_n1903), .A2(
        DP_OP_422J2_124_3477_n1906), .Y(DP_OP_422J2_124_3477_n1871) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1097 ( .A1(DP_OP_422J2_124_3477_n1902), .A2(
        DP_OP_422J2_124_3477_n1906), .Y(DP_OP_422J2_124_3477_n1870) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1096 ( .A1(DP_OP_424J2_126_3477_n2734), .A2(
        DP_OP_422J2_124_3477_n1906), .Y(DP_OP_422J2_124_3477_n1869) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1095 ( .A1(DP_OP_422J2_124_3477_n1900), .A2(
        DP_OP_422J2_124_3477_n1906), .Y(DP_OP_422J2_124_3477_n1868) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1094 ( .A1(DP_OP_422J2_124_3477_n1899), .A2(
        DP_OP_422J2_124_3477_n1906), .Y(DP_OP_422J2_124_3477_n1867) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1093 ( .A1(DP_OP_422J2_124_3477_n1898), 
        .A2(DP_OP_422J2_124_3477_n1906), .Y(DP_OP_422J2_124_3477_n1866) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1074 ( .A1(DP_OP_422J2_124_3477_n1855), 
        .A2(DP_OP_422J2_124_3477_n1865), .Y(DP_OP_422J2_124_3477_n1847) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1073 ( .A1(DP_OP_422J2_124_3477_n1854), .A2(
        DP_OP_422J2_124_3477_n1865), .Y(DP_OP_422J2_124_3477_n1846) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1066 ( .A1(DP_OP_422J2_124_3477_n1855), 
        .A2(DP_OP_422J2_124_3477_n1864), .Y(DP_OP_422J2_124_3477_n1839) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1065 ( .A1(DP_OP_422J2_124_3477_n1854), .A2(
        DP_OP_422J2_124_3477_n1864), .Y(DP_OP_422J2_124_3477_n1838) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1058 ( .A1(DP_OP_422J2_124_3477_n1855), 
        .A2(DP_OP_422J2_124_3477_n1863), .Y(DP_OP_422J2_124_3477_n1831) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1057 ( .A1(DP_OP_422J2_124_3477_n1854), .A2(
        DP_OP_422J2_124_3477_n1863), .Y(DP_OP_422J2_124_3477_n1830) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1056 ( .A1(DP_OP_422J2_124_3477_n1861), .A2(
        DP_OP_422J2_124_3477_n1862), .Y(DP_OP_422J2_124_3477_n1829) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1055 ( .A1(DP_OP_423J2_125_3477_n2864), .A2(
        DP_OP_422J2_124_3477_n1862), .Y(DP_OP_422J2_124_3477_n1828) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1054 ( .A1(DP_OP_422J2_124_3477_n1859), .A2(
        DP_OP_422J2_124_3477_n1862), .Y(DP_OP_422J2_124_3477_n1827) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1053 ( .A1(DP_OP_422J2_124_3477_n1858), .A2(
        DP_OP_422J2_124_3477_n1862), .Y(DP_OP_422J2_124_3477_n1826) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1052 ( .A1(DP_OP_423J2_125_3477_n2861), .A2(
        DP_OP_422J2_124_3477_n1862), .Y(DP_OP_422J2_124_3477_n1825) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1051 ( .A1(DP_OP_424J2_126_3477_n2777), .A2(
        DP_OP_422J2_124_3477_n1862), .Y(DP_OP_422J2_124_3477_n1824) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1050 ( .A1(DP_OP_422J2_124_3477_n1855), .A2(
        DP_OP_422J2_124_3477_n1862), .Y(DP_OP_422J2_124_3477_n1823) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1049 ( .A1(DP_OP_422J2_124_3477_n1854), 
        .A2(DP_OP_422J2_124_3477_n1862), .Y(DP_OP_422J2_124_3477_n1822) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1000 ( .A1(n372), .A2(
        DP_OP_424J2_126_3477_n2), .Y(DP_OP_422J2_124_3477_n1774) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U999 ( .A1(n298), .A2(n337), .Y(
        DP_OP_422J2_124_3477_n181) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U998 ( .A1(n423), .A2(
        DP_OP_425J2_127_3477_n2), .Y(DP_OP_422J2_124_3477_n179) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U997 ( .A1(n412), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_422J2_124_3477_n177) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U996 ( .A1(n377), .A2(n337), .Y(
        DP_OP_422J2_124_3477_n175) );
  HADDX1_HVT DP_OP_422J2_124_3477_U983 ( .A0(DP_OP_422J2_124_3477_n2644), .B0(
        DP_OP_422J2_124_3477_n2730), .C1(DP_OP_422J2_124_3477_n1771), .SO(
        DP_OP_422J2_124_3477_n1772) );
  FADDX1_HVT DP_OP_422J2_124_3477_U982 ( .A(DP_OP_422J2_124_3477_n2600), .B(
        DP_OP_422J2_124_3477_n1788), .CI(DP_OP_422J2_124_3477_n2292), .CO(
        DP_OP_422J2_124_3477_n1769), .S(DP_OP_422J2_124_3477_n1770) );
  FADDX1_HVT DP_OP_422J2_124_3477_U981 ( .A(DP_OP_422J2_124_3477_n1853), .B(
        DP_OP_422J2_124_3477_n2028), .CI(DP_OP_422J2_124_3477_n2072), .CO(
        DP_OP_422J2_124_3477_n1767), .S(DP_OP_422J2_124_3477_n1768) );
  FADDX1_HVT DP_OP_422J2_124_3477_U980 ( .A(DP_OP_422J2_124_3477_n2204), .B(
        DP_OP_422J2_124_3477_n1985), .CI(DP_OP_422J2_124_3477_n2512), .CO(
        DP_OP_422J2_124_3477_n1765), .S(DP_OP_422J2_124_3477_n1766) );
  FADDX1_HVT DP_OP_422J2_124_3477_U979 ( .A(DP_OP_422J2_124_3477_n2556), .B(
        DP_OP_422J2_124_3477_n2688), .CI(DP_OP_422J2_124_3477_n2774), .CO(
        DP_OP_422J2_124_3477_n1763), .S(DP_OP_422J2_124_3477_n1764) );
  FADDX1_HVT DP_OP_422J2_124_3477_U978 ( .A(DP_OP_422J2_124_3477_n2424), .B(
        DP_OP_422J2_124_3477_n2336), .CI(DP_OP_422J2_124_3477_n2862), .CO(
        DP_OP_422J2_124_3477_n1761), .S(DP_OP_422J2_124_3477_n1762) );
  FADDX1_HVT DP_OP_422J2_124_3477_U977 ( .A(DP_OP_422J2_124_3477_n2468), .B(
        DP_OP_422J2_124_3477_n2116), .CI(DP_OP_422J2_124_3477_n1897), .CO(
        DP_OP_422J2_124_3477_n1759), .S(DP_OP_422J2_124_3477_n1760) );
  FADDX1_HVT DP_OP_422J2_124_3477_U976 ( .A(DP_OP_422J2_124_3477_n2248), .B(
        DP_OP_422J2_124_3477_n1941), .CI(DP_OP_422J2_124_3477_n2906), .CO(
        DP_OP_422J2_124_3477_n1757), .S(DP_OP_422J2_124_3477_n1758) );
  FADDX1_HVT DP_OP_422J2_124_3477_U975 ( .A(DP_OP_422J2_124_3477_n2160), .B(
        DP_OP_422J2_124_3477_n2380), .CI(DP_OP_422J2_124_3477_n2818), .CO(
        DP_OP_422J2_124_3477_n1755), .S(DP_OP_422J2_124_3477_n1756) );
  FADDX1_HVT DP_OP_422J2_124_3477_U974 ( .A(DP_OP_422J2_124_3477_n1772), .B(
        DP_OP_422J2_124_3477_n1762), .CI(DP_OP_422J2_124_3477_n1764), .CO(
        DP_OP_422J2_124_3477_n1753), .S(DP_OP_422J2_124_3477_n1754) );
  FADDX1_HVT DP_OP_422J2_124_3477_U973 ( .A(DP_OP_422J2_124_3477_n1766), .B(
        DP_OP_422J2_124_3477_n1760), .CI(DP_OP_422J2_124_3477_n1768), .CO(
        DP_OP_422J2_124_3477_n1751), .S(DP_OP_422J2_124_3477_n1752) );
  FADDX1_HVT DP_OP_422J2_124_3477_U972 ( .A(DP_OP_422J2_124_3477_n1770), .B(
        DP_OP_422J2_124_3477_n1758), .CI(DP_OP_422J2_124_3477_n1756), .CO(
        DP_OP_422J2_124_3477_n1749), .S(DP_OP_422J2_124_3477_n1750) );
  HADDX1_HVT DP_OP_422J2_124_3477_U971 ( .A0(DP_OP_422J2_124_3477_n2555), .B0(
        DP_OP_422J2_124_3477_n2416), .C1(DP_OP_422J2_124_3477_n1747), .SO(
        DP_OP_422J2_124_3477_n1748) );
  FADDX1_HVT DP_OP_422J2_124_3477_U970 ( .A(DP_OP_422J2_124_3477_n1852), .B(
        DP_OP_422J2_124_3477_n2729), .CI(DP_OP_422J2_124_3477_n2071), .CO(
        DP_OP_422J2_124_3477_n1745), .S(DP_OP_422J2_124_3477_n1746) );
  FADDX1_HVT DP_OP_422J2_124_3477_U969 ( .A(DP_OP_422J2_124_3477_n2115), .B(
        DP_OP_422J2_124_3477_n2152), .CI(DP_OP_422J2_124_3477_n2291), .CO(
        DP_OP_422J2_124_3477_n1743), .S(DP_OP_422J2_124_3477_n1744) );
  FADDX1_HVT DP_OP_422J2_124_3477_U968 ( .A(DP_OP_422J2_124_3477_n2203), .B(
        DP_OP_422J2_124_3477_n1787), .CI(DP_OP_422J2_124_3477_n2511), .CO(
        DP_OP_422J2_124_3477_n1741), .S(DP_OP_422J2_124_3477_n1742) );
  FADDX1_HVT DP_OP_422J2_124_3477_U967 ( .A(DP_OP_422J2_124_3477_n2599), .B(
        DP_OP_422J2_124_3477_n2328), .CI(DP_OP_422J2_124_3477_n2773), .CO(
        DP_OP_422J2_124_3477_n1739), .S(DP_OP_422J2_124_3477_n1740) );
  FADDX1_HVT DP_OP_422J2_124_3477_U966 ( .A(DP_OP_422J2_124_3477_n2643), .B(
        DP_OP_422J2_124_3477_n2027), .CI(DP_OP_422J2_124_3477_n2861), .CO(
        DP_OP_422J2_124_3477_n1737), .S(DP_OP_422J2_124_3477_n1738) );
  FADDX1_HVT DP_OP_422J2_124_3477_U965 ( .A(DP_OP_422J2_124_3477_n2467), .B(
        DP_OP_422J2_124_3477_n1984), .CI(DP_OP_422J2_124_3477_n1896), .CO(
        DP_OP_422J2_124_3477_n1735), .S(DP_OP_422J2_124_3477_n1736) );
  FADDX1_HVT DP_OP_422J2_124_3477_U964 ( .A(DP_OP_422J2_124_3477_n2423), .B(
        DP_OP_422J2_124_3477_n2592), .CI(DP_OP_422J2_124_3477_n2636), .CO(
        DP_OP_422J2_124_3477_n1733), .S(DP_OP_422J2_124_3477_n1734) );
  FADDX1_HVT DP_OP_422J2_124_3477_U963 ( .A(DP_OP_422J2_124_3477_n2335), .B(
        DP_OP_422J2_124_3477_n2064), .CI(DP_OP_422J2_124_3477_n2504), .CO(
        DP_OP_422J2_124_3477_n1731), .S(DP_OP_422J2_124_3477_n1732) );
  FADDX1_HVT DP_OP_422J2_124_3477_U962 ( .A(DP_OP_422J2_124_3477_n1845), .B(
        DP_OP_422J2_124_3477_n2687), .CI(DP_OP_422J2_124_3477_n1889), .CO(
        DP_OP_422J2_124_3477_n1729), .S(DP_OP_422J2_124_3477_n1730) );
  FADDX1_HVT DP_OP_422J2_124_3477_U961 ( .A(DP_OP_422J2_124_3477_n2108), .B(
        DP_OP_422J2_124_3477_n2854), .CI(DP_OP_422J2_124_3477_n2240), .CO(
        DP_OP_422J2_124_3477_n1727), .S(DP_OP_422J2_124_3477_n1728) );
  FADDX1_HVT DP_OP_422J2_124_3477_U960 ( .A(DP_OP_422J2_124_3477_n2680), .B(
        DP_OP_422J2_124_3477_n1940), .CI(DP_OP_422J2_124_3477_n2196), .CO(
        DP_OP_422J2_124_3477_n1725), .S(DP_OP_422J2_124_3477_n1726) );
  FADDX1_HVT DP_OP_422J2_124_3477_U959 ( .A(DP_OP_422J2_124_3477_n2247), .B(
        DP_OP_422J2_124_3477_n2898), .CI(DP_OP_422J2_124_3477_n2372), .CO(
        DP_OP_422J2_124_3477_n1723), .S(DP_OP_422J2_124_3477_n1724) );
  FADDX1_HVT DP_OP_422J2_124_3477_U958 ( .A(DP_OP_422J2_124_3477_n2460), .B(
        DP_OP_422J2_124_3477_n2810), .CI(DP_OP_422J2_124_3477_n1977), .CO(
        DP_OP_422J2_124_3477_n1721), .S(DP_OP_422J2_124_3477_n1722) );
  FADDX1_HVT DP_OP_422J2_124_3477_U957 ( .A(DP_OP_422J2_124_3477_n2548), .B(
        DP_OP_422J2_124_3477_n2766), .CI(DP_OP_422J2_124_3477_n2379), .CO(
        DP_OP_422J2_124_3477_n1719), .S(DP_OP_422J2_124_3477_n1720) );
  FADDX1_HVT DP_OP_422J2_124_3477_U956 ( .A(DP_OP_422J2_124_3477_n2284), .B(
        DP_OP_422J2_124_3477_n1933), .CI(DP_OP_422J2_124_3477_n2817), .CO(
        DP_OP_422J2_124_3477_n1717), .S(DP_OP_422J2_124_3477_n1718) );
  FADDX1_HVT DP_OP_422J2_124_3477_U955 ( .A(DP_OP_422J2_124_3477_n2159), .B(
        DP_OP_422J2_124_3477_n2722), .CI(DP_OP_422J2_124_3477_n2905), .CO(
        DP_OP_422J2_124_3477_n1715), .S(DP_OP_422J2_124_3477_n1716) );
  FADDX1_HVT DP_OP_422J2_124_3477_U954 ( .A(DP_OP_422J2_124_3477_n2020), .B(
        DP_OP_422J2_124_3477_n1771), .CI(DP_OP_422J2_124_3477_n1748), .CO(
        DP_OP_422J2_124_3477_n1713), .S(DP_OP_422J2_124_3477_n1714) );
  FADDX1_HVT DP_OP_422J2_124_3477_U953 ( .A(DP_OP_422J2_124_3477_n1759), .B(
        DP_OP_422J2_124_3477_n1769), .CI(DP_OP_422J2_124_3477_n1767), .CO(
        DP_OP_422J2_124_3477_n1711), .S(DP_OP_422J2_124_3477_n1712) );
  FADDX1_HVT DP_OP_422J2_124_3477_U952 ( .A(DP_OP_422J2_124_3477_n1763), .B(
        DP_OP_422J2_124_3477_n1765), .CI(DP_OP_422J2_124_3477_n1761), .CO(
        DP_OP_422J2_124_3477_n1709), .S(DP_OP_422J2_124_3477_n1710) );
  FADDX1_HVT DP_OP_422J2_124_3477_U951 ( .A(DP_OP_422J2_124_3477_n1757), .B(
        DP_OP_422J2_124_3477_n1755), .CI(DP_OP_422J2_124_3477_n1738), .CO(
        DP_OP_422J2_124_3477_n1707), .S(DP_OP_422J2_124_3477_n1708) );
  FADDX1_HVT DP_OP_422J2_124_3477_U950 ( .A(DP_OP_422J2_124_3477_n1736), .B(
        DP_OP_422J2_124_3477_n1742), .CI(DP_OP_422J2_124_3477_n1730), .CO(
        DP_OP_422J2_124_3477_n1705), .S(DP_OP_422J2_124_3477_n1706) );
  FADDX1_HVT DP_OP_422J2_124_3477_U949 ( .A(DP_OP_422J2_124_3477_n1740), .B(
        DP_OP_422J2_124_3477_n1746), .CI(DP_OP_422J2_124_3477_n1734), .CO(
        DP_OP_422J2_124_3477_n1703), .S(DP_OP_422J2_124_3477_n1704) );
  FADDX1_HVT DP_OP_422J2_124_3477_U948 ( .A(DP_OP_422J2_124_3477_n1732), .B(
        DP_OP_422J2_124_3477_n1744), .CI(DP_OP_422J2_124_3477_n1728), .CO(
        DP_OP_422J2_124_3477_n1701), .S(DP_OP_422J2_124_3477_n1702) );
  FADDX1_HVT DP_OP_422J2_124_3477_U947 ( .A(DP_OP_422J2_124_3477_n1726), .B(
        DP_OP_422J2_124_3477_n1720), .CI(DP_OP_422J2_124_3477_n1716), .CO(
        DP_OP_422J2_124_3477_n1699), .S(DP_OP_422J2_124_3477_n1700) );
  FADDX1_HVT DP_OP_422J2_124_3477_U946 ( .A(DP_OP_422J2_124_3477_n1724), .B(
        DP_OP_422J2_124_3477_n1722), .CI(DP_OP_422J2_124_3477_n1718), .CO(
        DP_OP_422J2_124_3477_n1697), .S(DP_OP_422J2_124_3477_n1698) );
  FADDX1_HVT DP_OP_422J2_124_3477_U945 ( .A(DP_OP_422J2_124_3477_n1714), .B(
        DP_OP_422J2_124_3477_n1753), .CI(DP_OP_422J2_124_3477_n1751), .CO(
        DP_OP_422J2_124_3477_n1695), .S(DP_OP_422J2_124_3477_n1696) );
  FADDX1_HVT DP_OP_422J2_124_3477_U944 ( .A(DP_OP_422J2_124_3477_n1712), .B(
        DP_OP_422J2_124_3477_n1710), .CI(DP_OP_422J2_124_3477_n1749), .CO(
        DP_OP_422J2_124_3477_n1693), .S(DP_OP_422J2_124_3477_n1694) );
  FADDX1_HVT DP_OP_422J2_124_3477_U943 ( .A(DP_OP_422J2_124_3477_n1708), .B(
        DP_OP_422J2_124_3477_n1706), .CI(DP_OP_422J2_124_3477_n1704), .CO(
        DP_OP_422J2_124_3477_n1691), .S(DP_OP_422J2_124_3477_n1692) );
  FADDX1_HVT DP_OP_422J2_124_3477_U942 ( .A(DP_OP_422J2_124_3477_n1702), .B(
        DP_OP_422J2_124_3477_n1700), .CI(DP_OP_422J2_124_3477_n1698), .CO(
        DP_OP_422J2_124_3477_n1689), .S(DP_OP_422J2_124_3477_n1690) );
  FADDX1_HVT DP_OP_422J2_124_3477_U941 ( .A(DP_OP_422J2_124_3477_n1696), .B(
        DP_OP_422J2_124_3477_n1694), .CI(DP_OP_422J2_124_3477_n1692), .CO(
        DP_OP_422J2_124_3477_n1687), .S(DP_OP_422J2_124_3477_n1688) );
  HADDX1_HVT DP_OP_422J2_124_3477_U940 ( .A0(DP_OP_422J2_124_3477_n2554), .B0(
        DP_OP_422J2_124_3477_n2540), .C1(DP_OP_422J2_124_3477_n1685), .SO(
        DP_OP_422J2_124_3477_n1686) );
  FADDX1_HVT DP_OP_422J2_124_3477_U939 ( .A(DP_OP_422J2_124_3477_n2846), .B(
        DP_OP_422J2_124_3477_n2415), .CI(DP_OP_422J2_124_3477_n2290), .CO(
        DP_OP_422J2_124_3477_n1683), .S(DP_OP_422J2_124_3477_n1684) );
  FADDX1_HVT DP_OP_422J2_124_3477_U938 ( .A(DP_OP_422J2_124_3477_n2334), .B(
        DP_OP_422J2_124_3477_n2151), .CI(DP_OP_422J2_124_3477_n2070), .CO(
        DP_OP_422J2_124_3477_n1681), .S(DP_OP_422J2_124_3477_n1682) );
  FADDX1_HVT DP_OP_422J2_124_3477_U937 ( .A(DP_OP_422J2_124_3477_n2598), .B(
        DP_OP_422J2_124_3477_n1969), .CI(DP_OP_422J2_124_3477_n2276), .CO(
        DP_OP_422J2_124_3477_n1679), .S(DP_OP_422J2_124_3477_n1680) );
  FADDX1_HVT DP_OP_422J2_124_3477_U936 ( .A(DP_OP_422J2_124_3477_n2202), .B(
        DP_OP_422J2_124_3477_n2728), .CI(DP_OP_422J2_124_3477_n2144), .CO(
        DP_OP_422J2_124_3477_n1677), .S(DP_OP_422J2_124_3477_n1678) );
  FADDX1_HVT DP_OP_422J2_124_3477_U935 ( .A(DP_OP_422J2_124_3477_n2422), .B(
        DP_OP_422J2_124_3477_n1786), .CI(DP_OP_422J2_124_3477_n2584), .CO(
        DP_OP_422J2_124_3477_n1675), .S(DP_OP_422J2_124_3477_n1676) );
  FADDX1_HVT DP_OP_422J2_124_3477_U934 ( .A(DP_OP_422J2_124_3477_n2114), .B(
        DP_OP_422J2_124_3477_n2503), .CI(DP_OP_422J2_124_3477_n2510), .CO(
        DP_OP_422J2_124_3477_n1673), .S(DP_OP_422J2_124_3477_n1674) );
  FADDX1_HVT DP_OP_422J2_124_3477_U933 ( .A(DP_OP_422J2_124_3477_n2466), .B(
        DP_OP_422J2_124_3477_n2063), .CI(DP_OP_422J2_124_3477_n2452), .CO(
        DP_OP_422J2_124_3477_n1671), .S(DP_OP_422J2_124_3477_n1672) );
  FADDX1_HVT DP_OP_422J2_124_3477_U932 ( .A(DP_OP_422J2_124_3477_n1851), .B(
        DP_OP_422J2_124_3477_n2026), .CI(DP_OP_422J2_124_3477_n2100), .CO(
        DP_OP_422J2_124_3477_n1669), .S(DP_OP_422J2_124_3477_n1670) );
  FADDX1_HVT DP_OP_422J2_124_3477_U931 ( .A(DP_OP_422J2_124_3477_n2890), .B(
        DP_OP_422J2_124_3477_n2327), .CI(DP_OP_422J2_124_3477_n2232), .CO(
        DP_OP_422J2_124_3477_n1667), .S(DP_OP_422J2_124_3477_n1668) );
  FADDX1_HVT DP_OP_422J2_124_3477_U930 ( .A(DP_OP_422J2_124_3477_n2642), .B(
        DP_OP_422J2_124_3477_n2758), .CI(DP_OP_422J2_124_3477_n2860), .CO(
        DP_OP_422J2_124_3477_n1665), .S(DP_OP_422J2_124_3477_n1666) );
  FADDX1_HVT DP_OP_422J2_124_3477_U929 ( .A(DP_OP_422J2_124_3477_n1983), .B(
        DP_OP_422J2_124_3477_n2686), .CI(DP_OP_422J2_124_3477_n2772), .CO(
        DP_OP_422J2_124_3477_n1663), .S(DP_OP_422J2_124_3477_n1664) );
  FADDX1_HVT DP_OP_422J2_124_3477_U928 ( .A(DP_OP_422J2_124_3477_n2591), .B(
        DP_OP_422J2_124_3477_n2635), .CI(DP_OP_422J2_124_3477_n1895), .CO(
        DP_OP_422J2_124_3477_n1661), .S(DP_OP_422J2_124_3477_n1662) );
  FADDX1_HVT DP_OP_422J2_124_3477_U927 ( .A(DP_OP_422J2_124_3477_n1844), .B(
        DP_OP_422J2_124_3477_n1888), .CI(DP_OP_422J2_124_3477_n2107), .CO(
        DP_OP_422J2_124_3477_n1659), .S(DP_OP_422J2_124_3477_n1660) );
  FADDX1_HVT DP_OP_422J2_124_3477_U926 ( .A(DP_OP_422J2_124_3477_n2496), .B(
        DP_OP_422J2_124_3477_n2320), .CI(DP_OP_422J2_124_3477_n2188), .CO(
        DP_OP_422J2_124_3477_n1657), .S(DP_OP_422J2_124_3477_n1658) );
  FADDX1_HVT DP_OP_422J2_124_3477_U925 ( .A(DP_OP_422J2_124_3477_n2364), .B(
        DP_OP_422J2_124_3477_n2056), .CI(DP_OP_422J2_124_3477_n1925), .CO(
        DP_OP_422J2_124_3477_n1655), .S(DP_OP_422J2_124_3477_n1656) );
  FADDX1_HVT DP_OP_422J2_124_3477_U924 ( .A(DP_OP_422J2_124_3477_n2679), .B(
        DP_OP_422J2_124_3477_n2672), .CI(DP_OP_422J2_124_3477_n1837), .CO(
        DP_OP_422J2_124_3477_n1653), .S(DP_OP_422J2_124_3477_n1654) );
  FADDX1_HVT DP_OP_422J2_124_3477_U923 ( .A(DP_OP_422J2_124_3477_n2246), .B(
        DP_OP_422J2_124_3477_n2897), .CI(DP_OP_422J2_124_3477_n2239), .CO(
        DP_OP_422J2_124_3477_n1651), .S(DP_OP_422J2_124_3477_n1652) );
  FADDX1_HVT DP_OP_422J2_124_3477_U922 ( .A(DP_OP_422J2_124_3477_n2459), .B(
        DP_OP_422J2_124_3477_n2283), .CI(DP_OP_422J2_124_3477_n2195), .CO(
        DP_OP_422J2_124_3477_n1649), .S(DP_OP_422J2_124_3477_n1650) );
  FADDX1_HVT DP_OP_422J2_124_3477_U921 ( .A(DP_OP_422J2_124_3477_n2714), .B(
        DP_OP_422J2_124_3477_n2765), .CI(DP_OP_422J2_124_3477_n2371), .CO(
        DP_OP_422J2_124_3477_n1647), .S(DP_OP_422J2_124_3477_n1648) );
  FADDX1_HVT DP_OP_422J2_124_3477_U920 ( .A(DP_OP_422J2_124_3477_n2547), .B(
        DP_OP_422J2_124_3477_n2809), .CI(DP_OP_422J2_124_3477_n2012), .CO(
        DP_OP_422J2_124_3477_n1645), .S(DP_OP_422J2_124_3477_n1646) );
  FADDX1_HVT DP_OP_422J2_124_3477_U919 ( .A(DP_OP_422J2_124_3477_n1939), .B(
        DP_OP_422J2_124_3477_n2853), .CI(DP_OP_422J2_124_3477_n2802), .CO(
        DP_OP_422J2_124_3477_n1643), .S(DP_OP_422J2_124_3477_n1644) );
  FADDX1_HVT DP_OP_422J2_124_3477_U918 ( .A(DP_OP_422J2_124_3477_n2158), .B(
        DP_OP_422J2_124_3477_n1976), .CI(DP_OP_422J2_124_3477_n2816), .CO(
        DP_OP_422J2_124_3477_n1641), .S(DP_OP_422J2_124_3477_n1642) );
  FADDX1_HVT DP_OP_422J2_124_3477_U917 ( .A(DP_OP_422J2_124_3477_n2408), .B(
        DP_OP_422J2_124_3477_n2378), .CI(DP_OP_422J2_124_3477_n2628), .CO(
        DP_OP_422J2_124_3477_n1639), .S(DP_OP_422J2_124_3477_n1640) );
  FADDX1_HVT DP_OP_422J2_124_3477_U916 ( .A(DP_OP_422J2_124_3477_n2019), .B(
        DP_OP_422J2_124_3477_n2904), .CI(DP_OP_422J2_124_3477_n2721), .CO(
        DP_OP_422J2_124_3477_n1637), .S(DP_OP_422J2_124_3477_n1638) );
  FADDX1_HVT DP_OP_422J2_124_3477_U915 ( .A(DP_OP_422J2_124_3477_n1932), .B(
        DP_OP_422J2_124_3477_n1881), .CI(DP_OP_422J2_124_3477_n1747), .CO(
        DP_OP_422J2_124_3477_n1635), .S(DP_OP_422J2_124_3477_n1636) );
  FADDX1_HVT DP_OP_422J2_124_3477_U914 ( .A(DP_OP_422J2_124_3477_n1686), .B(
        DP_OP_422J2_124_3477_n1745), .CI(DP_OP_422J2_124_3477_n1729), .CO(
        DP_OP_422J2_124_3477_n1633), .S(DP_OP_422J2_124_3477_n1634) );
  FADDX1_HVT DP_OP_422J2_124_3477_U913 ( .A(DP_OP_422J2_124_3477_n1743), .B(
        DP_OP_422J2_124_3477_n1731), .CI(DP_OP_422J2_124_3477_n1741), .CO(
        DP_OP_422J2_124_3477_n1631), .S(DP_OP_422J2_124_3477_n1632) );
  FADDX1_HVT DP_OP_422J2_124_3477_U912 ( .A(DP_OP_422J2_124_3477_n1733), .B(
        DP_OP_422J2_124_3477_n1735), .CI(DP_OP_422J2_124_3477_n1737), .CO(
        DP_OP_422J2_124_3477_n1629), .S(DP_OP_422J2_124_3477_n1630) );
  FADDX1_HVT DP_OP_422J2_124_3477_U911 ( .A(DP_OP_422J2_124_3477_n1739), .B(
        DP_OP_422J2_124_3477_n1727), .CI(DP_OP_422J2_124_3477_n1725), .CO(
        DP_OP_422J2_124_3477_n1627), .S(DP_OP_422J2_124_3477_n1628) );
  FADDX1_HVT DP_OP_422J2_124_3477_U910 ( .A(DP_OP_422J2_124_3477_n1723), .B(
        DP_OP_422J2_124_3477_n1717), .CI(DP_OP_422J2_124_3477_n1715), .CO(
        DP_OP_422J2_124_3477_n1625), .S(DP_OP_422J2_124_3477_n1626) );
  FADDX1_HVT DP_OP_422J2_124_3477_U909 ( .A(DP_OP_422J2_124_3477_n1721), .B(
        DP_OP_422J2_124_3477_n1719), .CI(DP_OP_422J2_124_3477_n1668), .CO(
        DP_OP_422J2_124_3477_n1623), .S(DP_OP_422J2_124_3477_n1624) );
  FADDX1_HVT DP_OP_422J2_124_3477_U908 ( .A(DP_OP_422J2_124_3477_n1678), .B(
        DP_OP_422J2_124_3477_n1664), .CI(DP_OP_422J2_124_3477_n1660), .CO(
        DP_OP_422J2_124_3477_n1621), .S(DP_OP_422J2_124_3477_n1622) );
  FADDX1_HVT DP_OP_422J2_124_3477_U907 ( .A(DP_OP_422J2_124_3477_n1676), .B(
        DP_OP_422J2_124_3477_n1670), .CI(DP_OP_422J2_124_3477_n1662), .CO(
        DP_OP_422J2_124_3477_n1619), .S(DP_OP_422J2_124_3477_n1620) );
  FADDX1_HVT DP_OP_422J2_124_3477_U906 ( .A(DP_OP_422J2_124_3477_n1684), .B(
        DP_OP_422J2_124_3477_n1666), .CI(DP_OP_422J2_124_3477_n1672), .CO(
        DP_OP_422J2_124_3477_n1617), .S(DP_OP_422J2_124_3477_n1618) );
  FADDX1_HVT DP_OP_422J2_124_3477_U905 ( .A(DP_OP_422J2_124_3477_n1682), .B(
        DP_OP_422J2_124_3477_n1674), .CI(DP_OP_422J2_124_3477_n1680), .CO(
        DP_OP_422J2_124_3477_n1615), .S(DP_OP_422J2_124_3477_n1616) );
  FADDX1_HVT DP_OP_422J2_124_3477_U904 ( .A(DP_OP_422J2_124_3477_n1658), .B(
        DP_OP_422J2_124_3477_n1644), .CI(DP_OP_422J2_124_3477_n1713), .CO(
        DP_OP_422J2_124_3477_n1613), .S(DP_OP_422J2_124_3477_n1614) );
  FADDX1_HVT DP_OP_422J2_124_3477_U903 ( .A(DP_OP_422J2_124_3477_n1656), .B(
        DP_OP_422J2_124_3477_n1646), .CI(DP_OP_422J2_124_3477_n1642), .CO(
        DP_OP_422J2_124_3477_n1611), .S(DP_OP_422J2_124_3477_n1612) );
  FADDX1_HVT DP_OP_422J2_124_3477_U902 ( .A(DP_OP_422J2_124_3477_n1654), .B(
        DP_OP_422J2_124_3477_n1648), .CI(DP_OP_422J2_124_3477_n1640), .CO(
        DP_OP_422J2_124_3477_n1609), .S(DP_OP_422J2_124_3477_n1610) );
  FADDX1_HVT DP_OP_422J2_124_3477_U901 ( .A(DP_OP_422J2_124_3477_n1652), .B(
        DP_OP_422J2_124_3477_n1650), .CI(DP_OP_422J2_124_3477_n1638), .CO(
        DP_OP_422J2_124_3477_n1607), .S(DP_OP_422J2_124_3477_n1608) );
  FADDX1_HVT DP_OP_422J2_124_3477_U900 ( .A(DP_OP_422J2_124_3477_n1636), .B(
        DP_OP_422J2_124_3477_n1711), .CI(DP_OP_422J2_124_3477_n1709), .CO(
        DP_OP_422J2_124_3477_n1605), .S(DP_OP_422J2_124_3477_n1606) );
  FADDX1_HVT DP_OP_422J2_124_3477_U899 ( .A(DP_OP_422J2_124_3477_n1707), .B(
        DP_OP_422J2_124_3477_n1634), .CI(DP_OP_422J2_124_3477_n1632), .CO(
        DP_OP_422J2_124_3477_n1603), .S(DP_OP_422J2_124_3477_n1604) );
  FADDX1_HVT DP_OP_422J2_124_3477_U898 ( .A(DP_OP_422J2_124_3477_n1705), .B(
        DP_OP_422J2_124_3477_n1630), .CI(DP_OP_422J2_124_3477_n1628), .CO(
        DP_OP_422J2_124_3477_n1601), .S(DP_OP_422J2_124_3477_n1602) );
  FADDX1_HVT DP_OP_422J2_124_3477_U897 ( .A(DP_OP_422J2_124_3477_n1703), .B(
        DP_OP_422J2_124_3477_n1701), .CI(DP_OP_422J2_124_3477_n1699), .CO(
        DP_OP_422J2_124_3477_n1599), .S(DP_OP_422J2_124_3477_n1600) );
  FADDX1_HVT DP_OP_422J2_124_3477_U896 ( .A(DP_OP_422J2_124_3477_n1697), .B(
        DP_OP_422J2_124_3477_n1626), .CI(DP_OP_422J2_124_3477_n1624), .CO(
        DP_OP_422J2_124_3477_n1597), .S(DP_OP_422J2_124_3477_n1598) );
  FADDX1_HVT DP_OP_422J2_124_3477_U895 ( .A(DP_OP_422J2_124_3477_n1622), .B(
        DP_OP_422J2_124_3477_n1616), .CI(DP_OP_422J2_124_3477_n1618), .CO(
        DP_OP_422J2_124_3477_n1595), .S(DP_OP_422J2_124_3477_n1596) );
  FADDX1_HVT DP_OP_422J2_124_3477_U894 ( .A(DP_OP_422J2_124_3477_n1620), .B(
        DP_OP_422J2_124_3477_n1614), .CI(DP_OP_422J2_124_3477_n1612), .CO(
        DP_OP_422J2_124_3477_n1593), .S(DP_OP_422J2_124_3477_n1594) );
  FADDX1_HVT DP_OP_422J2_124_3477_U893 ( .A(DP_OP_422J2_124_3477_n1610), .B(
        DP_OP_422J2_124_3477_n1608), .CI(DP_OP_422J2_124_3477_n1695), .CO(
        DP_OP_422J2_124_3477_n1591), .S(DP_OP_422J2_124_3477_n1592) );
  FADDX1_HVT DP_OP_422J2_124_3477_U892 ( .A(DP_OP_422J2_124_3477_n1606), .B(
        DP_OP_422J2_124_3477_n1693), .CI(DP_OP_422J2_124_3477_n1604), .CO(
        DP_OP_422J2_124_3477_n1589), .S(DP_OP_422J2_124_3477_n1590) );
  FADDX1_HVT DP_OP_422J2_124_3477_U891 ( .A(DP_OP_422J2_124_3477_n1691), .B(
        DP_OP_422J2_124_3477_n1602), .CI(DP_OP_422J2_124_3477_n1600), .CO(
        DP_OP_422J2_124_3477_n1587), .S(DP_OP_422J2_124_3477_n1588) );
  FADDX1_HVT DP_OP_422J2_124_3477_U890 ( .A(DP_OP_422J2_124_3477_n1689), .B(
        DP_OP_422J2_124_3477_n1598), .CI(DP_OP_422J2_124_3477_n1596), .CO(
        DP_OP_422J2_124_3477_n1585), .S(DP_OP_422J2_124_3477_n1586) );
  FADDX1_HVT DP_OP_422J2_124_3477_U889 ( .A(DP_OP_422J2_124_3477_n1594), .B(
        DP_OP_422J2_124_3477_n1592), .CI(DP_OP_422J2_124_3477_n1590), .CO(
        DP_OP_422J2_124_3477_n1583), .S(DP_OP_422J2_124_3477_n1584) );
  FADDX1_HVT DP_OP_422J2_124_3477_U888 ( .A(DP_OP_422J2_124_3477_n1687), .B(
        DP_OP_422J2_124_3477_n1588), .CI(DP_OP_422J2_124_3477_n1586), .CO(
        DP_OP_422J2_124_3477_n1581), .S(DP_OP_422J2_124_3477_n1582) );
  FADDX1_HVT DP_OP_422J2_124_3477_U886 ( .A(DP_OP_422J2_124_3477_n2706), .B(
        DP_OP_422J2_124_3477_n1829), .CI(DP_OP_422J2_124_3477_n2750), .CO(
        DP_OP_422J2_124_3477_n1577), .S(DP_OP_422J2_124_3477_n1578) );
  FADDX1_HVT DP_OP_422J2_124_3477_U885 ( .A(DP_OP_422J2_124_3477_n2092), .B(
        DP_OP_422J2_124_3477_n2576), .CI(DP_OP_422J2_124_3477_n1961), .CO(
        DP_OP_422J2_124_3477_n1575), .S(DP_OP_422J2_124_3477_n1576) );
  FADDX1_HVT DP_OP_422J2_124_3477_U884 ( .A(DP_OP_422J2_124_3477_n2838), .B(
        DP_OP_422J2_124_3477_n2488), .CI(DP_OP_422J2_124_3477_n1917), .CO(
        DP_OP_422J2_124_3477_n1573), .S(DP_OP_422J2_124_3477_n1574) );
  FADDX1_HVT DP_OP_422J2_124_3477_U883 ( .A(DP_OP_422J2_124_3477_n2620), .B(
        DP_OP_422J2_124_3477_n2180), .CI(DP_OP_422J2_124_3477_n2532), .CO(
        DP_OP_422J2_124_3477_n1571), .S(DP_OP_422J2_124_3477_n1572) );
  FADDX1_HVT DP_OP_422J2_124_3477_U882 ( .A(DP_OP_422J2_124_3477_n2794), .B(
        DP_OP_422J2_124_3477_n2444), .CI(DP_OP_422J2_124_3477_n2048), .CO(
        DP_OP_422J2_124_3477_n1569), .S(DP_OP_422J2_124_3477_n1570) );
  FADDX1_HVT DP_OP_422J2_124_3477_U881 ( .A(DP_OP_422J2_124_3477_n1873), .B(
        DP_OP_422J2_124_3477_n2268), .CI(DP_OP_422J2_124_3477_n2882), .CO(
        DP_OP_422J2_124_3477_n1567), .S(DP_OP_422J2_124_3477_n1568) );
  FADDX1_HVT DP_OP_422J2_124_3477_U880 ( .A(DP_OP_422J2_124_3477_n2136), .B(
        DP_OP_422J2_124_3477_n2312), .CI(DP_OP_422J2_124_3477_n2664), .CO(
        DP_OP_422J2_124_3477_n1565), .S(DP_OP_422J2_124_3477_n1566) );
  FADDX1_HVT DP_OP_422J2_124_3477_U879 ( .A(DP_OP_422J2_124_3477_n2356), .B(
        DP_OP_422J2_124_3477_n2400), .CI(DP_OP_422J2_124_3477_n2201), .CO(
        DP_OP_422J2_124_3477_n1563), .S(DP_OP_422J2_124_3477_n1564) );
  FADDX1_HVT DP_OP_422J2_124_3477_U878 ( .A(DP_OP_422J2_124_3477_n2113), .B(
        DP_OP_422J2_124_3477_n1968), .CI(DP_OP_422J2_124_3477_n2275), .CO(
        DP_OP_422J2_124_3477_n1561), .S(DP_OP_422J2_124_3477_n1562) );
  FADDX1_HVT DP_OP_422J2_124_3477_U877 ( .A(DP_OP_422J2_124_3477_n2845), .B(
        DP_OP_422J2_124_3477_n2539), .CI(DP_OP_422J2_124_3477_n2069), .CO(
        DP_OP_422J2_124_3477_n1559), .S(DP_OP_422J2_124_3477_n1560) );
  FADDX1_HVT DP_OP_422J2_124_3477_U876 ( .A(DP_OP_422J2_124_3477_n2597), .B(
        DP_OP_422J2_124_3477_n2150), .CI(DP_OP_422J2_124_3477_n2143), .CO(
        DP_OP_422J2_124_3477_n1557), .S(DP_OP_422J2_124_3477_n1558) );
  FADDX1_HVT DP_OP_422J2_124_3477_U875 ( .A(DP_OP_422J2_124_3477_n2553), .B(
        DP_OP_422J2_124_3477_n2727), .CI(DP_OP_422J2_124_3477_n2289), .CO(
        DP_OP_422J2_124_3477_n1555), .S(DP_OP_422J2_124_3477_n1556) );
  FADDX1_HVT DP_OP_422J2_124_3477_U874 ( .A(DP_OP_422J2_124_3477_n2421), .B(
        DP_OP_422J2_124_3477_n2414), .CI(DP_OP_422J2_124_3477_n2583), .CO(
        DP_OP_422J2_124_3477_n1553), .S(DP_OP_422J2_124_3477_n1554) );
  FADDX1_HVT DP_OP_422J2_124_3477_U873 ( .A(DP_OP_422J2_124_3477_n2889), .B(
        DP_OP_422J2_124_3477_n1580), .CI(DP_OP_422J2_124_3477_n2509), .CO(
        DP_OP_422J2_124_3477_n1551), .S(DP_OP_422J2_124_3477_n1552) );
  FADDX1_HVT DP_OP_422J2_124_3477_U872 ( .A(DP_OP_422J2_124_3477_n2333), .B(
        DP_OP_422J2_124_3477_n2224), .CI(DP_OP_422J2_124_3477_n1894), .CO(
        DP_OP_422J2_124_3477_n1549), .S(DP_OP_422J2_124_3477_n1550) );
  FADDX1_HVT DP_OP_422J2_124_3477_U871 ( .A(DP_OP_422J2_124_3477_n2465), .B(
        DP_OP_422J2_124_3477_n1785), .CI(DP_OP_422J2_124_3477_n2771), .CO(
        DP_OP_422J2_124_3477_n1547), .S(DP_OP_422J2_124_3477_n1548) );
  FADDX1_HVT DP_OP_422J2_124_3477_U870 ( .A(DP_OP_422J2_124_3477_n1850), .B(
        DP_OP_422J2_124_3477_n2025), .CI(DP_OP_422J2_124_3477_n2451), .CO(
        DP_OP_422J2_124_3477_n1545), .S(DP_OP_422J2_124_3477_n1546) );
  FADDX1_HVT DP_OP_422J2_124_3477_U869 ( .A(DP_OP_422J2_124_3477_n2641), .B(
        DP_OP_422J2_124_3477_n2502), .CI(DP_OP_422J2_124_3477_n2859), .CO(
        DP_OP_422J2_124_3477_n1543), .S(DP_OP_422J2_124_3477_n1544) );
  FADDX1_HVT DP_OP_422J2_124_3477_U868 ( .A(DP_OP_422J2_124_3477_n2685), .B(
        DP_OP_422J2_124_3477_n2062), .CI(DP_OP_422J2_124_3477_n2231), .CO(
        DP_OP_422J2_124_3477_n1541), .S(DP_OP_422J2_124_3477_n1542) );
  FADDX1_HVT DP_OP_422J2_124_3477_U867 ( .A(DP_OP_422J2_124_3477_n2326), .B(
        DP_OP_422J2_124_3477_n1982), .CI(DP_OP_422J2_124_3477_n2099), .CO(
        DP_OP_422J2_124_3477_n1539), .S(DP_OP_422J2_124_3477_n1540) );
  FADDX1_HVT DP_OP_422J2_124_3477_U866 ( .A(DP_OP_422J2_124_3477_n2757), .B(
        DP_OP_422J2_124_3477_n2590), .CI(DP_OP_422J2_124_3477_n1843), .CO(
        DP_OP_422J2_124_3477_n1537), .S(DP_OP_422J2_124_3477_n1538) );
  FADDX1_HVT DP_OP_422J2_124_3477_U865 ( .A(DP_OP_422J2_124_3477_n2634), .B(
        DP_OP_422J2_124_3477_n2495), .CI(DP_OP_422J2_124_3477_n2106), .CO(
        DP_OP_422J2_124_3477_n1535), .S(DP_OP_422J2_124_3477_n1536) );
  FADDX1_HVT DP_OP_422J2_124_3477_U864 ( .A(DP_OP_422J2_124_3477_n1887), .B(
        DP_OP_422J2_124_3477_n2319), .CI(DP_OP_422J2_124_3477_n2187), .CO(
        DP_OP_422J2_124_3477_n1533), .S(DP_OP_422J2_124_3477_n1534) );
  FADDX1_HVT DP_OP_422J2_124_3477_U863 ( .A(DP_OP_422J2_124_3477_n2363), .B(
        DP_OP_422J2_124_3477_n2055), .CI(DP_OP_422J2_124_3477_n1924), .CO(
        DP_OP_422J2_124_3477_n1531), .S(DP_OP_422J2_124_3477_n1532) );
  FADDX1_HVT DP_OP_422J2_124_3477_U862 ( .A(DP_OP_422J2_124_3477_n2678), .B(
        DP_OP_422J2_124_3477_n2671), .CI(DP_OP_422J2_124_3477_n1836), .CO(
        DP_OP_422J2_124_3477_n1529), .S(DP_OP_422J2_124_3477_n1530) );
  FADDX1_HVT DP_OP_422J2_124_3477_U861 ( .A(DP_OP_422J2_124_3477_n2245), .B(
        DP_OP_422J2_124_3477_n2896), .CI(DP_OP_422J2_124_3477_n2238), .CO(
        DP_OP_422J2_124_3477_n1527), .S(DP_OP_422J2_124_3477_n1528) );
  FADDX1_HVT DP_OP_422J2_124_3477_U860 ( .A(DP_OP_422J2_124_3477_n2458), .B(
        DP_OP_422J2_124_3477_n2282), .CI(DP_OP_422J2_124_3477_n2370), .CO(
        DP_OP_422J2_124_3477_n1525), .S(DP_OP_422J2_124_3477_n1526) );
  FADDX1_HVT DP_OP_422J2_124_3477_U859 ( .A(DP_OP_422J2_124_3477_n2713), .B(
        DP_OP_422J2_124_3477_n2764), .CI(DP_OP_422J2_124_3477_n2011), .CO(
        DP_OP_422J2_124_3477_n1523), .S(DP_OP_422J2_124_3477_n1524) );
  FADDX1_HVT DP_OP_422J2_124_3477_U858 ( .A(DP_OP_422J2_124_3477_n2546), .B(
        DP_OP_422J2_124_3477_n2808), .CI(DP_OP_422J2_124_3477_n2194), .CO(
        DP_OP_422J2_124_3477_n1521), .S(DP_OP_422J2_124_3477_n1522) );
  FADDX1_HVT DP_OP_422J2_124_3477_U857 ( .A(DP_OP_422J2_124_3477_n1938), .B(
        DP_OP_422J2_124_3477_n2852), .CI(DP_OP_422J2_124_3477_n2627), .CO(
        DP_OP_422J2_124_3477_n1519), .S(DP_OP_422J2_124_3477_n1520) );
  FADDX1_HVT DP_OP_422J2_124_3477_U856 ( .A(DP_OP_422J2_124_3477_n2018), .B(
        DP_OP_422J2_124_3477_n1975), .CI(DP_OP_422J2_124_3477_n2815), .CO(
        DP_OP_422J2_124_3477_n1517), .S(DP_OP_422J2_124_3477_n1518) );
  FADDX1_HVT DP_OP_422J2_124_3477_U855 ( .A(DP_OP_422J2_124_3477_n2157), .B(
        DP_OP_422J2_124_3477_n2720), .CI(DP_OP_422J2_124_3477_n2801), .CO(
        DP_OP_422J2_124_3477_n1515), .S(DP_OP_422J2_124_3477_n1516) );
  FADDX1_HVT DP_OP_422J2_124_3477_U854 ( .A(DP_OP_422J2_124_3477_n2407), .B(
        DP_OP_422J2_124_3477_n2377), .CI(DP_OP_422J2_124_3477_n2903), .CO(
        DP_OP_422J2_124_3477_n1513), .S(DP_OP_422J2_124_3477_n1514) );
  FADDX1_HVT DP_OP_422J2_124_3477_U853 ( .A(DP_OP_422J2_124_3477_n1931), .B(
        DP_OP_422J2_124_3477_n1880), .CI(DP_OP_422J2_124_3477_n1685), .CO(
        DP_OP_422J2_124_3477_n1511), .S(DP_OP_422J2_124_3477_n1512) );
  FADDX1_HVT DP_OP_422J2_124_3477_U852 ( .A(DP_OP_422J2_124_3477_n1683), .B(
        DP_OP_422J2_124_3477_n1661), .CI(DP_OP_422J2_124_3477_n1659), .CO(
        DP_OP_422J2_124_3477_n1509), .S(DP_OP_422J2_124_3477_n1510) );
  FADDX1_HVT DP_OP_422J2_124_3477_U851 ( .A(DP_OP_422J2_124_3477_n1681), .B(
        DP_OP_422J2_124_3477_n1665), .CI(DP_OP_422J2_124_3477_n1663), .CO(
        DP_OP_422J2_124_3477_n1507), .S(DP_OP_422J2_124_3477_n1508) );
  FADDX1_HVT DP_OP_422J2_124_3477_U850 ( .A(DP_OP_422J2_124_3477_n1679), .B(
        DP_OP_422J2_124_3477_n1667), .CI(DP_OP_422J2_124_3477_n1669), .CO(
        DP_OP_422J2_124_3477_n1505), .S(DP_OP_422J2_124_3477_n1506) );
  FADDX1_HVT DP_OP_422J2_124_3477_U849 ( .A(DP_OP_422J2_124_3477_n1677), .B(
        DP_OP_422J2_124_3477_n1671), .CI(DP_OP_422J2_124_3477_n1673), .CO(
        DP_OP_422J2_124_3477_n1503), .S(DP_OP_422J2_124_3477_n1504) );
  FADDX1_HVT DP_OP_422J2_124_3477_U848 ( .A(DP_OP_422J2_124_3477_n1675), .B(
        DP_OP_422J2_124_3477_n1657), .CI(DP_OP_422J2_124_3477_n1655), .CO(
        DP_OP_422J2_124_3477_n1501), .S(DP_OP_422J2_124_3477_n1502) );
  FADDX1_HVT DP_OP_422J2_124_3477_U847 ( .A(DP_OP_422J2_124_3477_n1653), .B(
        DP_OP_422J2_124_3477_n1574), .CI(DP_OP_422J2_124_3477_n1564), .CO(
        DP_OP_422J2_124_3477_n1499), .S(DP_OP_422J2_124_3477_n1500) );
  FADDX1_HVT DP_OP_422J2_124_3477_U846 ( .A(DP_OP_422J2_124_3477_n1651), .B(
        DP_OP_422J2_124_3477_n1572), .CI(DP_OP_422J2_124_3477_n1639), .CO(
        DP_OP_422J2_124_3477_n1497), .S(DP_OP_422J2_124_3477_n1498) );
  FADDX1_HVT DP_OP_422J2_124_3477_U845 ( .A(DP_OP_422J2_124_3477_n1649), .B(
        DP_OP_422J2_124_3477_n1566), .CI(DP_OP_422J2_124_3477_n1637), .CO(
        DP_OP_422J2_124_3477_n1495), .S(DP_OP_422J2_124_3477_n1496) );
  FADDX1_HVT DP_OP_422J2_124_3477_U844 ( .A(DP_OP_422J2_124_3477_n1647), .B(
        DP_OP_422J2_124_3477_n1568), .CI(DP_OP_422J2_124_3477_n1641), .CO(
        DP_OP_422J2_124_3477_n1493), .S(DP_OP_422J2_124_3477_n1494) );
  FADDX1_HVT DP_OP_422J2_124_3477_U843 ( .A(DP_OP_422J2_124_3477_n1645), .B(
        DP_OP_422J2_124_3477_n1570), .CI(DP_OP_422J2_124_3477_n1576), .CO(
        DP_OP_422J2_124_3477_n1491), .S(DP_OP_422J2_124_3477_n1492) );
  FADDX1_HVT DP_OP_422J2_124_3477_U842 ( .A(DP_OP_422J2_124_3477_n1643), .B(
        DP_OP_422J2_124_3477_n1578), .CI(DP_OP_422J2_124_3477_n1635), .CO(
        DP_OP_422J2_124_3477_n1489), .S(DP_OP_422J2_124_3477_n1490) );
  FADDX1_HVT DP_OP_422J2_124_3477_U841 ( .A(DP_OP_422J2_124_3477_n1556), .B(
        DP_OP_422J2_124_3477_n1538), .CI(DP_OP_422J2_124_3477_n1536), .CO(
        DP_OP_422J2_124_3477_n1487), .S(DP_OP_422J2_124_3477_n1488) );
  FADDX1_HVT DP_OP_422J2_124_3477_U840 ( .A(DP_OP_422J2_124_3477_n1560), .B(
        DP_OP_422J2_124_3477_n1540), .CI(DP_OP_422J2_124_3477_n1542), .CO(
        DP_OP_422J2_124_3477_n1485), .S(DP_OP_422J2_124_3477_n1486) );
  FADDX1_HVT DP_OP_422J2_124_3477_U839 ( .A(DP_OP_422J2_124_3477_n1554), .B(
        DP_OP_422J2_124_3477_n1548), .CI(DP_OP_422J2_124_3477_n1546), .CO(
        DP_OP_422J2_124_3477_n1483), .S(DP_OP_422J2_124_3477_n1484) );
  FADDX1_HVT DP_OP_422J2_124_3477_U838 ( .A(DP_OP_422J2_124_3477_n1550), .B(
        DP_OP_422J2_124_3477_n1544), .CI(DP_OP_422J2_124_3477_n1562), .CO(
        DP_OP_422J2_124_3477_n1481), .S(DP_OP_422J2_124_3477_n1482) );
  FADDX1_HVT DP_OP_422J2_124_3477_U837 ( .A(DP_OP_422J2_124_3477_n1552), .B(
        DP_OP_422J2_124_3477_n1558), .CI(DP_OP_422J2_124_3477_n1534), .CO(
        DP_OP_422J2_124_3477_n1479), .S(DP_OP_422J2_124_3477_n1480) );
  FADDX1_HVT DP_OP_422J2_124_3477_U836 ( .A(DP_OP_422J2_124_3477_n1532), .B(
        DP_OP_422J2_124_3477_n1520), .CI(DP_OP_422J2_124_3477_n1516), .CO(
        DP_OP_422J2_124_3477_n1477), .S(DP_OP_422J2_124_3477_n1478) );
  FADDX1_HVT DP_OP_422J2_124_3477_U835 ( .A(DP_OP_422J2_124_3477_n1530), .B(
        DP_OP_422J2_124_3477_n1524), .CI(DP_OP_422J2_124_3477_n1514), .CO(
        DP_OP_422J2_124_3477_n1475), .S(DP_OP_422J2_124_3477_n1476) );
  FADDX1_HVT DP_OP_422J2_124_3477_U834 ( .A(DP_OP_422J2_124_3477_n1528), .B(
        DP_OP_422J2_124_3477_n1522), .CI(DP_OP_422J2_124_3477_n1518), .CO(
        DP_OP_422J2_124_3477_n1473), .S(DP_OP_422J2_124_3477_n1474) );
  FADDX1_HVT DP_OP_422J2_124_3477_U833 ( .A(DP_OP_422J2_124_3477_n1526), .B(
        DP_OP_422J2_124_3477_n1512), .CI(DP_OP_422J2_124_3477_n1633), .CO(
        DP_OP_422J2_124_3477_n1471), .S(DP_OP_422J2_124_3477_n1472) );
  FADDX1_HVT DP_OP_422J2_124_3477_U832 ( .A(DP_OP_422J2_124_3477_n1631), .B(
        DP_OP_422J2_124_3477_n1629), .CI(DP_OP_422J2_124_3477_n1627), .CO(
        DP_OP_422J2_124_3477_n1469), .S(DP_OP_422J2_124_3477_n1470) );
  FADDX1_HVT DP_OP_422J2_124_3477_U831 ( .A(DP_OP_422J2_124_3477_n1625), .B(
        DP_OP_422J2_124_3477_n1623), .CI(DP_OP_422J2_124_3477_n1621), .CO(
        DP_OP_422J2_124_3477_n1467), .S(DP_OP_422J2_124_3477_n1468) );
  FADDX1_HVT DP_OP_422J2_124_3477_U830 ( .A(DP_OP_422J2_124_3477_n1619), .B(
        DP_OP_422J2_124_3477_n1510), .CI(DP_OP_422J2_124_3477_n1502), .CO(
        DP_OP_422J2_124_3477_n1465), .S(DP_OP_422J2_124_3477_n1466) );
  FADDX1_HVT DP_OP_422J2_124_3477_U829 ( .A(DP_OP_422J2_124_3477_n1617), .B(
        DP_OP_422J2_124_3477_n1506), .CI(DP_OP_422J2_124_3477_n1504), .CO(
        DP_OP_422J2_124_3477_n1463), .S(DP_OP_422J2_124_3477_n1464) );
  FADDX1_HVT DP_OP_422J2_124_3477_U828 ( .A(DP_OP_422J2_124_3477_n1615), .B(
        DP_OP_422J2_124_3477_n1508), .CI(DP_OP_422J2_124_3477_n1613), .CO(
        DP_OP_422J2_124_3477_n1461), .S(DP_OP_422J2_124_3477_n1462) );
  FADDX1_HVT DP_OP_422J2_124_3477_U827 ( .A(DP_OP_422J2_124_3477_n1611), .B(
        DP_OP_422J2_124_3477_n1494), .CI(DP_OP_422J2_124_3477_n1490), .CO(
        DP_OP_422J2_124_3477_n1459), .S(DP_OP_422J2_124_3477_n1460) );
  FADDX1_HVT DP_OP_422J2_124_3477_U826 ( .A(DP_OP_422J2_124_3477_n1609), .B(
        DP_OP_422J2_124_3477_n1496), .CI(DP_OP_422J2_124_3477_n1492), .CO(
        DP_OP_422J2_124_3477_n1457), .S(DP_OP_422J2_124_3477_n1458) );
  FADDX1_HVT DP_OP_422J2_124_3477_U825 ( .A(DP_OP_422J2_124_3477_n1500), .B(
        DP_OP_422J2_124_3477_n1607), .CI(DP_OP_422J2_124_3477_n1498), .CO(
        DP_OP_422J2_124_3477_n1455), .S(DP_OP_422J2_124_3477_n1456) );
  FADDX1_HVT DP_OP_422J2_124_3477_U824 ( .A(DP_OP_422J2_124_3477_n1484), .B(
        DP_OP_422J2_124_3477_n1480), .CI(DP_OP_422J2_124_3477_n1605), .CO(
        DP_OP_422J2_124_3477_n1453), .S(DP_OP_422J2_124_3477_n1454) );
  FADDX1_HVT DP_OP_422J2_124_3477_U823 ( .A(DP_OP_422J2_124_3477_n1488), .B(
        DP_OP_422J2_124_3477_n1486), .CI(DP_OP_422J2_124_3477_n1482), .CO(
        DP_OP_422J2_124_3477_n1451), .S(DP_OP_422J2_124_3477_n1452) );
  FADDX1_HVT DP_OP_422J2_124_3477_U822 ( .A(DP_OP_422J2_124_3477_n1478), .B(
        DP_OP_422J2_124_3477_n1476), .CI(DP_OP_422J2_124_3477_n1474), .CO(
        DP_OP_422J2_124_3477_n1449), .S(DP_OP_422J2_124_3477_n1450) );
  FADDX1_HVT DP_OP_422J2_124_3477_U821 ( .A(DP_OP_422J2_124_3477_n1472), .B(
        DP_OP_422J2_124_3477_n1603), .CI(DP_OP_422J2_124_3477_n1601), .CO(
        DP_OP_422J2_124_3477_n1447), .S(DP_OP_422J2_124_3477_n1448) );
  FADDX1_HVT DP_OP_422J2_124_3477_U820 ( .A(DP_OP_422J2_124_3477_n1470), .B(
        DP_OP_422J2_124_3477_n1599), .CI(DP_OP_422J2_124_3477_n1597), .CO(
        DP_OP_422J2_124_3477_n1445), .S(DP_OP_422J2_124_3477_n1446) );
  FADDX1_HVT DP_OP_422J2_124_3477_U819 ( .A(DP_OP_422J2_124_3477_n1468), .B(
        DP_OP_422J2_124_3477_n1464), .CI(DP_OP_422J2_124_3477_n1466), .CO(
        DP_OP_422J2_124_3477_n1443), .S(DP_OP_422J2_124_3477_n1444) );
  FADDX1_HVT DP_OP_422J2_124_3477_U818 ( .A(DP_OP_422J2_124_3477_n1595), .B(
        DP_OP_422J2_124_3477_n1462), .CI(DP_OP_422J2_124_3477_n1593), .CO(
        DP_OP_422J2_124_3477_n1441), .S(DP_OP_422J2_124_3477_n1442) );
  FADDX1_HVT DP_OP_422J2_124_3477_U817 ( .A(DP_OP_422J2_124_3477_n1460), .B(
        DP_OP_422J2_124_3477_n1458), .CI(DP_OP_422J2_124_3477_n1591), .CO(
        DP_OP_422J2_124_3477_n1439), .S(DP_OP_422J2_124_3477_n1440) );
  FADDX1_HVT DP_OP_422J2_124_3477_U816 ( .A(DP_OP_422J2_124_3477_n1456), .B(
        DP_OP_422J2_124_3477_n1452), .CI(DP_OP_422J2_124_3477_n1454), .CO(
        DP_OP_422J2_124_3477_n1437), .S(DP_OP_422J2_124_3477_n1438) );
  FADDX1_HVT DP_OP_422J2_124_3477_U815 ( .A(DP_OP_422J2_124_3477_n1450), .B(
        DP_OP_422J2_124_3477_n1589), .CI(DP_OP_422J2_124_3477_n1448), .CO(
        DP_OP_422J2_124_3477_n1435), .S(DP_OP_422J2_124_3477_n1436) );
  FADDX1_HVT DP_OP_422J2_124_3477_U814 ( .A(DP_OP_422J2_124_3477_n1587), .B(
        DP_OP_422J2_124_3477_n1446), .CI(DP_OP_422J2_124_3477_n1585), .CO(
        DP_OP_422J2_124_3477_n1433), .S(DP_OP_422J2_124_3477_n1434) );
  FADDX1_HVT DP_OP_422J2_124_3477_U813 ( .A(DP_OP_422J2_124_3477_n1444), .B(
        DP_OP_422J2_124_3477_n1442), .CI(DP_OP_422J2_124_3477_n1440), .CO(
        DP_OP_422J2_124_3477_n1431), .S(DP_OP_422J2_124_3477_n1432) );
  FADDX1_HVT DP_OP_422J2_124_3477_U812 ( .A(DP_OP_422J2_124_3477_n1438), .B(
        DP_OP_422J2_124_3477_n1583), .CI(DP_OP_422J2_124_3477_n1436), .CO(
        DP_OP_422J2_124_3477_n1429), .S(DP_OP_422J2_124_3477_n1430) );
  FADDX1_HVT DP_OP_422J2_124_3477_U811 ( .A(DP_OP_422J2_124_3477_n1581), .B(
        DP_OP_422J2_124_3477_n1434), .CI(DP_OP_422J2_124_3477_n1432), .CO(
        DP_OP_422J2_124_3477_n1427), .S(DP_OP_422J2_124_3477_n1428) );
  FADDX1_HVT DP_OP_422J2_124_3477_U810 ( .A(DP_OP_422J2_124_3477_n1579), .B(
        DP_OP_422J2_124_3477_n1828), .CI(DP_OP_422J2_124_3477_n2749), .CO(
        DP_OP_422J2_124_3477_n1425), .S(DP_OP_422J2_124_3477_n1426) );
  FADDX1_HVT DP_OP_422J2_124_3477_U809 ( .A(DP_OP_422J2_124_3477_n2004), .B(
        DP_OP_422J2_124_3477_n2443), .CI(DP_OP_422J2_124_3477_n1960), .CO(
        DP_OP_422J2_124_3477_n1423), .S(DP_OP_422J2_124_3477_n1424) );
  FADDX1_HVT DP_OP_422J2_124_3477_U808 ( .A(DP_OP_422J2_124_3477_n2705), .B(
        DP_OP_422J2_124_3477_n2575), .CI(DP_OP_422J2_124_3477_n2531), .CO(
        DP_OP_422J2_124_3477_n1421), .S(DP_OP_422J2_124_3477_n1422) );
  FADDX1_HVT DP_OP_422J2_124_3477_U807 ( .A(DP_OP_422J2_124_3477_n2619), .B(
        DP_OP_422J2_124_3477_n2179), .CI(DP_OP_422J2_124_3477_n1916), .CO(
        DP_OP_422J2_124_3477_n1419), .S(DP_OP_422J2_124_3477_n1420) );
  FADDX1_HVT DP_OP_422J2_124_3477_U806 ( .A(DP_OP_422J2_124_3477_n2091), .B(
        DP_OP_422J2_124_3477_n2487), .CI(DP_OP_422J2_124_3477_n2047), .CO(
        DP_OP_422J2_124_3477_n1417), .S(DP_OP_422J2_124_3477_n1418) );
  FADDX1_HVT DP_OP_422J2_124_3477_U805 ( .A(DP_OP_422J2_124_3477_n2311), .B(
        DP_OP_422J2_124_3477_n2267), .CI(DP_OP_422J2_124_3477_n2881), .CO(
        DP_OP_422J2_124_3477_n1415), .S(DP_OP_422J2_124_3477_n1416) );
  FADDX1_HVT DP_OP_422J2_124_3477_U804 ( .A(DP_OP_422J2_124_3477_n2837), .B(
        DP_OP_422J2_124_3477_n2355), .CI(DP_OP_422J2_124_3477_n2135), .CO(
        DP_OP_422J2_124_3477_n1413), .S(DP_OP_422J2_124_3477_n1414) );
  FADDX1_HVT DP_OP_422J2_124_3477_U803 ( .A(DP_OP_422J2_124_3477_n1872), .B(
        DP_OP_422J2_124_3477_n2793), .CI(DP_OP_422J2_124_3477_n2663), .CO(
        DP_OP_422J2_124_3477_n1411), .S(DP_OP_422J2_124_3477_n1412) );
  FADDX1_HVT DP_OP_422J2_124_3477_U802 ( .A(DP_OP_422J2_124_3477_n2399), .B(
        DP_OP_422J2_124_3477_n1967), .CI(DP_OP_422J2_124_3477_n2582), .CO(
        DP_OP_422J2_124_3477_n1409), .S(DP_OP_422J2_124_3477_n1410) );
  FADDX1_HVT DP_OP_422J2_124_3477_U801 ( .A(DP_OP_422J2_124_3477_n2596), .B(
        DP_OP_422J2_124_3477_n2726), .CI(DP_OP_422J2_124_3477_n2274), .CO(
        DP_OP_422J2_124_3477_n1407), .S(DP_OP_422J2_124_3477_n1408) );
  FADDX1_HVT DP_OP_422J2_124_3477_U800 ( .A(DP_OP_422J2_124_3477_n2420), .B(
        DP_OP_422J2_124_3477_n2413), .CI(DP_OP_422J2_124_3477_n2068), .CO(
        DP_OP_422J2_124_3477_n1405), .S(DP_OP_422J2_124_3477_n1406) );
  FADDX1_HVT DP_OP_422J2_124_3477_U799 ( .A(DP_OP_422J2_124_3477_n2200), .B(
        DP_OP_422J2_124_3477_n2538), .CI(DP_OP_422J2_124_3477_n2142), .CO(
        DP_OP_422J2_124_3477_n1403), .S(DP_OP_422J2_124_3477_n1404) );
  FADDX1_HVT DP_OP_422J2_124_3477_U798 ( .A(DP_OP_422J2_124_3477_n2552), .B(
        DP_OP_422J2_124_3477_n2149), .CI(DP_OP_422J2_124_3477_n2288), .CO(
        DP_OP_422J2_124_3477_n1401), .S(DP_OP_422J2_124_3477_n1402) );
  FADDX1_HVT DP_OP_422J2_124_3477_U797 ( .A(DP_OP_422J2_124_3477_n2888), .B(
        DP_OP_422J2_124_3477_n2223), .CI(DP_OP_422J2_124_3477_n2508), .CO(
        DP_OP_422J2_124_3477_n1399), .S(DP_OP_422J2_124_3477_n1400) );
  FADDX1_HVT DP_OP_422J2_124_3477_U796 ( .A(DP_OP_422J2_124_3477_n2640), .B(
        DP_OP_422J2_124_3477_n1784), .CI(DP_OP_422J2_124_3477_n2858), .CO(
        DP_OP_422J2_124_3477_n1397), .S(DP_OP_422J2_124_3477_n1398) );
  FADDX1_HVT DP_OP_422J2_124_3477_U795 ( .A(DP_OP_422J2_124_3477_n2332), .B(
        DP_OP_422J2_124_3477_n2061), .CI(DP_OP_422J2_124_3477_n2098), .CO(
        DP_OP_422J2_124_3477_n1395), .S(DP_OP_422J2_124_3477_n1396) );
  FADDX1_HVT DP_OP_422J2_124_3477_U794 ( .A(DP_OP_422J2_124_3477_n2464), .B(
        DP_OP_422J2_124_3477_n1842), .CI(DP_OP_422J2_124_3477_n1893), .CO(
        DP_OP_422J2_124_3477_n1393), .S(DP_OP_422J2_124_3477_n1394) );
  FADDX1_HVT DP_OP_422J2_124_3477_U793 ( .A(DP_OP_422J2_124_3477_n2112), .B(
        DP_OP_422J2_124_3477_n1981), .CI(DP_OP_422J2_124_3477_n2770), .CO(
        DP_OP_422J2_124_3477_n1391), .S(DP_OP_422J2_124_3477_n1392) );
  FADDX1_HVT DP_OP_422J2_124_3477_U792 ( .A(DP_OP_422J2_124_3477_n1849), .B(
        DP_OP_422J2_124_3477_n2325), .CI(DP_OP_422J2_124_3477_n2230), .CO(
        DP_OP_422J2_124_3477_n1389), .S(DP_OP_422J2_124_3477_n1390) );
  FADDX1_HVT DP_OP_422J2_124_3477_U791 ( .A(DP_OP_422J2_124_3477_n2844), .B(
        DP_OP_422J2_124_3477_n2633), .CI(DP_OP_422J2_124_3477_n2450), .CO(
        DP_OP_422J2_124_3477_n1387), .S(DP_OP_422J2_124_3477_n1388) );
  FADDX1_HVT DP_OP_422J2_124_3477_U790 ( .A(DP_OP_422J2_124_3477_n2589), .B(
        DP_OP_422J2_124_3477_n2756), .CI(DP_OP_422J2_124_3477_n2684), .CO(
        DP_OP_422J2_124_3477_n1385), .S(DP_OP_422J2_124_3477_n1386) );
  FADDX1_HVT DP_OP_422J2_124_3477_U789 ( .A(DP_OP_422J2_124_3477_n2501), .B(
        DP_OP_422J2_124_3477_n2024), .CI(DP_OP_422J2_124_3477_n1886), .CO(
        DP_OP_422J2_124_3477_n1383), .S(DP_OP_422J2_124_3477_n1384) );
  FADDX1_HVT DP_OP_422J2_124_3477_U788 ( .A(DP_OP_422J2_124_3477_n2494), .B(
        DP_OP_422J2_124_3477_n2054), .CI(DP_OP_422J2_124_3477_n2186), .CO(
        DP_OP_422J2_124_3477_n1381), .S(DP_OP_422J2_124_3477_n1382) );
  FADDX1_HVT DP_OP_422J2_124_3477_U787 ( .A(DP_OP_422J2_124_3477_n2105), .B(
        DP_OP_422J2_124_3477_n2318), .CI(DP_OP_422J2_124_3477_n1923), .CO(
        DP_OP_422J2_124_3477_n1379), .S(DP_OP_422J2_124_3477_n1380) );
  FADDX1_HVT DP_OP_422J2_124_3477_U786 ( .A(DP_OP_422J2_124_3477_n2362), .B(
        DP_OP_422J2_124_3477_n2670), .CI(DP_OP_422J2_124_3477_n1835), .CO(
        DP_OP_422J2_124_3477_n1377), .S(DP_OP_422J2_124_3477_n1378) );
  FADDX1_HVT DP_OP_422J2_124_3477_U785 ( .A(DP_OP_422J2_124_3477_n2677), .B(
        DP_OP_422J2_124_3477_n2851), .CI(DP_OP_422J2_124_3477_n2237), .CO(
        DP_OP_422J2_124_3477_n1375), .S(DP_OP_422J2_124_3477_n1376) );
  FADDX1_HVT DP_OP_422J2_124_3477_U784 ( .A(DP_OP_422J2_124_3477_n2244), .B(
        DP_OP_422J2_124_3477_n2895), .CI(DP_OP_422J2_124_3477_n2193), .CO(
        DP_OP_422J2_124_3477_n1373), .S(DP_OP_422J2_124_3477_n1374) );
  FADDX1_HVT DP_OP_422J2_124_3477_U783 ( .A(DP_OP_422J2_124_3477_n2457), .B(
        DP_OP_422J2_124_3477_n2281), .CI(DP_OP_422J2_124_3477_n2369), .CO(
        DP_OP_422J2_124_3477_n1371), .S(DP_OP_422J2_124_3477_n1372) );
  FADDX1_HVT DP_OP_422J2_124_3477_U782 ( .A(DP_OP_422J2_124_3477_n2712), .B(
        DP_OP_422J2_124_3477_n2763), .CI(DP_OP_422J2_124_3477_n2010), .CO(
        DP_OP_422J2_124_3477_n1369), .S(DP_OP_422J2_124_3477_n1370) );
  FADDX1_HVT DP_OP_422J2_124_3477_U781 ( .A(DP_OP_422J2_124_3477_n2545), .B(
        DP_OP_422J2_124_3477_n2807), .CI(DP_OP_422J2_124_3477_n1974), .CO(
        DP_OP_422J2_124_3477_n1367), .S(DP_OP_422J2_124_3477_n1368) );
  FADDX1_HVT DP_OP_422J2_124_3477_U780 ( .A(DP_OP_422J2_124_3477_n1937), .B(
        DP_OP_422J2_124_3477_n2406), .CI(DP_OP_422J2_124_3477_n2626), .CO(
        DP_OP_422J2_124_3477_n1365), .S(DP_OP_422J2_124_3477_n1366) );
  FADDX1_HVT DP_OP_422J2_124_3477_U779 ( .A(DP_OP_422J2_124_3477_n2156), .B(
        DP_OP_422J2_124_3477_n2800), .CI(DP_OP_422J2_124_3477_n2814), .CO(
        DP_OP_422J2_124_3477_n1363), .S(DP_OP_422J2_124_3477_n1364) );
  FADDX1_HVT DP_OP_422J2_124_3477_U778 ( .A(DP_OP_422J2_124_3477_n2017), .B(
        DP_OP_422J2_124_3477_n2902), .CI(DP_OP_422J2_124_3477_n2376), .CO(
        DP_OP_422J2_124_3477_n1361), .S(DP_OP_422J2_124_3477_n1362) );
  FADDX1_HVT DP_OP_422J2_124_3477_U777 ( .A(DP_OP_422J2_124_3477_n1930), .B(
        DP_OP_422J2_124_3477_n1879), .CI(DP_OP_422J2_124_3477_n2719), .CO(
        DP_OP_422J2_124_3477_n1359), .S(DP_OP_422J2_124_3477_n1360) );
  FADDX1_HVT DP_OP_422J2_124_3477_U776 ( .A(DP_OP_422J2_124_3477_n1577), .B(
        DP_OP_422J2_124_3477_n1565), .CI(DP_OP_422J2_124_3477_n1563), .CO(
        DP_OP_422J2_124_3477_n1357), .S(DP_OP_422J2_124_3477_n1358) );
  FADDX1_HVT DP_OP_422J2_124_3477_U775 ( .A(DP_OP_422J2_124_3477_n1575), .B(
        DP_OP_422J2_124_3477_n1567), .CI(DP_OP_422J2_124_3477_n1569), .CO(
        DP_OP_422J2_124_3477_n1355), .S(DP_OP_422J2_124_3477_n1356) );
  FADDX1_HVT DP_OP_422J2_124_3477_U774 ( .A(DP_OP_422J2_124_3477_n1573), .B(
        DP_OP_422J2_124_3477_n1571), .CI(DP_OP_422J2_124_3477_n1561), .CO(
        DP_OP_422J2_124_3477_n1353), .S(DP_OP_422J2_124_3477_n1354) );
  FADDX1_HVT DP_OP_422J2_124_3477_U773 ( .A(DP_OP_422J2_124_3477_n1559), .B(
        DP_OP_422J2_124_3477_n1537), .CI(DP_OP_422J2_124_3477_n1535), .CO(
        DP_OP_422J2_124_3477_n1351), .S(DP_OP_422J2_124_3477_n1352) );
  FADDX1_HVT DP_OP_422J2_124_3477_U772 ( .A(DP_OP_422J2_124_3477_n1557), .B(
        DP_OP_422J2_124_3477_n1539), .CI(DP_OP_422J2_124_3477_n1541), .CO(
        DP_OP_422J2_124_3477_n1349), .S(DP_OP_422J2_124_3477_n1350) );
  FADDX1_HVT DP_OP_422J2_124_3477_U771 ( .A(DP_OP_422J2_124_3477_n1555), .B(
        DP_OP_422J2_124_3477_n1543), .CI(DP_OP_422J2_124_3477_n1545), .CO(
        DP_OP_422J2_124_3477_n1347), .S(DP_OP_422J2_124_3477_n1348) );
  FADDX1_HVT DP_OP_422J2_124_3477_U770 ( .A(DP_OP_422J2_124_3477_n1553), .B(
        DP_OP_422J2_124_3477_n1547), .CI(DP_OP_422J2_124_3477_n1549), .CO(
        DP_OP_422J2_124_3477_n1345), .S(DP_OP_422J2_124_3477_n1346) );
  FADDX1_HVT DP_OP_422J2_124_3477_U769 ( .A(DP_OP_422J2_124_3477_n1551), .B(
        DP_OP_422J2_124_3477_n1533), .CI(DP_OP_422J2_124_3477_n1531), .CO(
        DP_OP_422J2_124_3477_n1343), .S(DP_OP_422J2_124_3477_n1344) );
  FADDX1_HVT DP_OP_422J2_124_3477_U768 ( .A(DP_OP_422J2_124_3477_n1529), .B(
        DP_OP_422J2_124_3477_n1420), .CI(DP_OP_422J2_124_3477_n1515), .CO(
        DP_OP_422J2_124_3477_n1341), .S(DP_OP_422J2_124_3477_n1342) );
  FADDX1_HVT DP_OP_422J2_124_3477_U767 ( .A(DP_OP_422J2_124_3477_n1527), .B(
        DP_OP_422J2_124_3477_n1412), .CI(DP_OP_422J2_124_3477_n1513), .CO(
        DP_OP_422J2_124_3477_n1339), .S(DP_OP_422J2_124_3477_n1340) );
  FADDX1_HVT DP_OP_422J2_124_3477_U766 ( .A(DP_OP_422J2_124_3477_n1525), .B(
        DP_OP_422J2_124_3477_n1414), .CI(DP_OP_422J2_124_3477_n1517), .CO(
        DP_OP_422J2_124_3477_n1337), .S(DP_OP_422J2_124_3477_n1338) );
  FADDX1_HVT DP_OP_422J2_124_3477_U765 ( .A(DP_OP_422J2_124_3477_n1523), .B(
        DP_OP_422J2_124_3477_n1416), .CI(DP_OP_422J2_124_3477_n1418), .CO(
        DP_OP_422J2_124_3477_n1335), .S(DP_OP_422J2_124_3477_n1336) );
  FADDX1_HVT DP_OP_422J2_124_3477_U764 ( .A(DP_OP_422J2_124_3477_n1521), .B(
        DP_OP_422J2_124_3477_n1424), .CI(DP_OP_422J2_124_3477_n1426), .CO(
        DP_OP_422J2_124_3477_n1333), .S(DP_OP_422J2_124_3477_n1334) );
  FADDX1_HVT DP_OP_422J2_124_3477_U763 ( .A(DP_OP_422J2_124_3477_n1519), .B(
        DP_OP_422J2_124_3477_n1422), .CI(DP_OP_422J2_124_3477_n1511), .CO(
        DP_OP_422J2_124_3477_n1331), .S(DP_OP_422J2_124_3477_n1332) );
  FADDX1_HVT DP_OP_422J2_124_3477_U762 ( .A(DP_OP_422J2_124_3477_n1410), .B(
        DP_OP_422J2_124_3477_n1386), .CI(DP_OP_422J2_124_3477_n1384), .CO(
        DP_OP_422J2_124_3477_n1329), .S(DP_OP_422J2_124_3477_n1330) );
  FADDX1_HVT DP_OP_422J2_124_3477_U761 ( .A(DP_OP_422J2_124_3477_n1400), .B(
        DP_OP_422J2_124_3477_n1398), .CI(DP_OP_422J2_124_3477_n1394), .CO(
        DP_OP_422J2_124_3477_n1327), .S(DP_OP_422J2_124_3477_n1328) );
  FADDX1_HVT DP_OP_422J2_124_3477_U760 ( .A(DP_OP_422J2_124_3477_n1396), .B(
        DP_OP_422J2_124_3477_n1388), .CI(DP_OP_422J2_124_3477_n1390), .CO(
        DP_OP_422J2_124_3477_n1325), .S(DP_OP_422J2_124_3477_n1326) );
  FADDX1_HVT DP_OP_422J2_124_3477_U759 ( .A(DP_OP_422J2_124_3477_n1402), .B(
        DP_OP_422J2_124_3477_n1408), .CI(DP_OP_422J2_124_3477_n1404), .CO(
        DP_OP_422J2_124_3477_n1323), .S(DP_OP_422J2_124_3477_n1324) );
  FADDX1_HVT DP_OP_422J2_124_3477_U758 ( .A(DP_OP_422J2_124_3477_n1406), .B(
        DP_OP_422J2_124_3477_n1392), .CI(DP_OP_422J2_124_3477_n1382), .CO(
        DP_OP_422J2_124_3477_n1321), .S(DP_OP_422J2_124_3477_n1322) );
  FADDX1_HVT DP_OP_422J2_124_3477_U757 ( .A(DP_OP_422J2_124_3477_n1380), .B(
        DP_OP_422J2_124_3477_n1366), .CI(DP_OP_422J2_124_3477_n1360), .CO(
        DP_OP_422J2_124_3477_n1319), .S(DP_OP_422J2_124_3477_n1320) );
  FADDX1_HVT DP_OP_422J2_124_3477_U756 ( .A(DP_OP_422J2_124_3477_n1378), .B(
        DP_OP_422J2_124_3477_n1370), .CI(DP_OP_422J2_124_3477_n1364), .CO(
        DP_OP_422J2_124_3477_n1317), .S(DP_OP_422J2_124_3477_n1318) );
  FADDX1_HVT DP_OP_422J2_124_3477_U755 ( .A(DP_OP_422J2_124_3477_n1376), .B(
        DP_OP_422J2_124_3477_n1368), .CI(DP_OP_422J2_124_3477_n1362), .CO(
        DP_OP_422J2_124_3477_n1315), .S(DP_OP_422J2_124_3477_n1316) );
  FADDX1_HVT DP_OP_422J2_124_3477_U754 ( .A(DP_OP_422J2_124_3477_n1374), .B(
        DP_OP_422J2_124_3477_n1372), .CI(DP_OP_422J2_124_3477_n1509), .CO(
        DP_OP_422J2_124_3477_n1313), .S(DP_OP_422J2_124_3477_n1314) );
  FADDX1_HVT DP_OP_422J2_124_3477_U753 ( .A(DP_OP_422J2_124_3477_n1507), .B(
        DP_OP_422J2_124_3477_n1505), .CI(DP_OP_422J2_124_3477_n1501), .CO(
        DP_OP_422J2_124_3477_n1311), .S(DP_OP_422J2_124_3477_n1312) );
  FADDX1_HVT DP_OP_422J2_124_3477_U752 ( .A(DP_OP_422J2_124_3477_n1503), .B(
        DP_OP_422J2_124_3477_n1499), .CI(DP_OP_422J2_124_3477_n1497), .CO(
        DP_OP_422J2_124_3477_n1309), .S(DP_OP_422J2_124_3477_n1310) );
  FADDX1_HVT DP_OP_422J2_124_3477_U751 ( .A(DP_OP_422J2_124_3477_n1495), .B(
        DP_OP_422J2_124_3477_n1356), .CI(DP_OP_422J2_124_3477_n1354), .CO(
        DP_OP_422J2_124_3477_n1307), .S(DP_OP_422J2_124_3477_n1308) );
  FADDX1_HVT DP_OP_422J2_124_3477_U750 ( .A(DP_OP_422J2_124_3477_n1493), .B(
        DP_OP_422J2_124_3477_n1489), .CI(DP_OP_422J2_124_3477_n1358), .CO(
        DP_OP_422J2_124_3477_n1305), .S(DP_OP_422J2_124_3477_n1306) );
  FADDX1_HVT DP_OP_422J2_124_3477_U749 ( .A(DP_OP_422J2_124_3477_n1491), .B(
        DP_OP_422J2_124_3477_n1487), .CI(DP_OP_422J2_124_3477_n1485), .CO(
        DP_OP_422J2_124_3477_n1303), .S(DP_OP_422J2_124_3477_n1304) );
  FADDX1_HVT DP_OP_422J2_124_3477_U748 ( .A(DP_OP_422J2_124_3477_n1483), .B(
        DP_OP_422J2_124_3477_n1350), .CI(DP_OP_422J2_124_3477_n1344), .CO(
        DP_OP_422J2_124_3477_n1301), .S(DP_OP_422J2_124_3477_n1302) );
  FADDX1_HVT DP_OP_422J2_124_3477_U747 ( .A(DP_OP_422J2_124_3477_n1481), .B(
        DP_OP_422J2_124_3477_n1352), .CI(DP_OP_422J2_124_3477_n1348), .CO(
        DP_OP_422J2_124_3477_n1299), .S(DP_OP_422J2_124_3477_n1300) );
  FADDX1_HVT DP_OP_422J2_124_3477_U746 ( .A(DP_OP_422J2_124_3477_n1479), .B(
        DP_OP_422J2_124_3477_n1346), .CI(DP_OP_422J2_124_3477_n1477), .CO(
        DP_OP_422J2_124_3477_n1297), .S(DP_OP_422J2_124_3477_n1298) );
  FADDX1_HVT DP_OP_422J2_124_3477_U745 ( .A(DP_OP_422J2_124_3477_n1475), .B(
        DP_OP_422J2_124_3477_n1332), .CI(DP_OP_422J2_124_3477_n1471), .CO(
        DP_OP_422J2_124_3477_n1295), .S(DP_OP_422J2_124_3477_n1296) );
  FADDX1_HVT DP_OP_422J2_124_3477_U744 ( .A(DP_OP_422J2_124_3477_n1342), .B(
        DP_OP_422J2_124_3477_n1336), .CI(DP_OP_422J2_124_3477_n1334), .CO(
        DP_OP_422J2_124_3477_n1293), .S(DP_OP_422J2_124_3477_n1294) );
  FADDX1_HVT DP_OP_422J2_124_3477_U743 ( .A(DP_OP_422J2_124_3477_n1473), .B(
        DP_OP_422J2_124_3477_n1340), .CI(DP_OP_422J2_124_3477_n1338), .CO(
        DP_OP_422J2_124_3477_n1291), .S(DP_OP_422J2_124_3477_n1292) );
  FADDX1_HVT DP_OP_422J2_124_3477_U742 ( .A(DP_OP_422J2_124_3477_n1330), .B(
        DP_OP_422J2_124_3477_n1324), .CI(DP_OP_422J2_124_3477_n1322), .CO(
        DP_OP_422J2_124_3477_n1289), .S(DP_OP_422J2_124_3477_n1290) );
  FADDX1_HVT DP_OP_422J2_124_3477_U741 ( .A(DP_OP_422J2_124_3477_n1326), .B(
        DP_OP_422J2_124_3477_n1328), .CI(DP_OP_422J2_124_3477_n1320), .CO(
        DP_OP_422J2_124_3477_n1287), .S(DP_OP_422J2_124_3477_n1288) );
  FADDX1_HVT DP_OP_422J2_124_3477_U740 ( .A(DP_OP_422J2_124_3477_n1318), .B(
        DP_OP_422J2_124_3477_n1316), .CI(DP_OP_422J2_124_3477_n1469), .CO(
        DP_OP_422J2_124_3477_n1285), .S(DP_OP_422J2_124_3477_n1286) );
  FADDX1_HVT DP_OP_422J2_124_3477_U739 ( .A(DP_OP_422J2_124_3477_n1467), .B(
        DP_OP_422J2_124_3477_n1314), .CI(DP_OP_422J2_124_3477_n1465), .CO(
        DP_OP_422J2_124_3477_n1283), .S(DP_OP_422J2_124_3477_n1284) );
  FADDX1_HVT DP_OP_422J2_124_3477_U738 ( .A(DP_OP_422J2_124_3477_n1463), .B(
        DP_OP_422J2_124_3477_n1312), .CI(DP_OP_422J2_124_3477_n1310), .CO(
        DP_OP_422J2_124_3477_n1281), .S(DP_OP_422J2_124_3477_n1282) );
  FADDX1_HVT DP_OP_422J2_124_3477_U737 ( .A(DP_OP_422J2_124_3477_n1461), .B(
        DP_OP_422J2_124_3477_n1459), .CI(DP_OP_422J2_124_3477_n1457), .CO(
        DP_OP_422J2_124_3477_n1279), .S(DP_OP_422J2_124_3477_n1280) );
  FADDX1_HVT DP_OP_422J2_124_3477_U736 ( .A(DP_OP_422J2_124_3477_n1455), .B(
        DP_OP_422J2_124_3477_n1308), .CI(DP_OP_422J2_124_3477_n1306), .CO(
        DP_OP_422J2_124_3477_n1277), .S(DP_OP_422J2_124_3477_n1278) );
  FADDX1_HVT DP_OP_422J2_124_3477_U735 ( .A(DP_OP_422J2_124_3477_n1304), .B(
        DP_OP_422J2_124_3477_n1300), .CI(DP_OP_422J2_124_3477_n1298), .CO(
        DP_OP_422J2_124_3477_n1275), .S(DP_OP_422J2_124_3477_n1276) );
  FADDX1_HVT DP_OP_422J2_124_3477_U734 ( .A(DP_OP_422J2_124_3477_n1453), .B(
        DP_OP_422J2_124_3477_n1302), .CI(DP_OP_422J2_124_3477_n1451), .CO(
        DP_OP_422J2_124_3477_n1273), .S(DP_OP_422J2_124_3477_n1274) );
  FADDX1_HVT DP_OP_422J2_124_3477_U733 ( .A(DP_OP_422J2_124_3477_n1449), .B(
        DP_OP_422J2_124_3477_n1296), .CI(DP_OP_422J2_124_3477_n1292), .CO(
        DP_OP_422J2_124_3477_n1271), .S(DP_OP_422J2_124_3477_n1272) );
  FADDX1_HVT DP_OP_422J2_124_3477_U732 ( .A(DP_OP_422J2_124_3477_n1294), .B(
        DP_OP_422J2_124_3477_n1290), .CI(DP_OP_422J2_124_3477_n1447), .CO(
        DP_OP_422J2_124_3477_n1269), .S(DP_OP_422J2_124_3477_n1270) );
  FADDX1_HVT DP_OP_422J2_124_3477_U731 ( .A(DP_OP_422J2_124_3477_n1288), .B(
        DP_OP_422J2_124_3477_n1286), .CI(DP_OP_422J2_124_3477_n1445), .CO(
        DP_OP_422J2_124_3477_n1267), .S(DP_OP_422J2_124_3477_n1268) );
  FADDX1_HVT DP_OP_422J2_124_3477_U730 ( .A(DP_OP_422J2_124_3477_n1284), .B(
        DP_OP_422J2_124_3477_n1443), .CI(DP_OP_422J2_124_3477_n1441), .CO(
        DP_OP_422J2_124_3477_n1265), .S(DP_OP_422J2_124_3477_n1266) );
  FADDX1_HVT DP_OP_422J2_124_3477_U729 ( .A(DP_OP_422J2_124_3477_n1282), .B(
        DP_OP_422J2_124_3477_n1280), .CI(DP_OP_422J2_124_3477_n1439), .CO(
        DP_OP_422J2_124_3477_n1263), .S(DP_OP_422J2_124_3477_n1264) );
  FADDX1_HVT DP_OP_422J2_124_3477_U728 ( .A(DP_OP_422J2_124_3477_n1278), .B(
        DP_OP_422J2_124_3477_n1437), .CI(DP_OP_422J2_124_3477_n1276), .CO(
        DP_OP_422J2_124_3477_n1261), .S(DP_OP_422J2_124_3477_n1262) );
  FADDX1_HVT DP_OP_422J2_124_3477_U727 ( .A(DP_OP_422J2_124_3477_n1274), .B(
        DP_OP_422J2_124_3477_n1272), .CI(DP_OP_422J2_124_3477_n1435), .CO(
        DP_OP_422J2_124_3477_n1259), .S(DP_OP_422J2_124_3477_n1260) );
  FADDX1_HVT DP_OP_422J2_124_3477_U726 ( .A(DP_OP_422J2_124_3477_n1270), .B(
        DP_OP_422J2_124_3477_n1268), .CI(DP_OP_422J2_124_3477_n1433), .CO(
        DP_OP_422J2_124_3477_n1257), .S(DP_OP_422J2_124_3477_n1258) );
  FADDX1_HVT DP_OP_422J2_124_3477_U725 ( .A(DP_OP_422J2_124_3477_n1266), .B(
        DP_OP_422J2_124_3477_n1431), .CI(DP_OP_422J2_124_3477_n1264), .CO(
        DP_OP_422J2_124_3477_n1255), .S(DP_OP_422J2_124_3477_n1256) );
  FADDX1_HVT DP_OP_422J2_124_3477_U724 ( .A(DP_OP_422J2_124_3477_n1262), .B(
        DP_OP_422J2_124_3477_n1429), .CI(DP_OP_422J2_124_3477_n1260), .CO(
        DP_OP_422J2_124_3477_n1253), .S(DP_OP_422J2_124_3477_n1254) );
  FADDX1_HVT DP_OP_422J2_124_3477_U723 ( .A(DP_OP_422J2_124_3477_n1258), .B(
        DP_OP_422J2_124_3477_n1427), .CI(DP_OP_422J2_124_3477_n1256), .CO(
        DP_OP_422J2_124_3477_n1251), .S(DP_OP_422J2_124_3477_n1252) );
  HADDX1_HVT DP_OP_422J2_124_3477_U722 ( .A0(DP_OP_422J2_124_3477_n2704), .B0(
        DP_OP_422J2_124_3477_n1827), .C1(DP_OP_422J2_124_3477_n1249), .SO(
        DP_OP_422J2_124_3477_n1250) );
  FADDX1_HVT DP_OP_422J2_124_3477_U721 ( .A(DP_OP_422J2_124_3477_n2003), .B(
        DP_OP_422J2_124_3477_n2530), .CI(DP_OP_422J2_124_3477_n1959), .CO(
        DP_OP_422J2_124_3477_n1247), .S(DP_OP_422J2_124_3477_n1248) );
  FADDX1_HVT DP_OP_422J2_124_3477_U720 ( .A(DP_OP_422J2_124_3477_n2310), .B(
        DP_OP_422J2_124_3477_n2046), .CI(DP_OP_422J2_124_3477_n2748), .CO(
        DP_OP_422J2_124_3477_n1245), .S(DP_OP_422J2_124_3477_n1246) );
  FADDX1_HVT DP_OP_422J2_124_3477_U719 ( .A(DP_OP_422J2_124_3477_n2662), .B(
        DP_OP_422J2_124_3477_n2442), .CI(DP_OP_422J2_124_3477_n2178), .CO(
        DP_OP_422J2_124_3477_n1243), .S(DP_OP_422J2_124_3477_n1244) );
  FADDX1_HVT DP_OP_422J2_124_3477_U718 ( .A(DP_OP_422J2_124_3477_n1871), .B(
        DP_OP_422J2_124_3477_n1915), .CI(DP_OP_422J2_124_3477_n2574), .CO(
        DP_OP_422J2_124_3477_n1241), .S(DP_OP_422J2_124_3477_n1242) );
  FADDX1_HVT DP_OP_422J2_124_3477_U717 ( .A(DP_OP_422J2_124_3477_n2354), .B(
        DP_OP_422J2_124_3477_n2880), .CI(DP_OP_422J2_124_3477_n2486), .CO(
        DP_OP_422J2_124_3477_n1239), .S(DP_OP_422J2_124_3477_n1240) );
  FADDX1_HVT DP_OP_422J2_124_3477_U716 ( .A(DP_OP_422J2_124_3477_n2090), .B(
        DP_OP_422J2_124_3477_n2836), .CI(DP_OP_422J2_124_3477_n2266), .CO(
        DP_OP_422J2_124_3477_n1237), .S(DP_OP_422J2_124_3477_n1238) );
  FADDX1_HVT DP_OP_422J2_124_3477_U715 ( .A(DP_OP_422J2_124_3477_n2792), .B(
        DP_OP_422J2_124_3477_n2134), .CI(DP_OP_422J2_124_3477_n2618), .CO(
        DP_OP_422J2_124_3477_n1235), .S(DP_OP_422J2_124_3477_n1236) );
  FADDX1_HVT DP_OP_422J2_124_3477_U714 ( .A(DP_OP_422J2_124_3477_n2398), .B(
        DP_OP_422J2_124_3477_n1966), .CI(DP_OP_422J2_124_3477_n2581), .CO(
        DP_OP_422J2_124_3477_n1233), .S(DP_OP_422J2_124_3477_n1234) );
  FADDX1_HVT DP_OP_422J2_124_3477_U713 ( .A(DP_OP_422J2_124_3477_n2639), .B(
        DP_OP_422J2_124_3477_n2148), .CI(DP_OP_422J2_124_3477_n2067), .CO(
        DP_OP_422J2_124_3477_n1231), .S(DP_OP_422J2_124_3477_n1232) );
  FADDX1_HVT DP_OP_422J2_124_3477_U712 ( .A(DP_OP_422J2_124_3477_n2419), .B(
        DP_OP_422J2_124_3477_n2537), .CI(DP_OP_422J2_124_3477_n2141), .CO(
        DP_OP_422J2_124_3477_n1229), .S(DP_OP_422J2_124_3477_n1230) );
  FADDX1_HVT DP_OP_422J2_124_3477_U711 ( .A(DP_OP_422J2_124_3477_n1848), .B(
        DP_OP_422J2_124_3477_n2412), .CI(DP_OP_422J2_124_3477_n2273), .CO(
        DP_OP_422J2_124_3477_n1227), .S(DP_OP_422J2_124_3477_n1228) );
  FADDX1_HVT DP_OP_422J2_124_3477_U710 ( .A(DP_OP_422J2_124_3477_n2199), .B(
        DP_OP_422J2_124_3477_n2725), .CI(DP_OP_422J2_124_3477_n2287), .CO(
        DP_OP_422J2_124_3477_n1225), .S(DP_OP_422J2_124_3477_n1226) );
  FADDX1_HVT DP_OP_422J2_124_3477_U709 ( .A(DP_OP_422J2_124_3477_n2551), .B(
        DP_OP_422J2_124_3477_n2222), .CI(DP_OP_422J2_124_3477_n2507), .CO(
        DP_OP_422J2_124_3477_n1223), .S(DP_OP_422J2_124_3477_n1224) );
  FADDX1_HVT DP_OP_422J2_124_3477_U708 ( .A(DP_OP_422J2_124_3477_n2595), .B(
        DP_OP_422J2_124_3477_n1783), .CI(DP_OP_422J2_124_3477_n1892), .CO(
        DP_OP_422J2_124_3477_n1221), .S(DP_OP_422J2_124_3477_n1222) );
  FADDX1_HVT DP_OP_422J2_124_3477_U707 ( .A(DP_OP_422J2_124_3477_n2463), .B(
        DP_OP_422J2_124_3477_n2683), .CI(DP_OP_422J2_124_3477_n2769), .CO(
        DP_OP_422J2_124_3477_n1219), .S(DP_OP_422J2_124_3477_n1220) );
  FADDX1_HVT DP_OP_422J2_124_3477_U706 ( .A(DP_OP_422J2_124_3477_n2111), .B(
        DP_OP_422J2_124_3477_n2500), .CI(DP_OP_422J2_124_3477_n2229), .CO(
        DP_OP_422J2_124_3477_n1217), .S(DP_OP_422J2_124_3477_n1218) );
  FADDX1_HVT DP_OP_422J2_124_3477_U705 ( .A(DP_OP_422J2_124_3477_n2887), .B(
        DP_OP_422J2_124_3477_n2755), .CI(DP_OP_422J2_124_3477_n2449), .CO(
        DP_OP_422J2_124_3477_n1215), .S(DP_OP_422J2_124_3477_n1216) );
  FADDX1_HVT DP_OP_422J2_124_3477_U704 ( .A(DP_OP_422J2_124_3477_n2331), .B(
        DP_OP_422J2_124_3477_n1980), .CI(DP_OP_422J2_124_3477_n2097), .CO(
        DP_OP_422J2_124_3477_n1213), .S(DP_OP_422J2_124_3477_n1214) );
  FADDX1_HVT DP_OP_422J2_124_3477_U703 ( .A(DP_OP_422J2_124_3477_n2843), .B(
        DP_OP_422J2_124_3477_n2632), .CI(DP_OP_422J2_124_3477_n2857), .CO(
        DP_OP_422J2_124_3477_n1211), .S(DP_OP_422J2_124_3477_n1212) );
  FADDX1_HVT DP_OP_422J2_124_3477_U702 ( .A(DP_OP_422J2_124_3477_n1841), .B(
        DP_OP_422J2_124_3477_n2324), .CI(DP_OP_422J2_124_3477_n2588), .CO(
        DP_OP_422J2_124_3477_n1209), .S(DP_OP_422J2_124_3477_n1210) );
  FADDX1_HVT DP_OP_422J2_124_3477_U701 ( .A(DP_OP_422J2_124_3477_n2060), .B(
        DP_OP_422J2_124_3477_n2023), .CI(DP_OP_422J2_124_3477_n2104), .CO(
        DP_OP_422J2_124_3477_n1207), .S(DP_OP_422J2_124_3477_n1208) );
  FADDX1_HVT DP_OP_422J2_124_3477_U700 ( .A(DP_OP_422J2_124_3477_n1885), .B(
        DP_OP_422J2_124_3477_n2053), .CI(DP_OP_422J2_124_3477_n1922), .CO(
        DP_OP_422J2_124_3477_n1205), .S(DP_OP_422J2_124_3477_n1206) );
  FADDX1_HVT DP_OP_422J2_124_3477_U699 ( .A(DP_OP_422J2_124_3477_n2493), .B(
        DP_OP_422J2_124_3477_n2317), .CI(DP_OP_422J2_124_3477_n2185), .CO(
        DP_OP_422J2_124_3477_n1203), .S(DP_OP_422J2_124_3477_n1204) );
  FADDX1_HVT DP_OP_422J2_124_3477_U698 ( .A(DP_OP_422J2_124_3477_n2361), .B(
        DP_OP_422J2_124_3477_n2669), .CI(DP_OP_422J2_124_3477_n1834), .CO(
        DP_OP_422J2_124_3477_n1201), .S(DP_OP_422J2_124_3477_n1202) );
  FADDX1_HVT DP_OP_422J2_124_3477_U697 ( .A(DP_OP_422J2_124_3477_n2676), .B(
        DP_OP_422J2_124_3477_n2850), .CI(DP_OP_422J2_124_3477_n2236), .CO(
        DP_OP_422J2_124_3477_n1199), .S(DP_OP_422J2_124_3477_n1200) );
  FADDX1_HVT DP_OP_422J2_124_3477_U696 ( .A(DP_OP_422J2_124_3477_n2243), .B(
        DP_OP_422J2_124_3477_n2894), .CI(DP_OP_422J2_124_3477_n2192), .CO(
        DP_OP_422J2_124_3477_n1197), .S(DP_OP_422J2_124_3477_n1198) );
  FADDX1_HVT DP_OP_422J2_124_3477_U695 ( .A(DP_OP_422J2_124_3477_n2456), .B(
        DP_OP_422J2_124_3477_n2280), .CI(DP_OP_422J2_124_3477_n2368), .CO(
        DP_OP_422J2_124_3477_n1195), .S(DP_OP_422J2_124_3477_n1196) );
  FADDX1_HVT DP_OP_422J2_124_3477_U694 ( .A(DP_OP_422J2_124_3477_n2711), .B(
        DP_OP_422J2_124_3477_n2762), .CI(DP_OP_422J2_124_3477_n2009), .CO(
        DP_OP_422J2_124_3477_n1193), .S(DP_OP_422J2_124_3477_n1194) );
  FADDX1_HVT DP_OP_422J2_124_3477_U693 ( .A(DP_OP_422J2_124_3477_n2544), .B(
        DP_OP_422J2_124_3477_n2806), .CI(DP_OP_422J2_124_3477_n2625), .CO(
        DP_OP_422J2_124_3477_n1191), .S(DP_OP_422J2_124_3477_n1192) );
  FADDX1_HVT DP_OP_422J2_124_3477_U692 ( .A(DP_OP_422J2_124_3477_n1936), .B(
        DP_OP_422J2_124_3477_n2155), .CI(DP_OP_422J2_124_3477_n2799), .CO(
        DP_OP_422J2_124_3477_n1189), .S(DP_OP_422J2_124_3477_n1190) );
  FADDX1_HVT DP_OP_422J2_124_3477_U691 ( .A(DP_OP_422J2_124_3477_n2405), .B(
        DP_OP_422J2_124_3477_n1973), .CI(DP_OP_422J2_124_3477_n2813), .CO(
        DP_OP_422J2_124_3477_n1187), .S(DP_OP_422J2_124_3477_n1188) );
  FADDX1_HVT DP_OP_422J2_124_3477_U690 ( .A(DP_OP_422J2_124_3477_n2016), .B(
        DP_OP_422J2_124_3477_n2375), .CI(DP_OP_422J2_124_3477_n2718), .CO(
        DP_OP_422J2_124_3477_n1185), .S(DP_OP_422J2_124_3477_n1186) );
  FADDX1_HVT DP_OP_422J2_124_3477_U689 ( .A(DP_OP_422J2_124_3477_n1929), .B(
        DP_OP_422J2_124_3477_n1878), .CI(DP_OP_422J2_124_3477_n2901), .CO(
        DP_OP_422J2_124_3477_n1183), .S(DP_OP_422J2_124_3477_n1184) );
  FADDX1_HVT DP_OP_422J2_124_3477_U688 ( .A(DP_OP_422J2_124_3477_n1250), .B(
        DP_OP_422J2_124_3477_n1425), .CI(DP_OP_422J2_124_3477_n1411), .CO(
        DP_OP_422J2_124_3477_n1181), .S(DP_OP_422J2_124_3477_n1182) );
  FADDX1_HVT DP_OP_422J2_124_3477_U687 ( .A(DP_OP_422J2_124_3477_n1423), .B(
        DP_OP_422J2_124_3477_n1413), .CI(DP_OP_422J2_124_3477_n1415), .CO(
        DP_OP_422J2_124_3477_n1179), .S(DP_OP_422J2_124_3477_n1180) );
  FADDX1_HVT DP_OP_422J2_124_3477_U686 ( .A(DP_OP_422J2_124_3477_n1421), .B(
        DP_OP_422J2_124_3477_n1417), .CI(DP_OP_422J2_124_3477_n1419), .CO(
        DP_OP_422J2_124_3477_n1177), .S(DP_OP_422J2_124_3477_n1178) );
  FADDX1_HVT DP_OP_422J2_124_3477_U685 ( .A(DP_OP_422J2_124_3477_n1409), .B(
        DP_OP_422J2_124_3477_n1383), .CI(DP_OP_422J2_124_3477_n1385), .CO(
        DP_OP_422J2_124_3477_n1175), .S(DP_OP_422J2_124_3477_n1176) );
  FADDX1_HVT DP_OP_422J2_124_3477_U684 ( .A(DP_OP_422J2_124_3477_n1407), .B(
        DP_OP_422J2_124_3477_n1387), .CI(DP_OP_422J2_124_3477_n1389), .CO(
        DP_OP_422J2_124_3477_n1173), .S(DP_OP_422J2_124_3477_n1174) );
  FADDX1_HVT DP_OP_422J2_124_3477_U683 ( .A(DP_OP_422J2_124_3477_n1405), .B(
        DP_OP_422J2_124_3477_n1391), .CI(DP_OP_422J2_124_3477_n1393), .CO(
        DP_OP_422J2_124_3477_n1171), .S(DP_OP_422J2_124_3477_n1172) );
  FADDX1_HVT DP_OP_422J2_124_3477_U682 ( .A(DP_OP_422J2_124_3477_n1403), .B(
        DP_OP_422J2_124_3477_n1395), .CI(DP_OP_422J2_124_3477_n1397), .CO(
        DP_OP_422J2_124_3477_n1169), .S(DP_OP_422J2_124_3477_n1170) );
  FADDX1_HVT DP_OP_422J2_124_3477_U681 ( .A(DP_OP_422J2_124_3477_n1401), .B(
        DP_OP_422J2_124_3477_n1399), .CI(DP_OP_422J2_124_3477_n1381), .CO(
        DP_OP_422J2_124_3477_n1167), .S(DP_OP_422J2_124_3477_n1168) );
  FADDX1_HVT DP_OP_422J2_124_3477_U680 ( .A(DP_OP_422J2_124_3477_n1379), .B(
        DP_OP_422J2_124_3477_n1242), .CI(DP_OP_422J2_124_3477_n1359), .CO(
        DP_OP_422J2_124_3477_n1165), .S(DP_OP_422J2_124_3477_n1166) );
  FADDX1_HVT DP_OP_422J2_124_3477_U679 ( .A(DP_OP_422J2_124_3477_n1377), .B(
        DP_OP_422J2_124_3477_n1244), .CI(DP_OP_422J2_124_3477_n1361), .CO(
        DP_OP_422J2_124_3477_n1163), .S(DP_OP_422J2_124_3477_n1164) );
  FADDX1_HVT DP_OP_422J2_124_3477_U678 ( .A(DP_OP_422J2_124_3477_n1375), .B(
        DP_OP_422J2_124_3477_n1246), .CI(DP_OP_422J2_124_3477_n1363), .CO(
        DP_OP_422J2_124_3477_n1161), .S(DP_OP_422J2_124_3477_n1162) );
  FADDX1_HVT DP_OP_422J2_124_3477_U677 ( .A(DP_OP_422J2_124_3477_n1373), .B(
        DP_OP_422J2_124_3477_n1236), .CI(DP_OP_422J2_124_3477_n1238), .CO(
        DP_OP_422J2_124_3477_n1159), .S(DP_OP_422J2_124_3477_n1160) );
  FADDX1_HVT DP_OP_422J2_124_3477_U676 ( .A(DP_OP_422J2_124_3477_n1371), .B(
        DP_OP_422J2_124_3477_n1248), .CI(DP_OP_422J2_124_3477_n1240), .CO(
        DP_OP_422J2_124_3477_n1157), .S(DP_OP_422J2_124_3477_n1158) );
  FADDX1_HVT DP_OP_422J2_124_3477_U675 ( .A(DP_OP_422J2_124_3477_n1367), .B(
        DP_OP_422J2_124_3477_n1369), .CI(DP_OP_422J2_124_3477_n1365), .CO(
        DP_OP_422J2_124_3477_n1155), .S(DP_OP_422J2_124_3477_n1156) );
  FADDX1_HVT DP_OP_422J2_124_3477_U674 ( .A(DP_OP_422J2_124_3477_n1234), .B(
        DP_OP_422J2_124_3477_n1210), .CI(DP_OP_422J2_124_3477_n1208), .CO(
        DP_OP_422J2_124_3477_n1153), .S(DP_OP_422J2_124_3477_n1154) );
  FADDX1_HVT DP_OP_422J2_124_3477_U673 ( .A(DP_OP_422J2_124_3477_n1226), .B(
        DP_OP_422J2_124_3477_n1220), .CI(DP_OP_422J2_124_3477_n1222), .CO(
        DP_OP_422J2_124_3477_n1151), .S(DP_OP_422J2_124_3477_n1152) );
  FADDX1_HVT DP_OP_422J2_124_3477_U672 ( .A(DP_OP_422J2_124_3477_n1224), .B(
        DP_OP_422J2_124_3477_n1214), .CI(DP_OP_422J2_124_3477_n1216), .CO(
        DP_OP_422J2_124_3477_n1149), .S(DP_OP_422J2_124_3477_n1150) );
  FADDX1_HVT DP_OP_422J2_124_3477_U671 ( .A(DP_OP_422J2_124_3477_n1212), .B(
        DP_OP_422J2_124_3477_n1232), .CI(DP_OP_422J2_124_3477_n1228), .CO(
        DP_OP_422J2_124_3477_n1147), .S(DP_OP_422J2_124_3477_n1148) );
  FADDX1_HVT DP_OP_422J2_124_3477_U670 ( .A(DP_OP_422J2_124_3477_n1230), .B(
        DP_OP_422J2_124_3477_n1218), .CI(DP_OP_422J2_124_3477_n1206), .CO(
        DP_OP_422J2_124_3477_n1145), .S(DP_OP_422J2_124_3477_n1146) );
  FADDX1_HVT DP_OP_422J2_124_3477_U669 ( .A(DP_OP_422J2_124_3477_n1204), .B(
        DP_OP_422J2_124_3477_n1190), .CI(DP_OP_422J2_124_3477_n1184), .CO(
        DP_OP_422J2_124_3477_n1143), .S(DP_OP_422J2_124_3477_n1144) );
  FADDX1_HVT DP_OP_422J2_124_3477_U668 ( .A(DP_OP_422J2_124_3477_n1202), .B(
        DP_OP_422J2_124_3477_n1194), .CI(DP_OP_422J2_124_3477_n1188), .CO(
        DP_OP_422J2_124_3477_n1141), .S(DP_OP_422J2_124_3477_n1142) );
  FADDX1_HVT DP_OP_422J2_124_3477_U667 ( .A(DP_OP_422J2_124_3477_n1200), .B(
        DP_OP_422J2_124_3477_n1192), .CI(DP_OP_422J2_124_3477_n1186), .CO(
        DP_OP_422J2_124_3477_n1139), .S(DP_OP_422J2_124_3477_n1140) );
  FADDX1_HVT DP_OP_422J2_124_3477_U666 ( .A(DP_OP_422J2_124_3477_n1198), .B(
        DP_OP_422J2_124_3477_n1196), .CI(DP_OP_422J2_124_3477_n1357), .CO(
        DP_OP_422J2_124_3477_n1137), .S(DP_OP_422J2_124_3477_n1138) );
  FADDX1_HVT DP_OP_422J2_124_3477_U665 ( .A(DP_OP_422J2_124_3477_n1355), .B(
        DP_OP_422J2_124_3477_n1353), .CI(DP_OP_422J2_124_3477_n1351), .CO(
        DP_OP_422J2_124_3477_n1135), .S(DP_OP_422J2_124_3477_n1136) );
  FADDX1_HVT DP_OP_422J2_124_3477_U664 ( .A(DP_OP_422J2_124_3477_n1349), .B(
        DP_OP_422J2_124_3477_n1345), .CI(DP_OP_422J2_124_3477_n1343), .CO(
        DP_OP_422J2_124_3477_n1133), .S(DP_OP_422J2_124_3477_n1134) );
  FADDX1_HVT DP_OP_422J2_124_3477_U663 ( .A(DP_OP_422J2_124_3477_n1347), .B(
        DP_OP_422J2_124_3477_n1182), .CI(DP_OP_422J2_124_3477_n1341), .CO(
        DP_OP_422J2_124_3477_n1131), .S(DP_OP_422J2_124_3477_n1132) );
  FADDX1_HVT DP_OP_422J2_124_3477_U662 ( .A(DP_OP_422J2_124_3477_n1339), .B(
        DP_OP_422J2_124_3477_n1180), .CI(DP_OP_422J2_124_3477_n1178), .CO(
        DP_OP_422J2_124_3477_n1129), .S(DP_OP_422J2_124_3477_n1130) );
  FADDX1_HVT DP_OP_422J2_124_3477_U661 ( .A(DP_OP_422J2_124_3477_n1337), .B(
        DP_OP_422J2_124_3477_n1333), .CI(DP_OP_422J2_124_3477_n1331), .CO(
        DP_OP_422J2_124_3477_n1127), .S(DP_OP_422J2_124_3477_n1128) );
  FADDX1_HVT DP_OP_422J2_124_3477_U660 ( .A(DP_OP_422J2_124_3477_n1335), .B(
        DP_OP_422J2_124_3477_n1329), .CI(DP_OP_422J2_124_3477_n1176), .CO(
        DP_OP_422J2_124_3477_n1125), .S(DP_OP_422J2_124_3477_n1126) );
  FADDX1_HVT DP_OP_422J2_124_3477_U659 ( .A(DP_OP_422J2_124_3477_n1323), .B(
        DP_OP_422J2_124_3477_n1170), .CI(DP_OP_422J2_124_3477_n1168), .CO(
        DP_OP_422J2_124_3477_n1123), .S(DP_OP_422J2_124_3477_n1124) );
  FADDX1_HVT DP_OP_422J2_124_3477_U658 ( .A(DP_OP_422J2_124_3477_n1327), .B(
        DP_OP_422J2_124_3477_n1325), .CI(DP_OP_422J2_124_3477_n1321), .CO(
        DP_OP_422J2_124_3477_n1121), .S(DP_OP_422J2_124_3477_n1122) );
  FADDX1_HVT DP_OP_422J2_124_3477_U657 ( .A(DP_OP_422J2_124_3477_n1174), .B(
        DP_OP_422J2_124_3477_n1172), .CI(DP_OP_422J2_124_3477_n1319), .CO(
        DP_OP_422J2_124_3477_n1119), .S(DP_OP_422J2_124_3477_n1120) );
  FADDX1_HVT DP_OP_422J2_124_3477_U656 ( .A(DP_OP_422J2_124_3477_n1166), .B(
        DP_OP_422J2_124_3477_n1158), .CI(DP_OP_422J2_124_3477_n1156), .CO(
        DP_OP_422J2_124_3477_n1117), .S(DP_OP_422J2_124_3477_n1118) );
  FADDX1_HVT DP_OP_422J2_124_3477_U655 ( .A(DP_OP_422J2_124_3477_n1317), .B(
        DP_OP_422J2_124_3477_n1162), .CI(DP_OP_422J2_124_3477_n1160), .CO(
        DP_OP_422J2_124_3477_n1115), .S(DP_OP_422J2_124_3477_n1116) );
  FADDX1_HVT DP_OP_422J2_124_3477_U654 ( .A(DP_OP_422J2_124_3477_n1164), .B(
        DP_OP_422J2_124_3477_n1315), .CI(DP_OP_422J2_124_3477_n1154), .CO(
        DP_OP_422J2_124_3477_n1113), .S(DP_OP_422J2_124_3477_n1114) );
  FADDX1_HVT DP_OP_422J2_124_3477_U653 ( .A(DP_OP_422J2_124_3477_n1148), .B(
        DP_OP_422J2_124_3477_n1313), .CI(DP_OP_422J2_124_3477_n1146), .CO(
        DP_OP_422J2_124_3477_n1111), .S(DP_OP_422J2_124_3477_n1112) );
  FADDX1_HVT DP_OP_422J2_124_3477_U652 ( .A(DP_OP_422J2_124_3477_n1150), .B(
        DP_OP_422J2_124_3477_n1152), .CI(DP_OP_422J2_124_3477_n1144), .CO(
        DP_OP_422J2_124_3477_n1109), .S(DP_OP_422J2_124_3477_n1110) );
  FADDX1_HVT DP_OP_422J2_124_3477_U651 ( .A(DP_OP_422J2_124_3477_n1142), .B(
        DP_OP_422J2_124_3477_n1311), .CI(DP_OP_422J2_124_3477_n1309), .CO(
        DP_OP_422J2_124_3477_n1107), .S(DP_OP_422J2_124_3477_n1108) );
  FADDX1_HVT DP_OP_422J2_124_3477_U650 ( .A(DP_OP_422J2_124_3477_n1140), .B(
        DP_OP_422J2_124_3477_n1138), .CI(DP_OP_422J2_124_3477_n1307), .CO(
        DP_OP_422J2_124_3477_n1105), .S(DP_OP_422J2_124_3477_n1106) );
  FADDX1_HVT DP_OP_422J2_124_3477_U649 ( .A(DP_OP_422J2_124_3477_n1305), .B(
        DP_OP_422J2_124_3477_n1136), .CI(DP_OP_422J2_124_3477_n1303), .CO(
        DP_OP_422J2_124_3477_n1103), .S(DP_OP_422J2_124_3477_n1104) );
  FADDX1_HVT DP_OP_422J2_124_3477_U648 ( .A(DP_OP_422J2_124_3477_n1301), .B(
        DP_OP_422J2_124_3477_n1134), .CI(DP_OP_422J2_124_3477_n1132), .CO(
        DP_OP_422J2_124_3477_n1101), .S(DP_OP_422J2_124_3477_n1102) );
  FADDX1_HVT DP_OP_422J2_124_3477_U647 ( .A(DP_OP_422J2_124_3477_n1299), .B(
        DP_OP_422J2_124_3477_n1297), .CI(DP_OP_422J2_124_3477_n1295), .CO(
        DP_OP_422J2_124_3477_n1099), .S(DP_OP_422J2_124_3477_n1100) );
  FADDX1_HVT DP_OP_422J2_124_3477_U646 ( .A(DP_OP_422J2_124_3477_n1293), .B(
        DP_OP_422J2_124_3477_n1128), .CI(DP_OP_422J2_124_3477_n1126), .CO(
        DP_OP_422J2_124_3477_n1097), .S(DP_OP_422J2_124_3477_n1098) );
  FADDX1_HVT DP_OP_422J2_124_3477_U645 ( .A(DP_OP_422J2_124_3477_n1291), .B(
        DP_OP_422J2_124_3477_n1130), .CI(DP_OP_422J2_124_3477_n1289), .CO(
        DP_OP_422J2_124_3477_n1095), .S(DP_OP_422J2_124_3477_n1096) );
  FADDX1_HVT DP_OP_422J2_124_3477_U644 ( .A(DP_OP_422J2_124_3477_n1287), .B(
        DP_OP_422J2_124_3477_n1124), .CI(DP_OP_422J2_124_3477_n1120), .CO(
        DP_OP_422J2_124_3477_n1093), .S(DP_OP_422J2_124_3477_n1094) );
  FADDX1_HVT DP_OP_422J2_124_3477_U643 ( .A(DP_OP_422J2_124_3477_n1122), .B(
        DP_OP_422J2_124_3477_n1118), .CI(DP_OP_422J2_124_3477_n1285), .CO(
        DP_OP_422J2_124_3477_n1091), .S(DP_OP_422J2_124_3477_n1092) );
  FADDX1_HVT DP_OP_422J2_124_3477_U642 ( .A(DP_OP_422J2_124_3477_n1116), .B(
        DP_OP_422J2_124_3477_n1114), .CI(DP_OP_422J2_124_3477_n1112), .CO(
        DP_OP_422J2_124_3477_n1089), .S(DP_OP_422J2_124_3477_n1090) );
  FADDX1_HVT DP_OP_422J2_124_3477_U641 ( .A(DP_OP_422J2_124_3477_n1283), .B(
        DP_OP_422J2_124_3477_n1110), .CI(DP_OP_422J2_124_3477_n1108), .CO(
        DP_OP_422J2_124_3477_n1087), .S(DP_OP_422J2_124_3477_n1088) );
  FADDX1_HVT DP_OP_422J2_124_3477_U640 ( .A(DP_OP_422J2_124_3477_n1281), .B(
        DP_OP_422J2_124_3477_n1106), .CI(DP_OP_422J2_124_3477_n1279), .CO(
        DP_OP_422J2_124_3477_n1085), .S(DP_OP_422J2_124_3477_n1086) );
  FADDX1_HVT DP_OP_422J2_124_3477_U639 ( .A(DP_OP_422J2_124_3477_n1277), .B(
        DP_OP_422J2_124_3477_n1104), .CI(DP_OP_422J2_124_3477_n1275), .CO(
        DP_OP_422J2_124_3477_n1083), .S(DP_OP_422J2_124_3477_n1084) );
  FADDX1_HVT DP_OP_422J2_124_3477_U638 ( .A(DP_OP_422J2_124_3477_n1273), .B(
        DP_OP_422J2_124_3477_n1102), .CI(DP_OP_422J2_124_3477_n1100), .CO(
        DP_OP_422J2_124_3477_n1081), .S(DP_OP_422J2_124_3477_n1082) );
  FADDX1_HVT DP_OP_422J2_124_3477_U637 ( .A(DP_OP_422J2_124_3477_n1271), .B(
        DP_OP_422J2_124_3477_n1098), .CI(DP_OP_422J2_124_3477_n1269), .CO(
        DP_OP_422J2_124_3477_n1079), .S(DP_OP_422J2_124_3477_n1080) );
  FADDX1_HVT DP_OP_422J2_124_3477_U636 ( .A(DP_OP_422J2_124_3477_n1096), .B(
        DP_OP_422J2_124_3477_n1094), .CI(DP_OP_422J2_124_3477_n1267), .CO(
        DP_OP_422J2_124_3477_n1077), .S(DP_OP_422J2_124_3477_n1078) );
  FADDX1_HVT DP_OP_422J2_124_3477_U635 ( .A(DP_OP_422J2_124_3477_n1092), .B(
        DP_OP_422J2_124_3477_n1090), .CI(DP_OP_422J2_124_3477_n1088), .CO(
        DP_OP_422J2_124_3477_n1075), .S(DP_OP_422J2_124_3477_n1076) );
  FADDX1_HVT DP_OP_422J2_124_3477_U634 ( .A(DP_OP_422J2_124_3477_n1265), .B(
        DP_OP_422J2_124_3477_n1086), .CI(DP_OP_422J2_124_3477_n1263), .CO(
        DP_OP_422J2_124_3477_n1073), .S(DP_OP_422J2_124_3477_n1074) );
  FADDX1_HVT DP_OP_422J2_124_3477_U633 ( .A(DP_OP_422J2_124_3477_n1084), .B(
        DP_OP_422J2_124_3477_n1261), .CI(DP_OP_422J2_124_3477_n1082), .CO(
        DP_OP_422J2_124_3477_n1071), .S(DP_OP_422J2_124_3477_n1072) );
  FADDX1_HVT DP_OP_422J2_124_3477_U632 ( .A(DP_OP_422J2_124_3477_n1259), .B(
        DP_OP_422J2_124_3477_n1080), .CI(DP_OP_422J2_124_3477_n1078), .CO(
        DP_OP_422J2_124_3477_n1069), .S(DP_OP_422J2_124_3477_n1070) );
  FADDX1_HVT DP_OP_422J2_124_3477_U631 ( .A(DP_OP_422J2_124_3477_n1257), .B(
        DP_OP_422J2_124_3477_n1076), .CI(DP_OP_422J2_124_3477_n1255), .CO(
        DP_OP_422J2_124_3477_n1067), .S(DP_OP_422J2_124_3477_n1068) );
  FADDX1_HVT DP_OP_422J2_124_3477_U630 ( .A(DP_OP_422J2_124_3477_n1074), .B(
        DP_OP_422J2_124_3477_n1072), .CI(DP_OP_422J2_124_3477_n1253), .CO(
        DP_OP_422J2_124_3477_n1065), .S(DP_OP_422J2_124_3477_n1066) );
  FADDX1_HVT DP_OP_422J2_124_3477_U629 ( .A(DP_OP_422J2_124_3477_n1070), .B(
        DP_OP_422J2_124_3477_n1251), .CI(DP_OP_422J2_124_3477_n1068), .CO(
        DP_OP_422J2_124_3477_n1063), .S(DP_OP_422J2_124_3477_n1064) );
  OR2X1_HVT DP_OP_422J2_124_3477_U628 ( .A1(DP_OP_422J2_124_3477_n2703), .A2(
        DP_OP_422J2_124_3477_n2002), .Y(DP_OP_422J2_124_3477_n1061) );
  FADDX1_HVT DP_OP_422J2_124_3477_U626 ( .A(DP_OP_422J2_124_3477_n2835), .B(
        DP_OP_422J2_124_3477_n1826), .CI(DP_OP_422J2_124_3477_n2747), .CO(
        DP_OP_422J2_124_3477_n1059), .S(DP_OP_422J2_124_3477_n1060) );
  FADDX1_HVT DP_OP_422J2_124_3477_U625 ( .A(DP_OP_422J2_124_3477_n2617), .B(
        DP_OP_422J2_124_3477_n2441), .CI(DP_OP_422J2_124_3477_n1958), .CO(
        DP_OP_422J2_124_3477_n1057), .S(DP_OP_422J2_124_3477_n1058) );
  FADDX1_HVT DP_OP_422J2_124_3477_U624 ( .A(DP_OP_422J2_124_3477_n1870), .B(
        DP_OP_422J2_124_3477_n2485), .CI(DP_OP_422J2_124_3477_n2177), .CO(
        DP_OP_422J2_124_3477_n1055), .S(DP_OP_422J2_124_3477_n1056) );
  FADDX1_HVT DP_OP_422J2_124_3477_U623 ( .A(DP_OP_422J2_124_3477_n2353), .B(
        DP_OP_422J2_124_3477_n1914), .CI(DP_OP_422J2_124_3477_n2573), .CO(
        DP_OP_422J2_124_3477_n1053), .S(DP_OP_422J2_124_3477_n1054) );
  FADDX1_HVT DP_OP_422J2_124_3477_U622 ( .A(DP_OP_422J2_124_3477_n2133), .B(
        DP_OP_422J2_124_3477_n2529), .CI(DP_OP_422J2_124_3477_n2045), .CO(
        DP_OP_422J2_124_3477_n1051), .S(DP_OP_422J2_124_3477_n1052) );
  FADDX1_HVT DP_OP_422J2_124_3477_U621 ( .A(DP_OP_422J2_124_3477_n2089), .B(
        DP_OP_422J2_124_3477_n2265), .CI(DP_OP_422J2_124_3477_n2879), .CO(
        DP_OP_422J2_124_3477_n1049), .S(DP_OP_422J2_124_3477_n1050) );
  FADDX1_HVT DP_OP_422J2_124_3477_U620 ( .A(DP_OP_422J2_124_3477_n2661), .B(
        DP_OP_422J2_124_3477_n2309), .CI(DP_OP_422J2_124_3477_n2791), .CO(
        DP_OP_422J2_124_3477_n1047), .S(DP_OP_422J2_124_3477_n1048) );
  FADDX1_HVT DP_OP_422J2_124_3477_U619 ( .A(DP_OP_422J2_124_3477_n2397), .B(
        DP_OP_422J2_124_3477_n1965), .CI(DP_OP_422J2_124_3477_n2580), .CO(
        DP_OP_422J2_124_3477_n1045), .S(DP_OP_422J2_124_3477_n1046) );
  FADDX1_HVT DP_OP_422J2_124_3477_U618 ( .A(DP_OP_422J2_124_3477_n2638), .B(
        DP_OP_422J2_124_3477_n2147), .CI(DP_OP_422J2_124_3477_n2272), .CO(
        DP_OP_422J2_124_3477_n1043), .S(DP_OP_422J2_124_3477_n1044) );
  FADDX1_HVT DP_OP_422J2_124_3477_U617 ( .A(DP_OP_422J2_124_3477_n2198), .B(
        DP_OP_422J2_124_3477_n2411), .CI(DP_OP_422J2_124_3477_n2286), .CO(
        DP_OP_422J2_124_3477_n1041), .S(DP_OP_422J2_124_3477_n1042) );
  FADDX1_HVT DP_OP_422J2_124_3477_U616 ( .A(DP_OP_422J2_124_3477_n2550), .B(
        DP_OP_422J2_124_3477_n2536), .CI(DP_OP_422J2_124_3477_n2140), .CO(
        DP_OP_422J2_124_3477_n1039), .S(DP_OP_422J2_124_3477_n1040) );
  FADDX1_HVT DP_OP_422J2_124_3477_U615 ( .A(DP_OP_422J2_124_3477_n2330), .B(
        DP_OP_422J2_124_3477_n2724), .CI(DP_OP_422J2_124_3477_n2066), .CO(
        DP_OP_422J2_124_3477_n1037), .S(DP_OP_422J2_124_3477_n1038) );
  FADDX1_HVT DP_OP_422J2_124_3477_U614 ( .A(DP_OP_422J2_124_3477_n1847), .B(
        DP_OP_422J2_124_3477_n2221), .CI(DP_OP_422J2_124_3477_n2506), .CO(
        DP_OP_422J2_124_3477_n1035), .S(DP_OP_422J2_124_3477_n1036) );
  FADDX1_HVT DP_OP_422J2_124_3477_U613 ( .A(DP_OP_422J2_124_3477_n2462), .B(
        DP_OP_422J2_124_3477_n1782), .CI(DP_OP_422J2_124_3477_n2228), .CO(
        DP_OP_422J2_124_3477_n1033), .S(DP_OP_422J2_124_3477_n1034) );
  FADDX1_HVT DP_OP_422J2_124_3477_U612 ( .A(DP_OP_422J2_124_3477_n2418), .B(
        DP_OP_422J2_124_3477_n1840), .CI(DP_OP_422J2_124_3477_n2768), .CO(
        DP_OP_422J2_124_3477_n1031), .S(DP_OP_422J2_124_3477_n1032) );
  FADDX1_HVT DP_OP_422J2_124_3477_U611 ( .A(DP_OP_422J2_124_3477_n2110), .B(
        DP_OP_422J2_124_3477_n2499), .CI(DP_OP_422J2_124_3477_n2856), .CO(
        DP_OP_422J2_124_3477_n1029), .S(DP_OP_422J2_124_3477_n1030) );
  FADDX1_HVT DP_OP_422J2_124_3477_U610 ( .A(DP_OP_422J2_124_3477_n2594), .B(
        DP_OP_422J2_124_3477_n2682), .CI(DP_OP_422J2_124_3477_n1891), .CO(
        DP_OP_422J2_124_3477_n1027), .S(DP_OP_422J2_124_3477_n1028) );
  FADDX1_HVT DP_OP_422J2_124_3477_U609 ( .A(DP_OP_422J2_124_3477_n2842), .B(
        DP_OP_422J2_124_3477_n2587), .CI(DP_OP_422J2_124_3477_n2448), .CO(
        DP_OP_422J2_124_3477_n1025), .S(DP_OP_422J2_124_3477_n1026) );
  FADDX1_HVT DP_OP_422J2_124_3477_U608 ( .A(DP_OP_422J2_124_3477_n2886), .B(
        DP_OP_422J2_124_3477_n2754), .CI(DP_OP_422J2_124_3477_n2096), .CO(
        DP_OP_422J2_124_3477_n1023), .S(DP_OP_422J2_124_3477_n1024) );
  FADDX1_HVT DP_OP_422J2_124_3477_U607 ( .A(DP_OP_422J2_124_3477_n2631), .B(
        DP_OP_422J2_124_3477_n1979), .CI(DP_OP_422J2_124_3477_n2022), .CO(
        DP_OP_422J2_124_3477_n1021), .S(DP_OP_422J2_124_3477_n1022) );
  FADDX1_HVT DP_OP_422J2_124_3477_U606 ( .A(DP_OP_422J2_124_3477_n2323), .B(
        DP_OP_422J2_124_3477_n2059), .CI(DP_OP_422J2_124_3477_n2103), .CO(
        DP_OP_422J2_124_3477_n1019), .S(DP_OP_422J2_124_3477_n1020) );
  FADDX1_HVT DP_OP_422J2_124_3477_U605 ( .A(DP_OP_422J2_124_3477_n1884), .B(
        DP_OP_422J2_124_3477_n2052), .CI(DP_OP_422J2_124_3477_n1921), .CO(
        DP_OP_422J2_124_3477_n1017), .S(DP_OP_422J2_124_3477_n1018) );
  FADDX1_HVT DP_OP_422J2_124_3477_U604 ( .A(DP_OP_422J2_124_3477_n2492), .B(
        DP_OP_422J2_124_3477_n2316), .CI(DP_OP_422J2_124_3477_n2184), .CO(
        DP_OP_422J2_124_3477_n1015), .S(DP_OP_422J2_124_3477_n1016) );
  FADDX1_HVT DP_OP_422J2_124_3477_U603 ( .A(DP_OP_422J2_124_3477_n2360), .B(
        DP_OP_422J2_124_3477_n2668), .CI(DP_OP_422J2_124_3477_n1833), .CO(
        DP_OP_422J2_124_3477_n1013), .S(DP_OP_422J2_124_3477_n1014) );
  FADDX1_HVT DP_OP_422J2_124_3477_U602 ( .A(DP_OP_422J2_124_3477_n2675), .B(
        DP_OP_422J2_124_3477_n2849), .CI(DP_OP_422J2_124_3477_n2235), .CO(
        DP_OP_422J2_124_3477_n1011), .S(DP_OP_422J2_124_3477_n1012) );
  FADDX1_HVT DP_OP_422J2_124_3477_U601 ( .A(DP_OP_422J2_124_3477_n2242), .B(
        DP_OP_422J2_124_3477_n2893), .CI(DP_OP_422J2_124_3477_n2191), .CO(
        DP_OP_422J2_124_3477_n1009), .S(DP_OP_422J2_124_3477_n1010) );
  FADDX1_HVT DP_OP_422J2_124_3477_U600 ( .A(DP_OP_422J2_124_3477_n2455), .B(
        DP_OP_422J2_124_3477_n2279), .CI(DP_OP_422J2_124_3477_n2367), .CO(
        DP_OP_422J2_124_3477_n1007), .S(DP_OP_422J2_124_3477_n1008) );
  FADDX1_HVT DP_OP_422J2_124_3477_U599 ( .A(DP_OP_422J2_124_3477_n2710), .B(
        DP_OP_422J2_124_3477_n2761), .CI(DP_OP_422J2_124_3477_n2008), .CO(
        DP_OP_422J2_124_3477_n1005), .S(DP_OP_422J2_124_3477_n1006) );
  FADDX1_HVT DP_OP_422J2_124_3477_U598 ( .A(DP_OP_422J2_124_3477_n2543), .B(
        DP_OP_422J2_124_3477_n2805), .CI(DP_OP_422J2_124_3477_n2624), .CO(
        DP_OP_422J2_124_3477_n1003), .S(DP_OP_422J2_124_3477_n1004) );
  FADDX1_HVT DP_OP_422J2_124_3477_U597 ( .A(DP_OP_422J2_124_3477_n1935), .B(
        DP_OP_422J2_124_3477_n2154), .CI(DP_OP_422J2_124_3477_n2798), .CO(
        DP_OP_422J2_124_3477_n1001), .S(DP_OP_422J2_124_3477_n1002) );
  FADDX1_HVT DP_OP_422J2_124_3477_U596 ( .A(DP_OP_422J2_124_3477_n2404), .B(
        DP_OP_422J2_124_3477_n1972), .CI(DP_OP_422J2_124_3477_n1249), .CO(
        DP_OP_422J2_124_3477_n999), .S(DP_OP_422J2_124_3477_n1000) );
  FADDX1_HVT DP_OP_422J2_124_3477_U595 ( .A(DP_OP_422J2_124_3477_n2015), .B(
        DP_OP_422J2_124_3477_n2717), .CI(DP_OP_422J2_124_3477_n2812), .CO(
        DP_OP_422J2_124_3477_n997), .S(DP_OP_422J2_124_3477_n998) );
  FADDX1_HVT DP_OP_422J2_124_3477_U594 ( .A(DP_OP_422J2_124_3477_n1928), .B(
        DP_OP_422J2_124_3477_n2900), .CI(DP_OP_422J2_124_3477_n2374), .CO(
        DP_OP_422J2_124_3477_n995), .S(DP_OP_422J2_124_3477_n996) );
  FADDX1_HVT DP_OP_422J2_124_3477_U593 ( .A(DP_OP_422J2_124_3477_n1877), .B(
        DP_OP_422J2_124_3477_n1247), .CI(DP_OP_422J2_124_3477_n1245), .CO(
        DP_OP_422J2_124_3477_n993), .S(DP_OP_422J2_124_3477_n994) );
  FADDX1_HVT DP_OP_422J2_124_3477_U592 ( .A(DP_OP_422J2_124_3477_n1243), .B(
        DP_OP_422J2_124_3477_n1235), .CI(DP_OP_422J2_124_3477_n1062), .CO(
        DP_OP_422J2_124_3477_n991), .S(DP_OP_422J2_124_3477_n992) );
  FADDX1_HVT DP_OP_422J2_124_3477_U591 ( .A(DP_OP_422J2_124_3477_n1241), .B(
        DP_OP_422J2_124_3477_n1237), .CI(DP_OP_422J2_124_3477_n1239), .CO(
        DP_OP_422J2_124_3477_n989), .S(DP_OP_422J2_124_3477_n990) );
  FADDX1_HVT DP_OP_422J2_124_3477_U590 ( .A(DP_OP_422J2_124_3477_n1233), .B(
        DP_OP_422J2_124_3477_n1207), .CI(DP_OP_422J2_124_3477_n1209), .CO(
        DP_OP_422J2_124_3477_n987), .S(DP_OP_422J2_124_3477_n988) );
  FADDX1_HVT DP_OP_422J2_124_3477_U589 ( .A(DP_OP_422J2_124_3477_n1231), .B(
        DP_OP_422J2_124_3477_n1211), .CI(DP_OP_422J2_124_3477_n1213), .CO(
        DP_OP_422J2_124_3477_n985), .S(DP_OP_422J2_124_3477_n986) );
  FADDX1_HVT DP_OP_422J2_124_3477_U588 ( .A(DP_OP_422J2_124_3477_n1229), .B(
        DP_OP_422J2_124_3477_n1215), .CI(DP_OP_422J2_124_3477_n1217), .CO(
        DP_OP_422J2_124_3477_n983), .S(DP_OP_422J2_124_3477_n984) );
  FADDX1_HVT DP_OP_422J2_124_3477_U587 ( .A(DP_OP_422J2_124_3477_n1227), .B(
        DP_OP_422J2_124_3477_n1219), .CI(DP_OP_422J2_124_3477_n1221), .CO(
        DP_OP_422J2_124_3477_n981), .S(DP_OP_422J2_124_3477_n982) );
  FADDX1_HVT DP_OP_422J2_124_3477_U586 ( .A(DP_OP_422J2_124_3477_n1223), .B(
        DP_OP_422J2_124_3477_n1225), .CI(DP_OP_422J2_124_3477_n1203), .CO(
        DP_OP_422J2_124_3477_n979), .S(DP_OP_422J2_124_3477_n980) );
  FADDX1_HVT DP_OP_422J2_124_3477_U585 ( .A(DP_OP_422J2_124_3477_n1205), .B(
        DP_OP_422J2_124_3477_n1054), .CI(DP_OP_422J2_124_3477_n1183), .CO(
        DP_OP_422J2_124_3477_n977), .S(DP_OP_422J2_124_3477_n978) );
  FADDX1_HVT DP_OP_422J2_124_3477_U584 ( .A(DP_OP_422J2_124_3477_n1201), .B(
        DP_OP_422J2_124_3477_n1058), .CI(DP_OP_422J2_124_3477_n1185), .CO(
        DP_OP_422J2_124_3477_n975), .S(DP_OP_422J2_124_3477_n976) );
  FADDX1_HVT DP_OP_422J2_124_3477_U583 ( .A(DP_OP_422J2_124_3477_n1199), .B(
        DP_OP_422J2_124_3477_n1052), .CI(DP_OP_422J2_124_3477_n1187), .CO(
        DP_OP_422J2_124_3477_n973), .S(DP_OP_422J2_124_3477_n974) );
  FADDX1_HVT DP_OP_422J2_124_3477_U582 ( .A(DP_OP_422J2_124_3477_n1197), .B(
        DP_OP_422J2_124_3477_n1056), .CI(DP_OP_422J2_124_3477_n1048), .CO(
        DP_OP_422J2_124_3477_n971), .S(DP_OP_422J2_124_3477_n972) );
  FADDX1_HVT DP_OP_422J2_124_3477_U581 ( .A(DP_OP_422J2_124_3477_n1195), .B(
        DP_OP_422J2_124_3477_n1060), .CI(DP_OP_422J2_124_3477_n1050), .CO(
        DP_OP_422J2_124_3477_n969), .S(DP_OP_422J2_124_3477_n970) );
  FADDX1_HVT DP_OP_422J2_124_3477_U580 ( .A(DP_OP_422J2_124_3477_n1191), .B(
        DP_OP_422J2_124_3477_n1193), .CI(DP_OP_422J2_124_3477_n1189), .CO(
        DP_OP_422J2_124_3477_n967), .S(DP_OP_422J2_124_3477_n968) );
  FADDX1_HVT DP_OP_422J2_124_3477_U579 ( .A(DP_OP_422J2_124_3477_n1046), .B(
        DP_OP_422J2_124_3477_n1022), .CI(DP_OP_422J2_124_3477_n1020), .CO(
        DP_OP_422J2_124_3477_n965), .S(DP_OP_422J2_124_3477_n966) );
  FADDX1_HVT DP_OP_422J2_124_3477_U578 ( .A(DP_OP_422J2_124_3477_n1036), .B(
        DP_OP_422J2_124_3477_n1034), .CI(DP_OP_422J2_124_3477_n1030), .CO(
        DP_OP_422J2_124_3477_n963), .S(DP_OP_422J2_124_3477_n964) );
  FADDX1_HVT DP_OP_422J2_124_3477_U577 ( .A(DP_OP_422J2_124_3477_n1032), .B(
        DP_OP_422J2_124_3477_n1026), .CI(DP_OP_422J2_124_3477_n1028), .CO(
        DP_OP_422J2_124_3477_n961), .S(DP_OP_422J2_124_3477_n962) );
  FADDX1_HVT DP_OP_422J2_124_3477_U576 ( .A(DP_OP_422J2_124_3477_n1024), .B(
        DP_OP_422J2_124_3477_n1044), .CI(DP_OP_422J2_124_3477_n1042), .CO(
        DP_OP_422J2_124_3477_n959), .S(DP_OP_422J2_124_3477_n960) );
  FADDX1_HVT DP_OP_422J2_124_3477_U575 ( .A(DP_OP_422J2_124_3477_n1040), .B(
        DP_OP_422J2_124_3477_n1038), .CI(DP_OP_422J2_124_3477_n1018), .CO(
        DP_OP_422J2_124_3477_n957), .S(DP_OP_422J2_124_3477_n958) );
  FADDX1_HVT DP_OP_422J2_124_3477_U574 ( .A(DP_OP_422J2_124_3477_n1016), .B(
        DP_OP_422J2_124_3477_n1002), .CI(DP_OP_422J2_124_3477_n996), .CO(
        DP_OP_422J2_124_3477_n955), .S(DP_OP_422J2_124_3477_n956) );
  FADDX1_HVT DP_OP_422J2_124_3477_U573 ( .A(DP_OP_422J2_124_3477_n1014), .B(
        DP_OP_422J2_124_3477_n1006), .CI(DP_OP_422J2_124_3477_n1000), .CO(
        DP_OP_422J2_124_3477_n953), .S(DP_OP_422J2_124_3477_n954) );
  FADDX1_HVT DP_OP_422J2_124_3477_U572 ( .A(DP_OP_422J2_124_3477_n1012), .B(
        DP_OP_422J2_124_3477_n1004), .CI(DP_OP_422J2_124_3477_n998), .CO(
        DP_OP_422J2_124_3477_n951), .S(DP_OP_422J2_124_3477_n952) );
  FADDX1_HVT DP_OP_422J2_124_3477_U571 ( .A(DP_OP_422J2_124_3477_n1010), .B(
        DP_OP_422J2_124_3477_n1008), .CI(DP_OP_422J2_124_3477_n1181), .CO(
        DP_OP_422J2_124_3477_n949), .S(DP_OP_422J2_124_3477_n950) );
  FADDX1_HVT DP_OP_422J2_124_3477_U570 ( .A(DP_OP_422J2_124_3477_n1179), .B(
        DP_OP_422J2_124_3477_n1177), .CI(DP_OP_422J2_124_3477_n1175), .CO(
        DP_OP_422J2_124_3477_n947), .S(DP_OP_422J2_124_3477_n948) );
  FADDX1_HVT DP_OP_422J2_124_3477_U569 ( .A(DP_OP_422J2_124_3477_n1173), .B(
        DP_OP_422J2_124_3477_n1167), .CI(DP_OP_422J2_124_3477_n1169), .CO(
        DP_OP_422J2_124_3477_n945), .S(DP_OP_422J2_124_3477_n946) );
  FADDX1_HVT DP_OP_422J2_124_3477_U568 ( .A(DP_OP_422J2_124_3477_n1171), .B(
        DP_OP_422J2_124_3477_n994), .CI(DP_OP_422J2_124_3477_n1165), .CO(
        DP_OP_422J2_124_3477_n943), .S(DP_OP_422J2_124_3477_n944) );
  FADDX1_HVT DP_OP_422J2_124_3477_U567 ( .A(DP_OP_422J2_124_3477_n1163), .B(
        DP_OP_422J2_124_3477_n992), .CI(DP_OP_422J2_124_3477_n990), .CO(
        DP_OP_422J2_124_3477_n941), .S(DP_OP_422J2_124_3477_n942) );
  FADDX1_HVT DP_OP_422J2_124_3477_U566 ( .A(DP_OP_422J2_124_3477_n1161), .B(
        DP_OP_422J2_124_3477_n1157), .CI(DP_OP_422J2_124_3477_n1155), .CO(
        DP_OP_422J2_124_3477_n939), .S(DP_OP_422J2_124_3477_n940) );
  FADDX1_HVT DP_OP_422J2_124_3477_U565 ( .A(DP_OP_422J2_124_3477_n1159), .B(
        DP_OP_422J2_124_3477_n1153), .CI(DP_OP_422J2_124_3477_n988), .CO(
        DP_OP_422J2_124_3477_n937), .S(DP_OP_422J2_124_3477_n938) );
  FADDX1_HVT DP_OP_422J2_124_3477_U564 ( .A(DP_OP_422J2_124_3477_n1151), .B(
        DP_OP_422J2_124_3477_n984), .CI(DP_OP_422J2_124_3477_n980), .CO(
        DP_OP_422J2_124_3477_n935), .S(DP_OP_422J2_124_3477_n936) );
  FADDX1_HVT DP_OP_422J2_124_3477_U563 ( .A(DP_OP_422J2_124_3477_n1149), .B(
        DP_OP_422J2_124_3477_n982), .CI(DP_OP_422J2_124_3477_n986), .CO(
        DP_OP_422J2_124_3477_n933), .S(DP_OP_422J2_124_3477_n934) );
  FADDX1_HVT DP_OP_422J2_124_3477_U562 ( .A(DP_OP_422J2_124_3477_n1147), .B(
        DP_OP_422J2_124_3477_n1145), .CI(DP_OP_422J2_124_3477_n1143), .CO(
        DP_OP_422J2_124_3477_n931), .S(DP_OP_422J2_124_3477_n932) );
  FADDX1_HVT DP_OP_422J2_124_3477_U561 ( .A(DP_OP_422J2_124_3477_n978), .B(
        DP_OP_422J2_124_3477_n968), .CI(DP_OP_422J2_124_3477_n1137), .CO(
        DP_OP_422J2_124_3477_n929), .S(DP_OP_422J2_124_3477_n930) );
  FADDX1_HVT DP_OP_422J2_124_3477_U560 ( .A(DP_OP_422J2_124_3477_n1141), .B(
        DP_OP_422J2_124_3477_n972), .CI(DP_OP_422J2_124_3477_n970), .CO(
        DP_OP_422J2_124_3477_n927), .S(DP_OP_422J2_124_3477_n928) );
  FADDX1_HVT DP_OP_422J2_124_3477_U559 ( .A(DP_OP_422J2_124_3477_n976), .B(
        DP_OP_422J2_124_3477_n1139), .CI(DP_OP_422J2_124_3477_n974), .CO(
        DP_OP_422J2_124_3477_n925), .S(DP_OP_422J2_124_3477_n926) );
  FADDX1_HVT DP_OP_422J2_124_3477_U558 ( .A(DP_OP_422J2_124_3477_n966), .B(
        DP_OP_422J2_124_3477_n1135), .CI(DP_OP_422J2_124_3477_n958), .CO(
        DP_OP_422J2_124_3477_n923), .S(DP_OP_422J2_124_3477_n924) );
  FADDX1_HVT DP_OP_422J2_124_3477_U557 ( .A(DP_OP_422J2_124_3477_n960), .B(
        DP_OP_422J2_124_3477_n964), .CI(DP_OP_422J2_124_3477_n962), .CO(
        DP_OP_422J2_124_3477_n921), .S(DP_OP_422J2_124_3477_n922) );
  FADDX1_HVT DP_OP_422J2_124_3477_U556 ( .A(DP_OP_422J2_124_3477_n956), .B(
        DP_OP_422J2_124_3477_n950), .CI(DP_OP_422J2_124_3477_n1131), .CO(
        DP_OP_422J2_124_3477_n919), .S(DP_OP_422J2_124_3477_n920) );
  FADDX1_HVT DP_OP_422J2_124_3477_U555 ( .A(DP_OP_422J2_124_3477_n954), .B(
        DP_OP_422J2_124_3477_n952), .CI(DP_OP_422J2_124_3477_n1133), .CO(
        DP_OP_422J2_124_3477_n917), .S(DP_OP_422J2_124_3477_n918) );
  FADDX1_HVT DP_OP_422J2_124_3477_U554 ( .A(DP_OP_422J2_124_3477_n1129), .B(
        DP_OP_422J2_124_3477_n948), .CI(DP_OP_422J2_124_3477_n1125), .CO(
        DP_OP_422J2_124_3477_n915), .S(DP_OP_422J2_124_3477_n916) );
  FADDX1_HVT DP_OP_422J2_124_3477_U553 ( .A(DP_OP_422J2_124_3477_n1127), .B(
        DP_OP_422J2_124_3477_n1123), .CI(DP_OP_422J2_124_3477_n1121), .CO(
        DP_OP_422J2_124_3477_n913), .S(DP_OP_422J2_124_3477_n914) );
  FADDX1_HVT DP_OP_422J2_124_3477_U552 ( .A(DP_OP_422J2_124_3477_n1119), .B(
        DP_OP_422J2_124_3477_n946), .CI(DP_OP_422J2_124_3477_n944), .CO(
        DP_OP_422J2_124_3477_n911), .S(DP_OP_422J2_124_3477_n912) );
  FADDX1_HVT DP_OP_422J2_124_3477_U551 ( .A(DP_OP_422J2_124_3477_n1117), .B(
        DP_OP_422J2_124_3477_n940), .CI(DP_OP_422J2_124_3477_n1113), .CO(
        DP_OP_422J2_124_3477_n909), .S(DP_OP_422J2_124_3477_n910) );
  FADDX1_HVT DP_OP_422J2_124_3477_U550 ( .A(DP_OP_422J2_124_3477_n1115), .B(
        DP_OP_422J2_124_3477_n942), .CI(DP_OP_422J2_124_3477_n938), .CO(
        DP_OP_422J2_124_3477_n907), .S(DP_OP_422J2_124_3477_n908) );
  FADDX1_HVT DP_OP_422J2_124_3477_U549 ( .A(DP_OP_422J2_124_3477_n936), .B(
        DP_OP_422J2_124_3477_n934), .CI(DP_OP_422J2_124_3477_n932), .CO(
        DP_OP_422J2_124_3477_n905), .S(DP_OP_422J2_124_3477_n906) );
  FADDX1_HVT DP_OP_422J2_124_3477_U548 ( .A(DP_OP_422J2_124_3477_n1111), .B(
        DP_OP_422J2_124_3477_n1109), .CI(DP_OP_422J2_124_3477_n930), .CO(
        DP_OP_422J2_124_3477_n903), .S(DP_OP_422J2_124_3477_n904) );
  FADDX1_HVT DP_OP_422J2_124_3477_U547 ( .A(DP_OP_422J2_124_3477_n1107), .B(
        DP_OP_422J2_124_3477_n928), .CI(DP_OP_422J2_124_3477_n1105), .CO(
        DP_OP_422J2_124_3477_n901), .S(DP_OP_422J2_124_3477_n902) );
  FADDX1_HVT DP_OP_422J2_124_3477_U546 ( .A(DP_OP_422J2_124_3477_n926), .B(
        DP_OP_422J2_124_3477_n924), .CI(DP_OP_422J2_124_3477_n922), .CO(
        DP_OP_422J2_124_3477_n899), .S(DP_OP_422J2_124_3477_n900) );
  FADDX1_HVT DP_OP_422J2_124_3477_U545 ( .A(DP_OP_422J2_124_3477_n1103), .B(
        DP_OP_422J2_124_3477_n920), .CI(DP_OP_422J2_124_3477_n918), .CO(
        DP_OP_422J2_124_3477_n897), .S(DP_OP_422J2_124_3477_n898) );
  FADDX1_HVT DP_OP_422J2_124_3477_U544 ( .A(DP_OP_422J2_124_3477_n1101), .B(
        DP_OP_422J2_124_3477_n1099), .CI(DP_OP_422J2_124_3477_n1097), .CO(
        DP_OP_422J2_124_3477_n895), .S(DP_OP_422J2_124_3477_n896) );
  FADDX1_HVT DP_OP_422J2_124_3477_U543 ( .A(DP_OP_422J2_124_3477_n916), .B(
        DP_OP_422J2_124_3477_n1095), .CI(DP_OP_422J2_124_3477_n914), .CO(
        DP_OP_422J2_124_3477_n893), .S(DP_OP_422J2_124_3477_n894) );
  FADDX1_HVT DP_OP_422J2_124_3477_U542 ( .A(DP_OP_422J2_124_3477_n1093), .B(
        DP_OP_422J2_124_3477_n912), .CI(DP_OP_422J2_124_3477_n1091), .CO(
        DP_OP_422J2_124_3477_n891), .S(DP_OP_422J2_124_3477_n892) );
  FADDX1_HVT DP_OP_422J2_124_3477_U541 ( .A(DP_OP_422J2_124_3477_n910), .B(
        DP_OP_422J2_124_3477_n908), .CI(DP_OP_422J2_124_3477_n1089), .CO(
        DP_OP_422J2_124_3477_n889), .S(DP_OP_422J2_124_3477_n890) );
  FADDX1_HVT DP_OP_422J2_124_3477_U540 ( .A(DP_OP_422J2_124_3477_n906), .B(
        DP_OP_422J2_124_3477_n1087), .CI(DP_OP_422J2_124_3477_n904), .CO(
        DP_OP_422J2_124_3477_n887), .S(DP_OP_422J2_124_3477_n888) );
  FADDX1_HVT DP_OP_422J2_124_3477_U539 ( .A(DP_OP_422J2_124_3477_n902), .B(
        DP_OP_422J2_124_3477_n1085), .CI(DP_OP_422J2_124_3477_n900), .CO(
        DP_OP_422J2_124_3477_n885), .S(DP_OP_422J2_124_3477_n886) );
  FADDX1_HVT DP_OP_422J2_124_3477_U538 ( .A(DP_OP_422J2_124_3477_n1083), .B(
        DP_OP_422J2_124_3477_n898), .CI(DP_OP_422J2_124_3477_n1081), .CO(
        DP_OP_422J2_124_3477_n883), .S(DP_OP_422J2_124_3477_n884) );
  FADDX1_HVT DP_OP_422J2_124_3477_U537 ( .A(DP_OP_422J2_124_3477_n896), .B(
        DP_OP_422J2_124_3477_n1079), .CI(DP_OP_422J2_124_3477_n894), .CO(
        DP_OP_422J2_124_3477_n881), .S(DP_OP_422J2_124_3477_n882) );
  FADDX1_HVT DP_OP_422J2_124_3477_U536 ( .A(DP_OP_422J2_124_3477_n1077), .B(
        DP_OP_422J2_124_3477_n892), .CI(DP_OP_422J2_124_3477_n890), .CO(
        DP_OP_422J2_124_3477_n879), .S(DP_OP_422J2_124_3477_n880) );
  FADDX1_HVT DP_OP_422J2_124_3477_U535 ( .A(DP_OP_422J2_124_3477_n1075), .B(
        DP_OP_422J2_124_3477_n888), .CI(DP_OP_422J2_124_3477_n1073), .CO(
        DP_OP_422J2_124_3477_n877), .S(DP_OP_422J2_124_3477_n878) );
  FADDX1_HVT DP_OP_422J2_124_3477_U534 ( .A(DP_OP_422J2_124_3477_n886), .B(
        DP_OP_422J2_124_3477_n1071), .CI(DP_OP_422J2_124_3477_n884), .CO(
        DP_OP_422J2_124_3477_n875), .S(DP_OP_422J2_124_3477_n876) );
  FADDX1_HVT DP_OP_422J2_124_3477_U533 ( .A(DP_OP_422J2_124_3477_n882), .B(
        DP_OP_422J2_124_3477_n1069), .CI(DP_OP_422J2_124_3477_n880), .CO(
        DP_OP_422J2_124_3477_n873), .S(DP_OP_422J2_124_3477_n874) );
  FADDX1_HVT DP_OP_422J2_124_3477_U532 ( .A(DP_OP_422J2_124_3477_n1067), .B(
        DP_OP_422J2_124_3477_n878), .CI(DP_OP_422J2_124_3477_n876), .CO(
        DP_OP_422J2_124_3477_n871), .S(DP_OP_422J2_124_3477_n872) );
  FADDX1_HVT DP_OP_422J2_124_3477_U531 ( .A(DP_OP_422J2_124_3477_n1065), .B(
        DP_OP_422J2_124_3477_n874), .CI(DP_OP_422J2_124_3477_n1063), .CO(
        DP_OP_422J2_124_3477_n869), .S(DP_OP_422J2_124_3477_n870) );
  FADDX1_HVT DP_OP_422J2_124_3477_U530 ( .A(DP_OP_422J2_124_3477_n2001), .B(
        DP_OP_422J2_124_3477_n2723), .CI(DP_OP_422J2_124_3477_n2505), .CO(
        DP_OP_422J2_124_3477_n867), .S(DP_OP_422J2_124_3477_n868) );
  FADDX1_HVT DP_OP_422J2_124_3477_U529 ( .A(DP_OP_422J2_124_3477_n2702), .B(
        DP_OP_422J2_124_3477_n1825), .CI(DP_OP_422J2_124_3477_n2767), .CO(
        DP_OP_422J2_124_3477_n865), .S(DP_OP_422J2_124_3477_n866) );
  FADDX1_HVT DP_OP_422J2_124_3477_U528 ( .A(DP_OP_422J2_124_3477_n1869), .B(
        DP_OP_422J2_124_3477_n2528), .CI(DP_OP_422J2_124_3477_n2855), .CO(
        DP_OP_422J2_124_3477_n863), .S(DP_OP_422J2_124_3477_n864) );
  FADDX1_HVT DP_OP_422J2_124_3477_U527 ( .A(DP_OP_422J2_124_3477_n2660), .B(
        DP_OP_422J2_124_3477_n2572), .CI(DP_OP_422J2_124_3477_n1890), .CO(
        DP_OP_422J2_124_3477_n861), .S(DP_OP_422J2_124_3477_n862) );
  FADDX1_HVT DP_OP_422J2_124_3477_U526 ( .A(DP_OP_422J2_124_3477_n2088), .B(
        DP_OP_422J2_124_3477_n2440), .CI(DP_OP_422J2_124_3477_n2746), .CO(
        DP_OP_422J2_124_3477_n859), .S(DP_OP_422J2_124_3477_n860) );
  FADDX1_HVT DP_OP_422J2_124_3477_U525 ( .A(DP_OP_422J2_124_3477_n2132), .B(
        DP_OP_422J2_124_3477_n1913), .CI(DP_OP_422J2_124_3477_n1957), .CO(
        DP_OP_422J2_124_3477_n857), .S(DP_OP_422J2_124_3477_n858) );
  FADDX1_HVT DP_OP_422J2_124_3477_U524 ( .A(DP_OP_422J2_124_3477_n2308), .B(
        DP_OP_422J2_124_3477_n2176), .CI(DP_OP_422J2_124_3477_n2484), .CO(
        DP_OP_422J2_124_3477_n855), .S(DP_OP_422J2_124_3477_n856) );
  FADDX1_HVT DP_OP_422J2_124_3477_U523 ( .A(DP_OP_422J2_124_3477_n2834), .B(
        DP_OP_422J2_124_3477_n2878), .CI(DP_OP_422J2_124_3477_n2044), .CO(
        DP_OP_422J2_124_3477_n853), .S(DP_OP_422J2_124_3477_n854) );
  FADDX1_HVT DP_OP_422J2_124_3477_U522 ( .A(DP_OP_422J2_124_3477_n2790), .B(
        DP_OP_422J2_124_3477_n2681), .CI(DP_OP_422J2_124_3477_n1978), .CO(
        DP_OP_422J2_124_3477_n851), .S(DP_OP_422J2_124_3477_n852) );
  FADDX1_HVT DP_OP_422J2_124_3477_U521 ( .A(DP_OP_422J2_124_3477_n2616), .B(
        DP_OP_422J2_124_3477_n2109), .CI(DP_OP_422J2_124_3477_n2021), .CO(
        DP_OP_422J2_124_3477_n849), .S(DP_OP_422J2_124_3477_n850) );
  FADDX1_HVT DP_OP_422J2_124_3477_U520 ( .A(DP_OP_422J2_124_3477_n2352), .B(
        DP_OP_422J2_124_3477_n2461), .CI(DP_OP_422J2_124_3477_n2417), .CO(
        DP_OP_422J2_124_3477_n847), .S(DP_OP_422J2_124_3477_n848) );
  FADDX1_HVT DP_OP_422J2_124_3477_U519 ( .A(DP_OP_422J2_124_3477_n2264), .B(
        DP_OP_422J2_124_3477_n2637), .CI(DP_OP_422J2_124_3477_n2593), .CO(
        DP_OP_422J2_124_3477_n845), .S(DP_OP_422J2_124_3477_n846) );
  FADDX1_HVT DP_OP_422J2_124_3477_U518 ( .A(DP_OP_422J2_124_3477_n2329), .B(
        DP_OP_422J2_124_3477_n1846), .CI(DP_OP_422J2_124_3477_n2285), .CO(
        DP_OP_422J2_124_3477_n843), .S(DP_OP_422J2_124_3477_n844) );
  FADDX1_HVT DP_OP_422J2_124_3477_U517 ( .A(DP_OP_422J2_124_3477_n2197), .B(
        DP_OP_422J2_124_3477_n2549), .CI(DP_OP_422J2_124_3477_n2065), .CO(
        DP_OP_422J2_124_3477_n841), .S(DP_OP_422J2_124_3477_n842) );
  FADDX1_HVT DP_OP_422J2_124_3477_U516 ( .A(DP_OP_422J2_124_3477_n2396), .B(
        DP_OP_422J2_124_3477_n2241), .CI(DP_OP_422J2_124_3477_n2373), .CO(
        DP_OP_422J2_124_3477_n839), .S(DP_OP_422J2_124_3477_n840) );
  FADDX1_HVT DP_OP_422J2_124_3477_U515 ( .A(DP_OP_422J2_124_3477_n2841), .B(
        DP_OP_422J2_124_3477_n1934), .CI(DP_OP_422J2_124_3477_n2271), .CO(
        DP_OP_422J2_124_3477_n837), .S(DP_OP_422J2_124_3477_n838) );
  FADDX1_HVT DP_OP_422J2_124_3477_U514 ( .A(DP_OP_422J2_124_3477_n2885), .B(
        DP_OP_422J2_124_3477_n2535), .CI(DP_OP_422J2_124_3477_n2139), .CO(
        DP_OP_422J2_124_3477_n835), .S(DP_OP_422J2_124_3477_n836) );
  FADDX1_HVT DP_OP_422J2_124_3477_U513 ( .A(DP_OP_422J2_124_3477_n2322), .B(
        DP_OP_422J2_124_3477_n2410), .CI(DP_OP_422J2_124_3477_n2899), .CO(
        DP_OP_422J2_124_3477_n833), .S(DP_OP_422J2_124_3477_n834) );
  FADDX1_HVT DP_OP_422J2_124_3477_U512 ( .A(DP_OP_422J2_124_3477_n2058), .B(
        DP_OP_422J2_124_3477_n1964), .CI(DP_OP_422J2_124_3477_n2579), .CO(
        DP_OP_422J2_124_3477_n831), .S(DP_OP_422J2_124_3477_n832) );
  FADDX1_HVT DP_OP_422J2_124_3477_U511 ( .A(DP_OP_422J2_124_3477_n2586), .B(
        DP_OP_422J2_124_3477_n2146), .CI(DP_OP_422J2_124_3477_n2153), .CO(
        DP_OP_422J2_124_3477_n829), .S(DP_OP_422J2_124_3477_n830) );
  FADDX1_HVT DP_OP_422J2_124_3477_U510 ( .A(DP_OP_422J2_124_3477_n1839), .B(
        DP_OP_422J2_124_3477_n2220), .CI(DP_OP_422J2_124_3477_n2227), .CO(
        DP_OP_422J2_124_3477_n827), .S(DP_OP_422J2_124_3477_n828) );
  FADDX1_HVT DP_OP_422J2_124_3477_U509 ( .A(DP_OP_422J2_124_3477_n2630), .B(
        DP_OP_422J2_124_3477_n1781), .CI(DP_OP_422J2_124_3477_n2447), .CO(
        DP_OP_422J2_124_3477_n825), .S(DP_OP_422J2_124_3477_n826) );
  FADDX1_HVT DP_OP_422J2_124_3477_U508 ( .A(DP_OP_422J2_124_3477_n2753), .B(
        DP_OP_422J2_124_3477_n2498), .CI(DP_OP_422J2_124_3477_n2095), .CO(
        DP_OP_422J2_124_3477_n823), .S(DP_OP_422J2_124_3477_n824) );
  FADDX1_HVT DP_OP_422J2_124_3477_U507 ( .A(DP_OP_422J2_124_3477_n1883), .B(
        DP_OP_422J2_124_3477_n2051), .CI(DP_OP_422J2_124_3477_n1920), .CO(
        DP_OP_422J2_124_3477_n821), .S(DP_OP_422J2_124_3477_n822) );
  FADDX1_HVT DP_OP_422J2_124_3477_U506 ( .A(DP_OP_422J2_124_3477_n2491), .B(
        DP_OP_422J2_124_3477_n2315), .CI(DP_OP_422J2_124_3477_n2183), .CO(
        DP_OP_422J2_124_3477_n819), .S(DP_OP_422J2_124_3477_n820) );
  FADDX1_HVT DP_OP_422J2_124_3477_U505 ( .A(DP_OP_422J2_124_3477_n2102), .B(
        DP_OP_422J2_124_3477_n2667), .CI(DP_OP_422J2_124_3477_n1832), .CO(
        DP_OP_422J2_124_3477_n817), .S(DP_OP_422J2_124_3477_n818) );
  FADDX1_HVT DP_OP_422J2_124_3477_U504 ( .A(DP_OP_422J2_124_3477_n2359), .B(
        DP_OP_422J2_124_3477_n2848), .CI(DP_OP_422J2_124_3477_n2234), .CO(
        DP_OP_422J2_124_3477_n815), .S(DP_OP_422J2_124_3477_n816) );
  FADDX1_HVT DP_OP_422J2_124_3477_U503 ( .A(DP_OP_422J2_124_3477_n2674), .B(
        DP_OP_422J2_124_3477_n2542), .CI(DP_OP_422J2_124_3477_n2190), .CO(
        DP_OP_422J2_124_3477_n813), .S(DP_OP_422J2_124_3477_n814) );
  FADDX1_HVT DP_OP_422J2_124_3477_U502 ( .A(DP_OP_422J2_124_3477_n2811), .B(
        DP_OP_422J2_124_3477_n2892), .CI(DP_OP_422J2_124_3477_n2007), .CO(
        DP_OP_422J2_124_3477_n811), .S(DP_OP_422J2_124_3477_n812) );
  FADDX1_HVT DP_OP_422J2_124_3477_U501 ( .A(DP_OP_422J2_124_3477_n2454), .B(
        DP_OP_422J2_124_3477_n2278), .CI(DP_OP_422J2_124_3477_n2366), .CO(
        DP_OP_422J2_124_3477_n809), .S(DP_OP_422J2_124_3477_n810) );
  FADDX1_HVT DP_OP_422J2_124_3477_U500 ( .A(DP_OP_422J2_124_3477_n2709), .B(
        DP_OP_422J2_124_3477_n2760), .CI(DP_OP_422J2_124_3477_n2623), .CO(
        DP_OP_422J2_124_3477_n807), .S(DP_OP_422J2_124_3477_n808) );
  FADDX1_HVT DP_OP_422J2_124_3477_U499 ( .A(DP_OP_422J2_124_3477_n2804), .B(
        DP_OP_422J2_124_3477_n1061), .CI(DP_OP_422J2_124_3477_n2797), .CO(
        DP_OP_422J2_124_3477_n805), .S(DP_OP_422J2_124_3477_n806) );
  FADDX1_HVT DP_OP_422J2_124_3477_U498 ( .A(DP_OP_422J2_124_3477_n2014), .B(
        DP_OP_422J2_124_3477_n2716), .CI(DP_OP_422J2_124_3477_n1971), .CO(
        DP_OP_422J2_124_3477_n803), .S(DP_OP_422J2_124_3477_n804) );
  FADDX1_HVT DP_OP_422J2_124_3477_U497 ( .A(DP_OP_422J2_124_3477_n2403), .B(
        DP_OP_422J2_124_3477_n1927), .CI(DP_OP_422J2_124_3477_n1876), .CO(
        DP_OP_422J2_124_3477_n801), .S(DP_OP_422J2_124_3477_n802) );
  FADDX1_HVT DP_OP_422J2_124_3477_U496 ( .A(DP_OP_422J2_124_3477_n1051), .B(
        DP_OP_422J2_124_3477_n1059), .CI(DP_OP_422J2_124_3477_n1057), .CO(
        DP_OP_422J2_124_3477_n799), .S(DP_OP_422J2_124_3477_n800) );
  FADDX1_HVT DP_OP_422J2_124_3477_U495 ( .A(DP_OP_422J2_124_3477_n1053), .B(
        DP_OP_422J2_124_3477_n1047), .CI(DP_OP_422J2_124_3477_n1055), .CO(
        DP_OP_422J2_124_3477_n797), .S(DP_OP_422J2_124_3477_n798) );
  FADDX1_HVT DP_OP_422J2_124_3477_U494 ( .A(DP_OP_422J2_124_3477_n1049), .B(
        DP_OP_422J2_124_3477_n1045), .CI(DP_OP_422J2_124_3477_n1025), .CO(
        DP_OP_422J2_124_3477_n795), .S(DP_OP_422J2_124_3477_n796) );
  FADDX1_HVT DP_OP_422J2_124_3477_U493 ( .A(DP_OP_422J2_124_3477_n1043), .B(
        DP_OP_422J2_124_3477_n1019), .CI(DP_OP_422J2_124_3477_n1021), .CO(
        DP_OP_422J2_124_3477_n793), .S(DP_OP_422J2_124_3477_n794) );
  FADDX1_HVT DP_OP_422J2_124_3477_U492 ( .A(DP_OP_422J2_124_3477_n1041), .B(
        DP_OP_422J2_124_3477_n1023), .CI(DP_OP_422J2_124_3477_n1027), .CO(
        DP_OP_422J2_124_3477_n791), .S(DP_OP_422J2_124_3477_n792) );
  FADDX1_HVT DP_OP_422J2_124_3477_U491 ( .A(DP_OP_422J2_124_3477_n1033), .B(
        DP_OP_422J2_124_3477_n1029), .CI(DP_OP_422J2_124_3477_n1031), .CO(
        DP_OP_422J2_124_3477_n789), .S(DP_OP_422J2_124_3477_n790) );
  FADDX1_HVT DP_OP_422J2_124_3477_U490 ( .A(DP_OP_422J2_124_3477_n1039), .B(
        DP_OP_422J2_124_3477_n1037), .CI(DP_OP_422J2_124_3477_n1035), .CO(
        DP_OP_422J2_124_3477_n787), .S(DP_OP_422J2_124_3477_n788) );
  FADDX1_HVT DP_OP_422J2_124_3477_U489 ( .A(DP_OP_422J2_124_3477_n1015), .B(
        DP_OP_422J2_124_3477_n848), .CI(DP_OP_422J2_124_3477_n995), .CO(
        DP_OP_422J2_124_3477_n785), .S(DP_OP_422J2_124_3477_n786) );
  FADDX1_HVT DP_OP_422J2_124_3477_U488 ( .A(DP_OP_422J2_124_3477_n1017), .B(
        DP_OP_422J2_124_3477_n850), .CI(DP_OP_422J2_124_3477_n999), .CO(
        DP_OP_422J2_124_3477_n783), .S(DP_OP_422J2_124_3477_n784) );
  FADDX1_HVT DP_OP_422J2_124_3477_U487 ( .A(DP_OP_422J2_124_3477_n1013), .B(
        DP_OP_422J2_124_3477_n846), .CI(DP_OP_422J2_124_3477_n997), .CO(
        DP_OP_422J2_124_3477_n781), .S(DP_OP_422J2_124_3477_n782) );
  FADDX1_HVT DP_OP_422J2_124_3477_U486 ( .A(DP_OP_422J2_124_3477_n1011), .B(
        DP_OP_422J2_124_3477_n860), .CI(DP_OP_422J2_124_3477_n844), .CO(
        DP_OP_422J2_124_3477_n779), .S(DP_OP_422J2_124_3477_n780) );
  FADDX1_HVT DP_OP_422J2_124_3477_U485 ( .A(DP_OP_422J2_124_3477_n1009), .B(
        DP_OP_422J2_124_3477_n862), .CI(DP_OP_422J2_124_3477_n842), .CO(
        DP_OP_422J2_124_3477_n777), .S(DP_OP_422J2_124_3477_n778) );
  FADDX1_HVT DP_OP_422J2_124_3477_U484 ( .A(DP_OP_422J2_124_3477_n1007), .B(
        DP_OP_422J2_124_3477_n864), .CI(DP_OP_422J2_124_3477_n852), .CO(
        DP_OP_422J2_124_3477_n775), .S(DP_OP_422J2_124_3477_n776) );
  FADDX1_HVT DP_OP_422J2_124_3477_U483 ( .A(DP_OP_422J2_124_3477_n1005), .B(
        DP_OP_422J2_124_3477_n854), .CI(DP_OP_422J2_124_3477_n858), .CO(
        DP_OP_422J2_124_3477_n773), .S(DP_OP_422J2_124_3477_n774) );
  FADDX1_HVT DP_OP_422J2_124_3477_U482 ( .A(DP_OP_422J2_124_3477_n1003), .B(
        DP_OP_422J2_124_3477_n868), .CI(DP_OP_422J2_124_3477_n856), .CO(
        DP_OP_422J2_124_3477_n771), .S(DP_OP_422J2_124_3477_n772) );
  FADDX1_HVT DP_OP_422J2_124_3477_U481 ( .A(DP_OP_422J2_124_3477_n1001), .B(
        DP_OP_422J2_124_3477_n866), .CI(DP_OP_422J2_124_3477_n840), .CO(
        DP_OP_422J2_124_3477_n769), .S(DP_OP_422J2_124_3477_n770) );
  FADDX1_HVT DP_OP_422J2_124_3477_U480 ( .A(DP_OP_422J2_124_3477_n836), .B(
        DP_OP_422J2_124_3477_n828), .CI(DP_OP_422J2_124_3477_n824), .CO(
        DP_OP_422J2_124_3477_n767), .S(DP_OP_422J2_124_3477_n768) );
  FADDX1_HVT DP_OP_422J2_124_3477_U479 ( .A(DP_OP_422J2_124_3477_n838), .B(
        DP_OP_422J2_124_3477_n832), .CI(DP_OP_422J2_124_3477_n834), .CO(
        DP_OP_422J2_124_3477_n765), .S(DP_OP_422J2_124_3477_n766) );
  FADDX1_HVT DP_OP_422J2_124_3477_U478 ( .A(DP_OP_422J2_124_3477_n826), .B(
        DP_OP_422J2_124_3477_n830), .CI(DP_OP_422J2_124_3477_n820), .CO(
        DP_OP_422J2_124_3477_n763), .S(DP_OP_422J2_124_3477_n764) );
  FADDX1_HVT DP_OP_422J2_124_3477_U477 ( .A(DP_OP_422J2_124_3477_n818), .B(
        DP_OP_422J2_124_3477_n808), .CI(DP_OP_422J2_124_3477_n802), .CO(
        DP_OP_422J2_124_3477_n761), .S(DP_OP_422J2_124_3477_n762) );
  FADDX1_HVT DP_OP_422J2_124_3477_U476 ( .A(DP_OP_422J2_124_3477_n822), .B(
        DP_OP_422J2_124_3477_n810), .CI(DP_OP_422J2_124_3477_n804), .CO(
        DP_OP_422J2_124_3477_n759), .S(DP_OP_422J2_124_3477_n760) );
  FADDX1_HVT DP_OP_422J2_124_3477_U475 ( .A(DP_OP_422J2_124_3477_n816), .B(
        DP_OP_422J2_124_3477_n812), .CI(DP_OP_422J2_124_3477_n806), .CO(
        DP_OP_422J2_124_3477_n757), .S(DP_OP_422J2_124_3477_n758) );
  FADDX1_HVT DP_OP_422J2_124_3477_U474 ( .A(DP_OP_422J2_124_3477_n814), .B(
        DP_OP_422J2_124_3477_n993), .CI(DP_OP_422J2_124_3477_n991), .CO(
        DP_OP_422J2_124_3477_n755), .S(DP_OP_422J2_124_3477_n756) );
  FADDX1_HVT DP_OP_422J2_124_3477_U473 ( .A(DP_OP_422J2_124_3477_n989), .B(
        DP_OP_422J2_124_3477_n987), .CI(DP_OP_422J2_124_3477_n985), .CO(
        DP_OP_422J2_124_3477_n753), .S(DP_OP_422J2_124_3477_n754) );
  FADDX1_HVT DP_OP_422J2_124_3477_U472 ( .A(DP_OP_422J2_124_3477_n983), .B(
        DP_OP_422J2_124_3477_n979), .CI(DP_OP_422J2_124_3477_n981), .CO(
        DP_OP_422J2_124_3477_n751), .S(DP_OP_422J2_124_3477_n752) );
  FADDX1_HVT DP_OP_422J2_124_3477_U471 ( .A(DP_OP_422J2_124_3477_n977), .B(
        DP_OP_422J2_124_3477_n798), .CI(DP_OP_422J2_124_3477_n800), .CO(
        DP_OP_422J2_124_3477_n749), .S(DP_OP_422J2_124_3477_n750) );
  FADDX1_HVT DP_OP_422J2_124_3477_U470 ( .A(DP_OP_422J2_124_3477_n975), .B(
        DP_OP_422J2_124_3477_n969), .CI(DP_OP_422J2_124_3477_n967), .CO(
        DP_OP_422J2_124_3477_n747), .S(DP_OP_422J2_124_3477_n748) );
  FADDX1_HVT DP_OP_422J2_124_3477_U469 ( .A(DP_OP_422J2_124_3477_n973), .B(
        DP_OP_422J2_124_3477_n971), .CI(DP_OP_422J2_124_3477_n796), .CO(
        DP_OP_422J2_124_3477_n745), .S(DP_OP_422J2_124_3477_n746) );
  FADDX1_HVT DP_OP_422J2_124_3477_U468 ( .A(DP_OP_422J2_124_3477_n965), .B(
        DP_OP_422J2_124_3477_n792), .CI(DP_OP_422J2_124_3477_n790), .CO(
        DP_OP_422J2_124_3477_n743), .S(DP_OP_422J2_124_3477_n744) );
  FADDX1_HVT DP_OP_422J2_124_3477_U467 ( .A(DP_OP_422J2_124_3477_n959), .B(
        DP_OP_422J2_124_3477_n788), .CI(DP_OP_422J2_124_3477_n794), .CO(
        DP_OP_422J2_124_3477_n741), .S(DP_OP_422J2_124_3477_n742) );
  FADDX1_HVT DP_OP_422J2_124_3477_U466 ( .A(DP_OP_422J2_124_3477_n963), .B(
        DP_OP_422J2_124_3477_n957), .CI(DP_OP_422J2_124_3477_n961), .CO(
        DP_OP_422J2_124_3477_n739), .S(DP_OP_422J2_124_3477_n740) );
  FADDX1_HVT DP_OP_422J2_124_3477_U465 ( .A(DP_OP_422J2_124_3477_n955), .B(
        DP_OP_422J2_124_3477_n774), .CI(DP_OP_422J2_124_3477_n770), .CO(
        DP_OP_422J2_124_3477_n737), .S(DP_OP_422J2_124_3477_n738) );
  FADDX1_HVT DP_OP_422J2_124_3477_U464 ( .A(DP_OP_422J2_124_3477_n784), .B(
        DP_OP_422J2_124_3477_n776), .CI(DP_OP_422J2_124_3477_n772), .CO(
        DP_OP_422J2_124_3477_n735), .S(DP_OP_422J2_124_3477_n736) );
  FADDX1_HVT DP_OP_422J2_124_3477_U463 ( .A(DP_OP_422J2_124_3477_n786), .B(
        DP_OP_422J2_124_3477_n949), .CI(DP_OP_422J2_124_3477_n778), .CO(
        DP_OP_422J2_124_3477_n733), .S(DP_OP_422J2_124_3477_n734) );
  FADDX1_HVT DP_OP_422J2_124_3477_U462 ( .A(DP_OP_422J2_124_3477_n953), .B(
        DP_OP_422J2_124_3477_n951), .CI(DP_OP_422J2_124_3477_n780), .CO(
        DP_OP_422J2_124_3477_n731), .S(DP_OP_422J2_124_3477_n732) );
  FADDX1_HVT DP_OP_422J2_124_3477_U461 ( .A(DP_OP_422J2_124_3477_n782), .B(
        DP_OP_422J2_124_3477_n766), .CI(DP_OP_422J2_124_3477_n768), .CO(
        DP_OP_422J2_124_3477_n729), .S(DP_OP_422J2_124_3477_n730) );
  FADDX1_HVT DP_OP_422J2_124_3477_U460 ( .A(DP_OP_422J2_124_3477_n947), .B(
        DP_OP_422J2_124_3477_n764), .CI(DP_OP_422J2_124_3477_n760), .CO(
        DP_OP_422J2_124_3477_n727), .S(DP_OP_422J2_124_3477_n728) );
  FADDX1_HVT DP_OP_422J2_124_3477_U459 ( .A(DP_OP_422J2_124_3477_n762), .B(
        DP_OP_422J2_124_3477_n945), .CI(DP_OP_422J2_124_3477_n756), .CO(
        DP_OP_422J2_124_3477_n725), .S(DP_OP_422J2_124_3477_n726) );
  FADDX1_HVT DP_OP_422J2_124_3477_U458 ( .A(DP_OP_422J2_124_3477_n758), .B(
        DP_OP_422J2_124_3477_n943), .CI(DP_OP_422J2_124_3477_n941), .CO(
        DP_OP_422J2_124_3477_n723), .S(DP_OP_422J2_124_3477_n724) );
  FADDX1_HVT DP_OP_422J2_124_3477_U457 ( .A(DP_OP_422J2_124_3477_n939), .B(
        DP_OP_422J2_124_3477_n937), .CI(DP_OP_422J2_124_3477_n754), .CO(
        DP_OP_422J2_124_3477_n721), .S(DP_OP_422J2_124_3477_n722) );
  FADDX1_HVT DP_OP_422J2_124_3477_U456 ( .A(DP_OP_422J2_124_3477_n935), .B(
        DP_OP_422J2_124_3477_n931), .CI(DP_OP_422J2_124_3477_n752), .CO(
        DP_OP_422J2_124_3477_n719), .S(DP_OP_422J2_124_3477_n720) );
  FADDX1_HVT DP_OP_422J2_124_3477_U455 ( .A(DP_OP_422J2_124_3477_n933), .B(
        DP_OP_422J2_124_3477_n929), .CI(DP_OP_422J2_124_3477_n750), .CO(
        DP_OP_422J2_124_3477_n717), .S(DP_OP_422J2_124_3477_n718) );
  FADDX1_HVT DP_OP_422J2_124_3477_U454 ( .A(DP_OP_422J2_124_3477_n927), .B(
        DP_OP_422J2_124_3477_n925), .CI(DP_OP_422J2_124_3477_n746), .CO(
        DP_OP_422J2_124_3477_n715), .S(DP_OP_422J2_124_3477_n716) );
  FADDX1_HVT DP_OP_422J2_124_3477_U453 ( .A(DP_OP_422J2_124_3477_n748), .B(
        DP_OP_422J2_124_3477_n923), .CI(DP_OP_422J2_124_3477_n744), .CO(
        DP_OP_422J2_124_3477_n713), .S(DP_OP_422J2_124_3477_n714) );
  FADDX1_HVT DP_OP_422J2_124_3477_U452 ( .A(DP_OP_422J2_124_3477_n921), .B(
        DP_OP_422J2_124_3477_n740), .CI(DP_OP_422J2_124_3477_n742), .CO(
        DP_OP_422J2_124_3477_n711), .S(DP_OP_422J2_124_3477_n712) );
  FADDX1_HVT DP_OP_422J2_124_3477_U451 ( .A(DP_OP_422J2_124_3477_n919), .B(
        DP_OP_422J2_124_3477_n917), .CI(DP_OP_422J2_124_3477_n732), .CO(
        DP_OP_422J2_124_3477_n709), .S(DP_OP_422J2_124_3477_n710) );
  FADDX1_HVT DP_OP_422J2_124_3477_U450 ( .A(DP_OP_422J2_124_3477_n736), .B(
        DP_OP_422J2_124_3477_n734), .CI(DP_OP_422J2_124_3477_n738), .CO(
        DP_OP_422J2_124_3477_n707), .S(DP_OP_422J2_124_3477_n708) );
  FADDX1_HVT DP_OP_422J2_124_3477_U449 ( .A(DP_OP_422J2_124_3477_n730), .B(
        DP_OP_422J2_124_3477_n915), .CI(DP_OP_422J2_124_3477_n728), .CO(
        DP_OP_422J2_124_3477_n705), .S(DP_OP_422J2_124_3477_n706) );
  FADDX1_HVT DP_OP_422J2_124_3477_U448 ( .A(DP_OP_422J2_124_3477_n913), .B(
        DP_OP_422J2_124_3477_n726), .CI(DP_OP_422J2_124_3477_n724), .CO(
        DP_OP_422J2_124_3477_n703), .S(DP_OP_422J2_124_3477_n704) );
  FADDX1_HVT DP_OP_422J2_124_3477_U447 ( .A(DP_OP_422J2_124_3477_n911), .B(
        DP_OP_422J2_124_3477_n909), .CI(DP_OP_422J2_124_3477_n907), .CO(
        DP_OP_422J2_124_3477_n701), .S(DP_OP_422J2_124_3477_n702) );
  FADDX1_HVT DP_OP_422J2_124_3477_U446 ( .A(DP_OP_422J2_124_3477_n722), .B(
        DP_OP_422J2_124_3477_n905), .CI(DP_OP_422J2_124_3477_n720), .CO(
        DP_OP_422J2_124_3477_n699), .S(DP_OP_422J2_124_3477_n700) );
  FADDX1_HVT DP_OP_422J2_124_3477_U445 ( .A(DP_OP_422J2_124_3477_n903), .B(
        DP_OP_422J2_124_3477_n718), .CI(DP_OP_422J2_124_3477_n901), .CO(
        DP_OP_422J2_124_3477_n697), .S(DP_OP_422J2_124_3477_n698) );
  FADDX1_HVT DP_OP_422J2_124_3477_U444 ( .A(DP_OP_422J2_124_3477_n716), .B(
        DP_OP_422J2_124_3477_n899), .CI(DP_OP_422J2_124_3477_n714), .CO(
        DP_OP_422J2_124_3477_n695), .S(DP_OP_422J2_124_3477_n696) );
  FADDX1_HVT DP_OP_422J2_124_3477_U443 ( .A(DP_OP_422J2_124_3477_n712), .B(
        DP_OP_422J2_124_3477_n897), .CI(DP_OP_422J2_124_3477_n710), .CO(
        DP_OP_422J2_124_3477_n693), .S(DP_OP_422J2_124_3477_n694) );
  FADDX1_HVT DP_OP_422J2_124_3477_U442 ( .A(DP_OP_422J2_124_3477_n708), .B(
        DP_OP_422J2_124_3477_n895), .CI(DP_OP_422J2_124_3477_n706), .CO(
        DP_OP_422J2_124_3477_n691), .S(DP_OP_422J2_124_3477_n692) );
  FADDX1_HVT DP_OP_422J2_124_3477_U441 ( .A(DP_OP_422J2_124_3477_n893), .B(
        DP_OP_422J2_124_3477_n704), .CI(DP_OP_422J2_124_3477_n891), .CO(
        DP_OP_422J2_124_3477_n689), .S(DP_OP_422J2_124_3477_n690) );
  FADDX1_HVT DP_OP_422J2_124_3477_U440 ( .A(DP_OP_422J2_124_3477_n702), .B(
        DP_OP_422J2_124_3477_n889), .CI(DP_OP_422J2_124_3477_n700), .CO(
        DP_OP_422J2_124_3477_n687), .S(DP_OP_422J2_124_3477_n688) );
  FADDX1_HVT DP_OP_422J2_124_3477_U439 ( .A(DP_OP_422J2_124_3477_n887), .B(
        DP_OP_422J2_124_3477_n698), .CI(DP_OP_422J2_124_3477_n885), .CO(
        DP_OP_422J2_124_3477_n685), .S(DP_OP_422J2_124_3477_n686) );
  FADDX1_HVT DP_OP_422J2_124_3477_U438 ( .A(DP_OP_422J2_124_3477_n696), .B(
        DP_OP_422J2_124_3477_n883), .CI(DP_OP_422J2_124_3477_n694), .CO(
        DP_OP_422J2_124_3477_n683), .S(DP_OP_422J2_124_3477_n684) );
  FADDX1_HVT DP_OP_422J2_124_3477_U437 ( .A(DP_OP_422J2_124_3477_n692), .B(
        DP_OP_422J2_124_3477_n881), .CI(DP_OP_422J2_124_3477_n690), .CO(
        DP_OP_422J2_124_3477_n681), .S(DP_OP_422J2_124_3477_n682) );
  FADDX1_HVT DP_OP_422J2_124_3477_U436 ( .A(DP_OP_422J2_124_3477_n879), .B(
        DP_OP_422J2_124_3477_n688), .CI(DP_OP_422J2_124_3477_n877), .CO(
        DP_OP_422J2_124_3477_n679), .S(DP_OP_422J2_124_3477_n680) );
  FADDX1_HVT DP_OP_422J2_124_3477_U435 ( .A(DP_OP_422J2_124_3477_n686), .B(
        DP_OP_422J2_124_3477_n875), .CI(DP_OP_422J2_124_3477_n684), .CO(
        DP_OP_422J2_124_3477_n677), .S(DP_OP_422J2_124_3477_n678) );
  FADDX1_HVT DP_OP_422J2_124_3477_U434 ( .A(DP_OP_422J2_124_3477_n682), .B(
        DP_OP_422J2_124_3477_n873), .CI(DP_OP_422J2_124_3477_n680), .CO(
        DP_OP_422J2_124_3477_n675), .S(DP_OP_422J2_124_3477_n676) );
  FADDX1_HVT DP_OP_422J2_124_3477_U433 ( .A(DP_OP_422J2_124_3477_n871), .B(
        DP_OP_422J2_124_3477_n678), .CI(DP_OP_422J2_124_3477_n676), .CO(
        DP_OP_422J2_124_3477_n673), .S(DP_OP_422J2_124_3477_n674) );
  FADDX1_HVT DP_OP_422J2_124_3477_U431 ( .A(DP_OP_422J2_124_3477_n2000), .B(
        DP_OP_422J2_124_3477_n2145), .CI(DP_OP_422J2_124_3477_n1956), .CO(
        DP_OP_422J2_124_3477_n669), .S(DP_OP_422J2_124_3477_n670) );
  FADDX1_HVT DP_OP_422J2_124_3477_U430 ( .A(DP_OP_422J2_124_3477_n2351), .B(
        DP_OP_422J2_124_3477_n2409), .CI(DP_OP_422J2_124_3477_n2745), .CO(
        DP_OP_422J2_124_3477_n667), .S(DP_OP_422J2_124_3477_n668) );
  FADDX1_HVT DP_OP_422J2_124_3477_U429 ( .A(DP_OP_422J2_124_3477_n2307), .B(
        DP_OP_422J2_124_3477_n2571), .CI(DP_OP_422J2_124_3477_n1824), .CO(
        DP_OP_422J2_124_3477_n665), .S(DP_OP_422J2_124_3477_n666) );
  FADDX1_HVT DP_OP_422J2_124_3477_U428 ( .A(DP_OP_422J2_124_3477_n2131), .B(
        DP_OP_422J2_124_3477_n2175), .CI(DP_OP_422J2_124_3477_n2043), .CO(
        DP_OP_422J2_124_3477_n663), .S(DP_OP_422J2_124_3477_n664) );
  FADDX1_HVT DP_OP_422J2_124_3477_U427 ( .A(DP_OP_422J2_124_3477_n2087), .B(
        DP_OP_422J2_124_3477_n2439), .CI(DP_OP_422J2_124_3477_n2483), .CO(
        DP_OP_422J2_124_3477_n661), .S(DP_OP_422J2_124_3477_n662) );
  FADDX1_HVT DP_OP_422J2_124_3477_U426 ( .A(DP_OP_422J2_124_3477_n2789), .B(
        DP_OP_422J2_124_3477_n2527), .CI(DP_OP_422J2_124_3477_n1912), .CO(
        DP_OP_422J2_124_3477_n659), .S(DP_OP_422J2_124_3477_n660) );
  FADDX1_HVT DP_OP_422J2_124_3477_U425 ( .A(DP_OP_422J2_124_3477_n1868), .B(
        DP_OP_422J2_124_3477_n2057), .CI(DP_OP_422J2_124_3477_n2877), .CO(
        DP_OP_422J2_124_3477_n657), .S(DP_OP_422J2_124_3477_n658) );
  FADDX1_HVT DP_OP_422J2_124_3477_U424 ( .A(DP_OP_422J2_124_3477_n2615), .B(
        DP_OP_422J2_124_3477_n2497), .CI(DP_OP_422J2_124_3477_n2629), .CO(
        DP_OP_422J2_124_3477_n655), .S(DP_OP_422J2_124_3477_n656) );
  FADDX1_HVT DP_OP_422J2_124_3477_U423 ( .A(DP_OP_422J2_124_3477_n2659), .B(
        DP_OP_422J2_124_3477_n2321), .CI(DP_OP_422J2_124_3477_n1838), .CO(
        DP_OP_422J2_124_3477_n653), .S(DP_OP_422J2_124_3477_n654) );
  FADDX1_HVT DP_OP_422J2_124_3477_U422 ( .A(DP_OP_422J2_124_3477_n2833), .B(
        DP_OP_422J2_124_3477_n2263), .CI(DP_OP_422J2_124_3477_n2585), .CO(
        DP_OP_422J2_124_3477_n651), .S(DP_OP_422J2_124_3477_n652) );
  FADDX1_HVT DP_OP_422J2_124_3477_U421 ( .A(DP_OP_422J2_124_3477_n2395), .B(
        DP_OP_422J2_124_3477_n2534), .CI(DP_OP_422J2_124_3477_n2715), .CO(
        DP_OP_422J2_124_3477_n649), .S(DP_OP_422J2_124_3477_n650) );
  FADDX1_HVT DP_OP_422J2_124_3477_U420 ( .A(DP_OP_422J2_124_3477_n2840), .B(
        DP_OP_422J2_124_3477_n2541), .CI(DP_OP_422J2_124_3477_n2138), .CO(
        DP_OP_422J2_124_3477_n647), .S(DP_OP_422J2_124_3477_n648) );
  FADDX1_HVT DP_OP_422J2_124_3477_U419 ( .A(DP_OP_422J2_124_3477_n2884), .B(
        DP_OP_422J2_124_3477_n2453), .CI(DP_OP_422J2_124_3477_n2270), .CO(
        DP_OP_422J2_124_3477_n645), .S(DP_OP_422J2_124_3477_n646) );
  FADDX1_HVT DP_OP_422J2_124_3477_U418 ( .A(DP_OP_422J2_124_3477_n2752), .B(
        DP_OP_422J2_124_3477_n2847), .CI(DP_OP_422J2_124_3477_n2233), .CO(
        DP_OP_422J2_124_3477_n643), .S(DP_OP_422J2_124_3477_n644) );
  FADDX1_HVT DP_OP_422J2_124_3477_U417 ( .A(DP_OP_422J2_124_3477_n1780), .B(
        DP_OP_422J2_124_3477_n1963), .CI(DP_OP_422J2_124_3477_n2189), .CO(
        DP_OP_422J2_124_3477_n641), .S(DP_OP_422J2_124_3477_n642) );
  FADDX1_HVT DP_OP_422J2_124_3477_U416 ( .A(DP_OP_422J2_124_3477_n2219), .B(
        DP_OP_422J2_124_3477_n2673), .CI(DP_OP_422J2_124_3477_n2365), .CO(
        DP_OP_422J2_124_3477_n639), .S(DP_OP_422J2_124_3477_n640) );
  FADDX1_HVT DP_OP_422J2_124_3477_U415 ( .A(DP_OP_422J2_124_3477_n672), .B(
        DP_OP_422J2_124_3477_n2101), .CI(DP_OP_422J2_124_3477_n1970), .CO(
        DP_OP_422J2_124_3477_n637), .S(DP_OP_422J2_124_3477_n638) );
  FADDX1_HVT DP_OP_422J2_124_3477_U414 ( .A(DP_OP_422J2_124_3477_n1882), .B(
        DP_OP_422J2_124_3477_n2277), .CI(DP_OP_422J2_124_3477_n2578), .CO(
        DP_OP_422J2_124_3477_n635), .S(DP_OP_422J2_124_3477_n636) );
  FADDX1_HVT DP_OP_422J2_124_3477_U413 ( .A(DP_OP_422J2_124_3477_n2803), .B(
        DP_OP_422J2_124_3477_n1926), .CI(DP_OP_422J2_124_3477_n2314), .CO(
        DP_OP_422J2_124_3477_n633), .S(DP_OP_422J2_124_3477_n634) );
  FADDX1_HVT DP_OP_422J2_124_3477_U412 ( .A(DP_OP_422J2_124_3477_n2891), .B(
        DP_OP_422J2_124_3477_n2013), .CI(DP_OP_422J2_124_3477_n2050), .CO(
        DP_OP_422J2_124_3477_n631), .S(DP_OP_422J2_124_3477_n632) );
  FADDX1_HVT DP_OP_422J2_124_3477_U411 ( .A(DP_OP_422J2_124_3477_n2446), .B(
        DP_OP_422J2_124_3477_n2759), .CI(DP_OP_422J2_124_3477_n2666), .CO(
        DP_OP_422J2_124_3477_n629), .S(DP_OP_422J2_124_3477_n630) );
  FADDX1_HVT DP_OP_422J2_124_3477_U410 ( .A(DP_OP_422J2_124_3477_n2226), .B(
        DP_OP_422J2_124_3477_n2094), .CI(DP_OP_422J2_124_3477_n2708), .CO(
        DP_OP_422J2_124_3477_n627), .S(DP_OP_422J2_124_3477_n628) );
  FADDX1_HVT DP_OP_422J2_124_3477_U409 ( .A(DP_OP_422J2_124_3477_n2490), .B(
        DP_OP_422J2_124_3477_n2358), .CI(DP_OP_422J2_124_3477_n1919), .CO(
        DP_OP_422J2_124_3477_n625), .S(DP_OP_422J2_124_3477_n626) );
  FADDX1_HVT DP_OP_422J2_124_3477_U408 ( .A(DP_OP_422J2_124_3477_n2402), .B(
        DP_OP_422J2_124_3477_n1831), .CI(DP_OP_422J2_124_3477_n2182), .CO(
        DP_OP_422J2_124_3477_n623), .S(DP_OP_422J2_124_3477_n624) );
  FADDX1_HVT DP_OP_422J2_124_3477_U407 ( .A(DP_OP_422J2_124_3477_n1875), .B(
        DP_OP_422J2_124_3477_n2622), .CI(DP_OP_422J2_124_3477_n2006), .CO(
        DP_OP_422J2_124_3477_n621), .S(DP_OP_422J2_124_3477_n622) );
  FADDX1_HVT DP_OP_422J2_124_3477_U406 ( .A(DP_OP_422J2_124_3477_n2796), .B(
        DP_OP_422J2_124_3477_n867), .CI(DP_OP_422J2_124_3477_n865), .CO(
        DP_OP_422J2_124_3477_n619), .S(DP_OP_422J2_124_3477_n620) );
  FADDX1_HVT DP_OP_422J2_124_3477_U405 ( .A(DP_OP_422J2_124_3477_n863), .B(
        DP_OP_422J2_124_3477_n841), .CI(DP_OP_422J2_124_3477_n843), .CO(
        DP_OP_422J2_124_3477_n617), .S(DP_OP_422J2_124_3477_n618) );
  FADDX1_HVT DP_OP_422J2_124_3477_U404 ( .A(DP_OP_422J2_124_3477_n861), .B(
        DP_OP_422J2_124_3477_n847), .CI(DP_OP_422J2_124_3477_n845), .CO(
        DP_OP_422J2_124_3477_n615), .S(DP_OP_422J2_124_3477_n616) );
  FADDX1_HVT DP_OP_422J2_124_3477_U403 ( .A(DP_OP_422J2_124_3477_n859), .B(
        DP_OP_422J2_124_3477_n849), .CI(DP_OP_422J2_124_3477_n851), .CO(
        DP_OP_422J2_124_3477_n613), .S(DP_OP_422J2_124_3477_n614) );
  FADDX1_HVT DP_OP_422J2_124_3477_U402 ( .A(DP_OP_422J2_124_3477_n857), .B(
        DP_OP_422J2_124_3477_n853), .CI(DP_OP_422J2_124_3477_n855), .CO(
        DP_OP_422J2_124_3477_n611), .S(DP_OP_422J2_124_3477_n612) );
  FADDX1_HVT DP_OP_422J2_124_3477_U401 ( .A(DP_OP_422J2_124_3477_n839), .B(
        DP_OP_422J2_124_3477_n823), .CI(DP_OP_422J2_124_3477_n825), .CO(
        DP_OP_422J2_124_3477_n609), .S(DP_OP_422J2_124_3477_n610) );
  FADDX1_HVT DP_OP_422J2_124_3477_U400 ( .A(DP_OP_422J2_124_3477_n837), .B(
        DP_OP_422J2_124_3477_n827), .CI(DP_OP_422J2_124_3477_n829), .CO(
        DP_OP_422J2_124_3477_n607), .S(DP_OP_422J2_124_3477_n608) );
  FADDX1_HVT DP_OP_422J2_124_3477_U399 ( .A(DP_OP_422J2_124_3477_n835), .B(
        DP_OP_422J2_124_3477_n831), .CI(DP_OP_422J2_124_3477_n833), .CO(
        DP_OP_422J2_124_3477_n605), .S(DP_OP_422J2_124_3477_n606) );
  FADDX1_HVT DP_OP_422J2_124_3477_U398 ( .A(DP_OP_422J2_124_3477_n821), .B(
        DP_OP_422J2_124_3477_n668), .CI(DP_OP_422J2_124_3477_n803), .CO(
        DP_OP_422J2_124_3477_n603), .S(DP_OP_422J2_124_3477_n604) );
  FADDX1_HVT DP_OP_422J2_124_3477_U397 ( .A(DP_OP_422J2_124_3477_n819), .B(
        DP_OP_422J2_124_3477_n656), .CI(DP_OP_422J2_124_3477_n801), .CO(
        DP_OP_422J2_124_3477_n601), .S(DP_OP_422J2_124_3477_n602) );
  FADDX1_HVT DP_OP_422J2_124_3477_U396 ( .A(DP_OP_422J2_124_3477_n817), .B(
        DP_OP_422J2_124_3477_n666), .CI(DP_OP_422J2_124_3477_n805), .CO(
        DP_OP_422J2_124_3477_n599), .S(DP_OP_422J2_124_3477_n600) );
  FADDX1_HVT DP_OP_422J2_124_3477_U395 ( .A(DP_OP_422J2_124_3477_n815), .B(
        DP_OP_422J2_124_3477_n660), .CI(DP_OP_422J2_124_3477_n652), .CO(
        DP_OP_422J2_124_3477_n597), .S(DP_OP_422J2_124_3477_n598) );
  FADDX1_HVT DP_OP_422J2_124_3477_U394 ( .A(DP_OP_422J2_124_3477_n813), .B(
        DP_OP_422J2_124_3477_n658), .CI(DP_OP_422J2_124_3477_n654), .CO(
        DP_OP_422J2_124_3477_n595), .S(DP_OP_422J2_124_3477_n596) );
  FADDX1_HVT DP_OP_422J2_124_3477_U393 ( .A(DP_OP_422J2_124_3477_n811), .B(
        DP_OP_422J2_124_3477_n662), .CI(DP_OP_422J2_124_3477_n664), .CO(
        DP_OP_422J2_124_3477_n593), .S(DP_OP_422J2_124_3477_n594) );
  FADDX1_HVT DP_OP_422J2_124_3477_U392 ( .A(DP_OP_422J2_124_3477_n809), .B(
        DP_OP_422J2_124_3477_n807), .CI(DP_OP_422J2_124_3477_n670), .CO(
        DP_OP_422J2_124_3477_n591), .S(DP_OP_422J2_124_3477_n592) );
  FADDX1_HVT DP_OP_422J2_124_3477_U391 ( .A(DP_OP_422J2_124_3477_n650), .B(
        DP_OP_422J2_124_3477_n636), .CI(DP_OP_422J2_124_3477_n630), .CO(
        DP_OP_422J2_124_3477_n589), .S(DP_OP_422J2_124_3477_n590) );
  FADDX1_HVT DP_OP_422J2_124_3477_U390 ( .A(DP_OP_422J2_124_3477_n646), .B(
        DP_OP_422J2_124_3477_n638), .CI(DP_OP_422J2_124_3477_n628), .CO(
        DP_OP_422J2_124_3477_n587), .S(DP_OP_422J2_124_3477_n588) );
  FADDX1_HVT DP_OP_422J2_124_3477_U389 ( .A(DP_OP_422J2_124_3477_n648), .B(
        DP_OP_422J2_124_3477_n640), .CI(DP_OP_422J2_124_3477_n632), .CO(
        DP_OP_422J2_124_3477_n585), .S(DP_OP_422J2_124_3477_n586) );
  FADDX1_HVT DP_OP_422J2_124_3477_U388 ( .A(DP_OP_422J2_124_3477_n644), .B(
        DP_OP_422J2_124_3477_n642), .CI(DP_OP_422J2_124_3477_n634), .CO(
        DP_OP_422J2_124_3477_n583), .S(DP_OP_422J2_124_3477_n584) );
  FADDX1_HVT DP_OP_422J2_124_3477_U387 ( .A(DP_OP_422J2_124_3477_n626), .B(
        DP_OP_422J2_124_3477_n624), .CI(DP_OP_422J2_124_3477_n622), .CO(
        DP_OP_422J2_124_3477_n581), .S(DP_OP_422J2_124_3477_n582) );
  FADDX1_HVT DP_OP_422J2_124_3477_U386 ( .A(DP_OP_422J2_124_3477_n799), .B(
        DP_OP_422J2_124_3477_n797), .CI(DP_OP_422J2_124_3477_n795), .CO(
        DP_OP_422J2_124_3477_n579), .S(DP_OP_422J2_124_3477_n580) );
  FADDX1_HVT DP_OP_422J2_124_3477_U385 ( .A(DP_OP_422J2_124_3477_n793), .B(
        DP_OP_422J2_124_3477_n787), .CI(DP_OP_422J2_124_3477_n789), .CO(
        DP_OP_422J2_124_3477_n577), .S(DP_OP_422J2_124_3477_n578) );
  FADDX1_HVT DP_OP_422J2_124_3477_U384 ( .A(DP_OP_422J2_124_3477_n791), .B(
        DP_OP_422J2_124_3477_n620), .CI(DP_OP_422J2_124_3477_n785), .CO(
        DP_OP_422J2_124_3477_n575), .S(DP_OP_422J2_124_3477_n576) );
  FADDX1_HVT DP_OP_422J2_124_3477_U383 ( .A(DP_OP_422J2_124_3477_n783), .B(
        DP_OP_422J2_124_3477_n612), .CI(DP_OP_422J2_124_3477_n618), .CO(
        DP_OP_422J2_124_3477_n573), .S(DP_OP_422J2_124_3477_n574) );
  FADDX1_HVT DP_OP_422J2_124_3477_U382 ( .A(DP_OP_422J2_124_3477_n781), .B(
        DP_OP_422J2_124_3477_n616), .CI(DP_OP_422J2_124_3477_n614), .CO(
        DP_OP_422J2_124_3477_n571), .S(DP_OP_422J2_124_3477_n572) );
  FADDX1_HVT DP_OP_422J2_124_3477_U381 ( .A(DP_OP_422J2_124_3477_n779), .B(
        DP_OP_422J2_124_3477_n771), .CI(DP_OP_422J2_124_3477_n769), .CO(
        DP_OP_422J2_124_3477_n569), .S(DP_OP_422J2_124_3477_n570) );
  FADDX1_HVT DP_OP_422J2_124_3477_U380 ( .A(DP_OP_422J2_124_3477_n777), .B(
        DP_OP_422J2_124_3477_n775), .CI(DP_OP_422J2_124_3477_n773), .CO(
        DP_OP_422J2_124_3477_n567), .S(DP_OP_422J2_124_3477_n568) );
  FADDX1_HVT DP_OP_422J2_124_3477_U379 ( .A(DP_OP_422J2_124_3477_n610), .B(
        DP_OP_422J2_124_3477_n767), .CI(DP_OP_422J2_124_3477_n763), .CO(
        DP_OP_422J2_124_3477_n565), .S(DP_OP_422J2_124_3477_n566) );
  FADDX1_HVT DP_OP_422J2_124_3477_U378 ( .A(DP_OP_422J2_124_3477_n606), .B(
        DP_OP_422J2_124_3477_n608), .CI(DP_OP_422J2_124_3477_n765), .CO(
        DP_OP_422J2_124_3477_n563), .S(DP_OP_422J2_124_3477_n564) );
  FADDX1_HVT DP_OP_422J2_124_3477_U377 ( .A(DP_OP_422J2_124_3477_n761), .B(
        DP_OP_422J2_124_3477_n592), .CI(DP_OP_422J2_124_3477_n755), .CO(
        DP_OP_422J2_124_3477_n561), .S(DP_OP_422J2_124_3477_n562) );
  FADDX1_HVT DP_OP_422J2_124_3477_U376 ( .A(DP_OP_422J2_124_3477_n759), .B(
        DP_OP_422J2_124_3477_n596), .CI(DP_OP_422J2_124_3477_n594), .CO(
        DP_OP_422J2_124_3477_n559), .S(DP_OP_422J2_124_3477_n560) );
  FADDX1_HVT DP_OP_422J2_124_3477_U375 ( .A(DP_OP_422J2_124_3477_n600), .B(
        DP_OP_422J2_124_3477_n757), .CI(DP_OP_422J2_124_3477_n598), .CO(
        DP_OP_422J2_124_3477_n557), .S(DP_OP_422J2_124_3477_n558) );
  FADDX1_HVT DP_OP_422J2_124_3477_U374 ( .A(DP_OP_422J2_124_3477_n602), .B(
        DP_OP_422J2_124_3477_n604), .CI(DP_OP_422J2_124_3477_n590), .CO(
        DP_OP_422J2_124_3477_n555), .S(DP_OP_422J2_124_3477_n556) );
  FADDX1_HVT DP_OP_422J2_124_3477_U373 ( .A(DP_OP_422J2_124_3477_n586), .B(
        DP_OP_422J2_124_3477_n584), .CI(DP_OP_422J2_124_3477_n753), .CO(
        DP_OP_422J2_124_3477_n553), .S(DP_OP_422J2_124_3477_n554) );
  FADDX1_HVT DP_OP_422J2_124_3477_U372 ( .A(DP_OP_422J2_124_3477_n588), .B(
        DP_OP_422J2_124_3477_n751), .CI(DP_OP_422J2_124_3477_n582), .CO(
        DP_OP_422J2_124_3477_n551), .S(DP_OP_422J2_124_3477_n552) );
  FADDX1_HVT DP_OP_422J2_124_3477_U371 ( .A(DP_OP_422J2_124_3477_n749), .B(
        DP_OP_422J2_124_3477_n745), .CI(DP_OP_422J2_124_3477_n580), .CO(
        DP_OP_422J2_124_3477_n549), .S(DP_OP_422J2_124_3477_n550) );
  FADDX1_HVT DP_OP_422J2_124_3477_U370 ( .A(DP_OP_422J2_124_3477_n747), .B(
        DP_OP_422J2_124_3477_n743), .CI(DP_OP_422J2_124_3477_n741), .CO(
        DP_OP_422J2_124_3477_n547), .S(DP_OP_422J2_124_3477_n548) );
  FADDX1_HVT DP_OP_422J2_124_3477_U369 ( .A(DP_OP_422J2_124_3477_n739), .B(
        DP_OP_422J2_124_3477_n578), .CI(DP_OP_422J2_124_3477_n576), .CO(
        DP_OP_422J2_124_3477_n545), .S(DP_OP_422J2_124_3477_n546) );
  FADDX1_HVT DP_OP_422J2_124_3477_U368 ( .A(DP_OP_422J2_124_3477_n737), .B(
        DP_OP_422J2_124_3477_n568), .CI(DP_OP_422J2_124_3477_n729), .CO(
        DP_OP_422J2_124_3477_n543), .S(DP_OP_422J2_124_3477_n544) );
  FADDX1_HVT DP_OP_422J2_124_3477_U367 ( .A(DP_OP_422J2_124_3477_n735), .B(
        DP_OP_422J2_124_3477_n731), .CI(DP_OP_422J2_124_3477_n570), .CO(
        DP_OP_422J2_124_3477_n541), .S(DP_OP_422J2_124_3477_n542) );
  FADDX1_HVT DP_OP_422J2_124_3477_U366 ( .A(DP_OP_422J2_124_3477_n733), .B(
        DP_OP_422J2_124_3477_n574), .CI(DP_OP_422J2_124_3477_n572), .CO(
        DP_OP_422J2_124_3477_n539), .S(DP_OP_422J2_124_3477_n540) );
  FADDX1_HVT DP_OP_422J2_124_3477_U365 ( .A(DP_OP_422J2_124_3477_n566), .B(
        DP_OP_422J2_124_3477_n564), .CI(DP_OP_422J2_124_3477_n727), .CO(
        DP_OP_422J2_124_3477_n537), .S(DP_OP_422J2_124_3477_n538) );
  FADDX1_HVT DP_OP_422J2_124_3477_U364 ( .A(DP_OP_422J2_124_3477_n725), .B(
        DP_OP_422J2_124_3477_n723), .CI(DP_OP_422J2_124_3477_n556), .CO(
        DP_OP_422J2_124_3477_n535), .S(DP_OP_422J2_124_3477_n536) );
  FADDX1_HVT DP_OP_422J2_124_3477_U363 ( .A(DP_OP_422J2_124_3477_n560), .B(
        DP_OP_422J2_124_3477_n558), .CI(DP_OP_422J2_124_3477_n562), .CO(
        DP_OP_422J2_124_3477_n533), .S(DP_OP_422J2_124_3477_n534) );
  FADDX1_HVT DP_OP_422J2_124_3477_U362 ( .A(DP_OP_422J2_124_3477_n554), .B(
        DP_OP_422J2_124_3477_n721), .CI(DP_OP_422J2_124_3477_n552), .CO(
        DP_OP_422J2_124_3477_n531), .S(DP_OP_422J2_124_3477_n532) );
  FADDX1_HVT DP_OP_422J2_124_3477_U361 ( .A(DP_OP_422J2_124_3477_n719), .B(
        DP_OP_422J2_124_3477_n717), .CI(DP_OP_422J2_124_3477_n550), .CO(
        DP_OP_422J2_124_3477_n529), .S(DP_OP_422J2_124_3477_n530) );
  FADDX1_HVT DP_OP_422J2_124_3477_U360 ( .A(DP_OP_422J2_124_3477_n715), .B(
        DP_OP_422J2_124_3477_n713), .CI(DP_OP_422J2_124_3477_n548), .CO(
        DP_OP_422J2_124_3477_n527), .S(DP_OP_422J2_124_3477_n528) );
  FADDX1_HVT DP_OP_422J2_124_3477_U359 ( .A(DP_OP_422J2_124_3477_n711), .B(
        DP_OP_422J2_124_3477_n546), .CI(DP_OP_422J2_124_3477_n709), .CO(
        DP_OP_422J2_124_3477_n525), .S(DP_OP_422J2_124_3477_n526) );
  FADDX1_HVT DP_OP_422J2_124_3477_U358 ( .A(DP_OP_422J2_124_3477_n544), .B(
        DP_OP_422J2_124_3477_n542), .CI(DP_OP_422J2_124_3477_n540), .CO(
        DP_OP_422J2_124_3477_n523), .S(DP_OP_422J2_124_3477_n524) );
  FADDX1_HVT DP_OP_422J2_124_3477_U357 ( .A(DP_OP_422J2_124_3477_n707), .B(
        DP_OP_422J2_124_3477_n705), .CI(DP_OP_422J2_124_3477_n538), .CO(
        DP_OP_422J2_124_3477_n521), .S(DP_OP_422J2_124_3477_n522) );
  FADDX1_HVT DP_OP_422J2_124_3477_U356 ( .A(DP_OP_422J2_124_3477_n703), .B(
        DP_OP_422J2_124_3477_n534), .CI(DP_OP_422J2_124_3477_n536), .CO(
        DP_OP_422J2_124_3477_n519), .S(DP_OP_422J2_124_3477_n520) );
  FADDX1_HVT DP_OP_422J2_124_3477_U355 ( .A(DP_OP_422J2_124_3477_n701), .B(
        DP_OP_422J2_124_3477_n532), .CI(DP_OP_422J2_124_3477_n699), .CO(
        DP_OP_422J2_124_3477_n517), .S(DP_OP_422J2_124_3477_n518) );
  FADDX1_HVT DP_OP_422J2_124_3477_U354 ( .A(DP_OP_422J2_124_3477_n697), .B(
        DP_OP_422J2_124_3477_n530), .CI(DP_OP_422J2_124_3477_n695), .CO(
        DP_OP_422J2_124_3477_n515), .S(DP_OP_422J2_124_3477_n516) );
  FADDX1_HVT DP_OP_422J2_124_3477_U353 ( .A(DP_OP_422J2_124_3477_n528), .B(
        DP_OP_422J2_124_3477_n693), .CI(DP_OP_422J2_124_3477_n526), .CO(
        DP_OP_422J2_124_3477_n513), .S(DP_OP_422J2_124_3477_n514) );
  FADDX1_HVT DP_OP_422J2_124_3477_U352 ( .A(DP_OP_422J2_124_3477_n524), .B(
        DP_OP_422J2_124_3477_n691), .CI(DP_OP_422J2_124_3477_n522), .CO(
        DP_OP_422J2_124_3477_n511), .S(DP_OP_422J2_124_3477_n512) );
  FADDX1_HVT DP_OP_422J2_124_3477_U351 ( .A(DP_OP_422J2_124_3477_n689), .B(
        DP_OP_422J2_124_3477_n520), .CI(DP_OP_422J2_124_3477_n687), .CO(
        DP_OP_422J2_124_3477_n509), .S(DP_OP_422J2_124_3477_n510) );
  FADDX1_HVT DP_OP_422J2_124_3477_U350 ( .A(DP_OP_422J2_124_3477_n518), .B(
        DP_OP_422J2_124_3477_n685), .CI(DP_OP_422J2_124_3477_n516), .CO(
        DP_OP_422J2_124_3477_n507), .S(DP_OP_422J2_124_3477_n508) );
  FADDX1_HVT DP_OP_422J2_124_3477_U349 ( .A(DP_OP_422J2_124_3477_n683), .B(
        DP_OP_422J2_124_3477_n514), .CI(DP_OP_422J2_124_3477_n512), .CO(
        DP_OP_422J2_124_3477_n505), .S(DP_OP_422J2_124_3477_n506) );
  FADDX1_HVT DP_OP_422J2_124_3477_U348 ( .A(DP_OP_422J2_124_3477_n681), .B(
        DP_OP_422J2_124_3477_n510), .CI(DP_OP_422J2_124_3477_n679), .CO(
        DP_OP_422J2_124_3477_n503), .S(DP_OP_422J2_124_3477_n504) );
  FADDX1_HVT DP_OP_422J2_124_3477_U347 ( .A(DP_OP_422J2_124_3477_n508), .B(
        DP_OP_422J2_124_3477_n677), .CI(DP_OP_422J2_124_3477_n506), .CO(
        DP_OP_422J2_124_3477_n501), .S(DP_OP_422J2_124_3477_n502) );
  FADDX1_HVT DP_OP_422J2_124_3477_U346 ( .A(DP_OP_422J2_124_3477_n675), .B(
        DP_OP_422J2_124_3477_n504), .CI(DP_OP_422J2_124_3477_n502), .CO(
        DP_OP_422J2_124_3477_n499), .S(DP_OP_422J2_124_3477_n500) );
  FADDX1_HVT DP_OP_422J2_124_3477_U345 ( .A(DP_OP_422J2_124_3477_n671), .B(
        DP_OP_422J2_124_3477_n2533), .CI(DP_OP_422J2_124_3477_n2577), .CO(
        DP_OP_422J2_124_3477_n497), .S(DP_OP_422J2_124_3477_n498) );
  FADDX1_HVT DP_OP_422J2_124_3477_U344 ( .A(DP_OP_422J2_124_3477_n1999), .B(
        DP_OP_422J2_124_3477_n1962), .CI(DP_OP_422J2_124_3477_n2225), .CO(
        DP_OP_422J2_124_3477_n495), .S(DP_OP_422J2_124_3477_n496) );
  FADDX1_HVT DP_OP_422J2_124_3477_U343 ( .A(DP_OP_422J2_124_3477_n2701), .B(
        DP_OP_422J2_124_3477_n1823), .CI(DP_OP_422J2_124_3477_n2445), .CO(
        DP_OP_422J2_124_3477_n493), .S(DP_OP_422J2_124_3477_n494) );
  FADDX1_HVT DP_OP_422J2_124_3477_U342 ( .A(DP_OP_422J2_124_3477_n2614), .B(
        DP_OP_422J2_124_3477_n1911), .CI(DP_OP_422J2_124_3477_n2093), .CO(
        DP_OP_422J2_124_3477_n491), .S(DP_OP_422J2_124_3477_n492) );
  FADDX1_HVT DP_OP_422J2_124_3477_U341 ( .A(DP_OP_422J2_124_3477_n1867), .B(
        DP_OP_422J2_124_3477_n2438), .CI(DP_OP_422J2_124_3477_n1955), .CO(
        DP_OP_422J2_124_3477_n489), .S(DP_OP_422J2_124_3477_n490) );
  FADDX1_HVT DP_OP_422J2_124_3477_U340 ( .A(DP_OP_422J2_124_3477_n2788), .B(
        DP_OP_422J2_124_3477_n2482), .CI(DP_OP_422J2_124_3477_n2744), .CO(
        DP_OP_422J2_124_3477_n487), .S(DP_OP_422J2_124_3477_n488) );
  FADDX1_HVT DP_OP_422J2_124_3477_U339 ( .A(DP_OP_422J2_124_3477_n2086), .B(
        DP_OP_422J2_124_3477_n2526), .CI(DP_OP_422J2_124_3477_n2174), .CO(
        DP_OP_422J2_124_3477_n485), .S(DP_OP_422J2_124_3477_n486) );
  FADDX1_HVT DP_OP_422J2_124_3477_U338 ( .A(DP_OP_422J2_124_3477_n2658), .B(
        DP_OP_422J2_124_3477_n2042), .CI(DP_OP_422J2_124_3477_n2570), .CO(
        DP_OP_422J2_124_3477_n483), .S(DP_OP_422J2_124_3477_n484) );
  FADDX1_HVT DP_OP_422J2_124_3477_U337 ( .A(DP_OP_422J2_124_3477_n2306), .B(
        DP_OP_422J2_124_3477_n2751), .CI(DP_OP_422J2_124_3477_n2876), .CO(
        DP_OP_422J2_124_3477_n481), .S(DP_OP_422J2_124_3477_n482) );
  FADDX1_HVT DP_OP_422J2_124_3477_U336 ( .A(DP_OP_422J2_124_3477_n2130), .B(
        DP_OP_422J2_124_3477_n2839), .CI(DP_OP_422J2_124_3477_n2883), .CO(
        DP_OP_422J2_124_3477_n479), .S(DP_OP_422J2_124_3477_n480) );
  FADDX1_HVT DP_OP_422J2_124_3477_U335 ( .A(DP_OP_422J2_124_3477_n2832), .B(
        DP_OP_422J2_124_3477_n2350), .CI(DP_OP_422J2_124_3477_n2262), .CO(
        DP_OP_422J2_124_3477_n477), .S(DP_OP_422J2_124_3477_n478) );
  FADDX1_HVT DP_OP_422J2_124_3477_U334 ( .A(DP_OP_422J2_124_3477_n2394), .B(
        DP_OP_422J2_124_3477_n2357), .CI(DP_OP_422J2_124_3477_n1874), .CO(
        DP_OP_422J2_124_3477_n475), .S(DP_OP_422J2_124_3477_n476) );
  FADDX1_HVT DP_OP_422J2_124_3477_U333 ( .A(DP_OP_422J2_124_3477_n2137), .B(
        DP_OP_422J2_124_3477_n2489), .CI(DP_OP_422J2_124_3477_n2401), .CO(
        DP_OP_422J2_124_3477_n473), .S(DP_OP_422J2_124_3477_n474) );
  FADDX1_HVT DP_OP_422J2_124_3477_U332 ( .A(DP_OP_422J2_124_3477_n2269), .B(
        DP_OP_422J2_124_3477_n2218), .CI(DP_OP_422J2_124_3477_n2049), .CO(
        DP_OP_422J2_124_3477_n471), .S(DP_OP_422J2_124_3477_n472) );
  FADDX1_HVT DP_OP_422J2_124_3477_U331 ( .A(DP_OP_422J2_124_3477_n1779), .B(
        DP_OP_422J2_124_3477_n2707), .CI(DP_OP_422J2_124_3477_n1830), .CO(
        DP_OP_422J2_124_3477_n469), .S(DP_OP_422J2_124_3477_n470) );
  FADDX1_HVT DP_OP_422J2_124_3477_U330 ( .A(DP_OP_422J2_124_3477_n2665), .B(
        DP_OP_422J2_124_3477_n2313), .CI(DP_OP_422J2_124_3477_n1918), .CO(
        DP_OP_422J2_124_3477_n467), .S(DP_OP_422J2_124_3477_n468) );
  FADDX1_HVT DP_OP_422J2_124_3477_U329 ( .A(DP_OP_422J2_124_3477_n2795), .B(
        DP_OP_422J2_124_3477_n2005), .CI(DP_OP_422J2_124_3477_n2181), .CO(
        DP_OP_422J2_124_3477_n465), .S(DP_OP_422J2_124_3477_n466) );
  FADDX1_HVT DP_OP_422J2_124_3477_U328 ( .A(DP_OP_422J2_124_3477_n2621), .B(
        DP_OP_422J2_124_3477_n669), .CI(DP_OP_422J2_124_3477_n667), .CO(
        DP_OP_422J2_124_3477_n463), .S(DP_OP_422J2_124_3477_n464) );
  FADDX1_HVT DP_OP_422J2_124_3477_U327 ( .A(DP_OP_422J2_124_3477_n665), .B(
        DP_OP_422J2_124_3477_n651), .CI(DP_OP_422J2_124_3477_n653), .CO(
        DP_OP_422J2_124_3477_n461), .S(DP_OP_422J2_124_3477_n462) );
  FADDX1_HVT DP_OP_422J2_124_3477_U326 ( .A(DP_OP_422J2_124_3477_n663), .B(
        DP_OP_422J2_124_3477_n655), .CI(DP_OP_422J2_124_3477_n657), .CO(
        DP_OP_422J2_124_3477_n459), .S(DP_OP_422J2_124_3477_n460) );
  FADDX1_HVT DP_OP_422J2_124_3477_U325 ( .A(DP_OP_422J2_124_3477_n661), .B(
        DP_OP_422J2_124_3477_n659), .CI(DP_OP_422J2_124_3477_n649), .CO(
        DP_OP_422J2_124_3477_n457), .S(DP_OP_422J2_124_3477_n458) );
  FADDX1_HVT DP_OP_422J2_124_3477_U324 ( .A(DP_OP_422J2_124_3477_n647), .B(
        DP_OP_422J2_124_3477_n635), .CI(DP_OP_422J2_124_3477_n627), .CO(
        DP_OP_422J2_124_3477_n455), .S(DP_OP_422J2_124_3477_n456) );
  FADDX1_HVT DP_OP_422J2_124_3477_U323 ( .A(DP_OP_422J2_124_3477_n645), .B(
        DP_OP_422J2_124_3477_n637), .CI(DP_OP_422J2_124_3477_n629), .CO(
        DP_OP_422J2_124_3477_n453), .S(DP_OP_422J2_124_3477_n454) );
  FADDX1_HVT DP_OP_422J2_124_3477_U322 ( .A(DP_OP_422J2_124_3477_n643), .B(
        DP_OP_422J2_124_3477_n639), .CI(DP_OP_422J2_124_3477_n631), .CO(
        DP_OP_422J2_124_3477_n451), .S(DP_OP_422J2_124_3477_n452) );
  FADDX1_HVT DP_OP_422J2_124_3477_U321 ( .A(DP_OP_422J2_124_3477_n641), .B(
        DP_OP_422J2_124_3477_n633), .CI(DP_OP_422J2_124_3477_n625), .CO(
        DP_OP_422J2_124_3477_n449), .S(DP_OP_422J2_124_3477_n450) );
  FADDX1_HVT DP_OP_422J2_124_3477_U320 ( .A(DP_OP_422J2_124_3477_n496), .B(
        DP_OP_422J2_124_3477_n623), .CI(DP_OP_422J2_124_3477_n621), .CO(
        DP_OP_422J2_124_3477_n447), .S(DP_OP_422J2_124_3477_n448) );
  FADDX1_HVT DP_OP_422J2_124_3477_U319 ( .A(DP_OP_422J2_124_3477_n498), .B(
        DP_OP_422J2_124_3477_n486), .CI(DP_OP_422J2_124_3477_n488), .CO(
        DP_OP_422J2_124_3477_n445), .S(DP_OP_422J2_124_3477_n446) );
  FADDX1_HVT DP_OP_422J2_124_3477_U318 ( .A(DP_OP_422J2_124_3477_n494), .B(
        DP_OP_422J2_124_3477_n478), .CI(DP_OP_422J2_124_3477_n484), .CO(
        DP_OP_422J2_124_3477_n443), .S(DP_OP_422J2_124_3477_n444) );
  FADDX1_HVT DP_OP_422J2_124_3477_U317 ( .A(DP_OP_422J2_124_3477_n482), .B(
        DP_OP_422J2_124_3477_n480), .CI(DP_OP_422J2_124_3477_n490), .CO(
        DP_OP_422J2_124_3477_n441), .S(DP_OP_422J2_124_3477_n442) );
  FADDX1_HVT DP_OP_422J2_124_3477_U316 ( .A(DP_OP_422J2_124_3477_n492), .B(
        DP_OP_422J2_124_3477_n476), .CI(DP_OP_422J2_124_3477_n474), .CO(
        DP_OP_422J2_124_3477_n439), .S(DP_OP_422J2_124_3477_n440) );
  FADDX1_HVT DP_OP_422J2_124_3477_U315 ( .A(DP_OP_422J2_124_3477_n472), .B(
        DP_OP_422J2_124_3477_n470), .CI(DP_OP_422J2_124_3477_n468), .CO(
        DP_OP_422J2_124_3477_n437), .S(DP_OP_422J2_124_3477_n438) );
  FADDX1_HVT DP_OP_422J2_124_3477_U314 ( .A(DP_OP_422J2_124_3477_n466), .B(
        DP_OP_422J2_124_3477_n619), .CI(DP_OP_422J2_124_3477_n617), .CO(
        DP_OP_422J2_124_3477_n435), .S(DP_OP_422J2_124_3477_n436) );
  FADDX1_HVT DP_OP_422J2_124_3477_U313 ( .A(DP_OP_422J2_124_3477_n615), .B(
        DP_OP_422J2_124_3477_n611), .CI(DP_OP_422J2_124_3477_n613), .CO(
        DP_OP_422J2_124_3477_n433), .S(DP_OP_422J2_124_3477_n434) );
  FADDX1_HVT DP_OP_422J2_124_3477_U312 ( .A(DP_OP_422J2_124_3477_n609), .B(
        DP_OP_422J2_124_3477_n605), .CI(DP_OP_422J2_124_3477_n607), .CO(
        DP_OP_422J2_124_3477_n431), .S(DP_OP_422J2_124_3477_n432) );
  FADDX1_HVT DP_OP_422J2_124_3477_U311 ( .A(DP_OP_422J2_124_3477_n464), .B(
        DP_OP_422J2_124_3477_n591), .CI(DP_OP_422J2_124_3477_n458), .CO(
        DP_OP_422J2_124_3477_n429), .S(DP_OP_422J2_124_3477_n430) );
  FADDX1_HVT DP_OP_422J2_124_3477_U310 ( .A(DP_OP_422J2_124_3477_n603), .B(
        DP_OP_422J2_124_3477_n462), .CI(DP_OP_422J2_124_3477_n460), .CO(
        DP_OP_422J2_124_3477_n427), .S(DP_OP_422J2_124_3477_n428) );
  FADDX1_HVT DP_OP_422J2_124_3477_U309 ( .A(DP_OP_422J2_124_3477_n601), .B(
        DP_OP_422J2_124_3477_n595), .CI(DP_OP_422J2_124_3477_n593), .CO(
        DP_OP_422J2_124_3477_n425), .S(DP_OP_422J2_124_3477_n426) );
  FADDX1_HVT DP_OP_422J2_124_3477_U308 ( .A(DP_OP_422J2_124_3477_n599), .B(
        DP_OP_422J2_124_3477_n597), .CI(DP_OP_422J2_124_3477_n589), .CO(
        DP_OP_422J2_124_3477_n423), .S(DP_OP_422J2_124_3477_n424) );
  FADDX1_HVT DP_OP_422J2_124_3477_U307 ( .A(DP_OP_422J2_124_3477_n454), .B(
        DP_OP_422J2_124_3477_n583), .CI(DP_OP_422J2_124_3477_n450), .CO(
        DP_OP_422J2_124_3477_n421), .S(DP_OP_422J2_124_3477_n422) );
  FADDX1_HVT DP_OP_422J2_124_3477_U306 ( .A(DP_OP_422J2_124_3477_n587), .B(
        DP_OP_422J2_124_3477_n585), .CI(DP_OP_422J2_124_3477_n452), .CO(
        DP_OP_422J2_124_3477_n419), .S(DP_OP_422J2_124_3477_n420) );
  FADDX1_HVT DP_OP_422J2_124_3477_U305 ( .A(DP_OP_422J2_124_3477_n456), .B(
        DP_OP_422J2_124_3477_n581), .CI(DP_OP_422J2_124_3477_n444), .CO(
        DP_OP_422J2_124_3477_n417), .S(DP_OP_422J2_124_3477_n418) );
  FADDX1_HVT DP_OP_422J2_124_3477_U304 ( .A(DP_OP_422J2_124_3477_n446), .B(
        DP_OP_422J2_124_3477_n442), .CI(DP_OP_422J2_124_3477_n440), .CO(
        DP_OP_422J2_124_3477_n415), .S(DP_OP_422J2_124_3477_n416) );
  FADDX1_HVT DP_OP_422J2_124_3477_U303 ( .A(DP_OP_422J2_124_3477_n448), .B(
        DP_OP_422J2_124_3477_n438), .CI(DP_OP_422J2_124_3477_n579), .CO(
        DP_OP_422J2_124_3477_n413), .S(DP_OP_422J2_124_3477_n414) );
  FADDX1_HVT DP_OP_422J2_124_3477_U302 ( .A(DP_OP_422J2_124_3477_n577), .B(
        DP_OP_422J2_124_3477_n575), .CI(DP_OP_422J2_124_3477_n436), .CO(
        DP_OP_422J2_124_3477_n411), .S(DP_OP_422J2_124_3477_n412) );
  FADDX1_HVT DP_OP_422J2_124_3477_U301 ( .A(DP_OP_422J2_124_3477_n573), .B(
        DP_OP_422J2_124_3477_n567), .CI(DP_OP_422J2_124_3477_n434), .CO(
        DP_OP_422J2_124_3477_n409), .S(DP_OP_422J2_124_3477_n410) );
  FADDX1_HVT DP_OP_422J2_124_3477_U300 ( .A(DP_OP_422J2_124_3477_n571), .B(
        DP_OP_422J2_124_3477_n569), .CI(DP_OP_422J2_124_3477_n565), .CO(
        DP_OP_422J2_124_3477_n407), .S(DP_OP_422J2_124_3477_n408) );
  FADDX1_HVT DP_OP_422J2_124_3477_U299 ( .A(DP_OP_422J2_124_3477_n432), .B(
        DP_OP_422J2_124_3477_n563), .CI(DP_OP_422J2_124_3477_n430), .CO(
        DP_OP_422J2_124_3477_n405), .S(DP_OP_422J2_124_3477_n406) );
  FADDX1_HVT DP_OP_422J2_124_3477_U298 ( .A(DP_OP_422J2_124_3477_n561), .B(
        DP_OP_422J2_124_3477_n555), .CI(DP_OP_422J2_124_3477_n424), .CO(
        DP_OP_422J2_124_3477_n403), .S(DP_OP_422J2_124_3477_n404) );
  FADDX1_HVT DP_OP_422J2_124_3477_U297 ( .A(DP_OP_422J2_124_3477_n559), .B(
        DP_OP_422J2_124_3477_n426), .CI(DP_OP_422J2_124_3477_n428), .CO(
        DP_OP_422J2_124_3477_n401), .S(DP_OP_422J2_124_3477_n402) );
  FADDX1_HVT DP_OP_422J2_124_3477_U296 ( .A(DP_OP_422J2_124_3477_n557), .B(
        DP_OP_422J2_124_3477_n553), .CI(DP_OP_422J2_124_3477_n422), .CO(
        DP_OP_422J2_124_3477_n399), .S(DP_OP_422J2_124_3477_n400) );
  FADDX1_HVT DP_OP_422J2_124_3477_U295 ( .A(DP_OP_422J2_124_3477_n420), .B(
        DP_OP_422J2_124_3477_n551), .CI(DP_OP_422J2_124_3477_n418), .CO(
        DP_OP_422J2_124_3477_n397), .S(DP_OP_422J2_124_3477_n398) );
  FADDX1_HVT DP_OP_422J2_124_3477_U294 ( .A(DP_OP_422J2_124_3477_n416), .B(
        DP_OP_422J2_124_3477_n414), .CI(DP_OP_422J2_124_3477_n549), .CO(
        DP_OP_422J2_124_3477_n395), .S(DP_OP_422J2_124_3477_n396) );
  FADDX1_HVT DP_OP_422J2_124_3477_U293 ( .A(DP_OP_422J2_124_3477_n547), .B(
        DP_OP_422J2_124_3477_n545), .CI(DP_OP_422J2_124_3477_n412), .CO(
        DP_OP_422J2_124_3477_n393), .S(DP_OP_422J2_124_3477_n394) );
  FADDX1_HVT DP_OP_422J2_124_3477_U292 ( .A(DP_OP_422J2_124_3477_n543), .B(
        DP_OP_422J2_124_3477_n410), .CI(DP_OP_422J2_124_3477_n408), .CO(
        DP_OP_422J2_124_3477_n391), .S(DP_OP_422J2_124_3477_n392) );
  FADDX1_HVT DP_OP_422J2_124_3477_U291 ( .A(DP_OP_422J2_124_3477_n541), .B(
        DP_OP_422J2_124_3477_n539), .CI(DP_OP_422J2_124_3477_n537), .CO(
        DP_OP_422J2_124_3477_n389), .S(DP_OP_422J2_124_3477_n390) );
  FADDX1_HVT DP_OP_422J2_124_3477_U290 ( .A(DP_OP_422J2_124_3477_n406), .B(
        DP_OP_422J2_124_3477_n535), .CI(DP_OP_422J2_124_3477_n402), .CO(
        DP_OP_422J2_124_3477_n387), .S(DP_OP_422J2_124_3477_n388) );
  FADDX1_HVT DP_OP_422J2_124_3477_U289 ( .A(DP_OP_422J2_124_3477_n404), .B(
        DP_OP_422J2_124_3477_n533), .CI(DP_OP_422J2_124_3477_n400), .CO(
        DP_OP_422J2_124_3477_n385), .S(DP_OP_422J2_124_3477_n386) );
  FADDX1_HVT DP_OP_422J2_124_3477_U288 ( .A(DP_OP_422J2_124_3477_n531), .B(
        DP_OP_422J2_124_3477_n398), .CI(DP_OP_422J2_124_3477_n529), .CO(
        DP_OP_422J2_124_3477_n383), .S(DP_OP_422J2_124_3477_n384) );
  FADDX1_HVT DP_OP_422J2_124_3477_U287 ( .A(DP_OP_422J2_124_3477_n396), .B(
        DP_OP_422J2_124_3477_n527), .CI(DP_OP_422J2_124_3477_n394), .CO(
        DP_OP_422J2_124_3477_n381), .S(DP_OP_422J2_124_3477_n382) );
  FADDX1_HVT DP_OP_422J2_124_3477_U286 ( .A(DP_OP_422J2_124_3477_n525), .B(
        DP_OP_422J2_124_3477_n523), .CI(DP_OP_422J2_124_3477_n392), .CO(
        DP_OP_422J2_124_3477_n379), .S(DP_OP_422J2_124_3477_n380) );
  FADDX1_HVT DP_OP_422J2_124_3477_U285 ( .A(DP_OP_422J2_124_3477_n390), .B(
        DP_OP_422J2_124_3477_n521), .CI(DP_OP_422J2_124_3477_n519), .CO(
        DP_OP_422J2_124_3477_n377), .S(DP_OP_422J2_124_3477_n378) );
  FADDX1_HVT DP_OP_422J2_124_3477_U284 ( .A(DP_OP_422J2_124_3477_n388), .B(
        DP_OP_422J2_124_3477_n386), .CI(DP_OP_422J2_124_3477_n517), .CO(
        DP_OP_422J2_124_3477_n375), .S(DP_OP_422J2_124_3477_n376) );
  FADDX1_HVT DP_OP_422J2_124_3477_U283 ( .A(DP_OP_422J2_124_3477_n384), .B(
        DP_OP_422J2_124_3477_n515), .CI(DP_OP_422J2_124_3477_n382), .CO(
        DP_OP_422J2_124_3477_n373), .S(DP_OP_422J2_124_3477_n374) );
  FADDX1_HVT DP_OP_422J2_124_3477_U282 ( .A(DP_OP_422J2_124_3477_n513), .B(
        DP_OP_422J2_124_3477_n380), .CI(DP_OP_422J2_124_3477_n511), .CO(
        DP_OP_422J2_124_3477_n371), .S(DP_OP_422J2_124_3477_n372) );
  FADDX1_HVT DP_OP_422J2_124_3477_U281 ( .A(DP_OP_422J2_124_3477_n378), .B(
        DP_OP_422J2_124_3477_n509), .CI(DP_OP_422J2_124_3477_n376), .CO(
        DP_OP_422J2_124_3477_n369), .S(DP_OP_422J2_124_3477_n370) );
  FADDX1_HVT DP_OP_422J2_124_3477_U280 ( .A(DP_OP_422J2_124_3477_n507), .B(
        DP_OP_422J2_124_3477_n374), .CI(DP_OP_422J2_124_3477_n505), .CO(
        DP_OP_422J2_124_3477_n367), .S(DP_OP_422J2_124_3477_n368) );
  FADDX1_HVT DP_OP_422J2_124_3477_U279 ( .A(DP_OP_422J2_124_3477_n372), .B(
        DP_OP_422J2_124_3477_n370), .CI(DP_OP_422J2_124_3477_n503), .CO(
        DP_OP_422J2_124_3477_n365), .S(DP_OP_422J2_124_3477_n366) );
  FADDX1_HVT DP_OP_422J2_124_3477_U278 ( .A(DP_OP_422J2_124_3477_n501), .B(
        DP_OP_422J2_124_3477_n368), .CI(DP_OP_422J2_124_3477_n366), .CO(
        DP_OP_422J2_124_3477_n363), .S(DP_OP_422J2_124_3477_n364) );
  FADDX1_HVT DP_OP_422J2_124_3477_U276 ( .A(DP_OP_422J2_124_3477_n1998), .B(
        DP_OP_422J2_124_3477_n1822), .CI(DP_OP_422J2_124_3477_n2743), .CO(
        DP_OP_422J2_124_3477_n359), .S(DP_OP_422J2_124_3477_n360) );
  FADDX1_HVT DP_OP_422J2_124_3477_U275 ( .A(DP_OP_422J2_124_3477_n2613), .B(
        DP_OP_422J2_124_3477_n2437), .CI(DP_OP_422J2_124_3477_n1954), .CO(
        DP_OP_422J2_124_3477_n357), .S(DP_OP_422J2_124_3477_n358) );
  FADDX1_HVT DP_OP_422J2_124_3477_U274 ( .A(DP_OP_422J2_124_3477_n2305), .B(
        DP_OP_422J2_124_3477_n2569), .CI(DP_OP_422J2_124_3477_n2525), .CO(
        DP_OP_422J2_124_3477_n355), .S(DP_OP_422J2_124_3477_n356) );
  FADDX1_HVT DP_OP_422J2_124_3477_U273 ( .A(DP_OP_422J2_124_3477_n2831), .B(
        DP_OP_422J2_124_3477_n1910), .CI(DP_OP_422J2_124_3477_n2481), .CO(
        DP_OP_422J2_124_3477_n353), .S(DP_OP_422J2_124_3477_n354) );
  FADDX1_HVT DP_OP_422J2_124_3477_U272 ( .A(DP_OP_422J2_124_3477_n2085), .B(
        DP_OP_422J2_124_3477_n2041), .CI(DP_OP_422J2_124_3477_n2173), .CO(
        DP_OP_422J2_124_3477_n351), .S(DP_OP_422J2_124_3477_n352) );
  FADDX1_HVT DP_OP_422J2_124_3477_U271 ( .A(DP_OP_422J2_124_3477_n2349), .B(
        DP_OP_422J2_124_3477_n1778), .CI(DP_OP_422J2_124_3477_n2875), .CO(
        DP_OP_422J2_124_3477_n349), .S(DP_OP_422J2_124_3477_n350) );
  FADDX1_HVT DP_OP_422J2_124_3477_U270 ( .A(DP_OP_422J2_124_3477_n2657), .B(
        DP_OP_422J2_124_3477_n2129), .CI(DP_OP_422J2_124_3477_n2261), .CO(
        DP_OP_422J2_124_3477_n347), .S(DP_OP_422J2_124_3477_n348) );
  FADDX1_HVT DP_OP_422J2_124_3477_U269 ( .A(DP_OP_422J2_124_3477_n2787), .B(
        DP_OP_422J2_124_3477_n1866), .CI(DP_OP_422J2_124_3477_n2393), .CO(
        DP_OP_422J2_124_3477_n345), .S(DP_OP_422J2_124_3477_n346) );
  FADDX1_HVT DP_OP_422J2_124_3477_U268 ( .A(DP_OP_422J2_124_3477_n2217), .B(
        DP_OP_422J2_124_3477_n362), .CI(DP_OP_422J2_124_3477_n497), .CO(
        DP_OP_422J2_124_3477_n343), .S(DP_OP_422J2_124_3477_n344) );
  FADDX1_HVT DP_OP_422J2_124_3477_U267 ( .A(DP_OP_422J2_124_3477_n495), .B(
        DP_OP_422J2_124_3477_n477), .CI(DP_OP_422J2_124_3477_n479), .CO(
        DP_OP_422J2_124_3477_n341), .S(DP_OP_422J2_124_3477_n342) );
  FADDX1_HVT DP_OP_422J2_124_3477_U266 ( .A(DP_OP_422J2_124_3477_n493), .B(
        DP_OP_422J2_124_3477_n481), .CI(DP_OP_422J2_124_3477_n483), .CO(
        DP_OP_422J2_124_3477_n339), .S(DP_OP_422J2_124_3477_n340) );
  FADDX1_HVT DP_OP_422J2_124_3477_U265 ( .A(DP_OP_422J2_124_3477_n491), .B(
        DP_OP_422J2_124_3477_n485), .CI(DP_OP_422J2_124_3477_n487), .CO(
        DP_OP_422J2_124_3477_n337), .S(DP_OP_422J2_124_3477_n338) );
  FADDX1_HVT DP_OP_422J2_124_3477_U264 ( .A(DP_OP_422J2_124_3477_n489), .B(
        DP_OP_422J2_124_3477_n475), .CI(DP_OP_422J2_124_3477_n473), .CO(
        DP_OP_422J2_124_3477_n335), .S(DP_OP_422J2_124_3477_n336) );
  FADDX1_HVT DP_OP_422J2_124_3477_U263 ( .A(DP_OP_422J2_124_3477_n471), .B(
        DP_OP_422J2_124_3477_n469), .CI(DP_OP_422J2_124_3477_n467), .CO(
        DP_OP_422J2_124_3477_n333), .S(DP_OP_422J2_124_3477_n334) );
  FADDX1_HVT DP_OP_422J2_124_3477_U262 ( .A(DP_OP_422J2_124_3477_n465), .B(
        DP_OP_422J2_124_3477_n360), .CI(DP_OP_422J2_124_3477_n352), .CO(
        DP_OP_422J2_124_3477_n331), .S(DP_OP_422J2_124_3477_n332) );
  FADDX1_HVT DP_OP_422J2_124_3477_U261 ( .A(DP_OP_422J2_124_3477_n354), .B(
        DP_OP_422J2_124_3477_n348), .CI(DP_OP_422J2_124_3477_n346), .CO(
        DP_OP_422J2_124_3477_n329), .S(DP_OP_422J2_124_3477_n330) );
  FADDX1_HVT DP_OP_422J2_124_3477_U260 ( .A(DP_OP_422J2_124_3477_n350), .B(
        DP_OP_422J2_124_3477_n358), .CI(DP_OP_422J2_124_3477_n356), .CO(
        DP_OP_422J2_124_3477_n327), .S(DP_OP_422J2_124_3477_n328) );
  FADDX1_HVT DP_OP_422J2_124_3477_U259 ( .A(DP_OP_422J2_124_3477_n463), .B(
        DP_OP_422J2_124_3477_n461), .CI(DP_OP_422J2_124_3477_n457), .CO(
        DP_OP_422J2_124_3477_n325), .S(DP_OP_422J2_124_3477_n326) );
  FADDX1_HVT DP_OP_422J2_124_3477_U258 ( .A(DP_OP_422J2_124_3477_n459), .B(
        DP_OP_422J2_124_3477_n455), .CI(DP_OP_422J2_124_3477_n453), .CO(
        DP_OP_422J2_124_3477_n323), .S(DP_OP_422J2_124_3477_n324) );
  FADDX1_HVT DP_OP_422J2_124_3477_U257 ( .A(DP_OP_422J2_124_3477_n451), .B(
        DP_OP_422J2_124_3477_n449), .CI(DP_OP_422J2_124_3477_n344), .CO(
        DP_OP_422J2_124_3477_n321), .S(DP_OP_422J2_124_3477_n322) );
  FADDX1_HVT DP_OP_422J2_124_3477_U256 ( .A(DP_OP_422J2_124_3477_n447), .B(
        DP_OP_422J2_124_3477_n338), .CI(DP_OP_422J2_124_3477_n336), .CO(
        DP_OP_422J2_124_3477_n319), .S(DP_OP_422J2_124_3477_n320) );
  FADDX1_HVT DP_OP_422J2_124_3477_U255 ( .A(DP_OP_422J2_124_3477_n445), .B(
        DP_OP_422J2_124_3477_n441), .CI(DP_OP_422J2_124_3477_n439), .CO(
        DP_OP_422J2_124_3477_n317), .S(DP_OP_422J2_124_3477_n318) );
  FADDX1_HVT DP_OP_422J2_124_3477_U254 ( .A(DP_OP_422J2_124_3477_n443), .B(
        DP_OP_422J2_124_3477_n342), .CI(DP_OP_422J2_124_3477_n340), .CO(
        DP_OP_422J2_124_3477_n315), .S(DP_OP_422J2_124_3477_n316) );
  FADDX1_HVT DP_OP_422J2_124_3477_U253 ( .A(DP_OP_422J2_124_3477_n437), .B(
        DP_OP_422J2_124_3477_n334), .CI(DP_OP_422J2_124_3477_n435), .CO(
        DP_OP_422J2_124_3477_n313), .S(DP_OP_422J2_124_3477_n314) );
  FADDX1_HVT DP_OP_422J2_124_3477_U252 ( .A(DP_OP_422J2_124_3477_n332), .B(
        DP_OP_422J2_124_3477_n328), .CI(DP_OP_422J2_124_3477_n433), .CO(
        DP_OP_422J2_124_3477_n311), .S(DP_OP_422J2_124_3477_n312) );
  FADDX1_HVT DP_OP_422J2_124_3477_U251 ( .A(DP_OP_422J2_124_3477_n330), .B(
        DP_OP_422J2_124_3477_n431), .CI(DP_OP_422J2_124_3477_n429), .CO(
        DP_OP_422J2_124_3477_n309), .S(DP_OP_422J2_124_3477_n310) );
  FADDX1_HVT DP_OP_422J2_124_3477_U250 ( .A(DP_OP_422J2_124_3477_n326), .B(
        DP_OP_422J2_124_3477_n425), .CI(DP_OP_422J2_124_3477_n423), .CO(
        DP_OP_422J2_124_3477_n307), .S(DP_OP_422J2_124_3477_n308) );
  FADDX1_HVT DP_OP_422J2_124_3477_U249 ( .A(DP_OP_422J2_124_3477_n427), .B(
        DP_OP_422J2_124_3477_n324), .CI(DP_OP_422J2_124_3477_n421), .CO(
        DP_OP_422J2_124_3477_n305), .S(DP_OP_422J2_124_3477_n306) );
  FADDX1_HVT DP_OP_422J2_124_3477_U248 ( .A(DP_OP_422J2_124_3477_n419), .B(
        DP_OP_422J2_124_3477_n322), .CI(DP_OP_422J2_124_3477_n417), .CO(
        DP_OP_422J2_124_3477_n303), .S(DP_OP_422J2_124_3477_n304) );
  FADDX1_HVT DP_OP_422J2_124_3477_U247 ( .A(DP_OP_422J2_124_3477_n415), .B(
        DP_OP_422J2_124_3477_n318), .CI(DP_OP_422J2_124_3477_n413), .CO(
        DP_OP_422J2_124_3477_n301), .S(DP_OP_422J2_124_3477_n302) );
  FADDX1_HVT DP_OP_422J2_124_3477_U246 ( .A(DP_OP_422J2_124_3477_n316), .B(
        DP_OP_422J2_124_3477_n320), .CI(DP_OP_422J2_124_3477_n314), .CO(
        DP_OP_422J2_124_3477_n299), .S(DP_OP_422J2_124_3477_n300) );
  FADDX1_HVT DP_OP_422J2_124_3477_U245 ( .A(DP_OP_422J2_124_3477_n411), .B(
        DP_OP_422J2_124_3477_n312), .CI(DP_OP_422J2_124_3477_n409), .CO(
        DP_OP_422J2_124_3477_n297), .S(DP_OP_422J2_124_3477_n298) );
  FADDX1_HVT DP_OP_422J2_124_3477_U244 ( .A(DP_OP_422J2_124_3477_n407), .B(
        DP_OP_422J2_124_3477_n405), .CI(DP_OP_422J2_124_3477_n310), .CO(
        DP_OP_422J2_124_3477_n295), .S(DP_OP_422J2_124_3477_n296) );
  FADDX1_HVT DP_OP_422J2_124_3477_U243 ( .A(DP_OP_422J2_124_3477_n308), .B(
        DP_OP_422J2_124_3477_n401), .CI(DP_OP_422J2_124_3477_n399), .CO(
        DP_OP_422J2_124_3477_n293), .S(DP_OP_422J2_124_3477_n294) );
  FADDX1_HVT DP_OP_422J2_124_3477_U242 ( .A(DP_OP_422J2_124_3477_n403), .B(
        DP_OP_422J2_124_3477_n306), .CI(DP_OP_422J2_124_3477_n304), .CO(
        DP_OP_422J2_124_3477_n291), .S(DP_OP_422J2_124_3477_n292) );
  FADDX1_HVT DP_OP_422J2_124_3477_U241 ( .A(DP_OP_422J2_124_3477_n397), .B(
        DP_OP_422J2_124_3477_n302), .CI(DP_OP_422J2_124_3477_n395), .CO(
        DP_OP_422J2_124_3477_n289), .S(DP_OP_422J2_124_3477_n290) );
  FADDX1_HVT DP_OP_422J2_124_3477_U240 ( .A(DP_OP_422J2_124_3477_n300), .B(
        DP_OP_422J2_124_3477_n393), .CI(DP_OP_422J2_124_3477_n298), .CO(
        DP_OP_422J2_124_3477_n287), .S(DP_OP_422J2_124_3477_n288) );
  FADDX1_HVT DP_OP_422J2_124_3477_U239 ( .A(DP_OP_422J2_124_3477_n391), .B(
        DP_OP_422J2_124_3477_n389), .CI(DP_OP_422J2_124_3477_n296), .CO(
        DP_OP_422J2_124_3477_n285), .S(DP_OP_422J2_124_3477_n286) );
  FADDX1_HVT DP_OP_422J2_124_3477_U238 ( .A(DP_OP_422J2_124_3477_n387), .B(
        DP_OP_422J2_124_3477_n294), .CI(DP_OP_422J2_124_3477_n292), .CO(
        DP_OP_422J2_124_3477_n283), .S(DP_OP_422J2_124_3477_n284) );
  FADDX1_HVT DP_OP_422J2_124_3477_U237 ( .A(DP_OP_422J2_124_3477_n385), .B(
        DP_OP_422J2_124_3477_n383), .CI(DP_OP_422J2_124_3477_n290), .CO(
        DP_OP_422J2_124_3477_n281), .S(DP_OP_422J2_124_3477_n282) );
  FADDX1_HVT DP_OP_422J2_124_3477_U236 ( .A(DP_OP_422J2_124_3477_n381), .B(
        DP_OP_422J2_124_3477_n288), .CI(DP_OP_422J2_124_3477_n379), .CO(
        DP_OP_422J2_124_3477_n279), .S(DP_OP_422J2_124_3477_n280) );
  FADDX1_HVT DP_OP_422J2_124_3477_U235 ( .A(DP_OP_422J2_124_3477_n286), .B(
        DP_OP_422J2_124_3477_n377), .CI(DP_OP_422J2_124_3477_n284), .CO(
        DP_OP_422J2_124_3477_n277), .S(DP_OP_422J2_124_3477_n278) );
  FADDX1_HVT DP_OP_422J2_124_3477_U234 ( .A(DP_OP_422J2_124_3477_n375), .B(
        DP_OP_422J2_124_3477_n282), .CI(DP_OP_422J2_124_3477_n373), .CO(
        DP_OP_422J2_124_3477_n275), .S(DP_OP_422J2_124_3477_n276) );
  FADDX1_HVT DP_OP_422J2_124_3477_U233 ( .A(DP_OP_422J2_124_3477_n280), .B(
        DP_OP_422J2_124_3477_n371), .CI(DP_OP_422J2_124_3477_n278), .CO(
        DP_OP_422J2_124_3477_n273), .S(DP_OP_422J2_124_3477_n274) );
  FADDX1_HVT DP_OP_422J2_124_3477_U232 ( .A(DP_OP_422J2_124_3477_n369), .B(
        DP_OP_422J2_124_3477_n276), .CI(DP_OP_422J2_124_3477_n367), .CO(
        DP_OP_422J2_124_3477_n271), .S(DP_OP_422J2_124_3477_n272) );
  FADDX1_HVT DP_OP_422J2_124_3477_U231 ( .A(DP_OP_422J2_124_3477_n274), .B(
        DP_OP_422J2_124_3477_n365), .CI(DP_OP_422J2_124_3477_n272), .CO(
        DP_OP_422J2_124_3477_n269), .S(DP_OP_422J2_124_3477_n270) );
  FADDX1_HVT DP_OP_422J2_124_3477_U230 ( .A(DP_OP_422J2_124_3477_n361), .B(
        DP_OP_422J2_124_3477_n1777), .CI(DP_OP_422J2_124_3477_n359), .CO(
        DP_OP_422J2_124_3477_n267), .S(DP_OP_422J2_124_3477_n268) );
  FADDX1_HVT DP_OP_422J2_124_3477_U229 ( .A(DP_OP_422J2_124_3477_n349), .B(
        DP_OP_422J2_124_3477_n345), .CI(DP_OP_422J2_124_3477_n357), .CO(
        DP_OP_422J2_124_3477_n265), .S(DP_OP_422J2_124_3477_n266) );
  FADDX1_HVT DP_OP_422J2_124_3477_U228 ( .A(DP_OP_422J2_124_3477_n355), .B(
        DP_OP_422J2_124_3477_n353), .CI(DP_OP_422J2_124_3477_n351), .CO(
        DP_OP_422J2_124_3477_n263), .S(DP_OP_422J2_124_3477_n264) );
  FADDX1_HVT DP_OP_422J2_124_3477_U227 ( .A(DP_OP_422J2_124_3477_n347), .B(
        DP_OP_422J2_124_3477_n343), .CI(DP_OP_422J2_124_3477_n341), .CO(
        DP_OP_422J2_124_3477_n261), .S(DP_OP_422J2_124_3477_n262) );
  FADDX1_HVT DP_OP_422J2_124_3477_U226 ( .A(DP_OP_422J2_124_3477_n339), .B(
        DP_OP_422J2_124_3477_n337), .CI(DP_OP_422J2_124_3477_n335), .CO(
        DP_OP_422J2_124_3477_n259), .S(DP_OP_422J2_124_3477_n260) );
  FADDX1_HVT DP_OP_422J2_124_3477_U225 ( .A(DP_OP_422J2_124_3477_n333), .B(
        DP_OP_422J2_124_3477_n268), .CI(DP_OP_422J2_124_3477_n331), .CO(
        DP_OP_422J2_124_3477_n257), .S(DP_OP_422J2_124_3477_n258) );
  FADDX1_HVT DP_OP_422J2_124_3477_U224 ( .A(DP_OP_422J2_124_3477_n329), .B(
        DP_OP_422J2_124_3477_n264), .CI(DP_OP_422J2_124_3477_n266), .CO(
        DP_OP_422J2_124_3477_n255), .S(DP_OP_422J2_124_3477_n256) );
  FADDX1_HVT DP_OP_422J2_124_3477_U223 ( .A(DP_OP_422J2_124_3477_n327), .B(
        DP_OP_422J2_124_3477_n325), .CI(DP_OP_422J2_124_3477_n323), .CO(
        DP_OP_422J2_124_3477_n253), .S(DP_OP_422J2_124_3477_n254) );
  FADDX1_HVT DP_OP_422J2_124_3477_U222 ( .A(DP_OP_422J2_124_3477_n321), .B(
        DP_OP_422J2_124_3477_n262), .CI(DP_OP_422J2_124_3477_n319), .CO(
        DP_OP_422J2_124_3477_n251), .S(DP_OP_422J2_124_3477_n252) );
  FADDX1_HVT DP_OP_422J2_124_3477_U221 ( .A(DP_OP_422J2_124_3477_n317), .B(
        DP_OP_422J2_124_3477_n260), .CI(DP_OP_422J2_124_3477_n315), .CO(
        DP_OP_422J2_124_3477_n249), .S(DP_OP_422J2_124_3477_n250) );
  FADDX1_HVT DP_OP_422J2_124_3477_U220 ( .A(DP_OP_422J2_124_3477_n313), .B(
        DP_OP_422J2_124_3477_n258), .CI(DP_OP_422J2_124_3477_n311), .CO(
        DP_OP_422J2_124_3477_n247), .S(DP_OP_422J2_124_3477_n248) );
  FADDX1_HVT DP_OP_422J2_124_3477_U219 ( .A(DP_OP_422J2_124_3477_n256), .B(
        DP_OP_422J2_124_3477_n309), .CI(DP_OP_422J2_124_3477_n254), .CO(
        DP_OP_422J2_124_3477_n245), .S(DP_OP_422J2_124_3477_n246) );
  FADDX1_HVT DP_OP_422J2_124_3477_U218 ( .A(DP_OP_422J2_124_3477_n307), .B(
        DP_OP_422J2_124_3477_n305), .CI(DP_OP_422J2_124_3477_n303), .CO(
        DP_OP_422J2_124_3477_n243), .S(DP_OP_422J2_124_3477_n244) );
  FADDX1_HVT DP_OP_422J2_124_3477_U217 ( .A(DP_OP_422J2_124_3477_n252), .B(
        DP_OP_422J2_124_3477_n301), .CI(DP_OP_422J2_124_3477_n250), .CO(
        DP_OP_422J2_124_3477_n241), .S(DP_OP_422J2_124_3477_n242) );
  FADDX1_HVT DP_OP_422J2_124_3477_U216 ( .A(DP_OP_422J2_124_3477_n299), .B(
        DP_OP_422J2_124_3477_n248), .CI(DP_OP_422J2_124_3477_n297), .CO(
        DP_OP_422J2_124_3477_n239), .S(DP_OP_422J2_124_3477_n240) );
  FADDX1_HVT DP_OP_422J2_124_3477_U215 ( .A(DP_OP_422J2_124_3477_n295), .B(
        DP_OP_422J2_124_3477_n246), .CI(DP_OP_422J2_124_3477_n293), .CO(
        DP_OP_422J2_124_3477_n237), .S(DP_OP_422J2_124_3477_n238) );
  FADDX1_HVT DP_OP_422J2_124_3477_U214 ( .A(DP_OP_422J2_124_3477_n291), .B(
        DP_OP_422J2_124_3477_n244), .CI(DP_OP_422J2_124_3477_n289), .CO(
        DP_OP_422J2_124_3477_n235), .S(DP_OP_422J2_124_3477_n236) );
  FADDX1_HVT DP_OP_422J2_124_3477_U213 ( .A(DP_OP_422J2_124_3477_n242), .B(
        DP_OP_422J2_124_3477_n287), .CI(DP_OP_422J2_124_3477_n240), .CO(
        DP_OP_422J2_124_3477_n233), .S(DP_OP_422J2_124_3477_n234) );
  FADDX1_HVT DP_OP_422J2_124_3477_U212 ( .A(DP_OP_422J2_124_3477_n285), .B(
        DP_OP_422J2_124_3477_n238), .CI(DP_OP_422J2_124_3477_n283), .CO(
        DP_OP_422J2_124_3477_n231), .S(DP_OP_422J2_124_3477_n232) );
  FADDX1_HVT DP_OP_422J2_124_3477_U211 ( .A(DP_OP_422J2_124_3477_n281), .B(
        DP_OP_422J2_124_3477_n236), .CI(DP_OP_422J2_124_3477_n234), .CO(
        DP_OP_422J2_124_3477_n229), .S(DP_OP_422J2_124_3477_n230) );
  FADDX1_HVT DP_OP_422J2_124_3477_U210 ( .A(DP_OP_422J2_124_3477_n279), .B(
        DP_OP_422J2_124_3477_n277), .CI(DP_OP_422J2_124_3477_n232), .CO(
        DP_OP_422J2_124_3477_n227), .S(DP_OP_422J2_124_3477_n228) );
  FADDX1_HVT DP_OP_422J2_124_3477_U209 ( .A(DP_OP_422J2_124_3477_n275), .B(
        DP_OP_422J2_124_3477_n230), .CI(DP_OP_422J2_124_3477_n273), .CO(
        DP_OP_422J2_124_3477_n225), .S(DP_OP_422J2_124_3477_n226) );
  FADDX1_HVT DP_OP_422J2_124_3477_U208 ( .A(DP_OP_422J2_124_3477_n228), .B(
        DP_OP_422J2_124_3477_n271), .CI(DP_OP_422J2_124_3477_n226), .CO(
        DP_OP_422J2_124_3477_n223), .S(DP_OP_422J2_124_3477_n224) );
  FADDX1_HVT DP_OP_422J2_124_3477_U207 ( .A(DP_OP_422J2_124_3477_n1776), .B(
        DP_OP_422J2_124_3477_n267), .CI(DP_OP_422J2_124_3477_n265), .CO(
        DP_OP_422J2_124_3477_n221), .S(DP_OP_422J2_124_3477_n222) );
  FADDX1_HVT DP_OP_422J2_124_3477_U206 ( .A(DP_OP_422J2_124_3477_n263), .B(
        DP_OP_422J2_124_3477_n261), .CI(DP_OP_422J2_124_3477_n259), .CO(
        DP_OP_422J2_124_3477_n219), .S(DP_OP_422J2_124_3477_n220) );
  FADDX1_HVT DP_OP_422J2_124_3477_U205 ( .A(DP_OP_422J2_124_3477_n257), .B(
        DP_OP_422J2_124_3477_n222), .CI(DP_OP_422J2_124_3477_n255), .CO(
        DP_OP_422J2_124_3477_n217), .S(DP_OP_422J2_124_3477_n218) );
  FADDX1_HVT DP_OP_422J2_124_3477_U204 ( .A(DP_OP_422J2_124_3477_n253), .B(
        DP_OP_422J2_124_3477_n251), .CI(DP_OP_422J2_124_3477_n220), .CO(
        DP_OP_422J2_124_3477_n215), .S(DP_OP_422J2_124_3477_n216) );
  FADDX1_HVT DP_OP_422J2_124_3477_U203 ( .A(DP_OP_422J2_124_3477_n249), .B(
        DP_OP_422J2_124_3477_n247), .CI(DP_OP_422J2_124_3477_n218), .CO(
        DP_OP_422J2_124_3477_n213), .S(DP_OP_422J2_124_3477_n214) );
  FADDX1_HVT DP_OP_422J2_124_3477_U202 ( .A(DP_OP_422J2_124_3477_n245), .B(
        DP_OP_422J2_124_3477_n243), .CI(DP_OP_422J2_124_3477_n216), .CO(
        DP_OP_422J2_124_3477_n211), .S(DP_OP_422J2_124_3477_n212) );
  FADDX1_HVT DP_OP_422J2_124_3477_U201 ( .A(DP_OP_422J2_124_3477_n241), .B(
        DP_OP_422J2_124_3477_n214), .CI(DP_OP_422J2_124_3477_n239), .CO(
        DP_OP_422J2_124_3477_n209), .S(DP_OP_422J2_124_3477_n210) );
  FADDX1_HVT DP_OP_422J2_124_3477_U200 ( .A(DP_OP_422J2_124_3477_n237), .B(
        DP_OP_422J2_124_3477_n212), .CI(DP_OP_422J2_124_3477_n235), .CO(
        DP_OP_422J2_124_3477_n207), .S(DP_OP_422J2_124_3477_n208) );
  FADDX1_HVT DP_OP_422J2_124_3477_U199 ( .A(DP_OP_422J2_124_3477_n233), .B(
        DP_OP_422J2_124_3477_n210), .CI(DP_OP_422J2_124_3477_n231), .CO(
        DP_OP_422J2_124_3477_n205), .S(DP_OP_422J2_124_3477_n206) );
  FADDX1_HVT DP_OP_422J2_124_3477_U198 ( .A(DP_OP_422J2_124_3477_n208), .B(
        DP_OP_422J2_124_3477_n229), .CI(DP_OP_422J2_124_3477_n206), .CO(
        DP_OP_422J2_124_3477_n203), .S(DP_OP_422J2_124_3477_n204) );
  FADDX1_HVT DP_OP_422J2_124_3477_U197 ( .A(DP_OP_422J2_124_3477_n227), .B(
        DP_OP_422J2_124_3477_n225), .CI(DP_OP_422J2_124_3477_n204), .CO(
        DP_OP_422J2_124_3477_n201), .S(DP_OP_422J2_124_3477_n202) );
  FADDX1_HVT DP_OP_422J2_124_3477_U196 ( .A(DP_OP_422J2_124_3477_n1775), .B(
        DP_OP_422J2_124_3477_n221), .CI(DP_OP_422J2_124_3477_n219), .CO(
        DP_OP_422J2_124_3477_n199), .S(DP_OP_422J2_124_3477_n200) );
  FADDX1_HVT DP_OP_422J2_124_3477_U195 ( .A(DP_OP_422J2_124_3477_n217), .B(
        DP_OP_422J2_124_3477_n200), .CI(DP_OP_422J2_124_3477_n215), .CO(
        DP_OP_422J2_124_3477_n197), .S(DP_OP_422J2_124_3477_n198) );
  FADDX1_HVT DP_OP_422J2_124_3477_U194 ( .A(DP_OP_422J2_124_3477_n213), .B(
        DP_OP_422J2_124_3477_n211), .CI(DP_OP_422J2_124_3477_n198), .CO(
        DP_OP_422J2_124_3477_n195), .S(DP_OP_422J2_124_3477_n196) );
  FADDX1_HVT DP_OP_422J2_124_3477_U193 ( .A(DP_OP_422J2_124_3477_n209), .B(
        DP_OP_422J2_124_3477_n196), .CI(DP_OP_422J2_124_3477_n207), .CO(
        DP_OP_422J2_124_3477_n193), .S(DP_OP_422J2_124_3477_n194) );
  FADDX1_HVT DP_OP_422J2_124_3477_U192 ( .A(DP_OP_422J2_124_3477_n205), .B(
        DP_OP_422J2_124_3477_n194), .CI(DP_OP_422J2_124_3477_n203), .CO(
        DP_OP_422J2_124_3477_n191), .S(DP_OP_422J2_124_3477_n192) );
  FADDX1_HVT DP_OP_422J2_124_3477_U190 ( .A(DP_OP_422J2_124_3477_n190), .B(
        DP_OP_422J2_124_3477_n199), .CI(DP_OP_422J2_124_3477_n197), .CO(
        DP_OP_422J2_124_3477_n187), .S(DP_OP_422J2_124_3477_n188) );
  FADDX1_HVT DP_OP_422J2_124_3477_U189 ( .A(DP_OP_422J2_124_3477_n188), .B(
        DP_OP_422J2_124_3477_n195), .CI(DP_OP_422J2_124_3477_n193), .CO(
        DP_OP_422J2_124_3477_n185), .S(DP_OP_422J2_124_3477_n186) );
  FADDX1_HVT DP_OP_422J2_124_3477_U188 ( .A(DP_OP_422J2_124_3477_n1774), .B(
        DP_OP_422J2_124_3477_n189), .CI(DP_OP_422J2_124_3477_n187), .CO(
        DP_OP_422J2_124_3477_n183), .S(DP_OP_422J2_124_3477_n184) );
  FADDX1_HVT DP_OP_422J2_124_3477_U171 ( .A(DP_OP_422J2_124_3477_n1754), .B(
        DP_OP_422J2_124_3477_n1752), .CI(DP_OP_422J2_124_3477_n1750), .CO(
        DP_OP_422J2_124_3477_n131), .S(n_conv2_sum_a[0]) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U170 ( .A1(DP_OP_422J2_124_3477_n1688), 
        .A2(DP_OP_422J2_124_3477_n1690), .Y(DP_OP_422J2_124_3477_n130) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U169 ( .A1(DP_OP_422J2_124_3477_n1690), .A2(
        DP_OP_422J2_124_3477_n1688), .Y(DP_OP_422J2_124_3477_n129) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U163 ( .A1(DP_OP_422J2_124_3477_n1582), 
        .A2(DP_OP_422J2_124_3477_n1584), .Y(DP_OP_422J2_124_3477_n127) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U155 ( .A1(DP_OP_422J2_124_3477_n1428), 
        .A2(DP_OP_422J2_124_3477_n1430), .Y(DP_OP_422J2_124_3477_n122) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U154 ( .A1(DP_OP_422J2_124_3477_n1430), .A2(
        DP_OP_422J2_124_3477_n1428), .Y(DP_OP_422J2_124_3477_n121) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U149 ( .A1(DP_OP_422J2_124_3477_n1252), 
        .A2(DP_OP_422J2_124_3477_n1254), .Y(DP_OP_422J2_124_3477_n119) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U141 ( .A1(DP_OP_422J2_124_3477_n1064), 
        .A2(DP_OP_422J2_124_3477_n1066), .Y(DP_OP_422J2_124_3477_n114) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U140 ( .A1(DP_OP_422J2_124_3477_n1066), .A2(
        DP_OP_422J2_124_3477_n1064), .Y(DP_OP_422J2_124_3477_n113) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U135 ( .A1(DP_OP_422J2_124_3477_n870), .A2(
        DP_OP_422J2_124_3477_n872), .Y(DP_OP_422J2_124_3477_n111) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U127 ( .A1(DP_OP_422J2_124_3477_n674), .A2(
        DP_OP_422J2_124_3477_n869), .Y(DP_OP_422J2_124_3477_n106) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U126 ( .A1(DP_OP_422J2_124_3477_n869), .A2(
        DP_OP_422J2_124_3477_n674), .Y(DP_OP_422J2_124_3477_n105) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U120 ( .A1(DP_OP_422J2_124_3477_n500), .A2(
        DP_OP_422J2_124_3477_n673), .Y(DP_OP_422J2_124_3477_n102) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U119 ( .A1(DP_OP_422J2_124_3477_n673), .A2(
        DP_OP_422J2_124_3477_n500), .Y(DP_OP_422J2_124_3477_n101) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U114 ( .A1(DP_OP_422J2_124_3477_n364), .A2(
        DP_OP_422J2_124_3477_n499), .Y(DP_OP_422J2_124_3477_n99) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U113 ( .A1(DP_OP_422J2_124_3477_n499), .A2(
        DP_OP_422J2_124_3477_n364), .Y(DP_OP_422J2_124_3477_n98) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U105 ( .A1(DP_OP_422J2_124_3477_n270), .A2(
        DP_OP_422J2_124_3477_n363), .Y(DP_OP_422J2_124_3477_n93) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U104 ( .A1(DP_OP_422J2_124_3477_n363), .A2(
        DP_OP_422J2_124_3477_n270), .Y(DP_OP_422J2_124_3477_n92) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U97 ( .A1(DP_OP_422J2_124_3477_n224), .A2(
        DP_OP_422J2_124_3477_n269), .Y(DP_OP_422J2_124_3477_n88) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U96 ( .A1(DP_OP_422J2_124_3477_n269), .A2(
        DP_OP_422J2_124_3477_n224), .Y(DP_OP_422J2_124_3477_n87) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U92 ( .A1(DP_OP_422J2_124_3477_n87), .A2(
        DP_OP_422J2_124_3477_n92), .Y(DP_OP_422J2_124_3477_n85) );
  AOI21X1_HVT DP_OP_422J2_124_3477_U91 ( .A1(DP_OP_422J2_124_3477_n94), .A2(
        DP_OP_422J2_124_3477_n85), .A3(DP_OP_422J2_124_3477_n86), .Y(
        DP_OP_422J2_124_3477_n84) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U89 ( .A1(DP_OP_422J2_124_3477_n202), .A2(
        DP_OP_422J2_124_3477_n223), .Y(DP_OP_422J2_124_3477_n83) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U88 ( .A1(DP_OP_422J2_124_3477_n223), .A2(
        DP_OP_422J2_124_3477_n202), .Y(DP_OP_422J2_124_3477_n82) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U83 ( .A1(DP_OP_422J2_124_3477_n201), .A2(
        DP_OP_422J2_124_3477_n192), .Y(DP_OP_422J2_124_3477_n80) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U82 ( .A1(DP_OP_422J2_124_3477_n192), .A2(
        DP_OP_422J2_124_3477_n201), .Y(DP_OP_422J2_124_3477_n79) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U78 ( .A1(DP_OP_422J2_124_3477_n79), .A2(
        DP_OP_422J2_124_3477_n82), .Y(DP_OP_422J2_124_3477_n77) );
  AOI21X1_HVT DP_OP_422J2_124_3477_U77 ( .A1(DP_OP_422J2_124_3477_n86), .A2(
        DP_OP_422J2_124_3477_n77), .A3(DP_OP_422J2_124_3477_n78), .Y(
        DP_OP_422J2_124_3477_n76) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U76 ( .A1(DP_OP_422J2_124_3477_n85), .A2(
        DP_OP_422J2_124_3477_n77), .Y(DP_OP_422J2_124_3477_n75) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U72 ( .A1(DP_OP_422J2_124_3477_n191), .A2(
        DP_OP_422J2_124_3477_n186), .Y(DP_OP_422J2_124_3477_n68) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U62 ( .A1(DP_OP_422J2_124_3477_n185), .A2(
        DP_OP_422J2_124_3477_n184), .Y(DP_OP_422J2_124_3477_n65) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U61 ( .A1(DP_OP_422J2_124_3477_n184), .A2(
        DP_OP_422J2_124_3477_n185), .Y(DP_OP_422J2_124_3477_n64) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U54 ( .A1(DP_OP_422J2_124_3477_n183), .A2(
        DP_OP_422J2_124_3477_n182), .Y(DP_OP_422J2_124_3477_n60) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U53 ( .A1(DP_OP_422J2_124_3477_n182), .A2(
        DP_OP_422J2_124_3477_n183), .Y(DP_OP_422J2_124_3477_n59) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U49 ( .A1(DP_OP_422J2_124_3477_n59), .A2(
        DP_OP_422J2_124_3477_n64), .Y(DP_OP_422J2_124_3477_n57) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U47 ( .A1(DP_OP_422J2_124_3477_n69), .A2(
        DP_OP_422J2_124_3477_n57), .Y(DP_OP_422J2_124_3477_n55) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U44 ( .A1(DP_OP_422J2_124_3477_n180), .A2(
        DP_OP_422J2_124_3477_n181), .Y(DP_OP_422J2_124_3477_n53) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U43 ( .A1(DP_OP_422J2_124_3477_n181), .A2(
        DP_OP_422J2_124_3477_n180), .Y(DP_OP_422J2_124_3477_n52) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U39 ( .A1(DP_OP_422J2_124_3477_n52), .A2(
        DP_OP_422J2_124_3477_n55), .Y(DP_OP_422J2_124_3477_n50) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U34 ( .A1(DP_OP_422J2_124_3477_n178), .A2(
        DP_OP_422J2_124_3477_n179), .Y(DP_OP_422J2_124_3477_n46) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U27 ( .A1(DP_OP_422J2_124_3477_n50), .A2(
        DP_OP_422J2_124_3477_n45), .Y(DP_OP_422J2_124_3477_n41) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U24 ( .A1(DP_OP_422J2_124_3477_n176), .A2(
        DP_OP_422J2_124_3477_n177), .Y(DP_OP_422J2_124_3477_n39) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U23 ( .A1(DP_OP_422J2_124_3477_n177), .A2(
        DP_OP_422J2_124_3477_n176), .Y(DP_OP_422J2_124_3477_n38) );
  FADDX1_HVT DP_OP_422J2_124_3477_U15 ( .A(DP_OP_422J2_124_3477_n175), .B(
        DP_OP_422J2_124_3477_n174), .CI(DP_OP_422J2_124_3477_n35), .CO(
        DP_OP_422J2_124_3477_n34), .S(n_conv2_sum_a[20]) );
  FADDX1_HVT DP_OP_422J2_124_3477_U14 ( .A(DP_OP_422J2_124_3477_n173), .B(
        DP_OP_422J2_124_3477_n172), .CI(DP_OP_422J2_124_3477_n34), .CO(
        DP_OP_422J2_124_3477_n33), .S(n_conv2_sum_a[21]) );
  FADDX1_HVT DP_OP_422J2_124_3477_U13 ( .A(DP_OP_422J2_124_3477_n171), .B(
        DP_OP_422J2_124_3477_n170), .CI(DP_OP_422J2_124_3477_n33), .CO(
        DP_OP_422J2_124_3477_n32), .S(n_conv2_sum_a[22]) );
  FADDX1_HVT DP_OP_422J2_124_3477_U12 ( .A(DP_OP_422J2_124_3477_n169), .B(
        DP_OP_422J2_124_3477_n168), .CI(DP_OP_422J2_124_3477_n32), .CO(
        DP_OP_422J2_124_3477_n31), .S(n_conv2_sum_a[23]) );
  FADDX1_HVT DP_OP_422J2_124_3477_U11 ( .A(DP_OP_422J2_124_3477_n167), .B(
        DP_OP_422J2_124_3477_n166), .CI(DP_OP_422J2_124_3477_n31), .CO(
        DP_OP_422J2_124_3477_n30), .S(n_conv2_sum_a[24]) );
  FADDX1_HVT DP_OP_422J2_124_3477_U10 ( .A(DP_OP_422J2_124_3477_n165), .B(
        DP_OP_422J2_124_3477_n164), .CI(DP_OP_422J2_124_3477_n30), .CO(
        DP_OP_422J2_124_3477_n29), .S(n_conv2_sum_a[25]) );
  FADDX1_HVT DP_OP_422J2_124_3477_U9 ( .A(DP_OP_422J2_124_3477_n163), .B(
        DP_OP_422J2_124_3477_n162), .CI(DP_OP_422J2_124_3477_n29), .CO(
        DP_OP_422J2_124_3477_n28), .S(n_conv2_sum_a[26]) );
  FADDX1_HVT DP_OP_422J2_124_3477_U8 ( .A(DP_OP_422J2_124_3477_n161), .B(
        DP_OP_422J2_124_3477_n160), .CI(DP_OP_422J2_124_3477_n28), .CO(
        DP_OP_422J2_124_3477_n27), .S(n_conv2_sum_a[27]) );
  FADDX1_HVT DP_OP_422J2_124_3477_U7 ( .A(DP_OP_422J2_124_3477_n159), .B(
        DP_OP_422J2_124_3477_n158), .CI(DP_OP_422J2_124_3477_n27), .CO(
        DP_OP_422J2_124_3477_n26), .S(n_conv2_sum_a[28]) );
  FADDX1_HVT DP_OP_422J2_124_3477_U6 ( .A(DP_OP_422J2_124_3477_n157), .B(
        DP_OP_422J2_124_3477_n156), .CI(DP_OP_422J2_124_3477_n26), .CO(
        DP_OP_422J2_124_3477_n25), .S(n_conv2_sum_a[29]) );
  FADDX1_HVT DP_OP_422J2_124_3477_U5 ( .A(DP_OP_422J2_124_3477_n155), .B(
        DP_OP_422J2_124_3477_n154), .CI(DP_OP_422J2_124_3477_n25), .CO(
        DP_OP_422J2_124_3477_n24), .S(n_conv2_sum_a[30]) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2124 ( .A1(DP_OP_423J2_125_3477_n2903), 
        .A2(DP_OP_423J2_125_3477_n2913), .Y(DP_OP_423J2_125_3477_n2895) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2123 ( .A1(DP_OP_423J2_125_3477_n2902), .A2(
        DP_OP_423J2_125_3477_n2913), .Y(DP_OP_423J2_125_3477_n2894) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2115 ( .A1(DP_OP_423J2_125_3477_n2902), .A2(
        DP_OP_424J2_126_3477_n2917), .Y(DP_OP_423J2_125_3477_n2886) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2108 ( .A1(DP_OP_423J2_125_3477_n2903), 
        .A2(DP_OP_423J2_125_3477_n2911), .Y(DP_OP_423J2_125_3477_n2879) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2107 ( .A1(DP_OP_423J2_125_3477_n2902), .A2(
        DP_OP_423J2_125_3477_n2911), .Y(DP_OP_423J2_125_3477_n2878) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2106 ( .A1(DP_OP_423J2_125_3477_n2909), .A2(
        DP_OP_423J2_125_3477_n2910), .Y(DP_OP_423J2_125_3477_n2877) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2105 ( .A1(DP_OP_423J2_125_3477_n2908), .A2(
        DP_OP_423J2_125_3477_n2910), .Y(DP_OP_423J2_125_3477_n2876) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2104 ( .A1(DP_OP_423J2_125_3477_n2907), .A2(
        DP_OP_423J2_125_3477_n2910), .Y(DP_OP_423J2_125_3477_n2875) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2103 ( .A1(DP_OP_423J2_125_3477_n2906), .A2(
        DP_OP_423J2_125_3477_n2910), .Y(DP_OP_423J2_125_3477_n2874) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2102 ( .A1(DP_OP_425J2_127_3477_n1945), .A2(
        DP_OP_423J2_125_3477_n2910), .Y(DP_OP_423J2_125_3477_n2873) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2101 ( .A1(DP_OP_423J2_125_3477_n2904), .A2(
        DP_OP_423J2_125_3477_n2910), .Y(DP_OP_423J2_125_3477_n2872) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2100 ( .A1(DP_OP_423J2_125_3477_n2903), .A2(
        DP_OP_423J2_125_3477_n2910), .Y(DP_OP_423J2_125_3477_n2871) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2099 ( .A1(DP_OP_423J2_125_3477_n2902), 
        .A2(DP_OP_423J2_125_3477_n2910), .Y(DP_OP_423J2_125_3477_n2870) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2080 ( .A1(DP_OP_423J2_125_3477_n2859), 
        .A2(DP_OP_423J2_125_3477_n2869), .Y(DP_OP_423J2_125_3477_n2851) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2079 ( .A1(DP_OP_422J2_124_3477_n1854), .A2(
        DP_OP_423J2_125_3477_n2869), .Y(DP_OP_423J2_125_3477_n2850) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2072 ( .A1(DP_OP_423J2_125_3477_n2859), 
        .A2(DP_OP_423J2_125_3477_n2868), .Y(DP_OP_423J2_125_3477_n2843) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2071 ( .A1(DP_OP_422J2_124_3477_n1854), .A2(
        DP_OP_423J2_125_3477_n2868), .Y(DP_OP_423J2_125_3477_n2842) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2064 ( .A1(DP_OP_423J2_125_3477_n2859), 
        .A2(DP_OP_423J2_125_3477_n2867), .Y(DP_OP_423J2_125_3477_n2835) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2063 ( .A1(DP_OP_422J2_124_3477_n1854), .A2(
        DP_OP_423J2_125_3477_n2867), .Y(DP_OP_423J2_125_3477_n2834) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2062 ( .A1(DP_OP_423J2_125_3477_n2865), .A2(
        DP_OP_423J2_125_3477_n2866), .Y(DP_OP_423J2_125_3477_n2833) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2061 ( .A1(DP_OP_423J2_125_3477_n2864), .A2(
        DP_OP_423J2_125_3477_n2866), .Y(DP_OP_423J2_125_3477_n2832) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2060 ( .A1(DP_OP_425J2_127_3477_n1991), .A2(
        DP_OP_423J2_125_3477_n2866), .Y(DP_OP_423J2_125_3477_n2831) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2059 ( .A1(DP_OP_425J2_127_3477_n1990), .A2(
        DP_OP_423J2_125_3477_n2866), .Y(DP_OP_423J2_125_3477_n2830) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2058 ( .A1(DP_OP_423J2_125_3477_n2861), .A2(
        DP_OP_423J2_125_3477_n2866), .Y(DP_OP_423J2_125_3477_n2829) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2057 ( .A1(DP_OP_423J2_125_3477_n2860), .A2(
        DP_OP_423J2_125_3477_n2866), .Y(DP_OP_423J2_125_3477_n2828) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2056 ( .A1(DP_OP_423J2_125_3477_n2859), .A2(
        DP_OP_423J2_125_3477_n2866), .Y(DP_OP_423J2_125_3477_n2827) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2055 ( .A1(DP_OP_424J2_126_3477_n2775), 
        .A2(DP_OP_423J2_125_3477_n2866), .Y(DP_OP_423J2_125_3477_n2826) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2036 ( .A1(DP_OP_422J2_124_3477_n1899), 
        .A2(DP_OP_424J2_126_3477_n2830), .Y(DP_OP_423J2_125_3477_n2807) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2035 ( .A1(DP_OP_424J2_126_3477_n2731), .A2(
        DP_OP_424J2_126_3477_n2830), .Y(DP_OP_423J2_125_3477_n2806) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2027 ( .A1(DP_OP_422J2_124_3477_n1898), .A2(
        DP_OP_423J2_125_3477_n2824), .Y(DP_OP_423J2_125_3477_n2798) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2020 ( .A1(DP_OP_424J2_126_3477_n2732), 
        .A2(DP_OP_423J2_125_3477_n2823), .Y(DP_OP_423J2_125_3477_n2791) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2019 ( .A1(DP_OP_422J2_124_3477_n1898), .A2(
        DP_OP_423J2_125_3477_n2823), .Y(DP_OP_423J2_125_3477_n2790) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2018 ( .A1(DP_OP_424J2_126_3477_n2738), .A2(
        DP_OP_422J2_124_3477_n2827), .Y(DP_OP_423J2_125_3477_n2789) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2017 ( .A1(DP_OP_424J2_126_3477_n2737), .A2(
        DP_OP_424J2_126_3477_n2827), .Y(DP_OP_423J2_125_3477_n2788) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2016 ( .A1(DP_OP_424J2_126_3477_n2736), .A2(
        DP_OP_425J2_127_3477_n2827), .Y(DP_OP_423J2_125_3477_n2787) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2015 ( .A1(DP_OP_422J2_124_3477_n1902), .A2(
        DP_OP_425J2_127_3477_n2827), .Y(DP_OP_423J2_125_3477_n2786) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2014 ( .A1(DP_OP_424J2_126_3477_n2734), .A2(
        DP_OP_424J2_126_3477_n2827), .Y(DP_OP_423J2_125_3477_n2785) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2013 ( .A1(DP_OP_422J2_124_3477_n1900), .A2(
        DP_OP_422J2_124_3477_n2827), .Y(DP_OP_423J2_125_3477_n2784) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2012 ( .A1(DP_OP_424J2_126_3477_n2732), .A2(
        DP_OP_425J2_127_3477_n2827), .Y(DP_OP_423J2_125_3477_n2783) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2011 ( .A1(DP_OP_422J2_124_3477_n1898), 
        .A2(DP_OP_422J2_124_3477_n2827), .Y(DP_OP_423J2_125_3477_n2782) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1992 ( .A1(DP_OP_422J2_124_3477_n1943), 
        .A2(DP_OP_423J2_125_3477_n2781), .Y(DP_OP_423J2_125_3477_n2763) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1991 ( .A1(DP_OP_423J2_125_3477_n2770), .A2(
        DP_OP_423J2_125_3477_n2781), .Y(DP_OP_423J2_125_3477_n2762) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1984 ( .A1(DP_OP_425J2_127_3477_n2075), 
        .A2(DP_OP_424J2_126_3477_n2785), .Y(DP_OP_423J2_125_3477_n2755) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1983 ( .A1(DP_OP_423J2_125_3477_n2770), .A2(
        DP_OP_424J2_126_3477_n2785), .Y(DP_OP_423J2_125_3477_n2754) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1976 ( .A1(DP_OP_422J2_124_3477_n1943), 
        .A2(DP_OP_423J2_125_3477_n2779), .Y(DP_OP_423J2_125_3477_n2747) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1975 ( .A1(DP_OP_423J2_125_3477_n2770), .A2(
        DP_OP_423J2_125_3477_n2779), .Y(DP_OP_423J2_125_3477_n2746) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1974 ( .A1(DP_OP_423J2_125_3477_n2777), .A2(
        DP_OP_423J2_125_3477_n2778), .Y(DP_OP_423J2_125_3477_n2745) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1973 ( .A1(DP_OP_423J2_125_3477_n2776), .A2(
        DP_OP_423J2_125_3477_n2778), .Y(DP_OP_423J2_125_3477_n2744) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1972 ( .A1(DP_OP_423J2_125_3477_n2775), .A2(
        DP_OP_423J2_125_3477_n2778), .Y(DP_OP_423J2_125_3477_n2743) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1971 ( .A1(DP_OP_425J2_127_3477_n2078), .A2(
        DP_OP_423J2_125_3477_n2778), .Y(DP_OP_423J2_125_3477_n2742) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1970 ( .A1(DP_OP_422J2_124_3477_n1945), .A2(
        DP_OP_423J2_125_3477_n2778), .Y(DP_OP_423J2_125_3477_n2741) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1969 ( .A1(DP_OP_423J2_125_3477_n2772), .A2(
        DP_OP_423J2_125_3477_n2778), .Y(DP_OP_423J2_125_3477_n2740) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1968 ( .A1(DP_OP_422J2_124_3477_n1943), .A2(
        DP_OP_423J2_125_3477_n2778), .Y(DP_OP_423J2_125_3477_n2739) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1967 ( .A1(DP_OP_423J2_125_3477_n2770), 
        .A2(DP_OP_423J2_125_3477_n2778), .Y(DP_OP_423J2_125_3477_n2738) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1949 ( .A1(DP_OP_425J2_127_3477_n2120), 
        .A2(DP_OP_423J2_125_3477_n2737), .Y(DP_OP_423J2_125_3477_n2720) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1948 ( .A1(DP_OP_425J2_127_3477_n2119), 
        .A2(DP_OP_423J2_125_3477_n2737), .Y(DP_OP_423J2_125_3477_n2719) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1947 ( .A1(DP_OP_423J2_125_3477_n2726), .A2(
        DP_OP_423J2_125_3477_n2737), .Y(DP_OP_423J2_125_3477_n2718) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1939 ( .A1(DP_OP_423J2_125_3477_n2726), .A2(
        DP_OP_424J2_126_3477_n2741), .Y(DP_OP_423J2_125_3477_n2710) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1931 ( .A1(DP_OP_423J2_125_3477_n2726), .A2(
        DP_OP_424J2_126_3477_n2740), .Y(DP_OP_423J2_125_3477_n2702) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1930 ( .A1(DP_OP_423J2_125_3477_n2733), .A2(
        DP_OP_423J2_125_3477_n2734), .Y(DP_OP_423J2_125_3477_n1574) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1929 ( .A1(DP_OP_423J2_125_3477_n2732), .A2(
        DP_OP_423J2_125_3477_n2734), .Y(DP_OP_423J2_125_3477_n2701) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1928 ( .A1(DP_OP_423J2_125_3477_n2731), .A2(
        DP_OP_423J2_125_3477_n2734), .Y(DP_OP_423J2_125_3477_n2700) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1927 ( .A1(DP_OP_423J2_125_3477_n2730), .A2(
        DP_OP_423J2_125_3477_n2734), .Y(DP_OP_423J2_125_3477_n2699) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1926 ( .A1(DP_OP_423J2_125_3477_n2729), .A2(
        DP_OP_423J2_125_3477_n2734), .Y(DP_OP_423J2_125_3477_n2698) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1925 ( .A1(DP_OP_422J2_124_3477_n1988), .A2(
        DP_OP_423J2_125_3477_n2734), .Y(DP_OP_423J2_125_3477_n666) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1924 ( .A1(DP_OP_424J2_126_3477_n2644), .A2(
        DP_OP_423J2_125_3477_n2734), .Y(DP_OP_423J2_125_3477_n2697) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1923 ( .A1(DP_OP_423J2_125_3477_n2726), 
        .A2(DP_OP_423J2_125_3477_n2734), .Y(DP_OP_423J2_125_3477_n356) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1905 ( .A1(DP_OP_425J2_127_3477_n2164), 
        .A2(DP_OP_423J2_125_3477_n2696), .Y(DP_OP_423J2_125_3477_n2679) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1904 ( .A1(DP_OP_425J2_127_3477_n2163), 
        .A2(DP_OP_423J2_125_3477_n2696), .Y(DP_OP_423J2_125_3477_n2678) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1903 ( .A1(DP_OP_425J2_127_3477_n2162), .A2(
        DP_OP_423J2_125_3477_n2696), .Y(DP_OP_423J2_125_3477_n2677) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1896 ( .A1(DP_OP_425J2_127_3477_n2163), 
        .A2(DP_OP_423J2_125_3477_n2695), .Y(DP_OP_423J2_125_3477_n2670) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1895 ( .A1(DP_OP_425J2_127_3477_n2162), .A2(
        DP_OP_423J2_125_3477_n2695), .Y(DP_OP_423J2_125_3477_n2669) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1887 ( .A1(DP_OP_425J2_127_3477_n2162), .A2(
        DP_OP_422J2_124_3477_n2698), .Y(DP_OP_423J2_125_3477_n2661) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1886 ( .A1(DP_OP_425J2_127_3477_n2169), .A2(
        DP_OP_423J2_125_3477_n2693), .Y(DP_OP_423J2_125_3477_n2660) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1885 ( .A1(DP_OP_425J2_127_3477_n2168), .A2(
        DP_OP_423J2_125_3477_n2693), .Y(DP_OP_423J2_125_3477_n2659) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1884 ( .A1(DP_OP_423J2_125_3477_n2690), .A2(
        DP_OP_423J2_125_3477_n2693), .Y(DP_OP_423J2_125_3477_n2658) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1883 ( .A1(DP_OP_425J2_127_3477_n2166), .A2(
        DP_OP_423J2_125_3477_n2693), .Y(DP_OP_423J2_125_3477_n2657) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1882 ( .A1(DP_OP_423J2_125_3477_n2688), .A2(
        DP_OP_423J2_125_3477_n2693), .Y(DP_OP_423J2_125_3477_n2656) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1881 ( .A1(DP_OP_425J2_127_3477_n2164), .A2(
        DP_OP_423J2_125_3477_n2693), .Y(DP_OP_423J2_125_3477_n2655) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1880 ( .A1(DP_OP_425J2_127_3477_n2163), .A2(
        DP_OP_423J2_125_3477_n2693), .Y(DP_OP_423J2_125_3477_n2654) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1879 ( .A1(DP_OP_425J2_127_3477_n2162), 
        .A2(DP_OP_423J2_125_3477_n2693), .Y(DP_OP_423J2_125_3477_n2653) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1860 ( .A1(DP_OP_423J2_125_3477_n2642), 
        .A2(DP_OP_422J2_124_3477_n2656), .Y(DP_OP_423J2_125_3477_n2634) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1859 ( .A1(DP_OP_422J2_124_3477_n2073), .A2(
        DP_OP_424J2_126_3477_n2654), .Y(DP_OP_423J2_125_3477_n2633) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1852 ( .A1(DP_OP_423J2_125_3477_n2642), 
        .A2(DP_OP_423J2_125_3477_n2651), .Y(DP_OP_423J2_125_3477_n2626) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1851 ( .A1(DP_OP_422J2_124_3477_n2073), .A2(
        DP_OP_423J2_125_3477_n2651), .Y(DP_OP_423J2_125_3477_n2625) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1844 ( .A1(DP_OP_423J2_125_3477_n2642), 
        .A2(DP_OP_425J2_127_3477_n2652), .Y(DP_OP_423J2_125_3477_n2618) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1843 ( .A1(DP_OP_424J2_126_3477_n2555), .A2(
        DP_OP_424J2_126_3477_n2652), .Y(DP_OP_423J2_125_3477_n2617) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1842 ( .A1(DP_OP_423J2_125_3477_n2648), .A2(
        DP_OP_423J2_125_3477_n2649), .Y(DP_OP_423J2_125_3477_n2616) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1841 ( .A1(DP_OP_423J2_125_3477_n2647), .A2(
        DP_OP_423J2_125_3477_n2649), .Y(DP_OP_423J2_125_3477_n2615) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1840 ( .A1(DP_OP_423J2_125_3477_n2646), .A2(
        DP_OP_423J2_125_3477_n2649), .Y(DP_OP_423J2_125_3477_n2614) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1839 ( .A1(DP_OP_423J2_125_3477_n2645), .A2(
        DP_OP_423J2_125_3477_n2649), .Y(DP_OP_423J2_125_3477_n2613) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1838 ( .A1(DP_OP_422J2_124_3477_n2076), .A2(
        DP_OP_423J2_125_3477_n2649), .Y(DP_OP_423J2_125_3477_n2612) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1837 ( .A1(DP_OP_423J2_125_3477_n2643), .A2(
        DP_OP_423J2_125_3477_n2649), .Y(DP_OP_423J2_125_3477_n2611) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1836 ( .A1(DP_OP_423J2_125_3477_n2642), .A2(
        DP_OP_423J2_125_3477_n2649), .Y(DP_OP_423J2_125_3477_n2610) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1835 ( .A1(DP_OP_424J2_126_3477_n2555), 
        .A2(DP_OP_423J2_125_3477_n2649), .Y(DP_OP_423J2_125_3477_n2609) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1817 ( .A1(DP_OP_423J2_125_3477_n2599), 
        .A2(DP_OP_424J2_126_3477_n2610), .Y(DP_OP_423J2_125_3477_n2591) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1816 ( .A1(DP_OP_424J2_126_3477_n2512), 
        .A2(DP_OP_424J2_126_3477_n2610), .Y(DP_OP_423J2_125_3477_n2590) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1815 ( .A1(DP_OP_422J2_124_3477_n2117), .A2(
        DP_OP_424J2_126_3477_n2610), .Y(DP_OP_423J2_125_3477_n2589) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1808 ( .A1(DP_OP_422J2_124_3477_n2118), 
        .A2(DP_OP_423J2_125_3477_n2607), .Y(DP_OP_423J2_125_3477_n2582) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1807 ( .A1(DP_OP_425J2_127_3477_n2250), .A2(
        DP_OP_423J2_125_3477_n2607), .Y(DP_OP_423J2_125_3477_n2581) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1800 ( .A1(DP_OP_424J2_126_3477_n2512), 
        .A2(n451), .Y(DP_OP_423J2_125_3477_n2574) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1799 ( .A1(DP_OP_422J2_124_3477_n2117), .A2(
        n451), .Y(DP_OP_423J2_125_3477_n2573) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1798 ( .A1(DP_OP_423J2_125_3477_n2604), .A2(
        DP_OP_423J2_125_3477_n2605), .Y(DP_OP_423J2_125_3477_n2572) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1797 ( .A1(DP_OP_423J2_125_3477_n2603), .A2(
        DP_OP_423J2_125_3477_n2605), .Y(DP_OP_423J2_125_3477_n2571) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1796 ( .A1(DP_OP_423J2_125_3477_n2602), .A2(
        DP_OP_423J2_125_3477_n2605), .Y(DP_OP_423J2_125_3477_n2570) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1795 ( .A1(DP_OP_423J2_125_3477_n2601), .A2(
        DP_OP_423J2_125_3477_n2605), .Y(DP_OP_423J2_125_3477_n2569) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1794 ( .A1(DP_OP_423J2_125_3477_n2600), .A2(
        DP_OP_423J2_125_3477_n2605), .Y(DP_OP_423J2_125_3477_n2568) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1793 ( .A1(DP_OP_423J2_125_3477_n2599), .A2(
        DP_OP_423J2_125_3477_n2605), .Y(DP_OP_423J2_125_3477_n2567) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1792 ( .A1(DP_OP_422J2_124_3477_n2118), .A2(
        DP_OP_423J2_125_3477_n2605), .Y(DP_OP_423J2_125_3477_n2566) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1791 ( .A1(DP_OP_425J2_127_3477_n2250), 
        .A2(DP_OP_423J2_125_3477_n2605), .Y(DP_OP_423J2_125_3477_n2565) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1772 ( .A1(DP_OP_423J2_125_3477_n2554), 
        .A2(DP_OP_424J2_126_3477_n2566), .Y(DP_OP_423J2_125_3477_n2546) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1771 ( .A1(DP_OP_423J2_125_3477_n2553), .A2(
        DP_OP_425J2_127_3477_n2566), .Y(DP_OP_423J2_125_3477_n2545) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1764 ( .A1(DP_OP_423J2_125_3477_n2554), 
        .A2(DP_OP_422J2_124_3477_n2567), .Y(DP_OP_423J2_125_3477_n2538) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1763 ( .A1(DP_OP_423J2_125_3477_n2553), .A2(
        DP_OP_425J2_127_3477_n2565), .Y(DP_OP_423J2_125_3477_n2537) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1755 ( .A1(DP_OP_423J2_125_3477_n2553), .A2(
        DP_OP_423J2_125_3477_n2562), .Y(DP_OP_423J2_125_3477_n2529) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1754 ( .A1(DP_OP_422J2_124_3477_n2168), .A2(
        DP_OP_423J2_125_3477_n2561), .Y(DP_OP_423J2_125_3477_n2528) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1753 ( .A1(DP_OP_423J2_125_3477_n2559), .A2(
        DP_OP_423J2_125_3477_n2561), .Y(DP_OP_423J2_125_3477_n2527) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1752 ( .A1(DP_OP_423J2_125_3477_n2558), .A2(
        DP_OP_423J2_125_3477_n2561), .Y(DP_OP_423J2_125_3477_n2526) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1751 ( .A1(DP_OP_422J2_124_3477_n2165), .A2(
        DP_OP_423J2_125_3477_n2561), .Y(DP_OP_423J2_125_3477_n2525) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1750 ( .A1(DP_OP_422J2_124_3477_n2164), .A2(
        DP_OP_423J2_125_3477_n2561), .Y(DP_OP_423J2_125_3477_n2524) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1749 ( .A1(DP_OP_422J2_124_3477_n2163), .A2(
        DP_OP_423J2_125_3477_n2561), .Y(DP_OP_423J2_125_3477_n2523) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1748 ( .A1(DP_OP_423J2_125_3477_n2554), .A2(
        DP_OP_423J2_125_3477_n2561), .Y(DP_OP_423J2_125_3477_n2522) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1747 ( .A1(DP_OP_423J2_125_3477_n2553), 
        .A2(DP_OP_423J2_125_3477_n2561), .Y(DP_OP_423J2_125_3477_n2521) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1728 ( .A1(DP_OP_423J2_125_3477_n2510), 
        .A2(DP_OP_423J2_125_3477_n2520), .Y(DP_OP_423J2_125_3477_n2502) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1727 ( .A1(DP_OP_423J2_125_3477_n2509), .A2(
        DP_OP_423J2_125_3477_n2520), .Y(DP_OP_423J2_125_3477_n2501) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1719 ( .A1(DP_OP_423J2_125_3477_n2509), .A2(
        DP_OP_423J2_125_3477_n2519), .Y(DP_OP_423J2_125_3477_n2493) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1712 ( .A1(DP_OP_423J2_125_3477_n2510), 
        .A2(n444), .Y(DP_OP_423J2_125_3477_n2486) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1711 ( .A1(DP_OP_423J2_125_3477_n2509), .A2(
        n444), .Y(DP_OP_423J2_125_3477_n2485) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1710 ( .A1(DP_OP_423J2_125_3477_n2516), .A2(
        DP_OP_423J2_125_3477_n2517), .Y(DP_OP_423J2_125_3477_n2484) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1709 ( .A1(DP_OP_423J2_125_3477_n2515), .A2(
        DP_OP_423J2_125_3477_n2517), .Y(DP_OP_423J2_125_3477_n2483) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1708 ( .A1(DP_OP_422J2_124_3477_n2210), .A2(
        DP_OP_423J2_125_3477_n2517), .Y(DP_OP_423J2_125_3477_n2482) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1707 ( .A1(DP_OP_425J2_127_3477_n2342), .A2(
        DP_OP_423J2_125_3477_n2517), .Y(DP_OP_423J2_125_3477_n2481) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1706 ( .A1(DP_OP_425J2_127_3477_n2341), .A2(
        DP_OP_423J2_125_3477_n2517), .Y(DP_OP_423J2_125_3477_n2480) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1705 ( .A1(DP_OP_422J2_124_3477_n2207), .A2(
        DP_OP_423J2_125_3477_n2517), .Y(DP_OP_423J2_125_3477_n2479) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1704 ( .A1(DP_OP_423J2_125_3477_n2510), .A2(
        DP_OP_423J2_125_3477_n2517), .Y(DP_OP_423J2_125_3477_n2478) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1703 ( .A1(DP_OP_423J2_125_3477_n2509), 
        .A2(DP_OP_423J2_125_3477_n2517), .Y(DP_OP_423J2_125_3477_n2477) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1684 ( .A1(DP_OP_423J2_125_3477_n2466), 
        .A2(DP_OP_423J2_125_3477_n2476), .Y(DP_OP_423J2_125_3477_n2458) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1683 ( .A1(DP_OP_423J2_125_3477_n2465), .A2(
        DP_OP_423J2_125_3477_n2476), .Y(DP_OP_423J2_125_3477_n2457) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1676 ( .A1(DP_OP_423J2_125_3477_n2466), 
        .A2(DP_OP_423J2_125_3477_n2475), .Y(DP_OP_423J2_125_3477_n2450) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1675 ( .A1(DP_OP_423J2_125_3477_n2465), .A2(
        DP_OP_423J2_125_3477_n2475), .Y(DP_OP_423J2_125_3477_n2449) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1668 ( .A1(DP_OP_423J2_125_3477_n2466), 
        .A2(DP_OP_423J2_125_3477_n2474), .Y(DP_OP_423J2_125_3477_n2442) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1667 ( .A1(DP_OP_423J2_125_3477_n2465), .A2(
        DP_OP_423J2_125_3477_n2474), .Y(DP_OP_423J2_125_3477_n2441) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1666 ( .A1(DP_OP_423J2_125_3477_n2472), .A2(
        DP_OP_424J2_126_3477_n2475), .Y(DP_OP_423J2_125_3477_n2440) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1665 ( .A1(DP_OP_423J2_125_3477_n2471), .A2(
        DP_OP_424J2_126_3477_n2475), .Y(DP_OP_423J2_125_3477_n2439) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1664 ( .A1(DP_OP_423J2_125_3477_n2470), .A2(
        DP_OP_425J2_127_3477_n2475), .Y(DP_OP_423J2_125_3477_n2438) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1663 ( .A1(DP_OP_423J2_125_3477_n2469), .A2(
        DP_OP_424J2_126_3477_n2475), .Y(DP_OP_423J2_125_3477_n2437) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1662 ( .A1(DP_OP_423J2_125_3477_n2468), .A2(
        DP_OP_424J2_126_3477_n2475), .Y(DP_OP_423J2_125_3477_n2436) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1661 ( .A1(DP_OP_423J2_125_3477_n2467), .A2(
        DP_OP_422J2_124_3477_n2477), .Y(DP_OP_423J2_125_3477_n2435) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1660 ( .A1(DP_OP_423J2_125_3477_n2466), .A2(
        DP_OP_425J2_127_3477_n2475), .Y(DP_OP_423J2_125_3477_n2434) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1659 ( .A1(DP_OP_423J2_125_3477_n2465), 
        .A2(DP_OP_422J2_124_3477_n2477), .Y(DP_OP_423J2_125_3477_n2433) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1640 ( .A1(DP_OP_422J2_124_3477_n2294), 
        .A2(DP_OP_423J2_125_3477_n2432), .Y(DP_OP_423J2_125_3477_n2414) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1639 ( .A1(DP_OP_423J2_125_3477_n2421), .A2(
        DP_OP_423J2_125_3477_n2432), .Y(DP_OP_423J2_125_3477_n2413) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1631 ( .A1(DP_OP_423J2_125_3477_n2421), .A2(
        DP_OP_423J2_125_3477_n2431), .Y(DP_OP_423J2_125_3477_n2405) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1623 ( .A1(DP_OP_423J2_125_3477_n2421), .A2(
        DP_OP_423J2_125_3477_n2430), .Y(DP_OP_423J2_125_3477_n2397) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1622 ( .A1(DP_OP_423J2_125_3477_n2428), .A2(
        DP_OP_423J2_125_3477_n2429), .Y(DP_OP_423J2_125_3477_n2396) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1621 ( .A1(DP_OP_422J2_124_3477_n2299), .A2(
        DP_OP_423J2_125_3477_n2429), .Y(DP_OP_423J2_125_3477_n2395) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1620 ( .A1(DP_OP_422J2_124_3477_n2298), .A2(
        DP_OP_423J2_125_3477_n2429), .Y(DP_OP_423J2_125_3477_n2394) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1619 ( .A1(DP_OP_423J2_125_3477_n2425), .A2(
        DP_OP_423J2_125_3477_n2429), .Y(DP_OP_423J2_125_3477_n2393) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1618 ( .A1(DP_OP_423J2_125_3477_n2424), .A2(
        DP_OP_423J2_125_3477_n2429), .Y(DP_OP_423J2_125_3477_n2392) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1617 ( .A1(DP_OP_422J2_124_3477_n2295), .A2(
        DP_OP_423J2_125_3477_n2429), .Y(DP_OP_423J2_125_3477_n2391) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1616 ( .A1(DP_OP_422J2_124_3477_n2294), .A2(
        DP_OP_423J2_125_3477_n2429), .Y(DP_OP_423J2_125_3477_n2390) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1615 ( .A1(DP_OP_423J2_125_3477_n2421), 
        .A2(DP_OP_423J2_125_3477_n2429), .Y(DP_OP_423J2_125_3477_n2389) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1595 ( .A1(DP_OP_423J2_125_3477_n2377), .A2(
        DP_OP_423J2_125_3477_n2388), .Y(DP_OP_423J2_125_3477_n2369) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1588 ( .A1(DP_OP_422J2_124_3477_n2338), 
        .A2(DP_OP_423J2_125_3477_n2387), .Y(DP_OP_423J2_125_3477_n2362) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1587 ( .A1(DP_OP_423J2_125_3477_n2377), .A2(
        DP_OP_423J2_125_3477_n2387), .Y(DP_OP_423J2_125_3477_n2361) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1580 ( .A1(DP_OP_422J2_124_3477_n2338), 
        .A2(DP_OP_423J2_125_3477_n2386), .Y(DP_OP_423J2_125_3477_n2354) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1579 ( .A1(DP_OP_423J2_125_3477_n2377), .A2(
        DP_OP_423J2_125_3477_n2386), .Y(DP_OP_423J2_125_3477_n2353) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1578 ( .A1(DP_OP_422J2_124_3477_n2344), .A2(
        DP_OP_425J2_127_3477_n2387), .Y(DP_OP_423J2_125_3477_n2352) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1577 ( .A1(DP_OP_422J2_124_3477_n2343), .A2(
        DP_OP_424J2_126_3477_n2387), .Y(DP_OP_423J2_125_3477_n2351) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1576 ( .A1(DP_OP_422J2_124_3477_n2342), .A2(
        DP_OP_422J2_124_3477_n2389), .Y(DP_OP_423J2_125_3477_n2350) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1575 ( .A1(DP_OP_422J2_124_3477_n2341), .A2(
        DP_OP_425J2_127_3477_n2387), .Y(DP_OP_423J2_125_3477_n2349) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1574 ( .A1(DP_OP_422J2_124_3477_n2340), .A2(
        DP_OP_422J2_124_3477_n2389), .Y(DP_OP_423J2_125_3477_n2348) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1573 ( .A1(DP_OP_422J2_124_3477_n2339), .A2(
        DP_OP_422J2_124_3477_n2389), .Y(DP_OP_423J2_125_3477_n2347) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1572 ( .A1(DP_OP_422J2_124_3477_n2338), .A2(
        DP_OP_425J2_127_3477_n2387), .Y(DP_OP_423J2_125_3477_n2346) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1571 ( .A1(DP_OP_423J2_125_3477_n2377), 
        .A2(DP_OP_422J2_124_3477_n2389), .Y(DP_OP_423J2_125_3477_n2345) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1553 ( .A1(DP_OP_422J2_124_3477_n2427), 
        .A2(DP_OP_423J2_125_3477_n2344), .Y(DP_OP_423J2_125_3477_n2327) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1552 ( .A1(DP_OP_423J2_125_3477_n2334), 
        .A2(DP_OP_423J2_125_3477_n2344), .Y(DP_OP_423J2_125_3477_n2326) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1551 ( .A1(DP_OP_423J2_125_3477_n2333), .A2(
        DP_OP_423J2_125_3477_n2344), .Y(DP_OP_423J2_125_3477_n2325) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1544 ( .A1(DP_OP_423J2_125_3477_n2334), 
        .A2(DP_OP_423J2_125_3477_n2343), .Y(DP_OP_423J2_125_3477_n2318) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1543 ( .A1(DP_OP_423J2_125_3477_n2333), .A2(
        DP_OP_423J2_125_3477_n2343), .Y(DP_OP_423J2_125_3477_n2317) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1535 ( .A1(DP_OP_423J2_125_3477_n2333), .A2(
        n448), .Y(DP_OP_423J2_125_3477_n2309) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1534 ( .A1(DP_OP_422J2_124_3477_n2432), .A2(
        DP_OP_423J2_125_3477_n2341), .Y(DP_OP_423J2_125_3477_n2308) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1533 ( .A1(DP_OP_423J2_125_3477_n2339), .A2(
        DP_OP_423J2_125_3477_n2341), .Y(DP_OP_423J2_125_3477_n2307) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1532 ( .A1(DP_OP_422J2_124_3477_n2430), .A2(
        DP_OP_423J2_125_3477_n2341), .Y(DP_OP_423J2_125_3477_n2306) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1531 ( .A1(DP_OP_422J2_124_3477_n2429), .A2(
        DP_OP_423J2_125_3477_n2341), .Y(DP_OP_423J2_125_3477_n2305) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1530 ( .A1(DP_OP_422J2_124_3477_n2428), .A2(
        DP_OP_423J2_125_3477_n2341), .Y(DP_OP_423J2_125_3477_n2304) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1529 ( .A1(DP_OP_422J2_124_3477_n2427), .A2(
        DP_OP_423J2_125_3477_n2341), .Y(DP_OP_423J2_125_3477_n2303) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1528 ( .A1(DP_OP_423J2_125_3477_n2334), .A2(
        DP_OP_423J2_125_3477_n2341), .Y(DP_OP_423J2_125_3477_n2302) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1527 ( .A1(DP_OP_423J2_125_3477_n2333), 
        .A2(DP_OP_423J2_125_3477_n2341), .Y(DP_OP_423J2_125_3477_n2301) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1509 ( .A1(DP_OP_423J2_125_3477_n2291), 
        .A2(DP_OP_425J2_127_3477_n2305), .Y(DP_OP_423J2_125_3477_n2283) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1508 ( .A1(DP_OP_422J2_124_3477_n2470), 
        .A2(n446), .Y(DP_OP_423J2_125_3477_n2282) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1507 ( .A1(DP_OP_422J2_124_3477_n2469), .A2(
        n446), .Y(DP_OP_423J2_125_3477_n2281) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1500 ( .A1(DP_OP_422J2_124_3477_n2470), 
        .A2(DP_OP_423J2_125_3477_n2299), .Y(DP_OP_423J2_125_3477_n2274) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1499 ( .A1(DP_OP_422J2_124_3477_n2469), .A2(
        DP_OP_423J2_125_3477_n2299), .Y(DP_OP_423J2_125_3477_n2273) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1492 ( .A1(DP_OP_422J2_124_3477_n2470), 
        .A2(DP_OP_423J2_125_3477_n2298), .Y(DP_OP_423J2_125_3477_n2266) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1491 ( .A1(DP_OP_422J2_124_3477_n2469), .A2(
        DP_OP_423J2_125_3477_n2298), .Y(DP_OP_423J2_125_3477_n2265) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1490 ( .A1(DP_OP_422J2_124_3477_n2476), .A2(
        DP_OP_422J2_124_3477_n2301), .Y(DP_OP_423J2_125_3477_n2264) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1489 ( .A1(DP_OP_423J2_125_3477_n2295), .A2(
        DP_OP_422J2_124_3477_n2301), .Y(DP_OP_423J2_125_3477_n2263) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1488 ( .A1(DP_OP_423J2_125_3477_n2294), .A2(
        DP_OP_424J2_126_3477_n2302), .Y(DP_OP_423J2_125_3477_n2262) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1487 ( .A1(DP_OP_422J2_124_3477_n2473), .A2(
        DP_OP_422J2_124_3477_n2301), .Y(DP_OP_423J2_125_3477_n2261) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1486 ( .A1(DP_OP_422J2_124_3477_n2472), .A2(
        DP_OP_425J2_127_3477_n2302), .Y(DP_OP_423J2_125_3477_n2260) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1485 ( .A1(DP_OP_423J2_125_3477_n2291), .A2(
        DP_OP_424J2_126_3477_n2302), .Y(DP_OP_423J2_125_3477_n2259) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1484 ( .A1(DP_OP_422J2_124_3477_n2470), .A2(
        DP_OP_422J2_124_3477_n2301), .Y(DP_OP_423J2_125_3477_n2258) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1483 ( .A1(DP_OP_422J2_124_3477_n2469), 
        .A2(DP_OP_425J2_127_3477_n2302), .Y(DP_OP_423J2_125_3477_n2257) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1464 ( .A1(DP_OP_424J2_126_3477_n2339), 
        .A2(DP_OP_423J2_125_3477_n2256), .Y(DP_OP_423J2_125_3477_n2238) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1463 ( .A1(DP_OP_424J2_126_3477_n2338), .A2(
        DP_OP_423J2_125_3477_n2256), .Y(DP_OP_423J2_125_3477_n2237) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1456 ( .A1(DP_OP_422J2_124_3477_n2514), 
        .A2(DP_OP_424J2_126_3477_n2260), .Y(DP_OP_423J2_125_3477_n2230) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1455 ( .A1(DP_OP_424J2_126_3477_n2338), .A2(
        DP_OP_424J2_126_3477_n2260), .Y(DP_OP_423J2_125_3477_n2229) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1448 ( .A1(DP_OP_422J2_124_3477_n2514), 
        .A2(DP_OP_423J2_125_3477_n2254), .Y(DP_OP_423J2_125_3477_n2222) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1447 ( .A1(DP_OP_424J2_126_3477_n2338), .A2(
        DP_OP_423J2_125_3477_n2254), .Y(DP_OP_423J2_125_3477_n2221) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1446 ( .A1(DP_OP_422J2_124_3477_n2520), .A2(
        DP_OP_422J2_124_3477_n2257), .Y(DP_OP_423J2_125_3477_n2220) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1445 ( .A1(DP_OP_423J2_125_3477_n2251), .A2(
        n450), .Y(DP_OP_423J2_125_3477_n2219) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1444 ( .A1(DP_OP_425J2_127_3477_n2384), .A2(
        DP_OP_422J2_124_3477_n2257), .Y(DP_OP_423J2_125_3477_n2218) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1443 ( .A1(DP_OP_425J2_127_3477_n2383), .A2(
        DP_OP_422J2_124_3477_n2257), .Y(DP_OP_423J2_125_3477_n2217) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1442 ( .A1(DP_OP_425J2_127_3477_n2382), .A2(
        DP_OP_422J2_124_3477_n2257), .Y(DP_OP_423J2_125_3477_n2216) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1441 ( .A1(DP_OP_423J2_125_3477_n2247), .A2(
        n450), .Y(DP_OP_423J2_125_3477_n2215) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1440 ( .A1(DP_OP_424J2_126_3477_n2339), .A2(
        n450), .Y(DP_OP_423J2_125_3477_n2214) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1439 ( .A1(DP_OP_424J2_126_3477_n2338), 
        .A2(DP_OP_424J2_126_3477_n2258), .Y(DP_OP_423J2_125_3477_n2213) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1421 ( .A1(DP_OP_424J2_126_3477_n2296), 
        .A2(DP_OP_423J2_125_3477_n2212), .Y(DP_OP_423J2_125_3477_n2195) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1420 ( .A1(DP_OP_425J2_127_3477_n2424), 
        .A2(DP_OP_423J2_125_3477_n2212), .Y(DP_OP_423J2_125_3477_n2194) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1419 ( .A1(DP_OP_425J2_127_3477_n2423), .A2(
        DP_OP_423J2_125_3477_n2212), .Y(DP_OP_423J2_125_3477_n2193) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1412 ( .A1(DP_OP_425J2_127_3477_n2424), 
        .A2(DP_OP_423J2_125_3477_n2211), .Y(DP_OP_423J2_125_3477_n2186) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1411 ( .A1(DP_OP_425J2_127_3477_n2423), .A2(
        DP_OP_423J2_125_3477_n2211), .Y(DP_OP_423J2_125_3477_n2185) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1403 ( .A1(DP_OP_425J2_127_3477_n2423), .A2(
        DP_OP_425J2_127_3477_n2215), .Y(DP_OP_423J2_125_3477_n2177) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1402 ( .A1(DP_OP_425J2_127_3477_n2430), .A2(
        DP_OP_423J2_125_3477_n2209), .Y(DP_OP_423J2_125_3477_n2176) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1401 ( .A1(DP_OP_425J2_127_3477_n2429), .A2(
        DP_OP_423J2_125_3477_n2209), .Y(DP_OP_423J2_125_3477_n2175) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1400 ( .A1(DP_OP_422J2_124_3477_n2562), .A2(
        DP_OP_423J2_125_3477_n2209), .Y(DP_OP_423J2_125_3477_n2174) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1399 ( .A1(DP_OP_423J2_125_3477_n2205), .A2(
        DP_OP_423J2_125_3477_n2209), .Y(DP_OP_423J2_125_3477_n2173) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1398 ( .A1(DP_OP_423J2_125_3477_n2204), .A2(
        DP_OP_423J2_125_3477_n2209), .Y(DP_OP_423J2_125_3477_n2172) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1397 ( .A1(DP_OP_422J2_124_3477_n2559), .A2(
        DP_OP_423J2_125_3477_n2209), .Y(DP_OP_423J2_125_3477_n2171) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1396 ( .A1(DP_OP_425J2_127_3477_n2424), .A2(
        DP_OP_423J2_125_3477_n2209), .Y(DP_OP_423J2_125_3477_n2170) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1395 ( .A1(DP_OP_425J2_127_3477_n2423), 
        .A2(DP_OP_423J2_125_3477_n2209), .Y(DP_OP_423J2_125_3477_n2169) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1376 ( .A1(DP_OP_423J2_125_3477_n2158), 
        .A2(DP_OP_423J2_125_3477_n2168), .Y(DP_OP_423J2_125_3477_n2150) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1375 ( .A1(DP_OP_423J2_125_3477_n2157), .A2(
        DP_OP_423J2_125_3477_n2168), .Y(DP_OP_423J2_125_3477_n2149) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1368 ( .A1(DP_OP_423J2_125_3477_n2158), 
        .A2(DP_OP_423J2_125_3477_n2167), .Y(DP_OP_423J2_125_3477_n2142) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1367 ( .A1(DP_OP_423J2_125_3477_n2157), .A2(
        DP_OP_423J2_125_3477_n2167), .Y(DP_OP_423J2_125_3477_n2141) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1360 ( .A1(DP_OP_423J2_125_3477_n2158), 
        .A2(n452), .Y(DP_OP_423J2_125_3477_n2134) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1359 ( .A1(DP_OP_423J2_125_3477_n2157), .A2(
        DP_OP_422J2_124_3477_n2170), .Y(DP_OP_423J2_125_3477_n2133) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1358 ( .A1(DP_OP_423J2_125_3477_n2164), .A2(
        DP_OP_423J2_125_3477_n2165), .Y(DP_OP_423J2_125_3477_n2132) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1357 ( .A1(DP_OP_423J2_125_3477_n2163), .A2(
        DP_OP_423J2_125_3477_n2165), .Y(DP_OP_423J2_125_3477_n2131) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1356 ( .A1(DP_OP_425J2_127_3477_n2472), .A2(
        DP_OP_423J2_125_3477_n2165), .Y(DP_OP_423J2_125_3477_n2130) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1355 ( .A1(DP_OP_423J2_125_3477_n2161), .A2(
        DP_OP_423J2_125_3477_n2165), .Y(DP_OP_423J2_125_3477_n2129) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1354 ( .A1(DP_OP_423J2_125_3477_n2160), .A2(
        DP_OP_423J2_125_3477_n2165), .Y(DP_OP_423J2_125_3477_n2128) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1353 ( .A1(DP_OP_425J2_127_3477_n2469), .A2(
        DP_OP_423J2_125_3477_n2165), .Y(DP_OP_423J2_125_3477_n2127) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1352 ( .A1(DP_OP_423J2_125_3477_n2158), .A2(
        DP_OP_423J2_125_3477_n2165), .Y(DP_OP_423J2_125_3477_n2126) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1351 ( .A1(DP_OP_423J2_125_3477_n2157), 
        .A2(DP_OP_423J2_125_3477_n2165), .Y(DP_OP_423J2_125_3477_n2125) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1332 ( .A1(DP_OP_423J2_125_3477_n2114), 
        .A2(DP_OP_425J2_127_3477_n2129), .Y(DP_OP_423J2_125_3477_n2106) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1331 ( .A1(DP_OP_422J2_124_3477_n2645), .A2(
        DP_OP_424J2_126_3477_n2129), .Y(DP_OP_423J2_125_3477_n2105) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1324 ( .A1(DP_OP_423J2_125_3477_n2114), 
        .A2(DP_OP_422J2_124_3477_n2127), .Y(DP_OP_423J2_125_3477_n2098) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1323 ( .A1(DP_OP_422J2_124_3477_n2645), .A2(
        n440), .Y(DP_OP_423J2_125_3477_n2097) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1316 ( .A1(DP_OP_423J2_125_3477_n2114), 
        .A2(DP_OP_423J2_125_3477_n2122), .Y(DP_OP_423J2_125_3477_n2090) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1315 ( .A1(DP_OP_425J2_127_3477_n2511), .A2(
        DP_OP_423J2_125_3477_n2122), .Y(DP_OP_423J2_125_3477_n2089) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1314 ( .A1(DP_OP_425J2_127_3477_n2518), .A2(
        DP_OP_424J2_126_3477_n2126), .Y(DP_OP_423J2_125_3477_n2088) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1313 ( .A1(DP_OP_422J2_124_3477_n2651), .A2(
        DP_OP_424J2_126_3477_n2126), .Y(DP_OP_423J2_125_3477_n2087) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1312 ( .A1(DP_OP_422J2_124_3477_n2650), .A2(
        DP_OP_424J2_126_3477_n2126), .Y(DP_OP_423J2_125_3477_n2086) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1311 ( .A1(DP_OP_423J2_125_3477_n2117), .A2(
        DP_OP_424J2_126_3477_n2126), .Y(DP_OP_423J2_125_3477_n2085) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1310 ( .A1(DP_OP_423J2_125_3477_n2116), .A2(
        DP_OP_422J2_124_3477_n2125), .Y(DP_OP_423J2_125_3477_n2084) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1309 ( .A1(DP_OP_423J2_125_3477_n2115), .A2(
        DP_OP_424J2_126_3477_n2126), .Y(DP_OP_423J2_125_3477_n2083) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1308 ( .A1(DP_OP_423J2_125_3477_n2114), .A2(
        DP_OP_422J2_124_3477_n2125), .Y(DP_OP_423J2_125_3477_n2082) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1307 ( .A1(DP_OP_425J2_127_3477_n2511), 
        .A2(DP_OP_425J2_127_3477_n2126), .Y(DP_OP_423J2_125_3477_n2081) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1288 ( .A1(DP_OP_422J2_124_3477_n2690), 
        .A2(DP_OP_423J2_125_3477_n2080), .Y(DP_OP_423J2_125_3477_n2062) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1287 ( .A1(DP_OP_425J2_127_3477_n2555), .A2(
        DP_OP_423J2_125_3477_n2080), .Y(DP_OP_423J2_125_3477_n2061) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1280 ( .A1(DP_OP_422J2_124_3477_n2690), 
        .A2(DP_OP_422J2_124_3477_n2083), .Y(DP_OP_423J2_125_3477_n2054) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1279 ( .A1(DP_OP_425J2_127_3477_n2555), .A2(
        DP_OP_425J2_127_3477_n2084), .Y(DP_OP_423J2_125_3477_n2053) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1272 ( .A1(DP_OP_424J2_126_3477_n2163), 
        .A2(DP_OP_425J2_127_3477_n2083), .Y(DP_OP_423J2_125_3477_n2046) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1271 ( .A1(DP_OP_422J2_124_3477_n2689), .A2(
        n447), .Y(DP_OP_423J2_125_3477_n2045) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1270 ( .A1(DP_OP_423J2_125_3477_n2076), .A2(
        DP_OP_423J2_125_3477_n2077), .Y(DP_OP_423J2_125_3477_n2044) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1269 ( .A1(DP_OP_424J2_126_3477_n2168), .A2(
        DP_OP_423J2_125_3477_n2077), .Y(DP_OP_423J2_125_3477_n2043) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1268 ( .A1(DP_OP_423J2_125_3477_n2074), .A2(
        DP_OP_423J2_125_3477_n2077), .Y(DP_OP_423J2_125_3477_n2042) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1267 ( .A1(DP_OP_423J2_125_3477_n2073), .A2(
        DP_OP_423J2_125_3477_n2077), .Y(DP_OP_423J2_125_3477_n2041) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1266 ( .A1(DP_OP_422J2_124_3477_n2692), .A2(
        DP_OP_423J2_125_3477_n2077), .Y(DP_OP_423J2_125_3477_n2040) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1265 ( .A1(DP_OP_424J2_126_3477_n2164), .A2(
        DP_OP_423J2_125_3477_n2077), .Y(DP_OP_423J2_125_3477_n2039) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1264 ( .A1(DP_OP_422J2_124_3477_n2690), .A2(
        DP_OP_423J2_125_3477_n2077), .Y(DP_OP_423J2_125_3477_n2038) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1263 ( .A1(DP_OP_422J2_124_3477_n2689), 
        .A2(DP_OP_423J2_125_3477_n2077), .Y(DP_OP_423J2_125_3477_n2037) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1244 ( .A1(DP_OP_424J2_126_3477_n2119), 
        .A2(DP_OP_425J2_127_3477_n2041), .Y(DP_OP_423J2_125_3477_n2018) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1243 ( .A1(DP_OP_422J2_124_3477_n2731), .A2(
        DP_OP_422J2_124_3477_n2040), .Y(DP_OP_423J2_125_3477_n2017) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1237 ( .A1(DP_OP_424J2_126_3477_n2120), 
        .A2(DP_OP_425J2_127_3477_n2040), .Y(DP_OP_423J2_125_3477_n2011) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1236 ( .A1(DP_OP_424J2_126_3477_n2119), 
        .A2(DP_OP_424J2_126_3477_n2040), .Y(DP_OP_423J2_125_3477_n2010) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1235 ( .A1(DP_OP_424J2_126_3477_n2118), .A2(
        DP_OP_424J2_126_3477_n2040), .Y(DP_OP_423J2_125_3477_n2009) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1227 ( .A1(DP_OP_422J2_124_3477_n2731), .A2(
        DP_OP_423J2_125_3477_n2034), .Y(DP_OP_423J2_125_3477_n2001) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1226 ( .A1(DP_OP_423J2_125_3477_n2032), .A2(
        DP_OP_423J2_125_3477_n2033), .Y(DP_OP_423J2_125_3477_n2000) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1225 ( .A1(DP_OP_423J2_125_3477_n2031), .A2(
        DP_OP_423J2_125_3477_n2033), .Y(DP_OP_423J2_125_3477_n1999) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1224 ( .A1(DP_OP_423J2_125_3477_n2030), .A2(
        DP_OP_423J2_125_3477_n2033), .Y(DP_OP_423J2_125_3477_n1998) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1223 ( .A1(DP_OP_423J2_125_3477_n2029), .A2(
        DP_OP_423J2_125_3477_n2033), .Y(DP_OP_423J2_125_3477_n1997) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1222 ( .A1(DP_OP_423J2_125_3477_n2028), .A2(
        DP_OP_423J2_125_3477_n2033), .Y(DP_OP_423J2_125_3477_n1996) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1221 ( .A1(DP_OP_424J2_126_3477_n2120), .A2(
        DP_OP_423J2_125_3477_n2033), .Y(DP_OP_423J2_125_3477_n1995) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1220 ( .A1(DP_OP_422J2_124_3477_n2732), .A2(
        DP_OP_423J2_125_3477_n2033), .Y(DP_OP_423J2_125_3477_n1994) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1219 ( .A1(DP_OP_424J2_126_3477_n2118), 
        .A2(DP_OP_423J2_125_3477_n2033), .Y(DP_OP_423J2_125_3477_n1993) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1200 ( .A1(DP_OP_422J2_124_3477_n2776), 
        .A2(DP_OP_423J2_125_3477_n1992), .Y(DP_OP_423J2_125_3477_n1974) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1199 ( .A1(DP_OP_425J2_127_3477_n2643), .A2(
        DP_OP_423J2_125_3477_n1992), .Y(DP_OP_423J2_125_3477_n1973) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1192 ( .A1(DP_OP_422J2_124_3477_n2776), 
        .A2(DP_OP_423J2_125_3477_n1991), .Y(DP_OP_423J2_125_3477_n1966) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1191 ( .A1(DP_OP_425J2_127_3477_n2643), .A2(
        DP_OP_423J2_125_3477_n1991), .Y(DP_OP_423J2_125_3477_n1965) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1184 ( .A1(DP_OP_422J2_124_3477_n2776), 
        .A2(DP_OP_425J2_127_3477_n1995), .Y(DP_OP_423J2_125_3477_n1958) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1183 ( .A1(DP_OP_424J2_126_3477_n2074), .A2(
        DP_OP_425J2_127_3477_n1995), .Y(DP_OP_423J2_125_3477_n1957) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1182 ( .A1(DP_OP_422J2_124_3477_n2782), .A2(
        DP_OP_423J2_125_3477_n1989), .Y(DP_OP_423J2_125_3477_n1956) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1181 ( .A1(DP_OP_422J2_124_3477_n2781), .A2(
        DP_OP_423J2_125_3477_n1989), .Y(DP_OP_423J2_125_3477_n1955) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1180 ( .A1(DP_OP_423J2_125_3477_n1986), .A2(
        DP_OP_423J2_125_3477_n1989), .Y(DP_OP_423J2_125_3477_n1954) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1179 ( .A1(DP_OP_423J2_125_3477_n1985), .A2(
        DP_OP_423J2_125_3477_n1989), .Y(DP_OP_423J2_125_3477_n1953) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1178 ( .A1(DP_OP_424J2_126_3477_n2077), .A2(
        DP_OP_423J2_125_3477_n1989), .Y(DP_OP_423J2_125_3477_n1952) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1177 ( .A1(DP_OP_423J2_125_3477_n1983), .A2(
        DP_OP_423J2_125_3477_n1989), .Y(DP_OP_423J2_125_3477_n1951) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1176 ( .A1(DP_OP_425J2_127_3477_n2644), .A2(
        DP_OP_423J2_125_3477_n1989), .Y(DP_OP_423J2_125_3477_n1950) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1175 ( .A1(DP_OP_425J2_127_3477_n2643), 
        .A2(DP_OP_423J2_125_3477_n1989), .Y(DP_OP_423J2_125_3477_n1949) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1157 ( .A1(DP_OP_423J2_125_3477_n1939), 
        .A2(DP_OP_423J2_125_3477_n1948), .Y(DP_OP_423J2_125_3477_n1931) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1156 ( .A1(DP_OP_425J2_127_3477_n2688), 
        .A2(DP_OP_423J2_125_3477_n1948), .Y(DP_OP_423J2_125_3477_n1930) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1155 ( .A1(DP_OP_423J2_125_3477_n1937), .A2(
        DP_OP_423J2_125_3477_n1948), .Y(DP_OP_423J2_125_3477_n1929) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1148 ( .A1(DP_OP_425J2_127_3477_n2688), 
        .A2(DP_OP_423J2_125_3477_n1947), .Y(DP_OP_423J2_125_3477_n1922) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1147 ( .A1(DP_OP_423J2_125_3477_n1937), .A2(
        DP_OP_423J2_125_3477_n1947), .Y(DP_OP_423J2_125_3477_n1921) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1139 ( .A1(DP_OP_423J2_125_3477_n1937), .A2(
        n442), .Y(DP_OP_423J2_125_3477_n1913) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1138 ( .A1(DP_OP_425J2_127_3477_n2694), .A2(
        DP_OP_425J2_127_3477_n1950), .Y(DP_OP_423J2_125_3477_n1912) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1137 ( .A1(DP_OP_423J2_125_3477_n1943), .A2(
        DP_OP_425J2_127_3477_n1950), .Y(DP_OP_423J2_125_3477_n1911) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1136 ( .A1(DP_OP_425J2_127_3477_n2692), .A2(
        DP_OP_424J2_126_3477_n1950), .Y(DP_OP_423J2_125_3477_n1910) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1135 ( .A1(DP_OP_425J2_127_3477_n2691), .A2(
        DP_OP_424J2_126_3477_n1950), .Y(DP_OP_423J2_125_3477_n1909) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1134 ( .A1(DP_OP_425J2_127_3477_n2690), .A2(
        DP_OP_425J2_127_3477_n1950), .Y(DP_OP_423J2_125_3477_n1908) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1133 ( .A1(DP_OP_423J2_125_3477_n1939), .A2(
        DP_OP_425J2_127_3477_n1950), .Y(DP_OP_423J2_125_3477_n1907) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1132 ( .A1(DP_OP_425J2_127_3477_n2688), .A2(
        DP_OP_425J2_127_3477_n1950), .Y(DP_OP_423J2_125_3477_n1906) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1131 ( .A1(DP_OP_423J2_125_3477_n1937), 
        .A2(DP_OP_422J2_124_3477_n1950), .Y(DP_OP_423J2_125_3477_n1905) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1112 ( .A1(DP_OP_425J2_127_3477_n2732), 
        .A2(DP_OP_423J2_125_3477_n1904), .Y(DP_OP_423J2_125_3477_n1886) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1111 ( .A1(DP_OP_423J2_125_3477_n1893), .A2(
        DP_OP_423J2_125_3477_n1904), .Y(DP_OP_423J2_125_3477_n1885) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1104 ( .A1(DP_OP_425J2_127_3477_n2732), 
        .A2(n449), .Y(DP_OP_423J2_125_3477_n1878) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1103 ( .A1(DP_OP_423J2_125_3477_n1893), .A2(
        n449), .Y(DP_OP_423J2_125_3477_n1877) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1095 ( .A1(DP_OP_423J2_125_3477_n1893), .A2(
        DP_OP_424J2_126_3477_n1907), .Y(DP_OP_423J2_125_3477_n1869) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1094 ( .A1(DP_OP_425J2_127_3477_n2738), .A2(
        DP_OP_423J2_125_3477_n1901), .Y(DP_OP_423J2_125_3477_n1868) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1093 ( .A1(DP_OP_423J2_125_3477_n1899), .A2(
        DP_OP_423J2_125_3477_n1901), .Y(DP_OP_423J2_125_3477_n1867) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1092 ( .A1(DP_OP_423J2_125_3477_n1898), .A2(
        DP_OP_423J2_125_3477_n1901), .Y(DP_OP_423J2_125_3477_n1866) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1091 ( .A1(DP_OP_423J2_125_3477_n1897), .A2(
        DP_OP_423J2_125_3477_n1901), .Y(DP_OP_423J2_125_3477_n1865) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1090 ( .A1(DP_OP_423J2_125_3477_n1896), .A2(
        DP_OP_423J2_125_3477_n1901), .Y(DP_OP_423J2_125_3477_n1864) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1089 ( .A1(DP_OP_424J2_126_3477_n1988), .A2(
        DP_OP_423J2_125_3477_n1901), .Y(DP_OP_423J2_125_3477_n1863) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1088 ( .A1(DP_OP_425J2_127_3477_n2732), .A2(
        DP_OP_423J2_125_3477_n1901), .Y(DP_OP_423J2_125_3477_n1862) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1087 ( .A1(DP_OP_423J2_125_3477_n1893), 
        .A2(DP_OP_423J2_125_3477_n1901), .Y(DP_OP_423J2_125_3477_n1861) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1068 ( .A1(DP_OP_423J2_125_3477_n1850), 
        .A2(DP_OP_423J2_125_3477_n1860), .Y(DP_OP_423J2_125_3477_n1842) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1067 ( .A1(DP_OP_423J2_125_3477_n1849), .A2(
        DP_OP_423J2_125_3477_n1860), .Y(DP_OP_423J2_125_3477_n1841) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1059 ( .A1(DP_OP_423J2_125_3477_n1849), .A2(
        DP_OP_423J2_125_3477_n1859), .Y(DP_OP_423J2_125_3477_n1833) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1052 ( .A1(DP_OP_423J2_125_3477_n1850), 
        .A2(DP_OP_423J2_125_3477_n1858), .Y(DP_OP_423J2_125_3477_n1826) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1051 ( .A1(DP_OP_423J2_125_3477_n1849), .A2(
        DP_OP_423J2_125_3477_n1858), .Y(DP_OP_423J2_125_3477_n1825) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1050 ( .A1(DP_OP_423J2_125_3477_n1856), .A2(
        DP_OP_425J2_127_3477_n1862), .Y(DP_OP_423J2_125_3477_n1824) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1049 ( .A1(DP_OP_424J2_126_3477_n1948), .A2(
        DP_OP_424J2_126_3477_n1862), .Y(DP_OP_423J2_125_3477_n1823) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1048 ( .A1(DP_OP_422J2_124_3477_n2912), .A2(
        DP_OP_424J2_126_3477_n1862), .Y(DP_OP_423J2_125_3477_n1822) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1047 ( .A1(DP_OP_423J2_125_3477_n1853), .A2(
        DP_OP_425J2_127_3477_n1862), .Y(DP_OP_423J2_125_3477_n1821) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1046 ( .A1(DP_OP_423J2_125_3477_n1852), .A2(
        DP_OP_424J2_126_3477_n1862), .Y(DP_OP_423J2_125_3477_n1820) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1045 ( .A1(DP_OP_425J2_127_3477_n2777), .A2(
        DP_OP_425J2_127_3477_n1862), .Y(DP_OP_423J2_125_3477_n1819) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1044 ( .A1(DP_OP_423J2_125_3477_n1850), .A2(
        DP_OP_424J2_126_3477_n1862), .Y(DP_OP_423J2_125_3477_n1818) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1043 ( .A1(DP_OP_423J2_125_3477_n1849), 
        .A2(DP_OP_425J2_127_3477_n1862), .Y(DP_OP_423J2_125_3477_n1817) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U995 ( .A1(n296), .A2(n339), .Y(
        DP_OP_423J2_125_3477_n184) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U991 ( .A1(n313), .A2(n338), .Y(
        DP_OP_423J2_125_3477_n172) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U990 ( .A1(n304), .A2(
        DP_OP_423J2_125_3477_n2), .Y(DP_OP_423J2_125_3477_n170) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U989 ( .A1(n308), .A2(
        DP_OP_424J2_126_3477_n2), .Y(DP_OP_423J2_125_3477_n168) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U988 ( .A1(n311), .A2(n337), .Y(
        DP_OP_423J2_125_3477_n166) );
  HADDX1_HVT DP_OP_423J2_125_3477_U977 ( .A0(DP_OP_423J2_125_3477_n1783), .B0(
        DP_OP_423J2_125_3477_n2725), .C1(DP_OP_423J2_125_3477_n1766), .SO(
        DP_OP_423J2_125_3477_n1767) );
  FADDX1_HVT DP_OP_423J2_125_3477_U976 ( .A(DP_OP_423J2_125_3477_n1848), .B(
        DP_OP_423J2_125_3477_n2684), .CI(DP_OP_423J2_125_3477_n2508), .CO(
        DP_OP_423J2_125_3477_n1764), .S(DP_OP_423J2_125_3477_n1765) );
  FADDX1_HVT DP_OP_423J2_125_3477_U975 ( .A(DP_OP_423J2_125_3477_n2552), .B(
        DP_OP_423J2_125_3477_n2024), .CI(DP_OP_423J2_125_3477_n1892), .CO(
        DP_OP_423J2_125_3477_n1762), .S(DP_OP_423J2_125_3477_n1763) );
  FADDX1_HVT DP_OP_423J2_125_3477_U974 ( .A(DP_OP_423J2_125_3477_n2464), .B(
        DP_OP_423J2_125_3477_n1980), .CI(DP_OP_423J2_125_3477_n2769), .CO(
        DP_OP_423J2_125_3477_n1760), .S(DP_OP_423J2_125_3477_n1761) );
  FADDX1_HVT DP_OP_423J2_125_3477_U973 ( .A(DP_OP_423J2_125_3477_n2420), .B(
        DP_OP_423J2_125_3477_n2200), .CI(DP_OP_423J2_125_3477_n2857), .CO(
        DP_OP_423J2_125_3477_n1758), .S(DP_OP_423J2_125_3477_n1759) );
  FADDX1_HVT DP_OP_423J2_125_3477_U972 ( .A(DP_OP_423J2_125_3477_n2112), .B(
        DP_OP_423J2_125_3477_n2332), .CI(DP_OP_423J2_125_3477_n2640), .CO(
        DP_OP_423J2_125_3477_n1756), .S(DP_OP_423J2_125_3477_n1757) );
  FADDX1_HVT DP_OP_423J2_125_3477_U971 ( .A(DP_OP_423J2_125_3477_n2596), .B(
        DP_OP_423J2_125_3477_n2068), .CI(DP_OP_423J2_125_3477_n2288), .CO(
        DP_OP_423J2_125_3477_n1754), .S(DP_OP_423J2_125_3477_n1755) );
  FADDX1_HVT DP_OP_423J2_125_3477_U970 ( .A(DP_OP_423J2_125_3477_n2244), .B(
        DP_OP_423J2_125_3477_n1936), .CI(DP_OP_423J2_125_3477_n2376), .CO(
        DP_OP_423J2_125_3477_n1752), .S(DP_OP_423J2_125_3477_n1753) );
  FADDX1_HVT DP_OP_423J2_125_3477_U969 ( .A(DP_OP_423J2_125_3477_n2156), .B(
        DP_OP_423J2_125_3477_n2901), .CI(DP_OP_423J2_125_3477_n2813), .CO(
        DP_OP_423J2_125_3477_n1750), .S(DP_OP_423J2_125_3477_n1751) );
  FADDX1_HVT DP_OP_423J2_125_3477_U968 ( .A(DP_OP_423J2_125_3477_n1767), .B(
        DP_OP_423J2_125_3477_n1759), .CI(DP_OP_423J2_125_3477_n1761), .CO(
        DP_OP_423J2_125_3477_n1748), .S(DP_OP_423J2_125_3477_n1749) );
  FADDX1_HVT DP_OP_423J2_125_3477_U967 ( .A(DP_OP_423J2_125_3477_n1765), .B(
        DP_OP_423J2_125_3477_n1757), .CI(DP_OP_423J2_125_3477_n1755), .CO(
        DP_OP_423J2_125_3477_n1746), .S(DP_OP_423J2_125_3477_n1747) );
  FADDX1_HVT DP_OP_423J2_125_3477_U966 ( .A(DP_OP_423J2_125_3477_n1763), .B(
        DP_OP_423J2_125_3477_n1753), .CI(DP_OP_423J2_125_3477_n1751), .CO(
        DP_OP_423J2_125_3477_n1744), .S(DP_OP_423J2_125_3477_n1745) );
  HADDX1_HVT DP_OP_423J2_125_3477_U965 ( .A0(DP_OP_423J2_125_3477_n1782), .B0(
        DP_OP_423J2_125_3477_n2412), .C1(DP_OP_423J2_125_3477_n1742), .SO(
        DP_OP_423J2_125_3477_n1743) );
  FADDX1_HVT DP_OP_423J2_125_3477_U964 ( .A(DP_OP_423J2_125_3477_n2551), .B(
        DP_OP_423J2_125_3477_n2724), .CI(DP_OP_423J2_125_3477_n2768), .CO(
        DP_OP_423J2_125_3477_n1740), .S(DP_OP_423J2_125_3477_n1741) );
  FADDX1_HVT DP_OP_423J2_125_3477_U963 ( .A(DP_OP_423J2_125_3477_n2111), .B(
        DP_OP_423J2_125_3477_n2148), .CI(DP_OP_423J2_125_3477_n1891), .CO(
        DP_OP_423J2_125_3477_n1738), .S(DP_OP_423J2_125_3477_n1739) );
  FADDX1_HVT DP_OP_423J2_125_3477_U962 ( .A(DP_OP_423J2_125_3477_n2199), .B(
        DP_OP_423J2_125_3477_n2023), .CI(DP_OP_423J2_125_3477_n2507), .CO(
        DP_OP_423J2_125_3477_n1736), .S(DP_OP_423J2_125_3477_n1737) );
  FADDX1_HVT DP_OP_423J2_125_3477_U961 ( .A(DP_OP_423J2_125_3477_n2331), .B(
        DP_OP_423J2_125_3477_n2060), .CI(DP_OP_423J2_125_3477_n2856), .CO(
        DP_OP_423J2_125_3477_n1734), .S(DP_OP_423J2_125_3477_n1735) );
  FADDX1_HVT DP_OP_423J2_125_3477_U960 ( .A(DP_OP_423J2_125_3477_n2463), .B(
        DP_OP_423J2_125_3477_n2500), .CI(DP_OP_423J2_125_3477_n1979), .CO(
        DP_OP_423J2_125_3477_n1732), .S(DP_OP_423J2_125_3477_n1733) );
  FADDX1_HVT DP_OP_423J2_125_3477_U959 ( .A(DP_OP_423J2_125_3477_n2419), .B(
        DP_OP_423J2_125_3477_n2588), .CI(DP_OP_423J2_125_3477_n2632), .CO(
        DP_OP_423J2_125_3477_n1730), .S(DP_OP_423J2_125_3477_n1731) );
  FADDX1_HVT DP_OP_423J2_125_3477_U958 ( .A(DP_OP_423J2_125_3477_n2595), .B(
        DP_OP_423J2_125_3477_n2324), .CI(DP_OP_423J2_125_3477_n2683), .CO(
        DP_OP_423J2_125_3477_n1728), .S(DP_OP_423J2_125_3477_n1729) );
  FADDX1_HVT DP_OP_423J2_125_3477_U957 ( .A(DP_OP_423J2_125_3477_n2639), .B(
        DP_OP_423J2_125_3477_n1847), .CI(DP_OP_423J2_125_3477_n1840), .CO(
        DP_OP_423J2_125_3477_n1726), .S(DP_OP_423J2_125_3477_n1727) );
  FADDX1_HVT DP_OP_423J2_125_3477_U956 ( .A(DP_OP_423J2_125_3477_n2287), .B(
        DP_OP_423J2_125_3477_n2243), .CI(DP_OP_423J2_125_3477_n2893), .CO(
        DP_OP_423J2_125_3477_n1724), .S(DP_OP_423J2_125_3477_n1725) );
  FADDX1_HVT DP_OP_423J2_125_3477_U955 ( .A(DP_OP_423J2_125_3477_n2067), .B(
        DP_OP_423J2_125_3477_n1884), .CI(DP_OP_423J2_125_3477_n2280), .CO(
        DP_OP_423J2_125_3477_n1722), .S(DP_OP_423J2_125_3477_n1723) );
  FADDX1_HVT DP_OP_423J2_125_3477_U954 ( .A(DP_OP_423J2_125_3477_n2676), .B(
        DP_OP_423J2_125_3477_n2456), .CI(DP_OP_423J2_125_3477_n2761), .CO(
        DP_OP_423J2_125_3477_n1720), .S(DP_OP_423J2_125_3477_n1721) );
  FADDX1_HVT DP_OP_423J2_125_3477_U953 ( .A(DP_OP_423J2_125_3477_n2104), .B(
        DP_OP_423J2_125_3477_n2544), .CI(DP_OP_423J2_125_3477_n2900), .CO(
        DP_OP_423J2_125_3477_n1718), .S(DP_OP_423J2_125_3477_n1719) );
  FADDX1_HVT DP_OP_423J2_125_3477_U952 ( .A(DP_OP_423J2_125_3477_n1935), .B(
        DP_OP_423J2_125_3477_n2375), .CI(DP_OP_423J2_125_3477_n2812), .CO(
        DP_OP_423J2_125_3477_n1716), .S(DP_OP_423J2_125_3477_n1717) );
  FADDX1_HVT DP_OP_423J2_125_3477_U951 ( .A(DP_OP_423J2_125_3477_n2849), .B(
        DP_OP_423J2_125_3477_n2717), .CI(DP_OP_423J2_125_3477_n1972), .CO(
        DP_OP_423J2_125_3477_n1714), .S(DP_OP_423J2_125_3477_n1715) );
  FADDX1_HVT DP_OP_423J2_125_3477_U950 ( .A(DP_OP_423J2_125_3477_n2155), .B(
        DP_OP_423J2_125_3477_n2236), .CI(DP_OP_423J2_125_3477_n2192), .CO(
        DP_OP_423J2_125_3477_n1712), .S(DP_OP_423J2_125_3477_n1713) );
  FADDX1_HVT DP_OP_423J2_125_3477_U949 ( .A(DP_OP_423J2_125_3477_n2016), .B(
        DP_OP_423J2_125_3477_n2805), .CI(DP_OP_423J2_125_3477_n2368), .CO(
        DP_OP_423J2_125_3477_n1710), .S(DP_OP_423J2_125_3477_n1711) );
  FADDX1_HVT DP_OP_423J2_125_3477_U948 ( .A(DP_OP_423J2_125_3477_n1928), .B(
        DP_OP_423J2_125_3477_n1766), .CI(DP_OP_423J2_125_3477_n1743), .CO(
        DP_OP_423J2_125_3477_n1708), .S(DP_OP_423J2_125_3477_n1709) );
  FADDX1_HVT DP_OP_423J2_125_3477_U947 ( .A(DP_OP_423J2_125_3477_n1764), .B(
        DP_OP_423J2_125_3477_n1756), .CI(DP_OP_423J2_125_3477_n1754), .CO(
        DP_OP_423J2_125_3477_n1706), .S(DP_OP_423J2_125_3477_n1707) );
  FADDX1_HVT DP_OP_423J2_125_3477_U946 ( .A(DP_OP_423J2_125_3477_n1760), .B(
        DP_OP_423J2_125_3477_n1762), .CI(DP_OP_423J2_125_3477_n1758), .CO(
        DP_OP_423J2_125_3477_n1704), .S(DP_OP_423J2_125_3477_n1705) );
  FADDX1_HVT DP_OP_423J2_125_3477_U945 ( .A(DP_OP_423J2_125_3477_n1752), .B(
        DP_OP_423J2_125_3477_n1750), .CI(DP_OP_423J2_125_3477_n1733), .CO(
        DP_OP_423J2_125_3477_n1702), .S(DP_OP_423J2_125_3477_n1703) );
  FADDX1_HVT DP_OP_423J2_125_3477_U944 ( .A(DP_OP_423J2_125_3477_n1731), .B(
        DP_OP_423J2_125_3477_n1737), .CI(DP_OP_423J2_125_3477_n1735), .CO(
        DP_OP_423J2_125_3477_n1700), .S(DP_OP_423J2_125_3477_n1701) );
  FADDX1_HVT DP_OP_423J2_125_3477_U943 ( .A(DP_OP_423J2_125_3477_n1729), .B(
        DP_OP_423J2_125_3477_n1739), .CI(DP_OP_423J2_125_3477_n1741), .CO(
        DP_OP_423J2_125_3477_n1698), .S(DP_OP_423J2_125_3477_n1699) );
  FADDX1_HVT DP_OP_423J2_125_3477_U942 ( .A(DP_OP_423J2_125_3477_n1727), .B(
        DP_OP_423J2_125_3477_n1723), .CI(DP_OP_423J2_125_3477_n1725), .CO(
        DP_OP_423J2_125_3477_n1696), .S(DP_OP_423J2_125_3477_n1697) );
  FADDX1_HVT DP_OP_423J2_125_3477_U941 ( .A(DP_OP_423J2_125_3477_n1721), .B(
        DP_OP_423J2_125_3477_n1719), .CI(DP_OP_423J2_125_3477_n1711), .CO(
        DP_OP_423J2_125_3477_n1694), .S(DP_OP_423J2_125_3477_n1695) );
  FADDX1_HVT DP_OP_423J2_125_3477_U940 ( .A(DP_OP_423J2_125_3477_n1717), .B(
        DP_OP_423J2_125_3477_n1715), .CI(DP_OP_423J2_125_3477_n1713), .CO(
        DP_OP_423J2_125_3477_n1692), .S(DP_OP_423J2_125_3477_n1693) );
  FADDX1_HVT DP_OP_423J2_125_3477_U939 ( .A(DP_OP_423J2_125_3477_n1709), .B(
        DP_OP_423J2_125_3477_n1748), .CI(DP_OP_423J2_125_3477_n1746), .CO(
        DP_OP_423J2_125_3477_n1690), .S(DP_OP_423J2_125_3477_n1691) );
  FADDX1_HVT DP_OP_423J2_125_3477_U938 ( .A(DP_OP_423J2_125_3477_n1707), .B(
        DP_OP_423J2_125_3477_n1705), .CI(DP_OP_423J2_125_3477_n1744), .CO(
        DP_OP_423J2_125_3477_n1688), .S(DP_OP_423J2_125_3477_n1689) );
  FADDX1_HVT DP_OP_423J2_125_3477_U937 ( .A(DP_OP_423J2_125_3477_n1703), .B(
        DP_OP_423J2_125_3477_n1701), .CI(DP_OP_423J2_125_3477_n1699), .CO(
        DP_OP_423J2_125_3477_n1686), .S(DP_OP_423J2_125_3477_n1687) );
  FADDX1_HVT DP_OP_423J2_125_3477_U936 ( .A(DP_OP_423J2_125_3477_n1697), .B(
        DP_OP_423J2_125_3477_n1695), .CI(DP_OP_423J2_125_3477_n1693), .CO(
        DP_OP_423J2_125_3477_n1684), .S(DP_OP_423J2_125_3477_n1685) );
  FADDX1_HVT DP_OP_423J2_125_3477_U935 ( .A(DP_OP_423J2_125_3477_n1691), .B(
        DP_OP_423J2_125_3477_n1689), .CI(DP_OP_423J2_125_3477_n1687), .CO(
        DP_OP_423J2_125_3477_n1682), .S(DP_OP_423J2_125_3477_n1683) );
  HADDX1_HVT DP_OP_423J2_125_3477_U934 ( .A0(DP_OP_423J2_125_3477_n1781), .B0(
        DP_OP_423J2_125_3477_n2147), .C1(DP_OP_423J2_125_3477_n1680), .SO(
        DP_OP_423J2_125_3477_n1681) );
  FADDX1_HVT DP_OP_423J2_125_3477_U933 ( .A(DP_OP_423J2_125_3477_n2550), .B(
        DP_OP_423J2_125_3477_n2723), .CI(DP_OP_423J2_125_3477_n2096), .CO(
        DP_OP_423J2_125_3477_n1678), .S(DP_OP_423J2_125_3477_n1679) );
  FADDX1_HVT DP_OP_423J2_125_3477_U932 ( .A(DP_OP_423J2_125_3477_n2462), .B(
        DP_OP_423J2_125_3477_n2411), .CI(DP_OP_423J2_125_3477_n2506), .CO(
        DP_OP_423J2_125_3477_n1676), .S(DP_OP_423J2_125_3477_n1677) );
  FADDX1_HVT DP_OP_423J2_125_3477_U931 ( .A(DP_OP_423J2_125_3477_n2841), .B(
        DP_OP_423J2_125_3477_n2536), .CI(DP_OP_423J2_125_3477_n2855), .CO(
        DP_OP_423J2_125_3477_n1674), .S(DP_OP_423J2_125_3477_n1675) );
  FADDX1_HVT DP_OP_423J2_125_3477_U930 ( .A(DP_OP_423J2_125_3477_n2638), .B(
        DP_OP_423J2_125_3477_n1964), .CI(DP_OP_423J2_125_3477_n2767), .CO(
        DP_OP_423J2_125_3477_n1672), .S(DP_OP_423J2_125_3477_n1673) );
  FADDX1_HVT DP_OP_423J2_125_3477_U929 ( .A(DP_OP_423J2_125_3477_n2594), .B(
        DP_OP_423J2_125_3477_n2499), .CI(DP_OP_423J2_125_3477_n2448), .CO(
        DP_OP_423J2_125_3477_n1670), .S(DP_OP_423J2_125_3477_n1671) );
  FADDX1_HVT DP_OP_423J2_125_3477_U928 ( .A(DP_OP_423J2_125_3477_n2110), .B(
        DP_OP_423J2_125_3477_n2587), .CI(DP_OP_423J2_125_3477_n2228), .CO(
        DP_OP_423J2_125_3477_n1668), .S(DP_OP_423J2_125_3477_n1669) );
  FADDX1_HVT DP_OP_423J2_125_3477_U927 ( .A(DP_OP_423J2_125_3477_n2418), .B(
        DP_OP_423J2_125_3477_n2682), .CI(DP_OP_423J2_125_3477_n1890), .CO(
        DP_OP_423J2_125_3477_n1666), .S(DP_OP_423J2_125_3477_n1667) );
  FADDX1_HVT DP_OP_423J2_125_3477_U926 ( .A(DP_OP_423J2_125_3477_n2885), .B(
        DP_OP_423J2_125_3477_n2059), .CI(DP_OP_423J2_125_3477_n1978), .CO(
        DP_OP_423J2_125_3477_n1664), .S(DP_OP_423J2_125_3477_n1665) );
  FADDX1_HVT DP_OP_423J2_125_3477_U925 ( .A(DP_OP_423J2_125_3477_n2330), .B(
        DP_OP_423J2_125_3477_n2753), .CI(DP_OP_423J2_125_3477_n2631), .CO(
        DP_OP_423J2_125_3477_n1662), .S(DP_OP_423J2_125_3477_n1663) );
  FADDX1_HVT DP_OP_423J2_125_3477_U924 ( .A(DP_OP_423J2_125_3477_n2198), .B(
        DP_OP_423J2_125_3477_n2323), .CI(DP_OP_423J2_125_3477_n2022), .CO(
        DP_OP_423J2_125_3477_n1660), .S(DP_OP_423J2_125_3477_n1661) );
  FADDX1_HVT DP_OP_423J2_125_3477_U923 ( .A(DP_OP_423J2_125_3477_n1846), .B(
        DP_OP_423J2_125_3477_n1839), .CI(DP_OP_423J2_125_3477_n2066), .CO(
        DP_OP_423J2_125_3477_n1658), .S(DP_OP_423J2_125_3477_n1659) );
  FADDX1_HVT DP_OP_423J2_125_3477_U922 ( .A(DP_OP_423J2_125_3477_n2140), .B(
        DP_OP_423J2_125_3477_n2360), .CI(DP_OP_423J2_125_3477_n2892), .CO(
        DP_OP_423J2_125_3477_n1656), .S(DP_OP_423J2_125_3477_n1657) );
  FADDX1_HVT DP_OP_423J2_125_3477_U921 ( .A(DP_OP_423J2_125_3477_n2286), .B(
        DP_OP_423J2_125_3477_n2242), .CI(DP_OP_423J2_125_3477_n2804), .CO(
        DP_OP_423J2_125_3477_n1654), .S(DP_OP_423J2_125_3477_n1655) );
  FADDX1_HVT DP_OP_423J2_125_3477_U920 ( .A(DP_OP_423J2_125_3477_n2272), .B(
        DP_OP_423J2_125_3477_n2103), .CI(DP_OP_423J2_125_3477_n2279), .CO(
        DP_OP_423J2_125_3477_n1652), .S(DP_OP_423J2_125_3477_n1653) );
  FADDX1_HVT DP_OP_423J2_125_3477_U919 ( .A(DP_OP_423J2_125_3477_n2580), .B(
        DP_OP_423J2_125_3477_n2455), .CI(DP_OP_423J2_125_3477_n2716), .CO(
        DP_OP_423J2_125_3477_n1650), .S(DP_OP_423J2_125_3477_n1651) );
  FADDX1_HVT DP_OP_423J2_125_3477_U918 ( .A(DP_OP_423J2_125_3477_n2675), .B(
        DP_OP_423J2_125_3477_n2492), .CI(DP_OP_423J2_125_3477_n2760), .CO(
        DP_OP_423J2_125_3477_n1648), .S(DP_OP_423J2_125_3477_n1649) );
  FADDX1_HVT DP_OP_423J2_125_3477_U917 ( .A(DP_OP_423J2_125_3477_n1883), .B(
        DP_OP_423J2_125_3477_n2668), .CI(DP_OP_423J2_125_3477_n2899), .CO(
        DP_OP_423J2_125_3477_n1646), .S(DP_OP_423J2_125_3477_n1647) );
  FADDX1_HVT DP_OP_423J2_125_3477_U916 ( .A(DP_OP_423J2_125_3477_n2709), .B(
        DP_OP_423J2_125_3477_n2374), .CI(DP_OP_423J2_125_3477_n2811), .CO(
        DP_OP_423J2_125_3477_n1644), .S(DP_OP_423J2_125_3477_n1645) );
  FADDX1_HVT DP_OP_423J2_125_3477_U915 ( .A(DP_OP_423J2_125_3477_n2543), .B(
        DP_OP_423J2_125_3477_n2367), .CI(DP_OP_423J2_125_3477_n1832), .CO(
        DP_OP_423J2_125_3477_n1642), .S(DP_OP_423J2_125_3477_n1643) );
  FADDX1_HVT DP_OP_423J2_125_3477_U914 ( .A(DP_OP_423J2_125_3477_n2052), .B(
        DP_OP_423J2_125_3477_n2235), .CI(DP_OP_423J2_125_3477_n2184), .CO(
        DP_OP_423J2_125_3477_n1640), .S(DP_OP_423J2_125_3477_n1641) );
  FADDX1_HVT DP_OP_423J2_125_3477_U913 ( .A(DP_OP_423J2_125_3477_n2316), .B(
        DP_OP_423J2_125_3477_n2008), .CI(DP_OP_423J2_125_3477_n1920), .CO(
        DP_OP_423J2_125_3477_n1638), .S(DP_OP_423J2_125_3477_n1639) );
  FADDX1_HVT DP_OP_423J2_125_3477_U912 ( .A(DP_OP_423J2_125_3477_n1934), .B(
        DP_OP_423J2_125_3477_n2191), .CI(DP_OP_423J2_125_3477_n2624), .CO(
        DP_OP_423J2_125_3477_n1636), .S(DP_OP_423J2_125_3477_n1637) );
  FADDX1_HVT DP_OP_423J2_125_3477_U911 ( .A(DP_OP_423J2_125_3477_n2848), .B(
        DP_OP_423J2_125_3477_n1927), .CI(DP_OP_423J2_125_3477_n1971), .CO(
        DP_OP_423J2_125_3477_n1634), .S(DP_OP_423J2_125_3477_n1635) );
  FADDX1_HVT DP_OP_423J2_125_3477_U910 ( .A(DP_OP_423J2_125_3477_n2015), .B(
        DP_OP_423J2_125_3477_n1876), .CI(DP_OP_423J2_125_3477_n2797), .CO(
        DP_OP_423J2_125_3477_n1632), .S(DP_OP_423J2_125_3477_n1633) );
  FADDX1_HVT DP_OP_423J2_125_3477_U909 ( .A(DP_OP_423J2_125_3477_n2404), .B(
        DP_OP_423J2_125_3477_n2154), .CI(DP_OP_423J2_125_3477_n1742), .CO(
        DP_OP_423J2_125_3477_n1630), .S(DP_OP_423J2_125_3477_n1631) );
  FADDX1_HVT DP_OP_423J2_125_3477_U908 ( .A(DP_OP_423J2_125_3477_n1681), .B(
        DP_OP_423J2_125_3477_n1740), .CI(DP_OP_423J2_125_3477_n1726), .CO(
        DP_OP_423J2_125_3477_n1628), .S(DP_OP_423J2_125_3477_n1629) );
  FADDX1_HVT DP_OP_423J2_125_3477_U907 ( .A(DP_OP_423J2_125_3477_n1738), .B(
        DP_OP_423J2_125_3477_n1728), .CI(DP_OP_423J2_125_3477_n1736), .CO(
        DP_OP_423J2_125_3477_n1626), .S(DP_OP_423J2_125_3477_n1627) );
  FADDX1_HVT DP_OP_423J2_125_3477_U906 ( .A(DP_OP_423J2_125_3477_n1734), .B(
        DP_OP_423J2_125_3477_n1730), .CI(DP_OP_423J2_125_3477_n1732), .CO(
        DP_OP_423J2_125_3477_n1624), .S(DP_OP_423J2_125_3477_n1625) );
  FADDX1_HVT DP_OP_423J2_125_3477_U905 ( .A(DP_OP_423J2_125_3477_n1722), .B(
        DP_OP_423J2_125_3477_n1718), .CI(DP_OP_423J2_125_3477_n1710), .CO(
        DP_OP_423J2_125_3477_n1622), .S(DP_OP_423J2_125_3477_n1623) );
  FADDX1_HVT DP_OP_423J2_125_3477_U904 ( .A(DP_OP_423J2_125_3477_n1724), .B(
        DP_OP_423J2_125_3477_n1720), .CI(DP_OP_423J2_125_3477_n1712), .CO(
        DP_OP_423J2_125_3477_n1620), .S(DP_OP_423J2_125_3477_n1621) );
  FADDX1_HVT DP_OP_423J2_125_3477_U903 ( .A(DP_OP_423J2_125_3477_n1716), .B(
        DP_OP_423J2_125_3477_n1714), .CI(DP_OP_423J2_125_3477_n1659), .CO(
        DP_OP_423J2_125_3477_n1618), .S(DP_OP_423J2_125_3477_n1619) );
  FADDX1_HVT DP_OP_423J2_125_3477_U902 ( .A(DP_OP_423J2_125_3477_n1673), .B(
        DP_OP_423J2_125_3477_n1663), .CI(DP_OP_423J2_125_3477_n1665), .CO(
        DP_OP_423J2_125_3477_n1616), .S(DP_OP_423J2_125_3477_n1617) );
  FADDX1_HVT DP_OP_423J2_125_3477_U901 ( .A(DP_OP_423J2_125_3477_n1671), .B(
        DP_OP_423J2_125_3477_n1661), .CI(DP_OP_423J2_125_3477_n1677), .CO(
        DP_OP_423J2_125_3477_n1614), .S(DP_OP_423J2_125_3477_n1615) );
  FADDX1_HVT DP_OP_423J2_125_3477_U900 ( .A(DP_OP_423J2_125_3477_n1679), .B(
        DP_OP_423J2_125_3477_n1667), .CI(DP_OP_423J2_125_3477_n1669), .CO(
        DP_OP_423J2_125_3477_n1612), .S(DP_OP_423J2_125_3477_n1613) );
  FADDX1_HVT DP_OP_423J2_125_3477_U899 ( .A(DP_OP_423J2_125_3477_n1675), .B(
        DP_OP_423J2_125_3477_n1657), .CI(DP_OP_423J2_125_3477_n1655), .CO(
        DP_OP_423J2_125_3477_n1610), .S(DP_OP_423J2_125_3477_n1611) );
  FADDX1_HVT DP_OP_423J2_125_3477_U898 ( .A(DP_OP_423J2_125_3477_n1653), .B(
        DP_OP_423J2_125_3477_n1647), .CI(DP_OP_423J2_125_3477_n1708), .CO(
        DP_OP_423J2_125_3477_n1608), .S(DP_OP_423J2_125_3477_n1609) );
  FADDX1_HVT DP_OP_423J2_125_3477_U897 ( .A(DP_OP_423J2_125_3477_n1651), .B(
        DP_OP_423J2_125_3477_n1649), .CI(DP_OP_423J2_125_3477_n1633), .CO(
        DP_OP_423J2_125_3477_n1606), .S(DP_OP_423J2_125_3477_n1607) );
  FADDX1_HVT DP_OP_423J2_125_3477_U896 ( .A(DP_OP_423J2_125_3477_n1643), .B(
        DP_OP_423J2_125_3477_n1635), .CI(DP_OP_423J2_125_3477_n1631), .CO(
        DP_OP_423J2_125_3477_n1604), .S(DP_OP_423J2_125_3477_n1605) );
  FADDX1_HVT DP_OP_423J2_125_3477_U895 ( .A(DP_OP_423J2_125_3477_n1645), .B(
        DP_OP_423J2_125_3477_n1639), .CI(DP_OP_423J2_125_3477_n1637), .CO(
        DP_OP_423J2_125_3477_n1602), .S(DP_OP_423J2_125_3477_n1603) );
  FADDX1_HVT DP_OP_423J2_125_3477_U894 ( .A(DP_OP_423J2_125_3477_n1641), .B(
        DP_OP_423J2_125_3477_n1706), .CI(DP_OP_423J2_125_3477_n1704), .CO(
        DP_OP_423J2_125_3477_n1600), .S(DP_OP_423J2_125_3477_n1601) );
  FADDX1_HVT DP_OP_423J2_125_3477_U893 ( .A(DP_OP_423J2_125_3477_n1702), .B(
        DP_OP_423J2_125_3477_n1629), .CI(DP_OP_423J2_125_3477_n1700), .CO(
        DP_OP_423J2_125_3477_n1598), .S(DP_OP_423J2_125_3477_n1599) );
  FADDX1_HVT DP_OP_423J2_125_3477_U892 ( .A(DP_OP_423J2_125_3477_n1698), .B(
        DP_OP_423J2_125_3477_n1627), .CI(DP_OP_423J2_125_3477_n1696), .CO(
        DP_OP_423J2_125_3477_n1596), .S(DP_OP_423J2_125_3477_n1597) );
  FADDX1_HVT DP_OP_423J2_125_3477_U891 ( .A(DP_OP_423J2_125_3477_n1625), .B(
        DP_OP_423J2_125_3477_n1623), .CI(DP_OP_423J2_125_3477_n1621), .CO(
        DP_OP_423J2_125_3477_n1594), .S(DP_OP_423J2_125_3477_n1595) );
  FADDX1_HVT DP_OP_423J2_125_3477_U890 ( .A(DP_OP_423J2_125_3477_n1694), .B(
        DP_OP_423J2_125_3477_n1692), .CI(DP_OP_423J2_125_3477_n1619), .CO(
        DP_OP_423J2_125_3477_n1592), .S(DP_OP_423J2_125_3477_n1593) );
  FADDX1_HVT DP_OP_423J2_125_3477_U889 ( .A(DP_OP_423J2_125_3477_n1617), .B(
        DP_OP_423J2_125_3477_n1613), .CI(DP_OP_423J2_125_3477_n1611), .CO(
        DP_OP_423J2_125_3477_n1590), .S(DP_OP_423J2_125_3477_n1591) );
  FADDX1_HVT DP_OP_423J2_125_3477_U888 ( .A(DP_OP_423J2_125_3477_n1615), .B(
        DP_OP_423J2_125_3477_n1609), .CI(DP_OP_423J2_125_3477_n1607), .CO(
        DP_OP_423J2_125_3477_n1588), .S(DP_OP_423J2_125_3477_n1589) );
  FADDX1_HVT DP_OP_423J2_125_3477_U887 ( .A(DP_OP_423J2_125_3477_n1603), .B(
        DP_OP_423J2_125_3477_n1605), .CI(DP_OP_423J2_125_3477_n1690), .CO(
        DP_OP_423J2_125_3477_n1586), .S(DP_OP_423J2_125_3477_n1587) );
  FADDX1_HVT DP_OP_423J2_125_3477_U886 ( .A(DP_OP_423J2_125_3477_n1601), .B(
        DP_OP_423J2_125_3477_n1688), .CI(DP_OP_423J2_125_3477_n1599), .CO(
        DP_OP_423J2_125_3477_n1584), .S(DP_OP_423J2_125_3477_n1585) );
  FADDX1_HVT DP_OP_423J2_125_3477_U885 ( .A(DP_OP_423J2_125_3477_n1686), .B(
        DP_OP_423J2_125_3477_n1597), .CI(DP_OP_423J2_125_3477_n1595), .CO(
        DP_OP_423J2_125_3477_n1582), .S(DP_OP_423J2_125_3477_n1583) );
  FADDX1_HVT DP_OP_423J2_125_3477_U884 ( .A(DP_OP_423J2_125_3477_n1684), .B(
        DP_OP_423J2_125_3477_n1593), .CI(DP_OP_423J2_125_3477_n1591), .CO(
        DP_OP_423J2_125_3477_n1580), .S(DP_OP_423J2_125_3477_n1581) );
  FADDX1_HVT DP_OP_423J2_125_3477_U883 ( .A(DP_OP_423J2_125_3477_n1589), .B(
        DP_OP_423J2_125_3477_n1587), .CI(DP_OP_423J2_125_3477_n1585), .CO(
        DP_OP_423J2_125_3477_n1578), .S(DP_OP_423J2_125_3477_n1579) );
  FADDX1_HVT DP_OP_423J2_125_3477_U882 ( .A(DP_OP_423J2_125_3477_n1682), .B(
        DP_OP_423J2_125_3477_n1583), .CI(DP_OP_423J2_125_3477_n1581), .CO(
        DP_OP_423J2_125_3477_n1576), .S(DP_OP_423J2_125_3477_n1577) );
  FADDX1_HVT DP_OP_423J2_125_3477_U880 ( .A(DP_OP_423J2_125_3477_n2000), .B(
        DP_OP_423J2_125_3477_n2484), .CI(DP_OP_423J2_125_3477_n2745), .CO(
        DP_OP_423J2_125_3477_n1572), .S(DP_OP_423J2_125_3477_n1573) );
  FADDX1_HVT DP_OP_423J2_125_3477_U879 ( .A(DP_OP_423J2_125_3477_n2352), .B(
        DP_OP_423J2_125_3477_n1912), .CI(DP_OP_423J2_125_3477_n1956), .CO(
        DP_OP_423J2_125_3477_n1570), .S(DP_OP_423J2_125_3477_n1571) );
  FADDX1_HVT DP_OP_423J2_125_3477_U878 ( .A(DP_OP_423J2_125_3477_n2308), .B(
        DP_OP_423J2_125_3477_n2044), .CI(DP_OP_423J2_125_3477_n2440), .CO(
        DP_OP_423J2_125_3477_n1568), .S(DP_OP_423J2_125_3477_n1569) );
  FADDX1_HVT DP_OP_423J2_125_3477_U877 ( .A(DP_OP_423J2_125_3477_n2088), .B(
        DP_OP_423J2_125_3477_n2528), .CI(DP_OP_423J2_125_3477_n2176), .CO(
        DP_OP_423J2_125_3477_n1566), .S(DP_OP_423J2_125_3477_n1567) );
  FADDX1_HVT DP_OP_423J2_125_3477_U876 ( .A(DP_OP_423J2_125_3477_n2789), .B(
        DP_OP_423J2_125_3477_n2877), .CI(DP_OP_423J2_125_3477_n2572), .CO(
        DP_OP_423J2_125_3477_n1564), .S(DP_OP_423J2_125_3477_n1565) );
  FADDX1_HVT DP_OP_423J2_125_3477_U875 ( .A(DP_OP_423J2_125_3477_n2132), .B(
        DP_OP_423J2_125_3477_n2264), .CI(DP_OP_423J2_125_3477_n1824), .CO(
        DP_OP_423J2_125_3477_n1562), .S(DP_OP_423J2_125_3477_n1563) );
  FADDX1_HVT DP_OP_423J2_125_3477_U874 ( .A(DP_OP_423J2_125_3477_n2616), .B(
        DP_OP_423J2_125_3477_n2833), .CI(DP_OP_423J2_125_3477_n1868), .CO(
        DP_OP_423J2_125_3477_n1560), .S(DP_OP_423J2_125_3477_n1561) );
  FADDX1_HVT DP_OP_423J2_125_3477_U873 ( .A(DP_OP_423J2_125_3477_n2660), .B(
        DP_OP_423J2_125_3477_n1780), .CI(DP_OP_423J2_125_3477_n2417), .CO(
        DP_OP_423J2_125_3477_n1558), .S(DP_OP_423J2_125_3477_n1559) );
  FADDX1_HVT DP_OP_423J2_125_3477_U872 ( .A(DP_OP_423J2_125_3477_n2461), .B(
        DP_OP_423J2_125_3477_n2396), .CI(DP_OP_423J2_125_3477_n2447), .CO(
        DP_OP_423J2_125_3477_n1556), .S(DP_OP_423J2_125_3477_n1557) );
  FADDX1_HVT DP_OP_423J2_125_3477_U871 ( .A(DP_OP_423J2_125_3477_n2109), .B(
        DP_OP_423J2_125_3477_n2410), .CI(DP_OP_423J2_125_3477_n1889), .CO(
        DP_OP_423J2_125_3477_n1554), .S(DP_OP_423J2_125_3477_n1555) );
  FADDX1_HVT DP_OP_423J2_125_3477_U870 ( .A(DP_OP_423J2_125_3477_n2840), .B(
        DP_OP_423J2_125_3477_n2722), .CI(DP_OP_423J2_125_3477_n2227), .CO(
        DP_OP_423J2_125_3477_n1552), .S(DP_OP_423J2_125_3477_n1553) );
  FADDX1_HVT DP_OP_423J2_125_3477_U869 ( .A(DP_OP_423J2_125_3477_n2884), .B(
        DP_OP_423J2_125_3477_n2535), .CI(DP_OP_423J2_125_3477_n2505), .CO(
        DP_OP_423J2_125_3477_n1550), .S(DP_OP_423J2_125_3477_n1551) );
  FADDX1_HVT DP_OP_423J2_125_3477_U868 ( .A(DP_OP_423J2_125_3477_n2329), .B(
        DP_OP_423J2_125_3477_n2146), .CI(DP_OP_423J2_125_3477_n2854), .CO(
        DP_OP_423J2_125_3477_n1548), .S(DP_OP_423J2_125_3477_n1549) );
  FADDX1_HVT DP_OP_423J2_125_3477_U867 ( .A(DP_OP_423J2_125_3477_n2549), .B(
        DP_OP_423J2_125_3477_n1963), .CI(DP_OP_423J2_125_3477_n2766), .CO(
        DP_OP_423J2_125_3477_n1546), .S(DP_OP_423J2_125_3477_n1547) );
  FADDX1_HVT DP_OP_423J2_125_3477_U866 ( .A(DP_OP_423J2_125_3477_n2637), .B(
        DP_OP_423J2_125_3477_n2220), .CI(DP_OP_423J2_125_3477_n2095), .CO(
        DP_OP_423J2_125_3477_n1544), .S(DP_OP_423J2_125_3477_n1545) );
  FADDX1_HVT DP_OP_423J2_125_3477_U865 ( .A(DP_OP_423J2_125_3477_n2197), .B(
        DP_OP_423J2_125_3477_n1838), .CI(DP_OP_423J2_125_3477_n1575), .CO(
        DP_OP_423J2_125_3477_n1542), .S(DP_OP_423J2_125_3477_n1543) );
  FADDX1_HVT DP_OP_423J2_125_3477_U864 ( .A(DP_OP_423J2_125_3477_n2593), .B(
        DP_OP_423J2_125_3477_n2021), .CI(DP_OP_423J2_125_3477_n2681), .CO(
        DP_OP_423J2_125_3477_n1540), .S(DP_OP_423J2_125_3477_n1541) );
  FADDX1_HVT DP_OP_423J2_125_3477_U863 ( .A(DP_OP_423J2_125_3477_n1845), .B(
        DP_OP_423J2_125_3477_n2752), .CI(DP_OP_423J2_125_3477_n2498), .CO(
        DP_OP_423J2_125_3477_n1538), .S(DP_OP_423J2_125_3477_n1539) );
  FADDX1_HVT DP_OP_423J2_125_3477_U862 ( .A(DP_OP_423J2_125_3477_n1977), .B(
        DP_OP_423J2_125_3477_n2058), .CI(DP_OP_423J2_125_3477_n2586), .CO(
        DP_OP_423J2_125_3477_n1536), .S(DP_OP_423J2_125_3477_n1537) );
  FADDX1_HVT DP_OP_423J2_125_3477_U861 ( .A(DP_OP_423J2_125_3477_n2630), .B(
        DP_OP_423J2_125_3477_n2322), .CI(DP_OP_423J2_125_3477_n2285), .CO(
        DP_OP_423J2_125_3477_n1534), .S(DP_OP_423J2_125_3477_n1535) );
  FADDX1_HVT DP_OP_423J2_125_3477_U860 ( .A(DP_OP_423J2_125_3477_n2271), .B(
        DP_OP_423J2_125_3477_n2359), .CI(DP_OP_423J2_125_3477_n2891), .CO(
        DP_OP_423J2_125_3477_n1532), .S(DP_OP_423J2_125_3477_n1533) );
  FADDX1_HVT DP_OP_423J2_125_3477_U859 ( .A(DP_OP_423J2_125_3477_n2139), .B(
        DP_OP_423J2_125_3477_n2241), .CI(DP_OP_423J2_125_3477_n2803), .CO(
        DP_OP_423J2_125_3477_n1530), .S(DP_OP_423J2_125_3477_n1531) );
  FADDX1_HVT DP_OP_423J2_125_3477_U858 ( .A(DP_OP_423J2_125_3477_n2065), .B(
        DP_OP_423J2_125_3477_n1882), .CI(DP_OP_423J2_125_3477_n2278), .CO(
        DP_OP_423J2_125_3477_n1528), .S(DP_OP_423J2_125_3477_n1529) );
  FADDX1_HVT DP_OP_423J2_125_3477_U857 ( .A(DP_OP_423J2_125_3477_n2579), .B(
        DP_OP_423J2_125_3477_n2454), .CI(DP_OP_423J2_125_3477_n2898), .CO(
        DP_OP_423J2_125_3477_n1526), .S(DP_OP_423J2_125_3477_n1527) );
  FADDX1_HVT DP_OP_423J2_125_3477_U856 ( .A(DP_OP_423J2_125_3477_n2674), .B(
        DP_OP_423J2_125_3477_n2491), .CI(DP_OP_423J2_125_3477_n2759), .CO(
        DP_OP_423J2_125_3477_n1524), .S(DP_OP_423J2_125_3477_n1525) );
  FADDX1_HVT DP_OP_423J2_125_3477_U855 ( .A(DP_OP_423J2_125_3477_n2102), .B(
        DP_OP_423J2_125_3477_n2667), .CI(DP_OP_423J2_125_3477_n2373), .CO(
        DP_OP_423J2_125_3477_n1522), .S(DP_OP_423J2_125_3477_n1523) );
  FADDX1_HVT DP_OP_423J2_125_3477_U854 ( .A(DP_OP_423J2_125_3477_n2708), .B(
        DP_OP_423J2_125_3477_n2715), .CI(DP_OP_423J2_125_3477_n2810), .CO(
        DP_OP_423J2_125_3477_n1520), .S(DP_OP_423J2_125_3477_n1521) );
  FADDX1_HVT DP_OP_423J2_125_3477_U853 ( .A(DP_OP_423J2_125_3477_n2542), .B(
        DP_OP_423J2_125_3477_n2007), .CI(DP_OP_423J2_125_3477_n1831), .CO(
        DP_OP_423J2_125_3477_n1518), .S(DP_OP_423J2_125_3477_n1519) );
  FADDX1_HVT DP_OP_423J2_125_3477_U852 ( .A(DP_OP_423J2_125_3477_n2315), .B(
        DP_OP_423J2_125_3477_n2234), .CI(DP_OP_423J2_125_3477_n1919), .CO(
        DP_OP_423J2_125_3477_n1516), .S(DP_OP_423J2_125_3477_n1517) );
  FADDX1_HVT DP_OP_423J2_125_3477_U851 ( .A(DP_OP_423J2_125_3477_n2051), .B(
        DP_OP_423J2_125_3477_n2190), .CI(DP_OP_423J2_125_3477_n2183), .CO(
        DP_OP_423J2_125_3477_n1514), .S(DP_OP_423J2_125_3477_n1515) );
  FADDX1_HVT DP_OP_423J2_125_3477_U850 ( .A(DP_OP_423J2_125_3477_n1933), .B(
        DP_OP_423J2_125_3477_n2366), .CI(DP_OP_423J2_125_3477_n1970), .CO(
        DP_OP_423J2_125_3477_n1512), .S(DP_OP_423J2_125_3477_n1513) );
  FADDX1_HVT DP_OP_423J2_125_3477_U849 ( .A(DP_OP_423J2_125_3477_n2847), .B(
        DP_OP_423J2_125_3477_n1926), .CI(DP_OP_423J2_125_3477_n2623), .CO(
        DP_OP_423J2_125_3477_n1510), .S(DP_OP_423J2_125_3477_n1511) );
  FADDX1_HVT DP_OP_423J2_125_3477_U848 ( .A(DP_OP_423J2_125_3477_n2403), .B(
        DP_OP_423J2_125_3477_n1875), .CI(DP_OP_423J2_125_3477_n2796), .CO(
        DP_OP_423J2_125_3477_n1508), .S(DP_OP_423J2_125_3477_n1509) );
  FADDX1_HVT DP_OP_423J2_125_3477_U847 ( .A(DP_OP_423J2_125_3477_n2153), .B(
        DP_OP_423J2_125_3477_n2014), .CI(DP_OP_423J2_125_3477_n1680), .CO(
        DP_OP_423J2_125_3477_n1506), .S(DP_OP_423J2_125_3477_n1507) );
  FADDX1_HVT DP_OP_423J2_125_3477_U846 ( .A(DP_OP_423J2_125_3477_n1678), .B(
        DP_OP_423J2_125_3477_n1658), .CI(DP_OP_423J2_125_3477_n1660), .CO(
        DP_OP_423J2_125_3477_n1504), .S(DP_OP_423J2_125_3477_n1505) );
  FADDX1_HVT DP_OP_423J2_125_3477_U845 ( .A(DP_OP_423J2_125_3477_n1676), .B(
        DP_OP_423J2_125_3477_n1662), .CI(DP_OP_423J2_125_3477_n1664), .CO(
        DP_OP_423J2_125_3477_n1502), .S(DP_OP_423J2_125_3477_n1503) );
  FADDX1_HVT DP_OP_423J2_125_3477_U844 ( .A(DP_OP_423J2_125_3477_n1674), .B(
        DP_OP_423J2_125_3477_n1666), .CI(DP_OP_423J2_125_3477_n1668), .CO(
        DP_OP_423J2_125_3477_n1500), .S(DP_OP_423J2_125_3477_n1501) );
  FADDX1_HVT DP_OP_423J2_125_3477_U843 ( .A(DP_OP_423J2_125_3477_n1672), .B(
        DP_OP_423J2_125_3477_n1670), .CI(DP_OP_423J2_125_3477_n1656), .CO(
        DP_OP_423J2_125_3477_n1498), .S(DP_OP_423J2_125_3477_n1499) );
  FADDX1_HVT DP_OP_423J2_125_3477_U842 ( .A(DP_OP_423J2_125_3477_n1654), .B(
        DP_OP_423J2_125_3477_n1646), .CI(DP_OP_423J2_125_3477_n1632), .CO(
        DP_OP_423J2_125_3477_n1496), .S(DP_OP_423J2_125_3477_n1497) );
  FADDX1_HVT DP_OP_423J2_125_3477_U841 ( .A(DP_OP_423J2_125_3477_n1652), .B(
        DP_OP_423J2_125_3477_n1648), .CI(DP_OP_423J2_125_3477_n1634), .CO(
        DP_OP_423J2_125_3477_n1494), .S(DP_OP_423J2_125_3477_n1495) );
  FADDX1_HVT DP_OP_423J2_125_3477_U840 ( .A(DP_OP_423J2_125_3477_n1650), .B(
        DP_OP_423J2_125_3477_n1561), .CI(DP_OP_423J2_125_3477_n1636), .CO(
        DP_OP_423J2_125_3477_n1492), .S(DP_OP_423J2_125_3477_n1493) );
  FADDX1_HVT DP_OP_423J2_125_3477_U839 ( .A(DP_OP_423J2_125_3477_n1573), .B(
        DP_OP_423J2_125_3477_n1638), .CI(DP_OP_423J2_125_3477_n1630), .CO(
        DP_OP_423J2_125_3477_n1490), .S(DP_OP_423J2_125_3477_n1491) );
  FADDX1_HVT DP_OP_423J2_125_3477_U838 ( .A(DP_OP_423J2_125_3477_n1571), .B(
        DP_OP_423J2_125_3477_n1640), .CI(DP_OP_423J2_125_3477_n1559), .CO(
        DP_OP_423J2_125_3477_n1488), .S(DP_OP_423J2_125_3477_n1489) );
  FADDX1_HVT DP_OP_423J2_125_3477_U837 ( .A(DP_OP_423J2_125_3477_n1569), .B(
        DP_OP_423J2_125_3477_n1644), .CI(DP_OP_423J2_125_3477_n1642), .CO(
        DP_OP_423J2_125_3477_n1486), .S(DP_OP_423J2_125_3477_n1487) );
  FADDX1_HVT DP_OP_423J2_125_3477_U836 ( .A(DP_OP_423J2_125_3477_n1563), .B(
        DP_OP_423J2_125_3477_n1565), .CI(DP_OP_423J2_125_3477_n1567), .CO(
        DP_OP_423J2_125_3477_n1484), .S(DP_OP_423J2_125_3477_n1485) );
  FADDX1_HVT DP_OP_423J2_125_3477_U835 ( .A(DP_OP_423J2_125_3477_n1551), .B(
        DP_OP_423J2_125_3477_n1537), .CI(DP_OP_423J2_125_3477_n1535), .CO(
        DP_OP_423J2_125_3477_n1482), .S(DP_OP_423J2_125_3477_n1483) );
  FADDX1_HVT DP_OP_423J2_125_3477_U834 ( .A(DP_OP_423J2_125_3477_n1555), .B(
        DP_OP_423J2_125_3477_n1545), .CI(DP_OP_423J2_125_3477_n1543), .CO(
        DP_OP_423J2_125_3477_n1480), .S(DP_OP_423J2_125_3477_n1481) );
  FADDX1_HVT DP_OP_423J2_125_3477_U833 ( .A(DP_OP_423J2_125_3477_n1547), .B(
        DP_OP_423J2_125_3477_n1539), .CI(DP_OP_423J2_125_3477_n1557), .CO(
        DP_OP_423J2_125_3477_n1478), .S(DP_OP_423J2_125_3477_n1479) );
  FADDX1_HVT DP_OP_423J2_125_3477_U832 ( .A(DP_OP_423J2_125_3477_n1541), .B(
        DP_OP_423J2_125_3477_n1553), .CI(DP_OP_423J2_125_3477_n1549), .CO(
        DP_OP_423J2_125_3477_n1476), .S(DP_OP_423J2_125_3477_n1477) );
  FADDX1_HVT DP_OP_423J2_125_3477_U831 ( .A(DP_OP_423J2_125_3477_n1531), .B(
        DP_OP_423J2_125_3477_n1523), .CI(DP_OP_423J2_125_3477_n1509), .CO(
        DP_OP_423J2_125_3477_n1474), .S(DP_OP_423J2_125_3477_n1475) );
  FADDX1_HVT DP_OP_423J2_125_3477_U830 ( .A(DP_OP_423J2_125_3477_n1529), .B(
        DP_OP_423J2_125_3477_n1525), .CI(DP_OP_423J2_125_3477_n1511), .CO(
        DP_OP_423J2_125_3477_n1472), .S(DP_OP_423J2_125_3477_n1473) );
  FADDX1_HVT DP_OP_423J2_125_3477_U829 ( .A(DP_OP_423J2_125_3477_n1533), .B(
        DP_OP_423J2_125_3477_n1527), .CI(DP_OP_423J2_125_3477_n1513), .CO(
        DP_OP_423J2_125_3477_n1470), .S(DP_OP_423J2_125_3477_n1471) );
  FADDX1_HVT DP_OP_423J2_125_3477_U828 ( .A(DP_OP_423J2_125_3477_n1519), .B(
        DP_OP_423J2_125_3477_n1515), .CI(DP_OP_423J2_125_3477_n1507), .CO(
        DP_OP_423J2_125_3477_n1468), .S(DP_OP_423J2_125_3477_n1469) );
  FADDX1_HVT DP_OP_423J2_125_3477_U827 ( .A(DP_OP_423J2_125_3477_n1521), .B(
        DP_OP_423J2_125_3477_n1517), .CI(DP_OP_423J2_125_3477_n1628), .CO(
        DP_OP_423J2_125_3477_n1466), .S(DP_OP_423J2_125_3477_n1467) );
  FADDX1_HVT DP_OP_423J2_125_3477_U826 ( .A(DP_OP_423J2_125_3477_n1626), .B(
        DP_OP_423J2_125_3477_n1624), .CI(DP_OP_423J2_125_3477_n1622), .CO(
        DP_OP_423J2_125_3477_n1464), .S(DP_OP_423J2_125_3477_n1465) );
  FADDX1_HVT DP_OP_423J2_125_3477_U825 ( .A(DP_OP_423J2_125_3477_n1620), .B(
        DP_OP_423J2_125_3477_n1618), .CI(DP_OP_423J2_125_3477_n1616), .CO(
        DP_OP_423J2_125_3477_n1462), .S(DP_OP_423J2_125_3477_n1463) );
  FADDX1_HVT DP_OP_423J2_125_3477_U824 ( .A(DP_OP_423J2_125_3477_n1503), .B(
        DP_OP_423J2_125_3477_n1499), .CI(DP_OP_423J2_125_3477_n1610), .CO(
        DP_OP_423J2_125_3477_n1460), .S(DP_OP_423J2_125_3477_n1461) );
  FADDX1_HVT DP_OP_423J2_125_3477_U823 ( .A(DP_OP_423J2_125_3477_n1614), .B(
        DP_OP_423J2_125_3477_n1612), .CI(DP_OP_423J2_125_3477_n1501), .CO(
        DP_OP_423J2_125_3477_n1458), .S(DP_OP_423J2_125_3477_n1459) );
  FADDX1_HVT DP_OP_423J2_125_3477_U822 ( .A(DP_OP_423J2_125_3477_n1505), .B(
        DP_OP_423J2_125_3477_n1608), .CI(DP_OP_423J2_125_3477_n1497), .CO(
        DP_OP_423J2_125_3477_n1456), .S(DP_OP_423J2_125_3477_n1457) );
  FADDX1_HVT DP_OP_423J2_125_3477_U821 ( .A(DP_OP_423J2_125_3477_n1495), .B(
        DP_OP_423J2_125_3477_n1606), .CI(DP_OP_423J2_125_3477_n1604), .CO(
        DP_OP_423J2_125_3477_n1454), .S(DP_OP_423J2_125_3477_n1455) );
  FADDX1_HVT DP_OP_423J2_125_3477_U820 ( .A(DP_OP_423J2_125_3477_n1493), .B(
        DP_OP_423J2_125_3477_n1489), .CI(DP_OP_423J2_125_3477_n1602), .CO(
        DP_OP_423J2_125_3477_n1452), .S(DP_OP_423J2_125_3477_n1453) );
  FADDX1_HVT DP_OP_423J2_125_3477_U819 ( .A(DP_OP_423J2_125_3477_n1491), .B(
        DP_OP_423J2_125_3477_n1487), .CI(DP_OP_423J2_125_3477_n1485), .CO(
        DP_OP_423J2_125_3477_n1450), .S(DP_OP_423J2_125_3477_n1451) );
  FADDX1_HVT DP_OP_423J2_125_3477_U818 ( .A(DP_OP_423J2_125_3477_n1479), .B(
        DP_OP_423J2_125_3477_n1477), .CI(DP_OP_423J2_125_3477_n1600), .CO(
        DP_OP_423J2_125_3477_n1448), .S(DP_OP_423J2_125_3477_n1449) );
  FADDX1_HVT DP_OP_423J2_125_3477_U817 ( .A(DP_OP_423J2_125_3477_n1483), .B(
        DP_OP_423J2_125_3477_n1481), .CI(DP_OP_423J2_125_3477_n1475), .CO(
        DP_OP_423J2_125_3477_n1446), .S(DP_OP_423J2_125_3477_n1447) );
  FADDX1_HVT DP_OP_423J2_125_3477_U816 ( .A(DP_OP_423J2_125_3477_n1471), .B(
        DP_OP_423J2_125_3477_n1473), .CI(DP_OP_423J2_125_3477_n1469), .CO(
        DP_OP_423J2_125_3477_n1444), .S(DP_OP_423J2_125_3477_n1445) );
  FADDX1_HVT DP_OP_423J2_125_3477_U815 ( .A(DP_OP_423J2_125_3477_n1467), .B(
        DP_OP_423J2_125_3477_n1598), .CI(DP_OP_423J2_125_3477_n1596), .CO(
        DP_OP_423J2_125_3477_n1442), .S(DP_OP_423J2_125_3477_n1443) );
  FADDX1_HVT DP_OP_423J2_125_3477_U814 ( .A(DP_OP_423J2_125_3477_n1465), .B(
        DP_OP_423J2_125_3477_n1594), .CI(DP_OP_423J2_125_3477_n1592), .CO(
        DP_OP_423J2_125_3477_n1440), .S(DP_OP_423J2_125_3477_n1441) );
  FADDX1_HVT DP_OP_423J2_125_3477_U813 ( .A(DP_OP_423J2_125_3477_n1463), .B(
        DP_OP_423J2_125_3477_n1459), .CI(DP_OP_423J2_125_3477_n1461), .CO(
        DP_OP_423J2_125_3477_n1438), .S(DP_OP_423J2_125_3477_n1439) );
  FADDX1_HVT DP_OP_423J2_125_3477_U812 ( .A(DP_OP_423J2_125_3477_n1590), .B(
        DP_OP_423J2_125_3477_n1588), .CI(DP_OP_423J2_125_3477_n1457), .CO(
        DP_OP_423J2_125_3477_n1436), .S(DP_OP_423J2_125_3477_n1437) );
  FADDX1_HVT DP_OP_423J2_125_3477_U811 ( .A(DP_OP_423J2_125_3477_n1455), .B(
        DP_OP_423J2_125_3477_n1453), .CI(DP_OP_423J2_125_3477_n1586), .CO(
        DP_OP_423J2_125_3477_n1434), .S(DP_OP_423J2_125_3477_n1435) );
  FADDX1_HVT DP_OP_423J2_125_3477_U810 ( .A(DP_OP_423J2_125_3477_n1451), .B(
        DP_OP_423J2_125_3477_n1449), .CI(DP_OP_423J2_125_3477_n1447), .CO(
        DP_OP_423J2_125_3477_n1432), .S(DP_OP_423J2_125_3477_n1433) );
  FADDX1_HVT DP_OP_423J2_125_3477_U809 ( .A(DP_OP_423J2_125_3477_n1445), .B(
        DP_OP_423J2_125_3477_n1584), .CI(DP_OP_423J2_125_3477_n1443), .CO(
        DP_OP_423J2_125_3477_n1430), .S(DP_OP_423J2_125_3477_n1431) );
  FADDX1_HVT DP_OP_423J2_125_3477_U808 ( .A(DP_OP_423J2_125_3477_n1582), .B(
        DP_OP_423J2_125_3477_n1441), .CI(DP_OP_423J2_125_3477_n1580), .CO(
        DP_OP_423J2_125_3477_n1428), .S(DP_OP_423J2_125_3477_n1429) );
  FADDX1_HVT DP_OP_423J2_125_3477_U807 ( .A(DP_OP_423J2_125_3477_n1439), .B(
        DP_OP_423J2_125_3477_n1437), .CI(DP_OP_423J2_125_3477_n1435), .CO(
        DP_OP_423J2_125_3477_n1426), .S(DP_OP_423J2_125_3477_n1427) );
  FADDX1_HVT DP_OP_423J2_125_3477_U806 ( .A(DP_OP_423J2_125_3477_n1433), .B(
        DP_OP_423J2_125_3477_n1578), .CI(DP_OP_423J2_125_3477_n1431), .CO(
        DP_OP_423J2_125_3477_n1424), .S(DP_OP_423J2_125_3477_n1425) );
  FADDX1_HVT DP_OP_423J2_125_3477_U805 ( .A(DP_OP_423J2_125_3477_n1576), .B(
        DP_OP_423J2_125_3477_n1429), .CI(DP_OP_423J2_125_3477_n1427), .CO(
        DP_OP_423J2_125_3477_n1422), .S(DP_OP_423J2_125_3477_n1423) );
  FADDX1_HVT DP_OP_423J2_125_3477_U804 ( .A(DP_OP_423J2_125_3477_n1574), .B(
        DP_OP_423J2_125_3477_n2527), .CI(DP_OP_423J2_125_3477_n2744), .CO(
        DP_OP_423J2_125_3477_n1420), .S(DP_OP_423J2_125_3477_n1421) );
  FADDX1_HVT DP_OP_423J2_125_3477_U803 ( .A(DP_OP_423J2_125_3477_n1999), .B(
        DP_OP_423J2_125_3477_n1911), .CI(DP_OP_423J2_125_3477_n1955), .CO(
        DP_OP_423J2_125_3477_n1418), .S(DP_OP_423J2_125_3477_n1419) );
  FADDX1_HVT DP_OP_423J2_125_3477_U802 ( .A(DP_OP_423J2_125_3477_n2701), .B(
        DP_OP_423J2_125_3477_n2439), .CI(DP_OP_423J2_125_3477_n2571), .CO(
        DP_OP_423J2_125_3477_n1416), .S(DP_OP_423J2_125_3477_n1417) );
  FADDX1_HVT DP_OP_423J2_125_3477_U801 ( .A(DP_OP_423J2_125_3477_n2832), .B(
        DP_OP_423J2_125_3477_n2175), .CI(DP_OP_423J2_125_3477_n2483), .CO(
        DP_OP_423J2_125_3477_n1414), .S(DP_OP_423J2_125_3477_n1415) );
  FADDX1_HVT DP_OP_423J2_125_3477_U800 ( .A(DP_OP_423J2_125_3477_n1867), .B(
        DP_OP_423J2_125_3477_n2876), .CI(DP_OP_423J2_125_3477_n2043), .CO(
        DP_OP_423J2_125_3477_n1412), .S(DP_OP_423J2_125_3477_n1413) );
  FADDX1_HVT DP_OP_423J2_125_3477_U799 ( .A(DP_OP_423J2_125_3477_n2131), .B(
        DP_OP_423J2_125_3477_n2263), .CI(DP_OP_423J2_125_3477_n1823), .CO(
        DP_OP_423J2_125_3477_n1410), .S(DP_OP_423J2_125_3477_n1411) );
  FADDX1_HVT DP_OP_423J2_125_3477_U798 ( .A(DP_OP_423J2_125_3477_n2087), .B(
        DP_OP_423J2_125_3477_n2615), .CI(DP_OP_423J2_125_3477_n2351), .CO(
        DP_OP_423J2_125_3477_n1408), .S(DP_OP_423J2_125_3477_n1409) );
  FADDX1_HVT DP_OP_423J2_125_3477_U797 ( .A(DP_OP_423J2_125_3477_n2307), .B(
        DP_OP_423J2_125_3477_n2788), .CI(DP_OP_423J2_125_3477_n2659), .CO(
        DP_OP_423J2_125_3477_n1406), .S(DP_OP_423J2_125_3477_n1407) );
  FADDX1_HVT DP_OP_423J2_125_3477_U796 ( .A(DP_OP_423J2_125_3477_n1779), .B(
        DP_OP_423J2_125_3477_n2395), .CI(DP_OP_423J2_125_3477_n2226), .CO(
        DP_OP_423J2_125_3477_n1404), .S(DP_OP_423J2_125_3477_n1405) );
  FADDX1_HVT DP_OP_423J2_125_3477_U795 ( .A(DP_OP_423J2_125_3477_n2460), .B(
        DP_OP_423J2_125_3477_n2145), .CI(DP_OP_423J2_125_3477_n2853), .CO(
        DP_OP_423J2_125_3477_n1402), .S(DP_OP_423J2_125_3477_n1403) );
  FADDX1_HVT DP_OP_423J2_125_3477_U794 ( .A(DP_OP_423J2_125_3477_n2883), .B(
        DP_OP_423J2_125_3477_n2409), .CI(DP_OP_423J2_125_3477_n2765), .CO(
        DP_OP_423J2_125_3477_n1400), .S(DP_OP_423J2_125_3477_n1401) );
  FADDX1_HVT DP_OP_423J2_125_3477_U793 ( .A(DP_OP_423J2_125_3477_n2196), .B(
        DP_OP_423J2_125_3477_n2721), .CI(DP_OP_423J2_125_3477_n1888), .CO(
        DP_OP_423J2_125_3477_n1398), .S(DP_OP_423J2_125_3477_n1399) );
  FADDX1_HVT DP_OP_423J2_125_3477_U792 ( .A(DP_OP_423J2_125_3477_n2328), .B(
        DP_OP_423J2_125_3477_n1962), .CI(DP_OP_423J2_125_3477_n2504), .CO(
        DP_OP_423J2_125_3477_n1396), .S(DP_OP_423J2_125_3477_n1397) );
  FADDX1_HVT DP_OP_423J2_125_3477_U791 ( .A(DP_OP_423J2_125_3477_n2416), .B(
        DP_OP_423J2_125_3477_n2534), .CI(DP_OP_423J2_125_3477_n2446), .CO(
        DP_OP_423J2_125_3477_n1394), .S(DP_OP_423J2_125_3477_n1395) );
  FADDX1_HVT DP_OP_423J2_125_3477_U790 ( .A(DP_OP_423J2_125_3477_n2636), .B(
        DP_OP_423J2_125_3477_n2219), .CI(DP_OP_423J2_125_3477_n2094), .CO(
        DP_OP_423J2_125_3477_n1392), .S(DP_OP_423J2_125_3477_n1393) );
  FADDX1_HVT DP_OP_423J2_125_3477_U789 ( .A(DP_OP_423J2_125_3477_n2592), .B(
        DP_OP_423J2_125_3477_n1976), .CI(DP_OP_423J2_125_3477_n2057), .CO(
        DP_OP_423J2_125_3477_n1390), .S(DP_OP_423J2_125_3477_n1391) );
  FADDX1_HVT DP_OP_423J2_125_3477_U788 ( .A(DP_OP_423J2_125_3477_n2108), .B(
        DP_OP_423J2_125_3477_n2751), .CI(DP_OP_423J2_125_3477_n2629), .CO(
        DP_OP_423J2_125_3477_n1388), .S(DP_OP_423J2_125_3477_n1389) );
  FADDX1_HVT DP_OP_423J2_125_3477_U787 ( .A(DP_OP_423J2_125_3477_n1844), .B(
        DP_OP_423J2_125_3477_n2680), .CI(DP_OP_423J2_125_3477_n2585), .CO(
        DP_OP_423J2_125_3477_n1386), .S(DP_OP_423J2_125_3477_n1387) );
  FADDX1_HVT DP_OP_423J2_125_3477_U786 ( .A(DP_OP_423J2_125_3477_n2548), .B(
        DP_OP_423J2_125_3477_n2020), .CI(DP_OP_423J2_125_3477_n1837), .CO(
        DP_OP_423J2_125_3477_n1384), .S(DP_OP_423J2_125_3477_n1385) );
  FADDX1_HVT DP_OP_423J2_125_3477_U785 ( .A(DP_OP_423J2_125_3477_n2839), .B(
        DP_OP_423J2_125_3477_n2321), .CI(DP_OP_423J2_125_3477_n2497), .CO(
        DP_OP_423J2_125_3477_n1382), .S(DP_OP_423J2_125_3477_n1383) );
  FADDX1_HVT DP_OP_423J2_125_3477_U784 ( .A(DP_OP_423J2_125_3477_n2284), .B(
        DP_OP_423J2_125_3477_n2358), .CI(DP_OP_423J2_125_3477_n2890), .CO(
        DP_OP_423J2_125_3477_n1380), .S(DP_OP_423J2_125_3477_n1381) );
  FADDX1_HVT DP_OP_423J2_125_3477_U783 ( .A(DP_OP_423J2_125_3477_n2064), .B(
        DP_OP_423J2_125_3477_n2240), .CI(DP_OP_423J2_125_3477_n2277), .CO(
        DP_OP_423J2_125_3477_n1378), .S(DP_OP_423J2_125_3477_n1379) );
  FADDX1_HVT DP_OP_423J2_125_3477_U782 ( .A(DP_OP_423J2_125_3477_n2270), .B(
        DP_OP_423J2_125_3477_n2101), .CI(DP_OP_423J2_125_3477_n2802), .CO(
        DP_OP_423J2_125_3477_n1376), .S(DP_OP_423J2_125_3477_n1377) );
  FADDX1_HVT DP_OP_423J2_125_3477_U781 ( .A(DP_OP_423J2_125_3477_n2138), .B(
        DP_OP_423J2_125_3477_n1881), .CI(DP_OP_423J2_125_3477_n1925), .CO(
        DP_OP_423J2_125_3477_n1374), .S(DP_OP_423J2_125_3477_n1375) );
  FADDX1_HVT DP_OP_423J2_125_3477_U780 ( .A(DP_OP_423J2_125_3477_n2578), .B(
        DP_OP_423J2_125_3477_n2453), .CI(DP_OP_423J2_125_3477_n2897), .CO(
        DP_OP_423J2_125_3477_n1372), .S(DP_OP_423J2_125_3477_n1373) );
  FADDX1_HVT DP_OP_423J2_125_3477_U779 ( .A(DP_OP_423J2_125_3477_n2673), .B(
        DP_OP_423J2_125_3477_n2490), .CI(DP_OP_423J2_125_3477_n2758), .CO(
        DP_OP_423J2_125_3477_n1370), .S(DP_OP_423J2_125_3477_n1371) );
  FADDX1_HVT DP_OP_423J2_125_3477_U778 ( .A(DP_OP_423J2_125_3477_n2666), .B(
        DP_OP_423J2_125_3477_n2402), .CI(DP_OP_423J2_125_3477_n2809), .CO(
        DP_OP_423J2_125_3477_n1368), .S(DP_OP_423J2_125_3477_n1369) );
  FADDX1_HVT DP_OP_423J2_125_3477_U777 ( .A(DP_OP_423J2_125_3477_n2707), .B(
        DP_OP_423J2_125_3477_n2714), .CI(DP_OP_423J2_125_3477_n1830), .CO(
        DP_OP_423J2_125_3477_n1366), .S(DP_OP_423J2_125_3477_n1367) );
  FADDX1_HVT DP_OP_423J2_125_3477_U776 ( .A(DP_OP_423J2_125_3477_n2541), .B(
        DP_OP_423J2_125_3477_n2372), .CI(DP_OP_423J2_125_3477_n2182), .CO(
        DP_OP_423J2_125_3477_n1364), .S(DP_OP_423J2_125_3477_n1365) );
  FADDX1_HVT DP_OP_423J2_125_3477_U775 ( .A(DP_OP_423J2_125_3477_n2050), .B(
        DP_OP_423J2_125_3477_n2365), .CI(DP_OP_423J2_125_3477_n1918), .CO(
        DP_OP_423J2_125_3477_n1362), .S(DP_OP_423J2_125_3477_n1363) );
  FADDX1_HVT DP_OP_423J2_125_3477_U774 ( .A(DP_OP_423J2_125_3477_n2314), .B(
        DP_OP_423J2_125_3477_n2006), .CI(DP_OP_423J2_125_3477_n1969), .CO(
        DP_OP_423J2_125_3477_n1360), .S(DP_OP_423J2_125_3477_n1361) );
  FADDX1_HVT DP_OP_423J2_125_3477_U773 ( .A(DP_OP_423J2_125_3477_n1932), .B(
        DP_OP_423J2_125_3477_n2189), .CI(DP_OP_423J2_125_3477_n2622), .CO(
        DP_OP_423J2_125_3477_n1358), .S(DP_OP_423J2_125_3477_n1359) );
  FADDX1_HVT DP_OP_423J2_125_3477_U772 ( .A(DP_OP_423J2_125_3477_n2846), .B(
        DP_OP_423J2_125_3477_n2233), .CI(DP_OP_423J2_125_3477_n2795), .CO(
        DP_OP_423J2_125_3477_n1356), .S(DP_OP_423J2_125_3477_n1357) );
  FADDX1_HVT DP_OP_423J2_125_3477_U771 ( .A(DP_OP_423J2_125_3477_n2152), .B(
        DP_OP_423J2_125_3477_n2013), .CI(DP_OP_423J2_125_3477_n1874), .CO(
        DP_OP_423J2_125_3477_n1354), .S(DP_OP_423J2_125_3477_n1355) );
  FADDX1_HVT DP_OP_423J2_125_3477_U770 ( .A(DP_OP_423J2_125_3477_n1572), .B(
        DP_OP_423J2_125_3477_n1570), .CI(DP_OP_423J2_125_3477_n1558), .CO(
        DP_OP_423J2_125_3477_n1352), .S(DP_OP_423J2_125_3477_n1353) );
  FADDX1_HVT DP_OP_423J2_125_3477_U769 ( .A(DP_OP_423J2_125_3477_n1560), .B(
        DP_OP_423J2_125_3477_n1568), .CI(DP_OP_423J2_125_3477_n1566), .CO(
        DP_OP_423J2_125_3477_n1350), .S(DP_OP_423J2_125_3477_n1351) );
  FADDX1_HVT DP_OP_423J2_125_3477_U768 ( .A(DP_OP_423J2_125_3477_n1564), .B(
        DP_OP_423J2_125_3477_n1562), .CI(DP_OP_423J2_125_3477_n1556), .CO(
        DP_OP_423J2_125_3477_n1348), .S(DP_OP_423J2_125_3477_n1349) );
  FADDX1_HVT DP_OP_423J2_125_3477_U767 ( .A(DP_OP_423J2_125_3477_n1554), .B(
        DP_OP_423J2_125_3477_n1534), .CI(DP_OP_423J2_125_3477_n1536), .CO(
        DP_OP_423J2_125_3477_n1346), .S(DP_OP_423J2_125_3477_n1347) );
  FADDX1_HVT DP_OP_423J2_125_3477_U766 ( .A(DP_OP_423J2_125_3477_n1552), .B(
        DP_OP_423J2_125_3477_n1538), .CI(DP_OP_423J2_125_3477_n1540), .CO(
        DP_OP_423J2_125_3477_n1344), .S(DP_OP_423J2_125_3477_n1345) );
  FADDX1_HVT DP_OP_423J2_125_3477_U765 ( .A(DP_OP_423J2_125_3477_n1550), .B(
        DP_OP_423J2_125_3477_n1542), .CI(DP_OP_423J2_125_3477_n1544), .CO(
        DP_OP_423J2_125_3477_n1342), .S(DP_OP_423J2_125_3477_n1343) );
  FADDX1_HVT DP_OP_423J2_125_3477_U764 ( .A(DP_OP_423J2_125_3477_n1548), .B(
        DP_OP_423J2_125_3477_n1546), .CI(DP_OP_423J2_125_3477_n1532), .CO(
        DP_OP_423J2_125_3477_n1340), .S(DP_OP_423J2_125_3477_n1341) );
  FADDX1_HVT DP_OP_423J2_125_3477_U763 ( .A(DP_OP_423J2_125_3477_n1530), .B(
        DP_OP_423J2_125_3477_n1522), .CI(DP_OP_423J2_125_3477_n1508), .CO(
        DP_OP_423J2_125_3477_n1338), .S(DP_OP_423J2_125_3477_n1339) );
  FADDX1_HVT DP_OP_423J2_125_3477_U762 ( .A(DP_OP_423J2_125_3477_n1528), .B(
        DP_OP_423J2_125_3477_n1524), .CI(DP_OP_423J2_125_3477_n1510), .CO(
        DP_OP_423J2_125_3477_n1336), .S(DP_OP_423J2_125_3477_n1337) );
  FADDX1_HVT DP_OP_423J2_125_3477_U761 ( .A(DP_OP_423J2_125_3477_n1526), .B(
        DP_OP_423J2_125_3477_n1407), .CI(DP_OP_423J2_125_3477_n1512), .CO(
        DP_OP_423J2_125_3477_n1334), .S(DP_OP_423J2_125_3477_n1335) );
  FADDX1_HVT DP_OP_423J2_125_3477_U760 ( .A(DP_OP_423J2_125_3477_n1417), .B(
        DP_OP_423J2_125_3477_n1514), .CI(DP_OP_423J2_125_3477_n1506), .CO(
        DP_OP_423J2_125_3477_n1332), .S(DP_OP_423J2_125_3477_n1333) );
  FADDX1_HVT DP_OP_423J2_125_3477_U759 ( .A(DP_OP_423J2_125_3477_n1419), .B(
        DP_OP_423J2_125_3477_n1518), .CI(DP_OP_423J2_125_3477_n1516), .CO(
        DP_OP_423J2_125_3477_n1330), .S(DP_OP_423J2_125_3477_n1331) );
  FADDX1_HVT DP_OP_423J2_125_3477_U758 ( .A(DP_OP_423J2_125_3477_n1421), .B(
        DP_OP_423J2_125_3477_n1415), .CI(DP_OP_423J2_125_3477_n1520), .CO(
        DP_OP_423J2_125_3477_n1328), .S(DP_OP_423J2_125_3477_n1329) );
  FADDX1_HVT DP_OP_423J2_125_3477_U757 ( .A(DP_OP_423J2_125_3477_n1413), .B(
        DP_OP_423J2_125_3477_n1411), .CI(DP_OP_423J2_125_3477_n1409), .CO(
        DP_OP_423J2_125_3477_n1326), .S(DP_OP_423J2_125_3477_n1327) );
  FADDX1_HVT DP_OP_423J2_125_3477_U756 ( .A(DP_OP_423J2_125_3477_n1405), .B(
        DP_OP_423J2_125_3477_n1383), .CI(DP_OP_423J2_125_3477_n1393), .CO(
        DP_OP_423J2_125_3477_n1324), .S(DP_OP_423J2_125_3477_n1325) );
  FADDX1_HVT DP_OP_423J2_125_3477_U755 ( .A(DP_OP_423J2_125_3477_n1397), .B(
        DP_OP_423J2_125_3477_n1391), .CI(DP_OP_423J2_125_3477_n1385), .CO(
        DP_OP_423J2_125_3477_n1322), .S(DP_OP_423J2_125_3477_n1323) );
  FADDX1_HVT DP_OP_423J2_125_3477_U754 ( .A(DP_OP_423J2_125_3477_n1389), .B(
        DP_OP_423J2_125_3477_n1387), .CI(DP_OP_423J2_125_3477_n1403), .CO(
        DP_OP_423J2_125_3477_n1320), .S(DP_OP_423J2_125_3477_n1321) );
  FADDX1_HVT DP_OP_423J2_125_3477_U753 ( .A(DP_OP_423J2_125_3477_n1395), .B(
        DP_OP_423J2_125_3477_n1401), .CI(DP_OP_423J2_125_3477_n1399), .CO(
        DP_OP_423J2_125_3477_n1318), .S(DP_OP_423J2_125_3477_n1319) );
  FADDX1_HVT DP_OP_423J2_125_3477_U752 ( .A(DP_OP_423J2_125_3477_n1375), .B(
        DP_OP_423J2_125_3477_n1371), .CI(DP_OP_423J2_125_3477_n1355), .CO(
        DP_OP_423J2_125_3477_n1316), .S(DP_OP_423J2_125_3477_n1317) );
  FADDX1_HVT DP_OP_423J2_125_3477_U751 ( .A(DP_OP_423J2_125_3477_n1381), .B(
        DP_OP_423J2_125_3477_n1373), .CI(DP_OP_423J2_125_3477_n1357), .CO(
        DP_OP_423J2_125_3477_n1314), .S(DP_OP_423J2_125_3477_n1315) );
  FADDX1_HVT DP_OP_423J2_125_3477_U750 ( .A(DP_OP_423J2_125_3477_n1377), .B(
        DP_OP_423J2_125_3477_n1379), .CI(DP_OP_423J2_125_3477_n1359), .CO(
        DP_OP_423J2_125_3477_n1312), .S(DP_OP_423J2_125_3477_n1313) );
  FADDX1_HVT DP_OP_423J2_125_3477_U749 ( .A(DP_OP_423J2_125_3477_n1369), .B(
        DP_OP_423J2_125_3477_n1363), .CI(DP_OP_423J2_125_3477_n1361), .CO(
        DP_OP_423J2_125_3477_n1310), .S(DP_OP_423J2_125_3477_n1311) );
  FADDX1_HVT DP_OP_423J2_125_3477_U748 ( .A(DP_OP_423J2_125_3477_n1367), .B(
        DP_OP_423J2_125_3477_n1365), .CI(DP_OP_423J2_125_3477_n1504), .CO(
        DP_OP_423J2_125_3477_n1308), .S(DP_OP_423J2_125_3477_n1309) );
  FADDX1_HVT DP_OP_423J2_125_3477_U747 ( .A(DP_OP_423J2_125_3477_n1502), .B(
        DP_OP_423J2_125_3477_n1500), .CI(DP_OP_423J2_125_3477_n1498), .CO(
        DP_OP_423J2_125_3477_n1306), .S(DP_OP_423J2_125_3477_n1307) );
  FADDX1_HVT DP_OP_423J2_125_3477_U746 ( .A(DP_OP_423J2_125_3477_n1496), .B(
        DP_OP_423J2_125_3477_n1492), .CI(DP_OP_423J2_125_3477_n1349), .CO(
        DP_OP_423J2_125_3477_n1304), .S(DP_OP_423J2_125_3477_n1305) );
  FADDX1_HVT DP_OP_423J2_125_3477_U745 ( .A(DP_OP_423J2_125_3477_n1494), .B(
        DP_OP_423J2_125_3477_n1490), .CI(DP_OP_423J2_125_3477_n1351), .CO(
        DP_OP_423J2_125_3477_n1302), .S(DP_OP_423J2_125_3477_n1303) );
  FADDX1_HVT DP_OP_423J2_125_3477_U744 ( .A(DP_OP_423J2_125_3477_n1353), .B(
        DP_OP_423J2_125_3477_n1484), .CI(DP_OP_423J2_125_3477_n1486), .CO(
        DP_OP_423J2_125_3477_n1300), .S(DP_OP_423J2_125_3477_n1301) );
  FADDX1_HVT DP_OP_423J2_125_3477_U743 ( .A(DP_OP_423J2_125_3477_n1488), .B(
        DP_OP_423J2_125_3477_n1482), .CI(DP_OP_423J2_125_3477_n1480), .CO(
        DP_OP_423J2_125_3477_n1298), .S(DP_OP_423J2_125_3477_n1299) );
  FADDX1_HVT DP_OP_423J2_125_3477_U742 ( .A(DP_OP_423J2_125_3477_n1478), .B(
        DP_OP_423J2_125_3477_n1347), .CI(DP_OP_423J2_125_3477_n1341), .CO(
        DP_OP_423J2_125_3477_n1296), .S(DP_OP_423J2_125_3477_n1297) );
  FADDX1_HVT DP_OP_423J2_125_3477_U741 ( .A(DP_OP_423J2_125_3477_n1476), .B(
        DP_OP_423J2_125_3477_n1345), .CI(DP_OP_423J2_125_3477_n1343), .CO(
        DP_OP_423J2_125_3477_n1294), .S(DP_OP_423J2_125_3477_n1295) );
  FADDX1_HVT DP_OP_423J2_125_3477_U740 ( .A(DP_OP_423J2_125_3477_n1474), .B(
        DP_OP_423J2_125_3477_n1335), .CI(DP_OP_423J2_125_3477_n1468), .CO(
        DP_OP_423J2_125_3477_n1292), .S(DP_OP_423J2_125_3477_n1293) );
  FADDX1_HVT DP_OP_423J2_125_3477_U739 ( .A(DP_OP_423J2_125_3477_n1472), .B(
        DP_OP_423J2_125_3477_n1339), .CI(DP_OP_423J2_125_3477_n1327), .CO(
        DP_OP_423J2_125_3477_n1290), .S(DP_OP_423J2_125_3477_n1291) );
  FADDX1_HVT DP_OP_423J2_125_3477_U738 ( .A(DP_OP_423J2_125_3477_n1470), .B(
        DP_OP_423J2_125_3477_n1337), .CI(DP_OP_423J2_125_3477_n1333), .CO(
        DP_OP_423J2_125_3477_n1288), .S(DP_OP_423J2_125_3477_n1289) );
  FADDX1_HVT DP_OP_423J2_125_3477_U737 ( .A(DP_OP_423J2_125_3477_n1329), .B(
        DP_OP_423J2_125_3477_n1331), .CI(DP_OP_423J2_125_3477_n1466), .CO(
        DP_OP_423J2_125_3477_n1286), .S(DP_OP_423J2_125_3477_n1287) );
  FADDX1_HVT DP_OP_423J2_125_3477_U736 ( .A(DP_OP_423J2_125_3477_n1325), .B(
        DP_OP_423J2_125_3477_n1323), .CI(DP_OP_423J2_125_3477_n1321), .CO(
        DP_OP_423J2_125_3477_n1284), .S(DP_OP_423J2_125_3477_n1285) );
  FADDX1_HVT DP_OP_423J2_125_3477_U735 ( .A(DP_OP_423J2_125_3477_n1319), .B(
        DP_OP_423J2_125_3477_n1313), .CI(DP_OP_423J2_125_3477_n1315), .CO(
        DP_OP_423J2_125_3477_n1282), .S(DP_OP_423J2_125_3477_n1283) );
  FADDX1_HVT DP_OP_423J2_125_3477_U734 ( .A(DP_OP_423J2_125_3477_n1317), .B(
        DP_OP_423J2_125_3477_n1464), .CI(DP_OP_423J2_125_3477_n1311), .CO(
        DP_OP_423J2_125_3477_n1280), .S(DP_OP_423J2_125_3477_n1281) );
  FADDX1_HVT DP_OP_423J2_125_3477_U733 ( .A(DP_OP_423J2_125_3477_n1462), .B(
        DP_OP_423J2_125_3477_n1309), .CI(DP_OP_423J2_125_3477_n1460), .CO(
        DP_OP_423J2_125_3477_n1278), .S(DP_OP_423J2_125_3477_n1279) );
  FADDX1_HVT DP_OP_423J2_125_3477_U732 ( .A(DP_OP_423J2_125_3477_n1458), .B(
        DP_OP_423J2_125_3477_n1307), .CI(DP_OP_423J2_125_3477_n1456), .CO(
        DP_OP_423J2_125_3477_n1276), .S(DP_OP_423J2_125_3477_n1277) );
  FADDX1_HVT DP_OP_423J2_125_3477_U731 ( .A(DP_OP_423J2_125_3477_n1305), .B(
        DP_OP_423J2_125_3477_n1452), .CI(DP_OP_423J2_125_3477_n1301), .CO(
        DP_OP_423J2_125_3477_n1274), .S(DP_OP_423J2_125_3477_n1275) );
  FADDX1_HVT DP_OP_423J2_125_3477_U730 ( .A(DP_OP_423J2_125_3477_n1454), .B(
        DP_OP_423J2_125_3477_n1303), .CI(DP_OP_423J2_125_3477_n1450), .CO(
        DP_OP_423J2_125_3477_n1272), .S(DP_OP_423J2_125_3477_n1273) );
  FADDX1_HVT DP_OP_423J2_125_3477_U729 ( .A(DP_OP_423J2_125_3477_n1299), .B(
        DP_OP_423J2_125_3477_n1297), .CI(DP_OP_423J2_125_3477_n1448), .CO(
        DP_OP_423J2_125_3477_n1270), .S(DP_OP_423J2_125_3477_n1271) );
  FADDX1_HVT DP_OP_423J2_125_3477_U728 ( .A(DP_OP_423J2_125_3477_n1295), .B(
        DP_OP_423J2_125_3477_n1446), .CI(DP_OP_423J2_125_3477_n1444), .CO(
        DP_OP_423J2_125_3477_n1268), .S(DP_OP_423J2_125_3477_n1269) );
  FADDX1_HVT DP_OP_423J2_125_3477_U727 ( .A(DP_OP_423J2_125_3477_n1291), .B(
        DP_OP_423J2_125_3477_n1289), .CI(DP_OP_423J2_125_3477_n1287), .CO(
        DP_OP_423J2_125_3477_n1266), .S(DP_OP_423J2_125_3477_n1267) );
  FADDX1_HVT DP_OP_423J2_125_3477_U726 ( .A(DP_OP_423J2_125_3477_n1293), .B(
        DP_OP_423J2_125_3477_n1285), .CI(DP_OP_423J2_125_3477_n1442), .CO(
        DP_OP_423J2_125_3477_n1264), .S(DP_OP_423J2_125_3477_n1265) );
  FADDX1_HVT DP_OP_423J2_125_3477_U725 ( .A(DP_OP_423J2_125_3477_n1283), .B(
        DP_OP_423J2_125_3477_n1281), .CI(DP_OP_423J2_125_3477_n1440), .CO(
        DP_OP_423J2_125_3477_n1262), .S(DP_OP_423J2_125_3477_n1263) );
  FADDX1_HVT DP_OP_423J2_125_3477_U724 ( .A(DP_OP_423J2_125_3477_n1279), .B(
        DP_OP_423J2_125_3477_n1438), .CI(DP_OP_423J2_125_3477_n1277), .CO(
        DP_OP_423J2_125_3477_n1260), .S(DP_OP_423J2_125_3477_n1261) );
  FADDX1_HVT DP_OP_423J2_125_3477_U723 ( .A(DP_OP_423J2_125_3477_n1436), .B(
        DP_OP_423J2_125_3477_n1275), .CI(DP_OP_423J2_125_3477_n1434), .CO(
        DP_OP_423J2_125_3477_n1258), .S(DP_OP_423J2_125_3477_n1259) );
  FADDX1_HVT DP_OP_423J2_125_3477_U722 ( .A(DP_OP_423J2_125_3477_n1273), .B(
        DP_OP_423J2_125_3477_n1432), .CI(DP_OP_423J2_125_3477_n1271), .CO(
        DP_OP_423J2_125_3477_n1256), .S(DP_OP_423J2_125_3477_n1257) );
  FADDX1_HVT DP_OP_423J2_125_3477_U721 ( .A(DP_OP_423J2_125_3477_n1269), .B(
        DP_OP_423J2_125_3477_n1267), .CI(DP_OP_423J2_125_3477_n1430), .CO(
        DP_OP_423J2_125_3477_n1254), .S(DP_OP_423J2_125_3477_n1255) );
  FADDX1_HVT DP_OP_423J2_125_3477_U720 ( .A(DP_OP_423J2_125_3477_n1265), .B(
        DP_OP_423J2_125_3477_n1263), .CI(DP_OP_423J2_125_3477_n1428), .CO(
        DP_OP_423J2_125_3477_n1252), .S(DP_OP_423J2_125_3477_n1253) );
  FADDX1_HVT DP_OP_423J2_125_3477_U719 ( .A(DP_OP_423J2_125_3477_n1261), .B(
        DP_OP_423J2_125_3477_n1426), .CI(DP_OP_423J2_125_3477_n1259), .CO(
        DP_OP_423J2_125_3477_n1250), .S(DP_OP_423J2_125_3477_n1251) );
  FADDX1_HVT DP_OP_423J2_125_3477_U718 ( .A(DP_OP_423J2_125_3477_n1257), .B(
        DP_OP_423J2_125_3477_n1424), .CI(DP_OP_423J2_125_3477_n1255), .CO(
        DP_OP_423J2_125_3477_n1248), .S(DP_OP_423J2_125_3477_n1249) );
  FADDX1_HVT DP_OP_423J2_125_3477_U717 ( .A(DP_OP_423J2_125_3477_n1253), .B(
        DP_OP_423J2_125_3477_n1422), .CI(DP_OP_423J2_125_3477_n1251), .CO(
        DP_OP_423J2_125_3477_n1246), .S(DP_OP_423J2_125_3477_n1247) );
  HADDX1_HVT DP_OP_423J2_125_3477_U716 ( .A0(DP_OP_423J2_125_3477_n2700), .B0(
        DP_OP_423J2_125_3477_n2042), .C1(DP_OP_423J2_125_3477_n1244), .SO(
        DP_OP_423J2_125_3477_n1245) );
  FADDX1_HVT DP_OP_423J2_125_3477_U715 ( .A(DP_OP_423J2_125_3477_n1998), .B(
        DP_OP_423J2_125_3477_n2482), .CI(DP_OP_423J2_125_3477_n1954), .CO(
        DP_OP_423J2_125_3477_n1242), .S(DP_OP_423J2_125_3477_n1243) );
  FADDX1_HVT DP_OP_423J2_125_3477_U714 ( .A(DP_OP_423J2_125_3477_n2130), .B(
        DP_OP_423J2_125_3477_n2438), .CI(DP_OP_423J2_125_3477_n2743), .CO(
        DP_OP_423J2_125_3477_n1240), .S(DP_OP_423J2_125_3477_n1241) );
  FADDX1_HVT DP_OP_423J2_125_3477_U713 ( .A(DP_OP_423J2_125_3477_n2306), .B(
        DP_OP_423J2_125_3477_n1910), .CI(DP_OP_423J2_125_3477_n2174), .CO(
        DP_OP_423J2_125_3477_n1238), .S(DP_OP_423J2_125_3477_n1239) );
  FADDX1_HVT DP_OP_423J2_125_3477_U712 ( .A(DP_OP_423J2_125_3477_n2658), .B(
        DP_OP_423J2_125_3477_n2526), .CI(DP_OP_423J2_125_3477_n2570), .CO(
        DP_OP_423J2_125_3477_n1236), .S(DP_OP_423J2_125_3477_n1237) );
  FADDX1_HVT DP_OP_423J2_125_3477_U711 ( .A(DP_OP_423J2_125_3477_n2787), .B(
        DP_OP_423J2_125_3477_n1822), .CI(DP_OP_423J2_125_3477_n2875), .CO(
        DP_OP_423J2_125_3477_n1234), .S(DP_OP_423J2_125_3477_n1235) );
  FADDX1_HVT DP_OP_423J2_125_3477_U710 ( .A(DP_OP_423J2_125_3477_n1866), .B(
        DP_OP_423J2_125_3477_n2614), .CI(DP_OP_423J2_125_3477_n2262), .CO(
        DP_OP_423J2_125_3477_n1232), .S(DP_OP_423J2_125_3477_n1233) );
  FADDX1_HVT DP_OP_423J2_125_3477_U709 ( .A(DP_OP_423J2_125_3477_n2831), .B(
        DP_OP_423J2_125_3477_n2086), .CI(DP_OP_423J2_125_3477_n2350), .CO(
        DP_OP_423J2_125_3477_n1230), .S(DP_OP_423J2_125_3477_n1231) );
  FADDX1_HVT DP_OP_423J2_125_3477_U708 ( .A(DP_OP_423J2_125_3477_n1778), .B(
        DP_OP_423J2_125_3477_n2394), .CI(DP_OP_423J2_125_3477_n2764), .CO(
        DP_OP_423J2_125_3477_n1228), .S(DP_OP_423J2_125_3477_n1229) );
  FADDX1_HVT DP_OP_423J2_125_3477_U707 ( .A(DP_OP_423J2_125_3477_n1843), .B(
        DP_OP_423J2_125_3477_n1961), .CI(DP_OP_423J2_125_3477_n2225), .CO(
        DP_OP_423J2_125_3477_n1226), .S(DP_OP_423J2_125_3477_n1227) );
  FADDX1_HVT DP_OP_423J2_125_3477_U706 ( .A(DP_OP_423J2_125_3477_n2635), .B(
        DP_OP_423J2_125_3477_n2720), .CI(DP_OP_423J2_125_3477_n2093), .CO(
        DP_OP_423J2_125_3477_n1224), .S(DP_OP_423J2_125_3477_n1225) );
  FADDX1_HVT DP_OP_423J2_125_3477_U705 ( .A(DP_OP_423J2_125_3477_n2107), .B(
        DP_OP_423J2_125_3477_n2408), .CI(DP_OP_423J2_125_3477_n2852), .CO(
        DP_OP_423J2_125_3477_n1222), .S(DP_OP_423J2_125_3477_n1223) );
  FADDX1_HVT DP_OP_423J2_125_3477_U704 ( .A(DP_OP_423J2_125_3477_n2195), .B(
        DP_OP_423J2_125_3477_n2533), .CI(DP_OP_423J2_125_3477_n1887), .CO(
        DP_OP_423J2_125_3477_n1220), .S(DP_OP_423J2_125_3477_n1221) );
  FADDX1_HVT DP_OP_423J2_125_3477_U703 ( .A(DP_OP_423J2_125_3477_n2882), .B(
        DP_OP_423J2_125_3477_n2144), .CI(DP_OP_423J2_125_3477_n2445), .CO(
        DP_OP_423J2_125_3477_n1218), .S(DP_OP_423J2_125_3477_n1219) );
  FADDX1_HVT DP_OP_423J2_125_3477_U702 ( .A(DP_OP_423J2_125_3477_n2591), .B(
        DP_OP_423J2_125_3477_n2218), .CI(DP_OP_423J2_125_3477_n2503), .CO(
        DP_OP_423J2_125_3477_n1216), .S(DP_OP_423J2_125_3477_n1217) );
  FADDX1_HVT DP_OP_423J2_125_3477_U701 ( .A(DP_OP_423J2_125_3477_n2547), .B(
        DP_OP_423J2_125_3477_n2320), .CI(DP_OP_423J2_125_3477_n2496), .CO(
        DP_OP_423J2_125_3477_n1214), .S(DP_OP_423J2_125_3477_n1215) );
  FADDX1_HVT DP_OP_423J2_125_3477_U700 ( .A(DP_OP_423J2_125_3477_n2838), .B(
        DP_OP_423J2_125_3477_n2056), .CI(DP_OP_423J2_125_3477_n2628), .CO(
        DP_OP_423J2_125_3477_n1212), .S(DP_OP_423J2_125_3477_n1213) );
  FADDX1_HVT DP_OP_423J2_125_3477_U699 ( .A(DP_OP_423J2_125_3477_n2415), .B(
        DP_OP_423J2_125_3477_n2679), .CI(DP_OP_423J2_125_3477_n1836), .CO(
        DP_OP_423J2_125_3477_n1210), .S(DP_OP_423J2_125_3477_n1211) );
  FADDX1_HVT DP_OP_423J2_125_3477_U698 ( .A(DP_OP_423J2_125_3477_n2459), .B(
        DP_OP_423J2_125_3477_n2019), .CI(DP_OP_423J2_125_3477_n2584), .CO(
        DP_OP_423J2_125_3477_n1208), .S(DP_OP_423J2_125_3477_n1209) );
  FADDX1_HVT DP_OP_423J2_125_3477_U697 ( .A(DP_OP_423J2_125_3477_n2327), .B(
        DP_OP_423J2_125_3477_n1975), .CI(DP_OP_423J2_125_3477_n2750), .CO(
        DP_OP_423J2_125_3477_n1206), .S(DP_OP_423J2_125_3477_n1207) );
  FADDX1_HVT DP_OP_423J2_125_3477_U696 ( .A(DP_OP_423J2_125_3477_n2269), .B(
        DP_OP_423J2_125_3477_n2357), .CI(DP_OP_423J2_125_3477_n2889), .CO(
        DP_OP_423J2_125_3477_n1204), .S(DP_OP_423J2_125_3477_n1205) );
  FADDX1_HVT DP_OP_423J2_125_3477_U695 ( .A(DP_OP_423J2_125_3477_n2283), .B(
        DP_OP_423J2_125_3477_n2239), .CI(DP_OP_423J2_125_3477_n2801), .CO(
        DP_OP_423J2_125_3477_n1202), .S(DP_OP_423J2_125_3477_n1203) );
  FADDX1_HVT DP_OP_423J2_125_3477_U694 ( .A(DP_OP_423J2_125_3477_n2063), .B(
        DP_OP_423J2_125_3477_n1880), .CI(DP_OP_423J2_125_3477_n2276), .CO(
        DP_OP_423J2_125_3477_n1200), .S(DP_OP_423J2_125_3477_n1201) );
  FADDX1_HVT DP_OP_423J2_125_3477_U693 ( .A(DP_OP_423J2_125_3477_n2137), .B(
        DP_OP_423J2_125_3477_n2100), .CI(DP_OP_423J2_125_3477_n1924), .CO(
        DP_OP_423J2_125_3477_n1198), .S(DP_OP_423J2_125_3477_n1199) );
  FADDX1_HVT DP_OP_423J2_125_3477_U692 ( .A(DP_OP_423J2_125_3477_n2577), .B(
        DP_OP_423J2_125_3477_n2452), .CI(DP_OP_423J2_125_3477_n2896), .CO(
        DP_OP_423J2_125_3477_n1196), .S(DP_OP_423J2_125_3477_n1197) );
  FADDX1_HVT DP_OP_423J2_125_3477_U691 ( .A(DP_OP_423J2_125_3477_n2672), .B(
        DP_OP_423J2_125_3477_n2489), .CI(DP_OP_423J2_125_3477_n2757), .CO(
        DP_OP_423J2_125_3477_n1194), .S(DP_OP_423J2_125_3477_n1195) );
  FADDX1_HVT DP_OP_423J2_125_3477_U690 ( .A(DP_OP_423J2_125_3477_n2665), .B(
        DP_OP_423J2_125_3477_n2401), .CI(DP_OP_423J2_125_3477_n2808), .CO(
        DP_OP_423J2_125_3477_n1192), .S(DP_OP_423J2_125_3477_n1193) );
  FADDX1_HVT DP_OP_423J2_125_3477_U689 ( .A(DP_OP_423J2_125_3477_n2706), .B(
        DP_OP_423J2_125_3477_n2713), .CI(DP_OP_423J2_125_3477_n1829), .CO(
        DP_OP_423J2_125_3477_n1190), .S(DP_OP_423J2_125_3477_n1191) );
  FADDX1_HVT DP_OP_423J2_125_3477_U688 ( .A(DP_OP_423J2_125_3477_n2540), .B(
        DP_OP_423J2_125_3477_n2371), .CI(DP_OP_423J2_125_3477_n2181), .CO(
        DP_OP_423J2_125_3477_n1188), .S(DP_OP_423J2_125_3477_n1189) );
  FADDX1_HVT DP_OP_423J2_125_3477_U687 ( .A(DP_OP_423J2_125_3477_n2049), .B(
        DP_OP_423J2_125_3477_n2232), .CI(DP_OP_423J2_125_3477_n1917), .CO(
        DP_OP_423J2_125_3477_n1186), .S(DP_OP_423J2_125_3477_n1187) );
  FADDX1_HVT DP_OP_423J2_125_3477_U686 ( .A(DP_OP_423J2_125_3477_n2313), .B(
        DP_OP_423J2_125_3477_n2364), .CI(DP_OP_423J2_125_3477_n1968), .CO(
        DP_OP_423J2_125_3477_n1184), .S(DP_OP_423J2_125_3477_n1185) );
  FADDX1_HVT DP_OP_423J2_125_3477_U685 ( .A(DP_OP_423J2_125_3477_n1931), .B(
        DP_OP_423J2_125_3477_n2188), .CI(DP_OP_423J2_125_3477_n2794), .CO(
        DP_OP_423J2_125_3477_n1182), .S(DP_OP_423J2_125_3477_n1183) );
  FADDX1_HVT DP_OP_423J2_125_3477_U684 ( .A(DP_OP_423J2_125_3477_n2845), .B(
        DP_OP_423J2_125_3477_n2005), .CI(DP_OP_423J2_125_3477_n2621), .CO(
        DP_OP_423J2_125_3477_n1180), .S(DP_OP_423J2_125_3477_n1181) );
  FADDX1_HVT DP_OP_423J2_125_3477_U683 ( .A(DP_OP_423J2_125_3477_n2151), .B(
        DP_OP_423J2_125_3477_n2012), .CI(DP_OP_423J2_125_3477_n1873), .CO(
        DP_OP_423J2_125_3477_n1178), .S(DP_OP_423J2_125_3477_n1179) );
  FADDX1_HVT DP_OP_423J2_125_3477_U682 ( .A(DP_OP_423J2_125_3477_n1245), .B(
        DP_OP_423J2_125_3477_n1420), .CI(DP_OP_423J2_125_3477_n1406), .CO(
        DP_OP_423J2_125_3477_n1176), .S(DP_OP_423J2_125_3477_n1177) );
  FADDX1_HVT DP_OP_423J2_125_3477_U681 ( .A(DP_OP_423J2_125_3477_n1418), .B(
        DP_OP_423J2_125_3477_n1414), .CI(DP_OP_423J2_125_3477_n1408), .CO(
        DP_OP_423J2_125_3477_n1174), .S(DP_OP_423J2_125_3477_n1175) );
  FADDX1_HVT DP_OP_423J2_125_3477_U680 ( .A(DP_OP_423J2_125_3477_n1416), .B(
        DP_OP_423J2_125_3477_n1412), .CI(DP_OP_423J2_125_3477_n1410), .CO(
        DP_OP_423J2_125_3477_n1172), .S(DP_OP_423J2_125_3477_n1173) );
  FADDX1_HVT DP_OP_423J2_125_3477_U679 ( .A(DP_OP_423J2_125_3477_n1404), .B(
        DP_OP_423J2_125_3477_n1382), .CI(DP_OP_423J2_125_3477_n1384), .CO(
        DP_OP_423J2_125_3477_n1170), .S(DP_OP_423J2_125_3477_n1171) );
  FADDX1_HVT DP_OP_423J2_125_3477_U678 ( .A(DP_OP_423J2_125_3477_n1402), .B(
        DP_OP_423J2_125_3477_n1386), .CI(DP_OP_423J2_125_3477_n1388), .CO(
        DP_OP_423J2_125_3477_n1168), .S(DP_OP_423J2_125_3477_n1169) );
  FADDX1_HVT DP_OP_423J2_125_3477_U677 ( .A(DP_OP_423J2_125_3477_n1400), .B(
        DP_OP_423J2_125_3477_n1390), .CI(DP_OP_423J2_125_3477_n1392), .CO(
        DP_OP_423J2_125_3477_n1166), .S(DP_OP_423J2_125_3477_n1167) );
  FADDX1_HVT DP_OP_423J2_125_3477_U676 ( .A(DP_OP_423J2_125_3477_n1398), .B(
        DP_OP_423J2_125_3477_n1394), .CI(DP_OP_423J2_125_3477_n1396), .CO(
        DP_OP_423J2_125_3477_n1164), .S(DP_OP_423J2_125_3477_n1165) );
  FADDX1_HVT DP_OP_423J2_125_3477_U675 ( .A(DP_OP_423J2_125_3477_n1380), .B(
        DP_OP_423J2_125_3477_n1370), .CI(DP_OP_423J2_125_3477_n1354), .CO(
        DP_OP_423J2_125_3477_n1162), .S(DP_OP_423J2_125_3477_n1163) );
  FADDX1_HVT DP_OP_423J2_125_3477_U674 ( .A(DP_OP_423J2_125_3477_n1378), .B(
        DP_OP_423J2_125_3477_n1372), .CI(DP_OP_423J2_125_3477_n1356), .CO(
        DP_OP_423J2_125_3477_n1160), .S(DP_OP_423J2_125_3477_n1161) );
  FADDX1_HVT DP_OP_423J2_125_3477_U673 ( .A(DP_OP_423J2_125_3477_n1376), .B(
        DP_OP_423J2_125_3477_n1374), .CI(DP_OP_423J2_125_3477_n1358), .CO(
        DP_OP_423J2_125_3477_n1158), .S(DP_OP_423J2_125_3477_n1159) );
  FADDX1_HVT DP_OP_423J2_125_3477_U672 ( .A(DP_OP_423J2_125_3477_n1243), .B(
        DP_OP_423J2_125_3477_n1360), .CI(DP_OP_423J2_125_3477_n1362), .CO(
        DP_OP_423J2_125_3477_n1156), .S(DP_OP_423J2_125_3477_n1157) );
  FADDX1_HVT DP_OP_423J2_125_3477_U671 ( .A(DP_OP_423J2_125_3477_n1233), .B(
        DP_OP_423J2_125_3477_n1364), .CI(DP_OP_423J2_125_3477_n1366), .CO(
        DP_OP_423J2_125_3477_n1154), .S(DP_OP_423J2_125_3477_n1155) );
  FADDX1_HVT DP_OP_423J2_125_3477_U670 ( .A(DP_OP_423J2_125_3477_n1235), .B(
        DP_OP_423J2_125_3477_n1241), .CI(DP_OP_423J2_125_3477_n1368), .CO(
        DP_OP_423J2_125_3477_n1152), .S(DP_OP_423J2_125_3477_n1153) );
  FADDX1_HVT DP_OP_423J2_125_3477_U669 ( .A(DP_OP_423J2_125_3477_n1237), .B(
        DP_OP_423J2_125_3477_n1231), .CI(DP_OP_423J2_125_3477_n1239), .CO(
        DP_OP_423J2_125_3477_n1150), .S(DP_OP_423J2_125_3477_n1151) );
  FADDX1_HVT DP_OP_423J2_125_3477_U668 ( .A(DP_OP_423J2_125_3477_n1229), .B(
        DP_OP_423J2_125_3477_n1209), .CI(DP_OP_423J2_125_3477_n1207), .CO(
        DP_OP_423J2_125_3477_n1148), .S(DP_OP_423J2_125_3477_n1149) );
  FADDX1_HVT DP_OP_423J2_125_3477_U667 ( .A(DP_OP_423J2_125_3477_n1221), .B(
        DP_OP_423J2_125_3477_n1211), .CI(DP_OP_423J2_125_3477_n1217), .CO(
        DP_OP_423J2_125_3477_n1146), .S(DP_OP_423J2_125_3477_n1147) );
  FADDX1_HVT DP_OP_423J2_125_3477_U666 ( .A(DP_OP_423J2_125_3477_n1219), .B(
        DP_OP_423J2_125_3477_n1227), .CI(DP_OP_423J2_125_3477_n1225), .CO(
        DP_OP_423J2_125_3477_n1144), .S(DP_OP_423J2_125_3477_n1145) );
  FADDX1_HVT DP_OP_423J2_125_3477_U665 ( .A(DP_OP_423J2_125_3477_n1215), .B(
        DP_OP_423J2_125_3477_n1223), .CI(DP_OP_423J2_125_3477_n1213), .CO(
        DP_OP_423J2_125_3477_n1142), .S(DP_OP_423J2_125_3477_n1143) );
  FADDX1_HVT DP_OP_423J2_125_3477_U664 ( .A(DP_OP_423J2_125_3477_n1203), .B(
        DP_OP_423J2_125_3477_n1195), .CI(DP_OP_423J2_125_3477_n1179), .CO(
        DP_OP_423J2_125_3477_n1140), .S(DP_OP_423J2_125_3477_n1141) );
  FADDX1_HVT DP_OP_423J2_125_3477_U663 ( .A(DP_OP_423J2_125_3477_n1205), .B(
        DP_OP_423J2_125_3477_n1197), .CI(DP_OP_423J2_125_3477_n1181), .CO(
        DP_OP_423J2_125_3477_n1138), .S(DP_OP_423J2_125_3477_n1139) );
  FADDX1_HVT DP_OP_423J2_125_3477_U662 ( .A(DP_OP_423J2_125_3477_n1201), .B(
        DP_OP_423J2_125_3477_n1199), .CI(DP_OP_423J2_125_3477_n1183), .CO(
        DP_OP_423J2_125_3477_n1136), .S(DP_OP_423J2_125_3477_n1137) );
  FADDX1_HVT DP_OP_423J2_125_3477_U661 ( .A(DP_OP_423J2_125_3477_n1193), .B(
        DP_OP_423J2_125_3477_n1185), .CI(DP_OP_423J2_125_3477_n1352), .CO(
        DP_OP_423J2_125_3477_n1134), .S(DP_OP_423J2_125_3477_n1135) );
  FADDX1_HVT DP_OP_423J2_125_3477_U660 ( .A(DP_OP_423J2_125_3477_n1191), .B(
        DP_OP_423J2_125_3477_n1187), .CI(DP_OP_423J2_125_3477_n1350), .CO(
        DP_OP_423J2_125_3477_n1132), .S(DP_OP_423J2_125_3477_n1133) );
  FADDX1_HVT DP_OP_423J2_125_3477_U659 ( .A(DP_OP_423J2_125_3477_n1189), .B(
        DP_OP_423J2_125_3477_n1348), .CI(DP_OP_423J2_125_3477_n1346), .CO(
        DP_OP_423J2_125_3477_n1130), .S(DP_OP_423J2_125_3477_n1131) );
  FADDX1_HVT DP_OP_423J2_125_3477_U658 ( .A(DP_OP_423J2_125_3477_n1344), .B(
        DP_OP_423J2_125_3477_n1340), .CI(DP_OP_423J2_125_3477_n1342), .CO(
        DP_OP_423J2_125_3477_n1128), .S(DP_OP_423J2_125_3477_n1129) );
  FADDX1_HVT DP_OP_423J2_125_3477_U657 ( .A(DP_OP_423J2_125_3477_n1336), .B(
        DP_OP_423J2_125_3477_n1334), .CI(DP_OP_423J2_125_3477_n1326), .CO(
        DP_OP_423J2_125_3477_n1126), .S(DP_OP_423J2_125_3477_n1127) );
  FADDX1_HVT DP_OP_423J2_125_3477_U656 ( .A(DP_OP_423J2_125_3477_n1338), .B(
        DP_OP_423J2_125_3477_n1177), .CI(DP_OP_423J2_125_3477_n1175), .CO(
        DP_OP_423J2_125_3477_n1124), .S(DP_OP_423J2_125_3477_n1125) );
  FADDX1_HVT DP_OP_423J2_125_3477_U655 ( .A(DP_OP_423J2_125_3477_n1173), .B(
        DP_OP_423J2_125_3477_n1328), .CI(DP_OP_423J2_125_3477_n1330), .CO(
        DP_OP_423J2_125_3477_n1122), .S(DP_OP_423J2_125_3477_n1123) );
  FADDX1_HVT DP_OP_423J2_125_3477_U654 ( .A(DP_OP_423J2_125_3477_n1332), .B(
        DP_OP_423J2_125_3477_n1324), .CI(DP_OP_423J2_125_3477_n1171), .CO(
        DP_OP_423J2_125_3477_n1120), .S(DP_OP_423J2_125_3477_n1121) );
  FADDX1_HVT DP_OP_423J2_125_3477_U653 ( .A(DP_OP_423J2_125_3477_n1165), .B(
        DP_OP_423J2_125_3477_n1167), .CI(DP_OP_423J2_125_3477_n1169), .CO(
        DP_OP_423J2_125_3477_n1118), .S(DP_OP_423J2_125_3477_n1119) );
  FADDX1_HVT DP_OP_423J2_125_3477_U652 ( .A(DP_OP_423J2_125_3477_n1322), .B(
        DP_OP_423J2_125_3477_n1318), .CI(DP_OP_423J2_125_3477_n1320), .CO(
        DP_OP_423J2_125_3477_n1116), .S(DP_OP_423J2_125_3477_n1117) );
  FADDX1_HVT DP_OP_423J2_125_3477_U651 ( .A(DP_OP_423J2_125_3477_n1316), .B(
        DP_OP_423J2_125_3477_n1159), .CI(DP_OP_423J2_125_3477_n1310), .CO(
        DP_OP_423J2_125_3477_n1114), .S(DP_OP_423J2_125_3477_n1115) );
  FADDX1_HVT DP_OP_423J2_125_3477_U650 ( .A(DP_OP_423J2_125_3477_n1314), .B(
        DP_OP_423J2_125_3477_n1163), .CI(DP_OP_423J2_125_3477_n1153), .CO(
        DP_OP_423J2_125_3477_n1112), .S(DP_OP_423J2_125_3477_n1113) );
  FADDX1_HVT DP_OP_423J2_125_3477_U649 ( .A(DP_OP_423J2_125_3477_n1312), .B(
        DP_OP_423J2_125_3477_n1161), .CI(DP_OP_423J2_125_3477_n1155), .CO(
        DP_OP_423J2_125_3477_n1110), .S(DP_OP_423J2_125_3477_n1111) );
  FADDX1_HVT DP_OP_423J2_125_3477_U648 ( .A(DP_OP_423J2_125_3477_n1157), .B(
        DP_OP_423J2_125_3477_n1151), .CI(DP_OP_423J2_125_3477_n1149), .CO(
        DP_OP_423J2_125_3477_n1108), .S(DP_OP_423J2_125_3477_n1109) );
  FADDX1_HVT DP_OP_423J2_125_3477_U647 ( .A(DP_OP_423J2_125_3477_n1143), .B(
        DP_OP_423J2_125_3477_n1147), .CI(DP_OP_423J2_125_3477_n1308), .CO(
        DP_OP_423J2_125_3477_n1106), .S(DP_OP_423J2_125_3477_n1107) );
  FADDX1_HVT DP_OP_423J2_125_3477_U646 ( .A(DP_OP_423J2_125_3477_n1145), .B(
        DP_OP_423J2_125_3477_n1137), .CI(DP_OP_423J2_125_3477_n1139), .CO(
        DP_OP_423J2_125_3477_n1104), .S(DP_OP_423J2_125_3477_n1105) );
  FADDX1_HVT DP_OP_423J2_125_3477_U645 ( .A(DP_OP_423J2_125_3477_n1141), .B(
        DP_OP_423J2_125_3477_n1306), .CI(DP_OP_423J2_125_3477_n1133), .CO(
        DP_OP_423J2_125_3477_n1102), .S(DP_OP_423J2_125_3477_n1103) );
  FADDX1_HVT DP_OP_423J2_125_3477_U644 ( .A(DP_OP_423J2_125_3477_n1135), .B(
        DP_OP_423J2_125_3477_n1304), .CI(DP_OP_423J2_125_3477_n1300), .CO(
        DP_OP_423J2_125_3477_n1100), .S(DP_OP_423J2_125_3477_n1101) );
  FADDX1_HVT DP_OP_423J2_125_3477_U643 ( .A(DP_OP_423J2_125_3477_n1302), .B(
        DP_OP_423J2_125_3477_n1131), .CI(DP_OP_423J2_125_3477_n1298), .CO(
        DP_OP_423J2_125_3477_n1098), .S(DP_OP_423J2_125_3477_n1099) );
  FADDX1_HVT DP_OP_423J2_125_3477_U642 ( .A(DP_OP_423J2_125_3477_n1296), .B(
        DP_OP_423J2_125_3477_n1294), .CI(DP_OP_423J2_125_3477_n1129), .CO(
        DP_OP_423J2_125_3477_n1096), .S(DP_OP_423J2_125_3477_n1097) );
  FADDX1_HVT DP_OP_423J2_125_3477_U641 ( .A(DP_OP_423J2_125_3477_n1292), .B(
        DP_OP_423J2_125_3477_n1127), .CI(DP_OP_423J2_125_3477_n1123), .CO(
        DP_OP_423J2_125_3477_n1094), .S(DP_OP_423J2_125_3477_n1095) );
  FADDX1_HVT DP_OP_423J2_125_3477_U640 ( .A(DP_OP_423J2_125_3477_n1290), .B(
        DP_OP_423J2_125_3477_n1125), .CI(DP_OP_423J2_125_3477_n1286), .CO(
        DP_OP_423J2_125_3477_n1092), .S(DP_OP_423J2_125_3477_n1093) );
  FADDX1_HVT DP_OP_423J2_125_3477_U639 ( .A(DP_OP_423J2_125_3477_n1288), .B(
        DP_OP_423J2_125_3477_n1121), .CI(DP_OP_423J2_125_3477_n1284), .CO(
        DP_OP_423J2_125_3477_n1090), .S(DP_OP_423J2_125_3477_n1091) );
  FADDX1_HVT DP_OP_423J2_125_3477_U638 ( .A(DP_OP_423J2_125_3477_n1117), .B(
        DP_OP_423J2_125_3477_n1119), .CI(DP_OP_423J2_125_3477_n1282), .CO(
        DP_OP_423J2_125_3477_n1088), .S(DP_OP_423J2_125_3477_n1089) );
  FADDX1_HVT DP_OP_423J2_125_3477_U637 ( .A(DP_OP_423J2_125_3477_n1280), .B(
        DP_OP_423J2_125_3477_n1111), .CI(DP_OP_423J2_125_3477_n1109), .CO(
        DP_OP_423J2_125_3477_n1086), .S(DP_OP_423J2_125_3477_n1087) );
  FADDX1_HVT DP_OP_423J2_125_3477_U636 ( .A(DP_OP_423J2_125_3477_n1115), .B(
        DP_OP_423J2_125_3477_n1113), .CI(DP_OP_423J2_125_3477_n1107), .CO(
        DP_OP_423J2_125_3477_n1084), .S(DP_OP_423J2_125_3477_n1085) );
  FADDX1_HVT DP_OP_423J2_125_3477_U635 ( .A(DP_OP_423J2_125_3477_n1278), .B(
        DP_OP_423J2_125_3477_n1105), .CI(DP_OP_423J2_125_3477_n1103), .CO(
        DP_OP_423J2_125_3477_n1082), .S(DP_OP_423J2_125_3477_n1083) );
  FADDX1_HVT DP_OP_423J2_125_3477_U634 ( .A(DP_OP_423J2_125_3477_n1276), .B(
        DP_OP_423J2_125_3477_n1101), .CI(DP_OP_423J2_125_3477_n1274), .CO(
        DP_OP_423J2_125_3477_n1080), .S(DP_OP_423J2_125_3477_n1081) );
  FADDX1_HVT DP_OP_423J2_125_3477_U633 ( .A(DP_OP_423J2_125_3477_n1272), .B(
        DP_OP_423J2_125_3477_n1099), .CI(DP_OP_423J2_125_3477_n1270), .CO(
        DP_OP_423J2_125_3477_n1078), .S(DP_OP_423J2_125_3477_n1079) );
  FADDX1_HVT DP_OP_423J2_125_3477_U632 ( .A(DP_OP_423J2_125_3477_n1268), .B(
        DP_OP_423J2_125_3477_n1097), .CI(DP_OP_423J2_125_3477_n1093), .CO(
        DP_OP_423J2_125_3477_n1076), .S(DP_OP_423J2_125_3477_n1077) );
  FADDX1_HVT DP_OP_423J2_125_3477_U631 ( .A(DP_OP_423J2_125_3477_n1095), .B(
        DP_OP_423J2_125_3477_n1266), .CI(DP_OP_423J2_125_3477_n1091), .CO(
        DP_OP_423J2_125_3477_n1074), .S(DP_OP_423J2_125_3477_n1075) );
  FADDX1_HVT DP_OP_423J2_125_3477_U630 ( .A(DP_OP_423J2_125_3477_n1264), .B(
        DP_OP_423J2_125_3477_n1089), .CI(DP_OP_423J2_125_3477_n1262), .CO(
        DP_OP_423J2_125_3477_n1072), .S(DP_OP_423J2_125_3477_n1073) );
  FADDX1_HVT DP_OP_423J2_125_3477_U629 ( .A(DP_OP_423J2_125_3477_n1087), .B(
        DP_OP_423J2_125_3477_n1085), .CI(DP_OP_423J2_125_3477_n1260), .CO(
        DP_OP_423J2_125_3477_n1070), .S(DP_OP_423J2_125_3477_n1071) );
  FADDX1_HVT DP_OP_423J2_125_3477_U628 ( .A(DP_OP_423J2_125_3477_n1083), .B(
        DP_OP_423J2_125_3477_n1081), .CI(DP_OP_423J2_125_3477_n1258), .CO(
        DP_OP_423J2_125_3477_n1068), .S(DP_OP_423J2_125_3477_n1069) );
  FADDX1_HVT DP_OP_423J2_125_3477_U627 ( .A(DP_OP_423J2_125_3477_n1079), .B(
        DP_OP_423J2_125_3477_n1256), .CI(DP_OP_423J2_125_3477_n1077), .CO(
        DP_OP_423J2_125_3477_n1066), .S(DP_OP_423J2_125_3477_n1067) );
  FADDX1_HVT DP_OP_423J2_125_3477_U626 ( .A(DP_OP_423J2_125_3477_n1254), .B(
        DP_OP_423J2_125_3477_n1075), .CI(DP_OP_423J2_125_3477_n1073), .CO(
        DP_OP_423J2_125_3477_n1064), .S(DP_OP_423J2_125_3477_n1065) );
  FADDX1_HVT DP_OP_423J2_125_3477_U625 ( .A(DP_OP_423J2_125_3477_n1252), .B(
        DP_OP_423J2_125_3477_n1071), .CI(DP_OP_423J2_125_3477_n1250), .CO(
        DP_OP_423J2_125_3477_n1062), .S(DP_OP_423J2_125_3477_n1063) );
  FADDX1_HVT DP_OP_423J2_125_3477_U624 ( .A(DP_OP_423J2_125_3477_n1069), .B(
        DP_OP_423J2_125_3477_n1067), .CI(DP_OP_423J2_125_3477_n1248), .CO(
        DP_OP_423J2_125_3477_n1060), .S(DP_OP_423J2_125_3477_n1061) );
  FADDX1_HVT DP_OP_423J2_125_3477_U623 ( .A(DP_OP_423J2_125_3477_n1065), .B(
        DP_OP_423J2_125_3477_n1246), .CI(DP_OP_423J2_125_3477_n1063), .CO(
        DP_OP_423J2_125_3477_n1058), .S(DP_OP_423J2_125_3477_n1059) );
  OR2X1_HVT DP_OP_423J2_125_3477_U622 ( .A1(DP_OP_423J2_125_3477_n1997), .A2(
        DP_OP_423J2_125_3477_n2699), .Y(DP_OP_423J2_125_3477_n1056) );
  FADDX1_HVT DP_OP_423J2_125_3477_U620 ( .A(DP_OP_423J2_125_3477_n2085), .B(
        DP_OP_423J2_125_3477_n2041), .CI(DP_OP_423J2_125_3477_n2742), .CO(
        DP_OP_423J2_125_3477_n1054), .S(DP_OP_423J2_125_3477_n1055) );
  FADDX1_HVT DP_OP_423J2_125_3477_U619 ( .A(DP_OP_423J2_125_3477_n2786), .B(
        DP_OP_423J2_125_3477_n2437), .CI(DP_OP_423J2_125_3477_n1953), .CO(
        DP_OP_423J2_125_3477_n1052), .S(DP_OP_423J2_125_3477_n1053) );
  FADDX1_HVT DP_OP_423J2_125_3477_U618 ( .A(DP_OP_423J2_125_3477_n2657), .B(
        DP_OP_423J2_125_3477_n2569), .CI(DP_OP_423J2_125_3477_n2481), .CO(
        DP_OP_423J2_125_3477_n1050), .S(DP_OP_423J2_125_3477_n1051) );
  FADDX1_HVT DP_OP_423J2_125_3477_U617 ( .A(DP_OP_423J2_125_3477_n1865), .B(
        DP_OP_423J2_125_3477_n2173), .CI(DP_OP_423J2_125_3477_n2525), .CO(
        DP_OP_423J2_125_3477_n1048), .S(DP_OP_423J2_125_3477_n1049) );
  FADDX1_HVT DP_OP_423J2_125_3477_U616 ( .A(DP_OP_423J2_125_3477_n2129), .B(
        DP_OP_423J2_125_3477_n2874), .CI(DP_OP_423J2_125_3477_n1909), .CO(
        DP_OP_423J2_125_3477_n1046), .S(DP_OP_423J2_125_3477_n1047) );
  FADDX1_HVT DP_OP_423J2_125_3477_U615 ( .A(DP_OP_423J2_125_3477_n2349), .B(
        DP_OP_423J2_125_3477_n2261), .CI(DP_OP_423J2_125_3477_n1821), .CO(
        DP_OP_423J2_125_3477_n1044), .S(DP_OP_423J2_125_3477_n1045) );
  FADDX1_HVT DP_OP_423J2_125_3477_U614 ( .A(DP_OP_423J2_125_3477_n2613), .B(
        DP_OP_423J2_125_3477_n2305), .CI(DP_OP_423J2_125_3477_n2830), .CO(
        DP_OP_423J2_125_3477_n1042), .S(DP_OP_423J2_125_3477_n1043) );
  FADDX1_HVT DP_OP_423J2_125_3477_U613 ( .A(DP_OP_423J2_125_3477_n1777), .B(
        DP_OP_423J2_125_3477_n2393), .CI(DP_OP_423J2_125_3477_n2763), .CO(
        DP_OP_423J2_125_3477_n1040), .S(DP_OP_423J2_125_3477_n1041) );
  FADDX1_HVT DP_OP_423J2_125_3477_U612 ( .A(DP_OP_423J2_125_3477_n1842), .B(
        DP_OP_423J2_125_3477_n1960), .CI(DP_OP_423J2_125_3477_n1886), .CO(
        DP_OP_423J2_125_3477_n1038), .S(DP_OP_423J2_125_3477_n1039) );
  FADDX1_HVT DP_OP_423J2_125_3477_U611 ( .A(DP_OP_423J2_125_3477_n2634), .B(
        DP_OP_423J2_125_3477_n2719), .CI(DP_OP_423J2_125_3477_n2444), .CO(
        DP_OP_423J2_125_3477_n1036), .S(DP_OP_423J2_125_3477_n1037) );
  FADDX1_HVT DP_OP_423J2_125_3477_U610 ( .A(DP_OP_423J2_125_3477_n2106), .B(
        DP_OP_423J2_125_3477_n2407), .CI(DP_OP_423J2_125_3477_n2502), .CO(
        DP_OP_423J2_125_3477_n1034), .S(DP_OP_423J2_125_3477_n1035) );
  FADDX1_HVT DP_OP_423J2_125_3477_U609 ( .A(DP_OP_423J2_125_3477_n2590), .B(
        DP_OP_423J2_125_3477_n2143), .CI(DP_OP_423J2_125_3477_n2851), .CO(
        DP_OP_423J2_125_3477_n1032), .S(DP_OP_423J2_125_3477_n1033) );
  FADDX1_HVT DP_OP_423J2_125_3477_U608 ( .A(DP_OP_423J2_125_3477_n2458), .B(
        DP_OP_423J2_125_3477_n2532), .CI(DP_OP_423J2_125_3477_n2092), .CO(
        DP_OP_423J2_125_3477_n1030), .S(DP_OP_423J2_125_3477_n1031) );
  FADDX1_HVT DP_OP_423J2_125_3477_U607 ( .A(DP_OP_423J2_125_3477_n2414), .B(
        DP_OP_423J2_125_3477_n2217), .CI(DP_OP_423J2_125_3477_n2224), .CO(
        DP_OP_423J2_125_3477_n1028), .S(DP_OP_423J2_125_3477_n1029) );
  FADDX1_HVT DP_OP_423J2_125_3477_U606 ( .A(DP_OP_423J2_125_3477_n2194), .B(
        DP_OP_423J2_125_3477_n2627), .CI(DP_OP_423J2_125_3477_n2495), .CO(
        DP_OP_423J2_125_3477_n1026), .S(DP_OP_423J2_125_3477_n1027) );
  FADDX1_HVT DP_OP_423J2_125_3477_U605 ( .A(DP_OP_423J2_125_3477_n2546), .B(
        DP_OP_423J2_125_3477_n1974), .CI(DP_OP_423J2_125_3477_n1835), .CO(
        DP_OP_423J2_125_3477_n1024), .S(DP_OP_423J2_125_3477_n1025) );
  FADDX1_HVT DP_OP_423J2_125_3477_U604 ( .A(DP_OP_423J2_125_3477_n2837), .B(
        DP_OP_423J2_125_3477_n2678), .CI(DP_OP_423J2_125_3477_n2583), .CO(
        DP_OP_423J2_125_3477_n1022), .S(DP_OP_423J2_125_3477_n1023) );
  FADDX1_HVT DP_OP_423J2_125_3477_U603 ( .A(DP_OP_423J2_125_3477_n2326), .B(
        DP_OP_423J2_125_3477_n2749), .CI(DP_OP_423J2_125_3477_n2018), .CO(
        DP_OP_423J2_125_3477_n1020), .S(DP_OP_423J2_125_3477_n1021) );
  FADDX1_HVT DP_OP_423J2_125_3477_U602 ( .A(DP_OP_423J2_125_3477_n2881), .B(
        DP_OP_423J2_125_3477_n2055), .CI(DP_OP_423J2_125_3477_n2319), .CO(
        DP_OP_423J2_125_3477_n1018), .S(DP_OP_423J2_125_3477_n1019) );
  FADDX1_HVT DP_OP_423J2_125_3477_U601 ( .A(DP_OP_423J2_125_3477_n2062), .B(
        DP_OP_423J2_125_3477_n2356), .CI(DP_OP_423J2_125_3477_n2888), .CO(
        DP_OP_423J2_125_3477_n1016), .S(DP_OP_423J2_125_3477_n1017) );
  FADDX1_HVT DP_OP_423J2_125_3477_U600 ( .A(DP_OP_423J2_125_3477_n2282), .B(
        DP_OP_423J2_125_3477_n2238), .CI(DP_OP_423J2_125_3477_n2275), .CO(
        DP_OP_423J2_125_3477_n1014), .S(DP_OP_423J2_125_3477_n1015) );
  FADDX1_HVT DP_OP_423J2_125_3477_U599 ( .A(DP_OP_423J2_125_3477_n2136), .B(
        DP_OP_423J2_125_3477_n2099), .CI(DP_OP_423J2_125_3477_n2800), .CO(
        DP_OP_423J2_125_3477_n1012), .S(DP_OP_423J2_125_3477_n1013) );
  FADDX1_HVT DP_OP_423J2_125_3477_U598 ( .A(DP_OP_423J2_125_3477_n2268), .B(
        DP_OP_423J2_125_3477_n2488), .CI(DP_OP_423J2_125_3477_n1923), .CO(
        DP_OP_423J2_125_3477_n1010), .S(DP_OP_423J2_125_3477_n1011) );
  FADDX1_HVT DP_OP_423J2_125_3477_U597 ( .A(DP_OP_423J2_125_3477_n2576), .B(
        DP_OP_423J2_125_3477_n2451), .CI(DP_OP_423J2_125_3477_n2370), .CO(
        DP_OP_423J2_125_3477_n1008), .S(DP_OP_423J2_125_3477_n1009) );
  FADDX1_HVT DP_OP_423J2_125_3477_U596 ( .A(DP_OP_423J2_125_3477_n2671), .B(
        DP_OP_423J2_125_3477_n1879), .CI(DP_OP_423J2_125_3477_n2756), .CO(
        DP_OP_423J2_125_3477_n1006), .S(DP_OP_423J2_125_3477_n1007) );
  FADDX1_HVT DP_OP_423J2_125_3477_U595 ( .A(DP_OP_423J2_125_3477_n2664), .B(
        DP_OP_423J2_125_3477_n2150), .CI(DP_OP_423J2_125_3477_n1244), .CO(
        DP_OP_423J2_125_3477_n1004), .S(DP_OP_423J2_125_3477_n1005) );
  FADDX1_HVT DP_OP_423J2_125_3477_U594 ( .A(DP_OP_423J2_125_3477_n2539), .B(
        DP_OP_423J2_125_3477_n2895), .CI(DP_OP_423J2_125_3477_n2807), .CO(
        DP_OP_423J2_125_3477_n1002), .S(DP_OP_423J2_125_3477_n1003) );
  FADDX1_HVT DP_OP_423J2_125_3477_U593 ( .A(DP_OP_423J2_125_3477_n2705), .B(
        DP_OP_423J2_125_3477_n2712), .CI(DP_OP_423J2_125_3477_n1828), .CO(
        DP_OP_423J2_125_3477_n1000), .S(DP_OP_423J2_125_3477_n1001) );
  FADDX1_HVT DP_OP_423J2_125_3477_U592 ( .A(DP_OP_423J2_125_3477_n2048), .B(
        DP_OP_423J2_125_3477_n2231), .CI(DP_OP_423J2_125_3477_n2180), .CO(
        DP_OP_423J2_125_3477_n998), .S(DP_OP_423J2_125_3477_n999) );
  FADDX1_HVT DP_OP_423J2_125_3477_U591 ( .A(DP_OP_423J2_125_3477_n2312), .B(
        DP_OP_423J2_125_3477_n2187), .CI(DP_OP_423J2_125_3477_n1916), .CO(
        DP_OP_423J2_125_3477_n996), .S(DP_OP_423J2_125_3477_n997) );
  FADDX1_HVT DP_OP_423J2_125_3477_U590 ( .A(DP_OP_423J2_125_3477_n1930), .B(
        DP_OP_423J2_125_3477_n2004), .CI(DP_OP_423J2_125_3477_n2793), .CO(
        DP_OP_423J2_125_3477_n994), .S(DP_OP_423J2_125_3477_n995) );
  FADDX1_HVT DP_OP_423J2_125_3477_U589 ( .A(DP_OP_423J2_125_3477_n2844), .B(
        DP_OP_423J2_125_3477_n2363), .CI(DP_OP_423J2_125_3477_n2620), .CO(
        DP_OP_423J2_125_3477_n992), .S(DP_OP_423J2_125_3477_n993) );
  FADDX1_HVT DP_OP_423J2_125_3477_U588 ( .A(DP_OP_423J2_125_3477_n2400), .B(
        DP_OP_423J2_125_3477_n1872), .CI(DP_OP_423J2_125_3477_n1967), .CO(
        DP_OP_423J2_125_3477_n990), .S(DP_OP_423J2_125_3477_n991) );
  FADDX1_HVT DP_OP_423J2_125_3477_U587 ( .A(DP_OP_423J2_125_3477_n2011), .B(
        DP_OP_423J2_125_3477_n1242), .CI(DP_OP_423J2_125_3477_n1240), .CO(
        DP_OP_423J2_125_3477_n988), .S(DP_OP_423J2_125_3477_n989) );
  FADDX1_HVT DP_OP_423J2_125_3477_U586 ( .A(DP_OP_423J2_125_3477_n1238), .B(
        DP_OP_423J2_125_3477_n1230), .CI(DP_OP_423J2_125_3477_n1057), .CO(
        DP_OP_423J2_125_3477_n986), .S(DP_OP_423J2_125_3477_n987) );
  FADDX1_HVT DP_OP_423J2_125_3477_U585 ( .A(DP_OP_423J2_125_3477_n1236), .B(
        DP_OP_423J2_125_3477_n1234), .CI(DP_OP_423J2_125_3477_n1232), .CO(
        DP_OP_423J2_125_3477_n984), .S(DP_OP_423J2_125_3477_n985) );
  FADDX1_HVT DP_OP_423J2_125_3477_U584 ( .A(DP_OP_423J2_125_3477_n1228), .B(
        DP_OP_423J2_125_3477_n1226), .CI(DP_OP_423J2_125_3477_n1224), .CO(
        DP_OP_423J2_125_3477_n982), .S(DP_OP_423J2_125_3477_n983) );
  FADDX1_HVT DP_OP_423J2_125_3477_U583 ( .A(DP_OP_423J2_125_3477_n1222), .B(
        DP_OP_423J2_125_3477_n1206), .CI(DP_OP_423J2_125_3477_n1208), .CO(
        DP_OP_423J2_125_3477_n980), .S(DP_OP_423J2_125_3477_n981) );
  FADDX1_HVT DP_OP_423J2_125_3477_U582 ( .A(DP_OP_423J2_125_3477_n1220), .B(
        DP_OP_423J2_125_3477_n1210), .CI(DP_OP_423J2_125_3477_n1212), .CO(
        DP_OP_423J2_125_3477_n978), .S(DP_OP_423J2_125_3477_n979) );
  FADDX1_HVT DP_OP_423J2_125_3477_U581 ( .A(DP_OP_423J2_125_3477_n1218), .B(
        DP_OP_423J2_125_3477_n1214), .CI(DP_OP_423J2_125_3477_n1216), .CO(
        DP_OP_423J2_125_3477_n976), .S(DP_OP_423J2_125_3477_n977) );
  FADDX1_HVT DP_OP_423J2_125_3477_U580 ( .A(DP_OP_423J2_125_3477_n1202), .B(
        DP_OP_423J2_125_3477_n1194), .CI(DP_OP_423J2_125_3477_n1178), .CO(
        DP_OP_423J2_125_3477_n974), .S(DP_OP_423J2_125_3477_n975) );
  FADDX1_HVT DP_OP_423J2_125_3477_U579 ( .A(DP_OP_423J2_125_3477_n1200), .B(
        DP_OP_423J2_125_3477_n1196), .CI(DP_OP_423J2_125_3477_n1180), .CO(
        DP_OP_423J2_125_3477_n972), .S(DP_OP_423J2_125_3477_n973) );
  FADDX1_HVT DP_OP_423J2_125_3477_U578 ( .A(DP_OP_423J2_125_3477_n1204), .B(
        DP_OP_423J2_125_3477_n1198), .CI(DP_OP_423J2_125_3477_n1182), .CO(
        DP_OP_423J2_125_3477_n970), .S(DP_OP_423J2_125_3477_n971) );
  FADDX1_HVT DP_OP_423J2_125_3477_U577 ( .A(DP_OP_423J2_125_3477_n1047), .B(
        DP_OP_423J2_125_3477_n1186), .CI(DP_OP_423J2_125_3477_n1184), .CO(
        DP_OP_423J2_125_3477_n968), .S(DP_OP_423J2_125_3477_n969) );
  FADDX1_HVT DP_OP_423J2_125_3477_U576 ( .A(DP_OP_423J2_125_3477_n1043), .B(
        DP_OP_423J2_125_3477_n1190), .CI(DP_OP_423J2_125_3477_n1188), .CO(
        DP_OP_423J2_125_3477_n966), .S(DP_OP_423J2_125_3477_n967) );
  FADDX1_HVT DP_OP_423J2_125_3477_U575 ( .A(DP_OP_423J2_125_3477_n1045), .B(
        DP_OP_423J2_125_3477_n1055), .CI(DP_OP_423J2_125_3477_n1192), .CO(
        DP_OP_423J2_125_3477_n964), .S(DP_OP_423J2_125_3477_n965) );
  FADDX1_HVT DP_OP_423J2_125_3477_U574 ( .A(DP_OP_423J2_125_3477_n1053), .B(
        DP_OP_423J2_125_3477_n1051), .CI(DP_OP_423J2_125_3477_n1049), .CO(
        DP_OP_423J2_125_3477_n962), .S(DP_OP_423J2_125_3477_n963) );
  FADDX1_HVT DP_OP_423J2_125_3477_U573 ( .A(DP_OP_423J2_125_3477_n1041), .B(
        DP_OP_423J2_125_3477_n1019), .CI(DP_OP_423J2_125_3477_n1021), .CO(
        DP_OP_423J2_125_3477_n960), .S(DP_OP_423J2_125_3477_n961) );
  FADDX1_HVT DP_OP_423J2_125_3477_U572 ( .A(DP_OP_423J2_125_3477_n1033), .B(
        DP_OP_423J2_125_3477_n1027), .CI(DP_OP_423J2_125_3477_n1029), .CO(
        DP_OP_423J2_125_3477_n958), .S(DP_OP_423J2_125_3477_n959) );
  FADDX1_HVT DP_OP_423J2_125_3477_U571 ( .A(DP_OP_423J2_125_3477_n1025), .B(
        DP_OP_423J2_125_3477_n1039), .CI(DP_OP_423J2_125_3477_n1037), .CO(
        DP_OP_423J2_125_3477_n956), .S(DP_OP_423J2_125_3477_n957) );
  FADDX1_HVT DP_OP_423J2_125_3477_U570 ( .A(DP_OP_423J2_125_3477_n1031), .B(
        DP_OP_423J2_125_3477_n1023), .CI(DP_OP_423J2_125_3477_n1035), .CO(
        DP_OP_423J2_125_3477_n954), .S(DP_OP_423J2_125_3477_n955) );
  FADDX1_HVT DP_OP_423J2_125_3477_U569 ( .A(DP_OP_423J2_125_3477_n1013), .B(
        DP_OP_423J2_125_3477_n1007), .CI(DP_OP_423J2_125_3477_n991), .CO(
        DP_OP_423J2_125_3477_n952), .S(DP_OP_423J2_125_3477_n953) );
  FADDX1_HVT DP_OP_423J2_125_3477_U568 ( .A(DP_OP_423J2_125_3477_n1017), .B(
        DP_OP_423J2_125_3477_n1009), .CI(DP_OP_423J2_125_3477_n993), .CO(
        DP_OP_423J2_125_3477_n950), .S(DP_OP_423J2_125_3477_n951) );
  FADDX1_HVT DP_OP_423J2_125_3477_U567 ( .A(DP_OP_423J2_125_3477_n1011), .B(
        DP_OP_423J2_125_3477_n1015), .CI(DP_OP_423J2_125_3477_n995), .CO(
        DP_OP_423J2_125_3477_n948), .S(DP_OP_423J2_125_3477_n949) );
  FADDX1_HVT DP_OP_423J2_125_3477_U566 ( .A(DP_OP_423J2_125_3477_n1005), .B(
        DP_OP_423J2_125_3477_n997), .CI(DP_OP_423J2_125_3477_n1174), .CO(
        DP_OP_423J2_125_3477_n946), .S(DP_OP_423J2_125_3477_n947) );
  FADDX1_HVT DP_OP_423J2_125_3477_U565 ( .A(DP_OP_423J2_125_3477_n1003), .B(
        DP_OP_423J2_125_3477_n999), .CI(DP_OP_423J2_125_3477_n1172), .CO(
        DP_OP_423J2_125_3477_n944), .S(DP_OP_423J2_125_3477_n945) );
  FADDX1_HVT DP_OP_423J2_125_3477_U564 ( .A(DP_OP_423J2_125_3477_n1001), .B(
        DP_OP_423J2_125_3477_n1176), .CI(DP_OP_423J2_125_3477_n1170), .CO(
        DP_OP_423J2_125_3477_n942), .S(DP_OP_423J2_125_3477_n943) );
  FADDX1_HVT DP_OP_423J2_125_3477_U563 ( .A(DP_OP_423J2_125_3477_n1168), .B(
        DP_OP_423J2_125_3477_n1164), .CI(DP_OP_423J2_125_3477_n1166), .CO(
        DP_OP_423J2_125_3477_n940), .S(DP_OP_423J2_125_3477_n941) );
  FADDX1_HVT DP_OP_423J2_125_3477_U562 ( .A(DP_OP_423J2_125_3477_n1158), .B(
        DP_OP_423J2_125_3477_n989), .CI(DP_OP_423J2_125_3477_n985), .CO(
        DP_OP_423J2_125_3477_n938), .S(DP_OP_423J2_125_3477_n939) );
  FADDX1_HVT DP_OP_423J2_125_3477_U561 ( .A(DP_OP_423J2_125_3477_n1162), .B(
        DP_OP_423J2_125_3477_n1160), .CI(DP_OP_423J2_125_3477_n987), .CO(
        DP_OP_423J2_125_3477_n936), .S(DP_OP_423J2_125_3477_n937) );
  FADDX1_HVT DP_OP_423J2_125_3477_U560 ( .A(DP_OP_423J2_125_3477_n1156), .B(
        DP_OP_423J2_125_3477_n1150), .CI(DP_OP_423J2_125_3477_n1152), .CO(
        DP_OP_423J2_125_3477_n934), .S(DP_OP_423J2_125_3477_n935) );
  FADDX1_HVT DP_OP_423J2_125_3477_U559 ( .A(DP_OP_423J2_125_3477_n1154), .B(
        DP_OP_423J2_125_3477_n1148), .CI(DP_OP_423J2_125_3477_n983), .CO(
        DP_OP_423J2_125_3477_n932), .S(DP_OP_423J2_125_3477_n933) );
  FADDX1_HVT DP_OP_423J2_125_3477_U558 ( .A(DP_OP_423J2_125_3477_n1146), .B(
        DP_OP_423J2_125_3477_n979), .CI(DP_OP_423J2_125_3477_n981), .CO(
        DP_OP_423J2_125_3477_n930), .S(DP_OP_423J2_125_3477_n931) );
  FADDX1_HVT DP_OP_423J2_125_3477_U557 ( .A(DP_OP_423J2_125_3477_n1144), .B(
        DP_OP_423J2_125_3477_n1142), .CI(DP_OP_423J2_125_3477_n977), .CO(
        DP_OP_423J2_125_3477_n928), .S(DP_OP_423J2_125_3477_n929) );
  FADDX1_HVT DP_OP_423J2_125_3477_U556 ( .A(DP_OP_423J2_125_3477_n1140), .B(
        DP_OP_423J2_125_3477_n971), .CI(DP_OP_423J2_125_3477_n1132), .CO(
        DP_OP_423J2_125_3477_n926), .S(DP_OP_423J2_125_3477_n927) );
  FADDX1_HVT DP_OP_423J2_125_3477_U555 ( .A(DP_OP_423J2_125_3477_n1138), .B(
        DP_OP_423J2_125_3477_n973), .CI(DP_OP_423J2_125_3477_n1134), .CO(
        DP_OP_423J2_125_3477_n924), .S(DP_OP_423J2_125_3477_n925) );
  FADDX1_HVT DP_OP_423J2_125_3477_U554 ( .A(DP_OP_423J2_125_3477_n1136), .B(
        DP_OP_423J2_125_3477_n975), .CI(DP_OP_423J2_125_3477_n963), .CO(
        DP_OP_423J2_125_3477_n922), .S(DP_OP_423J2_125_3477_n923) );
  FADDX1_HVT DP_OP_423J2_125_3477_U553 ( .A(DP_OP_423J2_125_3477_n965), .B(
        DP_OP_423J2_125_3477_n969), .CI(DP_OP_423J2_125_3477_n967), .CO(
        DP_OP_423J2_125_3477_n920), .S(DP_OP_423J2_125_3477_n921) );
  FADDX1_HVT DP_OP_423J2_125_3477_U552 ( .A(DP_OP_423J2_125_3477_n961), .B(
        DP_OP_423J2_125_3477_n959), .CI(DP_OP_423J2_125_3477_n1130), .CO(
        DP_OP_423J2_125_3477_n918), .S(DP_OP_423J2_125_3477_n919) );
  FADDX1_HVT DP_OP_423J2_125_3477_U551 ( .A(DP_OP_423J2_125_3477_n955), .B(
        DP_OP_423J2_125_3477_n957), .CI(DP_OP_423J2_125_3477_n951), .CO(
        DP_OP_423J2_125_3477_n916), .S(DP_OP_423J2_125_3477_n917) );
  FADDX1_HVT DP_OP_423J2_125_3477_U550 ( .A(DP_OP_423J2_125_3477_n949), .B(
        DP_OP_423J2_125_3477_n1128), .CI(DP_OP_423J2_125_3477_n945), .CO(
        DP_OP_423J2_125_3477_n914), .S(DP_OP_423J2_125_3477_n915) );
  FADDX1_HVT DP_OP_423J2_125_3477_U549 ( .A(DP_OP_423J2_125_3477_n953), .B(
        DP_OP_423J2_125_3477_n947), .CI(DP_OP_423J2_125_3477_n1124), .CO(
        DP_OP_423J2_125_3477_n912), .S(DP_OP_423J2_125_3477_n913) );
  FADDX1_HVT DP_OP_423J2_125_3477_U548 ( .A(DP_OP_423J2_125_3477_n1126), .B(
        DP_OP_423J2_125_3477_n1122), .CI(DP_OP_423J2_125_3477_n943), .CO(
        DP_OP_423J2_125_3477_n910), .S(DP_OP_423J2_125_3477_n911) );
  FADDX1_HVT DP_OP_423J2_125_3477_U547 ( .A(DP_OP_423J2_125_3477_n1120), .B(
        DP_OP_423J2_125_3477_n1118), .CI(DP_OP_423J2_125_3477_n941), .CO(
        DP_OP_423J2_125_3477_n908), .S(DP_OP_423J2_125_3477_n909) );
  FADDX1_HVT DP_OP_423J2_125_3477_U546 ( .A(DP_OP_423J2_125_3477_n1116), .B(
        DP_OP_423J2_125_3477_n1114), .CI(DP_OP_423J2_125_3477_n1112), .CO(
        DP_OP_423J2_125_3477_n906), .S(DP_OP_423J2_125_3477_n907) );
  FADDX1_HVT DP_OP_423J2_125_3477_U545 ( .A(DP_OP_423J2_125_3477_n1110), .B(
        DP_OP_423J2_125_3477_n939), .CI(DP_OP_423J2_125_3477_n935), .CO(
        DP_OP_423J2_125_3477_n904), .S(DP_OP_423J2_125_3477_n905) );
  FADDX1_HVT DP_OP_423J2_125_3477_U544 ( .A(DP_OP_423J2_125_3477_n937), .B(
        DP_OP_423J2_125_3477_n1108), .CI(DP_OP_423J2_125_3477_n933), .CO(
        DP_OP_423J2_125_3477_n902), .S(DP_OP_423J2_125_3477_n903) );
  FADDX1_HVT DP_OP_423J2_125_3477_U543 ( .A(DP_OP_423J2_125_3477_n931), .B(
        DP_OP_423J2_125_3477_n1106), .CI(DP_OP_423J2_125_3477_n1104), .CO(
        DP_OP_423J2_125_3477_n900), .S(DP_OP_423J2_125_3477_n901) );
  FADDX1_HVT DP_OP_423J2_125_3477_U542 ( .A(DP_OP_423J2_125_3477_n929), .B(
        DP_OP_423J2_125_3477_n1102), .CI(DP_OP_423J2_125_3477_n923), .CO(
        DP_OP_423J2_125_3477_n898), .S(DP_OP_423J2_125_3477_n899) );
  FADDX1_HVT DP_OP_423J2_125_3477_U541 ( .A(DP_OP_423J2_125_3477_n925), .B(
        DP_OP_423J2_125_3477_n927), .CI(DP_OP_423J2_125_3477_n1100), .CO(
        DP_OP_423J2_125_3477_n896), .S(DP_OP_423J2_125_3477_n897) );
  FADDX1_HVT DP_OP_423J2_125_3477_U540 ( .A(DP_OP_423J2_125_3477_n921), .B(
        DP_OP_423J2_125_3477_n1098), .CI(DP_OP_423J2_125_3477_n919), .CO(
        DP_OP_423J2_125_3477_n894), .S(DP_OP_423J2_125_3477_n895) );
  FADDX1_HVT DP_OP_423J2_125_3477_U539 ( .A(DP_OP_423J2_125_3477_n917), .B(
        DP_OP_423J2_125_3477_n915), .CI(DP_OP_423J2_125_3477_n1096), .CO(
        DP_OP_423J2_125_3477_n892), .S(DP_OP_423J2_125_3477_n893) );
  FADDX1_HVT DP_OP_423J2_125_3477_U538 ( .A(DP_OP_423J2_125_3477_n913), .B(
        DP_OP_423J2_125_3477_n1094), .CI(DP_OP_423J2_125_3477_n911), .CO(
        DP_OP_423J2_125_3477_n890), .S(DP_OP_423J2_125_3477_n891) );
  FADDX1_HVT DP_OP_423J2_125_3477_U537 ( .A(DP_OP_423J2_125_3477_n1092), .B(
        DP_OP_423J2_125_3477_n1090), .CI(DP_OP_423J2_125_3477_n909), .CO(
        DP_OP_423J2_125_3477_n888), .S(DP_OP_423J2_125_3477_n889) );
  FADDX1_HVT DP_OP_423J2_125_3477_U536 ( .A(DP_OP_423J2_125_3477_n1088), .B(
        DP_OP_423J2_125_3477_n907), .CI(DP_OP_423J2_125_3477_n1086), .CO(
        DP_OP_423J2_125_3477_n886), .S(DP_OP_423J2_125_3477_n887) );
  FADDX1_HVT DP_OP_423J2_125_3477_U535 ( .A(DP_OP_423J2_125_3477_n905), .B(
        DP_OP_423J2_125_3477_n903), .CI(DP_OP_423J2_125_3477_n1084), .CO(
        DP_OP_423J2_125_3477_n884), .S(DP_OP_423J2_125_3477_n885) );
  FADDX1_HVT DP_OP_423J2_125_3477_U534 ( .A(DP_OP_423J2_125_3477_n901), .B(
        DP_OP_423J2_125_3477_n1082), .CI(DP_OP_423J2_125_3477_n899), .CO(
        DP_OP_423J2_125_3477_n882), .S(DP_OP_423J2_125_3477_n883) );
  FADDX1_HVT DP_OP_423J2_125_3477_U533 ( .A(DP_OP_423J2_125_3477_n897), .B(
        DP_OP_423J2_125_3477_n1080), .CI(DP_OP_423J2_125_3477_n895), .CO(
        DP_OP_423J2_125_3477_n880), .S(DP_OP_423J2_125_3477_n881) );
  FADDX1_HVT DP_OP_423J2_125_3477_U532 ( .A(DP_OP_423J2_125_3477_n1078), .B(
        DP_OP_423J2_125_3477_n893), .CI(DP_OP_423J2_125_3477_n1076), .CO(
        DP_OP_423J2_125_3477_n878), .S(DP_OP_423J2_125_3477_n879) );
  FADDX1_HVT DP_OP_423J2_125_3477_U531 ( .A(DP_OP_423J2_125_3477_n891), .B(
        DP_OP_423J2_125_3477_n1074), .CI(DP_OP_423J2_125_3477_n889), .CO(
        DP_OP_423J2_125_3477_n876), .S(DP_OP_423J2_125_3477_n877) );
  FADDX1_HVT DP_OP_423J2_125_3477_U530 ( .A(DP_OP_423J2_125_3477_n1072), .B(
        DP_OP_423J2_125_3477_n887), .CI(DP_OP_423J2_125_3477_n885), .CO(
        DP_OP_423J2_125_3477_n874), .S(DP_OP_423J2_125_3477_n875) );
  FADDX1_HVT DP_OP_423J2_125_3477_U529 ( .A(DP_OP_423J2_125_3477_n1070), .B(
        DP_OP_423J2_125_3477_n883), .CI(DP_OP_423J2_125_3477_n1068), .CO(
        DP_OP_423J2_125_3477_n872), .S(DP_OP_423J2_125_3477_n873) );
  FADDX1_HVT DP_OP_423J2_125_3477_U528 ( .A(DP_OP_423J2_125_3477_n881), .B(
        DP_OP_423J2_125_3477_n1066), .CI(DP_OP_423J2_125_3477_n879), .CO(
        DP_OP_423J2_125_3477_n870), .S(DP_OP_423J2_125_3477_n871) );
  FADDX1_HVT DP_OP_423J2_125_3477_U527 ( .A(DP_OP_423J2_125_3477_n877), .B(
        DP_OP_423J2_125_3477_n1064), .CI(DP_OP_423J2_125_3477_n875), .CO(
        DP_OP_423J2_125_3477_n868), .S(DP_OP_423J2_125_3477_n869) );
  FADDX1_HVT DP_OP_423J2_125_3477_U526 ( .A(DP_OP_423J2_125_3477_n1062), .B(
        DP_OP_423J2_125_3477_n873), .CI(DP_OP_423J2_125_3477_n871), .CO(
        DP_OP_423J2_125_3477_n866), .S(DP_OP_423J2_125_3477_n867) );
  FADDX1_HVT DP_OP_423J2_125_3477_U525 ( .A(DP_OP_423J2_125_3477_n1060), .B(
        DP_OP_423J2_125_3477_n869), .CI(DP_OP_423J2_125_3477_n1058), .CO(
        DP_OP_423J2_125_3477_n864), .S(DP_OP_423J2_125_3477_n865) );
  FADDX1_HVT DP_OP_423J2_125_3477_U524 ( .A(DP_OP_423J2_125_3477_n1996), .B(
        DP_OP_423J2_125_3477_n2718), .CI(DP_OP_423J2_125_3477_n1885), .CO(
        DP_OP_423J2_125_3477_n862), .S(DP_OP_423J2_125_3477_n863) );
  FADDX1_HVT DP_OP_423J2_125_3477_U523 ( .A(DP_OP_423J2_125_3477_n2698), .B(
        DP_OP_423J2_125_3477_n2172), .CI(DP_OP_423J2_125_3477_n2501), .CO(
        DP_OP_423J2_125_3477_n860), .S(DP_OP_423J2_125_3477_n861) );
  FADDX1_HVT DP_OP_423J2_125_3477_U522 ( .A(DP_OP_423J2_125_3477_n2348), .B(
        DP_OP_423J2_125_3477_n2040), .CI(DP_OP_423J2_125_3477_n2850), .CO(
        DP_OP_423J2_125_3477_n858), .S(DP_OP_423J2_125_3477_n859) );
  FADDX1_HVT DP_OP_423J2_125_3477_U521 ( .A(DP_OP_423J2_125_3477_n1864), .B(
        DP_OP_423J2_125_3477_n2524), .CI(DP_OP_423J2_125_3477_n2762), .CO(
        DP_OP_423J2_125_3477_n856), .S(DP_OP_423J2_125_3477_n857) );
  FADDX1_HVT DP_OP_423J2_125_3477_U520 ( .A(DP_OP_423J2_125_3477_n2084), .B(
        DP_OP_423J2_125_3477_n2568), .CI(DP_OP_423J2_125_3477_n1952), .CO(
        DP_OP_423J2_125_3477_n854), .S(DP_OP_423J2_125_3477_n855) );
  FADDX1_HVT DP_OP_423J2_125_3477_U519 ( .A(DP_OP_423J2_125_3477_n2656), .B(
        DP_OP_423J2_125_3477_n1908), .CI(DP_OP_423J2_125_3477_n2741), .CO(
        DP_OP_423J2_125_3477_n852), .S(DP_OP_423J2_125_3477_n853) );
  FADDX1_HVT DP_OP_423J2_125_3477_U518 ( .A(DP_OP_423J2_125_3477_n2304), .B(
        DP_OP_423J2_125_3477_n2436), .CI(DP_OP_423J2_125_3477_n2480), .CO(
        DP_OP_423J2_125_3477_n850), .S(DP_OP_423J2_125_3477_n851) );
  FADDX1_HVT DP_OP_423J2_125_3477_U517 ( .A(DP_OP_423J2_125_3477_n2829), .B(
        DP_OP_423J2_125_3477_n1820), .CI(DP_OP_423J2_125_3477_n2873), .CO(
        DP_OP_423J2_125_3477_n848), .S(DP_OP_423J2_125_3477_n849) );
  FADDX1_HVT DP_OP_423J2_125_3477_U516 ( .A(DP_OP_423J2_125_3477_n2785), .B(
        DP_OP_423J2_125_3477_n2677), .CI(DP_OP_423J2_125_3477_n1973), .CO(
        DP_OP_423J2_125_3477_n846), .S(DP_OP_423J2_125_3477_n847) );
  FADDX1_HVT DP_OP_423J2_125_3477_U515 ( .A(DP_OP_423J2_125_3477_n2612), .B(
        DP_OP_423J2_125_3477_n2457), .CI(DP_OP_423J2_125_3477_n2017), .CO(
        DP_OP_423J2_125_3477_n844), .S(DP_OP_423J2_125_3477_n845) );
  FADDX1_HVT DP_OP_423J2_125_3477_U514 ( .A(DP_OP_423J2_125_3477_n2128), .B(
        DP_OP_423J2_125_3477_n2413), .CI(DP_OP_423J2_125_3477_n2633), .CO(
        DP_OP_423J2_125_3477_n842), .S(DP_OP_423J2_125_3477_n843) );
  FADDX1_HVT DP_OP_423J2_125_3477_U513 ( .A(DP_OP_423J2_125_3477_n2260), .B(
        DP_OP_423J2_125_3477_n2589), .CI(DP_OP_423J2_125_3477_n2105), .CO(
        DP_OP_423J2_125_3477_n840), .S(DP_OP_423J2_125_3477_n841) );
  FADDX1_HVT DP_OP_423J2_125_3477_U512 ( .A(DP_OP_423J2_125_3477_n2325), .B(
        DP_OP_423J2_125_3477_n1841), .CI(DP_OP_423J2_125_3477_n2193), .CO(
        DP_OP_423J2_125_3477_n838), .S(DP_OP_423J2_125_3477_n839) );
  FADDX1_HVT DP_OP_423J2_125_3477_U511 ( .A(DP_OP_423J2_125_3477_n2545), .B(
        DP_OP_423J2_125_3477_n2061), .CI(DP_OP_423J2_125_3477_n2281), .CO(
        DP_OP_423J2_125_3477_n836), .S(DP_OP_423J2_125_3477_n837) );
  FADDX1_HVT DP_OP_423J2_125_3477_U510 ( .A(DP_OP_423J2_125_3477_n1776), .B(
        DP_OP_423J2_125_3477_n2392), .CI(DP_OP_423J2_125_3477_n2149), .CO(
        DP_OP_423J2_125_3477_n834), .S(DP_OP_423J2_125_3477_n835) );
  FADDX1_HVT DP_OP_423J2_125_3477_U509 ( .A(DP_OP_423J2_125_3477_n2836), .B(
        DP_OP_423J2_125_3477_n2237), .CI(DP_OP_423J2_125_3477_n1929), .CO(
        DP_OP_423J2_125_3477_n832), .S(DP_OP_423J2_125_3477_n833) );
  FADDX1_HVT DP_OP_423J2_125_3477_U508 ( .A(DP_OP_423J2_125_3477_n2880), .B(
        DP_OP_423J2_125_3477_n2142), .CI(DP_OP_423J2_125_3477_n2091), .CO(
        DP_OP_423J2_125_3477_n830), .S(DP_OP_423J2_125_3477_n831) );
  FADDX1_HVT DP_OP_423J2_125_3477_U507 ( .A(DP_OP_423J2_125_3477_n2054), .B(
        DP_OP_423J2_125_3477_n2531), .CI(DP_OP_423J2_125_3477_n2223), .CO(
        DP_OP_423J2_125_3477_n828), .S(DP_OP_423J2_125_3477_n829) );
  FADDX1_HVT DP_OP_423J2_125_3477_U506 ( .A(DP_OP_423J2_125_3477_n2582), .B(
        DP_OP_423J2_125_3477_n1959), .CI(DP_OP_423J2_125_3477_n2443), .CO(
        DP_OP_423J2_125_3477_n826), .S(DP_OP_423J2_125_3477_n827) );
  FADDX1_HVT DP_OP_423J2_125_3477_U505 ( .A(DP_OP_423J2_125_3477_n2318), .B(
        DP_OP_423J2_125_3477_n2216), .CI(DP_OP_423J2_125_3477_n2406), .CO(
        DP_OP_423J2_125_3477_n824), .S(DP_OP_423J2_125_3477_n825) );
  FADDX1_HVT DP_OP_423J2_125_3477_U504 ( .A(DP_OP_423J2_125_3477_n2494), .B(
        DP_OP_423J2_125_3477_n2748), .CI(DP_OP_423J2_125_3477_n1834), .CO(
        DP_OP_423J2_125_3477_n822), .S(DP_OP_423J2_125_3477_n823) );
  FADDX1_HVT DP_OP_423J2_125_3477_U503 ( .A(DP_OP_423J2_125_3477_n2626), .B(
        DP_OP_423J2_125_3477_n2135), .CI(DP_OP_423J2_125_3477_n2267), .CO(
        DP_OP_423J2_125_3477_n820), .S(DP_OP_423J2_125_3477_n821) );
  FADDX1_HVT DP_OP_423J2_125_3477_U502 ( .A(DP_OP_423J2_125_3477_n2894), .B(
        DP_OP_423J2_125_3477_n2450), .CI(DP_OP_423J2_125_3477_n2887), .CO(
        DP_OP_423J2_125_3477_n818), .S(DP_OP_423J2_125_3477_n819) );
  FADDX1_HVT DP_OP_423J2_125_3477_U501 ( .A(DP_OP_423J2_125_3477_n2369), .B(
        DP_OP_423J2_125_3477_n2355), .CI(DP_OP_423J2_125_3477_n2799), .CO(
        DP_OP_423J2_125_3477_n816), .S(DP_OP_423J2_125_3477_n817) );
  FADDX1_HVT DP_OP_423J2_125_3477_U500 ( .A(DP_OP_423J2_125_3477_n2575), .B(
        DP_OP_423J2_125_3477_n2806), .CI(DP_OP_423J2_125_3477_n2711), .CO(
        DP_OP_423J2_125_3477_n814), .S(DP_OP_423J2_125_3477_n815) );
  FADDX1_HVT DP_OP_423J2_125_3477_U499 ( .A(DP_OP_423J2_125_3477_n2670), .B(
        DP_OP_423J2_125_3477_n1878), .CI(DP_OP_423J2_125_3477_n2755), .CO(
        DP_OP_423J2_125_3477_n812), .S(DP_OP_423J2_125_3477_n813) );
  FADDX1_HVT DP_OP_423J2_125_3477_U498 ( .A(DP_OP_423J2_125_3477_n2098), .B(
        DP_OP_423J2_125_3477_n2487), .CI(DP_OP_423J2_125_3477_n2362), .CO(
        DP_OP_423J2_125_3477_n810), .S(DP_OP_423J2_125_3477_n811) );
  FADDX1_HVT DP_OP_423J2_125_3477_U497 ( .A(DP_OP_423J2_125_3477_n2663), .B(
        DP_OP_423J2_125_3477_n2274), .CI(DP_OP_423J2_125_3477_n1827), .CO(
        DP_OP_423J2_125_3477_n808), .S(DP_OP_423J2_125_3477_n809) );
  FADDX1_HVT DP_OP_423J2_125_3477_U496 ( .A(DP_OP_423J2_125_3477_n2704), .B(
        DP_OP_423J2_125_3477_n2186), .CI(DP_OP_423J2_125_3477_n1915), .CO(
        DP_OP_423J2_125_3477_n806), .S(DP_OP_423J2_125_3477_n807) );
  FADDX1_HVT DP_OP_423J2_125_3477_U495 ( .A(DP_OP_423J2_125_3477_n2538), .B(
        DP_OP_423J2_125_3477_n2230), .CI(DP_OP_423J2_125_3477_n2179), .CO(
        DP_OP_423J2_125_3477_n804), .S(DP_OP_423J2_125_3477_n805) );
  FADDX1_HVT DP_OP_423J2_125_3477_U494 ( .A(DP_OP_423J2_125_3477_n2311), .B(
        DP_OP_423J2_125_3477_n2003), .CI(DP_OP_423J2_125_3477_n2792), .CO(
        DP_OP_423J2_125_3477_n802), .S(DP_OP_423J2_125_3477_n803) );
  FADDX1_HVT DP_OP_423J2_125_3477_U493 ( .A(DP_OP_423J2_125_3477_n2047), .B(
        DP_OP_423J2_125_3477_n1056), .CI(DP_OP_423J2_125_3477_n1966), .CO(
        DP_OP_423J2_125_3477_n800), .S(DP_OP_423J2_125_3477_n801) );
  FADDX1_HVT DP_OP_423J2_125_3477_U492 ( .A(DP_OP_423J2_125_3477_n2843), .B(
        DP_OP_423J2_125_3477_n1922), .CI(DP_OP_423J2_125_3477_n2619), .CO(
        DP_OP_423J2_125_3477_n798), .S(DP_OP_423J2_125_3477_n799) );
  FADDX1_HVT DP_OP_423J2_125_3477_U491 ( .A(DP_OP_423J2_125_3477_n2399), .B(
        DP_OP_423J2_125_3477_n2010), .CI(DP_OP_423J2_125_3477_n1871), .CO(
        DP_OP_423J2_125_3477_n796), .S(DP_OP_423J2_125_3477_n797) );
  FADDX1_HVT DP_OP_423J2_125_3477_U490 ( .A(DP_OP_423J2_125_3477_n1046), .B(
        DP_OP_423J2_125_3477_n1042), .CI(DP_OP_423J2_125_3477_n1044), .CO(
        DP_OP_423J2_125_3477_n794), .S(DP_OP_423J2_125_3477_n795) );
  FADDX1_HVT DP_OP_423J2_125_3477_U489 ( .A(DP_OP_423J2_125_3477_n1054), .B(
        DP_OP_423J2_125_3477_n1048), .CI(DP_OP_423J2_125_3477_n1050), .CO(
        DP_OP_423J2_125_3477_n792), .S(DP_OP_423J2_125_3477_n793) );
  FADDX1_HVT DP_OP_423J2_125_3477_U488 ( .A(DP_OP_423J2_125_3477_n1052), .B(
        DP_OP_423J2_125_3477_n1040), .CI(DP_OP_423J2_125_3477_n1038), .CO(
        DP_OP_423J2_125_3477_n790), .S(DP_OP_423J2_125_3477_n791) );
  FADDX1_HVT DP_OP_423J2_125_3477_U487 ( .A(DP_OP_423J2_125_3477_n1036), .B(
        DP_OP_423J2_125_3477_n1018), .CI(DP_OP_423J2_125_3477_n1020), .CO(
        DP_OP_423J2_125_3477_n788), .S(DP_OP_423J2_125_3477_n789) );
  FADDX1_HVT DP_OP_423J2_125_3477_U486 ( .A(DP_OP_423J2_125_3477_n1034), .B(
        DP_OP_423J2_125_3477_n1022), .CI(DP_OP_423J2_125_3477_n1024), .CO(
        DP_OP_423J2_125_3477_n786), .S(DP_OP_423J2_125_3477_n787) );
  FADDX1_HVT DP_OP_423J2_125_3477_U485 ( .A(DP_OP_423J2_125_3477_n1032), .B(
        DP_OP_423J2_125_3477_n1026), .CI(DP_OP_423J2_125_3477_n1028), .CO(
        DP_OP_423J2_125_3477_n784), .S(DP_OP_423J2_125_3477_n785) );
  FADDX1_HVT DP_OP_423J2_125_3477_U484 ( .A(DP_OP_423J2_125_3477_n1030), .B(
        DP_OP_423J2_125_3477_n1014), .CI(DP_OP_423J2_125_3477_n1012), .CO(
        DP_OP_423J2_125_3477_n782), .S(DP_OP_423J2_125_3477_n783) );
  FADDX1_HVT DP_OP_423J2_125_3477_U483 ( .A(DP_OP_423J2_125_3477_n1010), .B(
        DP_OP_423J2_125_3477_n1006), .CI(DP_OP_423J2_125_3477_n990), .CO(
        DP_OP_423J2_125_3477_n780), .S(DP_OP_423J2_125_3477_n781) );
  FADDX1_HVT DP_OP_423J2_125_3477_U482 ( .A(DP_OP_423J2_125_3477_n1016), .B(
        DP_OP_423J2_125_3477_n1008), .CI(DP_OP_423J2_125_3477_n992), .CO(
        DP_OP_423J2_125_3477_n778), .S(DP_OP_423J2_125_3477_n779) );
  FADDX1_HVT DP_OP_423J2_125_3477_U481 ( .A(DP_OP_423J2_125_3477_n863), .B(
        DP_OP_423J2_125_3477_n994), .CI(DP_OP_423J2_125_3477_n837), .CO(
        DP_OP_423J2_125_3477_n776), .S(DP_OP_423J2_125_3477_n777) );
  FADDX1_HVT DP_OP_423J2_125_3477_U480 ( .A(DP_OP_423J2_125_3477_n861), .B(
        DP_OP_423J2_125_3477_n996), .CI(DP_OP_423J2_125_3477_n998), .CO(
        DP_OP_423J2_125_3477_n774), .S(DP_OP_423J2_125_3477_n775) );
  FADDX1_HVT DP_OP_423J2_125_3477_U479 ( .A(DP_OP_423J2_125_3477_n851), .B(
        DP_OP_423J2_125_3477_n1000), .CI(DP_OP_423J2_125_3477_n1002), .CO(
        DP_OP_423J2_125_3477_n772), .S(DP_OP_423J2_125_3477_n773) );
  FADDX1_HVT DP_OP_423J2_125_3477_U478 ( .A(DP_OP_423J2_125_3477_n853), .B(
        DP_OP_423J2_125_3477_n839), .CI(DP_OP_423J2_125_3477_n1004), .CO(
        DP_OP_423J2_125_3477_n770), .S(DP_OP_423J2_125_3477_n771) );
  FADDX1_HVT DP_OP_423J2_125_3477_U477 ( .A(DP_OP_423J2_125_3477_n847), .B(
        DP_OP_423J2_125_3477_n843), .CI(DP_OP_423J2_125_3477_n841), .CO(
        DP_OP_423J2_125_3477_n768), .S(DP_OP_423J2_125_3477_n769) );
  FADDX1_HVT DP_OP_423J2_125_3477_U476 ( .A(DP_OP_423J2_125_3477_n849), .B(
        DP_OP_423J2_125_3477_n857), .CI(DP_OP_423J2_125_3477_n859), .CO(
        DP_OP_423J2_125_3477_n766), .S(DP_OP_423J2_125_3477_n767) );
  FADDX1_HVT DP_OP_423J2_125_3477_U475 ( .A(DP_OP_423J2_125_3477_n855), .B(
        DP_OP_423J2_125_3477_n845), .CI(DP_OP_423J2_125_3477_n835), .CO(
        DP_OP_423J2_125_3477_n764), .S(DP_OP_423J2_125_3477_n765) );
  FADDX1_HVT DP_OP_423J2_125_3477_U474 ( .A(DP_OP_423J2_125_3477_n833), .B(
        DP_OP_423J2_125_3477_n825), .CI(DP_OP_423J2_125_3477_n821), .CO(
        DP_OP_423J2_125_3477_n762), .S(DP_OP_423J2_125_3477_n763) );
  FADDX1_HVT DP_OP_423J2_125_3477_U473 ( .A(DP_OP_423J2_125_3477_n831), .B(
        DP_OP_423J2_125_3477_n829), .CI(DP_OP_423J2_125_3477_n827), .CO(
        DP_OP_423J2_125_3477_n760), .S(DP_OP_423J2_125_3477_n761) );
  FADDX1_HVT DP_OP_423J2_125_3477_U472 ( .A(DP_OP_423J2_125_3477_n823), .B(
        DP_OP_423J2_125_3477_n819), .CI(DP_OP_423J2_125_3477_n817), .CO(
        DP_OP_423J2_125_3477_n758), .S(DP_OP_423J2_125_3477_n759) );
  FADDX1_HVT DP_OP_423J2_125_3477_U471 ( .A(DP_OP_423J2_125_3477_n815), .B(
        DP_OP_423J2_125_3477_n811), .CI(DP_OP_423J2_125_3477_n797), .CO(
        DP_OP_423J2_125_3477_n756), .S(DP_OP_423J2_125_3477_n757) );
  FADDX1_HVT DP_OP_423J2_125_3477_U470 ( .A(DP_OP_423J2_125_3477_n813), .B(
        DP_OP_423J2_125_3477_n809), .CI(DP_OP_423J2_125_3477_n799), .CO(
        DP_OP_423J2_125_3477_n754), .S(DP_OP_423J2_125_3477_n755) );
  FADDX1_HVT DP_OP_423J2_125_3477_U469 ( .A(DP_OP_423J2_125_3477_n805), .B(
        DP_OP_423J2_125_3477_n801), .CI(DP_OP_423J2_125_3477_n986), .CO(
        DP_OP_423J2_125_3477_n752), .S(DP_OP_423J2_125_3477_n753) );
  FADDX1_HVT DP_OP_423J2_125_3477_U468 ( .A(DP_OP_423J2_125_3477_n807), .B(
        DP_OP_423J2_125_3477_n803), .CI(DP_OP_423J2_125_3477_n984), .CO(
        DP_OP_423J2_125_3477_n750), .S(DP_OP_423J2_125_3477_n751) );
  FADDX1_HVT DP_OP_423J2_125_3477_U467 ( .A(DP_OP_423J2_125_3477_n988), .B(
        DP_OP_423J2_125_3477_n982), .CI(DP_OP_423J2_125_3477_n976), .CO(
        DP_OP_423J2_125_3477_n748), .S(DP_OP_423J2_125_3477_n749) );
  FADDX1_HVT DP_OP_423J2_125_3477_U466 ( .A(DP_OP_423J2_125_3477_n980), .B(
        DP_OP_423J2_125_3477_n978), .CI(DP_OP_423J2_125_3477_n974), .CO(
        DP_OP_423J2_125_3477_n746), .S(DP_OP_423J2_125_3477_n747) );
  FADDX1_HVT DP_OP_423J2_125_3477_U465 ( .A(DP_OP_423J2_125_3477_n972), .B(
        DP_OP_423J2_125_3477_n970), .CI(DP_OP_423J2_125_3477_n793), .CO(
        DP_OP_423J2_125_3477_n744), .S(DP_OP_423J2_125_3477_n745) );
  FADDX1_HVT DP_OP_423J2_125_3477_U464 ( .A(DP_OP_423J2_125_3477_n968), .B(
        DP_OP_423J2_125_3477_n795), .CI(DP_OP_423J2_125_3477_n791), .CO(
        DP_OP_423J2_125_3477_n742), .S(DP_OP_423J2_125_3477_n743) );
  FADDX1_HVT DP_OP_423J2_125_3477_U463 ( .A(DP_OP_423J2_125_3477_n966), .B(
        DP_OP_423J2_125_3477_n962), .CI(DP_OP_423J2_125_3477_n964), .CO(
        DP_OP_423J2_125_3477_n740), .S(DP_OP_423J2_125_3477_n741) );
  FADDX1_HVT DP_OP_423J2_125_3477_U462 ( .A(DP_OP_423J2_125_3477_n960), .B(
        DP_OP_423J2_125_3477_n785), .CI(DP_OP_423J2_125_3477_n783), .CO(
        DP_OP_423J2_125_3477_n738), .S(DP_OP_423J2_125_3477_n739) );
  FADDX1_HVT DP_OP_423J2_125_3477_U461 ( .A(DP_OP_423J2_125_3477_n787), .B(
        DP_OP_423J2_125_3477_n789), .CI(DP_OP_423J2_125_3477_n954), .CO(
        DP_OP_423J2_125_3477_n736), .S(DP_OP_423J2_125_3477_n737) );
  FADDX1_HVT DP_OP_423J2_125_3477_U460 ( .A(DP_OP_423J2_125_3477_n958), .B(
        DP_OP_423J2_125_3477_n956), .CI(DP_OP_423J2_125_3477_n952), .CO(
        DP_OP_423J2_125_3477_n734), .S(DP_OP_423J2_125_3477_n735) );
  FADDX1_HVT DP_OP_423J2_125_3477_U459 ( .A(DP_OP_423J2_125_3477_n950), .B(
        DP_OP_423J2_125_3477_n781), .CI(DP_OP_423J2_125_3477_n944), .CO(
        DP_OP_423J2_125_3477_n732), .S(DP_OP_423J2_125_3477_n733) );
  FADDX1_HVT DP_OP_423J2_125_3477_U458 ( .A(DP_OP_423J2_125_3477_n948), .B(
        DP_OP_423J2_125_3477_n779), .CI(DP_OP_423J2_125_3477_n946), .CO(
        DP_OP_423J2_125_3477_n730), .S(DP_OP_423J2_125_3477_n731) );
  FADDX1_HVT DP_OP_423J2_125_3477_U457 ( .A(DP_OP_423J2_125_3477_n775), .B(
        DP_OP_423J2_125_3477_n771), .CI(DP_OP_423J2_125_3477_n765), .CO(
        DP_OP_423J2_125_3477_n728), .S(DP_OP_423J2_125_3477_n729) );
  FADDX1_HVT DP_OP_423J2_125_3477_U456 ( .A(DP_OP_423J2_125_3477_n777), .B(
        DP_OP_423J2_125_3477_n773), .CI(DP_OP_423J2_125_3477_n769), .CO(
        DP_OP_423J2_125_3477_n726), .S(DP_OP_423J2_125_3477_n727) );
  FADDX1_HVT DP_OP_423J2_125_3477_U455 ( .A(DP_OP_423J2_125_3477_n767), .B(
        DP_OP_423J2_125_3477_n761), .CI(DP_OP_423J2_125_3477_n763), .CO(
        DP_OP_423J2_125_3477_n724), .S(DP_OP_423J2_125_3477_n725) );
  FADDX1_HVT DP_OP_423J2_125_3477_U454 ( .A(DP_OP_423J2_125_3477_n942), .B(
        DP_OP_423J2_125_3477_n759), .CI(DP_OP_423J2_125_3477_n757), .CO(
        DP_OP_423J2_125_3477_n722), .S(DP_OP_423J2_125_3477_n723) );
  FADDX1_HVT DP_OP_423J2_125_3477_U453 ( .A(DP_OP_423J2_125_3477_n940), .B(
        DP_OP_423J2_125_3477_n755), .CI(DP_OP_423J2_125_3477_n753), .CO(
        DP_OP_423J2_125_3477_n720), .S(DP_OP_423J2_125_3477_n721) );
  FADDX1_HVT DP_OP_423J2_125_3477_U452 ( .A(DP_OP_423J2_125_3477_n751), .B(
        DP_OP_423J2_125_3477_n938), .CI(DP_OP_423J2_125_3477_n934), .CO(
        DP_OP_423J2_125_3477_n718), .S(DP_OP_423J2_125_3477_n719) );
  FADDX1_HVT DP_OP_423J2_125_3477_U451 ( .A(DP_OP_423J2_125_3477_n936), .B(
        DP_OP_423J2_125_3477_n932), .CI(DP_OP_423J2_125_3477_n749), .CO(
        DP_OP_423J2_125_3477_n716), .S(DP_OP_423J2_125_3477_n717) );
  FADDX1_HVT DP_OP_423J2_125_3477_U450 ( .A(DP_OP_423J2_125_3477_n930), .B(
        DP_OP_423J2_125_3477_n928), .CI(DP_OP_423J2_125_3477_n747), .CO(
        DP_OP_423J2_125_3477_n714), .S(DP_OP_423J2_125_3477_n715) );
  FADDX1_HVT DP_OP_423J2_125_3477_U449 ( .A(DP_OP_423J2_125_3477_n926), .B(
        DP_OP_423J2_125_3477_n745), .CI(DP_OP_423J2_125_3477_n920), .CO(
        DP_OP_423J2_125_3477_n712), .S(DP_OP_423J2_125_3477_n713) );
  FADDX1_HVT DP_OP_423J2_125_3477_U448 ( .A(DP_OP_423J2_125_3477_n924), .B(
        DP_OP_423J2_125_3477_n922), .CI(DP_OP_423J2_125_3477_n743), .CO(
        DP_OP_423J2_125_3477_n710), .S(DP_OP_423J2_125_3477_n711) );
  FADDX1_HVT DP_OP_423J2_125_3477_U447 ( .A(DP_OP_423J2_125_3477_n741), .B(
        DP_OP_423J2_125_3477_n918), .CI(DP_OP_423J2_125_3477_n739), .CO(
        DP_OP_423J2_125_3477_n708), .S(DP_OP_423J2_125_3477_n709) );
  FADDX1_HVT DP_OP_423J2_125_3477_U446 ( .A(DP_OP_423J2_125_3477_n737), .B(
        DP_OP_423J2_125_3477_n916), .CI(DP_OP_423J2_125_3477_n735), .CO(
        DP_OP_423J2_125_3477_n706), .S(DP_OP_423J2_125_3477_n707) );
  FADDX1_HVT DP_OP_423J2_125_3477_U445 ( .A(DP_OP_423J2_125_3477_n914), .B(
        DP_OP_423J2_125_3477_n912), .CI(DP_OP_423J2_125_3477_n727), .CO(
        DP_OP_423J2_125_3477_n704), .S(DP_OP_423J2_125_3477_n705) );
  FADDX1_HVT DP_OP_423J2_125_3477_U444 ( .A(DP_OP_423J2_125_3477_n731), .B(
        DP_OP_423J2_125_3477_n733), .CI(DP_OP_423J2_125_3477_n729), .CO(
        DP_OP_423J2_125_3477_n702), .S(DP_OP_423J2_125_3477_n703) );
  FADDX1_HVT DP_OP_423J2_125_3477_U443 ( .A(DP_OP_423J2_125_3477_n725), .B(
        DP_OP_423J2_125_3477_n910), .CI(DP_OP_423J2_125_3477_n723), .CO(
        DP_OP_423J2_125_3477_n700), .S(DP_OP_423J2_125_3477_n701) );
  FADDX1_HVT DP_OP_423J2_125_3477_U442 ( .A(DP_OP_423J2_125_3477_n908), .B(
        DP_OP_423J2_125_3477_n721), .CI(DP_OP_423J2_125_3477_n906), .CO(
        DP_OP_423J2_125_3477_n698), .S(DP_OP_423J2_125_3477_n699) );
  FADDX1_HVT DP_OP_423J2_125_3477_U441 ( .A(DP_OP_423J2_125_3477_n719), .B(
        DP_OP_423J2_125_3477_n904), .CI(DP_OP_423J2_125_3477_n902), .CO(
        DP_OP_423J2_125_3477_n696), .S(DP_OP_423J2_125_3477_n697) );
  FADDX1_HVT DP_OP_423J2_125_3477_U440 ( .A(DP_OP_423J2_125_3477_n717), .B(
        DP_OP_423J2_125_3477_n900), .CI(DP_OP_423J2_125_3477_n715), .CO(
        DP_OP_423J2_125_3477_n694), .S(DP_OP_423J2_125_3477_n695) );
  FADDX1_HVT DP_OP_423J2_125_3477_U439 ( .A(DP_OP_423J2_125_3477_n898), .B(
        DP_OP_423J2_125_3477_n711), .CI(DP_OP_423J2_125_3477_n896), .CO(
        DP_OP_423J2_125_3477_n692), .S(DP_OP_423J2_125_3477_n693) );
  FADDX1_HVT DP_OP_423J2_125_3477_U438 ( .A(DP_OP_423J2_125_3477_n713), .B(
        DP_OP_423J2_125_3477_n894), .CI(DP_OP_423J2_125_3477_n709), .CO(
        DP_OP_423J2_125_3477_n690), .S(DP_OP_423J2_125_3477_n691) );
  FADDX1_HVT DP_OP_423J2_125_3477_U437 ( .A(DP_OP_423J2_125_3477_n707), .B(
        DP_OP_423J2_125_3477_n892), .CI(DP_OP_423J2_125_3477_n705), .CO(
        DP_OP_423J2_125_3477_n688), .S(DP_OP_423J2_125_3477_n689) );
  FADDX1_HVT DP_OP_423J2_125_3477_U436 ( .A(DP_OP_423J2_125_3477_n703), .B(
        DP_OP_423J2_125_3477_n890), .CI(DP_OP_423J2_125_3477_n701), .CO(
        DP_OP_423J2_125_3477_n686), .S(DP_OP_423J2_125_3477_n687) );
  FADDX1_HVT DP_OP_423J2_125_3477_U435 ( .A(DP_OP_423J2_125_3477_n888), .B(
        DP_OP_423J2_125_3477_n699), .CI(DP_OP_423J2_125_3477_n886), .CO(
        DP_OP_423J2_125_3477_n684), .S(DP_OP_423J2_125_3477_n685) );
  FADDX1_HVT DP_OP_423J2_125_3477_U434 ( .A(DP_OP_423J2_125_3477_n697), .B(
        DP_OP_423J2_125_3477_n884), .CI(DP_OP_423J2_125_3477_n695), .CO(
        DP_OP_423J2_125_3477_n682), .S(DP_OP_423J2_125_3477_n683) );
  FADDX1_HVT DP_OP_423J2_125_3477_U433 ( .A(DP_OP_423J2_125_3477_n882), .B(
        DP_OP_423J2_125_3477_n693), .CI(DP_OP_423J2_125_3477_n880), .CO(
        DP_OP_423J2_125_3477_n680), .S(DP_OP_423J2_125_3477_n681) );
  FADDX1_HVT DP_OP_423J2_125_3477_U432 ( .A(DP_OP_423J2_125_3477_n691), .B(
        DP_OP_423J2_125_3477_n878), .CI(DP_OP_423J2_125_3477_n689), .CO(
        DP_OP_423J2_125_3477_n678), .S(DP_OP_423J2_125_3477_n679) );
  FADDX1_HVT DP_OP_423J2_125_3477_U431 ( .A(DP_OP_423J2_125_3477_n687), .B(
        DP_OP_423J2_125_3477_n876), .CI(DP_OP_423J2_125_3477_n685), .CO(
        DP_OP_423J2_125_3477_n676), .S(DP_OP_423J2_125_3477_n677) );
  FADDX1_HVT DP_OP_423J2_125_3477_U430 ( .A(DP_OP_423J2_125_3477_n874), .B(
        DP_OP_423J2_125_3477_n683), .CI(DP_OP_423J2_125_3477_n872), .CO(
        DP_OP_423J2_125_3477_n674), .S(DP_OP_423J2_125_3477_n675) );
  FADDX1_HVT DP_OP_423J2_125_3477_U429 ( .A(DP_OP_423J2_125_3477_n681), .B(
        DP_OP_423J2_125_3477_n870), .CI(DP_OP_423J2_125_3477_n679), .CO(
        DP_OP_423J2_125_3477_n672), .S(DP_OP_423J2_125_3477_n673) );
  FADDX1_HVT DP_OP_423J2_125_3477_U428 ( .A(DP_OP_423J2_125_3477_n677), .B(
        DP_OP_423J2_125_3477_n868), .CI(DP_OP_423J2_125_3477_n675), .CO(
        DP_OP_423J2_125_3477_n670), .S(DP_OP_423J2_125_3477_n671) );
  FADDX1_HVT DP_OP_423J2_125_3477_U427 ( .A(DP_OP_423J2_125_3477_n866), .B(
        DP_OP_423J2_125_3477_n673), .CI(DP_OP_423J2_125_3477_n671), .CO(
        DP_OP_423J2_125_3477_n668), .S(DP_OP_423J2_125_3477_n669) );
  FADDX1_HVT DP_OP_423J2_125_3477_U425 ( .A(DP_OP_423J2_125_3477_n1995), .B(
        DP_OP_423J2_125_3477_n2141), .CI(DP_OP_423J2_125_3477_n1951), .CO(
        DP_OP_423J2_125_3477_n664), .S(DP_OP_423J2_125_3477_n665) );
  FADDX1_HVT DP_OP_423J2_125_3477_U424 ( .A(DP_OP_423J2_125_3477_n2347), .B(
        DP_OP_423J2_125_3477_n2405), .CI(DP_OP_423J2_125_3477_n2740), .CO(
        DP_OP_423J2_125_3477_n662), .S(DP_OP_423J2_125_3477_n663) );
  FADDX1_HVT DP_OP_423J2_125_3477_U423 ( .A(DP_OP_423J2_125_3477_n2303), .B(
        DP_OP_423J2_125_3477_n2567), .CI(DP_OP_423J2_125_3477_n2435), .CO(
        DP_OP_423J2_125_3477_n660), .S(DP_OP_423J2_125_3477_n661) );
  FADDX1_HVT DP_OP_423J2_125_3477_U422 ( .A(DP_OP_423J2_125_3477_n2127), .B(
        DP_OP_423J2_125_3477_n2523), .CI(DP_OP_423J2_125_3477_n2039), .CO(
        DP_OP_423J2_125_3477_n658), .S(DP_OP_423J2_125_3477_n659) );
  FADDX1_HVT DP_OP_423J2_125_3477_U421 ( .A(DP_OP_423J2_125_3477_n1863), .B(
        DP_OP_423J2_125_3477_n1907), .CI(DP_OP_423J2_125_3477_n2479), .CO(
        DP_OP_423J2_125_3477_n656), .S(DP_OP_423J2_125_3477_n657) );
  FADDX1_HVT DP_OP_423J2_125_3477_U420 ( .A(DP_OP_423J2_125_3477_n2083), .B(
        DP_OP_423J2_125_3477_n2872), .CI(DP_OP_423J2_125_3477_n2171), .CO(
        DP_OP_423J2_125_3477_n654), .S(DP_OP_423J2_125_3477_n655) );
  FADDX1_HVT DP_OP_423J2_125_3477_U419 ( .A(DP_OP_423J2_125_3477_n2784), .B(
        DP_OP_423J2_125_3477_n2053), .CI(DP_OP_423J2_125_3477_n1819), .CO(
        DP_OP_423J2_125_3477_n652), .S(DP_OP_423J2_125_3477_n653) );
  FADDX1_HVT DP_OP_423J2_125_3477_U418 ( .A(DP_OP_423J2_125_3477_n2611), .B(
        DP_OP_423J2_125_3477_n2493), .CI(DP_OP_423J2_125_3477_n2317), .CO(
        DP_OP_423J2_125_3477_n650), .S(DP_OP_423J2_125_3477_n651) );
  FADDX1_HVT DP_OP_423J2_125_3477_U417 ( .A(DP_OP_423J2_125_3477_n2828), .B(
        DP_OP_423J2_125_3477_n1833), .CI(DP_OP_423J2_125_3477_n2581), .CO(
        DP_OP_423J2_125_3477_n648), .S(DP_OP_423J2_125_3477_n649) );
  FADDX1_HVT DP_OP_423J2_125_3477_U416 ( .A(DP_OP_423J2_125_3477_n2655), .B(
        DP_OP_423J2_125_3477_n2259), .CI(DP_OP_423J2_125_3477_n2625), .CO(
        DP_OP_423J2_125_3477_n646), .S(DP_OP_423J2_125_3477_n647) );
  FADDX1_HVT DP_OP_423J2_125_3477_U415 ( .A(DP_OP_423J2_125_3477_n1775), .B(
        DP_OP_423J2_125_3477_n2391), .CI(DP_OP_423J2_125_3477_n2886), .CO(
        DP_OP_423J2_125_3477_n644), .S(DP_OP_423J2_125_3477_n645) );
  FADDX1_HVT DP_OP_423J2_125_3477_U414 ( .A(DP_OP_423J2_125_3477_n2879), .B(
        DP_OP_423J2_125_3477_n2530), .CI(DP_OP_423J2_125_3477_n2798), .CO(
        DP_OP_423J2_125_3477_n642), .S(DP_OP_423J2_125_3477_n643) );
  FADDX1_HVT DP_OP_423J2_125_3477_U413 ( .A(DP_OP_423J2_125_3477_n2835), .B(
        DP_OP_423J2_125_3477_n1958), .CI(DP_OP_423J2_125_3477_n2273), .CO(
        DP_OP_423J2_125_3477_n640), .S(DP_OP_423J2_125_3477_n641) );
  FADDX1_HVT DP_OP_423J2_125_3477_U412 ( .A(DP_OP_423J2_125_3477_n2747), .B(
        DP_OP_423J2_125_3477_n2097), .CI(DP_OP_423J2_125_3477_n1921), .CO(
        DP_OP_423J2_125_3477_n638), .S(DP_OP_423J2_125_3477_n639) );
  FADDX1_HVT DP_OP_423J2_125_3477_U411 ( .A(DP_OP_423J2_125_3477_n667), .B(
        DP_OP_423J2_125_3477_n2449), .CI(DP_OP_423J2_125_3477_n2266), .CO(
        DP_OP_423J2_125_3477_n636), .S(DP_OP_423J2_125_3477_n637) );
  FADDX1_HVT DP_OP_423J2_125_3477_U410 ( .A(DP_OP_423J2_125_3477_n2215), .B(
        DP_OP_423J2_125_3477_n1877), .CI(DP_OP_423J2_125_3477_n2710), .CO(
        DP_OP_423J2_125_3477_n634), .S(DP_OP_423J2_125_3477_n635) );
  FADDX1_HVT DP_OP_423J2_125_3477_U409 ( .A(DP_OP_423J2_125_3477_n2669), .B(
        DP_OP_423J2_125_3477_n2442), .CI(DP_OP_423J2_125_3477_n2754), .CO(
        DP_OP_423J2_125_3477_n632), .S(DP_OP_423J2_125_3477_n633) );
  FADDX1_HVT DP_OP_423J2_125_3477_U408 ( .A(DP_OP_423J2_125_3477_n2090), .B(
        DP_OP_423J2_125_3477_n2009), .CI(DP_OP_423J2_125_3477_n1965), .CO(
        DP_OP_423J2_125_3477_n630), .S(DP_OP_423J2_125_3477_n631) );
  FADDX1_HVT DP_OP_423J2_125_3477_U407 ( .A(DP_OP_423J2_125_3477_n2222), .B(
        DP_OP_423J2_125_3477_n2842), .CI(DP_OP_423J2_125_3477_n2354), .CO(
        DP_OP_423J2_125_3477_n628), .S(DP_OP_423J2_125_3477_n629) );
  FADDX1_HVT DP_OP_423J2_125_3477_U406 ( .A(DP_OP_423J2_125_3477_n2537), .B(
        DP_OP_423J2_125_3477_n2229), .CI(DP_OP_423J2_125_3477_n2662), .CO(
        DP_OP_423J2_125_3477_n626), .S(DP_OP_423J2_125_3477_n627) );
  FADDX1_HVT DP_OP_423J2_125_3477_U405 ( .A(DP_OP_423J2_125_3477_n2134), .B(
        DP_OP_423J2_125_3477_n2486), .CI(DP_OP_423J2_125_3477_n2398), .CO(
        DP_OP_423J2_125_3477_n624), .S(DP_OP_423J2_125_3477_n625) );
  FADDX1_HVT DP_OP_423J2_125_3477_U404 ( .A(DP_OP_423J2_125_3477_n2361), .B(
        DP_OP_423J2_125_3477_n2574), .CI(DP_OP_423J2_125_3477_n2310), .CO(
        DP_OP_423J2_125_3477_n622), .S(DP_OP_423J2_125_3477_n623) );
  FADDX1_HVT DP_OP_423J2_125_3477_U403 ( .A(DP_OP_423J2_125_3477_n2185), .B(
        DP_OP_423J2_125_3477_n2703), .CI(DP_OP_423J2_125_3477_n2046), .CO(
        DP_OP_423J2_125_3477_n620), .S(DP_OP_423J2_125_3477_n621) );
  FADDX1_HVT DP_OP_423J2_125_3477_U402 ( .A(DP_OP_423J2_125_3477_n2002), .B(
        DP_OP_423J2_125_3477_n2178), .CI(DP_OP_423J2_125_3477_n1826), .CO(
        DP_OP_423J2_125_3477_n618), .S(DP_OP_423J2_125_3477_n619) );
  FADDX1_HVT DP_OP_423J2_125_3477_U401 ( .A(DP_OP_423J2_125_3477_n1870), .B(
        DP_OP_423J2_125_3477_n2618), .CI(DP_OP_423J2_125_3477_n1914), .CO(
        DP_OP_423J2_125_3477_n616), .S(DP_OP_423J2_125_3477_n617) );
  FADDX1_HVT DP_OP_423J2_125_3477_U400 ( .A(DP_OP_423J2_125_3477_n2791), .B(
        DP_OP_423J2_125_3477_n862), .CI(DP_OP_423J2_125_3477_n860), .CO(
        DP_OP_423J2_125_3477_n614), .S(DP_OP_423J2_125_3477_n615) );
  FADDX1_HVT DP_OP_423J2_125_3477_U399 ( .A(DP_OP_423J2_125_3477_n858), .B(
        DP_OP_423J2_125_3477_n838), .CI(DP_OP_423J2_125_3477_n836), .CO(
        DP_OP_423J2_125_3477_n612), .S(DP_OP_423J2_125_3477_n613) );
  FADDX1_HVT DP_OP_423J2_125_3477_U398 ( .A(DP_OP_423J2_125_3477_n856), .B(
        DP_OP_423J2_125_3477_n842), .CI(DP_OP_423J2_125_3477_n840), .CO(
        DP_OP_423J2_125_3477_n610), .S(DP_OP_423J2_125_3477_n611) );
  FADDX1_HVT DP_OP_423J2_125_3477_U397 ( .A(DP_OP_423J2_125_3477_n854), .B(
        DP_OP_423J2_125_3477_n844), .CI(DP_OP_423J2_125_3477_n846), .CO(
        DP_OP_423J2_125_3477_n608), .S(DP_OP_423J2_125_3477_n609) );
  FADDX1_HVT DP_OP_423J2_125_3477_U396 ( .A(DP_OP_423J2_125_3477_n852), .B(
        DP_OP_423J2_125_3477_n848), .CI(DP_OP_423J2_125_3477_n850), .CO(
        DP_OP_423J2_125_3477_n606), .S(DP_OP_423J2_125_3477_n607) );
  FADDX1_HVT DP_OP_423J2_125_3477_U395 ( .A(DP_OP_423J2_125_3477_n834), .B(
        DP_OP_423J2_125_3477_n822), .CI(DP_OP_423J2_125_3477_n820), .CO(
        DP_OP_423J2_125_3477_n604), .S(DP_OP_423J2_125_3477_n605) );
  FADDX1_HVT DP_OP_423J2_125_3477_U394 ( .A(DP_OP_423J2_125_3477_n832), .B(
        DP_OP_423J2_125_3477_n824), .CI(DP_OP_423J2_125_3477_n826), .CO(
        DP_OP_423J2_125_3477_n602), .S(DP_OP_423J2_125_3477_n603) );
  FADDX1_HVT DP_OP_423J2_125_3477_U393 ( .A(DP_OP_423J2_125_3477_n830), .B(
        DP_OP_423J2_125_3477_n828), .CI(DP_OP_423J2_125_3477_n818), .CO(
        DP_OP_423J2_125_3477_n600), .S(DP_OP_423J2_125_3477_n601) );
  FADDX1_HVT DP_OP_423J2_125_3477_U392 ( .A(DP_OP_423J2_125_3477_n816), .B(
        DP_OP_423J2_125_3477_n810), .CI(DP_OP_423J2_125_3477_n796), .CO(
        DP_OP_423J2_125_3477_n598), .S(DP_OP_423J2_125_3477_n599) );
  FADDX1_HVT DP_OP_423J2_125_3477_U391 ( .A(DP_OP_423J2_125_3477_n814), .B(
        DP_OP_423J2_125_3477_n651), .CI(DP_OP_423J2_125_3477_n798), .CO(
        DP_OP_423J2_125_3477_n596), .S(DP_OP_423J2_125_3477_n597) );
  FADDX1_HVT DP_OP_423J2_125_3477_U390 ( .A(DP_OP_423J2_125_3477_n812), .B(
        DP_OP_423J2_125_3477_n657), .CI(DP_OP_423J2_125_3477_n802), .CO(
        DP_OP_423J2_125_3477_n594), .S(DP_OP_423J2_125_3477_n595) );
  FADDX1_HVT DP_OP_423J2_125_3477_U389 ( .A(DP_OP_423J2_125_3477_n665), .B(
        DP_OP_423J2_125_3477_n806), .CI(DP_OP_423J2_125_3477_n800), .CO(
        DP_OP_423J2_125_3477_n592), .S(DP_OP_423J2_125_3477_n593) );
  FADDX1_HVT DP_OP_423J2_125_3477_U388 ( .A(DP_OP_423J2_125_3477_n655), .B(
        DP_OP_423J2_125_3477_n808), .CI(DP_OP_423J2_125_3477_n804), .CO(
        DP_OP_423J2_125_3477_n590), .S(DP_OP_423J2_125_3477_n591) );
  FADDX1_HVT DP_OP_423J2_125_3477_U387 ( .A(DP_OP_423J2_125_3477_n653), .B(
        DP_OP_423J2_125_3477_n663), .CI(DP_OP_423J2_125_3477_n661), .CO(
        DP_OP_423J2_125_3477_n588), .S(DP_OP_423J2_125_3477_n589) );
  FADDX1_HVT DP_OP_423J2_125_3477_U386 ( .A(DP_OP_423J2_125_3477_n647), .B(
        DP_OP_423J2_125_3477_n659), .CI(DP_OP_423J2_125_3477_n649), .CO(
        DP_OP_423J2_125_3477_n586), .S(DP_OP_423J2_125_3477_n587) );
  FADDX1_HVT DP_OP_423J2_125_3477_U385 ( .A(DP_OP_423J2_125_3477_n645), .B(
        DP_OP_423J2_125_3477_n633), .CI(DP_OP_423J2_125_3477_n627), .CO(
        DP_OP_423J2_125_3477_n584), .S(DP_OP_423J2_125_3477_n585) );
  FADDX1_HVT DP_OP_423J2_125_3477_U384 ( .A(DP_OP_423J2_125_3477_n643), .B(
        DP_OP_423J2_125_3477_n635), .CI(DP_OP_423J2_125_3477_n629), .CO(
        DP_OP_423J2_125_3477_n582), .S(DP_OP_423J2_125_3477_n583) );
  FADDX1_HVT DP_OP_423J2_125_3477_U383 ( .A(DP_OP_423J2_125_3477_n641), .B(
        DP_OP_423J2_125_3477_n637), .CI(DP_OP_423J2_125_3477_n631), .CO(
        DP_OP_423J2_125_3477_n580), .S(DP_OP_423J2_125_3477_n581) );
  FADDX1_HVT DP_OP_423J2_125_3477_U382 ( .A(DP_OP_423J2_125_3477_n639), .B(
        DP_OP_423J2_125_3477_n625), .CI(DP_OP_423J2_125_3477_n623), .CO(
        DP_OP_423J2_125_3477_n578), .S(DP_OP_423J2_125_3477_n579) );
  FADDX1_HVT DP_OP_423J2_125_3477_U381 ( .A(DP_OP_423J2_125_3477_n621), .B(
        DP_OP_423J2_125_3477_n619), .CI(DP_OP_423J2_125_3477_n617), .CO(
        DP_OP_423J2_125_3477_n576), .S(DP_OP_423J2_125_3477_n577) );
  FADDX1_HVT DP_OP_423J2_125_3477_U380 ( .A(DP_OP_423J2_125_3477_n794), .B(
        DP_OP_423J2_125_3477_n792), .CI(DP_OP_423J2_125_3477_n790), .CO(
        DP_OP_423J2_125_3477_n574), .S(DP_OP_423J2_125_3477_n575) );
  FADDX1_HVT DP_OP_423J2_125_3477_U379 ( .A(DP_OP_423J2_125_3477_n788), .B(
        DP_OP_423J2_125_3477_n784), .CI(DP_OP_423J2_125_3477_n782), .CO(
        DP_OP_423J2_125_3477_n572), .S(DP_OP_423J2_125_3477_n573) );
  FADDX1_HVT DP_OP_423J2_125_3477_U378 ( .A(DP_OP_423J2_125_3477_n786), .B(
        DP_OP_423J2_125_3477_n780), .CI(DP_OP_423J2_125_3477_n778), .CO(
        DP_OP_423J2_125_3477_n570), .S(DP_OP_423J2_125_3477_n571) );
  FADDX1_HVT DP_OP_423J2_125_3477_U377 ( .A(DP_OP_423J2_125_3477_n615), .B(
        DP_OP_423J2_125_3477_n776), .CI(DP_OP_423J2_125_3477_n607), .CO(
        DP_OP_423J2_125_3477_n568), .S(DP_OP_423J2_125_3477_n569) );
  FADDX1_HVT DP_OP_423J2_125_3477_U376 ( .A(DP_OP_423J2_125_3477_n774), .B(
        DP_OP_423J2_125_3477_n613), .CI(DP_OP_423J2_125_3477_n611), .CO(
        DP_OP_423J2_125_3477_n566), .S(DP_OP_423J2_125_3477_n567) );
  FADDX1_HVT DP_OP_423J2_125_3477_U375 ( .A(DP_OP_423J2_125_3477_n772), .B(
        DP_OP_423J2_125_3477_n609), .CI(DP_OP_423J2_125_3477_n764), .CO(
        DP_OP_423J2_125_3477_n564), .S(DP_OP_423J2_125_3477_n565) );
  FADDX1_HVT DP_OP_423J2_125_3477_U374 ( .A(DP_OP_423J2_125_3477_n770), .B(
        DP_OP_423J2_125_3477_n766), .CI(DP_OP_423J2_125_3477_n768), .CO(
        DP_OP_423J2_125_3477_n562), .S(DP_OP_423J2_125_3477_n563) );
  FADDX1_HVT DP_OP_423J2_125_3477_U373 ( .A(DP_OP_423J2_125_3477_n605), .B(
        DP_OP_423J2_125_3477_n601), .CI(DP_OP_423J2_125_3477_n758), .CO(
        DP_OP_423J2_125_3477_n560), .S(DP_OP_423J2_125_3477_n561) );
  FADDX1_HVT DP_OP_423J2_125_3477_U372 ( .A(DP_OP_423J2_125_3477_n762), .B(
        DP_OP_423J2_125_3477_n603), .CI(DP_OP_423J2_125_3477_n760), .CO(
        DP_OP_423J2_125_3477_n558), .S(DP_OP_423J2_125_3477_n559) );
  FADDX1_HVT DP_OP_423J2_125_3477_U371 ( .A(DP_OP_423J2_125_3477_n599), .B(
        DP_OP_423J2_125_3477_n754), .CI(DP_OP_423J2_125_3477_n752), .CO(
        DP_OP_423J2_125_3477_n556), .S(DP_OP_423J2_125_3477_n557) );
  FADDX1_HVT DP_OP_423J2_125_3477_U370 ( .A(DP_OP_423J2_125_3477_n756), .B(
        DP_OP_423J2_125_3477_n591), .CI(DP_OP_423J2_125_3477_n750), .CO(
        DP_OP_423J2_125_3477_n554), .S(DP_OP_423J2_125_3477_n555) );
  FADDX1_HVT DP_OP_423J2_125_3477_U369 ( .A(DP_OP_423J2_125_3477_n597), .B(
        DP_OP_423J2_125_3477_n589), .CI(DP_OP_423J2_125_3477_n587), .CO(
        DP_OP_423J2_125_3477_n552), .S(DP_OP_423J2_125_3477_n553) );
  FADDX1_HVT DP_OP_423J2_125_3477_U368 ( .A(DP_OP_423J2_125_3477_n595), .B(
        DP_OP_423J2_125_3477_n593), .CI(DP_OP_423J2_125_3477_n585), .CO(
        DP_OP_423J2_125_3477_n550), .S(DP_OP_423J2_125_3477_n551) );
  FADDX1_HVT DP_OP_423J2_125_3477_U367 ( .A(DP_OP_423J2_125_3477_n581), .B(
        DP_OP_423J2_125_3477_n583), .CI(DP_OP_423J2_125_3477_n748), .CO(
        DP_OP_423J2_125_3477_n548), .S(DP_OP_423J2_125_3477_n549) );
  FADDX1_HVT DP_OP_423J2_125_3477_U366 ( .A(DP_OP_423J2_125_3477_n579), .B(
        DP_OP_423J2_125_3477_n746), .CI(DP_OP_423J2_125_3477_n577), .CO(
        DP_OP_423J2_125_3477_n546), .S(DP_OP_423J2_125_3477_n547) );
  FADDX1_HVT DP_OP_423J2_125_3477_U365 ( .A(DP_OP_423J2_125_3477_n744), .B(
        DP_OP_423J2_125_3477_n742), .CI(DP_OP_423J2_125_3477_n575), .CO(
        DP_OP_423J2_125_3477_n544), .S(DP_OP_423J2_125_3477_n545) );
  FADDX1_HVT DP_OP_423J2_125_3477_U364 ( .A(DP_OP_423J2_125_3477_n740), .B(
        DP_OP_423J2_125_3477_n738), .CI(DP_OP_423J2_125_3477_n736), .CO(
        DP_OP_423J2_125_3477_n542), .S(DP_OP_423J2_125_3477_n543) );
  FADDX1_HVT DP_OP_423J2_125_3477_U363 ( .A(DP_OP_423J2_125_3477_n734), .B(
        DP_OP_423J2_125_3477_n573), .CI(DP_OP_423J2_125_3477_n571), .CO(
        DP_OP_423J2_125_3477_n540), .S(DP_OP_423J2_125_3477_n541) );
  FADDX1_HVT DP_OP_423J2_125_3477_U362 ( .A(DP_OP_423J2_125_3477_n732), .B(
        DP_OP_423J2_125_3477_n569), .CI(DP_OP_423J2_125_3477_n563), .CO(
        DP_OP_423J2_125_3477_n538), .S(DP_OP_423J2_125_3477_n539) );
  FADDX1_HVT DP_OP_423J2_125_3477_U361 ( .A(DP_OP_423J2_125_3477_n730), .B(
        DP_OP_423J2_125_3477_n728), .CI(DP_OP_423J2_125_3477_n565), .CO(
        DP_OP_423J2_125_3477_n536), .S(DP_OP_423J2_125_3477_n537) );
  FADDX1_HVT DP_OP_423J2_125_3477_U360 ( .A(DP_OP_423J2_125_3477_n726), .B(
        DP_OP_423J2_125_3477_n567), .CI(DP_OP_423J2_125_3477_n724), .CO(
        DP_OP_423J2_125_3477_n534), .S(DP_OP_423J2_125_3477_n535) );
  FADDX1_HVT DP_OP_423J2_125_3477_U359 ( .A(DP_OP_423J2_125_3477_n561), .B(
        DP_OP_423J2_125_3477_n559), .CI(DP_OP_423J2_125_3477_n722), .CO(
        DP_OP_423J2_125_3477_n532), .S(DP_OP_423J2_125_3477_n533) );
  FADDX1_HVT DP_OP_423J2_125_3477_U358 ( .A(DP_OP_423J2_125_3477_n557), .B(
        DP_OP_423J2_125_3477_n720), .CI(DP_OP_423J2_125_3477_n718), .CO(
        DP_OP_423J2_125_3477_n530), .S(DP_OP_423J2_125_3477_n531) );
  FADDX1_HVT DP_OP_423J2_125_3477_U357 ( .A(DP_OP_423J2_125_3477_n553), .B(
        DP_OP_423J2_125_3477_n555), .CI(DP_OP_423J2_125_3477_n551), .CO(
        DP_OP_423J2_125_3477_n528), .S(DP_OP_423J2_125_3477_n529) );
  FADDX1_HVT DP_OP_423J2_125_3477_U356 ( .A(DP_OP_423J2_125_3477_n549), .B(
        DP_OP_423J2_125_3477_n716), .CI(DP_OP_423J2_125_3477_n547), .CO(
        DP_OP_423J2_125_3477_n526), .S(DP_OP_423J2_125_3477_n527) );
  FADDX1_HVT DP_OP_423J2_125_3477_U355 ( .A(DP_OP_423J2_125_3477_n714), .B(
        DP_OP_423J2_125_3477_n712), .CI(DP_OP_423J2_125_3477_n710), .CO(
        DP_OP_423J2_125_3477_n524), .S(DP_OP_423J2_125_3477_n525) );
  FADDX1_HVT DP_OP_423J2_125_3477_U354 ( .A(DP_OP_423J2_125_3477_n545), .B(
        DP_OP_423J2_125_3477_n708), .CI(DP_OP_423J2_125_3477_n543), .CO(
        DP_OP_423J2_125_3477_n522), .S(DP_OP_423J2_125_3477_n523) );
  FADDX1_HVT DP_OP_423J2_125_3477_U353 ( .A(DP_OP_423J2_125_3477_n706), .B(
        DP_OP_423J2_125_3477_n541), .CI(DP_OP_423J2_125_3477_n704), .CO(
        DP_OP_423J2_125_3477_n520), .S(DP_OP_423J2_125_3477_n521) );
  FADDX1_HVT DP_OP_423J2_125_3477_U352 ( .A(DP_OP_423J2_125_3477_n539), .B(
        DP_OP_423J2_125_3477_n537), .CI(DP_OP_423J2_125_3477_n535), .CO(
        DP_OP_423J2_125_3477_n518), .S(DP_OP_423J2_125_3477_n519) );
  FADDX1_HVT DP_OP_423J2_125_3477_U351 ( .A(DP_OP_423J2_125_3477_n702), .B(
        DP_OP_423J2_125_3477_n700), .CI(DP_OP_423J2_125_3477_n533), .CO(
        DP_OP_423J2_125_3477_n516), .S(DP_OP_423J2_125_3477_n517) );
  FADDX1_HVT DP_OP_423J2_125_3477_U350 ( .A(DP_OP_423J2_125_3477_n698), .B(
        DP_OP_423J2_125_3477_n531), .CI(DP_OP_423J2_125_3477_n529), .CO(
        DP_OP_423J2_125_3477_n514), .S(DP_OP_423J2_125_3477_n515) );
  FADDX1_HVT DP_OP_423J2_125_3477_U349 ( .A(DP_OP_423J2_125_3477_n696), .B(
        DP_OP_423J2_125_3477_n527), .CI(DP_OP_423J2_125_3477_n694), .CO(
        DP_OP_423J2_125_3477_n512), .S(DP_OP_423J2_125_3477_n513) );
  FADDX1_HVT DP_OP_423J2_125_3477_U348 ( .A(DP_OP_423J2_125_3477_n692), .B(
        DP_OP_423J2_125_3477_n525), .CI(DP_OP_423J2_125_3477_n690), .CO(
        DP_OP_423J2_125_3477_n510), .S(DP_OP_423J2_125_3477_n511) );
  FADDX1_HVT DP_OP_423J2_125_3477_U347 ( .A(DP_OP_423J2_125_3477_n523), .B(
        DP_OP_423J2_125_3477_n688), .CI(DP_OP_423J2_125_3477_n521), .CO(
        DP_OP_423J2_125_3477_n508), .S(DP_OP_423J2_125_3477_n509) );
  FADDX1_HVT DP_OP_423J2_125_3477_U346 ( .A(DP_OP_423J2_125_3477_n519), .B(
        DP_OP_423J2_125_3477_n686), .CI(DP_OP_423J2_125_3477_n517), .CO(
        DP_OP_423J2_125_3477_n506), .S(DP_OP_423J2_125_3477_n507) );
  FADDX1_HVT DP_OP_423J2_125_3477_U345 ( .A(DP_OP_423J2_125_3477_n684), .B(
        DP_OP_423J2_125_3477_n515), .CI(DP_OP_423J2_125_3477_n682), .CO(
        DP_OP_423J2_125_3477_n504), .S(DP_OP_423J2_125_3477_n505) );
  FADDX1_HVT DP_OP_423J2_125_3477_U344 ( .A(DP_OP_423J2_125_3477_n513), .B(
        DP_OP_423J2_125_3477_n680), .CI(DP_OP_423J2_125_3477_n511), .CO(
        DP_OP_423J2_125_3477_n502), .S(DP_OP_423J2_125_3477_n503) );
  FADDX1_HVT DP_OP_423J2_125_3477_U343 ( .A(DP_OP_423J2_125_3477_n678), .B(
        DP_OP_423J2_125_3477_n509), .CI(DP_OP_423J2_125_3477_n507), .CO(
        DP_OP_423J2_125_3477_n500), .S(DP_OP_423J2_125_3477_n501) );
  FADDX1_HVT DP_OP_423J2_125_3477_U342 ( .A(DP_OP_423J2_125_3477_n676), .B(
        DP_OP_423J2_125_3477_n505), .CI(DP_OP_423J2_125_3477_n674), .CO(
        DP_OP_423J2_125_3477_n498), .S(DP_OP_423J2_125_3477_n499) );
  FADDX1_HVT DP_OP_423J2_125_3477_U341 ( .A(DP_OP_423J2_125_3477_n503), .B(
        DP_OP_423J2_125_3477_n672), .CI(DP_OP_423J2_125_3477_n501), .CO(
        DP_OP_423J2_125_3477_n496), .S(DP_OP_423J2_125_3477_n497) );
  FADDX1_HVT DP_OP_423J2_125_3477_U340 ( .A(DP_OP_423J2_125_3477_n670), .B(
        DP_OP_423J2_125_3477_n499), .CI(DP_OP_423J2_125_3477_n497), .CO(
        DP_OP_423J2_125_3477_n494), .S(DP_OP_423J2_125_3477_n495) );
  FADDX1_HVT DP_OP_423J2_125_3477_U339 ( .A(DP_OP_423J2_125_3477_n666), .B(
        DP_OP_423J2_125_3477_n2529), .CI(DP_OP_423J2_125_3477_n2221), .CO(
        DP_OP_423J2_125_3477_n492), .S(DP_OP_423J2_125_3477_n493) );
  FADDX1_HVT DP_OP_423J2_125_3477_U338 ( .A(DP_OP_423J2_125_3477_n1994), .B(
        DP_OP_423J2_125_3477_n1957), .CI(DP_OP_423J2_125_3477_n2441), .CO(
        DP_OP_423J2_125_3477_n490), .S(DP_OP_423J2_125_3477_n491) );
  FADDX1_HVT DP_OP_423J2_125_3477_U337 ( .A(DP_OP_423J2_125_3477_n2697), .B(
        DP_OP_423J2_125_3477_n2170), .CI(DP_OP_423J2_125_3477_n2089), .CO(
        DP_OP_423J2_125_3477_n488), .S(DP_OP_423J2_125_3477_n489) );
  FADDX1_HVT DP_OP_423J2_125_3477_U336 ( .A(DP_OP_423J2_125_3477_n2082), .B(
        DP_OP_423J2_125_3477_n1906), .CI(DP_OP_423J2_125_3477_n2739), .CO(
        DP_OP_423J2_125_3477_n486), .S(DP_OP_423J2_125_3477_n487) );
  FADDX1_HVT DP_OP_423J2_125_3477_U335 ( .A(DP_OP_423J2_125_3477_n1862), .B(
        DP_OP_423J2_125_3477_n2478), .CI(DP_OP_423J2_125_3477_n1950), .CO(
        DP_OP_423J2_125_3477_n484), .S(DP_OP_423J2_125_3477_n485) );
  FADDX1_HVT DP_OP_423J2_125_3477_U334 ( .A(DP_OP_423J2_125_3477_n2783), .B(
        DP_OP_423J2_125_3477_n2434), .CI(DP_OP_423J2_125_3477_n2038), .CO(
        DP_OP_423J2_125_3477_n482), .S(DP_OP_423J2_125_3477_n483) );
  FADDX1_HVT DP_OP_423J2_125_3477_U333 ( .A(DP_OP_423J2_125_3477_n2126), .B(
        DP_OP_423J2_125_3477_n2566), .CI(DP_OP_423J2_125_3477_n2522), .CO(
        DP_OP_423J2_125_3477_n480), .S(DP_OP_423J2_125_3477_n481) );
  FADDX1_HVT DP_OP_423J2_125_3477_U332 ( .A(DP_OP_423J2_125_3477_n2346), .B(
        DP_OP_423J2_125_3477_n1818), .CI(DP_OP_423J2_125_3477_n2871), .CO(
        DP_OP_423J2_125_3477_n478), .S(DP_OP_423J2_125_3477_n479) );
  FADDX1_HVT DP_OP_423J2_125_3477_U331 ( .A(DP_OP_423J2_125_3477_n2827), .B(
        DP_OP_423J2_125_3477_n2878), .CI(DP_OP_423J2_125_3477_n2746), .CO(
        DP_OP_423J2_125_3477_n476), .S(DP_OP_423J2_125_3477_n477) );
  FADDX1_HVT DP_OP_423J2_125_3477_U330 ( .A(DP_OP_423J2_125_3477_n2610), .B(
        DP_OP_423J2_125_3477_n2258), .CI(DP_OP_423J2_125_3477_n2834), .CO(
        DP_OP_423J2_125_3477_n474), .S(DP_OP_423J2_125_3477_n475) );
  FADDX1_HVT DP_OP_423J2_125_3477_U329 ( .A(DP_OP_423J2_125_3477_n2654), .B(
        DP_OP_423J2_125_3477_n2302), .CI(DP_OP_423J2_125_3477_n2133), .CO(
        DP_OP_423J2_125_3477_n472), .S(DP_OP_423J2_125_3477_n473) );
  FADDX1_HVT DP_OP_423J2_125_3477_U328 ( .A(DP_OP_423J2_125_3477_n2265), .B(
        DP_OP_423J2_125_3477_n2390), .CI(DP_OP_423J2_125_3477_n2397), .CO(
        DP_OP_423J2_125_3477_n470), .S(DP_OP_423J2_125_3477_n471) );
  FADDX1_HVT DP_OP_423J2_125_3477_U327 ( .A(DP_OP_423J2_125_3477_n1774), .B(
        DP_OP_423J2_125_3477_n2353), .CI(DP_OP_423J2_125_3477_n2309), .CO(
        DP_OP_423J2_125_3477_n468), .S(DP_OP_423J2_125_3477_n469) );
  FADDX1_HVT DP_OP_423J2_125_3477_U326 ( .A(DP_OP_423J2_125_3477_n2214), .B(
        DP_OP_423J2_125_3477_n2485), .CI(DP_OP_423J2_125_3477_n2001), .CO(
        DP_OP_423J2_125_3477_n466), .S(DP_OP_423J2_125_3477_n467) );
  FADDX1_HVT DP_OP_423J2_125_3477_U325 ( .A(DP_OP_423J2_125_3477_n2573), .B(
        DP_OP_423J2_125_3477_n2661), .CI(DP_OP_423J2_125_3477_n2045), .CO(
        DP_OP_423J2_125_3477_n464), .S(DP_OP_423J2_125_3477_n465) );
  FADDX1_HVT DP_OP_423J2_125_3477_U324 ( .A(DP_OP_423J2_125_3477_n2702), .B(
        DP_OP_423J2_125_3477_n1869), .CI(DP_OP_423J2_125_3477_n1825), .CO(
        DP_OP_423J2_125_3477_n462), .S(DP_OP_423J2_125_3477_n463) );
  FADDX1_HVT DP_OP_423J2_125_3477_U323 ( .A(DP_OP_423J2_125_3477_n2790), .B(
        DP_OP_423J2_125_3477_n1913), .CI(DP_OP_423J2_125_3477_n2177), .CO(
        DP_OP_423J2_125_3477_n460), .S(DP_OP_423J2_125_3477_n461) );
  FADDX1_HVT DP_OP_423J2_125_3477_U322 ( .A(DP_OP_423J2_125_3477_n2617), .B(
        DP_OP_423J2_125_3477_n664), .CI(DP_OP_423J2_125_3477_n662), .CO(
        DP_OP_423J2_125_3477_n458), .S(DP_OP_423J2_125_3477_n459) );
  FADDX1_HVT DP_OP_423J2_125_3477_U321 ( .A(DP_OP_423J2_125_3477_n660), .B(
        DP_OP_423J2_125_3477_n646), .CI(DP_OP_423J2_125_3477_n648), .CO(
        DP_OP_423J2_125_3477_n456), .S(DP_OP_423J2_125_3477_n457) );
  FADDX1_HVT DP_OP_423J2_125_3477_U320 ( .A(DP_OP_423J2_125_3477_n658), .B(
        DP_OP_423J2_125_3477_n650), .CI(DP_OP_423J2_125_3477_n652), .CO(
        DP_OP_423J2_125_3477_n454), .S(DP_OP_423J2_125_3477_n455) );
  FADDX1_HVT DP_OP_423J2_125_3477_U319 ( .A(DP_OP_423J2_125_3477_n656), .B(
        DP_OP_423J2_125_3477_n654), .CI(DP_OP_423J2_125_3477_n644), .CO(
        DP_OP_423J2_125_3477_n452), .S(DP_OP_423J2_125_3477_n453) );
  FADDX1_HVT DP_OP_423J2_125_3477_U318 ( .A(DP_OP_423J2_125_3477_n642), .B(
        DP_OP_423J2_125_3477_n632), .CI(DP_OP_423J2_125_3477_n626), .CO(
        DP_OP_423J2_125_3477_n450), .S(DP_OP_423J2_125_3477_n451) );
  FADDX1_HVT DP_OP_423J2_125_3477_U317 ( .A(DP_OP_423J2_125_3477_n640), .B(
        DP_OP_423J2_125_3477_n634), .CI(DP_OP_423J2_125_3477_n628), .CO(
        DP_OP_423J2_125_3477_n448), .S(DP_OP_423J2_125_3477_n449) );
  FADDX1_HVT DP_OP_423J2_125_3477_U316 ( .A(DP_OP_423J2_125_3477_n638), .B(
        DP_OP_423J2_125_3477_n636), .CI(DP_OP_423J2_125_3477_n630), .CO(
        DP_OP_423J2_125_3477_n446), .S(DP_OP_423J2_125_3477_n447) );
  FADDX1_HVT DP_OP_423J2_125_3477_U315 ( .A(DP_OP_423J2_125_3477_n624), .B(
        DP_OP_423J2_125_3477_n620), .CI(DP_OP_423J2_125_3477_n473), .CO(
        DP_OP_423J2_125_3477_n444), .S(DP_OP_423J2_125_3477_n445) );
  FADDX1_HVT DP_OP_423J2_125_3477_U314 ( .A(DP_OP_423J2_125_3477_n622), .B(
        DP_OP_423J2_125_3477_n491), .CI(DP_OP_423J2_125_3477_n485), .CO(
        DP_OP_423J2_125_3477_n442), .S(DP_OP_423J2_125_3477_n443) );
  FADDX1_HVT DP_OP_423J2_125_3477_U313 ( .A(DP_OP_423J2_125_3477_n489), .B(
        DP_OP_423J2_125_3477_n475), .CI(DP_OP_423J2_125_3477_n616), .CO(
        DP_OP_423J2_125_3477_n440), .S(DP_OP_423J2_125_3477_n441) );
  FADDX1_HVT DP_OP_423J2_125_3477_U312 ( .A(DP_OP_423J2_125_3477_n493), .B(
        DP_OP_423J2_125_3477_n481), .CI(DP_OP_423J2_125_3477_n618), .CO(
        DP_OP_423J2_125_3477_n438), .S(DP_OP_423J2_125_3477_n439) );
  FADDX1_HVT DP_OP_423J2_125_3477_U311 ( .A(DP_OP_423J2_125_3477_n479), .B(
        DP_OP_423J2_125_3477_n483), .CI(DP_OP_423J2_125_3477_n487), .CO(
        DP_OP_423J2_125_3477_n436), .S(DP_OP_423J2_125_3477_n437) );
  FADDX1_HVT DP_OP_423J2_125_3477_U310 ( .A(DP_OP_423J2_125_3477_n477), .B(
        DP_OP_423J2_125_3477_n471), .CI(DP_OP_423J2_125_3477_n469), .CO(
        DP_OP_423J2_125_3477_n434), .S(DP_OP_423J2_125_3477_n435) );
  FADDX1_HVT DP_OP_423J2_125_3477_U309 ( .A(DP_OP_423J2_125_3477_n467), .B(
        DP_OP_423J2_125_3477_n465), .CI(DP_OP_423J2_125_3477_n463), .CO(
        DP_OP_423J2_125_3477_n432), .S(DP_OP_423J2_125_3477_n433) );
  FADDX1_HVT DP_OP_423J2_125_3477_U308 ( .A(DP_OP_423J2_125_3477_n461), .B(
        DP_OP_423J2_125_3477_n614), .CI(DP_OP_423J2_125_3477_n612), .CO(
        DP_OP_423J2_125_3477_n430), .S(DP_OP_423J2_125_3477_n431) );
  FADDX1_HVT DP_OP_423J2_125_3477_U307 ( .A(DP_OP_423J2_125_3477_n610), .B(
        DP_OP_423J2_125_3477_n606), .CI(DP_OP_423J2_125_3477_n608), .CO(
        DP_OP_423J2_125_3477_n428), .S(DP_OP_423J2_125_3477_n429) );
  FADDX1_HVT DP_OP_423J2_125_3477_U306 ( .A(DP_OP_423J2_125_3477_n604), .B(
        DP_OP_423J2_125_3477_n600), .CI(DP_OP_423J2_125_3477_n602), .CO(
        DP_OP_423J2_125_3477_n426), .S(DP_OP_423J2_125_3477_n427) );
  FADDX1_HVT DP_OP_423J2_125_3477_U305 ( .A(DP_OP_423J2_125_3477_n598), .B(
        DP_OP_423J2_125_3477_n594), .CI(DP_OP_423J2_125_3477_n453), .CO(
        DP_OP_423J2_125_3477_n424), .S(DP_OP_423J2_125_3477_n425) );
  FADDX1_HVT DP_OP_423J2_125_3477_U304 ( .A(DP_OP_423J2_125_3477_n459), .B(
        DP_OP_423J2_125_3477_n596), .CI(DP_OP_423J2_125_3477_n457), .CO(
        DP_OP_423J2_125_3477_n422), .S(DP_OP_423J2_125_3477_n423) );
  FADDX1_HVT DP_OP_423J2_125_3477_U303 ( .A(DP_OP_423J2_125_3477_n592), .B(
        DP_OP_423J2_125_3477_n455), .CI(DP_OP_423J2_125_3477_n586), .CO(
        DP_OP_423J2_125_3477_n420), .S(DP_OP_423J2_125_3477_n421) );
  FADDX1_HVT DP_OP_423J2_125_3477_U302 ( .A(DP_OP_423J2_125_3477_n590), .B(
        DP_OP_423J2_125_3477_n588), .CI(DP_OP_423J2_125_3477_n584), .CO(
        DP_OP_423J2_125_3477_n418), .S(DP_OP_423J2_125_3477_n419) );
  FADDX1_HVT DP_OP_423J2_125_3477_U301 ( .A(DP_OP_423J2_125_3477_n449), .B(
        DP_OP_423J2_125_3477_n447), .CI(DP_OP_423J2_125_3477_n578), .CO(
        DP_OP_423J2_125_3477_n416), .S(DP_OP_423J2_125_3477_n417) );
  FADDX1_HVT DP_OP_423J2_125_3477_U300 ( .A(DP_OP_423J2_125_3477_n582), .B(
        DP_OP_423J2_125_3477_n451), .CI(DP_OP_423J2_125_3477_n580), .CO(
        DP_OP_423J2_125_3477_n414), .S(DP_OP_423J2_125_3477_n415) );
  FADDX1_HVT DP_OP_423J2_125_3477_U299 ( .A(DP_OP_423J2_125_3477_n445), .B(
        DP_OP_423J2_125_3477_n443), .CI(DP_OP_423J2_125_3477_n576), .CO(
        DP_OP_423J2_125_3477_n412), .S(DP_OP_423J2_125_3477_n413) );
  FADDX1_HVT DP_OP_423J2_125_3477_U298 ( .A(DP_OP_423J2_125_3477_n441), .B(
        DP_OP_423J2_125_3477_n437), .CI(DP_OP_423J2_125_3477_n435), .CO(
        DP_OP_423J2_125_3477_n410), .S(DP_OP_423J2_125_3477_n411) );
  FADDX1_HVT DP_OP_423J2_125_3477_U297 ( .A(DP_OP_423J2_125_3477_n439), .B(
        DP_OP_423J2_125_3477_n433), .CI(DP_OP_423J2_125_3477_n574), .CO(
        DP_OP_423J2_125_3477_n408), .S(DP_OP_423J2_125_3477_n409) );
  FADDX1_HVT DP_OP_423J2_125_3477_U296 ( .A(DP_OP_423J2_125_3477_n572), .B(
        DP_OP_423J2_125_3477_n570), .CI(DP_OP_423J2_125_3477_n431), .CO(
        DP_OP_423J2_125_3477_n406), .S(DP_OP_423J2_125_3477_n407) );
  FADDX1_HVT DP_OP_423J2_125_3477_U295 ( .A(DP_OP_423J2_125_3477_n568), .B(
        DP_OP_423J2_125_3477_n566), .CI(DP_OP_423J2_125_3477_n429), .CO(
        DP_OP_423J2_125_3477_n404), .S(DP_OP_423J2_125_3477_n405) );
  FADDX1_HVT DP_OP_423J2_125_3477_U294 ( .A(DP_OP_423J2_125_3477_n564), .B(
        DP_OP_423J2_125_3477_n562), .CI(DP_OP_423J2_125_3477_n560), .CO(
        DP_OP_423J2_125_3477_n402), .S(DP_OP_423J2_125_3477_n403) );
  FADDX1_HVT DP_OP_423J2_125_3477_U293 ( .A(DP_OP_423J2_125_3477_n427), .B(
        DP_OP_423J2_125_3477_n558), .CI(DP_OP_423J2_125_3477_n425), .CO(
        DP_OP_423J2_125_3477_n400), .S(DP_OP_423J2_125_3477_n401) );
  FADDX1_HVT DP_OP_423J2_125_3477_U292 ( .A(DP_OP_423J2_125_3477_n556), .B(
        DP_OP_423J2_125_3477_n550), .CI(DP_OP_423J2_125_3477_n419), .CO(
        DP_OP_423J2_125_3477_n398), .S(DP_OP_423J2_125_3477_n399) );
  FADDX1_HVT DP_OP_423J2_125_3477_U291 ( .A(DP_OP_423J2_125_3477_n423), .B(
        DP_OP_423J2_125_3477_n552), .CI(DP_OP_423J2_125_3477_n421), .CO(
        DP_OP_423J2_125_3477_n396), .S(DP_OP_423J2_125_3477_n397) );
  FADDX1_HVT DP_OP_423J2_125_3477_U290 ( .A(DP_OP_423J2_125_3477_n554), .B(
        DP_OP_423J2_125_3477_n417), .CI(DP_OP_423J2_125_3477_n415), .CO(
        DP_OP_423J2_125_3477_n394), .S(DP_OP_423J2_125_3477_n395) );
  FADDX1_HVT DP_OP_423J2_125_3477_U289 ( .A(DP_OP_423J2_125_3477_n548), .B(
        DP_OP_423J2_125_3477_n546), .CI(DP_OP_423J2_125_3477_n413), .CO(
        DP_OP_423J2_125_3477_n392), .S(DP_OP_423J2_125_3477_n393) );
  FADDX1_HVT DP_OP_423J2_125_3477_U288 ( .A(DP_OP_423J2_125_3477_n411), .B(
        DP_OP_423J2_125_3477_n544), .CI(DP_OP_423J2_125_3477_n409), .CO(
        DP_OP_423J2_125_3477_n390), .S(DP_OP_423J2_125_3477_n391) );
  FADDX1_HVT DP_OP_423J2_125_3477_U287 ( .A(DP_OP_423J2_125_3477_n542), .B(
        DP_OP_423J2_125_3477_n540), .CI(DP_OP_423J2_125_3477_n407), .CO(
        DP_OP_423J2_125_3477_n388), .S(DP_OP_423J2_125_3477_n389) );
  FADDX1_HVT DP_OP_423J2_125_3477_U286 ( .A(DP_OP_423J2_125_3477_n538), .B(
        DP_OP_423J2_125_3477_n405), .CI(DP_OP_423J2_125_3477_n403), .CO(
        DP_OP_423J2_125_3477_n386), .S(DP_OP_423J2_125_3477_n387) );
  FADDX1_HVT DP_OP_423J2_125_3477_U285 ( .A(DP_OP_423J2_125_3477_n536), .B(
        DP_OP_423J2_125_3477_n534), .CI(DP_OP_423J2_125_3477_n532), .CO(
        DP_OP_423J2_125_3477_n384), .S(DP_OP_423J2_125_3477_n385) );
  FADDX1_HVT DP_OP_423J2_125_3477_U284 ( .A(DP_OP_423J2_125_3477_n401), .B(
        DP_OP_423J2_125_3477_n530), .CI(DP_OP_423J2_125_3477_n399), .CO(
        DP_OP_423J2_125_3477_n382), .S(DP_OP_423J2_125_3477_n383) );
  FADDX1_HVT DP_OP_423J2_125_3477_U283 ( .A(DP_OP_423J2_125_3477_n397), .B(
        DP_OP_423J2_125_3477_n528), .CI(DP_OP_423J2_125_3477_n395), .CO(
        DP_OP_423J2_125_3477_n380), .S(DP_OP_423J2_125_3477_n381) );
  FADDX1_HVT DP_OP_423J2_125_3477_U282 ( .A(DP_OP_423J2_125_3477_n526), .B(
        DP_OP_423J2_125_3477_n393), .CI(DP_OP_423J2_125_3477_n524), .CO(
        DP_OP_423J2_125_3477_n378), .S(DP_OP_423J2_125_3477_n379) );
  FADDX1_HVT DP_OP_423J2_125_3477_U281 ( .A(DP_OP_423J2_125_3477_n391), .B(
        DP_OP_423J2_125_3477_n522), .CI(DP_OP_423J2_125_3477_n389), .CO(
        DP_OP_423J2_125_3477_n376), .S(DP_OP_423J2_125_3477_n377) );
  FADDX1_HVT DP_OP_423J2_125_3477_U280 ( .A(DP_OP_423J2_125_3477_n520), .B(
        DP_OP_423J2_125_3477_n518), .CI(DP_OP_423J2_125_3477_n387), .CO(
        DP_OP_423J2_125_3477_n374), .S(DP_OP_423J2_125_3477_n375) );
  FADDX1_HVT DP_OP_423J2_125_3477_U279 ( .A(DP_OP_423J2_125_3477_n385), .B(
        DP_OP_423J2_125_3477_n516), .CI(DP_OP_423J2_125_3477_n514), .CO(
        DP_OP_423J2_125_3477_n372), .S(DP_OP_423J2_125_3477_n373) );
  FADDX1_HVT DP_OP_423J2_125_3477_U278 ( .A(DP_OP_423J2_125_3477_n383), .B(
        DP_OP_423J2_125_3477_n381), .CI(DP_OP_423J2_125_3477_n512), .CO(
        DP_OP_423J2_125_3477_n370), .S(DP_OP_423J2_125_3477_n371) );
  FADDX1_HVT DP_OP_423J2_125_3477_U277 ( .A(DP_OP_423J2_125_3477_n379), .B(
        DP_OP_423J2_125_3477_n510), .CI(DP_OP_423J2_125_3477_n377), .CO(
        DP_OP_423J2_125_3477_n368), .S(DP_OP_423J2_125_3477_n369) );
  FADDX1_HVT DP_OP_423J2_125_3477_U276 ( .A(DP_OP_423J2_125_3477_n508), .B(
        DP_OP_423J2_125_3477_n375), .CI(DP_OP_423J2_125_3477_n506), .CO(
        DP_OP_423J2_125_3477_n366), .S(DP_OP_423J2_125_3477_n367) );
  FADDX1_HVT DP_OP_423J2_125_3477_U275 ( .A(DP_OP_423J2_125_3477_n373), .B(
        DP_OP_423J2_125_3477_n504), .CI(DP_OP_423J2_125_3477_n371), .CO(
        DP_OP_423J2_125_3477_n364), .S(DP_OP_423J2_125_3477_n365) );
  FADDX1_HVT DP_OP_423J2_125_3477_U274 ( .A(DP_OP_423J2_125_3477_n502), .B(
        DP_OP_423J2_125_3477_n369), .CI(DP_OP_423J2_125_3477_n500), .CO(
        DP_OP_423J2_125_3477_n362), .S(DP_OP_423J2_125_3477_n363) );
  FADDX1_HVT DP_OP_423J2_125_3477_U273 ( .A(DP_OP_423J2_125_3477_n367), .B(
        DP_OP_423J2_125_3477_n365), .CI(DP_OP_423J2_125_3477_n498), .CO(
        DP_OP_423J2_125_3477_n360), .S(DP_OP_423J2_125_3477_n361) );
  FADDX1_HVT DP_OP_423J2_125_3477_U272 ( .A(DP_OP_423J2_125_3477_n496), .B(
        DP_OP_423J2_125_3477_n363), .CI(DP_OP_423J2_125_3477_n361), .CO(
        DP_OP_423J2_125_3477_n358), .S(DP_OP_423J2_125_3477_n359) );
  FADDX1_HVT DP_OP_423J2_125_3477_U270 ( .A(DP_OP_423J2_125_3477_n1993), .B(
        DP_OP_423J2_125_3477_n2477), .CI(DP_OP_423J2_125_3477_n1949), .CO(
        DP_OP_423J2_125_3477_n354), .S(DP_OP_423J2_125_3477_n355) );
  FADDX1_HVT DP_OP_423J2_125_3477_U269 ( .A(DP_OP_423J2_125_3477_n2653), .B(
        DP_OP_423J2_125_3477_n2521), .CI(DP_OP_423J2_125_3477_n2738), .CO(
        DP_OP_423J2_125_3477_n352), .S(DP_OP_423J2_125_3477_n353) );
  FADDX1_HVT DP_OP_423J2_125_3477_U268 ( .A(DP_OP_423J2_125_3477_n2081), .B(
        DP_OP_423J2_125_3477_n2565), .CI(DP_OP_423J2_125_3477_n2433), .CO(
        DP_OP_423J2_125_3477_n350), .S(DP_OP_423J2_125_3477_n351) );
  FADDX1_HVT DP_OP_423J2_125_3477_U267 ( .A(DP_OP_423J2_125_3477_n1861), .B(
        DP_OP_423J2_125_3477_n2037), .CI(DP_OP_423J2_125_3477_n1905), .CO(
        DP_OP_423J2_125_3477_n348), .S(DP_OP_423J2_125_3477_n349) );
  FADDX1_HVT DP_OP_423J2_125_3477_U266 ( .A(DP_OP_423J2_125_3477_n2826), .B(
        DP_OP_423J2_125_3477_n2870), .CI(DP_OP_423J2_125_3477_n2169), .CO(
        DP_OP_423J2_125_3477_n346), .S(DP_OP_423J2_125_3477_n347) );
  FADDX1_HVT DP_OP_423J2_125_3477_U265 ( .A(DP_OP_423J2_125_3477_n2782), .B(
        DP_OP_423J2_125_3477_n1773), .CI(DP_OP_423J2_125_3477_n1817), .CO(
        DP_OP_423J2_125_3477_n344), .S(DP_OP_423J2_125_3477_n345) );
  FADDX1_HVT DP_OP_423J2_125_3477_U264 ( .A(DP_OP_423J2_125_3477_n2345), .B(
        DP_OP_423J2_125_3477_n2301), .CI(DP_OP_423J2_125_3477_n2257), .CO(
        DP_OP_423J2_125_3477_n342), .S(DP_OP_423J2_125_3477_n343) );
  FADDX1_HVT DP_OP_423J2_125_3477_U263 ( .A(DP_OP_423J2_125_3477_n2609), .B(
        DP_OP_423J2_125_3477_n2125), .CI(DP_OP_423J2_125_3477_n357), .CO(
        DP_OP_423J2_125_3477_n340), .S(DP_OP_423J2_125_3477_n341) );
  FADDX1_HVT DP_OP_423J2_125_3477_U262 ( .A(DP_OP_423J2_125_3477_n2213), .B(
        DP_OP_423J2_125_3477_n2389), .CI(DP_OP_423J2_125_3477_n492), .CO(
        DP_OP_423J2_125_3477_n338), .S(DP_OP_423J2_125_3477_n339) );
  FADDX1_HVT DP_OP_423J2_125_3477_U261 ( .A(DP_OP_423J2_125_3477_n490), .B(
        DP_OP_423J2_125_3477_n472), .CI(DP_OP_423J2_125_3477_n474), .CO(
        DP_OP_423J2_125_3477_n336), .S(DP_OP_423J2_125_3477_n337) );
  FADDX1_HVT DP_OP_423J2_125_3477_U260 ( .A(DP_OP_423J2_125_3477_n488), .B(
        DP_OP_423J2_125_3477_n476), .CI(DP_OP_423J2_125_3477_n478), .CO(
        DP_OP_423J2_125_3477_n334), .S(DP_OP_423J2_125_3477_n335) );
  FADDX1_HVT DP_OP_423J2_125_3477_U259 ( .A(DP_OP_423J2_125_3477_n486), .B(
        DP_OP_423J2_125_3477_n480), .CI(DP_OP_423J2_125_3477_n482), .CO(
        DP_OP_423J2_125_3477_n332), .S(DP_OP_423J2_125_3477_n333) );
  FADDX1_HVT DP_OP_423J2_125_3477_U258 ( .A(DP_OP_423J2_125_3477_n484), .B(
        DP_OP_423J2_125_3477_n470), .CI(DP_OP_423J2_125_3477_n468), .CO(
        DP_OP_423J2_125_3477_n330), .S(DP_OP_423J2_125_3477_n331) );
  FADDX1_HVT DP_OP_423J2_125_3477_U257 ( .A(DP_OP_423J2_125_3477_n466), .B(
        DP_OP_423J2_125_3477_n464), .CI(DP_OP_423J2_125_3477_n462), .CO(
        DP_OP_423J2_125_3477_n328), .S(DP_OP_423J2_125_3477_n329) );
  FADDX1_HVT DP_OP_423J2_125_3477_U256 ( .A(DP_OP_423J2_125_3477_n460), .B(
        DP_OP_423J2_125_3477_n355), .CI(DP_OP_423J2_125_3477_n349), .CO(
        DP_OP_423J2_125_3477_n326), .S(DP_OP_423J2_125_3477_n327) );
  FADDX1_HVT DP_OP_423J2_125_3477_U255 ( .A(DP_OP_423J2_125_3477_n347), .B(
        DP_OP_423J2_125_3477_n343), .CI(DP_OP_423J2_125_3477_n341), .CO(
        DP_OP_423J2_125_3477_n324), .S(DP_OP_423J2_125_3477_n325) );
  FADDX1_HVT DP_OP_423J2_125_3477_U254 ( .A(DP_OP_423J2_125_3477_n345), .B(
        DP_OP_423J2_125_3477_n353), .CI(DP_OP_423J2_125_3477_n351), .CO(
        DP_OP_423J2_125_3477_n322), .S(DP_OP_423J2_125_3477_n323) );
  FADDX1_HVT DP_OP_423J2_125_3477_U253 ( .A(DP_OP_423J2_125_3477_n458), .B(
        DP_OP_423J2_125_3477_n456), .CI(DP_OP_423J2_125_3477_n452), .CO(
        DP_OP_423J2_125_3477_n320), .S(DP_OP_423J2_125_3477_n321) );
  FADDX1_HVT DP_OP_423J2_125_3477_U252 ( .A(DP_OP_423J2_125_3477_n454), .B(
        DP_OP_423J2_125_3477_n450), .CI(DP_OP_423J2_125_3477_n448), .CO(
        DP_OP_423J2_125_3477_n318), .S(DP_OP_423J2_125_3477_n319) );
  FADDX1_HVT DP_OP_423J2_125_3477_U251 ( .A(DP_OP_423J2_125_3477_n446), .B(
        DP_OP_423J2_125_3477_n339), .CI(DP_OP_423J2_125_3477_n444), .CO(
        DP_OP_423J2_125_3477_n316), .S(DP_OP_423J2_125_3477_n317) );
  FADDX1_HVT DP_OP_423J2_125_3477_U250 ( .A(DP_OP_423J2_125_3477_n442), .B(
        DP_OP_423J2_125_3477_n440), .CI(DP_OP_423J2_125_3477_n333), .CO(
        DP_OP_423J2_125_3477_n314), .S(DP_OP_423J2_125_3477_n315) );
  FADDX1_HVT DP_OP_423J2_125_3477_U249 ( .A(DP_OP_423J2_125_3477_n438), .B(
        DP_OP_423J2_125_3477_n436), .CI(DP_OP_423J2_125_3477_n331), .CO(
        DP_OP_423J2_125_3477_n312), .S(DP_OP_423J2_125_3477_n313) );
  FADDX1_HVT DP_OP_423J2_125_3477_U248 ( .A(DP_OP_423J2_125_3477_n335), .B(
        DP_OP_423J2_125_3477_n337), .CI(DP_OP_423J2_125_3477_n434), .CO(
        DP_OP_423J2_125_3477_n310), .S(DP_OP_423J2_125_3477_n311) );
  FADDX1_HVT DP_OP_423J2_125_3477_U247 ( .A(DP_OP_423J2_125_3477_n432), .B(
        DP_OP_423J2_125_3477_n329), .CI(DP_OP_423J2_125_3477_n430), .CO(
        DP_OP_423J2_125_3477_n308), .S(DP_OP_423J2_125_3477_n309) );
  FADDX1_HVT DP_OP_423J2_125_3477_U246 ( .A(DP_OP_423J2_125_3477_n327), .B(
        DP_OP_423J2_125_3477_n323), .CI(DP_OP_423J2_125_3477_n428), .CO(
        DP_OP_423J2_125_3477_n306), .S(DP_OP_423J2_125_3477_n307) );
  FADDX1_HVT DP_OP_423J2_125_3477_U245 ( .A(DP_OP_423J2_125_3477_n325), .B(
        DP_OP_423J2_125_3477_n426), .CI(DP_OP_423J2_125_3477_n424), .CO(
        DP_OP_423J2_125_3477_n304), .S(DP_OP_423J2_125_3477_n305) );
  FADDX1_HVT DP_OP_423J2_125_3477_U244 ( .A(DP_OP_423J2_125_3477_n422), .B(
        DP_OP_423J2_125_3477_n321), .CI(DP_OP_423J2_125_3477_n418), .CO(
        DP_OP_423J2_125_3477_n302), .S(DP_OP_423J2_125_3477_n303) );
  FADDX1_HVT DP_OP_423J2_125_3477_U243 ( .A(DP_OP_423J2_125_3477_n420), .B(
        DP_OP_423J2_125_3477_n319), .CI(DP_OP_423J2_125_3477_n416), .CO(
        DP_OP_423J2_125_3477_n300), .S(DP_OP_423J2_125_3477_n301) );
  FADDX1_HVT DP_OP_423J2_125_3477_U242 ( .A(DP_OP_423J2_125_3477_n414), .B(
        DP_OP_423J2_125_3477_n317), .CI(DP_OP_423J2_125_3477_n412), .CO(
        DP_OP_423J2_125_3477_n298), .S(DP_OP_423J2_125_3477_n299) );
  FADDX1_HVT DP_OP_423J2_125_3477_U241 ( .A(DP_OP_423J2_125_3477_n315), .B(
        DP_OP_423J2_125_3477_n410), .CI(DP_OP_423J2_125_3477_n311), .CO(
        DP_OP_423J2_125_3477_n296), .S(DP_OP_423J2_125_3477_n297) );
  FADDX1_HVT DP_OP_423J2_125_3477_U240 ( .A(DP_OP_423J2_125_3477_n313), .B(
        DP_OP_423J2_125_3477_n408), .CI(DP_OP_423J2_125_3477_n309), .CO(
        DP_OP_423J2_125_3477_n294), .S(DP_OP_423J2_125_3477_n295) );
  FADDX1_HVT DP_OP_423J2_125_3477_U239 ( .A(DP_OP_423J2_125_3477_n406), .B(
        DP_OP_423J2_125_3477_n307), .CI(DP_OP_423J2_125_3477_n404), .CO(
        DP_OP_423J2_125_3477_n292), .S(DP_OP_423J2_125_3477_n293) );
  FADDX1_HVT DP_OP_423J2_125_3477_U238 ( .A(DP_OP_423J2_125_3477_n402), .B(
        DP_OP_423J2_125_3477_n400), .CI(DP_OP_423J2_125_3477_n305), .CO(
        DP_OP_423J2_125_3477_n290), .S(DP_OP_423J2_125_3477_n291) );
  FADDX1_HVT DP_OP_423J2_125_3477_U237 ( .A(DP_OP_423J2_125_3477_n398), .B(
        DP_OP_423J2_125_3477_n396), .CI(DP_OP_423J2_125_3477_n394), .CO(
        DP_OP_423J2_125_3477_n288), .S(DP_OP_423J2_125_3477_n289) );
  FADDX1_HVT DP_OP_423J2_125_3477_U236 ( .A(DP_OP_423J2_125_3477_n303), .B(
        DP_OP_423J2_125_3477_n301), .CI(DP_OP_423J2_125_3477_n299), .CO(
        DP_OP_423J2_125_3477_n286), .S(DP_OP_423J2_125_3477_n287) );
  FADDX1_HVT DP_OP_423J2_125_3477_U235 ( .A(DP_OP_423J2_125_3477_n392), .B(
        DP_OP_423J2_125_3477_n297), .CI(DP_OP_423J2_125_3477_n390), .CO(
        DP_OP_423J2_125_3477_n284), .S(DP_OP_423J2_125_3477_n285) );
  FADDX1_HVT DP_OP_423J2_125_3477_U234 ( .A(DP_OP_423J2_125_3477_n295), .B(
        DP_OP_423J2_125_3477_n388), .CI(DP_OP_423J2_125_3477_n293), .CO(
        DP_OP_423J2_125_3477_n282), .S(DP_OP_423J2_125_3477_n283) );
  FADDX1_HVT DP_OP_423J2_125_3477_U233 ( .A(DP_OP_423J2_125_3477_n386), .B(
        DP_OP_423J2_125_3477_n384), .CI(DP_OP_423J2_125_3477_n291), .CO(
        DP_OP_423J2_125_3477_n280), .S(DP_OP_423J2_125_3477_n281) );
  FADDX1_HVT DP_OP_423J2_125_3477_U232 ( .A(DP_OP_423J2_125_3477_n382), .B(
        DP_OP_423J2_125_3477_n289), .CI(DP_OP_423J2_125_3477_n380), .CO(
        DP_OP_423J2_125_3477_n278), .S(DP_OP_423J2_125_3477_n279) );
  FADDX1_HVT DP_OP_423J2_125_3477_U231 ( .A(DP_OP_423J2_125_3477_n287), .B(
        DP_OP_423J2_125_3477_n378), .CI(DP_OP_423J2_125_3477_n285), .CO(
        DP_OP_423J2_125_3477_n276), .S(DP_OP_423J2_125_3477_n277) );
  FADDX1_HVT DP_OP_423J2_125_3477_U230 ( .A(DP_OP_423J2_125_3477_n376), .B(
        DP_OP_423J2_125_3477_n283), .CI(DP_OP_423J2_125_3477_n374), .CO(
        DP_OP_423J2_125_3477_n274), .S(DP_OP_423J2_125_3477_n275) );
  FADDX1_HVT DP_OP_423J2_125_3477_U229 ( .A(DP_OP_423J2_125_3477_n281), .B(
        DP_OP_423J2_125_3477_n372), .CI(DP_OP_423J2_125_3477_n279), .CO(
        DP_OP_423J2_125_3477_n272), .S(DP_OP_423J2_125_3477_n273) );
  FADDX1_HVT DP_OP_423J2_125_3477_U228 ( .A(DP_OP_423J2_125_3477_n370), .B(
        DP_OP_423J2_125_3477_n277), .CI(DP_OP_423J2_125_3477_n368), .CO(
        DP_OP_423J2_125_3477_n270), .S(DP_OP_423J2_125_3477_n271) );
  FADDX1_HVT DP_OP_423J2_125_3477_U227 ( .A(DP_OP_423J2_125_3477_n275), .B(
        DP_OP_423J2_125_3477_n366), .CI(DP_OP_423J2_125_3477_n273), .CO(
        DP_OP_423J2_125_3477_n268), .S(DP_OP_423J2_125_3477_n269) );
  FADDX1_HVT DP_OP_423J2_125_3477_U226 ( .A(DP_OP_423J2_125_3477_n364), .B(
        DP_OP_423J2_125_3477_n271), .CI(DP_OP_423J2_125_3477_n362), .CO(
        DP_OP_423J2_125_3477_n266), .S(DP_OP_423J2_125_3477_n267) );
  FADDX1_HVT DP_OP_423J2_125_3477_U225 ( .A(DP_OP_423J2_125_3477_n269), .B(
        DP_OP_423J2_125_3477_n360), .CI(DP_OP_423J2_125_3477_n267), .CO(
        DP_OP_423J2_125_3477_n264), .S(DP_OP_423J2_125_3477_n265) );
  FADDX1_HVT DP_OP_423J2_125_3477_U224 ( .A(DP_OP_423J2_125_3477_n356), .B(
        DP_OP_423J2_125_3477_n1772), .CI(DP_OP_423J2_125_3477_n354), .CO(
        DP_OP_423J2_125_3477_n262), .S(DP_OP_423J2_125_3477_n263) );
  FADDX1_HVT DP_OP_423J2_125_3477_U223 ( .A(DP_OP_423J2_125_3477_n344), .B(
        DP_OP_423J2_125_3477_n340), .CI(DP_OP_423J2_125_3477_n352), .CO(
        DP_OP_423J2_125_3477_n260), .S(DP_OP_423J2_125_3477_n261) );
  FADDX1_HVT DP_OP_423J2_125_3477_U222 ( .A(DP_OP_423J2_125_3477_n350), .B(
        DP_OP_423J2_125_3477_n348), .CI(DP_OP_423J2_125_3477_n346), .CO(
        DP_OP_423J2_125_3477_n258), .S(DP_OP_423J2_125_3477_n259) );
  FADDX1_HVT DP_OP_423J2_125_3477_U221 ( .A(DP_OP_423J2_125_3477_n342), .B(
        DP_OP_423J2_125_3477_n338), .CI(DP_OP_423J2_125_3477_n336), .CO(
        DP_OP_423J2_125_3477_n256), .S(DP_OP_423J2_125_3477_n257) );
  FADDX1_HVT DP_OP_423J2_125_3477_U220 ( .A(DP_OP_423J2_125_3477_n334), .B(
        DP_OP_423J2_125_3477_n332), .CI(DP_OP_423J2_125_3477_n330), .CO(
        DP_OP_423J2_125_3477_n254), .S(DP_OP_423J2_125_3477_n255) );
  FADDX1_HVT DP_OP_423J2_125_3477_U219 ( .A(DP_OP_423J2_125_3477_n328), .B(
        DP_OP_423J2_125_3477_n263), .CI(DP_OP_423J2_125_3477_n326), .CO(
        DP_OP_423J2_125_3477_n252), .S(DP_OP_423J2_125_3477_n253) );
  FADDX1_HVT DP_OP_423J2_125_3477_U218 ( .A(DP_OP_423J2_125_3477_n324), .B(
        DP_OP_423J2_125_3477_n259), .CI(DP_OP_423J2_125_3477_n261), .CO(
        DP_OP_423J2_125_3477_n250), .S(DP_OP_423J2_125_3477_n251) );
  FADDX1_HVT DP_OP_423J2_125_3477_U217 ( .A(DP_OP_423J2_125_3477_n322), .B(
        DP_OP_423J2_125_3477_n320), .CI(DP_OP_423J2_125_3477_n318), .CO(
        DP_OP_423J2_125_3477_n248), .S(DP_OP_423J2_125_3477_n249) );
  FADDX1_HVT DP_OP_423J2_125_3477_U216 ( .A(DP_OP_423J2_125_3477_n316), .B(
        DP_OP_423J2_125_3477_n257), .CI(DP_OP_423J2_125_3477_n314), .CO(
        DP_OP_423J2_125_3477_n246), .S(DP_OP_423J2_125_3477_n247) );
  FADDX1_HVT DP_OP_423J2_125_3477_U215 ( .A(DP_OP_423J2_125_3477_n312), .B(
        DP_OP_423J2_125_3477_n255), .CI(DP_OP_423J2_125_3477_n310), .CO(
        DP_OP_423J2_125_3477_n244), .S(DP_OP_423J2_125_3477_n245) );
  FADDX1_HVT DP_OP_423J2_125_3477_U214 ( .A(DP_OP_423J2_125_3477_n308), .B(
        DP_OP_423J2_125_3477_n253), .CI(DP_OP_423J2_125_3477_n306), .CO(
        DP_OP_423J2_125_3477_n242), .S(DP_OP_423J2_125_3477_n243) );
  FADDX1_HVT DP_OP_423J2_125_3477_U213 ( .A(DP_OP_423J2_125_3477_n251), .B(
        DP_OP_423J2_125_3477_n304), .CI(DP_OP_423J2_125_3477_n249), .CO(
        DP_OP_423J2_125_3477_n240), .S(DP_OP_423J2_125_3477_n241) );
  FADDX1_HVT DP_OP_423J2_125_3477_U212 ( .A(DP_OP_423J2_125_3477_n302), .B(
        DP_OP_423J2_125_3477_n300), .CI(DP_OP_423J2_125_3477_n298), .CO(
        DP_OP_423J2_125_3477_n238), .S(DP_OP_423J2_125_3477_n239) );
  FADDX1_HVT DP_OP_423J2_125_3477_U211 ( .A(DP_OP_423J2_125_3477_n247), .B(
        DP_OP_423J2_125_3477_n296), .CI(DP_OP_423J2_125_3477_n245), .CO(
        DP_OP_423J2_125_3477_n236), .S(DP_OP_423J2_125_3477_n237) );
  FADDX1_HVT DP_OP_423J2_125_3477_U210 ( .A(DP_OP_423J2_125_3477_n294), .B(
        DP_OP_423J2_125_3477_n243), .CI(DP_OP_423J2_125_3477_n292), .CO(
        DP_OP_423J2_125_3477_n234), .S(DP_OP_423J2_125_3477_n235) );
  FADDX1_HVT DP_OP_423J2_125_3477_U209 ( .A(DP_OP_423J2_125_3477_n290), .B(
        DP_OP_423J2_125_3477_n241), .CI(DP_OP_423J2_125_3477_n288), .CO(
        DP_OP_423J2_125_3477_n232), .S(DP_OP_423J2_125_3477_n233) );
  FADDX1_HVT DP_OP_423J2_125_3477_U208 ( .A(DP_OP_423J2_125_3477_n286), .B(
        DP_OP_423J2_125_3477_n239), .CI(DP_OP_423J2_125_3477_n284), .CO(
        DP_OP_423J2_125_3477_n230), .S(DP_OP_423J2_125_3477_n231) );
  FADDX1_HVT DP_OP_423J2_125_3477_U207 ( .A(DP_OP_423J2_125_3477_n237), .B(
        DP_OP_423J2_125_3477_n282), .CI(DP_OP_423J2_125_3477_n235), .CO(
        DP_OP_423J2_125_3477_n228), .S(DP_OP_423J2_125_3477_n229) );
  FADDX1_HVT DP_OP_423J2_125_3477_U206 ( .A(DP_OP_423J2_125_3477_n280), .B(
        DP_OP_423J2_125_3477_n233), .CI(DP_OP_423J2_125_3477_n278), .CO(
        DP_OP_423J2_125_3477_n226), .S(DP_OP_423J2_125_3477_n227) );
  FADDX1_HVT DP_OP_423J2_125_3477_U205 ( .A(DP_OP_423J2_125_3477_n231), .B(
        DP_OP_423J2_125_3477_n276), .CI(DP_OP_423J2_125_3477_n229), .CO(
        DP_OP_423J2_125_3477_n224), .S(DP_OP_423J2_125_3477_n225) );
  FADDX1_HVT DP_OP_423J2_125_3477_U204 ( .A(DP_OP_423J2_125_3477_n274), .B(
        DP_OP_423J2_125_3477_n272), .CI(DP_OP_423J2_125_3477_n227), .CO(
        DP_OP_423J2_125_3477_n222), .S(DP_OP_423J2_125_3477_n223) );
  FADDX1_HVT DP_OP_423J2_125_3477_U203 ( .A(DP_OP_423J2_125_3477_n270), .B(
        DP_OP_423J2_125_3477_n225), .CI(DP_OP_423J2_125_3477_n268), .CO(
        DP_OP_423J2_125_3477_n220), .S(DP_OP_423J2_125_3477_n221) );
  FADDX1_HVT DP_OP_423J2_125_3477_U202 ( .A(DP_OP_423J2_125_3477_n223), .B(
        DP_OP_423J2_125_3477_n266), .CI(DP_OP_423J2_125_3477_n221), .CO(
        DP_OP_423J2_125_3477_n218), .S(DP_OP_423J2_125_3477_n219) );
  FADDX1_HVT DP_OP_423J2_125_3477_U201 ( .A(DP_OP_423J2_125_3477_n1771), .B(
        DP_OP_423J2_125_3477_n262), .CI(DP_OP_423J2_125_3477_n260), .CO(
        DP_OP_423J2_125_3477_n216), .S(DP_OP_423J2_125_3477_n217) );
  FADDX1_HVT DP_OP_423J2_125_3477_U200 ( .A(DP_OP_423J2_125_3477_n258), .B(
        DP_OP_423J2_125_3477_n256), .CI(DP_OP_423J2_125_3477_n254), .CO(
        DP_OP_423J2_125_3477_n214), .S(DP_OP_423J2_125_3477_n215) );
  FADDX1_HVT DP_OP_423J2_125_3477_U199 ( .A(DP_OP_423J2_125_3477_n252), .B(
        DP_OP_423J2_125_3477_n217), .CI(DP_OP_423J2_125_3477_n250), .CO(
        DP_OP_423J2_125_3477_n212), .S(DP_OP_423J2_125_3477_n213) );
  FADDX1_HVT DP_OP_423J2_125_3477_U198 ( .A(DP_OP_423J2_125_3477_n248), .B(
        DP_OP_423J2_125_3477_n246), .CI(DP_OP_423J2_125_3477_n215), .CO(
        DP_OP_423J2_125_3477_n210), .S(DP_OP_423J2_125_3477_n211) );
  FADDX1_HVT DP_OP_423J2_125_3477_U197 ( .A(DP_OP_423J2_125_3477_n244), .B(
        DP_OP_423J2_125_3477_n242), .CI(DP_OP_423J2_125_3477_n213), .CO(
        DP_OP_423J2_125_3477_n208), .S(DP_OP_423J2_125_3477_n209) );
  FADDX1_HVT DP_OP_423J2_125_3477_U196 ( .A(DP_OP_423J2_125_3477_n240), .B(
        DP_OP_423J2_125_3477_n238), .CI(DP_OP_423J2_125_3477_n211), .CO(
        DP_OP_423J2_125_3477_n206), .S(DP_OP_423J2_125_3477_n207) );
  FADDX1_HVT DP_OP_423J2_125_3477_U195 ( .A(DP_OP_423J2_125_3477_n236), .B(
        DP_OP_423J2_125_3477_n209), .CI(DP_OP_423J2_125_3477_n234), .CO(
        DP_OP_423J2_125_3477_n204), .S(DP_OP_423J2_125_3477_n205) );
  FADDX1_HVT DP_OP_423J2_125_3477_U194 ( .A(DP_OP_423J2_125_3477_n232), .B(
        DP_OP_423J2_125_3477_n207), .CI(DP_OP_423J2_125_3477_n230), .CO(
        DP_OP_423J2_125_3477_n202), .S(DP_OP_423J2_125_3477_n203) );
  FADDX1_HVT DP_OP_423J2_125_3477_U193 ( .A(DP_OP_423J2_125_3477_n228), .B(
        DP_OP_423J2_125_3477_n205), .CI(DP_OP_423J2_125_3477_n226), .CO(
        DP_OP_423J2_125_3477_n200), .S(DP_OP_423J2_125_3477_n201) );
  FADDX1_HVT DP_OP_423J2_125_3477_U192 ( .A(DP_OP_423J2_125_3477_n203), .B(
        DP_OP_423J2_125_3477_n224), .CI(DP_OP_423J2_125_3477_n201), .CO(
        DP_OP_423J2_125_3477_n198), .S(DP_OP_423J2_125_3477_n199) );
  FADDX1_HVT DP_OP_423J2_125_3477_U191 ( .A(DP_OP_423J2_125_3477_n222), .B(
        DP_OP_423J2_125_3477_n220), .CI(DP_OP_423J2_125_3477_n199), .CO(
        DP_OP_423J2_125_3477_n196), .S(DP_OP_423J2_125_3477_n197) );
  FADDX1_HVT DP_OP_423J2_125_3477_U190 ( .A(DP_OP_423J2_125_3477_n1770), .B(
        DP_OP_423J2_125_3477_n216), .CI(DP_OP_423J2_125_3477_n214), .CO(
        DP_OP_423J2_125_3477_n194), .S(DP_OP_423J2_125_3477_n195) );
  FADDX1_HVT DP_OP_423J2_125_3477_U189 ( .A(DP_OP_423J2_125_3477_n212), .B(
        DP_OP_423J2_125_3477_n195), .CI(DP_OP_423J2_125_3477_n210), .CO(
        DP_OP_423J2_125_3477_n192), .S(DP_OP_423J2_125_3477_n193) );
  FADDX1_HVT DP_OP_423J2_125_3477_U188 ( .A(DP_OP_423J2_125_3477_n208), .B(
        DP_OP_423J2_125_3477_n206), .CI(DP_OP_423J2_125_3477_n193), .CO(
        DP_OP_423J2_125_3477_n190), .S(DP_OP_423J2_125_3477_n191) );
  FADDX1_HVT DP_OP_423J2_125_3477_U187 ( .A(DP_OP_423J2_125_3477_n204), .B(
        DP_OP_423J2_125_3477_n191), .CI(DP_OP_423J2_125_3477_n202), .CO(
        DP_OP_423J2_125_3477_n188), .S(DP_OP_423J2_125_3477_n189) );
  FADDX1_HVT DP_OP_423J2_125_3477_U186 ( .A(DP_OP_423J2_125_3477_n200), .B(
        DP_OP_423J2_125_3477_n189), .CI(DP_OP_423J2_125_3477_n198), .CO(
        DP_OP_423J2_125_3477_n186), .S(DP_OP_423J2_125_3477_n187) );
  FADDX1_HVT DP_OP_423J2_125_3477_U184 ( .A(DP_OP_423J2_125_3477_n185), .B(
        DP_OP_423J2_125_3477_n194), .CI(DP_OP_423J2_125_3477_n192), .CO(
        DP_OP_423J2_125_3477_n182), .S(DP_OP_423J2_125_3477_n183) );
  FADDX1_HVT DP_OP_423J2_125_3477_U183 ( .A(DP_OP_423J2_125_3477_n183), .B(
        DP_OP_423J2_125_3477_n190), .CI(DP_OP_423J2_125_3477_n188), .CO(
        DP_OP_423J2_125_3477_n180), .S(DP_OP_423J2_125_3477_n181) );
  FADDX1_HVT DP_OP_423J2_125_3477_U182 ( .A(DP_OP_423J2_125_3477_n1769), .B(
        DP_OP_423J2_125_3477_n184), .CI(DP_OP_423J2_125_3477_n182), .CO(
        DP_OP_423J2_125_3477_n178), .S(DP_OP_423J2_125_3477_n179) );
  FADDX1_HVT DP_OP_423J2_125_3477_U165 ( .A(DP_OP_423J2_125_3477_n1749), .B(
        DP_OP_423J2_125_3477_n1747), .CI(DP_OP_423J2_125_3477_n1745), .CO(
        DP_OP_423J2_125_3477_n127), .S(n_conv2_sum_b[0]) );
  FADDX1_HVT DP_OP_423J2_125_3477_U164 ( .A(DP_OP_423J2_125_3477_n127), .B(
        DP_OP_423J2_125_3477_n1685), .CI(DP_OP_423J2_125_3477_n1683), .CO(
        DP_OP_423J2_125_3477_n126), .S(n_conv2_sum_b[1]) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U163 ( .A1(DP_OP_423J2_125_3477_n1577), 
        .A2(DP_OP_423J2_125_3477_n1579), .Y(DP_OP_423J2_125_3477_n125) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U155 ( .A1(DP_OP_423J2_125_3477_n1423), 
        .A2(DP_OP_423J2_125_3477_n1425), .Y(DP_OP_423J2_125_3477_n120) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U154 ( .A1(DP_OP_423J2_125_3477_n1425), .A2(
        DP_OP_423J2_125_3477_n1423), .Y(DP_OP_423J2_125_3477_n119) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U149 ( .A1(DP_OP_423J2_125_3477_n1247), 
        .A2(DP_OP_423J2_125_3477_n1249), .Y(DP_OP_423J2_125_3477_n117) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U141 ( .A1(DP_OP_423J2_125_3477_n1059), 
        .A2(DP_OP_423J2_125_3477_n1061), .Y(DP_OP_423J2_125_3477_n112) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U140 ( .A1(DP_OP_423J2_125_3477_n1061), .A2(
        DP_OP_423J2_125_3477_n1059), .Y(DP_OP_423J2_125_3477_n111) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U135 ( .A1(DP_OP_423J2_125_3477_n865), .A2(
        DP_OP_423J2_125_3477_n867), .Y(DP_OP_423J2_125_3477_n109) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U127 ( .A1(DP_OP_423J2_125_3477_n669), .A2(
        DP_OP_423J2_125_3477_n864), .Y(DP_OP_423J2_125_3477_n104) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U126 ( .A1(DP_OP_423J2_125_3477_n864), .A2(
        DP_OP_423J2_125_3477_n669), .Y(DP_OP_423J2_125_3477_n103) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U120 ( .A1(DP_OP_423J2_125_3477_n495), .A2(
        DP_OP_423J2_125_3477_n668), .Y(DP_OP_423J2_125_3477_n100) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U119 ( .A1(DP_OP_423J2_125_3477_n668), .A2(
        DP_OP_423J2_125_3477_n495), .Y(DP_OP_423J2_125_3477_n99) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U114 ( .A1(DP_OP_423J2_125_3477_n359), .A2(
        DP_OP_423J2_125_3477_n494), .Y(DP_OP_423J2_125_3477_n97) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U113 ( .A1(DP_OP_423J2_125_3477_n494), .A2(
        DP_OP_423J2_125_3477_n359), .Y(DP_OP_423J2_125_3477_n96) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U105 ( .A1(DP_OP_423J2_125_3477_n265), .A2(
        DP_OP_423J2_125_3477_n358), .Y(DP_OP_423J2_125_3477_n91) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U104 ( .A1(DP_OP_423J2_125_3477_n358), .A2(
        DP_OP_423J2_125_3477_n265), .Y(DP_OP_423J2_125_3477_n90) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U97 ( .A1(DP_OP_423J2_125_3477_n219), .A2(
        DP_OP_423J2_125_3477_n264), .Y(DP_OP_423J2_125_3477_n86) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U96 ( .A1(DP_OP_423J2_125_3477_n264), .A2(
        DP_OP_423J2_125_3477_n219), .Y(DP_OP_423J2_125_3477_n85) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U92 ( .A1(DP_OP_423J2_125_3477_n85), .A2(
        DP_OP_423J2_125_3477_n90), .Y(DP_OP_423J2_125_3477_n83) );
  AOI21X1_HVT DP_OP_423J2_125_3477_U91 ( .A1(DP_OP_423J2_125_3477_n92), .A2(
        DP_OP_423J2_125_3477_n83), .A3(DP_OP_423J2_125_3477_n84), .Y(
        DP_OP_423J2_125_3477_n82) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U89 ( .A1(DP_OP_423J2_125_3477_n197), .A2(
        DP_OP_423J2_125_3477_n218), .Y(DP_OP_423J2_125_3477_n81) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U88 ( .A1(DP_OP_423J2_125_3477_n218), .A2(
        DP_OP_423J2_125_3477_n197), .Y(DP_OP_423J2_125_3477_n80) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U83 ( .A1(DP_OP_423J2_125_3477_n196), .A2(
        DP_OP_423J2_125_3477_n187), .Y(DP_OP_423J2_125_3477_n78) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U82 ( .A1(DP_OP_423J2_125_3477_n187), .A2(
        DP_OP_423J2_125_3477_n196), .Y(DP_OP_423J2_125_3477_n77) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U78 ( .A1(DP_OP_423J2_125_3477_n77), .A2(
        DP_OP_423J2_125_3477_n80), .Y(DP_OP_423J2_125_3477_n75) );
  AOI21X1_HVT DP_OP_423J2_125_3477_U77 ( .A1(DP_OP_423J2_125_3477_n84), .A2(
        DP_OP_423J2_125_3477_n75), .A3(DP_OP_423J2_125_3477_n76), .Y(
        DP_OP_423J2_125_3477_n74) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U76 ( .A1(DP_OP_423J2_125_3477_n83), .A2(
        DP_OP_423J2_125_3477_n75), .Y(DP_OP_423J2_125_3477_n73) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U72 ( .A1(DP_OP_423J2_125_3477_n186), .A2(
        DP_OP_423J2_125_3477_n181), .Y(DP_OP_423J2_125_3477_n66) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U62 ( .A1(DP_OP_423J2_125_3477_n180), .A2(
        DP_OP_423J2_125_3477_n179), .Y(DP_OP_423J2_125_3477_n63) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U61 ( .A1(DP_OP_423J2_125_3477_n179), .A2(
        DP_OP_423J2_125_3477_n180), .Y(DP_OP_423J2_125_3477_n62) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U54 ( .A1(DP_OP_423J2_125_3477_n178), .A2(
        DP_OP_423J2_125_3477_n177), .Y(DP_OP_423J2_125_3477_n58) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U53 ( .A1(DP_OP_423J2_125_3477_n177), .A2(
        DP_OP_423J2_125_3477_n178), .Y(DP_OP_423J2_125_3477_n57) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U49 ( .A1(DP_OP_423J2_125_3477_n57), .A2(
        DP_OP_423J2_125_3477_n62), .Y(DP_OP_423J2_125_3477_n55) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U47 ( .A1(DP_OP_423J2_125_3477_n67), .A2(
        DP_OP_423J2_125_3477_n55), .Y(DP_OP_423J2_125_3477_n53) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U44 ( .A1(DP_OP_423J2_125_3477_n175), .A2(
        DP_OP_423J2_125_3477_n176), .Y(DP_OP_423J2_125_3477_n51) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U43 ( .A1(DP_OP_423J2_125_3477_n176), .A2(
        DP_OP_423J2_125_3477_n175), .Y(DP_OP_423J2_125_3477_n50) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U39 ( .A1(DP_OP_423J2_125_3477_n50), .A2(
        DP_OP_423J2_125_3477_n53), .Y(DP_OP_423J2_125_3477_n48) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U34 ( .A1(DP_OP_423J2_125_3477_n173), .A2(
        DP_OP_423J2_125_3477_n174), .Y(DP_OP_423J2_125_3477_n44) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U27 ( .A1(DP_OP_423J2_125_3477_n48), .A2(
        DP_OP_423J2_125_3477_n43), .Y(DP_OP_423J2_125_3477_n39) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U24 ( .A1(DP_OP_423J2_125_3477_n171), .A2(
        DP_OP_423J2_125_3477_n172), .Y(DP_OP_423J2_125_3477_n37) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U23 ( .A1(DP_OP_423J2_125_3477_n172), .A2(
        DP_OP_423J2_125_3477_n171), .Y(DP_OP_423J2_125_3477_n36) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U19 ( .A1(DP_OP_423J2_125_3477_n36), .A2(
        DP_OP_423J2_125_3477_n39), .Y(DP_OP_423J2_125_3477_n34) );
  FADDX1_HVT DP_OP_423J2_125_3477_U15 ( .A(DP_OP_423J2_125_3477_n170), .B(
        DP_OP_423J2_125_3477_n169), .CI(DP_OP_423J2_125_3477_n33), .CO(
        DP_OP_423J2_125_3477_n32), .S(n_conv2_sum_b[20]) );
  FADDX1_HVT DP_OP_423J2_125_3477_U14 ( .A(DP_OP_423J2_125_3477_n168), .B(
        DP_OP_423J2_125_3477_n167), .CI(DP_OP_423J2_125_3477_n32), .CO(
        DP_OP_423J2_125_3477_n31), .S(n_conv2_sum_b[21]) );
  FADDX1_HVT DP_OP_423J2_125_3477_U13 ( .A(DP_OP_423J2_125_3477_n166), .B(
        DP_OP_423J2_125_3477_n165), .CI(DP_OP_423J2_125_3477_n31), .CO(
        DP_OP_423J2_125_3477_n30), .S(n_conv2_sum_b[22]) );
  FADDX1_HVT DP_OP_423J2_125_3477_U12 ( .A(DP_OP_423J2_125_3477_n164), .B(
        DP_OP_423J2_125_3477_n163), .CI(DP_OP_423J2_125_3477_n30), .CO(
        DP_OP_423J2_125_3477_n29), .S(n_conv2_sum_b[23]) );
  FADDX1_HVT DP_OP_423J2_125_3477_U11 ( .A(DP_OP_423J2_125_3477_n162), .B(
        DP_OP_423J2_125_3477_n161), .CI(DP_OP_423J2_125_3477_n29), .CO(
        DP_OP_423J2_125_3477_n28), .S(n_conv2_sum_b[24]) );
  FADDX1_HVT DP_OP_423J2_125_3477_U10 ( .A(DP_OP_423J2_125_3477_n160), .B(
        DP_OP_423J2_125_3477_n159), .CI(DP_OP_423J2_125_3477_n28), .CO(
        DP_OP_423J2_125_3477_n27), .S(n_conv2_sum_b[25]) );
  FADDX1_HVT DP_OP_423J2_125_3477_U9 ( .A(DP_OP_423J2_125_3477_n158), .B(
        DP_OP_423J2_125_3477_n157), .CI(DP_OP_423J2_125_3477_n27), .CO(
        DP_OP_423J2_125_3477_n26), .S(n_conv2_sum_b[26]) );
  FADDX1_HVT DP_OP_423J2_125_3477_U8 ( .A(DP_OP_423J2_125_3477_n156), .B(
        DP_OP_423J2_125_3477_n155), .CI(DP_OP_423J2_125_3477_n26), .CO(
        DP_OP_423J2_125_3477_n25), .S(n_conv2_sum_b[27]) );
  FADDX1_HVT DP_OP_423J2_125_3477_U7 ( .A(DP_OP_423J2_125_3477_n154), .B(
        DP_OP_423J2_125_3477_n153), .CI(DP_OP_423J2_125_3477_n25), .CO(
        DP_OP_423J2_125_3477_n24), .S(n_conv2_sum_b[28]) );
  FADDX1_HVT DP_OP_423J2_125_3477_U6 ( .A(DP_OP_423J2_125_3477_n152), .B(
        DP_OP_423J2_125_3477_n151), .CI(DP_OP_423J2_125_3477_n24), .CO(
        DP_OP_423J2_125_3477_n23), .S(n_conv2_sum_b[29]) );
  FADDX1_HVT DP_OP_423J2_125_3477_U5 ( .A(DP_OP_423J2_125_3477_n150), .B(
        DP_OP_423J2_125_3477_n149), .CI(DP_OP_423J2_125_3477_n23), .CO(
        DP_OP_423J2_125_3477_n22), .S(n_conv2_sum_b[30]) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1955 ( .A1(DP_OP_424J2_126_3477_n1988), 
        .A2(DP_OP_422J2_124_3477_n2742), .Y(DP_OP_425J2_127_3477_n2725) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1337 ( .A1(DP_OP_422J2_124_3477_n2651), 
        .A2(DP_OP_422J2_124_3477_n2128), .Y(DP_OP_423J2_125_3477_n2111) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1195 ( .A1(DP_OP_422J2_124_3477_n2869), 
        .A2(DP_OP_424J2_126_3477_n1995), .Y(DP_OP_424J2_126_3477_n1968) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1636 ( .A1(DP_OP_422J2_124_3477_n2298), 
        .A2(DP_OP_423J2_125_3477_n2431), .Y(DP_OP_423J2_125_3477_n2410) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1759 ( .A1(DP_OP_424J2_126_3477_n2471), 
        .A2(DP_OP_423J2_125_3477_n2562), .Y(DP_OP_423J2_125_3477_n2533) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1767 ( .A1(DP_OP_424J2_126_3477_n2561), 
        .A2(DP_OP_425J2_127_3477_n2564), .Y(DP_OP_424J2_126_3477_n2537) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1001 ( .A1(n386), .A2(
        DP_OP_424J2_126_3477_n2), .Y(DP_OP_423J2_125_3477_n1775) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2119 ( .A1(DP_OP_425J2_127_3477_n1860), 
        .A2(DP_OP_423J2_125_3477_n2911), .Y(DP_OP_424J2_126_3477_n2889) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1429 ( .A1(DP_OP_422J2_124_3477_n2649), 
        .A2(DP_OP_425J2_127_3477_n2217), .Y(DP_OP_424J2_126_3477_n2202) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1825 ( .A1(DP_OP_422J2_124_3477_n2033), 
        .A2(DP_OP_424J2_126_3477_n2610), .Y(DP_OP_424J2_126_3477_n2595) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1335 ( .A1(DP_OP_423J2_125_3477_n2117), 
        .A2(DP_OP_425J2_127_3477_n2129), .Y(DP_OP_423J2_125_3477_n2109) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2074 ( .A1(DP_OP_422J2_124_3477_n2868), 
        .A2(DP_OP_422J2_124_3477_n2872), .Y(DP_OP_422J2_124_3477_n2844) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1339 ( .A1(DP_OP_425J2_127_3477_n2120), 
        .A2(DP_OP_425J2_127_3477_n2129), .Y(DP_OP_425J2_127_3477_n2112) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1080 ( .A1(DP_OP_422J2_124_3477_n1861), 
        .A2(DP_OP_422J2_124_3477_n1865), .Y(DP_OP_422J2_124_3477_n1853) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1193 ( .A1(DP_OP_425J2_127_3477_n1990), 
        .A2(DP_OP_425J2_127_3477_n1995), .Y(DP_OP_425J2_127_3477_n1966) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2117 ( .A1(DP_OP_425J2_127_3477_n1858), 
        .A2(DP_OP_422J2_124_3477_n2916), .Y(DP_OP_424J2_126_3477_n2887) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1011 ( .A1(n388), .A2(n337), .Y(
        DP_OP_422J2_124_3477_n1784) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2115 ( .A1(DP_OP_425J2_127_3477_n2909), 
        .A2(DP_OP_425J2_127_3477_n2916), .Y(DP_OP_425J2_127_3477_n2885) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2069 ( .A1(DP_OP_423J2_125_3477_n2864), 
        .A2(DP_OP_423J2_125_3477_n2867), .Y(DP_OP_423J2_125_3477_n2840) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1868 ( .A1(DP_OP_422J2_124_3477_n2648), 
        .A2(DP_OP_422J2_124_3477_n2656), .Y(DP_OP_422J2_124_3477_n2640) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1951 ( .A1(DP_OP_423J2_125_3477_n2730), 
        .A2(DP_OP_423J2_125_3477_n2737), .Y(DP_OP_423J2_125_3477_n2722) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1344 ( .A1(DP_OP_422J2_124_3477_n2124), 
        .A2(DP_OP_422J2_124_3477_n2128), .Y(DP_OP_422J2_124_3477_n2116) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2118 ( .A1(DP_OP_422J2_124_3477_n2912), 
        .A2(DP_OP_422J2_124_3477_n2916), .Y(DP_OP_422J2_124_3477_n2888) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1333 ( .A1(DP_OP_423J2_125_3477_n2115), 
        .A2(DP_OP_424J2_126_3477_n2129), .Y(DP_OP_423J2_125_3477_n2107) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1378 ( .A1(DP_OP_423J2_125_3477_n2074), 
        .A2(DP_OP_422J2_124_3477_n2171), .Y(DP_OP_424J2_126_3477_n2151) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1339 ( .A1(DP_OP_425J2_127_3477_n2252), 
        .A2(DP_OP_422J2_124_3477_n2128), .Y(DP_OP_422J2_124_3477_n2111) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1195 ( .A1(DP_OP_423J2_125_3477_n2732), 
        .A2(DP_OP_422J2_124_3477_n1995), .Y(DP_OP_422J2_124_3477_n1968) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1071 ( .A1(DP_OP_423J2_125_3477_n1853), 
        .A2(DP_OP_423J2_125_3477_n1860), .Y(DP_OP_423J2_125_3477_n1845) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1863 ( .A1(DP_OP_423J2_125_3477_n2645), 
        .A2(DP_OP_422J2_124_3477_n2656), .Y(DP_OP_423J2_125_3477_n2637) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1007 ( .A1(n277), .A2(
        DP_OP_425J2_127_3477_n2), .Y(DP_OP_422J2_124_3477_n1780) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1869 ( .A1(DP_OP_425J2_127_3477_n2122), 
        .A2(DP_OP_424J2_126_3477_n2654), .Y(DP_OP_424J2_126_3477_n2639) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1341 ( .A1(DP_OP_422J2_124_3477_n2121), 
        .A2(DP_OP_422J2_124_3477_n2128), .Y(DP_OP_422J2_124_3477_n2113) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1423 ( .A1(DP_OP_423J2_125_3477_n2205), 
        .A2(DP_OP_423J2_125_3477_n2212), .Y(DP_OP_423J2_125_3477_n2197) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1819 ( .A1(DP_OP_423J2_125_3477_n2601), 
        .A2(DP_OP_425J2_127_3477_n2610), .Y(DP_OP_423J2_125_3477_n2593) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2111 ( .A1(DP_OP_423J2_125_3477_n2906), 
        .A2(DP_OP_423J2_125_3477_n2911), .Y(DP_OP_423J2_125_3477_n2882) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1765 ( .A1(DP_OP_425J2_127_3477_n2427), 
        .A2(DP_OP_422J2_124_3477_n2566), .Y(DP_OP_422J2_124_3477_n2537) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1696 ( .A1(DP_OP_422J2_124_3477_n2476), 
        .A2(DP_OP_422J2_124_3477_n2480), .Y(DP_OP_422J2_124_3477_n2468) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1761 ( .A1(DP_OP_423J2_125_3477_n2559), 
        .A2(DP_OP_423J2_125_3477_n2562), .Y(DP_OP_423J2_125_3477_n2535) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2113 ( .A1(DP_OP_423J2_125_3477_n2908), 
        .A2(DP_OP_423J2_125_3477_n2911), .Y(DP_OP_423J2_125_3477_n2884) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1370 ( .A1(DP_OP_423J2_125_3477_n2160), 
        .A2(DP_OP_423J2_125_3477_n2167), .Y(DP_OP_423J2_125_3477_n2144) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1077 ( .A1(DP_OP_424J2_126_3477_n1858), 
        .A2(DP_OP_424J2_126_3477_n1865), .Y(DP_OP_424J2_126_3477_n1850) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1872 ( .A1(DP_OP_422J2_124_3477_n2652), 
        .A2(DP_OP_422J2_124_3477_n2656), .Y(DP_OP_422J2_124_3477_n2644) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1766 ( .A1(DP_OP_422J2_124_3477_n2562), 
        .A2(DP_OP_422J2_124_3477_n2566), .Y(DP_OP_422J2_124_3477_n2538) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1960 ( .A1(DP_OP_423J2_125_3477_n2032), 
        .A2(DP_OP_422J2_124_3477_n2742), .Y(DP_OP_422J2_124_3477_n2730) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2073 ( .A1(DP_OP_424J2_126_3477_n2867), 
        .A2(DP_OP_422J2_124_3477_n2872), .Y(DP_OP_424J2_126_3477_n2843) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1555 ( .A1(DP_OP_422J2_124_3477_n2429), 
        .A2(DP_OP_423J2_125_3477_n2344), .Y(DP_OP_423J2_125_3477_n2329) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1428 ( .A1(DP_OP_422J2_124_3477_n2208), 
        .A2(DP_OP_422J2_124_3477_n2216), .Y(DP_OP_422J2_124_3477_n2200) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1372 ( .A1(DP_OP_425J2_127_3477_n2472), 
        .A2(DP_OP_423J2_125_3477_n2167), .Y(DP_OP_423J2_125_3477_n2146) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2117 ( .A1(DP_OP_425J2_127_3477_n2779), 
        .A2(DP_OP_422J2_124_3477_n2916), .Y(DP_OP_422J2_124_3477_n2887) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1763 ( .A1(DP_OP_425J2_127_3477_n2557), 
        .A2(DP_OP_425J2_127_3477_n2564), .Y(DP_OP_425J2_127_3477_n2533) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1775 ( .A1(DP_OP_424J2_126_3477_n2471), 
        .A2(DP_OP_424J2_126_3477_n2566), .Y(DP_OP_423J2_125_3477_n2549) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1189 ( .A1(DP_OP_422J2_124_3477_n2781), 
        .A2(DP_OP_424J2_126_3477_n1995), .Y(DP_OP_423J2_125_3477_n1963) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1015 ( .A1(n279), .A2(
        DP_OP_423J2_125_3477_n2), .Y(DP_OP_422J2_124_3477_n1788) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1649 ( .A1(DP_OP_425J2_127_3477_n2342), 
        .A2(DP_OP_423J2_125_3477_n2432), .Y(DP_OP_424J2_126_3477_n2419) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1779 ( .A1(DP_OP_422J2_124_3477_n2559), 
        .A2(DP_OP_422J2_124_3477_n2568), .Y(DP_OP_422J2_124_3477_n2551) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1691 ( .A1(DP_OP_422J2_124_3477_n2163), 
        .A2(DP_OP_424J2_126_3477_n2478), .Y(DP_OP_424J2_126_3477_n2461) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1957 ( .A1(DP_OP_424J2_126_3477_n2735), 
        .A2(DP_OP_424J2_126_3477_n2742), .Y(DP_OP_424J2_126_3477_n2727) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1765 ( .A1(DP_OP_424J2_126_3477_n2559), 
        .A2(DP_OP_423J2_125_3477_n2562), .Y(DP_OP_424J2_126_3477_n2535) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1561 ( .A1(DP_OP_424J2_126_3477_n2342), 
        .A2(DP_OP_424J2_126_3477_n2349), .Y(DP_OP_424J2_126_3477_n2334) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1692 ( .A1(DP_OP_422J2_124_3477_n2472), 
        .A2(DP_OP_422J2_124_3477_n2480), .Y(DP_OP_422J2_124_3477_n2464) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1193 ( .A1(DP_OP_423J2_125_3477_n1897), 
        .A2(DP_OP_424J2_126_3477_n1995), .Y(DP_OP_424J2_126_3477_n1966) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1828 ( .A1(DP_OP_422J2_124_3477_n2608), 
        .A2(DP_OP_422J2_124_3477_n2612), .Y(DP_OP_422J2_124_3477_n2600) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U985 ( .A1(n321), .A2(
        DP_OP_423J2_125_3477_n2), .Y(DP_OP_425J2_127_3477_n153) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1640 ( .A1(DP_OP_425J2_127_3477_n2341), 
        .A2(DP_OP_422J2_124_3477_n2435), .Y(DP_OP_424J2_126_3477_n2410) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1187 ( .A1(DP_OP_423J2_125_3477_n1985), 
        .A2(DP_OP_424J2_126_3477_n1995), .Y(DP_OP_423J2_125_3477_n1961) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2071 ( .A1(DP_OP_425J2_127_3477_n2865), 
        .A2(DP_OP_425J2_127_3477_n2872), .Y(DP_OP_425J2_127_3477_n2841) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1191 ( .A1(DP_OP_424J2_126_3477_n2777), 
        .A2(DP_OP_425J2_127_3477_n1995), .Y(DP_OP_425J2_127_3477_n1964) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1076 ( .A1(DP_OP_425J2_127_3477_n1989), 
        .A2(DP_OP_422J2_124_3477_n1865), .Y(DP_OP_422J2_124_3477_n1849) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1642 ( .A1(DP_OP_424J2_126_3477_n2428), 
        .A2(DP_OP_423J2_125_3477_n2431), .Y(DP_OP_424J2_126_3477_n2412) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1341 ( .A1(DP_OP_423J2_125_3477_n2029), 
        .A2(DP_OP_424J2_126_3477_n2129), .Y(DP_OP_424J2_126_3477_n2114) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1008 ( .A1(n265), .A2(
        DP_OP_424J2_126_3477_n2), .Y(DP_OP_425J2_127_3477_n1781) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1641 ( .A1(DP_OP_422J2_124_3477_n2429), 
        .A2(DP_OP_422J2_124_3477_n2435), .Y(DP_OP_422J2_124_3477_n2413) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1780 ( .A1(DP_OP_422J2_124_3477_n2560), 
        .A2(DP_OP_422J2_124_3477_n2568), .Y(DP_OP_422J2_124_3477_n2552) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1376 ( .A1(DP_OP_422J2_124_3477_n2692), 
        .A2(DP_OP_423J2_125_3477_n2167), .Y(DP_OP_424J2_126_3477_n2149) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1767 ( .A1(DP_OP_422J2_124_3477_n2563), 
        .A2(DP_OP_422J2_124_3477_n2566), .Y(DP_OP_422J2_124_3477_n2539) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2075 ( .A1(DP_OP_422J2_124_3477_n2869), 
        .A2(DP_OP_422J2_124_3477_n2872), .Y(DP_OP_422J2_124_3477_n2845) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1648 ( .A1(DP_OP_422J2_124_3477_n2428), 
        .A2(DP_OP_422J2_124_3477_n2436), .Y(DP_OP_422J2_124_3477_n2420) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1339 ( .A1(DP_OP_424J2_126_3477_n2120), 
        .A2(DP_OP_424J2_126_3477_n2129), .Y(DP_OP_424J2_126_3477_n2112) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1069 ( .A1(DP_OP_425J2_127_3477_n2777), 
        .A2(DP_OP_423J2_125_3477_n1860), .Y(DP_OP_423J2_125_3477_n1843) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1781 ( .A1(DP_OP_424J2_126_3477_n2559), 
        .A2(DP_OP_424J2_126_3477_n2566), .Y(DP_OP_424J2_126_3477_n2551) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1377 ( .A1(DP_OP_422J2_124_3477_n2165), 
        .A2(DP_OP_422J2_124_3477_n2171), .Y(DP_OP_422J2_124_3477_n2149) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1634 ( .A1(DP_OP_423J2_125_3477_n2424), 
        .A2(DP_OP_423J2_125_3477_n2431), .Y(DP_OP_423J2_125_3477_n2408) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1341 ( .A1(DP_OP_425J2_127_3477_n2122), 
        .A2(DP_OP_425J2_127_3477_n2129), .Y(DP_OP_425J2_127_3477_n2114) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1694 ( .A1(DP_OP_423J2_125_3477_n2294), 
        .A2(DP_OP_422J2_124_3477_n2480), .Y(DP_OP_422J2_124_3477_n2466) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1954 ( .A1(DP_OP_423J2_125_3477_n2733), 
        .A2(DP_OP_423J2_125_3477_n2737), .Y(DP_OP_423J2_125_3477_n2725) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1375 ( .A1(DP_OP_424J2_126_3477_n2164), 
        .A2(DP_OP_422J2_124_3477_n2171), .Y(DP_OP_424J2_126_3477_n2148) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1074 ( .A1(DP_OP_423J2_125_3477_n1856), 
        .A2(DP_OP_423J2_125_3477_n1860), .Y(DP_OP_423J2_125_3477_n1848) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1783 ( .A1(DP_OP_422J2_124_3477_n2563), 
        .A2(DP_OP_422J2_124_3477_n2568), .Y(DP_OP_422J2_124_3477_n2555) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1009 ( .A1(n395), .A2(
        DP_OP_423J2_125_3477_n2), .Y(DP_OP_424J2_126_3477_n1782) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2119 ( .A1(DP_OP_425J2_127_3477_n2913), 
        .A2(DP_OP_425J2_127_3477_n2916), .Y(DP_OP_425J2_127_3477_n2889) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2115 ( .A1(DP_OP_422J2_124_3477_n2909), 
        .A2(DP_OP_422J2_124_3477_n2916), .Y(DP_OP_422J2_124_3477_n2885) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2072 ( .A1(DP_OP_424J2_126_3477_n1857), 
        .A2(DP_OP_425J2_127_3477_n2872), .Y(DP_OP_425J2_127_3477_n2842) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1763 ( .A1(DP_OP_422J2_124_3477_n2559), 
        .A2(DP_OP_422J2_124_3477_n2566), .Y(DP_OP_422J2_124_3477_n2535) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1338 ( .A1(DP_OP_425J2_127_3477_n2518), 
        .A2(DP_OP_424J2_126_3477_n2129), .Y(DP_OP_423J2_125_3477_n2112) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1644 ( .A1(DP_OP_422J2_124_3477_n2432), 
        .A2(DP_OP_422J2_124_3477_n2435), .Y(DP_OP_422J2_124_3477_n2416) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1558 ( .A1(DP_OP_422J2_124_3477_n2432), 
        .A2(DP_OP_423J2_125_3477_n2344), .Y(DP_OP_423J2_125_3477_n2332) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1866 ( .A1(DP_OP_423J2_125_3477_n2648), 
        .A2(DP_OP_422J2_124_3477_n2656), .Y(DP_OP_423J2_125_3477_n2640) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2072 ( .A1(DP_OP_425J2_127_3477_n1901), 
        .A2(DP_OP_423J2_125_3477_n2867), .Y(DP_OP_424J2_126_3477_n2842) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1822 ( .A1(DP_OP_423J2_125_3477_n2604), 
        .A2(DP_OP_425J2_127_3477_n2610), .Y(DP_OP_423J2_125_3477_n2596) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1191 ( .A1(DP_OP_422J2_124_3477_n1988), 
        .A2(DP_OP_422J2_124_3477_n1995), .Y(DP_OP_422J2_124_3477_n1964) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1639 ( .A1(DP_OP_425J2_127_3477_n2340), 
        .A2(DP_OP_423J2_125_3477_n2431), .Y(DP_OP_424J2_126_3477_n2409) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2116 ( .A1(DP_OP_424J2_126_3477_n2910), 
        .A2(DP_OP_423J2_125_3477_n2911), .Y(DP_OP_424J2_126_3477_n2886) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1690 ( .A1(DP_OP_423J2_125_3477_n2472), 
        .A2(DP_OP_423J2_125_3477_n2476), .Y(DP_OP_423J2_125_3477_n2464) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2075 ( .A1(DP_OP_425J2_127_3477_n2869), 
        .A2(DP_OP_425J2_127_3477_n2872), .Y(DP_OP_425J2_127_3477_n2845) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2071 ( .A1(DP_OP_422J2_124_3477_n2865), 
        .A2(DP_OP_422J2_124_3477_n2872), .Y(DP_OP_422J2_124_3477_n2841) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1195 ( .A1(DP_OP_425J2_127_3477_n1992), 
        .A2(DP_OP_425J2_127_3477_n1995), .Y(DP_OP_425J2_127_3477_n1968) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1778 ( .A1(DP_OP_422J2_124_3477_n2168), 
        .A2(DP_OP_425J2_127_3477_n2566), .Y(DP_OP_423J2_125_3477_n2552) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1646 ( .A1(DP_OP_423J2_125_3477_n2428), 
        .A2(DP_OP_423J2_125_3477_n2432), .Y(DP_OP_423J2_125_3477_n2420) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1426 ( .A1(DP_OP_425J2_127_3477_n2430), 
        .A2(DP_OP_423J2_125_3477_n2212), .Y(DP_OP_423J2_125_3477_n2200) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1781 ( .A1(DP_OP_425J2_127_3477_n2559), 
        .A2(DP_OP_425J2_127_3477_n2566), .Y(DP_OP_425J2_127_3477_n2551) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1777 ( .A1(DP_OP_423J2_125_3477_n2559), 
        .A2(DP_OP_422J2_124_3477_n2568), .Y(DP_OP_423J2_125_3477_n2551) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1953 ( .A1(DP_OP_423J2_125_3477_n2732), 
        .A2(DP_OP_423J2_125_3477_n2737), .Y(DP_OP_423J2_125_3477_n2724) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1642 ( .A1(DP_OP_425J2_127_3477_n2428), 
        .A2(DP_OP_425J2_127_3477_n2433), .Y(DP_OP_425J2_127_3477_n2412) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1865 ( .A1(DP_OP_423J2_125_3477_n2647), 
        .A2(DP_OP_425J2_127_3477_n2654), .Y(DP_OP_423J2_125_3477_n2639) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1073 ( .A1(DP_OP_424J2_126_3477_n1948), 
        .A2(DP_OP_423J2_125_3477_n1860), .Y(DP_OP_423J2_125_3477_n1847) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1958 ( .A1(DP_OP_422J2_124_3477_n2736), 
        .A2(DP_OP_422J2_124_3477_n2742), .Y(DP_OP_422J2_124_3477_n2728) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1186 ( .A1(DP_OP_425J2_127_3477_n2646), 
        .A2(DP_OP_422J2_124_3477_n1995), .Y(DP_OP_423J2_125_3477_n1960) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1430 ( .A1(DP_OP_422J2_124_3477_n2210), 
        .A2(DP_OP_422J2_124_3477_n2216), .Y(DP_OP_422J2_124_3477_n2202) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1776 ( .A1(DP_OP_423J2_125_3477_n2558), 
        .A2(DP_OP_424J2_126_3477_n2566), .Y(DP_OP_423J2_125_3477_n2550) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1952 ( .A1(DP_OP_423J2_125_3477_n2731), 
        .A2(DP_OP_423J2_125_3477_n2737), .Y(DP_OP_423J2_125_3477_n2723) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1072 ( .A1(DP_OP_425J2_127_3477_n2780), 
        .A2(DP_OP_423J2_125_3477_n1860), .Y(DP_OP_423J2_125_3477_n1846) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1079 ( .A1(DP_OP_425J2_127_3477_n1860), 
        .A2(DP_OP_422J2_124_3477_n1865), .Y(DP_OP_425J2_127_3477_n1852) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1424 ( .A1(DP_OP_425J2_127_3477_n2428), 
        .A2(DP_OP_423J2_125_3477_n2212), .Y(DP_OP_423J2_125_3477_n2198) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1688 ( .A1(DP_OP_423J2_125_3477_n2470), 
        .A2(DP_OP_423J2_125_3477_n2476), .Y(DP_OP_423J2_125_3477_n2462) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1637 ( .A1(DP_OP_422J2_124_3477_n2299), 
        .A2(DP_OP_423J2_125_3477_n2431), .Y(DP_OP_423J2_125_3477_n2411) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1374 ( .A1(DP_OP_423J2_125_3477_n2164), 
        .A2(DP_OP_423J2_125_3477_n2167), .Y(DP_OP_423J2_125_3477_n2148) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1692 ( .A1(DP_OP_425J2_127_3477_n2297), 
        .A2(DP_OP_424J2_126_3477_n2478), .Y(DP_OP_424J2_126_3477_n2462) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1193 ( .A1(DP_OP_423J2_125_3477_n2730), 
        .A2(DP_OP_422J2_124_3477_n1995), .Y(DP_OP_422J2_124_3477_n1966) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1194 ( .A1(DP_OP_423J2_125_3477_n1898), 
        .A2(DP_OP_424J2_126_3477_n1995), .Y(DP_OP_424J2_126_3477_n1967) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1824 ( .A1(DP_OP_422J2_124_3477_n2032), 
        .A2(DP_OP_424J2_126_3477_n2610), .Y(DP_OP_424J2_126_3477_n2594) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1956 ( .A1(DP_OP_424J2_126_3477_n2734), 
        .A2(DP_OP_424J2_126_3477_n2742), .Y(DP_OP_424J2_126_3477_n2726) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U992 ( .A1(n303), .A2(n338), .Y(
        DP_OP_425J2_127_3477_n167) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1560 ( .A1(DP_OP_424J2_126_3477_n2341), 
        .A2(DP_OP_424J2_126_3477_n2349), .Y(DP_OP_424J2_126_3477_n2333) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1641 ( .A1(DP_OP_425J2_127_3477_n2342), 
        .A2(DP_OP_423J2_125_3477_n2431), .Y(DP_OP_424J2_126_3477_n2411) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2118 ( .A1(DP_OP_424J2_126_3477_n2912), 
        .A2(DP_OP_423J2_125_3477_n2911), .Y(DP_OP_424J2_126_3477_n2888) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1377 ( .A1(DP_OP_425J2_127_3477_n2559), 
        .A2(DP_OP_425J2_127_3477_n2172), .Y(DP_OP_424J2_126_3477_n2150) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1821 ( .A1(DP_OP_423J2_125_3477_n2603), 
        .A2(DP_OP_424J2_126_3477_n2610), .Y(DP_OP_423J2_125_3477_n2595) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1076 ( .A1(DP_OP_424J2_126_3477_n1857), 
        .A2(DP_OP_424J2_126_3477_n1865), .Y(DP_OP_424J2_126_3477_n1849) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1825 ( .A1(DP_OP_423J2_125_3477_n2029), 
        .A2(DP_OP_425J2_127_3477_n2610), .Y(DP_OP_425J2_127_3477_n2595) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U990 ( .A1(n329), .A2(
        DP_OP_424J2_126_3477_n2), .Y(DP_OP_425J2_127_3477_n163) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1429 ( .A1(DP_OP_424J2_126_3477_n2559), 
        .A2(DP_OP_425J2_127_3477_n2217), .Y(DP_OP_425J2_127_3477_n2202) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1378 ( .A1(DP_OP_423J2_125_3477_n2690), 
        .A2(DP_OP_425J2_127_3477_n2172), .Y(DP_OP_425J2_127_3477_n2151) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U988 ( .A1(n317), .A2(n337), .Y(
        DP_OP_425J2_127_3477_n159) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U987 ( .A1(n325), .A2(
        DP_OP_425J2_127_3477_n2), .Y(DP_OP_425J2_127_3477_n157) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1561 ( .A1(DP_OP_425J2_127_3477_n2342), 
        .A2(DP_OP_425J2_127_3477_n2349), .Y(DP_OP_425J2_127_3477_n2334) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1425 ( .A1(DP_OP_425J2_127_3477_n2429), 
        .A2(DP_OP_423J2_125_3477_n2212), .Y(DP_OP_423J2_125_3477_n2199) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1557 ( .A1(DP_OP_423J2_125_3477_n2339), 
        .A2(DP_OP_423J2_125_3477_n2344), .Y(DP_OP_423J2_125_3477_n2331) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U985 ( .A1(n324), .A2(n337), .Y(
        DP_OP_423J2_125_3477_n160) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1645 ( .A1(DP_OP_422J2_124_3477_n2299), 
        .A2(DP_OP_423J2_125_3477_n2432), .Y(DP_OP_423J2_125_3477_n2419) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1192 ( .A1(DP_OP_425J2_127_3477_n2734), 
        .A2(DP_OP_424J2_126_3477_n1995), .Y(DP_OP_424J2_126_3477_n1965) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U984 ( .A1(n328), .A2(
        DP_OP_425J2_127_3477_n2), .Y(DP_OP_423J2_125_3477_n158) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U986 ( .A1(n327), .A2(n338), .Y(
        DP_OP_425J2_127_3477_n155) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U983 ( .A1(n319), .A2(n338), .Y(
        DP_OP_423J2_125_3477_n156) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1077 ( .A1(DP_OP_425J2_127_3477_n1858), 
        .A2(DP_OP_424J2_126_3477_n1865), .Y(DP_OP_425J2_127_3477_n1850) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1428 ( .A1(DP_OP_422J2_124_3477_n2648), 
        .A2(DP_OP_425J2_127_3477_n2217), .Y(DP_OP_424J2_126_3477_n2201) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1766 ( .A1(DP_OP_422J2_124_3477_n2078), 
        .A2(DP_OP_423J2_125_3477_n2562), .Y(DP_OP_424J2_126_3477_n2536) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1012 ( .A1(n267), .A2(n338), .Y(
        DP_OP_425J2_127_3477_n1785) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1693 ( .A1(DP_OP_423J2_125_3477_n2161), 
        .A2(DP_OP_424J2_126_3477_n2478), .Y(DP_OP_425J2_127_3477_n2463) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1689 ( .A1(DP_OP_423J2_125_3477_n2471), 
        .A2(DP_OP_423J2_125_3477_n2476), .Y(DP_OP_423J2_125_3477_n2463) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1004 ( .A1(n282), .A2(
        DP_OP_423J2_125_3477_n2), .Y(DP_OP_425J2_127_3477_n1777) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1648 ( .A1(DP_OP_425J2_127_3477_n2341), 
        .A2(DP_OP_425J2_127_3477_n2434), .Y(DP_OP_424J2_126_3477_n2418) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1868 ( .A1(DP_OP_422J2_124_3477_n1989), 
        .A2(DP_OP_424J2_126_3477_n2654), .Y(DP_OP_424J2_126_3477_n2638) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1867 ( .A1(DP_OP_422J2_124_3477_n2647), 
        .A2(DP_OP_422J2_124_3477_n2656), .Y(DP_OP_422J2_124_3477_n2639) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1376 ( .A1(DP_OP_422J2_124_3477_n2164), 
        .A2(DP_OP_422J2_124_3477_n2171), .Y(DP_OP_422J2_124_3477_n2148) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1780 ( .A1(DP_OP_425J2_127_3477_n2209), 
        .A2(DP_OP_424J2_126_3477_n2566), .Y(DP_OP_424J2_126_3477_n2550) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1011 ( .A1(n389), .A2(
        DP_OP_424J2_126_3477_n2), .Y(DP_OP_424J2_126_3477_n1784) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1342 ( .A1(DP_OP_425J2_127_3477_n2255), 
        .A2(DP_OP_422J2_124_3477_n2128), .Y(DP_OP_422J2_124_3477_n2114) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1340 ( .A1(DP_OP_423J2_125_3477_n2028), 
        .A2(DP_OP_424J2_126_3477_n2129), .Y(DP_OP_424J2_126_3477_n2113) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1649 ( .A1(DP_OP_425J2_127_3477_n2427), 
        .A2(DP_OP_425J2_127_3477_n2434), .Y(DP_OP_425J2_127_3477_n2419) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2074 ( .A1(DP_OP_425J2_127_3477_n1903), 
        .A2(DP_OP_423J2_125_3477_n2867), .Y(DP_OP_424J2_126_3477_n2844) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2073 ( .A1(DP_OP_423J2_125_3477_n1897), 
        .A2(DP_OP_422J2_124_3477_n2872), .Y(DP_OP_422J2_124_3477_n2843) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1957 ( .A1(DP_OP_425J2_127_3477_n2735), 
        .A2(DP_OP_424J2_126_3477_n2742), .Y(DP_OP_425J2_127_3477_n2727) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1869 ( .A1(DP_OP_424J2_126_3477_n2078), 
        .A2(DP_OP_425J2_127_3477_n2654), .Y(DP_OP_425J2_127_3477_n2639) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1767 ( .A1(DP_OP_422J2_124_3477_n2695), 
        .A2(DP_OP_425J2_127_3477_n2564), .Y(DP_OP_425J2_127_3477_n2537) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1376 ( .A1(DP_OP_423J2_125_3477_n2688), 
        .A2(DP_OP_425J2_127_3477_n2172), .Y(DP_OP_425J2_127_3477_n2149) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1075 ( .A1(DP_OP_424J2_126_3477_n2909), 
        .A2(DP_OP_422J2_124_3477_n1865), .Y(DP_OP_425J2_127_3477_n1848) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1764 ( .A1(DP_OP_422J2_124_3477_n2560), 
        .A2(DP_OP_422J2_124_3477_n2566), .Y(DP_OP_422J2_124_3477_n2536) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1638 ( .A1(DP_OP_423J2_125_3477_n2428), 
        .A2(DP_OP_423J2_125_3477_n2431), .Y(DP_OP_423J2_125_3477_n2412) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1342 ( .A1(DP_OP_422J2_124_3477_n1991), 
        .A2(DP_OP_425J2_127_3477_n2129), .Y(DP_OP_425J2_127_3477_n2115) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1784 ( .A1(DP_OP_422J2_124_3477_n2696), 
        .A2(DP_OP_425J2_127_3477_n2566), .Y(DP_OP_425J2_127_3477_n2554) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1379 ( .A1(DP_OP_425J2_127_3477_n2168), 
        .A2(DP_OP_425J2_127_3477_n2172), .Y(DP_OP_425J2_127_3477_n2152) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1763 ( .A1(DP_OP_424J2_126_3477_n2557), 
        .A2(DP_OP_425J2_127_3477_n2564), .Y(DP_OP_424J2_126_3477_n2533) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1008 ( .A1(n375), .A2(
        DP_OP_423J2_125_3477_n2), .Y(DP_OP_424J2_126_3477_n1781) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1959 ( .A1(DP_OP_424J2_126_3477_n2737), 
        .A2(DP_OP_424J2_126_3477_n2742), .Y(DP_OP_424J2_126_3477_n2729) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1079 ( .A1(DP_OP_425J2_127_3477_n2869), 
        .A2(DP_OP_424J2_126_3477_n1865), .Y(DP_OP_424J2_126_3477_n1852) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1643 ( .A1(DP_OP_423J2_125_3477_n2339), 
        .A2(DP_OP_422J2_124_3477_n2435), .Y(DP_OP_422J2_124_3477_n2415) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2067 ( .A1(DP_OP_425J2_127_3477_n1990), 
        .A2(DP_OP_423J2_125_3477_n2867), .Y(DP_OP_423J2_125_3477_n2838) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2076 ( .A1(DP_OP_422J2_124_3477_n2870), 
        .A2(DP_OP_422J2_124_3477_n2872), .Y(DP_OP_422J2_124_3477_n2846) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1564 ( .A1(DP_OP_422J2_124_3477_n2344), 
        .A2(DP_OP_423J2_125_3477_n2344), .Y(DP_OP_422J2_124_3477_n2336) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1652 ( .A1(DP_OP_422J2_124_3477_n2432), 
        .A2(DP_OP_422J2_124_3477_n2436), .Y(DP_OP_422J2_124_3477_n2424) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1432 ( .A1(DP_OP_423J2_125_3477_n2516), 
        .A2(DP_OP_422J2_124_3477_n2216), .Y(DP_OP_422J2_124_3477_n2204) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1687 ( .A1(DP_OP_423J2_125_3477_n2469), 
        .A2(DP_OP_423J2_125_3477_n2476), .Y(DP_OP_423J2_125_3477_n2461) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1375 ( .A1(DP_OP_422J2_124_3477_n2163), 
        .A2(DP_OP_422J2_124_3477_n2171), .Y(DP_OP_422J2_124_3477_n2147) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1693 ( .A1(DP_OP_424J2_126_3477_n2471), 
        .A2(DP_OP_424J2_126_3477_n2478), .Y(DP_OP_424J2_126_3477_n2463) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1784 ( .A1(DP_OP_422J2_124_3477_n2564), 
        .A2(DP_OP_422J2_124_3477_n2568), .Y(DP_OP_422J2_124_3477_n2556) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2075 ( .A1(DP_OP_424J2_126_3477_n2869), 
        .A2(DP_OP_423J2_125_3477_n2867), .Y(DP_OP_424J2_126_3477_n2845) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1556 ( .A1(DP_OP_422J2_124_3477_n2430), 
        .A2(DP_OP_423J2_125_3477_n2344), .Y(DP_OP_423J2_125_3477_n2330) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1013 ( .A1(n391), .A2(n338), .Y(
        DP_OP_422J2_124_3477_n1786) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1650 ( .A1(DP_OP_422J2_124_3477_n2430), 
        .A2(DP_OP_422J2_124_3477_n2436), .Y(DP_OP_422J2_124_3477_n2422) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2114 ( .A1(DP_OP_423J2_125_3477_n2909), 
        .A2(DP_OP_423J2_125_3477_n2911), .Y(DP_OP_423J2_125_3477_n2885) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2070 ( .A1(DP_OP_423J2_125_3477_n2865), 
        .A2(DP_OP_423J2_125_3477_n2867), .Y(DP_OP_423J2_125_3477_n2841) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1762 ( .A1(DP_OP_422J2_124_3477_n2168), 
        .A2(DP_OP_423J2_125_3477_n2562), .Y(DP_OP_423J2_125_3477_n2536) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1644 ( .A1(DP_OP_422J2_124_3477_n2298), 
        .A2(DP_OP_423J2_125_3477_n2432), .Y(DP_OP_423J2_125_3477_n2418) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1336 ( .A1(DP_OP_424J2_126_3477_n2211), 
        .A2(DP_OP_425J2_127_3477_n2129), .Y(DP_OP_423J2_125_3477_n2110) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1078 ( .A1(DP_OP_422J2_124_3477_n1859), 
        .A2(DP_OP_422J2_124_3477_n1865), .Y(DP_OP_422J2_124_3477_n1851) );
  OR2X1_HVT DP_OP_422J2_124_3477_U984 ( .A1(n315), .A2(DP_OP_424J2_126_3477_n2), .Y(DP_OP_422J2_124_3477_n1773) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1640 ( .A1(DP_OP_423J2_125_3477_n2204), 
        .A2(DP_OP_425J2_127_3477_n2433), .Y(DP_OP_425J2_127_3477_n2410) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1864 ( .A1(DP_OP_423J2_125_3477_n2646), 
        .A2(DP_OP_422J2_124_3477_n2656), .Y(DP_OP_423J2_125_3477_n2638) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1190 ( .A1(DP_OP_422J2_124_3477_n2782), 
        .A2(DP_OP_424J2_126_3477_n1995), .Y(DP_OP_423J2_125_3477_n1964) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1820 ( .A1(DP_OP_423J2_125_3477_n2602), 
        .A2(DP_OP_425J2_127_3477_n2610), .Y(DP_OP_423J2_125_3477_n2594) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U997 ( .A1(n288), .A2(n338), .Y(
        DP_OP_423J2_125_3477_n1771) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2120 ( .A1(DP_OP_424J2_126_3477_n1949), 
        .A2(DP_OP_422J2_124_3477_n2916), .Y(DP_OP_422J2_124_3477_n2890) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1196 ( .A1(DP_OP_424J2_126_3477_n2650), 
        .A2(DP_OP_422J2_124_3477_n1995), .Y(DP_OP_422J2_124_3477_n1969) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1826 ( .A1(DP_OP_422J2_124_3477_n2606), 
        .A2(DP_OP_422J2_124_3477_n2612), .Y(DP_OP_422J2_124_3477_n2598) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2071 ( .A1(DP_OP_424J2_126_3477_n2865), 
        .A2(DP_OP_425J2_127_3477_n2872), .Y(DP_OP_424J2_126_3477_n2841) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2115 ( .A1(DP_OP_424J2_126_3477_n2909), 
        .A2(DP_OP_423J2_125_3477_n2911), .Y(DP_OP_424J2_126_3477_n2885) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1765 ( .A1(DP_OP_425J2_127_3477_n2559), 
        .A2(DP_OP_425J2_127_3477_n2564), .Y(DP_OP_425J2_127_3477_n2535) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2116 ( .A1(DP_OP_425J2_127_3477_n2778), 
        .A2(DP_OP_422J2_124_3477_n2916), .Y(DP_OP_422J2_124_3477_n2886) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1639 ( .A1(DP_OP_422J2_124_3477_n2427), 
        .A2(DP_OP_422J2_124_3477_n2435), .Y(DP_OP_422J2_124_3477_n2411) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2073 ( .A1(DP_OP_424J2_126_3477_n1858), 
        .A2(DP_OP_425J2_127_3477_n2872), .Y(DP_OP_425J2_127_3477_n2843) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1191 ( .A1(DP_OP_424J2_126_3477_n1988), 
        .A2(DP_OP_424J2_126_3477_n1995), .Y(DP_OP_424J2_126_3477_n1964) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1870 ( .A1(DP_OP_422J2_124_3477_n2650), 
        .A2(DP_OP_422J2_124_3477_n2656), .Y(DP_OP_422J2_124_3477_n2642) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1379 ( .A1(DP_OP_424J2_126_3477_n2168), 
        .A2(DP_OP_425J2_127_3477_n2172), .Y(DP_OP_424J2_126_3477_n2152) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1694 ( .A1(DP_OP_424J2_126_3477_n2472), 
        .A2(DP_OP_424J2_126_3477_n2478), .Y(DP_OP_424J2_126_3477_n2464) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1379 ( .A1(DP_OP_425J2_127_3477_n2300), 
        .A2(DP_OP_422J2_124_3477_n2171), .Y(DP_OP_422J2_124_3477_n2151) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1562 ( .A1(DP_OP_422J2_124_3477_n2342), 
        .A2(DP_OP_425J2_127_3477_n2349), .Y(DP_OP_422J2_124_3477_n2334) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1009 ( .A1(n392), .A2(
        DP_OP_425J2_127_3477_n2), .Y(DP_OP_422J2_124_3477_n1782) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2117 ( .A1(DP_OP_425J2_127_3477_n2911), 
        .A2(DP_OP_425J2_127_3477_n2916), .Y(DP_OP_425J2_127_3477_n2887) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1867 ( .A1(DP_OP_425J2_127_3477_n2120), 
        .A2(DP_OP_424J2_126_3477_n2654), .Y(DP_OP_424J2_126_3477_n2637) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2109 ( .A1(DP_OP_423J2_125_3477_n2904), 
        .A2(DP_OP_423J2_125_3477_n2911), .Y(DP_OP_423J2_125_3477_n2880) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1960 ( .A1(DP_OP_424J2_126_3477_n2738), 
        .A2(DP_OP_424J2_126_3477_n2742), .Y(DP_OP_424J2_126_3477_n2730) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1196 ( .A1(DP_OP_425J2_127_3477_n2738), 
        .A2(DP_OP_424J2_126_3477_n1995), .Y(DP_OP_424J2_126_3477_n1969) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1640 ( .A1(DP_OP_422J2_124_3477_n2428), 
        .A2(DP_OP_422J2_124_3477_n2435), .Y(DP_OP_422J2_124_3477_n2412) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2074 ( .A1(DP_OP_425J2_127_3477_n2868), 
        .A2(DP_OP_425J2_127_3477_n2872), .Y(DP_OP_425J2_127_3477_n2844) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1870 ( .A1(DP_OP_422J2_124_3477_n1991), 
        .A2(DP_OP_424J2_126_3477_n2654), .Y(DP_OP_424J2_126_3477_n2640) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1429 ( .A1(DP_OP_422J2_124_3477_n2209), 
        .A2(DP_OP_422J2_124_3477_n2216), .Y(DP_OP_422J2_124_3477_n2201) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1633 ( .A1(DP_OP_422J2_124_3477_n2295), 
        .A2(DP_OP_423J2_125_3477_n2431), .Y(DP_OP_423J2_125_3477_n2407) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1562 ( .A1(DP_OP_422J2_124_3477_n2518), 
        .A2(DP_OP_424J2_126_3477_n2349), .Y(DP_OP_424J2_126_3477_n2335) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1648 ( .A1(DP_OP_422J2_124_3477_n2560), 
        .A2(DP_OP_425J2_127_3477_n2434), .Y(DP_OP_425J2_127_3477_n2418) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1950 ( .A1(DP_OP_423J2_125_3477_n2729), 
        .A2(DP_OP_423J2_125_3477_n2737), .Y(DP_OP_423J2_125_3477_n2721) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1643 ( .A1(DP_OP_423J2_125_3477_n2425), 
        .A2(DP_OP_423J2_125_3477_n2432), .Y(DP_OP_423J2_125_3477_n2417) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1872 ( .A1(DP_OP_424J2_126_3477_n2650), 
        .A2(DP_OP_424J2_126_3477_n2654), .Y(DP_OP_424J2_126_3477_n2642) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1342 ( .A1(DP_OP_423J2_125_3477_n2030), 
        .A2(DP_OP_424J2_126_3477_n2129), .Y(DP_OP_424J2_126_3477_n2115) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1643 ( .A1(DP_OP_425J2_127_3477_n2429), 
        .A2(DP_OP_425J2_127_3477_n2433), .Y(DP_OP_425J2_127_3477_n2413) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1768 ( .A1(DP_OP_425J2_127_3477_n2213), 
        .A2(DP_OP_425J2_127_3477_n2564), .Y(DP_OP_424J2_126_3477_n2538) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1422 ( .A1(DP_OP_423J2_125_3477_n2204), 
        .A2(DP_OP_423J2_125_3477_n2212), .Y(DP_OP_423J2_125_3477_n2196) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2120 ( .A1(DP_OP_425J2_127_3477_n1861), 
        .A2(DP_OP_422J2_124_3477_n2916), .Y(DP_OP_424J2_126_3477_n2890) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2066 ( .A1(DP_OP_423J2_125_3477_n2861), 
        .A2(DP_OP_423J2_125_3477_n2867), .Y(DP_OP_423J2_125_3477_n2837) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1650 ( .A1(DP_OP_425J2_127_3477_n2428), 
        .A2(DP_OP_425J2_127_3477_n2434), .Y(DP_OP_425J2_127_3477_n2420) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1185 ( .A1(DP_OP_423J2_125_3477_n1983), 
        .A2(DP_OP_422J2_124_3477_n1995), .Y(DP_OP_423J2_125_3477_n1959) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1635 ( .A1(DP_OP_423J2_125_3477_n2425), 
        .A2(DP_OP_423J2_125_3477_n2431), .Y(DP_OP_423J2_125_3477_n2409) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2112 ( .A1(DP_OP_423J2_125_3477_n2907), 
        .A2(DP_OP_423J2_125_3477_n2911), .Y(DP_OP_423J2_125_3477_n2883) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1758 ( .A1(DP_OP_422J2_124_3477_n2164), 
        .A2(DP_OP_423J2_125_3477_n2562), .Y(DP_OP_423J2_125_3477_n2532) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1650 ( .A1(DP_OP_424J2_126_3477_n2428), 
        .A2(DP_OP_423J2_125_3477_n2432), .Y(DP_OP_424J2_126_3477_n2420) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1652 ( .A1(DP_OP_424J2_126_3477_n2430), 
        .A2(DP_OP_422J2_124_3477_n2436), .Y(DP_OP_424J2_126_3477_n2422) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1004 ( .A1(n370), .A2(
        DP_OP_424J2_126_3477_n2), .Y(DP_OP_424J2_126_3477_n1777) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1078 ( .A1(DP_OP_425J2_127_3477_n2868), 
        .A2(DP_OP_424J2_126_3477_n1865), .Y(DP_OP_424J2_126_3477_n1851) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1188 ( .A1(DP_OP_423J2_125_3477_n1986), 
        .A2(DP_OP_424J2_126_3477_n1995), .Y(DP_OP_423J2_125_3477_n1962) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1432 ( .A1(DP_OP_425J2_127_3477_n2213), 
        .A2(DP_OP_425J2_127_3477_n2217), .Y(DP_OP_425J2_127_3477_n2205) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1958 ( .A1(DP_OP_424J2_126_3477_n2736), 
        .A2(DP_OP_424J2_126_3477_n2742), .Y(DP_OP_424J2_126_3477_n2728) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1826 ( .A1(DP_OP_424J2_126_3477_n2604), 
        .A2(DP_OP_424J2_126_3477_n2610), .Y(DP_OP_424J2_126_3477_n2596) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1005 ( .A1(n393), .A2(
        DP_OP_425J2_127_3477_n2), .Y(DP_OP_424J2_126_3477_n1778) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2065 ( .A1(DP_OP_423J2_125_3477_n2860), 
        .A2(DP_OP_423J2_125_3477_n2867), .Y(DP_OP_423J2_125_3477_n2836) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2120 ( .A1(DP_OP_425J2_127_3477_n2914), 
        .A2(DP_OP_425J2_127_3477_n2916), .Y(DP_OP_425J2_127_3477_n2890) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1760 ( .A1(DP_OP_423J2_125_3477_n2558), 
        .A2(DP_OP_423J2_125_3477_n2562), .Y(DP_OP_423J2_125_3477_n2534) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1642 ( .A1(DP_OP_423J2_125_3477_n2424), 
        .A2(DP_OP_423J2_125_3477_n2432), .Y(DP_OP_423J2_125_3477_n2416) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1564 ( .A1(DP_OP_425J2_127_3477_n2386), 
        .A2(DP_OP_424J2_126_3477_n2349), .Y(DP_OP_424J2_126_3477_n2337) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1958 ( .A1(DP_OP_423J2_125_3477_n1898), 
        .A2(DP_OP_424J2_126_3477_n2742), .Y(DP_OP_425J2_127_3477_n2728) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1757 ( .A1(DP_OP_425J2_127_3477_n2296), 
        .A2(DP_OP_423J2_125_3477_n2562), .Y(DP_OP_423J2_125_3477_n2531) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1870 ( .A1(DP_OP_422J2_124_3477_n2780), 
        .A2(DP_OP_425J2_127_3477_n2654), .Y(DP_OP_425J2_127_3477_n2640) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2076 ( .A1(DP_OP_425J2_127_3477_n2870), 
        .A2(DP_OP_425J2_127_3477_n2872), .Y(DP_OP_425J2_127_3477_n2846) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1375 ( .A1(DP_OP_425J2_127_3477_n2164), 
        .A2(DP_OP_425J2_127_3477_n2172), .Y(DP_OP_425J2_127_3477_n2148) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2076 ( .A1(DP_OP_425J2_127_3477_n1905), 
        .A2(DP_OP_425J2_127_3477_n2872), .Y(DP_OP_424J2_126_3477_n2846) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1562 ( .A1(DP_OP_424J2_126_3477_n2428), 
        .A2(DP_OP_425J2_127_3477_n2349), .Y(DP_OP_425J2_127_3477_n2335) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1371 ( .A1(DP_OP_423J2_125_3477_n2161), 
        .A2(DP_OP_423J2_125_3477_n2167), .Y(DP_OP_423J2_125_3477_n2145) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1639 ( .A1(DP_OP_424J2_126_3477_n2296), 
        .A2(DP_OP_425J2_127_3477_n2433), .Y(DP_OP_425J2_127_3477_n2409) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1768 ( .A1(DP_OP_423J2_125_3477_n2076), 
        .A2(DP_OP_425J2_127_3477_n2564), .Y(DP_OP_425J2_127_3477_n2538) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1004 ( .A1(n368), .A2(
        DP_OP_425J2_127_3477_n2), .Y(DP_OP_422J2_124_3477_n1777) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1686 ( .A1(DP_OP_423J2_125_3477_n2468), 
        .A2(DP_OP_423J2_125_3477_n2476), .Y(DP_OP_423J2_125_3477_n2460) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1764 ( .A1(DP_OP_425J2_127_3477_n2558), 
        .A2(DP_OP_425J2_127_3477_n2564), .Y(DP_OP_425J2_127_3477_n2534) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1078 ( .A1(DP_OP_424J2_126_3477_n2912), 
        .A2(DP_OP_422J2_124_3477_n1865), .Y(DP_OP_425J2_127_3477_n1851) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1340 ( .A1(DP_OP_422J2_124_3477_n1989), 
        .A2(DP_OP_425J2_127_3477_n2129), .Y(DP_OP_425J2_127_3477_n2113) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1774 ( .A1(DP_OP_422J2_124_3477_n2164), 
        .A2(DP_OP_425J2_127_3477_n2566), .Y(DP_OP_423J2_125_3477_n2548) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1196 ( .A1(DP_OP_422J2_124_3477_n1861), 
        .A2(DP_OP_425J2_127_3477_n1995), .Y(DP_OP_425J2_127_3477_n1969) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1694 ( .A1(DP_OP_425J2_127_3477_n2472), 
        .A2(DP_OP_424J2_126_3477_n2478), .Y(DP_OP_425J2_127_3477_n2464) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2068 ( .A1(DP_OP_425J2_127_3477_n1991), 
        .A2(DP_OP_423J2_125_3477_n2867), .Y(DP_OP_423J2_125_3477_n2839) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1868 ( .A1(DP_OP_425J2_127_3477_n2646), 
        .A2(DP_OP_425J2_127_3477_n2654), .Y(DP_OP_425J2_127_3477_n2638) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1006 ( .A1(n266), .A2(n337), .Y(
        DP_OP_423J2_125_3477_n1780) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2116 ( .A1(DP_OP_425J2_127_3477_n2910), 
        .A2(DP_OP_425J2_127_3477_n2916), .Y(DP_OP_425J2_127_3477_n2886) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1194 ( .A1(DP_OP_425J2_127_3477_n1991), 
        .A2(DP_OP_425J2_127_3477_n1995), .Y(DP_OP_425J2_127_3477_n1967) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1692 ( .A1(DP_OP_423J2_125_3477_n2160), 
        .A2(DP_OP_424J2_126_3477_n2478), .Y(DP_OP_425J2_127_3477_n2462) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1959 ( .A1(DP_OP_423J2_125_3477_n2031), 
        .A2(DP_OP_422J2_124_3477_n2742), .Y(DP_OP_422J2_124_3477_n2729) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1960 ( .A1(DP_OP_425J2_127_3477_n2738), 
        .A2(DP_OP_423J2_125_3477_n2737), .Y(DP_OP_425J2_127_3477_n2730) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1005 ( .A1(n390), .A2(n337), .Y(
        DP_OP_422J2_124_3477_n1778) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1782 ( .A1(DP_OP_423J2_125_3477_n2646), 
        .A2(DP_OP_424J2_126_3477_n2566), .Y(DP_OP_424J2_126_3477_n2552) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1377 ( .A1(DP_OP_425J2_127_3477_n2166), 
        .A2(DP_OP_425J2_127_3477_n2172), .Y(DP_OP_425J2_127_3477_n2150) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1344 ( .A1(DP_OP_423J2_125_3477_n2733), 
        .A2(DP_OP_425J2_127_3477_n2129), .Y(DP_OP_425J2_127_3477_n2117) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1430 ( .A1(DP_OP_424J2_126_3477_n2211), 
        .A2(DP_OP_422J2_124_3477_n2216), .Y(DP_OP_424J2_126_3477_n2203) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1009 ( .A1(n275), .A2(
        DP_OP_425J2_127_3477_n2), .Y(DP_OP_425J2_127_3477_n1782) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1643 ( .A1(DP_OP_422J2_124_3477_n2211), 
        .A2(DP_OP_422J2_124_3477_n2435), .Y(DP_OP_424J2_126_3477_n2413) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1334 ( .A1(DP_OP_423J2_125_3477_n2116), 
        .A2(DP_OP_424J2_126_3477_n2129), .Y(DP_OP_423J2_125_3477_n2108) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1766 ( .A1(DP_OP_423J2_125_3477_n2074), 
        .A2(DP_OP_425J2_127_3477_n2564), .Y(DP_OP_425J2_127_3477_n2536) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1823 ( .A1(DP_OP_422J2_124_3477_n2603), 
        .A2(DP_OP_422J2_124_3477_n2612), .Y(DP_OP_422J2_124_3477_n2595) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1079 ( .A1(DP_OP_425J2_127_3477_n1992), 
        .A2(DP_OP_422J2_124_3477_n1865), .Y(DP_OP_422J2_124_3477_n1852) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1076 ( .A1(DP_OP_424J2_126_3477_n2910), 
        .A2(DP_OP_424J2_126_3477_n1865), .Y(DP_OP_425J2_127_3477_n1849) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1192 ( .A1(DP_OP_425J2_127_3477_n1989), 
        .A2(DP_OP_425J2_127_3477_n1995), .Y(DP_OP_425J2_127_3477_n1965) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1010 ( .A1(n366), .A2(n338), .Y(
        DP_OP_422J2_124_3477_n1783) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1070 ( .A1(DP_OP_423J2_125_3477_n1852), 
        .A2(DP_OP_423J2_125_3477_n1860), .Y(DP_OP_423J2_125_3477_n1844) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1828 ( .A1(DP_OP_423J2_125_3477_n2032), 
        .A2(DP_OP_425J2_127_3477_n2610), .Y(DP_OP_425J2_127_3477_n2598) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2119 ( .A1(DP_OP_422J2_124_3477_n2913), 
        .A2(DP_OP_422J2_124_3477_n2916), .Y(DP_OP_422J2_124_3477_n2889) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1430 ( .A1(DP_OP_422J2_124_3477_n2078), 
        .A2(DP_OP_425J2_127_3477_n2217), .Y(DP_OP_425J2_127_3477_n2203) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1827 ( .A1(DP_OP_424J2_126_3477_n2124), 
        .A2(DP_OP_425J2_127_3477_n2610), .Y(DP_OP_425J2_127_3477_n2597) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1828 ( .A1(DP_OP_422J2_124_3477_n2036), 
        .A2(DP_OP_424J2_126_3477_n2610), .Y(DP_OP_424J2_126_3477_n2598) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1644 ( .A1(DP_OP_425J2_127_3477_n2430), 
        .A2(DP_OP_425J2_127_3477_n2433), .Y(DP_OP_425J2_127_3477_n2414) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U985 ( .A1(n414), .A2(
        DP_OP_425J2_127_3477_n2), .Y(DP_OP_424J2_126_3477_n153) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1871 ( .A1(DP_OP_424J2_126_3477_n2649), 
        .A2(DP_OP_424J2_126_3477_n2654), .Y(DP_OP_424J2_126_3477_n2641) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1695 ( .A1(DP_OP_423J2_125_3477_n2295), 
        .A2(DP_OP_422J2_124_3477_n2480), .Y(DP_OP_422J2_124_3477_n2467) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1695 ( .A1(DP_OP_423J2_125_3477_n2163), 
        .A2(DP_OP_423J2_125_3477_n2476), .Y(DP_OP_425J2_127_3477_n2465) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1000 ( .A1(n292), .A2(
        DP_OP_423J2_125_3477_n2), .Y(DP_OP_423J2_125_3477_n1774) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1825 ( .A1(DP_OP_422J2_124_3477_n2605), 
        .A2(DP_OP_422J2_124_3477_n2612), .Y(DP_OP_422J2_124_3477_n2597) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1378 ( .A1(DP_OP_423J2_125_3477_n2558), 
        .A2(DP_OP_422J2_124_3477_n2171), .Y(DP_OP_422J2_124_3477_n2150) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1644 ( .A1(DP_OP_424J2_126_3477_n2430), 
        .A2(DP_OP_423J2_125_3477_n2431), .Y(DP_OP_424J2_126_3477_n2414) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1783 ( .A1(DP_OP_424J2_126_3477_n2561), 
        .A2(DP_OP_424J2_126_3477_n2566), .Y(DP_OP_424J2_126_3477_n2553) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1695 ( .A1(DP_OP_425J2_127_3477_n2300), 
        .A2(DP_OP_424J2_126_3477_n2478), .Y(DP_OP_424J2_126_3477_n2465) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1192 ( .A1(DP_OP_422J2_124_3477_n1989), 
        .A2(DP_OP_422J2_124_3477_n1995), .Y(DP_OP_422J2_124_3477_n1965) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1696 ( .A1(DP_OP_423J2_125_3477_n2164), 
        .A2(DP_OP_422J2_124_3477_n2480), .Y(DP_OP_425J2_127_3477_n2466) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1956 ( .A1(DP_OP_425J2_127_3477_n2734), 
        .A2(DP_OP_423J2_125_3477_n2737), .Y(DP_OP_425J2_127_3477_n2726) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1007 ( .A1(n271), .A2(n337), .Y(
        DP_OP_423J2_125_3477_n1781) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1651 ( .A1(DP_OP_423J2_125_3477_n2339), 
        .A2(DP_OP_422J2_124_3477_n2436), .Y(DP_OP_422J2_124_3477_n2423) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1563 ( .A1(DP_OP_423J2_125_3477_n2515), 
        .A2(DP_OP_425J2_127_3477_n2349), .Y(DP_OP_425J2_127_3477_n2336) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1373 ( .A1(DP_OP_423J2_125_3477_n2163), 
        .A2(DP_OP_423J2_125_3477_n2167), .Y(DP_OP_423J2_125_3477_n2147) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1764 ( .A1(DP_OP_425J2_127_3477_n2209), 
        .A2(DP_OP_422J2_124_3477_n2566), .Y(DP_OP_424J2_126_3477_n2534) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1824 ( .A1(DP_OP_423J2_125_3477_n2028), 
        .A2(DP_OP_425J2_127_3477_n2610), .Y(DP_OP_425J2_127_3477_n2594) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1956 ( .A1(DP_OP_422J2_124_3477_n2734), 
        .A2(DP_OP_422J2_124_3477_n2742), .Y(DP_OP_422J2_124_3477_n2726) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1651 ( .A1(DP_OP_423J2_125_3477_n2515), 
        .A2(DP_OP_422J2_124_3477_n2436), .Y(DP_OP_424J2_126_3477_n2421) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1781 ( .A1(DP_OP_425J2_127_3477_n2427), 
        .A2(DP_OP_422J2_124_3477_n2568), .Y(DP_OP_422J2_124_3477_n2553) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1824 ( .A1(DP_OP_422J2_124_3477_n2604), 
        .A2(DP_OP_422J2_124_3477_n2612), .Y(DP_OP_422J2_124_3477_n2596) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1380 ( .A1(DP_OP_422J2_124_3477_n2696), 
        .A2(DP_OP_425J2_127_3477_n2172), .Y(DP_OP_424J2_126_3477_n2153) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1957 ( .A1(DP_OP_422J2_124_3477_n2735), 
        .A2(DP_OP_422J2_124_3477_n2742), .Y(DP_OP_422J2_124_3477_n2727) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1563 ( .A1(DP_OP_424J2_126_3477_n2344), 
        .A2(DP_OP_424J2_126_3477_n2349), .Y(DP_OP_424J2_126_3477_n2336) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1768 ( .A1(DP_OP_422J2_124_3477_n2564), 
        .A2(DP_OP_422J2_124_3477_n2566), .Y(DP_OP_422J2_124_3477_n2540) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1564 ( .A1(DP_OP_423J2_125_3477_n2516), 
        .A2(DP_OP_425J2_127_3477_n2349), .Y(DP_OP_425J2_127_3477_n2337) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1783 ( .A1(DP_OP_424J2_126_3477_n2168), 
        .A2(DP_OP_425J2_127_3477_n2566), .Y(DP_OP_425J2_127_3477_n2553) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1782 ( .A1(DP_OP_422J2_124_3477_n2562), 
        .A2(DP_OP_422J2_124_3477_n2568), .Y(DP_OP_422J2_124_3477_n2554) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1869 ( .A1(DP_OP_422J2_124_3477_n2649), 
        .A2(DP_OP_422J2_124_3477_n2656), .Y(DP_OP_422J2_124_3477_n2641) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1343 ( .A1(DP_OP_424J2_126_3477_n2124), 
        .A2(DP_OP_424J2_126_3477_n2129), .Y(DP_OP_424J2_126_3477_n2116) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1380 ( .A1(DP_OP_425J2_127_3477_n2169), 
        .A2(DP_OP_425J2_127_3477_n2172), .Y(DP_OP_425J2_127_3477_n2153) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1014 ( .A1(n286), .A2(n337), .Y(
        DP_OP_424J2_126_3477_n1787) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1826 ( .A1(DP_OP_423J2_125_3477_n2030), 
        .A2(DP_OP_425J2_127_3477_n2610), .Y(DP_OP_425J2_127_3477_n2596) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1652 ( .A1(DP_OP_425J2_127_3477_n2430), 
        .A2(DP_OP_425J2_127_3477_n2434), .Y(DP_OP_425J2_127_3477_n2422) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1077 ( .A1(DP_OP_422J2_124_3477_n1858), 
        .A2(DP_OP_422J2_124_3477_n1865), .Y(DP_OP_422J2_124_3477_n1850) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1827 ( .A1(DP_OP_422J2_124_3477_n2607), 
        .A2(DP_OP_422J2_124_3477_n2612), .Y(DP_OP_422J2_124_3477_n2599) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1696 ( .A1(DP_OP_424J2_126_3477_n2474), 
        .A2(DP_OP_424J2_126_3477_n2478), .Y(DP_OP_424J2_126_3477_n2466) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1959 ( .A1(DP_OP_422J2_124_3477_n2869), 
        .A2(DP_OP_423J2_125_3477_n2737), .Y(DP_OP_425J2_127_3477_n2729) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1343 ( .A1(DP_OP_423J2_125_3477_n2732), 
        .A2(DP_OP_425J2_127_3477_n2129), .Y(DP_OP_425J2_127_3477_n2116) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1344 ( .A1(DP_OP_424J2_126_3477_n2125), 
        .A2(DP_OP_424J2_126_3477_n2129), .Y(DP_OP_424J2_126_3477_n2117) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1871 ( .A1(DP_OP_422J2_124_3477_n2651), 
        .A2(DP_OP_422J2_124_3477_n2656), .Y(DP_OP_422J2_124_3477_n2643) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1871 ( .A1(DP_OP_425J2_127_3477_n2649), 
        .A2(DP_OP_425J2_127_3477_n2654), .Y(DP_OP_425J2_127_3477_n2641) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1827 ( .A1(DP_OP_422J2_124_3477_n2035), 
        .A2(DP_OP_424J2_126_3477_n2610), .Y(DP_OP_424J2_126_3477_n2597) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1014 ( .A1(n385), .A2(n338), .Y(
        DP_OP_425J2_127_3477_n1787) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1642 ( .A1(DP_OP_422J2_124_3477_n2430), 
        .A2(DP_OP_422J2_124_3477_n2435), .Y(DP_OP_422J2_124_3477_n2414) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1432 ( .A1(DP_OP_425J2_127_3477_n2518), 
        .A2(DP_OP_425J2_127_3477_n2217), .Y(DP_OP_424J2_126_3477_n2205) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1649 ( .A1(DP_OP_422J2_124_3477_n2429), 
        .A2(DP_OP_422J2_124_3477_n2436), .Y(DP_OP_422J2_124_3477_n2421) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1343 ( .A1(DP_OP_424J2_126_3477_n2517), 
        .A2(DP_OP_422J2_124_3477_n2128), .Y(DP_OP_422J2_124_3477_n2115) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1194 ( .A1(DP_OP_422J2_124_3477_n1991), 
        .A2(DP_OP_422J2_124_3477_n1995), .Y(DP_OP_422J2_124_3477_n1967) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1428 ( .A1(DP_OP_425J2_127_3477_n2209), 
        .A2(DP_OP_425J2_127_3477_n2217), .Y(DP_OP_425J2_127_3477_n2201) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2118 ( .A1(DP_OP_425J2_127_3477_n2912), 
        .A2(DP_OP_425J2_127_3477_n2916), .Y(DP_OP_425J2_127_3477_n2888) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1782 ( .A1(DP_OP_422J2_124_3477_n2694), 
        .A2(DP_OP_425J2_127_3477_n2566), .Y(DP_OP_425J2_127_3477_n2552) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1380 ( .A1(DP_OP_422J2_124_3477_n2168), 
        .A2(DP_OP_422J2_124_3477_n2171), .Y(DP_OP_422J2_124_3477_n2152) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1006 ( .A1(n402), .A2(
        DP_OP_424J2_126_3477_n2), .Y(DP_OP_424J2_126_3477_n1779) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1784 ( .A1(DP_OP_425J2_127_3477_n2213), 
        .A2(DP_OP_424J2_126_3477_n2566), .Y(DP_OP_424J2_126_3477_n2554) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1872 ( .A1(DP_OP_425J2_127_3477_n2650), 
        .A2(DP_OP_425J2_127_3477_n2654), .Y(DP_OP_425J2_127_3477_n2642) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1080 ( .A1(DP_OP_425J2_127_3477_n2870), 
        .A2(DP_OP_424J2_126_3477_n1865), .Y(DP_OP_424J2_126_3477_n1853) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U986 ( .A1(n424), .A2(n337), .Y(
        DP_OP_424J2_126_3477_n155) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1431 ( .A1(DP_OP_424J2_126_3477_n2212), 
        .A2(DP_OP_423J2_125_3477_n2212), .Y(DP_OP_424J2_126_3477_n2204) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1651 ( .A1(DP_OP_425J2_127_3477_n2429), 
        .A2(DP_OP_425J2_127_3477_n2434), .Y(DP_OP_425J2_127_3477_n2421) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2110 ( .A1(DP_OP_425J2_127_3477_n1945), 
        .A2(DP_OP_423J2_125_3477_n2911), .Y(DP_OP_423J2_125_3477_n2881) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1431 ( .A1(DP_OP_422J2_124_3477_n2211), 
        .A2(DP_OP_422J2_124_3477_n2216), .Y(DP_OP_422J2_124_3477_n2203) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U987 ( .A1(n407), .A2(
        DP_OP_424J2_126_3477_n2), .Y(DP_OP_424J2_126_3477_n157) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2072 ( .A1(DP_OP_423J2_125_3477_n1896), 
        .A2(DP_OP_422J2_124_3477_n2872), .Y(DP_OP_422J2_124_3477_n2842) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1563 ( .A1(DP_OP_422J2_124_3477_n2343), 
        .A2(DP_OP_423J2_125_3477_n2344), .Y(DP_OP_422J2_124_3477_n2335) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1431 ( .A1(DP_OP_423J2_125_3477_n2647), 
        .A2(DP_OP_425J2_127_3477_n2217), .Y(DP_OP_425J2_127_3477_n2204) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1862 ( .A1(DP_OP_425J2_127_3477_n2209), 
        .A2(DP_OP_424J2_126_3477_n2654), .Y(DP_OP_423J2_125_3477_n2636) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1075 ( .A1(DP_OP_424J2_126_3477_n2777), 
        .A2(DP_OP_422J2_124_3477_n1865), .Y(DP_OP_422J2_124_3477_n1848) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1561 ( .A1(DP_OP_422J2_124_3477_n2341), 
        .A2(DP_OP_425J2_127_3477_n2349), .Y(DP_OP_422J2_124_3477_n2333) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1080 ( .A1(DP_OP_425J2_127_3477_n1861), 
        .A2(DP_OP_422J2_124_3477_n1865), .Y(DP_OP_425J2_127_3477_n1853) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1641 ( .A1(DP_OP_425J2_127_3477_n2427), 
        .A2(DP_OP_425J2_127_3477_n2433), .Y(DP_OP_425J2_127_3477_n2411) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1369 ( .A1(DP_OP_425J2_127_3477_n2469), 
        .A2(DP_OP_423J2_125_3477_n2167), .Y(DP_OP_423J2_125_3477_n2143) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U988 ( .A1(n378), .A2(
        DP_OP_423J2_125_3477_n2), .Y(DP_OP_424J2_126_3477_n159) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1693 ( .A1(DP_OP_422J2_124_3477_n2473), 
        .A2(DP_OP_422J2_124_3477_n2480), .Y(DP_OP_422J2_124_3477_n2465) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2117 ( .A1(DP_OP_423J2_125_3477_n2904), 
        .A2(DP_OP_424J2_126_3477_n2917), .Y(DP_OP_423J2_125_3477_n2888) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1232 ( .A1(DP_OP_423J2_125_3477_n2030), 
        .A2(DP_OP_423J2_125_3477_n2034), .Y(DP_OP_423J2_125_3477_n2006) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2126 ( .A1(DP_OP_422J2_124_3477_n2912), 
        .A2(DP_OP_422J2_124_3477_n2917), .Y(DP_OP_422J2_124_3477_n2896) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1070 ( .A1(DP_OP_424J2_126_3477_n2912), 
        .A2(DP_OP_425J2_127_3477_n1864), .Y(DP_OP_425J2_127_3477_n1843) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1591 ( .A1(DP_OP_422J2_124_3477_n2341), 
        .A2(DP_OP_423J2_125_3477_n2387), .Y(DP_OP_423J2_125_3477_n2365) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1502 ( .A1(DP_OP_423J2_125_3477_n2558), 
        .A2(DP_OP_423J2_125_3477_n2298), .Y(DP_OP_425J2_127_3477_n2275) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1599 ( .A1(DP_OP_422J2_124_3477_n2387), 
        .A2(DP_OP_422J2_124_3477_n2391), .Y(DP_OP_422J2_124_3477_n2371) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1165 ( .A1(DP_OP_425J2_127_3477_n2078), 
        .A2(DP_OP_425J2_127_3477_n1953), .Y(DP_OP_422J2_124_3477_n1938) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1815 ( .A1(DP_OP_424J2_126_3477_n2120), 
        .A2(DP_OP_423J2_125_3477_n2607), .Y(DP_OP_425J2_127_3477_n2585) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1166 ( .A1(DP_OP_423J2_125_3477_n2907), 
        .A2(DP_OP_425J2_127_3477_n1953), .Y(DP_OP_425J2_127_3477_n1939) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1724 ( .A1(DP_OP_425J2_127_3477_n2518), 
        .A2(DP_OP_424J2_126_3477_n2520), .Y(DP_OP_425J2_127_3477_n2494) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2037 ( .A1(DP_OP_425J2_127_3477_n2823), 
        .A2(DP_OP_425J2_127_3477_n2829), .Y(DP_OP_425J2_127_3477_n2807) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1422 ( .A1(DP_OP_422J2_124_3477_n2210), 
        .A2(DP_OP_422J2_124_3477_n2215), .Y(DP_OP_422J2_124_3477_n2194) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1802 ( .A1(DP_OP_423J2_125_3477_n2600), 
        .A2(n451), .Y(DP_OP_423J2_125_3477_n2576) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1072 ( .A1(DP_OP_422J2_124_3477_n1861), 
        .A2(DP_OP_422J2_124_3477_n1864), .Y(DP_OP_422J2_124_3477_n1845) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1415 ( .A1(DP_OP_423J2_125_3477_n2205), 
        .A2(DP_OP_423J2_125_3477_n2211), .Y(DP_OP_423J2_125_3477_n2189) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1423 ( .A1(DP_OP_423J2_125_3477_n2647), 
        .A2(DP_OP_422J2_124_3477_n2215), .Y(DP_OP_425J2_127_3477_n2196) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1511 ( .A1(DP_OP_422J2_124_3477_n2299), 
        .A2(DP_OP_423J2_125_3477_n2299), .Y(DP_OP_422J2_124_3477_n2283) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1466 ( .A1(DP_OP_424J2_126_3477_n2384), 
        .A2(DP_OP_422J2_124_3477_n2259), .Y(DP_OP_422J2_124_3477_n2238) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1386 ( .A1(DP_OP_424J2_126_3477_n2472), 
        .A2(DP_OP_425J2_127_3477_n2173), .Y(DP_OP_422J2_124_3477_n2158) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1809 ( .A1(DP_OP_423J2_125_3477_n2599), 
        .A2(DP_OP_423J2_125_3477_n2607), .Y(DP_OP_423J2_125_3477_n2583) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1554 ( .A1(DP_OP_424J2_126_3477_n2428), 
        .A2(DP_OP_425J2_127_3477_n2348), .Y(DP_OP_425J2_127_3477_n2327) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1808 ( .A1(DP_OP_423J2_125_3477_n2028), 
        .A2(n451), .Y(DP_OP_425J2_127_3477_n2578) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1626 ( .A1(DP_OP_423J2_125_3477_n2424), 
        .A2(DP_OP_423J2_125_3477_n2430), .Y(DP_OP_423J2_125_3477_n2400) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1635 ( .A1(DP_OP_423J2_125_3477_n2339), 
        .A2(DP_OP_422J2_124_3477_n2434), .Y(DP_OP_422J2_124_3477_n2407) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2126 ( .A1(DP_OP_425J2_127_3477_n2912), 
        .A2(DP_OP_425J2_127_3477_n2917), .Y(DP_OP_425J2_127_3477_n2896) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1818 ( .A1(DP_OP_423J2_125_3477_n2030), 
        .A2(DP_OP_424J2_126_3477_n2609), .Y(DP_OP_425J2_127_3477_n2588) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1067 ( .A1(DP_OP_424J2_126_3477_n2909), 
        .A2(DP_OP_425J2_127_3477_n1864), .Y(DP_OP_425J2_127_3477_n1840) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1299 ( .A1(DP_OP_423J2_125_3477_n2647), 
        .A2(n441), .Y(DP_OP_422J2_124_3477_n2071) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1231 ( .A1(DP_OP_423J2_125_3477_n2029), 
        .A2(DP_OP_423J2_125_3477_n2034), .Y(DP_OP_423J2_125_3477_n2005) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1105 ( .A1(DP_OP_422J2_124_3477_n2865), 
        .A2(n449), .Y(DP_OP_423J2_125_3477_n1879) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1636 ( .A1(DP_OP_422J2_124_3477_n2432), 
        .A2(DP_OP_422J2_124_3477_n2434), .Y(DP_OP_422J2_124_3477_n2408) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1290 ( .A1(DP_OP_425J2_127_3477_n2079), 
        .A2(DP_OP_425J2_127_3477_n2084), .Y(DP_OP_425J2_127_3477_n2063) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1516 ( .A1(DP_OP_425J2_127_3477_n2297), 
        .A2(DP_OP_425J2_127_3477_n2305), .Y(DP_OP_425J2_127_3477_n2289) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1458 ( .A1(DP_OP_425J2_127_3477_n2382), 
        .A2(DP_OP_422J2_124_3477_n2259), .Y(DP_OP_423J2_125_3477_n2232) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1253 ( .A1(DP_OP_422J2_124_3477_n1902), 
        .A2(DP_OP_425J2_127_3477_n2041), .Y(DP_OP_425J2_127_3477_n2026) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1714 ( .A1(DP_OP_422J2_124_3477_n2208), 
        .A2(n444), .Y(DP_OP_423J2_125_3477_n2488) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1553 ( .A1(DP_OP_425J2_127_3477_n2342), 
        .A2(DP_OP_425J2_127_3477_n2348), .Y(DP_OP_425J2_127_3477_n2326) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1165 ( .A1(DP_OP_423J2_125_3477_n2906), 
        .A2(DP_OP_425J2_127_3477_n1953), .Y(DP_OP_425J2_127_3477_n1938) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1474 ( .A1(DP_OP_424J2_126_3477_n2384), 
        .A2(DP_OP_422J2_124_3477_n2260), .Y(DP_OP_422J2_124_3477_n2246) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1239 ( .A1(DP_OP_422J2_124_3477_n2035), 
        .A2(DP_OP_423J2_125_3477_n2034), .Y(DP_OP_422J2_124_3477_n2011) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1209 ( .A1(DP_OP_425J2_127_3477_n1990), 
        .A2(DP_OP_425J2_127_3477_n1997), .Y(DP_OP_425J2_127_3477_n1982) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1252 ( .A1(DP_OP_425J2_127_3477_n2033), 
        .A2(DP_OP_425J2_127_3477_n2041), .Y(DP_OP_425J2_127_3477_n2025) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1494 ( .A1(DP_OP_422J2_124_3477_n2472), 
        .A2(DP_OP_423J2_125_3477_n2298), .Y(DP_OP_423J2_125_3477_n2268) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1370 ( .A1(DP_OP_423J2_125_3477_n2690), 
        .A2(DP_OP_424J2_126_3477_n2171), .Y(DP_OP_425J2_127_3477_n2143) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1372 ( .A1(DP_OP_422J2_124_3477_n2168), 
        .A2(DP_OP_422J2_124_3477_n2170), .Y(DP_OP_422J2_124_3477_n2144) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1208 ( .A1(DP_OP_425J2_127_3477_n1989), 
        .A2(DP_OP_425J2_127_3477_n1997), .Y(DP_OP_425J2_127_3477_n1981) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1061 ( .A1(DP_OP_425J2_127_3477_n2777), 
        .A2(DP_OP_423J2_125_3477_n1859), .Y(DP_OP_423J2_125_3477_n1835) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1326 ( .A1(DP_OP_423J2_125_3477_n2116), 
        .A2(n440), .Y(DP_OP_423J2_125_3477_n2100) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1247 ( .A1(DP_OP_422J2_124_3477_n2035), 
        .A2(DP_OP_422J2_124_3477_n2039), .Y(DP_OP_422J2_124_3477_n2019) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1363 ( .A1(DP_OP_423J2_125_3477_n2161), 
        .A2(n452), .Y(DP_OP_423J2_125_3477_n2137) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1729 ( .A1(DP_OP_423J2_125_3477_n2117), 
        .A2(DP_OP_424J2_126_3477_n2521), .Y(DP_OP_425J2_127_3477_n2499) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1517 ( .A1(DP_OP_422J2_124_3477_n2165), 
        .A2(DP_OP_425J2_127_3477_n2305), .Y(DP_OP_425J2_127_3477_n2290) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1168 ( .A1(DP_OP_424J2_126_3477_n1949), 
        .A2(DP_OP_424J2_126_3477_n1953), .Y(DP_OP_424J2_126_3477_n1941) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1372 ( .A1(DP_OP_425J2_127_3477_n2169), 
        .A2(DP_OP_424J2_126_3477_n2171), .Y(DP_OP_425J2_127_3477_n2145) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1914 ( .A1(DP_OP_425J2_127_3477_n2692), 
        .A2(DP_OP_424J2_126_3477_n2698), .Y(DP_OP_425J2_127_3477_n2684) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1503 ( .A1(DP_OP_425J2_127_3477_n2300), 
        .A2(DP_OP_422J2_124_3477_n2302), .Y(DP_OP_425J2_127_3477_n2276) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1465 ( .A1(DP_OP_422J2_124_3477_n2121), 
        .A2(DP_OP_425J2_127_3477_n2260), .Y(DP_OP_425J2_127_3477_n2238) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2118 ( .A1(DP_OP_425J2_127_3477_n1945), 
        .A2(DP_OP_422J2_124_3477_n2917), .Y(DP_OP_423J2_125_3477_n2889) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1071 ( .A1(DP_OP_425J2_127_3477_n1860), 
        .A2(DP_OP_425J2_127_3477_n1864), .Y(DP_OP_425J2_127_3477_n1844) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2125 ( .A1(DP_OP_425J2_127_3477_n2911), 
        .A2(DP_OP_425J2_127_3477_n2917), .Y(DP_OP_425J2_127_3477_n2895) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1423 ( .A1(DP_OP_422J2_124_3477_n2211), 
        .A2(DP_OP_422J2_124_3477_n2215), .Y(DP_OP_422J2_124_3477_n2195) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2127 ( .A1(DP_OP_425J2_127_3477_n2913), 
        .A2(DP_OP_425J2_127_3477_n2917), .Y(DP_OP_425J2_127_3477_n2897) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1913 ( .A1(DP_OP_425J2_127_3477_n2691), 
        .A2(DP_OP_422J2_124_3477_n2700), .Y(DP_OP_425J2_127_3477_n2683) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1590 ( .A1(DP_OP_422J2_124_3477_n2340), 
        .A2(DP_OP_423J2_125_3477_n2387), .Y(DP_OP_423J2_125_3477_n2364) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1476 ( .A1(DP_OP_422J2_124_3477_n2608), 
        .A2(DP_OP_423J2_125_3477_n2256), .Y(DP_OP_424J2_126_3477_n2249) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1861 ( .A1(DP_OP_423J2_125_3477_n1985), 
        .A2(DP_OP_424J2_126_3477_n2653), .Y(DP_OP_425J2_127_3477_n2631) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1812 ( .A1(DP_OP_424J2_126_3477_n2125), 
        .A2(DP_OP_424J2_126_3477_n2608), .Y(DP_OP_425J2_127_3477_n2582) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2127 ( .A1(DP_OP_422J2_124_3477_n2913), 
        .A2(DP_OP_422J2_124_3477_n2917), .Y(DP_OP_422J2_124_3477_n2897) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1721 ( .A1(DP_OP_422J2_124_3477_n2207), 
        .A2(DP_OP_423J2_125_3477_n2519), .Y(DP_OP_423J2_125_3477_n2495) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1457 ( .A1(DP_OP_423J2_125_3477_n2247), 
        .A2(DP_OP_424J2_126_3477_n2260), .Y(DP_OP_423J2_125_3477_n2231) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1853 ( .A1(DP_OP_423J2_125_3477_n2643), 
        .A2(DP_OP_423J2_125_3477_n2651), .Y(DP_OP_423J2_125_3477_n2627) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1986 ( .A1(DP_OP_425J2_127_3477_n2780), 
        .A2(DP_OP_423J2_125_3477_n2779), .Y(DP_OP_425J2_127_3477_n2756) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1385 ( .A1(DP_OP_422J2_124_3477_n2165), 
        .A2(DP_OP_425J2_127_3477_n2173), .Y(DP_OP_422J2_124_3477_n2157) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1817 ( .A1(DP_OP_423J2_125_3477_n2029), 
        .A2(DP_OP_422J2_124_3477_n2611), .Y(DP_OP_425J2_127_3477_n2587) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1291 ( .A1(DP_OP_423J2_125_3477_n2647), 
        .A2(DP_OP_422J2_124_3477_n2083), .Y(DP_OP_422J2_124_3477_n2063) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1731 ( .A1(DP_OP_424J2_126_3477_n2212), 
        .A2(DP_OP_423J2_125_3477_n2519), .Y(DP_OP_425J2_127_3477_n2501) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1388 ( .A1(DP_OP_423J2_125_3477_n2076), 
        .A2(DP_OP_424J2_126_3477_n2173), .Y(DP_OP_424J2_126_3477_n2161) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1291 ( .A1(DP_OP_424J2_126_3477_n2693), 
        .A2(DP_OP_425J2_127_3477_n2084), .Y(DP_OP_425J2_127_3477_n2064) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2038 ( .A1(DP_OP_424J2_126_3477_n1903), 
        .A2(DP_OP_425J2_127_3477_n2829), .Y(DP_OP_425J2_127_3477_n2808) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1501 ( .A1(DP_OP_423J2_125_3477_n2291), 
        .A2(DP_OP_423J2_125_3477_n2299), .Y(DP_OP_423J2_125_3477_n2275) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1413 ( .A1(DP_OP_424J2_126_3477_n2296), 
        .A2(DP_OP_423J2_125_3477_n2211), .Y(DP_OP_423J2_125_3477_n2187) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1289 ( .A1(DP_OP_425J2_127_3477_n2078), 
        .A2(DP_OP_425J2_127_3477_n2084), .Y(DP_OP_425J2_127_3477_n2062) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2038 ( .A1(DP_OP_424J2_126_3477_n2035), 
        .A2(DP_OP_424J2_126_3477_n2829), .Y(DP_OP_422J2_124_3477_n2808) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1978 ( .A1(DP_OP_422J2_124_3477_n1945), 
        .A2(DP_OP_423J2_125_3477_n2779), .Y(DP_OP_423J2_125_3477_n2749) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1362 ( .A1(DP_OP_423J2_125_3477_n2160), 
        .A2(n452), .Y(DP_OP_423J2_125_3477_n2136) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1495 ( .A1(DP_OP_422J2_124_3477_n2473), 
        .A2(DP_OP_423J2_125_3477_n2298), .Y(DP_OP_423J2_125_3477_n2269) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1598 ( .A1(DP_OP_425J2_127_3477_n2384), 
        .A2(DP_OP_423J2_125_3477_n2387), .Y(DP_OP_425J2_127_3477_n2368) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1164 ( .A1(DP_OP_425J2_127_3477_n1945), 
        .A2(DP_OP_425J2_127_3477_n1953), .Y(DP_OP_425J2_127_3477_n1937) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1545 ( .A1(DP_OP_422J2_124_3477_n2427), 
        .A2(DP_OP_423J2_125_3477_n2343), .Y(DP_OP_423J2_125_3477_n2319) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1238 ( .A1(DP_OP_424J2_126_3477_n2736), 
        .A2(DP_OP_425J2_127_3477_n2039), .Y(DP_OP_425J2_127_3477_n2011) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1862 ( .A1(DP_OP_423J2_125_3477_n1986), 
        .A2(DP_OP_423J2_125_3477_n2651), .Y(DP_OP_425J2_127_3477_n2632) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1325 ( .A1(DP_OP_423J2_125_3477_n2115), 
        .A2(n440), .Y(DP_OP_423J2_125_3477_n2099) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1467 ( .A1(DP_OP_424J2_126_3477_n2385), 
        .A2(DP_OP_422J2_124_3477_n2259), .Y(DP_OP_422J2_124_3477_n2239) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1166 ( .A1(DP_OP_425J2_127_3477_n2079), 
        .A2(DP_OP_423J2_125_3477_n1948), .Y(DP_OP_422J2_124_3477_n1939) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1731 ( .A1(DP_OP_424J2_126_3477_n2344), 
        .A2(DP_OP_422J2_124_3477_n2523), .Y(DP_OP_422J2_124_3477_n2503) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1069 ( .A1(DP_OP_425J2_127_3477_n1858), 
        .A2(DP_OP_425J2_127_3477_n1864), .Y(DP_OP_425J2_127_3477_n1842) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1510 ( .A1(DP_OP_422J2_124_3477_n2298), 
        .A2(DP_OP_425J2_127_3477_n2304), .Y(DP_OP_422J2_124_3477_n2282) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1281 ( .A1(DP_OP_424J2_126_3477_n2164), 
        .A2(DP_OP_422J2_124_3477_n2083), .Y(DP_OP_423J2_125_3477_n2055) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1730 ( .A1(DP_OP_424J2_126_3477_n2211), 
        .A2(DP_OP_424J2_126_3477_n2521), .Y(DP_OP_425J2_127_3477_n2500) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2029 ( .A1(DP_OP_424J2_126_3477_n2733), 
        .A2(DP_OP_423J2_125_3477_n2824), .Y(DP_OP_423J2_125_3477_n2800) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1254 ( .A1(DP_OP_424J2_126_3477_n2736), 
        .A2(DP_OP_425J2_127_3477_n2041), .Y(DP_OP_425J2_127_3477_n2027) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1912 ( .A1(DP_OP_425J2_127_3477_n2690), 
        .A2(DP_OP_424J2_126_3477_n2698), .Y(DP_OP_425J2_127_3477_n2682) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1987 ( .A1(DP_OP_424J2_126_3477_n1948), 
        .A2(DP_OP_424J2_126_3477_n2784), .Y(DP_OP_425J2_127_3477_n2757) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2039 ( .A1(DP_OP_424J2_126_3477_n1904), 
        .A2(DP_OP_425J2_127_3477_n2829), .Y(DP_OP_425J2_127_3477_n2809) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1245 ( .A1(DP_OP_422J2_124_3477_n1902), 
        .A2(DP_OP_425J2_127_3477_n2040), .Y(DP_OP_425J2_127_3477_n2018) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1230 ( .A1(DP_OP_423J2_125_3477_n2028), 
        .A2(DP_OP_423J2_125_3477_n2034), .Y(DP_OP_423J2_125_3477_n2004) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1863 ( .A1(DP_OP_425J2_127_3477_n2649), 
        .A2(DP_OP_423J2_125_3477_n2651), .Y(DP_OP_425J2_127_3477_n2633) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1598 ( .A1(DP_OP_422J2_124_3477_n2386), 
        .A2(DP_OP_422J2_124_3477_n2391), .Y(DP_OP_422J2_124_3477_n2370) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1116 ( .A1(DP_OP_422J2_124_3477_n1905), 
        .A2(DP_OP_422J2_124_3477_n1908), .Y(DP_OP_422J2_124_3477_n1889) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1296 ( .A1(DP_OP_425J2_127_3477_n2077), 
        .A2(DP_OP_423J2_125_3477_n2080), .Y(DP_OP_425J2_127_3477_n2069) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1509 ( .A1(DP_OP_422J2_124_3477_n2165), 
        .A2(DP_OP_425J2_127_3477_n2304), .Y(DP_OP_425J2_127_3477_n2282) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1414 ( .A1(DP_OP_423J2_125_3477_n2204), 
        .A2(DP_OP_423J2_125_3477_n2211), .Y(DP_OP_423J2_125_3477_n2188) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1589 ( .A1(DP_OP_422J2_124_3477_n2339), 
        .A2(DP_OP_423J2_125_3477_n2387), .Y(DP_OP_423J2_125_3477_n2363) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1246 ( .A1(DP_OP_424J2_126_3477_n2604), 
        .A2(DP_OP_422J2_124_3477_n2039), .Y(DP_OP_422J2_124_3477_n2018) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1240 ( .A1(DP_OP_424J2_126_3477_n2738), 
        .A2(DP_OP_425J2_127_3477_n2039), .Y(DP_OP_425J2_127_3477_n2013) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1810 ( .A1(DP_OP_423J2_125_3477_n2030), 
        .A2(DP_OP_424J2_126_3477_n2608), .Y(DP_OP_425J2_127_3477_n2580) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1628 ( .A1(DP_OP_422J2_124_3477_n2298), 
        .A2(DP_OP_423J2_125_3477_n2430), .Y(DP_OP_423J2_125_3477_n2402) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1915 ( .A1(DP_OP_422J2_124_3477_n2695), 
        .A2(DP_OP_422J2_124_3477_n2700), .Y(DP_OP_422J2_124_3477_n2687) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1473 ( .A1(DP_OP_424J2_126_3477_n2383), 
        .A2(DP_OP_422J2_124_3477_n2260), .Y(DP_OP_422J2_124_3477_n2245) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1985 ( .A1(DP_OP_425J2_127_3477_n2779), 
        .A2(DP_OP_424J2_126_3477_n2784), .Y(DP_OP_425J2_127_3477_n2755) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1297 ( .A1(DP_OP_423J2_125_3477_n2645), 
        .A2(n441), .Y(DP_OP_422J2_124_3477_n2069) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2040 ( .A1(DP_OP_424J2_126_3477_n2037), 
        .A2(DP_OP_423J2_125_3477_n2824), .Y(DP_OP_422J2_124_3477_n2810) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1987 ( .A1(DP_OP_422J2_124_3477_n2781), 
        .A2(DP_OP_422J2_124_3477_n2784), .Y(DP_OP_422J2_124_3477_n2757) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1367 ( .A1(DP_OP_425J2_127_3477_n2164), 
        .A2(DP_OP_422J2_124_3477_n2170), .Y(DP_OP_425J2_127_3477_n2140) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1387 ( .A1(DP_OP_423J2_125_3477_n2559), 
        .A2(DP_OP_424J2_126_3477_n2173), .Y(DP_OP_422J2_124_3477_n2159) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1369 ( .A1(DP_OP_425J2_127_3477_n2166), 
        .A2(n452), .Y(DP_OP_425J2_127_3477_n2142) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1818 ( .A1(DP_OP_422J2_124_3477_n2606), 
        .A2(DP_OP_422J2_124_3477_n2611), .Y(DP_OP_422J2_124_3477_n2590) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1728 ( .A1(DP_OP_422J2_124_3477_n2648), 
        .A2(DP_OP_424J2_126_3477_n2521), .Y(DP_OP_425J2_127_3477_n2498) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1512 ( .A1(DP_OP_423J2_125_3477_n2428), 
        .A2(DP_OP_423J2_125_3477_n2299), .Y(DP_OP_422J2_124_3477_n2284) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1070 ( .A1(DP_OP_422J2_124_3477_n1859), 
        .A2(DP_OP_422J2_124_3477_n1864), .Y(DP_OP_422J2_124_3477_n1843) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1862 ( .A1(DP_OP_422J2_124_3477_n2650), 
        .A2(DP_OP_422J2_124_3477_n2655), .Y(DP_OP_422J2_124_3477_n2634) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1600 ( .A1(DP_OP_422J2_124_3477_n2388), 
        .A2(DP_OP_422J2_124_3477_n2391), .Y(DP_OP_422J2_124_3477_n2372) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1807 ( .A1(DP_OP_424J2_126_3477_n2120), 
        .A2(DP_OP_424J2_126_3477_n2608), .Y(DP_OP_425J2_127_3477_n2577) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1422 ( .A1(DP_OP_423J2_125_3477_n2646), 
        .A2(DP_OP_422J2_124_3477_n2215), .Y(DP_OP_425J2_127_3477_n2195) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1115 ( .A1(DP_OP_422J2_124_3477_n1904), 
        .A2(DP_OP_422J2_124_3477_n1908), .Y(DP_OP_422J2_124_3477_n1888) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1723 ( .A1(DP_OP_424J2_126_3477_n2344), 
        .A2(DP_OP_422J2_124_3477_n2522), .Y(DP_OP_422J2_124_3477_n2495) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2128 ( .A1(DP_OP_423J2_125_3477_n1856), 
        .A2(DP_OP_422J2_124_3477_n2917), .Y(DP_OP_422J2_124_3477_n2898) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1475 ( .A1(DP_OP_424J2_126_3477_n2385), 
        .A2(DP_OP_422J2_124_3477_n2260), .Y(DP_OP_422J2_124_3477_n2247) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1114 ( .A1(DP_OP_425J2_127_3477_n1903), 
        .A2(n449), .Y(DP_OP_425J2_127_3477_n1887) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1334 ( .A1(DP_OP_425J2_127_3477_n2255), 
        .A2(DP_OP_422J2_124_3477_n2127), .Y(DP_OP_422J2_124_3477_n2106) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1335 ( .A1(DP_OP_424J2_126_3477_n2517), 
        .A2(DP_OP_422J2_124_3477_n2127), .Y(DP_OP_422J2_124_3477_n2107) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1424 ( .A1(DP_OP_424J2_126_3477_n2430), 
        .A2(DP_OP_422J2_124_3477_n2215), .Y(DP_OP_422J2_124_3477_n2196) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1288 ( .A1(DP_OP_425J2_127_3477_n2077), 
        .A2(DP_OP_425J2_127_3477_n2084), .Y(DP_OP_425J2_127_3477_n2061) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1167 ( .A1(DP_OP_424J2_126_3477_n2693), 
        .A2(DP_OP_425J2_127_3477_n1953), .Y(DP_OP_422J2_124_3477_n1940) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1517 ( .A1(DP_OP_423J2_125_3477_n2425), 
        .A2(DP_OP_422J2_124_3477_n2304), .Y(DP_OP_422J2_124_3477_n2289) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1468 ( .A1(DP_OP_424J2_126_3477_n2386), 
        .A2(DP_OP_422J2_124_3477_n2259), .Y(DP_OP_422J2_124_3477_n2240) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1552 ( .A1(DP_OP_425J2_127_3477_n2341), 
        .A2(DP_OP_425J2_127_3477_n2348), .Y(DP_OP_425J2_127_3477_n2325) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1336 ( .A1(DP_OP_422J2_124_3477_n2124), 
        .A2(DP_OP_422J2_124_3477_n2127), .Y(DP_OP_422J2_124_3477_n2108) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1730 ( .A1(DP_OP_422J2_124_3477_n2518), 
        .A2(DP_OP_422J2_124_3477_n2523), .Y(DP_OP_422J2_124_3477_n2502) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2124 ( .A1(DP_OP_425J2_127_3477_n2910), 
        .A2(DP_OP_425J2_127_3477_n2917), .Y(DP_OP_425J2_127_3477_n2894) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1474 ( .A1(DP_OP_425J2_127_3477_n2255), 
        .A2(DP_OP_425J2_127_3477_n2261), .Y(DP_OP_425J2_127_3477_n2247) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1556 ( .A1(DP_OP_422J2_124_3477_n2344), 
        .A2(DP_OP_422J2_124_3477_n2347), .Y(DP_OP_422J2_124_3477_n2328) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1253 ( .A1(DP_OP_422J2_124_3477_n2033), 
        .A2(DP_OP_422J2_124_3477_n2040), .Y(DP_OP_422J2_124_3477_n2025) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1298 ( .A1(DP_OP_422J2_124_3477_n2078), 
        .A2(n441), .Y(DP_OP_422J2_124_3477_n2070) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1255 ( .A1(DP_OP_422J2_124_3477_n2035), 
        .A2(DP_OP_422J2_124_3477_n2040), .Y(DP_OP_422J2_124_3477_n2027) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1246 ( .A1(DP_OP_422J2_124_3477_n1903), 
        .A2(DP_OP_425J2_127_3477_n2040), .Y(DP_OP_425J2_127_3477_n2019) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1247 ( .A1(DP_OP_424J2_126_3477_n2737), 
        .A2(DP_OP_425J2_127_3477_n2040), .Y(DP_OP_425J2_127_3477_n2020) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1332 ( .A1(DP_OP_423J2_125_3477_n2729), 
        .A2(DP_OP_425J2_127_3477_n2128), .Y(DP_OP_425J2_127_3477_n2105) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1211 ( .A1(DP_OP_423J2_125_3477_n2732), 
        .A2(DP_OP_422J2_124_3477_n1997), .Y(DP_OP_422J2_124_3477_n1984) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1464 ( .A1(DP_OP_422J2_124_3477_n2120), 
        .A2(DP_OP_425J2_127_3477_n2260), .Y(DP_OP_425J2_127_3477_n2237) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1816 ( .A1(DP_OP_423J2_125_3477_n2028), 
        .A2(DP_OP_423J2_125_3477_n2607), .Y(DP_OP_425J2_127_3477_n2586) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1386 ( .A1(DP_OP_423J2_125_3477_n2690), 
        .A2(DP_OP_425J2_127_3477_n2173), .Y(DP_OP_425J2_127_3477_n2159) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1988 ( .A1(DP_OP_422J2_124_3477_n2782), 
        .A2(DP_OP_422J2_124_3477_n2784), .Y(DP_OP_422J2_124_3477_n2758) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1466 ( .A1(DP_OP_425J2_127_3477_n2255), 
        .A2(DP_OP_425J2_127_3477_n2260), .Y(DP_OP_425J2_127_3477_n2239) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1864 ( .A1(DP_OP_422J2_124_3477_n2652), 
        .A2(DP_OP_422J2_124_3477_n2655), .Y(DP_OP_422J2_124_3477_n2636) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1820 ( .A1(DP_OP_422J2_124_3477_n2608), 
        .A2(DP_OP_422J2_124_3477_n2611), .Y(DP_OP_422J2_124_3477_n2592) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1383 ( .A1(DP_OP_425J2_127_3477_n2164), 
        .A2(DP_OP_425J2_127_3477_n2173), .Y(DP_OP_425J2_127_3477_n2156) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1508 ( .A1(DP_OP_425J2_127_3477_n2297), 
        .A2(DP_OP_425J2_127_3477_n2304), .Y(DP_OP_425J2_127_3477_n2281) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1801 ( .A1(DP_OP_423J2_125_3477_n2599), 
        .A2(n451), .Y(DP_OP_423J2_125_3477_n2575) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1636 ( .A1(DP_OP_425J2_127_3477_n2430), 
        .A2(DP_OP_423J2_125_3477_n2430), .Y(DP_OP_425J2_127_3477_n2406) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1334 ( .A1(DP_OP_423J2_125_3477_n2731), 
        .A2(DP_OP_425J2_127_3477_n2128), .Y(DP_OP_425J2_127_3477_n2107) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2030 ( .A1(DP_OP_425J2_127_3477_n2033), 
        .A2(DP_OP_423J2_125_3477_n2824), .Y(DP_OP_423J2_125_3477_n2801) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1229 ( .A1(DP_OP_424J2_126_3477_n2120), 
        .A2(DP_OP_423J2_125_3477_n2034), .Y(DP_OP_423J2_125_3477_n2003) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1071 ( .A1(DP_OP_425J2_127_3477_n1992), 
        .A2(DP_OP_422J2_124_3477_n1864), .Y(DP_OP_422J2_124_3477_n1844) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1501 ( .A1(DP_OP_424J2_126_3477_n2471), 
        .A2(DP_OP_423J2_125_3477_n2298), .Y(DP_OP_425J2_127_3477_n2274) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1113 ( .A1(DP_OP_424J2_126_3477_n2867), 
        .A2(n449), .Y(DP_OP_425J2_127_3477_n1886) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1554 ( .A1(DP_OP_422J2_124_3477_n2342), 
        .A2(DP_OP_422J2_124_3477_n2347), .Y(DP_OP_422J2_124_3477_n2326) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1209 ( .A1(DP_OP_423J2_125_3477_n2730), 
        .A2(DP_OP_422J2_124_3477_n1997), .Y(DP_OP_422J2_124_3477_n1982) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1810 ( .A1(DP_OP_423J2_125_3477_n2600), 
        .A2(DP_OP_423J2_125_3477_n2607), .Y(DP_OP_423J2_125_3477_n2584) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1913 ( .A1(DP_OP_423J2_125_3477_n2073), 
        .A2(DP_OP_422J2_124_3477_n2700), .Y(DP_OP_422J2_124_3477_n2685) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1295 ( .A1(DP_OP_423J2_125_3477_n2772), 
        .A2(n441), .Y(DP_OP_425J2_127_3477_n2068) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1520 ( .A1(DP_OP_423J2_125_3477_n2428), 
        .A2(DP_OP_422J2_124_3477_n2304), .Y(DP_OP_422J2_124_3477_n2292) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1290 ( .A1(DP_OP_422J2_124_3477_n2078), 
        .A2(DP_OP_422J2_124_3477_n2083), .Y(DP_OP_422J2_124_3477_n2062) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1597 ( .A1(DP_OP_425J2_127_3477_n2383), 
        .A2(DP_OP_424J2_126_3477_n2389), .Y(DP_OP_425J2_127_3477_n2367) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1256 ( .A1(DP_OP_422J2_124_3477_n2036), 
        .A2(DP_OP_422J2_124_3477_n2040), .Y(DP_OP_422J2_124_3477_n2028) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1515 ( .A1(DP_OP_425J2_127_3477_n2296), 
        .A2(DP_OP_425J2_127_3477_n2305), .Y(DP_OP_425J2_127_3477_n2288) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1809 ( .A1(DP_OP_423J2_125_3477_n2029), 
        .A2(DP_OP_422J2_124_3477_n2610), .Y(DP_OP_425J2_127_3477_n2579) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1300 ( .A1(DP_OP_425J2_127_3477_n2213), 
        .A2(n441), .Y(DP_OP_422J2_124_3477_n2072) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1916 ( .A1(DP_OP_422J2_124_3477_n2696), 
        .A2(DP_OP_422J2_124_3477_n2700), .Y(DP_OP_422J2_124_3477_n2688) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1979 ( .A1(DP_OP_424J2_126_3477_n2691), 
        .A2(DP_OP_423J2_125_3477_n2779), .Y(DP_OP_423J2_125_3477_n2750) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1333 ( .A1(DP_OP_425J2_127_3477_n2122), 
        .A2(DP_OP_425J2_127_3477_n2128), .Y(DP_OP_425J2_127_3477_n2106) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1062 ( .A1(DP_OP_423J2_125_3477_n1852), 
        .A2(DP_OP_423J2_125_3477_n1859), .Y(DP_OP_423J2_125_3477_n1836) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1631 ( .A1(DP_OP_422J2_124_3477_n2559), 
        .A2(DP_OP_424J2_126_3477_n2432), .Y(DP_OP_425J2_127_3477_n2401) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1212 ( .A1(DP_OP_423J2_125_3477_n2733), 
        .A2(DP_OP_422J2_124_3477_n1997), .Y(DP_OP_422J2_124_3477_n1985) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1472 ( .A1(DP_OP_423J2_125_3477_n2600), 
        .A2(DP_OP_425J2_127_3477_n2261), .Y(DP_OP_425J2_127_3477_n2245) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1384 ( .A1(DP_OP_423J2_125_3477_n2688), 
        .A2(DP_OP_425J2_127_3477_n2173), .Y(DP_OP_425J2_127_3477_n2157) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1983 ( .A1(DP_OP_425J2_127_3477_n2777), 
        .A2(DP_OP_424J2_126_3477_n2784), .Y(DP_OP_425J2_127_3477_n2753) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1722 ( .A1(DP_OP_422J2_124_3477_n2650), 
        .A2(DP_OP_424J2_126_3477_n2520), .Y(DP_OP_425J2_127_3477_n2492) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1722 ( .A1(DP_OP_422J2_124_3477_n2208), 
        .A2(DP_OP_423J2_125_3477_n2519), .Y(DP_OP_423J2_125_3477_n2496) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1282 ( .A1(DP_OP_425J2_127_3477_n2558), 
        .A2(DP_OP_425J2_127_3477_n2084), .Y(DP_OP_423J2_125_3477_n2056) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1421 ( .A1(DP_OP_423J2_125_3477_n2645), 
        .A2(DP_OP_423J2_125_3477_n2211), .Y(DP_OP_425J2_127_3477_n2194) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1518 ( .A1(DP_OP_422J2_124_3477_n2298), 
        .A2(DP_OP_422J2_124_3477_n2304), .Y(DP_OP_422J2_124_3477_n2290) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1546 ( .A1(DP_OP_422J2_124_3477_n2428), 
        .A2(DP_OP_423J2_125_3477_n2343), .Y(DP_OP_423J2_125_3477_n2320) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1819 ( .A1(DP_OP_422J2_124_3477_n2607), 
        .A2(DP_OP_422J2_124_3477_n2611), .Y(DP_OP_422J2_124_3477_n2591) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1248 ( .A1(DP_OP_422J2_124_3477_n2036), 
        .A2(DP_OP_422J2_124_3477_n2039), .Y(DP_OP_422J2_124_3477_n2020) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1863 ( .A1(DP_OP_422J2_124_3477_n2651), 
        .A2(DP_OP_422J2_124_3477_n2655), .Y(DP_OP_422J2_124_3477_n2635) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1634 ( .A1(DP_OP_425J2_127_3477_n2428), 
        .A2(DP_OP_422J2_124_3477_n2434), .Y(DP_OP_425J2_127_3477_n2404) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1235 ( .A1(DP_OP_424J2_126_3477_n2733), 
        .A2(DP_OP_425J2_127_3477_n2039), .Y(DP_OP_425J2_127_3477_n2008) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1719 ( .A1(DP_OP_422J2_124_3477_n2647), 
        .A2(DP_OP_424J2_126_3477_n2520), .Y(DP_OP_425J2_127_3477_n2489) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1499 ( .A1(DP_OP_425J2_127_3477_n2296), 
        .A2(DP_OP_423J2_125_3477_n2298), .Y(DP_OP_425J2_127_3477_n2272) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1503 ( .A1(DP_OP_422J2_124_3477_n2299), 
        .A2(DP_OP_422J2_124_3477_n2302), .Y(DP_OP_422J2_124_3477_n2275) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1854 ( .A1(DP_OP_425J2_127_3477_n2209), 
        .A2(DP_OP_423J2_125_3477_n2651), .Y(DP_OP_423J2_125_3477_n2628) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1812 ( .A1(DP_OP_422J2_124_3477_n2608), 
        .A2(DP_OP_422J2_124_3477_n2610), .Y(DP_OP_422J2_124_3477_n2584) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1977 ( .A1(DP_OP_423J2_125_3477_n2772), 
        .A2(DP_OP_423J2_125_3477_n2779), .Y(DP_OP_423J2_125_3477_n2748) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1633 ( .A1(DP_OP_425J2_127_3477_n2427), 
        .A2(DP_OP_424J2_126_3477_n2432), .Y(DP_OP_425J2_127_3477_n2403) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1915 ( .A1(DP_OP_423J2_125_3477_n1943), 
        .A2(DP_OP_422J2_124_3477_n2700), .Y(DP_OP_425J2_127_3477_n2685) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1112 ( .A1(DP_OP_425J2_127_3477_n1901), 
        .A2(DP_OP_424J2_126_3477_n1908), .Y(DP_OP_425J2_127_3477_n1885) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1240 ( .A1(DP_OP_422J2_124_3477_n2036), 
        .A2(DP_OP_423J2_125_3477_n2034), .Y(DP_OP_422J2_124_3477_n2012) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1596 ( .A1(DP_OP_425J2_127_3477_n2382), 
        .A2(DP_OP_422J2_124_3477_n2391), .Y(DP_OP_425J2_127_3477_n2366) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2039 ( .A1(DP_OP_422J2_124_3477_n2825), 
        .A2(DP_OP_424J2_126_3477_n2829), .Y(DP_OP_422J2_124_3477_n2809) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1724 ( .A1(DP_OP_422J2_124_3477_n2520), 
        .A2(DP_OP_422J2_124_3477_n2522), .Y(DP_OP_422J2_124_3477_n2496) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1555 ( .A1(DP_OP_423J2_125_3477_n2515), 
        .A2(DP_OP_425J2_127_3477_n2348), .Y(DP_OP_425J2_127_3477_n2328) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1371 ( .A1(DP_OP_425J2_127_3477_n2168), 
        .A2(n452), .Y(DP_OP_425J2_127_3477_n2144) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1210 ( .A1(DP_OP_425J2_127_3477_n1991), 
        .A2(DP_OP_425J2_127_3477_n1997), .Y(DP_OP_425J2_127_3477_n1983) );
  XNOR2X1_HVT DP_OP_423J2_125_3477_U621 ( .A1(DP_OP_423J2_125_3477_n2699), 
        .A2(DP_OP_423J2_125_3477_n1997), .Y(DP_OP_423J2_125_3477_n1057) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1500 ( .A1(DP_OP_425J2_127_3477_n2297), 
        .A2(n445), .Y(DP_OP_425J2_127_3477_n2273) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1504 ( .A1(DP_OP_422J2_124_3477_n2168), 
        .A2(n445), .Y(DP_OP_425J2_127_3477_n2277) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1727 ( .A1(DP_OP_423J2_125_3477_n2115), 
        .A2(DP_OP_422J2_124_3477_n2523), .Y(DP_OP_425J2_127_3477_n2497) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1287 ( .A1(DP_OP_424J2_126_3477_n2689), 
        .A2(DP_OP_425J2_127_3477_n2084), .Y(DP_OP_425J2_127_3477_n2060) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2035 ( .A1(DP_OP_425J2_127_3477_n2821), 
        .A2(DP_OP_425J2_127_3477_n2829), .Y(DP_OP_425J2_127_3477_n2805) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1106 ( .A1(DP_OP_423J2_125_3477_n1896), 
        .A2(n449), .Y(DP_OP_423J2_125_3477_n1880) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1368 ( .A1(DP_OP_423J2_125_3477_n2688), 
        .A2(DP_OP_422J2_124_3477_n2170), .Y(DP_OP_425J2_127_3477_n2141) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1984 ( .A1(DP_OP_425J2_127_3477_n2778), 
        .A2(DP_OP_422J2_124_3477_n2784), .Y(DP_OP_425J2_127_3477_n2754) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1502 ( .A1(DP_OP_422J2_124_3477_n2472), 
        .A2(DP_OP_423J2_125_3477_n2299), .Y(DP_OP_423J2_125_3477_n2276) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1297 ( .A1(DP_OP_425J2_127_3477_n2078), 
        .A2(DP_OP_423J2_125_3477_n2080), .Y(DP_OP_425J2_127_3477_n2070) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1419 ( .A1(DP_OP_424J2_126_3477_n2557), 
        .A2(DP_OP_422J2_124_3477_n2215), .Y(DP_OP_425J2_127_3477_n2192) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1988 ( .A1(DP_OP_424J2_126_3477_n1949), 
        .A2(DP_OP_423J2_125_3477_n2779), .Y(DP_OP_425J2_127_3477_n2758) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1720 ( .A1(DP_OP_422J2_124_3477_n2648), 
        .A2(n444), .Y(DP_OP_425J2_127_3477_n2490) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1803 ( .A1(DP_OP_423J2_125_3477_n2601), 
        .A2(n451), .Y(DP_OP_423J2_125_3477_n2577) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1236 ( .A1(DP_OP_425J2_127_3477_n2033), 
        .A2(DP_OP_425J2_127_3477_n2039), .Y(DP_OP_425J2_127_3477_n2009) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1819 ( .A1(DP_OP_424J2_126_3477_n2124), 
        .A2(DP_OP_424J2_126_3477_n2609), .Y(DP_OP_425J2_127_3477_n2589) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2123 ( .A1(DP_OP_425J2_127_3477_n2909), 
        .A2(DP_OP_425J2_127_3477_n2917), .Y(DP_OP_425J2_127_3477_n2893) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1551 ( .A1(DP_OP_425J2_127_3477_n2340), 
        .A2(DP_OP_425J2_127_3477_n2348), .Y(DP_OP_425J2_127_3477_n2324) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1518 ( .A1(DP_OP_424J2_126_3477_n2472), 
        .A2(DP_OP_425J2_127_3477_n2305), .Y(DP_OP_425J2_127_3477_n2291) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1507 ( .A1(DP_OP_425J2_127_3477_n2296), 
        .A2(DP_OP_425J2_127_3477_n2304), .Y(DP_OP_425J2_127_3477_n2280) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1068 ( .A1(DP_OP_424J2_126_3477_n2910), 
        .A2(DP_OP_425J2_127_3477_n1864), .Y(DP_OP_425J2_127_3477_n1841) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1371 ( .A1(DP_OP_425J2_127_3477_n2300), 
        .A2(DP_OP_422J2_124_3477_n2170), .Y(DP_OP_422J2_124_3477_n2143) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1732 ( .A1(DP_OP_422J2_124_3477_n2520), 
        .A2(DP_OP_422J2_124_3477_n2523), .Y(DP_OP_422J2_124_3477_n2504) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1292 ( .A1(DP_OP_425J2_127_3477_n2213), 
        .A2(DP_OP_422J2_124_3477_n2083), .Y(DP_OP_422J2_124_3477_n2064) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1210 ( .A1(DP_OP_422J2_124_3477_n1991), 
        .A2(DP_OP_422J2_124_3477_n1997), .Y(DP_OP_422J2_124_3477_n1983) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1467 ( .A1(DP_OP_423J2_125_3477_n2603), 
        .A2(DP_OP_425J2_127_3477_n2260), .Y(DP_OP_425J2_127_3477_n2240) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1914 ( .A1(DP_OP_422J2_124_3477_n2694), 
        .A2(DP_OP_422J2_124_3477_n2700), .Y(DP_OP_422J2_124_3477_n2686) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1715 ( .A1(DP_OP_422J2_124_3477_n2209), 
        .A2(n444), .Y(DP_OP_423J2_125_3477_n2489) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1114 ( .A1(DP_OP_422J2_124_3477_n1903), 
        .A2(DP_OP_422J2_124_3477_n1908), .Y(DP_OP_422J2_124_3477_n1887) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1115 ( .A1(DP_OP_424J2_126_3477_n2869), 
        .A2(DP_OP_422J2_124_3477_n1908), .Y(DP_OP_425J2_127_3477_n1888) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1519 ( .A1(DP_OP_422J2_124_3477_n2299), 
        .A2(DP_OP_422J2_124_3477_n2304), .Y(DP_OP_422J2_124_3477_n2291) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1811 ( .A1(DP_OP_423J2_125_3477_n2031), 
        .A2(n451), .Y(DP_OP_425J2_127_3477_n2581) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1111 ( .A1(DP_OP_424J2_126_3477_n2865), 
        .A2(DP_OP_422J2_124_3477_n1908), .Y(DP_OP_425J2_127_3477_n1884) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1504 ( .A1(DP_OP_423J2_125_3477_n2428), 
        .A2(DP_OP_422J2_124_3477_n2302), .Y(DP_OP_422J2_124_3477_n2276) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1625 ( .A1(DP_OP_422J2_124_3477_n2295), 
        .A2(DP_OP_423J2_125_3477_n2430), .Y(DP_OP_423J2_125_3477_n2399) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1510 ( .A1(DP_OP_424J2_126_3477_n2472), 
        .A2(DP_OP_425J2_127_3477_n2304), .Y(DP_OP_425J2_127_3477_n2283) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1555 ( .A1(DP_OP_422J2_124_3477_n2343), 
        .A2(DP_OP_422J2_124_3477_n2347), .Y(DP_OP_422J2_124_3477_n2327) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1811 ( .A1(DP_OP_422J2_124_3477_n2607), 
        .A2(DP_OP_422J2_124_3477_n2610), .Y(DP_OP_422J2_124_3477_n2583) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1713 ( .A1(DP_OP_422J2_124_3477_n2207), 
        .A2(DP_OP_424J2_126_3477_n2520), .Y(DP_OP_423J2_125_3477_n2487) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1635 ( .A1(DP_OP_425J2_127_3477_n2429), 
        .A2(DP_OP_424J2_126_3477_n2432), .Y(DP_OP_425J2_127_3477_n2405) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1473 ( .A1(DP_OP_423J2_125_3477_n2601), 
        .A2(DP_OP_425J2_127_3477_n2261), .Y(DP_OP_425J2_127_3477_n2246) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1599 ( .A1(DP_OP_423J2_125_3477_n2251), 
        .A2(DP_OP_423J2_125_3477_n2387), .Y(DP_OP_425J2_127_3477_n2369) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1335 ( .A1(DP_OP_423J2_125_3477_n2732), 
        .A2(DP_OP_425J2_127_3477_n2128), .Y(DP_OP_425J2_127_3477_n2108) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2036 ( .A1(DP_OP_424J2_126_3477_n1901), 
        .A2(DP_OP_425J2_127_3477_n2829), .Y(DP_OP_425J2_127_3477_n2806) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1377 ( .A1(DP_OP_425J2_127_3477_n2469), 
        .A2(DP_OP_423J2_125_3477_n2168), .Y(DP_OP_423J2_125_3477_n2151) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1385 ( .A1(DP_OP_425J2_127_3477_n2166), 
        .A2(DP_OP_425J2_127_3477_n2173), .Y(DP_OP_425J2_127_3477_n2158) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1860 ( .A1(DP_OP_425J2_127_3477_n2646), 
        .A2(DP_OP_423J2_125_3477_n2651), .Y(DP_OP_425J2_127_3477_n2630) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1632 ( .A1(DP_OP_422J2_124_3477_n2560), 
        .A2(DP_OP_424J2_126_3477_n2432), .Y(DP_OP_425J2_127_3477_n2402) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1388 ( .A1(DP_OP_422J2_124_3477_n2168), 
        .A2(DP_OP_425J2_127_3477_n2173), .Y(DP_OP_422J2_124_3477_n2160) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1254 ( .A1(DP_OP_424J2_126_3477_n2604), 
        .A2(DP_OP_422J2_124_3477_n2040), .Y(DP_OP_422J2_124_3477_n2026) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1463 ( .A1(DP_OP_425J2_127_3477_n2252), 
        .A2(DP_OP_425J2_127_3477_n2260), .Y(DP_OP_425J2_127_3477_n2236) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1168 ( .A1(DP_OP_422J2_124_3477_n1949), 
        .A2(DP_OP_424J2_126_3477_n1953), .Y(DP_OP_422J2_124_3477_n1941) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1331 ( .A1(DP_OP_425J2_127_3477_n2120), 
        .A2(DP_OP_425J2_127_3477_n2128), .Y(DP_OP_425J2_127_3477_n2104) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1476 ( .A1(DP_OP_424J2_126_3477_n2386), 
        .A2(DP_OP_422J2_124_3477_n2260), .Y(DP_OP_422J2_124_3477_n2248) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1239 ( .A1(DP_OP_422J2_124_3477_n1904), 
        .A2(DP_OP_425J2_127_3477_n2039), .Y(DP_OP_425J2_127_3477_n2012) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1237 ( .A1(DP_OP_424J2_126_3477_n2735), 
        .A2(DP_OP_425J2_127_3477_n2039), .Y(DP_OP_425J2_127_3477_n2010) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1723 ( .A1(DP_OP_422J2_124_3477_n2651), 
        .A2(n444), .Y(DP_OP_425J2_127_3477_n2493) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1511 ( .A1(DP_OP_425J2_127_3477_n2300), 
        .A2(DP_OP_425J2_127_3477_n2304), .Y(DP_OP_425J2_127_3477_n2284) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1238 ( .A1(DP_OP_423J2_125_3477_n2028), 
        .A2(DP_OP_425J2_127_3477_n2040), .Y(DP_OP_423J2_125_3477_n2012) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1244 ( .A1(DP_OP_425J2_127_3477_n2033), 
        .A2(DP_OP_425J2_127_3477_n2040), .Y(DP_OP_425J2_127_3477_n2017) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1864 ( .A1(DP_OP_425J2_127_3477_n2650), 
        .A2(DP_OP_424J2_126_3477_n2653), .Y(DP_OP_425J2_127_3477_n2634) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1721 ( .A1(DP_OP_423J2_125_3477_n2117), 
        .A2(n444), .Y(DP_OP_425J2_127_3477_n2491) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1420 ( .A1(DP_OP_425J2_127_3477_n2209), 
        .A2(DP_OP_423J2_125_3477_n2211), .Y(DP_OP_425J2_127_3477_n2193) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1820 ( .A1(DP_OP_424J2_126_3477_n2125), 
        .A2(DP_OP_422J2_124_3477_n2611), .Y(DP_OP_425J2_127_3477_n2590) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1298 ( .A1(DP_OP_425J2_127_3477_n2079), 
        .A2(DP_OP_424J2_126_3477_n2085), .Y(DP_OP_425J2_127_3477_n2071) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1493 ( .A1(DP_OP_423J2_125_3477_n2291), 
        .A2(DP_OP_423J2_125_3477_n2298), .Y(DP_OP_423J2_125_3477_n2267) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1361 ( .A1(DP_OP_425J2_127_3477_n2469), 
        .A2(n452), .Y(DP_OP_423J2_125_3477_n2135) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1519 ( .A1(DP_OP_422J2_124_3477_n2563), 
        .A2(DP_OP_425J2_127_3477_n2305), .Y(DP_OP_424J2_126_3477_n2292) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1116 ( .A1(DP_OP_425J2_127_3477_n1905), 
        .A2(n449), .Y(DP_OP_425J2_127_3477_n1889) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1518 ( .A1(DP_OP_425J2_127_3477_n2428), 
        .A2(n446), .Y(DP_OP_424J2_126_3477_n2291) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1459 ( .A1(DP_OP_424J2_126_3477_n2342), 
        .A2(DP_OP_422J2_124_3477_n2259), .Y(DP_OP_423J2_125_3477_n2233) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1988 ( .A1(DP_OP_423J2_125_3477_n2865), 
        .A2(DP_OP_424J2_126_3477_n2784), .Y(DP_OP_424J2_126_3477_n2758) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1600 ( .A1(DP_OP_425J2_127_3477_n2386), 
        .A2(DP_OP_422J2_124_3477_n2391), .Y(DP_OP_425J2_127_3477_n2370) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1499 ( .A1(DP_OP_424J2_126_3477_n2296), 
        .A2(DP_OP_422J2_124_3477_n2302), .Y(DP_OP_424J2_126_3477_n2272) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1501 ( .A1(DP_OP_423J2_125_3477_n2425), 
        .A2(DP_OP_422J2_124_3477_n2302), .Y(DP_OP_422J2_124_3477_n2273) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1250 ( .A1(DP_OP_423J2_125_3477_n2032), 
        .A2(DP_OP_424J2_126_3477_n2041), .Y(DP_OP_423J2_125_3477_n2024) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1235 ( .A1(DP_OP_422J2_124_3477_n2031), 
        .A2(DP_OP_424J2_126_3477_n2039), .Y(DP_OP_422J2_124_3477_n2007) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1335 ( .A1(DP_OP_424J2_126_3477_n2124), 
        .A2(n440), .Y(DP_OP_424J2_126_3477_n2108) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1818 ( .A1(DP_OP_424J2_126_3477_n2604), 
        .A2(DP_OP_424J2_126_3477_n2609), .Y(DP_OP_424J2_126_3477_n2588) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1511 ( .A1(DP_OP_425J2_127_3477_n2429), 
        .A2(DP_OP_424J2_126_3477_n2304), .Y(DP_OP_424J2_126_3477_n2284) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1599 ( .A1(DP_OP_424J2_126_3477_n2385), 
        .A2(DP_OP_424J2_126_3477_n2389), .Y(DP_OP_424J2_126_3477_n2369) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1804 ( .A1(DP_OP_423J2_125_3477_n2602), 
        .A2(n451), .Y(DP_OP_423J2_125_3477_n2578) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1503 ( .A1(DP_OP_422J2_124_3477_n2473), 
        .A2(DP_OP_423J2_125_3477_n2299), .Y(DP_OP_423J2_125_3477_n2277) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1517 ( .A1(DP_OP_423J2_125_3477_n2205), 
        .A2(n446), .Y(DP_OP_424J2_126_3477_n2290) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1466 ( .A1(DP_OP_424J2_126_3477_n2341), 
        .A2(DP_OP_423J2_125_3477_n2256), .Y(DP_OP_423J2_125_3477_n2240) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1245 ( .A1(DP_OP_422J2_124_3477_n2033), 
        .A2(DP_OP_422J2_124_3477_n2039), .Y(DP_OP_422J2_124_3477_n2017) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1724 ( .A1(DP_OP_423J2_125_3477_n2604), 
        .A2(DP_OP_424J2_126_3477_n2520), .Y(DP_OP_424J2_126_3477_n2494) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1290 ( .A1(DP_OP_425J2_127_3477_n2558), 
        .A2(DP_OP_423J2_125_3477_n2080), .Y(DP_OP_423J2_125_3477_n2064) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1239 ( .A1(DP_OP_423J2_125_3477_n2029), 
        .A2(DP_OP_425J2_127_3477_n2040), .Y(DP_OP_423J2_125_3477_n2013) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1598 ( .A1(DP_OP_424J2_126_3477_n2384), 
        .A2(DP_OP_424J2_126_3477_n2389), .Y(DP_OP_424J2_126_3477_n2368) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1386 ( .A1(DP_OP_423J2_125_3477_n2074), 
        .A2(DP_OP_424J2_126_3477_n2173), .Y(DP_OP_424J2_126_3477_n2159) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1378 ( .A1(DP_OP_423J2_125_3477_n2160), 
        .A2(DP_OP_423J2_125_3477_n2168), .Y(DP_OP_423J2_125_3477_n2152) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1716 ( .A1(DP_OP_422J2_124_3477_n2210), 
        .A2(n444), .Y(DP_OP_423J2_125_3477_n2490) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1206 ( .A1(DP_OP_422J2_124_3477_n2782), 
        .A2(DP_OP_423J2_125_3477_n1992), .Y(DP_OP_423J2_125_3477_n1980) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1115 ( .A1(DP_OP_424J2_126_3477_n1904), 
        .A2(DP_OP_424J2_126_3477_n1908), .Y(DP_OP_424J2_126_3477_n1888) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1596 ( .A1(DP_OP_424J2_126_3477_n2382), 
        .A2(DP_OP_424J2_126_3477_n2389), .Y(DP_OP_424J2_126_3477_n2366) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2039 ( .A1(DP_OP_424J2_126_3477_n2825), 
        .A2(DP_OP_424J2_126_3477_n2829), .Y(DP_OP_424J2_126_3477_n2809) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1423 ( .A1(DP_OP_424J2_126_3477_n2212), 
        .A2(DP_OP_424J2_126_3477_n2216), .Y(DP_OP_424J2_126_3477_n2196) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1810 ( .A1(DP_OP_422J2_124_3477_n2606), 
        .A2(DP_OP_422J2_124_3477_n2610), .Y(DP_OP_422J2_124_3477_n2582) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2119 ( .A1(DP_OP_423J2_125_3477_n2906), 
        .A2(DP_OP_422J2_124_3477_n2917), .Y(DP_OP_423J2_125_3477_n2890) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1636 ( .A1(DP_OP_424J2_126_3477_n2430), 
        .A2(DP_OP_424J2_126_3477_n2432), .Y(DP_OP_424J2_126_3477_n2406) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1247 ( .A1(DP_OP_422J2_124_3477_n2825), 
        .A2(DP_OP_424J2_126_3477_n2040), .Y(DP_OP_424J2_126_3477_n2020) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1729 ( .A1(DP_OP_424J2_126_3477_n2342), 
        .A2(DP_OP_422J2_124_3477_n2523), .Y(DP_OP_422J2_124_3477_n2501) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1510 ( .A1(DP_OP_422J2_124_3477_n2472), 
        .A2(n446), .Y(DP_OP_423J2_125_3477_n2284) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1244 ( .A1(DP_OP_424J2_126_3477_n2033), 
        .A2(DP_OP_424J2_126_3477_n2040), .Y(DP_OP_424J2_126_3477_n2017) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1556 ( .A1(DP_OP_424J2_126_3477_n2430), 
        .A2(DP_OP_425J2_127_3477_n2348), .Y(DP_OP_425J2_127_3477_n2329) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1550 ( .A1(DP_OP_422J2_124_3477_n2432), 
        .A2(DP_OP_423J2_125_3477_n2343), .Y(DP_OP_423J2_125_3477_n2324) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1167 ( .A1(DP_OP_423J2_125_3477_n2908), 
        .A2(DP_OP_425J2_127_3477_n1953), .Y(DP_OP_425J2_127_3477_n1940) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1255 ( .A1(DP_OP_422J2_124_3477_n1904), 
        .A2(DP_OP_425J2_127_3477_n2041), .Y(DP_OP_425J2_127_3477_n2028) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1291 ( .A1(DP_OP_425J2_127_3477_n2649), 
        .A2(DP_OP_424J2_126_3477_n2084), .Y(DP_OP_424J2_126_3477_n2064) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1331 ( .A1(DP_OP_423J2_125_3477_n2599), 
        .A2(DP_OP_422J2_124_3477_n2127), .Y(DP_OP_422J2_124_3477_n2103) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1071 ( .A1(DP_OP_425J2_127_3477_n2869), 
        .A2(DP_OP_422J2_124_3477_n1864), .Y(DP_OP_424J2_126_3477_n1844) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1812 ( .A1(DP_OP_422J2_124_3477_n2036), 
        .A2(DP_OP_424J2_126_3477_n2608), .Y(DP_OP_424J2_126_3477_n2582) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1245 ( .A1(DP_OP_424J2_126_3477_n2034), 
        .A2(DP_OP_424J2_126_3477_n2040), .Y(DP_OP_424J2_126_3477_n2018) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1254 ( .A1(DP_OP_424J2_126_3477_n2035), 
        .A2(DP_OP_424J2_126_3477_n2041), .Y(DP_OP_424J2_126_3477_n2027) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1166 ( .A1(DP_OP_422J2_124_3477_n2912), 
        .A2(DP_OP_424J2_126_3477_n1953), .Y(DP_OP_424J2_126_3477_n1939) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1066 ( .A1(DP_OP_423J2_125_3477_n1856), 
        .A2(DP_OP_423J2_125_3477_n1859), .Y(DP_OP_423J2_125_3477_n1840) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1728 ( .A1(DP_OP_425J2_127_3477_n2382), 
        .A2(DP_OP_422J2_124_3477_n2523), .Y(DP_OP_422J2_124_3477_n2500) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1421 ( .A1(DP_OP_422J2_124_3477_n2649), 
        .A2(DP_OP_424J2_126_3477_n2216), .Y(DP_OP_424J2_126_3477_n2194) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1239 ( .A1(DP_OP_422J2_124_3477_n2825), 
        .A2(DP_OP_424J2_126_3477_n2039), .Y(DP_OP_424J2_126_3477_n2012) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1252 ( .A1(DP_OP_424J2_126_3477_n2033), 
        .A2(DP_OP_424J2_126_3477_n2041), .Y(DP_OP_424J2_126_3477_n2025) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1863 ( .A1(DP_OP_424J2_126_3477_n2649), 
        .A2(DP_OP_424J2_126_3477_n2653), .Y(DP_OP_424J2_126_3477_n2633) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2038 ( .A1(DP_OP_424J2_126_3477_n2824), 
        .A2(DP_OP_424J2_126_3477_n2829), .Y(DP_OP_424J2_126_3477_n2808) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1069 ( .A1(DP_OP_424J2_126_3477_n1858), 
        .A2(DP_OP_422J2_124_3477_n1864), .Y(DP_OP_424J2_126_3477_n1842) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1388 ( .A1(DP_OP_425J2_127_3477_n2169), 
        .A2(DP_OP_425J2_127_3477_n2173), .Y(DP_OP_425J2_127_3477_n2161) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1470 ( .A1(DP_OP_425J2_127_3477_n2386), 
        .A2(DP_OP_423J2_125_3477_n2256), .Y(DP_OP_423J2_125_3477_n2244) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1334 ( .A1(DP_OP_423J2_125_3477_n2030), 
        .A2(n440), .Y(DP_OP_424J2_126_3477_n2107) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1914 ( .A1(DP_OP_425J2_127_3477_n2079), 
        .A2(DP_OP_424J2_126_3477_n2698), .Y(DP_OP_424J2_126_3477_n2684) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1162 ( .A1(DP_OP_425J2_127_3477_n2694), 
        .A2(DP_OP_423J2_125_3477_n1948), .Y(DP_OP_423J2_125_3477_n1936) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1382 ( .A1(DP_OP_423J2_125_3477_n2164), 
        .A2(DP_OP_423J2_125_3477_n2168), .Y(DP_OP_423J2_125_3477_n2156) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1731 ( .A1(DP_OP_424J2_126_3477_n2517), 
        .A2(DP_OP_424J2_126_3477_n2521), .Y(DP_OP_424J2_126_3477_n2501) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1819 ( .A1(DP_OP_422J2_124_3477_n2035), 
        .A2(DP_OP_424J2_126_3477_n2609), .Y(DP_OP_424J2_126_3477_n2589) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1635 ( .A1(DP_OP_422J2_124_3477_n2211), 
        .A2(DP_OP_424J2_126_3477_n2432), .Y(DP_OP_424J2_126_3477_n2405) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1296 ( .A1(DP_OP_424J2_126_3477_n2077), 
        .A2(DP_OP_424J2_126_3477_n2085), .Y(DP_OP_424J2_126_3477_n2069) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1288 ( .A1(DP_OP_422J2_124_3477_n2076), 
        .A2(DP_OP_422J2_124_3477_n2083), .Y(DP_OP_422J2_124_3477_n2060) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1504 ( .A1(DP_OP_425J2_127_3477_n2430), 
        .A2(n445), .Y(DP_OP_424J2_126_3477_n2277) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1287 ( .A1(DP_OP_423J2_125_3477_n2643), 
        .A2(DP_OP_422J2_124_3477_n2083), .Y(DP_OP_422J2_124_3477_n2059) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1385 ( .A1(DP_OP_423J2_125_3477_n2073), 
        .A2(DP_OP_424J2_126_3477_n2173), .Y(DP_OP_424J2_126_3477_n2158) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1210 ( .A1(DP_OP_423J2_125_3477_n1898), 
        .A2(DP_OP_422J2_124_3477_n1997), .Y(DP_OP_424J2_126_3477_n1983) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1424 ( .A1(DP_OP_425J2_127_3477_n2213), 
        .A2(DP_OP_422J2_124_3477_n2215), .Y(DP_OP_425J2_127_3477_n2197) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1555 ( .A1(DP_OP_424J2_126_3477_n2344), 
        .A2(DP_OP_422J2_124_3477_n2347), .Y(DP_OP_424J2_126_3477_n2328) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1475 ( .A1(DP_OP_424J2_126_3477_n2517), 
        .A2(DP_OP_425J2_127_3477_n2261), .Y(DP_OP_425J2_127_3477_n2248) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1336 ( .A1(DP_OP_423J2_125_3477_n2733), 
        .A2(DP_OP_425J2_127_3477_n2128), .Y(DP_OP_425J2_127_3477_n2109) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1367 ( .A1(DP_OP_424J2_126_3477_n2164), 
        .A2(DP_OP_424J2_126_3477_n2171), .Y(DP_OP_424J2_126_3477_n2140) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1387 ( .A1(DP_OP_425J2_127_3477_n2168), 
        .A2(DP_OP_425J2_127_3477_n2173), .Y(DP_OP_425J2_127_3477_n2160) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1466 ( .A1(DP_OP_422J2_124_3477_n2606), 
        .A2(DP_OP_424J2_126_3477_n2260), .Y(DP_OP_424J2_126_3477_n2239) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1809 ( .A1(DP_OP_422J2_124_3477_n2605), 
        .A2(DP_OP_422J2_124_3477_n2610), .Y(DP_OP_422J2_124_3477_n2581) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1372 ( .A1(DP_OP_423J2_125_3477_n2076), 
        .A2(DP_OP_424J2_126_3477_n2171), .Y(DP_OP_424J2_126_3477_n2145) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1248 ( .A1(DP_OP_422J2_124_3477_n1905), 
        .A2(DP_OP_425J2_127_3477_n2040), .Y(DP_OP_425J2_127_3477_n2021) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1240 ( .A1(DP_OP_424J2_126_3477_n2037), 
        .A2(DP_OP_424J2_126_3477_n2039), .Y(DP_OP_424J2_126_3477_n2013) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1370 ( .A1(DP_OP_423J2_125_3477_n2074), 
        .A2(DP_OP_424J2_126_3477_n2171), .Y(DP_OP_424J2_126_3477_n2143) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1468 ( .A1(DP_OP_423J2_125_3477_n2604), 
        .A2(DP_OP_425J2_127_3477_n2260), .Y(DP_OP_425J2_127_3477_n2241) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1500 ( .A1(DP_OP_423J2_125_3477_n2424), 
        .A2(DP_OP_422J2_124_3477_n2302), .Y(DP_OP_422J2_124_3477_n2272) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1467 ( .A1(DP_OP_422J2_124_3477_n2607), 
        .A2(DP_OP_424J2_126_3477_n2260), .Y(DP_OP_424J2_126_3477_n2240) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1502 ( .A1(DP_OP_422J2_124_3477_n2562), 
        .A2(n445), .Y(DP_OP_424J2_126_3477_n2275) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1981 ( .A1(DP_OP_423J2_125_3477_n2776), 
        .A2(DP_OP_423J2_125_3477_n2779), .Y(DP_OP_423J2_125_3477_n2752) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1504 ( .A1(DP_OP_423J2_125_3477_n2294), 
        .A2(DP_OP_423J2_125_3477_n2299), .Y(DP_OP_423J2_125_3477_n2278) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1242 ( .A1(DP_OP_423J2_125_3477_n2032), 
        .A2(DP_OP_424J2_126_3477_n2040), .Y(DP_OP_423J2_125_3477_n2016) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1108 ( .A1(DP_OP_423J2_125_3477_n1898), 
        .A2(DP_OP_424J2_126_3477_n1908), .Y(DP_OP_423J2_125_3477_n1882) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1203 ( .A1(DP_OP_423J2_125_3477_n1985), 
        .A2(DP_OP_423J2_125_3477_n1992), .Y(DP_OP_423J2_125_3477_n1977) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1291 ( .A1(DP_OP_423J2_125_3477_n2073), 
        .A2(DP_OP_423J2_125_3477_n2080), .Y(DP_OP_423J2_125_3477_n2065) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2034 ( .A1(DP_OP_422J2_124_3477_n1905), 
        .A2(DP_OP_423J2_125_3477_n2824), .Y(DP_OP_423J2_125_3477_n2805) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1629 ( .A1(DP_OP_422J2_124_3477_n2299), 
        .A2(DP_OP_423J2_125_3477_n2430), .Y(DP_OP_423J2_125_3477_n2403) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1594 ( .A1(DP_OP_422J2_124_3477_n2344), 
        .A2(DP_OP_423J2_125_3477_n2387), .Y(DP_OP_423J2_125_3477_n2368) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1328 ( .A1(DP_OP_424J2_126_3477_n2211), 
        .A2(n440), .Y(DP_OP_423J2_125_3477_n2102) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1910 ( .A1(DP_OP_425J2_127_3477_n2169), 
        .A2(DP_OP_423J2_125_3477_n2696), .Y(DP_OP_423J2_125_3477_n2684) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1513 ( .A1(DP_OP_423J2_125_3477_n2295), 
        .A2(n446), .Y(DP_OP_423J2_125_3477_n2287) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2032 ( .A1(DP_OP_422J2_124_3477_n1903), 
        .A2(DP_OP_423J2_125_3477_n2824), .Y(DP_OP_423J2_125_3477_n2803) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1332 ( .A1(DP_OP_423J2_125_3477_n2028), 
        .A2(n440), .Y(DP_OP_424J2_126_3477_n2105) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1209 ( .A1(DP_OP_423J2_125_3477_n1897), 
        .A2(DP_OP_422J2_124_3477_n1997), .Y(DP_OP_424J2_126_3477_n1982) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1467 ( .A1(DP_OP_424J2_126_3477_n2342), 
        .A2(DP_OP_423J2_125_3477_n2256), .Y(DP_OP_423J2_125_3477_n2241) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1469 ( .A1(DP_OP_423J2_125_3477_n2251), 
        .A2(DP_OP_423J2_125_3477_n2256), .Y(DP_OP_423J2_125_3477_n2243) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1502 ( .A1(DP_OP_422J2_124_3477_n2298), 
        .A2(DP_OP_422J2_124_3477_n2302), .Y(DP_OP_422J2_124_3477_n2274) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1515 ( .A1(DP_OP_422J2_124_3477_n2295), 
        .A2(DP_OP_422J2_124_3477_n2304), .Y(DP_OP_422J2_124_3477_n2287) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2122 ( .A1(DP_OP_423J2_125_3477_n2909), 
        .A2(DP_OP_424J2_126_3477_n2917), .Y(DP_OP_423J2_125_3477_n2893) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1253 ( .A1(DP_OP_424J2_126_3477_n2034), 
        .A2(DP_OP_424J2_126_3477_n2041), .Y(DP_OP_424J2_126_3477_n2026) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1861 ( .A1(DP_OP_422J2_124_3477_n2649), 
        .A2(DP_OP_422J2_124_3477_n2655), .Y(DP_OP_422J2_124_3477_n2633) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1862 ( .A1(DP_OP_422J2_124_3477_n1991), 
        .A2(DP_OP_424J2_126_3477_n2653), .Y(DP_OP_424J2_126_3477_n2632) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2036 ( .A1(DP_OP_424J2_126_3477_n2822), 
        .A2(DP_OP_424J2_126_3477_n2829), .Y(DP_OP_424J2_126_3477_n2806) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1365 ( .A1(DP_OP_423J2_125_3477_n2163), 
        .A2(n452), .Y(DP_OP_423J2_125_3477_n2139) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1553 ( .A1(DP_OP_422J2_124_3477_n2341), 
        .A2(DP_OP_422J2_124_3477_n2347), .Y(DP_OP_422J2_124_3477_n2325) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1371 ( .A1(DP_OP_424J2_126_3477_n2168), 
        .A2(DP_OP_424J2_126_3477_n2171), .Y(DP_OP_424J2_126_3477_n2144) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1237 ( .A1(DP_OP_424J2_126_3477_n2034), 
        .A2(DP_OP_424J2_126_3477_n2039), .Y(DP_OP_424J2_126_3477_n2010) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1296 ( .A1(DP_OP_422J2_124_3477_n2076), 
        .A2(DP_OP_424J2_126_3477_n2085), .Y(DP_OP_422J2_124_3477_n2068) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1381 ( .A1(DP_OP_423J2_125_3477_n2163), 
        .A2(DP_OP_423J2_125_3477_n2168), .Y(DP_OP_423J2_125_3477_n2155) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1284 ( .A1(DP_OP_423J2_125_3477_n2074), 
        .A2(DP_OP_425J2_127_3477_n2084), .Y(DP_OP_423J2_125_3477_n2058) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1516 ( .A1(DP_OP_423J2_125_3477_n2424), 
        .A2(DP_OP_422J2_124_3477_n2304), .Y(DP_OP_422J2_124_3477_n2288) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1462 ( .A1(DP_OP_422J2_124_3477_n2520), 
        .A2(DP_OP_424J2_126_3477_n2260), .Y(DP_OP_423J2_125_3477_n2236) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1719 ( .A1(DP_OP_423J2_125_3477_n2599), 
        .A2(DP_OP_424J2_126_3477_n2520), .Y(DP_OP_424J2_126_3477_n2489) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1418 ( .A1(DP_OP_425J2_127_3477_n2430), 
        .A2(DP_OP_423J2_125_3477_n2211), .Y(DP_OP_423J2_125_3477_n2192) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1503 ( .A1(DP_OP_425J2_127_3477_n2429), 
        .A2(DP_OP_422J2_124_3477_n2302), .Y(DP_OP_424J2_126_3477_n2276) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2035 ( .A1(DP_OP_424J2_126_3477_n2032), 
        .A2(DP_OP_424J2_126_3477_n2829), .Y(DP_OP_422J2_124_3477_n2805) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1633 ( .A1(DP_OP_422J2_124_3477_n2209), 
        .A2(DP_OP_424J2_126_3477_n2432), .Y(DP_OP_424J2_126_3477_n2403) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1064 ( .A1(DP_OP_425J2_127_3477_n2780), 
        .A2(DP_OP_423J2_125_3477_n1859), .Y(DP_OP_423J2_125_3477_n1838) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1161 ( .A1(DP_OP_423J2_125_3477_n1943), 
        .A2(DP_OP_423J2_125_3477_n1948), .Y(DP_OP_423J2_125_3477_n1935) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1987 ( .A1(DP_OP_425J2_127_3477_n1992), 
        .A2(DP_OP_424J2_126_3477_n2784), .Y(DP_OP_424J2_126_3477_n2757) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2120 ( .A1(DP_OP_423J2_125_3477_n2907), 
        .A2(DP_OP_424J2_126_3477_n2917), .Y(DP_OP_423J2_125_3477_n2891) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1722 ( .A1(DP_OP_422J2_124_3477_n2518), 
        .A2(DP_OP_422J2_124_3477_n2522), .Y(DP_OP_422J2_124_3477_n2494) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1497 ( .A1(DP_OP_423J2_125_3477_n2295), 
        .A2(DP_OP_423J2_125_3477_n2298), .Y(DP_OP_423J2_125_3477_n2271) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1812 ( .A1(DP_OP_423J2_125_3477_n2602), 
        .A2(DP_OP_423J2_125_3477_n2607), .Y(DP_OP_423J2_125_3477_n2586) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1420 ( .A1(DP_OP_422J2_124_3477_n2648), 
        .A2(DP_OP_424J2_126_3477_n2216), .Y(DP_OP_424J2_126_3477_n2193) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1463 ( .A1(DP_OP_424J2_126_3477_n2381), 
        .A2(DP_OP_422J2_124_3477_n2259), .Y(DP_OP_422J2_124_3477_n2235) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1508 ( .A1(DP_OP_423J2_125_3477_n2204), 
        .A2(DP_OP_424J2_126_3477_n2304), .Y(DP_OP_424J2_126_3477_n2281) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1907 ( .A1(DP_OP_425J2_127_3477_n2166), 
        .A2(DP_OP_423J2_125_3477_n2696), .Y(DP_OP_423J2_125_3477_n2681) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1235 ( .A1(DP_OP_424J2_126_3477_n2032), 
        .A2(DP_OP_424J2_126_3477_n2039), .Y(DP_OP_424J2_126_3477_n2008) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1247 ( .A1(DP_OP_423J2_125_3477_n2029), 
        .A2(DP_OP_424J2_126_3477_n2041), .Y(DP_OP_423J2_125_3477_n2021) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1721 ( .A1(DP_OP_423J2_125_3477_n2601), 
        .A2(DP_OP_424J2_126_3477_n2520), .Y(DP_OP_424J2_126_3477_n2491) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1112 ( .A1(DP_OP_424J2_126_3477_n1901), 
        .A2(DP_OP_424J2_126_3477_n1908), .Y(DP_OP_424J2_126_3477_n1885) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2124 ( .A1(DP_OP_424J2_126_3477_n2910), 
        .A2(DP_OP_424J2_126_3477_n2917), .Y(DP_OP_424J2_126_3477_n2894) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1913 ( .A1(DP_OP_424J2_126_3477_n2691), 
        .A2(DP_OP_424J2_126_3477_n2698), .Y(DP_OP_424J2_126_3477_n2683) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1811 ( .A1(DP_OP_422J2_124_3477_n2035), 
        .A2(DP_OP_424J2_126_3477_n2608), .Y(DP_OP_424J2_126_3477_n2581) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1370 ( .A1(DP_OP_423J2_125_3477_n2558), 
        .A2(DP_OP_422J2_124_3477_n2170), .Y(DP_OP_422J2_124_3477_n2142) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1289 ( .A1(DP_OP_423J2_125_3477_n2645), 
        .A2(DP_OP_422J2_124_3477_n2083), .Y(DP_OP_422J2_124_3477_n2061) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1730 ( .A1(DP_OP_423J2_125_3477_n2602), 
        .A2(DP_OP_424J2_126_3477_n2521), .Y(DP_OP_424J2_126_3477_n2500) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1724 ( .A1(DP_OP_424J2_126_3477_n2428), 
        .A2(DP_OP_423J2_125_3477_n2519), .Y(DP_OP_423J2_125_3477_n2498) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1909 ( .A1(DP_OP_425J2_127_3477_n2168), 
        .A2(DP_OP_423J2_125_3477_n2696), .Y(DP_OP_423J2_125_3477_n2683) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2127 ( .A1(DP_OP_425J2_127_3477_n1860), 
        .A2(DP_OP_424J2_126_3477_n2917), .Y(DP_OP_424J2_126_3477_n2897) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2128 ( .A1(DP_OP_425J2_127_3477_n2914), 
        .A2(DP_OP_425J2_127_3477_n2917), .Y(DP_OP_425J2_127_3477_n2898) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1249 ( .A1(DP_OP_423J2_125_3477_n2031), 
        .A2(DP_OP_422J2_124_3477_n2040), .Y(DP_OP_423J2_125_3477_n2023) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1292 ( .A1(DP_OP_423J2_125_3477_n2777), 
        .A2(DP_OP_425J2_127_3477_n2084), .Y(DP_OP_425J2_127_3477_n2065) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1631 ( .A1(DP_OP_422J2_124_3477_n2207), 
        .A2(DP_OP_424J2_126_3477_n2432), .Y(DP_OP_424J2_126_3477_n2401) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1252 ( .A1(DP_OP_422J2_124_3477_n2032), 
        .A2(DP_OP_422J2_124_3477_n2040), .Y(DP_OP_422J2_124_3477_n2024) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1856 ( .A1(DP_OP_423J2_125_3477_n2646), 
        .A2(DP_OP_423J2_125_3477_n2651), .Y(DP_OP_423J2_125_3477_n2630) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1240 ( .A1(DP_OP_423J2_125_3477_n2030), 
        .A2(DP_OP_424J2_126_3477_n2040), .Y(DP_OP_423J2_125_3477_n2014) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1286 ( .A1(DP_OP_423J2_125_3477_n2076), 
        .A2(DP_OP_422J2_124_3477_n2083), .Y(DP_OP_423J2_125_3477_n2060) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1333 ( .A1(DP_OP_422J2_124_3477_n2121), 
        .A2(DP_OP_422J2_124_3477_n2127), .Y(DP_OP_422J2_124_3477_n2105) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2040 ( .A1(DP_OP_425J2_127_3477_n2826), 
        .A2(DP_OP_425J2_127_3477_n2829), .Y(DP_OP_425J2_127_3477_n2810) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1379 ( .A1(DP_OP_423J2_125_3477_n2161), 
        .A2(DP_OP_423J2_125_3477_n2168), .Y(DP_OP_423J2_125_3477_n2153) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1732 ( .A1(DP_OP_425J2_127_3477_n2518), 
        .A2(DP_OP_423J2_125_3477_n2519), .Y(DP_OP_425J2_127_3477_n2502) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1416 ( .A1(DP_OP_422J2_124_3477_n2562), 
        .A2(DP_OP_423J2_125_3477_n2211), .Y(DP_OP_423J2_125_3477_n2190) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1814 ( .A1(DP_OP_423J2_125_3477_n2604), 
        .A2(DP_OP_423J2_125_3477_n2607), .Y(DP_OP_423J2_125_3477_n2588) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1070 ( .A1(DP_OP_425J2_127_3477_n2868), 
        .A2(DP_OP_425J2_127_3477_n1864), .Y(DP_OP_424J2_126_3477_n1843) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1474 ( .A1(DP_OP_422J2_124_3477_n2606), 
        .A2(DP_OP_423J2_125_3477_n2256), .Y(DP_OP_424J2_126_3477_n2247) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1519 ( .A1(DP_OP_425J2_127_3477_n2300), 
        .A2(DP_OP_425J2_127_3477_n2305), .Y(DP_OP_425J2_127_3477_n2292) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1512 ( .A1(DP_OP_422J2_124_3477_n2168), 
        .A2(DP_OP_425J2_127_3477_n2304), .Y(DP_OP_425J2_127_3477_n2285) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1460 ( .A1(DP_OP_422J2_124_3477_n2518), 
        .A2(DP_OP_425J2_127_3477_n2260), .Y(DP_OP_423J2_125_3477_n2234) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1113 ( .A1(DP_OP_422J2_124_3477_n1902), 
        .A2(DP_OP_422J2_124_3477_n1908), .Y(DP_OP_422J2_124_3477_n1886) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1233 ( .A1(DP_OP_423J2_125_3477_n2031), 
        .A2(DP_OP_423J2_125_3477_n2034), .Y(DP_OP_423J2_125_3477_n2007) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1983 ( .A1(DP_OP_424J2_126_3477_n2777), 
        .A2(DP_OP_424J2_126_3477_n2784), .Y(DP_OP_424J2_126_3477_n2753) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1548 ( .A1(DP_OP_422J2_124_3477_n2430), 
        .A2(DP_OP_423J2_125_3477_n2343), .Y(DP_OP_423J2_125_3477_n2322) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1069 ( .A1(DP_OP_422J2_124_3477_n1858), 
        .A2(DP_OP_422J2_124_3477_n1864), .Y(DP_OP_422J2_124_3477_n1842) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1514 ( .A1(DP_OP_422J2_124_3477_n2476), 
        .A2(DP_OP_422J2_124_3477_n2304), .Y(DP_OP_423J2_125_3477_n2288) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1554 ( .A1(DP_OP_422J2_124_3477_n2518), 
        .A2(DP_OP_423J2_125_3477_n2343), .Y(DP_OP_424J2_126_3477_n2327) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1817 ( .A1(DP_OP_422J2_124_3477_n2605), 
        .A2(DP_OP_422J2_124_3477_n2611), .Y(DP_OP_422J2_124_3477_n2589) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1511 ( .A1(DP_OP_422J2_124_3477_n2473), 
        .A2(DP_OP_425J2_127_3477_n2305), .Y(DP_OP_423J2_125_3477_n2285) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1986 ( .A1(DP_OP_422J2_124_3477_n2780), 
        .A2(DP_OP_422J2_124_3477_n2784), .Y(DP_OP_422J2_124_3477_n2756) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1297 ( .A1(DP_OP_424J2_126_3477_n2078), 
        .A2(DP_OP_424J2_126_3477_n2085), .Y(DP_OP_424J2_126_3477_n2070) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1294 ( .A1(DP_OP_423J2_125_3477_n2076), 
        .A2(DP_OP_423J2_125_3477_n2080), .Y(DP_OP_423J2_125_3477_n2068) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1211 ( .A1(DP_OP_425J2_127_3477_n1992), 
        .A2(DP_OP_425J2_127_3477_n1997), .Y(DP_OP_425J2_127_3477_n1984) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1592 ( .A1(DP_OP_422J2_124_3477_n2342), 
        .A2(DP_OP_423J2_125_3477_n2387), .Y(DP_OP_423J2_125_3477_n2366) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1807 ( .A1(DP_OP_422J2_124_3477_n2031), 
        .A2(DP_OP_424J2_126_3477_n2608), .Y(DP_OP_424J2_126_3477_n2577) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1159 ( .A1(DP_OP_425J2_127_3477_n2691), 
        .A2(DP_OP_423J2_125_3477_n1948), .Y(DP_OP_423J2_125_3477_n1933) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1858 ( .A1(DP_OP_423J2_125_3477_n2648), 
        .A2(DP_OP_423J2_125_3477_n2651), .Y(DP_OP_423J2_125_3477_n2632) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1726 ( .A1(DP_OP_423J2_125_3477_n2516), 
        .A2(DP_OP_423J2_125_3477_n2519), .Y(DP_OP_423J2_125_3477_n2500) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1205 ( .A1(DP_OP_425J2_127_3477_n2649), 
        .A2(DP_OP_423J2_125_3477_n1992), .Y(DP_OP_423J2_125_3477_n1979) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1072 ( .A1(DP_OP_425J2_127_3477_n1861), 
        .A2(DP_OP_425J2_127_3477_n1864), .Y(DP_OP_425J2_127_3477_n1845) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1293 ( .A1(DP_OP_422J2_124_3477_n2695), 
        .A2(DP_OP_423J2_125_3477_n2080), .Y(DP_OP_423J2_125_3477_n2067) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1912 ( .A1(DP_OP_422J2_124_3477_n2692), 
        .A2(DP_OP_422J2_124_3477_n2700), .Y(DP_OP_422J2_124_3477_n2684) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1805 ( .A1(DP_OP_423J2_125_3477_n2603), 
        .A2(DP_OP_422J2_124_3477_n2610), .Y(DP_OP_423J2_125_3477_n2579) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1299 ( .A1(DP_OP_423J2_125_3477_n2776), 
        .A2(n441), .Y(DP_OP_425J2_127_3477_n2072) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1208 ( .A1(DP_OP_422J2_124_3477_n1989), 
        .A2(DP_OP_422J2_124_3477_n1997), .Y(DP_OP_422J2_124_3477_n1981) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1110 ( .A1(DP_OP_425J2_127_3477_n2738), 
        .A2(n449), .Y(DP_OP_423J2_125_3477_n1884) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1165 ( .A1(DP_OP_423J2_125_3477_n1853), 
        .A2(DP_OP_424J2_126_3477_n1953), .Y(DP_OP_424J2_126_3477_n1938) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1506 ( .A1(DP_OP_422J2_124_3477_n2476), 
        .A2(DP_OP_423J2_125_3477_n2299), .Y(DP_OP_423J2_125_3477_n2280) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1721 ( .A1(DP_OP_425J2_127_3477_n2383), 
        .A2(DP_OP_422J2_124_3477_n2522), .Y(DP_OP_422J2_124_3477_n2493) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1330 ( .A1(DP_OP_422J2_124_3477_n2652), 
        .A2(n440), .Y(DP_OP_423J2_125_3477_n2104) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1717 ( .A1(DP_OP_423J2_125_3477_n2515), 
        .A2(DP_OP_422J2_124_3477_n2522), .Y(DP_OP_423J2_125_3477_n2491) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1290 ( .A1(DP_OP_422J2_124_3477_n2780), 
        .A2(DP_OP_424J2_126_3477_n2084), .Y(DP_OP_424J2_126_3477_n2063) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1366 ( .A1(DP_OP_423J2_125_3477_n2164), 
        .A2(n452), .Y(DP_OP_423J2_125_3477_n2140) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1507 ( .A1(DP_OP_422J2_124_3477_n2295), 
        .A2(DP_OP_424J2_126_3477_n2304), .Y(DP_OP_422J2_124_3477_n2279) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1424 ( .A1(DP_OP_425J2_127_3477_n2518), 
        .A2(DP_OP_424J2_126_3477_n2216), .Y(DP_OP_424J2_126_3477_n2197) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1475 ( .A1(DP_OP_422J2_124_3477_n2607), 
        .A2(DP_OP_423J2_125_3477_n2256), .Y(DP_OP_424J2_126_3477_n2248) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1634 ( .A1(DP_OP_422J2_124_3477_n2430), 
        .A2(DP_OP_422J2_124_3477_n2434), .Y(DP_OP_422J2_124_3477_n2406) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1984 ( .A1(DP_OP_424J2_126_3477_n2077), 
        .A2(DP_OP_422J2_124_3477_n2784), .Y(DP_OP_422J2_124_3477_n2754) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1983 ( .A1(DP_OP_422J2_124_3477_n2777), 
        .A2(DP_OP_422J2_124_3477_n2784), .Y(DP_OP_422J2_124_3477_n2753) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1246 ( .A1(DP_OP_424J2_126_3477_n2035), 
        .A2(DP_OP_424J2_126_3477_n2040), .Y(DP_OP_424J2_126_3477_n2019) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1808 ( .A1(DP_OP_422J2_124_3477_n2032), 
        .A2(DP_OP_424J2_126_3477_n2608), .Y(DP_OP_424J2_126_3477_n2578) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1387 ( .A1(DP_OP_424J2_126_3477_n2168), 
        .A2(DP_OP_424J2_126_3477_n2173), .Y(DP_OP_424J2_126_3477_n2160) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1472 ( .A1(DP_OP_424J2_126_3477_n2382), 
        .A2(DP_OP_422J2_124_3477_n2260), .Y(DP_OP_422J2_124_3477_n2244) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1595 ( .A1(DP_OP_422J2_124_3477_n2383), 
        .A2(DP_OP_422J2_124_3477_n2391), .Y(DP_OP_422J2_124_3477_n2367) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1855 ( .A1(DP_OP_423J2_125_3477_n2645), 
        .A2(DP_OP_423J2_125_3477_n2651), .Y(DP_OP_423J2_125_3477_n2629) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1980 ( .A1(DP_OP_423J2_125_3477_n2775), 
        .A2(DP_OP_423J2_125_3477_n2779), .Y(DP_OP_423J2_125_3477_n2751) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1116 ( .A1(DP_OP_425J2_127_3477_n2826), 
        .A2(DP_OP_424J2_126_3477_n1908), .Y(DP_OP_424J2_126_3477_n1889) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1287 ( .A1(DP_OP_423J2_125_3477_n1983), 
        .A2(DP_OP_424J2_126_3477_n2084), .Y(DP_OP_424J2_126_3477_n2060) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1512 ( .A1(DP_OP_425J2_127_3477_n2430), 
        .A2(DP_OP_424J2_126_3477_n2304), .Y(DP_OP_424J2_126_3477_n2285) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1288 ( .A1(DP_OP_424J2_126_3477_n2077), 
        .A2(DP_OP_424J2_126_3477_n2084), .Y(DP_OP_424J2_126_3477_n2061) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2125 ( .A1(DP_OP_425J2_127_3477_n2779), 
        .A2(DP_OP_422J2_124_3477_n2917), .Y(DP_OP_422J2_124_3477_n2895) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1204 ( .A1(DP_OP_423J2_125_3477_n1986), 
        .A2(DP_OP_423J2_125_3477_n1992), .Y(DP_OP_423J2_125_3477_n1978) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1421 ( .A1(DP_OP_422J2_124_3477_n2209), 
        .A2(DP_OP_422J2_124_3477_n2215), .Y(DP_OP_422J2_124_3477_n2193) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2128 ( .A1(DP_OP_425J2_127_3477_n1861), 
        .A2(DP_OP_424J2_126_3477_n2917), .Y(DP_OP_424J2_126_3477_n2898) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1285 ( .A1(DP_OP_424J2_126_3477_n2168), 
        .A2(DP_OP_424J2_126_3477_n2084), .Y(DP_OP_423J2_125_3477_n2059) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1811 ( .A1(DP_OP_423J2_125_3477_n2601), 
        .A2(DP_OP_423J2_125_3477_n2607), .Y(DP_OP_423J2_125_3477_n2585) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1500 ( .A1(DP_OP_422J2_124_3477_n2560), 
        .A2(n445), .Y(DP_OP_424J2_126_3477_n2273) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1857 ( .A1(DP_OP_423J2_125_3477_n2647), 
        .A2(DP_OP_423J2_125_3477_n2651), .Y(DP_OP_423J2_125_3477_n2631) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1816 ( .A1(DP_OP_422J2_124_3477_n2032), 
        .A2(DP_OP_424J2_126_3477_n2609), .Y(DP_OP_424J2_126_3477_n2586) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1982 ( .A1(DP_OP_423J2_125_3477_n2777), 
        .A2(DP_OP_423J2_125_3477_n2779), .Y(DP_OP_423J2_125_3477_n2753) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1906 ( .A1(DP_OP_423J2_125_3477_n2688), 
        .A2(DP_OP_423J2_125_3477_n2696), .Y(DP_OP_423J2_125_3477_n2680) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1067 ( .A1(DP_OP_423J2_125_3477_n2860), 
        .A2(DP_OP_422J2_124_3477_n1864), .Y(DP_OP_422J2_124_3477_n1840) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1505 ( .A1(DP_OP_423J2_125_3477_n2295), 
        .A2(DP_OP_423J2_125_3477_n2299), .Y(DP_OP_423J2_125_3477_n2279) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1723 ( .A1(DP_OP_424J2_126_3477_n2517), 
        .A2(DP_OP_424J2_126_3477_n2520), .Y(DP_OP_424J2_126_3477_n2493) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1063 ( .A1(DP_OP_423J2_125_3477_n1853), 
        .A2(DP_OP_423J2_125_3477_n1859), .Y(DP_OP_423J2_125_3477_n1837) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1246 ( .A1(DP_OP_423J2_125_3477_n2028), 
        .A2(DP_OP_425J2_127_3477_n2041), .Y(DP_OP_423J2_125_3477_n2020) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1593 ( .A1(DP_OP_422J2_124_3477_n2343), 
        .A2(DP_OP_423J2_125_3477_n2387), .Y(DP_OP_423J2_125_3477_n2367) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1723 ( .A1(DP_OP_422J2_124_3477_n2209), 
        .A2(DP_OP_423J2_125_3477_n2519), .Y(DP_OP_423J2_125_3477_n2497) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1547 ( .A1(DP_OP_422J2_124_3477_n2429), 
        .A2(DP_OP_423J2_125_3477_n2343), .Y(DP_OP_423J2_125_3477_n2321) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1333 ( .A1(DP_OP_422J2_124_3477_n2735), 
        .A2(DP_OP_422J2_124_3477_n2127), .Y(DP_OP_424J2_126_3477_n2106) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1727 ( .A1(DP_OP_423J2_125_3477_n2247), 
        .A2(DP_OP_422J2_124_3477_n2523), .Y(DP_OP_422J2_124_3477_n2499) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1911 ( .A1(DP_OP_424J2_126_3477_n2689), 
        .A2(DP_OP_424J2_126_3477_n2698), .Y(DP_OP_424J2_126_3477_n2681) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1498 ( .A1(DP_OP_422J2_124_3477_n2476), 
        .A2(DP_OP_423J2_125_3477_n2298), .Y(DP_OP_423J2_125_3477_n2272) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1329 ( .A1(DP_OP_422J2_124_3477_n2651), 
        .A2(n440), .Y(DP_OP_423J2_125_3477_n2103) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1369 ( .A1(DP_OP_425J2_127_3477_n2559), 
        .A2(DP_OP_424J2_126_3477_n2171), .Y(DP_OP_424J2_126_3477_n2142) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1808 ( .A1(DP_OP_422J2_124_3477_n2604), 
        .A2(DP_OP_422J2_124_3477_n2610), .Y(DP_OP_422J2_124_3477_n2580) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1420 ( .A1(DP_OP_422J2_124_3477_n2208), 
        .A2(DP_OP_422J2_124_3477_n2215), .Y(DP_OP_422J2_124_3477_n2192) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1476 ( .A1(DP_OP_423J2_125_3477_n2604), 
        .A2(DP_OP_425J2_127_3477_n2261), .Y(DP_OP_425J2_127_3477_n2249) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1068 ( .A1(DP_OP_424J2_126_3477_n1857), 
        .A2(DP_OP_423J2_125_3477_n1859), .Y(DP_OP_424J2_126_3477_n1841) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1520 ( .A1(DP_OP_422J2_124_3477_n2168), 
        .A2(DP_OP_425J2_127_3477_n2305), .Y(DP_OP_425J2_127_3477_n2293) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1860 ( .A1(DP_OP_422J2_124_3477_n2648), 
        .A2(DP_OP_422J2_124_3477_n2655), .Y(DP_OP_422J2_124_3477_n2632) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1815 ( .A1(DP_OP_422J2_124_3477_n2603), 
        .A2(DP_OP_422J2_124_3477_n2611), .Y(DP_OP_422J2_124_3477_n2587) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1248 ( .A1(DP_OP_424J2_126_3477_n2037), 
        .A2(DP_OP_424J2_126_3477_n2040), .Y(DP_OP_424J2_126_3477_n2021) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1208 ( .A1(DP_OP_425J2_127_3477_n2734), 
        .A2(DP_OP_423J2_125_3477_n1992), .Y(DP_OP_424J2_126_3477_n1981) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2040 ( .A1(DP_OP_424J2_126_3477_n2826), 
        .A2(DP_OP_424J2_126_3477_n2829), .Y(DP_OP_424J2_126_3477_n2810) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1499 ( .A1(DP_OP_422J2_124_3477_n2295), 
        .A2(DP_OP_422J2_124_3477_n2302), .Y(DP_OP_422J2_124_3477_n2271) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1864 ( .A1(DP_OP_424J2_126_3477_n2650), 
        .A2(DP_OP_424J2_126_3477_n2653), .Y(DP_OP_424J2_126_3477_n2634) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1463 ( .A1(DP_OP_422J2_124_3477_n2603), 
        .A2(DP_OP_424J2_126_3477_n2260), .Y(DP_OP_424J2_126_3477_n2236) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1915 ( .A1(DP_OP_424J2_126_3477_n2693), 
        .A2(DP_OP_424J2_126_3477_n2698), .Y(DP_OP_424J2_126_3477_n2685) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1107 ( .A1(DP_OP_423J2_125_3477_n1897), 
        .A2(DP_OP_422J2_124_3477_n1908), .Y(DP_OP_423J2_125_3477_n1881) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2121 ( .A1(DP_OP_423J2_125_3477_n2908), 
        .A2(DP_OP_425J2_127_3477_n2917), .Y(DP_OP_423J2_125_3477_n2892) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1364 ( .A1(DP_OP_425J2_127_3477_n2472), 
        .A2(n452), .Y(DP_OP_423J2_125_3477_n2138) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1632 ( .A1(DP_OP_422J2_124_3477_n2428), 
        .A2(DP_OP_422J2_124_3477_n2434), .Y(DP_OP_422J2_124_3477_n2404) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1512 ( .A1(DP_OP_423J2_125_3477_n2294), 
        .A2(n446), .Y(DP_OP_423J2_125_3477_n2286) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1725 ( .A1(DP_OP_423J2_125_3477_n2515), 
        .A2(DP_OP_423J2_125_3477_n2519), .Y(DP_OP_423J2_125_3477_n2499) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1820 ( .A1(DP_OP_422J2_124_3477_n2036), 
        .A2(DP_OP_424J2_126_3477_n2609), .Y(DP_OP_424J2_126_3477_n2590) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1468 ( .A1(DP_OP_422J2_124_3477_n2518), 
        .A2(DP_OP_423J2_125_3477_n2256), .Y(DP_OP_423J2_125_3477_n2242) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1556 ( .A1(DP_OP_425J2_127_3477_n2386), 
        .A2(DP_OP_422J2_124_3477_n2347), .Y(DP_OP_424J2_126_3477_n2329) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1984 ( .A1(DP_OP_423J2_125_3477_n2861), 
        .A2(DP_OP_424J2_126_3477_n2784), .Y(DP_OP_424J2_126_3477_n2754) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2031 ( .A1(DP_OP_422J2_124_3477_n1902), 
        .A2(DP_OP_423J2_125_3477_n2824), .Y(DP_OP_423J2_125_3477_n2802) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1815 ( .A1(DP_OP_422J2_124_3477_n2031), 
        .A2(DP_OP_424J2_126_3477_n2609), .Y(DP_OP_424J2_126_3477_n2585) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2033 ( .A1(DP_OP_424J2_126_3477_n2737), 
        .A2(DP_OP_423J2_125_3477_n2824), .Y(DP_OP_423J2_125_3477_n2804) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1255 ( .A1(DP_OP_422J2_124_3477_n2825), 
        .A2(DP_OP_424J2_126_3477_n2041), .Y(DP_OP_424J2_126_3477_n2028) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1368 ( .A1(DP_OP_422J2_124_3477_n2692), 
        .A2(DP_OP_424J2_126_3477_n2171), .Y(DP_OP_424J2_126_3477_n2141) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1109 ( .A1(DP_OP_423J2_125_3477_n1899), 
        .A2(n449), .Y(DP_OP_423J2_125_3477_n1883) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1327 ( .A1(DP_OP_423J2_125_3477_n2117), 
        .A2(DP_OP_425J2_127_3477_n2128), .Y(DP_OP_423J2_125_3477_n2101) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1211 ( .A1(DP_OP_422J2_124_3477_n2869), 
        .A2(DP_OP_425J2_127_3477_n1997), .Y(DP_OP_424J2_126_3477_n1984) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1111 ( .A1(DP_OP_422J2_124_3477_n1900), 
        .A2(DP_OP_422J2_124_3477_n1908), .Y(DP_OP_422J2_124_3477_n1884) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1465 ( .A1(DP_OP_424J2_126_3477_n2383), 
        .A2(DP_OP_422J2_124_3477_n2259), .Y(DP_OP_422J2_124_3477_n2237) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1496 ( .A1(DP_OP_423J2_125_3477_n2294), 
        .A2(DP_OP_423J2_125_3477_n2298), .Y(DP_OP_423J2_125_3477_n2270) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1292 ( .A1(DP_OP_425J2_127_3477_n2650), 
        .A2(DP_OP_424J2_126_3477_n2084), .Y(DP_OP_424J2_126_3477_n2065) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1807 ( .A1(DP_OP_422J2_124_3477_n2603), 
        .A2(DP_OP_422J2_124_3477_n2610), .Y(DP_OP_422J2_124_3477_n2579) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1241 ( .A1(DP_OP_423J2_125_3477_n2031), 
        .A2(DP_OP_425J2_127_3477_n2040), .Y(DP_OP_423J2_125_3477_n2015) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1067 ( .A1(DP_OP_425J2_127_3477_n2865), 
        .A2(DP_OP_423J2_125_3477_n1859), .Y(DP_OP_424J2_126_3477_n1840) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1384 ( .A1(DP_OP_422J2_124_3477_n2164), 
        .A2(DP_OP_424J2_126_3477_n2173), .Y(DP_OP_422J2_124_3477_n2156) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2123 ( .A1(DP_OP_422J2_124_3477_n2909), 
        .A2(DP_OP_422J2_124_3477_n2917), .Y(DP_OP_422J2_124_3477_n2893) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1813 ( .A1(DP_OP_423J2_125_3477_n2603), 
        .A2(DP_OP_423J2_125_3477_n2607), .Y(DP_OP_423J2_125_3477_n2587) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1509 ( .A1(DP_OP_423J2_125_3477_n2425), 
        .A2(DP_OP_424J2_126_3477_n2304), .Y(DP_OP_422J2_124_3477_n2281) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1600 ( .A1(DP_OP_424J2_126_3477_n2386), 
        .A2(DP_OP_424J2_126_3477_n2389), .Y(DP_OP_424J2_126_3477_n2370) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1806 ( .A1(DP_OP_423J2_125_3477_n2604), 
        .A2(DP_OP_424J2_126_3477_n2608), .Y(DP_OP_423J2_125_3477_n2580) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1597 ( .A1(DP_OP_422J2_124_3477_n2385), 
        .A2(DP_OP_422J2_124_3477_n2391), .Y(DP_OP_422J2_124_3477_n2369) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1720 ( .A1(DP_OP_425J2_127_3477_n2382), 
        .A2(DP_OP_422J2_124_3477_n2522), .Y(DP_OP_422J2_124_3477_n2492) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1809 ( .A1(DP_OP_422J2_124_3477_n2033), 
        .A2(DP_OP_424J2_126_3477_n2608), .Y(DP_OP_424J2_126_3477_n2579) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1419 ( .A1(DP_OP_422J2_124_3477_n2207), 
        .A2(DP_OP_422J2_124_3477_n2215), .Y(DP_OP_422J2_124_3477_n2191) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1908 ( .A1(DP_OP_423J2_125_3477_n2690), 
        .A2(DP_OP_423J2_125_3477_n2696), .Y(DP_OP_423J2_125_3477_n2682) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1468 ( .A1(DP_OP_422J2_124_3477_n2608), 
        .A2(DP_OP_424J2_126_3477_n2260), .Y(DP_OP_424J2_126_3477_n2241) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1720 ( .A1(DP_OP_423J2_125_3477_n2600), 
        .A2(DP_OP_424J2_126_3477_n2520), .Y(DP_OP_424J2_126_3477_n2490) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1367 ( .A1(DP_OP_422J2_124_3477_n2163), 
        .A2(DP_OP_422J2_124_3477_n2170), .Y(DP_OP_422J2_124_3477_n2139) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1283 ( .A1(DP_OP_423J2_125_3477_n2073), 
        .A2(DP_OP_422J2_124_3477_n2083), .Y(DP_OP_423J2_125_3477_n2057) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2123 ( .A1(DP_OP_424J2_126_3477_n2909), 
        .A2(DP_OP_424J2_126_3477_n2917), .Y(DP_OP_424J2_126_3477_n2893) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1202 ( .A1(DP_OP_424J2_126_3477_n2077), 
        .A2(DP_OP_423J2_125_3477_n1992), .Y(DP_OP_423J2_125_3477_n1976) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2037 ( .A1(DP_OP_424J2_126_3477_n2034), 
        .A2(DP_OP_423J2_125_3477_n2824), .Y(DP_OP_422J2_124_3477_n2807) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1369 ( .A1(DP_OP_422J2_124_3477_n2165), 
        .A2(DP_OP_422J2_124_3477_n2170), .Y(DP_OP_422J2_124_3477_n2141) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1860 ( .A1(DP_OP_423J2_125_3477_n2729), 
        .A2(DP_OP_424J2_126_3477_n2653), .Y(DP_OP_424J2_126_3477_n2630) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1160 ( .A1(DP_OP_425J2_127_3477_n2692), 
        .A2(DP_OP_423J2_125_3477_n1948), .Y(DP_OP_423J2_125_3477_n1934) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1331 ( .A1(DP_OP_424J2_126_3477_n2120), 
        .A2(DP_OP_422J2_124_3477_n2127), .Y(DP_OP_424J2_126_3477_n2104) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1295 ( .A1(DP_OP_423J2_125_3477_n1983), 
        .A2(DP_OP_424J2_126_3477_n2085), .Y(DP_OP_424J2_126_3477_n2068) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1417 ( .A1(DP_OP_425J2_127_3477_n2429), 
        .A2(DP_OP_423J2_125_3477_n2211), .Y(DP_OP_423J2_125_3477_n2191) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1473 ( .A1(DP_OP_422J2_124_3477_n2605), 
        .A2(DP_OP_425J2_127_3477_n2261), .Y(DP_OP_424J2_126_3477_n2246) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1238 ( .A1(DP_OP_424J2_126_3477_n2604), 
        .A2(DP_OP_424J2_126_3477_n2039), .Y(DP_OP_422J2_124_3477_n2010) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1552 ( .A1(DP_OP_424J2_126_3477_n2341), 
        .A2(DP_OP_423J2_125_3477_n2343), .Y(DP_OP_424J2_126_3477_n2325) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1336 ( .A1(DP_OP_424J2_126_3477_n2125), 
        .A2(DP_OP_425J2_127_3477_n2128), .Y(DP_OP_424J2_126_3477_n2109) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1985 ( .A1(DP_OP_423J2_125_3477_n1985), 
        .A2(DP_OP_422J2_124_3477_n2784), .Y(DP_OP_422J2_124_3477_n2755) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1464 ( .A1(DP_OP_424J2_126_3477_n2382), 
        .A2(DP_OP_422J2_124_3477_n2259), .Y(DP_OP_422J2_124_3477_n2236) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1248 ( .A1(DP_OP_423J2_125_3477_n2030), 
        .A2(DP_OP_424J2_126_3477_n2041), .Y(DP_OP_423J2_125_3477_n2022) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1212 ( .A1(DP_OP_425J2_127_3477_n2738), 
        .A2(DP_OP_423J2_125_3477_n1992), .Y(DP_OP_424J2_126_3477_n1985) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1510 ( .A1(DP_OP_425J2_127_3477_n2428), 
        .A2(DP_OP_424J2_126_3477_n2304), .Y(DP_OP_424J2_126_3477_n2283) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1114 ( .A1(DP_OP_424J2_126_3477_n1903), 
        .A2(DP_OP_424J2_126_3477_n1908), .Y(DP_OP_424J2_126_3477_n1887) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1549 ( .A1(DP_OP_423J2_125_3477_n2339), 
        .A2(DP_OP_423J2_125_3477_n2343), .Y(DP_OP_423J2_125_3477_n2323) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1810 ( .A1(DP_OP_424J2_126_3477_n2604), 
        .A2(DP_OP_424J2_126_3477_n2608), .Y(DP_OP_424J2_126_3477_n2580) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2035 ( .A1(DP_OP_424J2_126_3477_n2821), 
        .A2(DP_OP_424J2_126_3477_n2829), .Y(DP_OP_424J2_126_3477_n2805) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1368 ( .A1(DP_OP_422J2_124_3477_n2164), 
        .A2(DP_OP_422J2_124_3477_n2170), .Y(DP_OP_422J2_124_3477_n2140) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1861 ( .A1(DP_OP_425J2_127_3477_n2122), 
        .A2(DP_OP_424J2_126_3477_n2653), .Y(DP_OP_424J2_126_3477_n2631) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1515 ( .A1(DP_OP_424J2_126_3477_n2296), 
        .A2(n446), .Y(DP_OP_424J2_126_3477_n2288) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1552 ( .A1(DP_OP_422J2_124_3477_n2340), 
        .A2(DP_OP_422J2_124_3477_n2347), .Y(DP_OP_422J2_124_3477_n2324) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1912 ( .A1(DP_OP_425J2_127_3477_n2077), 
        .A2(DP_OP_424J2_126_3477_n2698), .Y(DP_OP_424J2_126_3477_n2682) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1236 ( .A1(DP_OP_424J2_126_3477_n2033), 
        .A2(DP_OP_424J2_126_3477_n2039), .Y(DP_OP_424J2_126_3477_n2009) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1244 ( .A1(DP_OP_422J2_124_3477_n2032), 
        .A2(DP_OP_422J2_124_3477_n2039), .Y(DP_OP_422J2_124_3477_n2016) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1164 ( .A1(DP_OP_425J2_127_3477_n2778), 
        .A2(DP_OP_424J2_126_3477_n1953), .Y(DP_OP_424J2_126_3477_n1937) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1464 ( .A1(DP_OP_422J2_124_3477_n2604), 
        .A2(DP_OP_424J2_126_3477_n2260), .Y(DP_OP_424J2_126_3477_n2237) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1630 ( .A1(DP_OP_423J2_125_3477_n2428), 
        .A2(DP_OP_423J2_125_3477_n2430), .Y(DP_OP_423J2_125_3477_n2404) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1729 ( .A1(DP_OP_422J2_124_3477_n2121), 
        .A2(DP_OP_424J2_126_3477_n2521), .Y(DP_OP_424J2_126_3477_n2499) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1722 ( .A1(DP_OP_423J2_125_3477_n2602), 
        .A2(DP_OP_424J2_126_3477_n2520), .Y(DP_OP_424J2_126_3477_n2492) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1508 ( .A1(DP_OP_423J2_125_3477_n2424), 
        .A2(DP_OP_423J2_125_3477_n2299), .Y(DP_OP_422J2_124_3477_n2280) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1380 ( .A1(DP_OP_425J2_127_3477_n2472), 
        .A2(DP_OP_423J2_125_3477_n2168), .Y(DP_OP_423J2_125_3477_n2154) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1986 ( .A1(DP_OP_425J2_127_3477_n1991), 
        .A2(DP_OP_424J2_126_3477_n2784), .Y(DP_OP_424J2_126_3477_n2756) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1596 ( .A1(DP_OP_422J2_124_3477_n2384), 
        .A2(DP_OP_422J2_124_3477_n2391), .Y(DP_OP_422J2_124_3477_n2368) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1627 ( .A1(DP_OP_423J2_125_3477_n2425), 
        .A2(DP_OP_423J2_125_3477_n2430), .Y(DP_OP_423J2_125_3477_n2401) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1516 ( .A1(DP_OP_422J2_124_3477_n2560), 
        .A2(n446), .Y(DP_OP_424J2_126_3477_n2289) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2125 ( .A1(DP_OP_425J2_127_3477_n1858), 
        .A2(DP_OP_424J2_126_3477_n2917), .Y(DP_OP_424J2_126_3477_n2895) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2036 ( .A1(DP_OP_424J2_126_3477_n2033), 
        .A2(DP_OP_423J2_125_3477_n2824), .Y(DP_OP_422J2_124_3477_n2806) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1632 ( .A1(DP_OP_422J2_124_3477_n2208), 
        .A2(DP_OP_424J2_126_3477_n2432), .Y(DP_OP_424J2_126_3477_n2402) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1461 ( .A1(DP_OP_423J2_125_3477_n2251), 
        .A2(DP_OP_425J2_127_3477_n2260), .Y(DP_OP_423J2_125_3477_n2235) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1292 ( .A1(DP_OP_423J2_125_3477_n2074), 
        .A2(DP_OP_423J2_125_3477_n2080), .Y(DP_OP_423J2_125_3477_n2066) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1985 ( .A1(DP_OP_425J2_127_3477_n1990), 
        .A2(DP_OP_424J2_126_3477_n2784), .Y(DP_OP_424J2_126_3477_n2755) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1237 ( .A1(DP_OP_422J2_124_3477_n2033), 
        .A2(DP_OP_424J2_126_3477_n2039), .Y(DP_OP_422J2_124_3477_n2009) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1383 ( .A1(DP_OP_422J2_124_3477_n2163), 
        .A2(DP_OP_425J2_127_3477_n2173), .Y(DP_OP_422J2_124_3477_n2155) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1112 ( .A1(DP_OP_425J2_127_3477_n2033), 
        .A2(DP_OP_422J2_124_3477_n1908), .Y(DP_OP_422J2_124_3477_n1885) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1859 ( .A1(DP_OP_422J2_124_3477_n2647), 
        .A2(DP_OP_422J2_124_3477_n2655), .Y(DP_OP_422J2_124_3477_n2631) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1068 ( .A1(DP_OP_425J2_127_3477_n1989), 
        .A2(DP_OP_422J2_124_3477_n1864), .Y(DP_OP_422J2_124_3477_n1841) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1212 ( .A1(DP_OP_422J2_124_3477_n1861), 
        .A2(DP_OP_425J2_127_3477_n1997), .Y(DP_OP_425J2_127_3477_n1985) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1065 ( .A1(DP_OP_424J2_126_3477_n1948), 
        .A2(DP_OP_423J2_125_3477_n1859), .Y(DP_OP_423J2_125_3477_n1839) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1472 ( .A1(DP_OP_422J2_124_3477_n2604), 
        .A2(DP_OP_425J2_127_3477_n2261), .Y(DP_OP_424J2_126_3477_n2245) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1634 ( .A1(DP_OP_424J2_126_3477_n2428), 
        .A2(DP_OP_424J2_126_3477_n2432), .Y(DP_OP_424J2_126_3477_n2404) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1728 ( .A1(DP_OP_423J2_125_3477_n2600), 
        .A2(DP_OP_424J2_126_3477_n2521), .Y(DP_OP_424J2_126_3477_n2498) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1167 ( .A1(DP_OP_424J2_126_3477_n1948), 
        .A2(DP_OP_424J2_126_3477_n1953), .Y(DP_OP_424J2_126_3477_n1940) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1732 ( .A1(DP_OP_423J2_125_3477_n2604), 
        .A2(DP_OP_424J2_126_3477_n2521), .Y(DP_OP_424J2_126_3477_n2502) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1111 ( .A1(DP_OP_425J2_127_3477_n2821), 
        .A2(DP_OP_424J2_126_3477_n1908), .Y(DP_OP_424J2_126_3477_n1884) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1072 ( .A1(DP_OP_425J2_127_3477_n2870), 
        .A2(DP_OP_422J2_124_3477_n1864), .Y(DP_OP_424J2_126_3477_n1845) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1507 ( .A1(DP_OP_424J2_126_3477_n2296), 
        .A2(DP_OP_424J2_126_3477_n2304), .Y(DP_OP_424J2_126_3477_n2280) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1238 ( .A1(DP_OP_424J2_126_3477_n2035), 
        .A2(DP_OP_424J2_126_3477_n2039), .Y(DP_OP_424J2_126_3477_n2011) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2037 ( .A1(DP_OP_424J2_126_3477_n2823), 
        .A2(DP_OP_424J2_126_3477_n2829), .Y(DP_OP_424J2_126_3477_n2807) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1419 ( .A1(DP_OP_422J2_124_3477_n2647), 
        .A2(DP_OP_424J2_126_3477_n2216), .Y(DP_OP_424J2_126_3477_n2192) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1332 ( .A1(DP_OP_422J2_124_3477_n2120), 
        .A2(DP_OP_422J2_124_3477_n2127), .Y(DP_OP_422J2_124_3477_n2104) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1299 ( .A1(DP_OP_422J2_124_3477_n2781), 
        .A2(DP_OP_424J2_126_3477_n2085), .Y(DP_OP_424J2_126_3477_n2072) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1298 ( .A1(DP_OP_422J2_124_3477_n2780), 
        .A2(DP_OP_424J2_126_3477_n2085), .Y(DP_OP_424J2_126_3477_n2071) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1465 ( .A1(DP_OP_422J2_124_3477_n2605), 
        .A2(DP_OP_424J2_126_3477_n2260), .Y(DP_OP_424J2_126_3477_n2238) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1384 ( .A1(DP_OP_425J2_127_3477_n2558), 
        .A2(DP_OP_424J2_126_3477_n2173), .Y(DP_OP_424J2_126_3477_n2157) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1501 ( .A1(DP_OP_425J2_127_3477_n2427), 
        .A2(n445), .Y(DP_OP_424J2_126_3477_n2274) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2126 ( .A1(DP_OP_424J2_126_3477_n2912), 
        .A2(DP_OP_424J2_126_3477_n2917), .Y(DP_OP_424J2_126_3477_n2896) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1719 ( .A1(DP_OP_423J2_125_3477_n2247), 
        .A2(DP_OP_422J2_124_3477_n2522), .Y(DP_OP_422J2_124_3477_n2491) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1300 ( .A1(DP_OP_422J2_124_3477_n1949), 
        .A2(n441), .Y(DP_OP_425J2_127_3477_n2073) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1916 ( .A1(DP_OP_425J2_127_3477_n2694), 
        .A2(DP_OP_424J2_126_3477_n2698), .Y(DP_OP_425J2_127_3477_n2686) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1633 ( .A1(DP_OP_422J2_124_3477_n2429), 
        .A2(DP_OP_422J2_124_3477_n2434), .Y(DP_OP_422J2_124_3477_n2405) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1113 ( .A1(DP_OP_425J2_127_3477_n2823), 
        .A2(DP_OP_424J2_126_3477_n1908), .Y(DP_OP_424J2_126_3477_n1886) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1718 ( .A1(DP_OP_423J2_125_3477_n2516), 
        .A2(n444), .Y(DP_OP_423J2_125_3477_n2492) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1520 ( .A1(DP_OP_425J2_127_3477_n2430), 
        .A2(DP_OP_422J2_124_3477_n2304), .Y(DP_OP_424J2_126_3477_n2293) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1509 ( .A1(DP_OP_423J2_125_3477_n2205), 
        .A2(DP_OP_424J2_126_3477_n2304), .Y(DP_OP_424J2_126_3477_n2282) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1234 ( .A1(DP_OP_423J2_125_3477_n2032), 
        .A2(DP_OP_423J2_125_3477_n2034), .Y(DP_OP_423J2_125_3477_n2008) );
  XNOR2X1_HVT DP_OP_422J2_124_3477_U627 ( .A1(DP_OP_422J2_124_3477_n2002), 
        .A2(DP_OP_422J2_124_3477_n2703), .Y(DP_OP_422J2_124_3477_n1062) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1816 ( .A1(DP_OP_422J2_124_3477_n2604), 
        .A2(DP_OP_422J2_124_3477_n2611), .Y(DP_OP_422J2_124_3477_n2588) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1817 ( .A1(DP_OP_422J2_124_3477_n2033), 
        .A2(DP_OP_424J2_126_3477_n2609), .Y(DP_OP_424J2_126_3477_n2587) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1553 ( .A1(DP_OP_424J2_126_3477_n2342), 
        .A2(DP_OP_422J2_124_3477_n2347), .Y(DP_OP_424J2_126_3477_n2326) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1256 ( .A1(DP_OP_424J2_126_3477_n2037), 
        .A2(DP_OP_424J2_126_3477_n2041), .Y(DP_OP_424J2_126_3477_n2029) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2124 ( .A1(DP_OP_425J2_127_3477_n2778), 
        .A2(DP_OP_422J2_124_3477_n2917), .Y(DP_OP_422J2_124_3477_n2894) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1168 ( .A1(DP_OP_423J2_125_3477_n2909), 
        .A2(DP_OP_425J2_127_3477_n1953), .Y(DP_OP_425J2_127_3477_n1941) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1236 ( .A1(DP_OP_422J2_124_3477_n2032), 
        .A2(DP_OP_423J2_125_3477_n2034), .Y(DP_OP_422J2_124_3477_n2008) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1422 ( .A1(DP_OP_424J2_126_3477_n2211), 
        .A2(DP_OP_424J2_126_3477_n2216), .Y(DP_OP_424J2_126_3477_n2195) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1289 ( .A1(DP_OP_424J2_126_3477_n2078), 
        .A2(DP_OP_424J2_126_3477_n2084), .Y(DP_OP_424J2_126_3477_n2062) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1300 ( .A1(DP_OP_422J2_124_3477_n2782), 
        .A2(DP_OP_424J2_126_3477_n2085), .Y(DP_OP_424J2_126_3477_n2073) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1631 ( .A1(DP_OP_422J2_124_3477_n2427), 
        .A2(DP_OP_422J2_124_3477_n2434), .Y(DP_OP_422J2_124_3477_n2403) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1916 ( .A1(DP_OP_423J2_125_3477_n2777), 
        .A2(DP_OP_424J2_126_3477_n2698), .Y(DP_OP_424J2_126_3477_n2686) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1256 ( .A1(DP_OP_422J2_124_3477_n1905), 
        .A2(DP_OP_425J2_127_3477_n2041), .Y(DP_OP_425J2_127_3477_n2029) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1597 ( .A1(DP_OP_424J2_126_3477_n2383), 
        .A2(DP_OP_424J2_126_3477_n2389), .Y(DP_OP_424J2_126_3477_n2367) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1325 ( .A1(DP_OP_422J2_124_3477_n2121), 
        .A2(DP_OP_425J2_127_3477_n2127), .Y(DP_OP_422J2_124_3477_n2097) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1156 ( .A1(DP_OP_422J2_124_3477_n1945), 
        .A2(DP_OP_422J2_124_3477_n1952), .Y(DP_OP_422J2_124_3477_n1929) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1943 ( .A1(DP_OP_423J2_125_3477_n2031), 
        .A2(DP_OP_422J2_124_3477_n2740), .Y(DP_OP_422J2_124_3477_n2713) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1772 ( .A1(DP_OP_422J2_124_3477_n2560), 
        .A2(DP_OP_422J2_124_3477_n2567), .Y(DP_OP_422J2_124_3477_n2544) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1774 ( .A1(DP_OP_422J2_124_3477_n2562), 
        .A2(DP_OP_422J2_124_3477_n2567), .Y(DP_OP_422J2_124_3477_n2546) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2081 ( .A1(DP_OP_423J2_125_3477_n1897), 
        .A2(DP_OP_422J2_124_3477_n2873), .Y(DP_OP_422J2_124_3477_n2851) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1013 ( .A1(n270), .A2(n343), .Y(
        DP_OP_425J2_127_3477_n1786) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2082 ( .A1(DP_OP_422J2_124_3477_n2868), 
        .A2(DP_OP_422J2_124_3477_n2873), .Y(DP_OP_422J2_124_3477_n2852) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1687 ( .A1(DP_OP_423J2_125_3477_n2163), 
        .A2(DP_OP_425J2_127_3477_n2477), .Y(DP_OP_425J2_127_3477_n2457) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1941 ( .A1(DP_OP_422J2_124_3477_n2735), 
        .A2(DP_OP_422J2_124_3477_n2740), .Y(DP_OP_422J2_124_3477_n2711) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1149 ( .A1(DP_OP_425J2_127_3477_n2078), 
        .A2(DP_OP_422J2_124_3477_n1951), .Y(DP_OP_422J2_124_3477_n1922) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1455 ( .A1(DP_OP_424J2_126_3477_n2381), 
        .A2(DP_OP_422J2_124_3477_n2258), .Y(DP_OP_422J2_124_3477_n2227) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U989 ( .A1(n318), .A2(n342), .Y(
        DP_OP_425J2_127_3477_n161) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1905 ( .A1(DP_OP_423J2_125_3477_n2073), 
        .A2(DP_OP_422J2_124_3477_n2699), .Y(DP_OP_422J2_124_3477_n2677) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1992 ( .A1(DP_OP_424J2_126_3477_n2077), 
        .A2(DP_OP_422J2_124_3477_n2785), .Y(DP_OP_422J2_124_3477_n2762) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1776 ( .A1(DP_OP_423J2_125_3477_n2076), 
        .A2(DP_OP_425J2_127_3477_n2565), .Y(DP_OP_425J2_127_3477_n2546) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1158 ( .A1(DP_OP_425J2_127_3477_n2079), 
        .A2(DP_OP_422J2_124_3477_n1952), .Y(DP_OP_422J2_124_3477_n1931) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1680 ( .A1(DP_OP_422J2_124_3477_n2476), 
        .A2(DP_OP_422J2_124_3477_n2478), .Y(DP_OP_422J2_124_3477_n2452) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1994 ( .A1(DP_OP_422J2_124_3477_n2780), 
        .A2(DP_OP_422J2_124_3477_n2785), .Y(DP_OP_422J2_124_3477_n2764) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2087 ( .A1(DP_OP_422J2_124_3477_n2865), 
        .A2(DP_OP_424J2_126_3477_n2874), .Y(DP_OP_422J2_124_3477_n2857) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2002 ( .A1(DP_OP_422J2_124_3477_n2780), 
        .A2(DP_OP_422J2_124_3477_n2786), .Y(DP_OP_422J2_124_3477_n2772) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1152 ( .A1(DP_OP_422J2_124_3477_n1949), 
        .A2(DP_OP_422J2_124_3477_n1951), .Y(DP_OP_422J2_124_3477_n1925) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1993 ( .A1(DP_OP_423J2_125_3477_n1985), 
        .A2(DP_OP_422J2_124_3477_n2785), .Y(DP_OP_422J2_124_3477_n2763) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1592 ( .A1(DP_OP_422J2_124_3477_n2388), 
        .A2(DP_OP_422J2_124_3477_n2390), .Y(DP_OP_422J2_124_3477_n2364) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1328 ( .A1(DP_OP_422J2_124_3477_n2124), 
        .A2(DP_OP_423J2_125_3477_n2122), .Y(DP_OP_422J2_124_3477_n2100) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1008 ( .A1(n373), .A2(n342), .Y(
        DP_OP_422J2_124_3477_n1781) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1323 ( .A1(DP_OP_423J2_125_3477_n2599), 
        .A2(DP_OP_424J2_126_3477_n2127), .Y(DP_OP_422J2_124_3477_n2095) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1906 ( .A1(DP_OP_425J2_127_3477_n2692), 
        .A2(DP_OP_424J2_126_3477_n2697), .Y(DP_OP_425J2_127_3477_n2676) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1124 ( .A1(DP_OP_425J2_127_3477_n1905), 
        .A2(DP_OP_423J2_125_3477_n1904), .Y(DP_OP_425J2_127_3477_n1897) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1942 ( .A1(DP_OP_422J2_124_3477_n2736), 
        .A2(DP_OP_422J2_124_3477_n2740), .Y(DP_OP_422J2_124_3477_n2712) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1416 ( .A1(DP_OP_423J2_125_3477_n2516), 
        .A2(DP_OP_422J2_124_3477_n2214), .Y(DP_OP_422J2_124_3477_n2188) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1158 ( .A1(DP_OP_423J2_125_3477_n2907), 
        .A2(DP_OP_424J2_126_3477_n1952), .Y(DP_OP_425J2_127_3477_n1931) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1675 ( .A1(DP_OP_423J2_125_3477_n2291), 
        .A2(DP_OP_422J2_124_3477_n2478), .Y(DP_OP_422J2_124_3477_n2447) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2004 ( .A1(DP_OP_423J2_125_3477_n1856), 
        .A2(DP_OP_425J2_127_3477_n2786), .Y(DP_OP_425J2_127_3477_n2774) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1907 ( .A1(DP_OP_422J2_124_3477_n2695), 
        .A2(DP_OP_422J2_124_3477_n2699), .Y(DP_OP_422J2_124_3477_n2679) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1906 ( .A1(DP_OP_422J2_124_3477_n2694), 
        .A2(DP_OP_422J2_124_3477_n2699), .Y(DP_OP_422J2_124_3477_n2678) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1015 ( .A1(n280), .A2(n338), .Y(
        DP_OP_425J2_127_3477_n1788) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1995 ( .A1(DP_OP_424J2_126_3477_n1948), 
        .A2(DP_OP_425J2_127_3477_n2785), .Y(DP_OP_425J2_127_3477_n2765) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1994 ( .A1(DP_OP_425J2_127_3477_n2780), 
        .A2(DP_OP_425J2_127_3477_n2785), .Y(DP_OP_425J2_127_3477_n2764) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1676 ( .A1(DP_OP_422J2_124_3477_n2472), 
        .A2(DP_OP_422J2_124_3477_n2478), .Y(DP_OP_422J2_124_3477_n2448) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U985 ( .A1(n409), .A2(n339), .Y(
        DP_OP_422J2_124_3477_n153) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1773 ( .A1(DP_OP_423J2_125_3477_n2205), 
        .A2(DP_OP_422J2_124_3477_n2567), .Y(DP_OP_422J2_124_3477_n2545) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1411 ( .A1(DP_OP_422J2_124_3477_n2207), 
        .A2(DP_OP_422J2_124_3477_n2214), .Y(DP_OP_422J2_124_3477_n2183) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1738 ( .A1(DP_OP_422J2_124_3477_n2518), 
        .A2(DP_OP_422J2_124_3477_n2524), .Y(DP_OP_422J2_124_3477_n2510) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2083 ( .A1(DP_OP_425J2_127_3477_n2869), 
        .A2(DP_OP_422J2_124_3477_n2873), .Y(DP_OP_425J2_127_3477_n2853) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2082 ( .A1(DP_OP_425J2_127_3477_n2868), 
        .A2(DP_OP_423J2_125_3477_n2868), .Y(DP_OP_425J2_127_3477_n2852) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1460 ( .A1(DP_OP_424J2_126_3477_n2386), 
        .A2(DP_OP_422J2_124_3477_n2258), .Y(DP_OP_422J2_124_3477_n2232) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1591 ( .A1(DP_OP_423J2_125_3477_n2251), 
        .A2(DP_OP_423J2_125_3477_n2386), .Y(DP_OP_425J2_127_3477_n2361) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1685 ( .A1(DP_OP_422J2_124_3477_n2473), 
        .A2(DP_OP_422J2_124_3477_n2479), .Y(DP_OP_422J2_124_3477_n2457) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1686 ( .A1(DP_OP_423J2_125_3477_n2294), 
        .A2(DP_OP_422J2_124_3477_n2479), .Y(DP_OP_422J2_124_3477_n2458) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1943 ( .A1(DP_OP_423J2_125_3477_n1899), 
        .A2(DP_OP_425J2_127_3477_n2740), .Y(DP_OP_425J2_127_3477_n2713) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2092 ( .A1(DP_OP_425J2_127_3477_n2870), 
        .A2(DP_OP_425J2_127_3477_n2874), .Y(DP_OP_425J2_127_3477_n2862) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1739 ( .A1(DP_OP_424J2_126_3477_n2212), 
        .A2(DP_OP_422J2_124_3477_n2524), .Y(DP_OP_425J2_127_3477_n2509) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1328 ( .A1(DP_OP_423J2_125_3477_n2733), 
        .A2(DP_OP_425J2_127_3477_n2127), .Y(DP_OP_425J2_127_3477_n2101) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1589 ( .A1(DP_OP_422J2_124_3477_n2385), 
        .A2(DP_OP_422J2_124_3477_n2390), .Y(DP_OP_422J2_124_3477_n2361) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1939 ( .A1(DP_OP_422J2_124_3477_n2733), 
        .A2(DP_OP_422J2_124_3477_n2740), .Y(DP_OP_422J2_124_3477_n2709) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2080 ( .A1(DP_OP_423J2_125_3477_n1896), 
        .A2(DP_OP_422J2_124_3477_n2873), .Y(DP_OP_422J2_124_3477_n2850) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1006 ( .A1(n400), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_422J2_124_3477_n1779) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1904 ( .A1(DP_OP_422J2_124_3477_n2692), 
        .A2(DP_OP_422J2_124_3477_n2699), .Y(DP_OP_422J2_124_3477_n2676) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1684 ( .A1(DP_OP_422J2_124_3477_n2472), 
        .A2(DP_OP_422J2_124_3477_n2479), .Y(DP_OP_422J2_124_3477_n2456) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1120 ( .A1(DP_OP_424J2_126_3477_n2734), 
        .A2(DP_OP_422J2_124_3477_n1909), .Y(DP_OP_422J2_124_3477_n1893) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1735 ( .A1(DP_OP_423J2_125_3477_n2247), 
        .A2(DP_OP_422J2_124_3477_n2524), .Y(DP_OP_422J2_124_3477_n2507) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1940 ( .A1(DP_OP_422J2_124_3477_n2734), 
        .A2(DP_OP_422J2_124_3477_n2740), .Y(DP_OP_422J2_124_3477_n2710) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1991 ( .A1(DP_OP_422J2_124_3477_n2777), 
        .A2(DP_OP_422J2_124_3477_n2785), .Y(DP_OP_422J2_124_3477_n2761) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1459 ( .A1(DP_OP_424J2_126_3477_n2385), 
        .A2(DP_OP_422J2_124_3477_n2258), .Y(DP_OP_422J2_124_3477_n2231) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1908 ( .A1(DP_OP_422J2_124_3477_n2696), 
        .A2(DP_OP_422J2_124_3477_n2699), .Y(DP_OP_422J2_124_3477_n2680) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2000 ( .A1(DP_OP_424J2_126_3477_n2077), 
        .A2(DP_OP_422J2_124_3477_n2786), .Y(DP_OP_422J2_124_3477_n2770) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2084 ( .A1(DP_OP_422J2_124_3477_n2870), 
        .A2(DP_OP_422J2_124_3477_n2873), .Y(DP_OP_422J2_124_3477_n2854) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2003 ( .A1(DP_OP_422J2_124_3477_n2781), 
        .A2(DP_OP_422J2_124_3477_n2786), .Y(DP_OP_422J2_124_3477_n2773) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1775 ( .A1(DP_OP_422J2_124_3477_n2563), 
        .A2(DP_OP_422J2_124_3477_n2567), .Y(DP_OP_422J2_124_3477_n2547) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2088 ( .A1(DP_OP_425J2_127_3477_n2734), 
        .A2(DP_OP_425J2_127_3477_n2874), .Y(DP_OP_422J2_124_3477_n2858) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2091 ( .A1(DP_OP_422J2_124_3477_n2869), 
        .A2(DP_OP_425J2_127_3477_n2874), .Y(DP_OP_422J2_124_3477_n2861) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1326 ( .A1(DP_OP_423J2_125_3477_n2602), 
        .A2(DP_OP_423J2_125_3477_n2122), .Y(DP_OP_422J2_124_3477_n2098) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1123 ( .A1(DP_OP_422J2_124_3477_n1904), 
        .A2(DP_OP_422J2_124_3477_n1909), .Y(DP_OP_422J2_124_3477_n1896) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1588 ( .A1(DP_OP_422J2_124_3477_n2384), 
        .A2(DP_OP_422J2_124_3477_n2390), .Y(DP_OP_422J2_124_3477_n2360) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1414 ( .A1(DP_OP_422J2_124_3477_n2210), 
        .A2(DP_OP_422J2_124_3477_n2214), .Y(DP_OP_422J2_124_3477_n2186) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1740 ( .A1(DP_OP_422J2_124_3477_n2520), 
        .A2(DP_OP_422J2_124_3477_n2524), .Y(DP_OP_422J2_124_3477_n2512) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1736 ( .A1(DP_OP_425J2_127_3477_n2382), 
        .A2(DP_OP_422J2_124_3477_n2524), .Y(DP_OP_422J2_124_3477_n2508) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1904 ( .A1(DP_OP_425J2_127_3477_n2690), 
        .A2(DP_OP_422J2_124_3477_n2699), .Y(DP_OP_425J2_127_3477_n2674) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1156 ( .A1(DP_OP_425J2_127_3477_n1945), 
        .A2(DP_OP_424J2_126_3477_n1952), .Y(DP_OP_425J2_127_3477_n1929) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1589 ( .A1(DP_OP_425J2_127_3477_n2383), 
        .A2(DP_OP_423J2_125_3477_n2386), .Y(DP_OP_425J2_127_3477_n2359) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1458 ( .A1(DP_OP_424J2_126_3477_n2384), 
        .A2(DP_OP_422J2_124_3477_n2258), .Y(DP_OP_422J2_124_3477_n2230) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1678 ( .A1(DP_OP_423J2_125_3477_n2294), 
        .A2(DP_OP_422J2_124_3477_n2478), .Y(DP_OP_422J2_124_3477_n2450) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1739 ( .A1(DP_OP_424J2_126_3477_n2344), 
        .A2(DP_OP_422J2_124_3477_n2524), .Y(DP_OP_422J2_124_3477_n2511) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1587 ( .A1(DP_OP_422J2_124_3477_n2383), 
        .A2(DP_OP_422J2_124_3477_n2390), .Y(DP_OP_422J2_124_3477_n2359) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2004 ( .A1(DP_OP_422J2_124_3477_n2782), 
        .A2(DP_OP_422J2_124_3477_n2786), .Y(DP_OP_422J2_124_3477_n2774) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1014 ( .A1(n285), .A2(n343), .Y(
        DP_OP_422J2_124_3477_n1787) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1456 ( .A1(DP_OP_424J2_126_3477_n2382), 
        .A2(DP_OP_422J2_124_3477_n2258), .Y(DP_OP_422J2_124_3477_n2228) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1677 ( .A1(DP_OP_422J2_124_3477_n2473), 
        .A2(DP_OP_422J2_124_3477_n2478), .Y(DP_OP_422J2_124_3477_n2449) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1324 ( .A1(DP_OP_422J2_124_3477_n2120), 
        .A2(DP_OP_425J2_127_3477_n2127), .Y(DP_OP_422J2_124_3477_n2096) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1996 ( .A1(DP_OP_422J2_124_3477_n2782), 
        .A2(DP_OP_422J2_124_3477_n2785), .Y(DP_OP_422J2_124_3477_n2766) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1412 ( .A1(DP_OP_422J2_124_3477_n2208), 
        .A2(DP_OP_422J2_124_3477_n2214), .Y(DP_OP_422J2_124_3477_n2184) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1740 ( .A1(DP_OP_425J2_127_3477_n2518), 
        .A2(DP_OP_422J2_124_3477_n2524), .Y(DP_OP_425J2_127_3477_n2510) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1155 ( .A1(DP_OP_423J2_125_3477_n2772), 
        .A2(DP_OP_422J2_124_3477_n1952), .Y(DP_OP_422J2_124_3477_n1928) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1776 ( .A1(DP_OP_422J2_124_3477_n2564), 
        .A2(DP_OP_422J2_124_3477_n2567), .Y(DP_OP_422J2_124_3477_n2548) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1148 ( .A1(DP_OP_422J2_124_3477_n1945), 
        .A2(DP_OP_422J2_124_3477_n1951), .Y(DP_OP_422J2_124_3477_n1921) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1688 ( .A1(DP_OP_422J2_124_3477_n2476), 
        .A2(DP_OP_422J2_124_3477_n2479), .Y(DP_OP_422J2_124_3477_n2460) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1590 ( .A1(DP_OP_425J2_127_3477_n2384), 
        .A2(DP_OP_424J2_126_3477_n2388), .Y(DP_OP_425J2_127_3477_n2360) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1457 ( .A1(DP_OP_424J2_126_3477_n2383), 
        .A2(DP_OP_422J2_124_3477_n2258), .Y(DP_OP_422J2_124_3477_n2229) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1160 ( .A1(DP_OP_422J2_124_3477_n1949), 
        .A2(DP_OP_422J2_124_3477_n1952), .Y(DP_OP_422J2_124_3477_n1933) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1157 ( .A1(DP_OP_423J2_125_3477_n2906), 
        .A2(DP_OP_422J2_124_3477_n1952), .Y(DP_OP_425J2_127_3477_n1930) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1905 ( .A1(DP_OP_425J2_127_3477_n2691), 
        .A2(DP_OP_422J2_124_3477_n2699), .Y(DP_OP_425J2_127_3477_n2675) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1124 ( .A1(DP_OP_422J2_124_3477_n1905), 
        .A2(DP_OP_422J2_124_3477_n1909), .Y(DP_OP_422J2_124_3477_n1897) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1683 ( .A1(DP_OP_423J2_125_3477_n2291), 
        .A2(DP_OP_422J2_124_3477_n2479), .Y(DP_OP_422J2_124_3477_n2455) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1590 ( .A1(DP_OP_422J2_124_3477_n2386), 
        .A2(DP_OP_422J2_124_3477_n2390), .Y(DP_OP_422J2_124_3477_n2362) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1157 ( .A1(DP_OP_425J2_127_3477_n2078), 
        .A2(DP_OP_422J2_124_3477_n1952), .Y(DP_OP_422J2_124_3477_n1930) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1147 ( .A1(DP_OP_423J2_125_3477_n2772), 
        .A2(DP_OP_422J2_124_3477_n1951), .Y(DP_OP_422J2_124_3477_n1920) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1150 ( .A1(DP_OP_425J2_127_3477_n2079), 
        .A2(DP_OP_422J2_124_3477_n1951), .Y(DP_OP_422J2_124_3477_n1923) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1327 ( .A1(DP_OP_424J2_126_3477_n2517), 
        .A2(DP_OP_424J2_126_3477_n2127), .Y(DP_OP_422J2_124_3477_n2099) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1995 ( .A1(DP_OP_422J2_124_3477_n2781), 
        .A2(DP_OP_422J2_124_3477_n2785), .Y(DP_OP_422J2_124_3477_n2765) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1416 ( .A1(DP_OP_425J2_127_3477_n2213), 
        .A2(DP_OP_425J2_127_3477_n2215), .Y(DP_OP_425J2_127_3477_n2189) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1738 ( .A1(DP_OP_422J2_124_3477_n2650), 
        .A2(DP_OP_423J2_125_3477_n2520), .Y(DP_OP_425J2_127_3477_n2508) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U992 ( .A1(n382), .A2(n339), .Y(
        DP_OP_422J2_124_3477_n167) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2090 ( .A1(DP_OP_425J2_127_3477_n2868), 
        .A2(DP_OP_425J2_127_3477_n2874), .Y(DP_OP_425J2_127_3477_n2860) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U991 ( .A1(n418), .A2(n340), .Y(
        DP_OP_422J2_124_3477_n165) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1944 ( .A1(DP_OP_423J2_125_3477_n2032), 
        .A2(DP_OP_422J2_124_3477_n2740), .Y(DP_OP_422J2_124_3477_n2714) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1996 ( .A1(DP_OP_424J2_126_3477_n1949), 
        .A2(DP_OP_425J2_127_3477_n2785), .Y(DP_OP_425J2_127_3477_n2766) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1908 ( .A1(DP_OP_425J2_127_3477_n2694), 
        .A2(DP_OP_423J2_125_3477_n2695), .Y(DP_OP_425J2_127_3477_n2678) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1774 ( .A1(DP_OP_422J2_124_3477_n2694), 
        .A2(DP_OP_425J2_127_3477_n2565), .Y(DP_OP_425J2_127_3477_n2544) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1999 ( .A1(DP_OP_422J2_124_3477_n2777), 
        .A2(DP_OP_422J2_124_3477_n2786), .Y(DP_OP_422J2_124_3477_n2769) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1687 ( .A1(DP_OP_423J2_125_3477_n2295), 
        .A2(DP_OP_422J2_124_3477_n2479), .Y(DP_OP_422J2_124_3477_n2459) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1160 ( .A1(DP_OP_423J2_125_3477_n2909), 
        .A2(DP_OP_422J2_124_3477_n1952), .Y(DP_OP_425J2_127_3477_n1933) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1121 ( .A1(DP_OP_422J2_124_3477_n1902), 
        .A2(DP_OP_422J2_124_3477_n1909), .Y(DP_OP_422J2_124_3477_n1894) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U990 ( .A1(n421), .A2(n341), .Y(
        DP_OP_422J2_124_3477_n163) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1152 ( .A1(DP_OP_423J2_125_3477_n2909), 
        .A2(DP_OP_425J2_127_3477_n1951), .Y(DP_OP_425J2_127_3477_n1925) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U989 ( .A1(n410), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_422J2_124_3477_n161) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U988 ( .A1(n376), .A2(n339), .Y(
        DP_OP_422J2_124_3477_n159) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1122 ( .A1(DP_OP_425J2_127_3477_n1903), 
        .A2(DP_OP_422J2_124_3477_n1909), .Y(DP_OP_425J2_127_3477_n1895) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2002 ( .A1(DP_OP_425J2_127_3477_n2780), 
        .A2(DP_OP_425J2_127_3477_n2786), .Y(DP_OP_425J2_127_3477_n2772) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1737 ( .A1(DP_OP_423J2_125_3477_n2117), 
        .A2(DP_OP_424J2_126_3477_n2522), .Y(DP_OP_425J2_127_3477_n2507) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U987 ( .A1(n405), .A2(n343), .Y(
        DP_OP_422J2_124_3477_n157) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U986 ( .A1(n420), .A2(n342), .Y(
        DP_OP_422J2_124_3477_n155) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1775 ( .A1(DP_OP_424J2_126_3477_n2168), 
        .A2(DP_OP_425J2_127_3477_n2565), .Y(DP_OP_425J2_127_3477_n2545) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1686 ( .A1(DP_OP_425J2_127_3477_n2472), 
        .A2(DP_OP_425J2_127_3477_n2477), .Y(DP_OP_425J2_127_3477_n2456) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2001 ( .A1(DP_OP_425J2_127_3477_n2779), 
        .A2(DP_OP_425J2_127_3477_n2786), .Y(DP_OP_425J2_127_3477_n2771) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1679 ( .A1(DP_OP_423J2_125_3477_n2163), 
        .A2(DP_OP_425J2_127_3477_n2476), .Y(DP_OP_425J2_127_3477_n2449) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1591 ( .A1(DP_OP_422J2_124_3477_n2387), 
        .A2(DP_OP_422J2_124_3477_n2390), .Y(DP_OP_422J2_124_3477_n2363) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1415 ( .A1(DP_OP_423J2_125_3477_n2647), 
        .A2(DP_OP_425J2_127_3477_n2215), .Y(DP_OP_425J2_127_3477_n2188) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2090 ( .A1(DP_OP_422J2_124_3477_n2868), 
        .A2(DP_OP_425J2_127_3477_n2874), .Y(DP_OP_422J2_124_3477_n2860) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1680 ( .A1(DP_OP_423J2_125_3477_n2164), 
        .A2(DP_OP_425J2_127_3477_n2476), .Y(DP_OP_425J2_127_3477_n2450) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1003 ( .A1(n403), .A2(n339), .Y(
        DP_OP_422J2_124_3477_n1776) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1460 ( .A1(DP_OP_423J2_125_3477_n2604), 
        .A2(DP_OP_425J2_127_3477_n2259), .Y(DP_OP_425J2_127_3477_n2233) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1151 ( .A1(DP_OP_423J2_125_3477_n2776), 
        .A2(DP_OP_422J2_124_3477_n1951), .Y(DP_OP_422J2_124_3477_n1924) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1944 ( .A1(DP_OP_425J2_127_3477_n2738), 
        .A2(DP_OP_425J2_127_3477_n2740), .Y(DP_OP_425J2_127_3477_n2714) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1159 ( .A1(DP_OP_423J2_125_3477_n2908), 
        .A2(DP_OP_423J2_125_3477_n1947), .Y(DP_OP_425J2_127_3477_n1932) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1903 ( .A1(DP_OP_425J2_127_3477_n2557), 
        .A2(DP_OP_422J2_124_3477_n2699), .Y(DP_OP_422J2_124_3477_n2675) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2079 ( .A1(DP_OP_422J2_124_3477_n2865), 
        .A2(DP_OP_422J2_124_3477_n2873), .Y(DP_OP_422J2_124_3477_n2849) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1413 ( .A1(DP_OP_422J2_124_3477_n2209), 
        .A2(DP_OP_422J2_124_3477_n2214), .Y(DP_OP_422J2_124_3477_n2185) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1907 ( .A1(DP_OP_423J2_125_3477_n1943), 
        .A2(DP_OP_424J2_126_3477_n2697), .Y(DP_OP_425J2_127_3477_n2677) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2089 ( .A1(DP_OP_423J2_125_3477_n1897), 
        .A2(DP_OP_424J2_126_3477_n2874), .Y(DP_OP_422J2_124_3477_n2859) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1123 ( .A1(DP_OP_424J2_126_3477_n2869), 
        .A2(DP_OP_424J2_126_3477_n1909), .Y(DP_OP_425J2_127_3477_n1896) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1159 ( .A1(DP_OP_424J2_126_3477_n2693), 
        .A2(DP_OP_422J2_124_3477_n1952), .Y(DP_OP_422J2_124_3477_n1932) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2091 ( .A1(DP_OP_425J2_127_3477_n2869), 
        .A2(DP_OP_425J2_127_3477_n2874), .Y(DP_OP_425J2_127_3477_n2861) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2092 ( .A1(DP_OP_422J2_124_3477_n2870), 
        .A2(DP_OP_424J2_126_3477_n2874), .Y(DP_OP_422J2_124_3477_n2862) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2003 ( .A1(DP_OP_422J2_124_3477_n2913), 
        .A2(DP_OP_425J2_127_3477_n2786), .Y(DP_OP_425J2_127_3477_n2773) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1688 ( .A1(DP_OP_423J2_125_3477_n2164), 
        .A2(DP_OP_425J2_127_3477_n2477), .Y(DP_OP_425J2_127_3477_n2458) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1679 ( .A1(DP_OP_423J2_125_3477_n2295), 
        .A2(DP_OP_422J2_124_3477_n2478), .Y(DP_OP_422J2_124_3477_n2451) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1771 ( .A1(DP_OP_422J2_124_3477_n2559), 
        .A2(DP_OP_422J2_124_3477_n2567), .Y(DP_OP_422J2_124_3477_n2543) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1327 ( .A1(DP_OP_423J2_125_3477_n2732), 
        .A2(DP_OP_425J2_127_3477_n2127), .Y(DP_OP_425J2_127_3477_n2100) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1121 ( .A1(DP_OP_424J2_126_3477_n2867), 
        .A2(DP_OP_423J2_125_3477_n1904), .Y(DP_OP_425J2_127_3477_n1894) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1737 ( .A1(DP_OP_424J2_126_3477_n2342), 
        .A2(DP_OP_422J2_124_3477_n2524), .Y(DP_OP_422J2_124_3477_n2509) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1459 ( .A1(DP_OP_424J2_126_3477_n2517), 
        .A2(DP_OP_425J2_127_3477_n2259), .Y(DP_OP_425J2_127_3477_n2232) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2089 ( .A1(DP_OP_424J2_126_3477_n1858), 
        .A2(DP_OP_425J2_127_3477_n2874), .Y(DP_OP_425J2_127_3477_n2859) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1592 ( .A1(DP_OP_425J2_127_3477_n2386), 
        .A2(DP_OP_424J2_126_3477_n2388), .Y(DP_OP_425J2_127_3477_n2362) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1151 ( .A1(DP_OP_423J2_125_3477_n2908), 
        .A2(DP_OP_425J2_127_3477_n1951), .Y(DP_OP_425J2_127_3477_n1924) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2083 ( .A1(DP_OP_422J2_124_3477_n2869), 
        .A2(DP_OP_422J2_124_3477_n2873), .Y(DP_OP_422J2_124_3477_n2853) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2084 ( .A1(DP_OP_425J2_127_3477_n2870), 
        .A2(DP_OP_422J2_124_3477_n2873), .Y(DP_OP_425J2_127_3477_n2854) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1415 ( .A1(DP_OP_422J2_124_3477_n2211), 
        .A2(DP_OP_422J2_124_3477_n2214), .Y(DP_OP_422J2_124_3477_n2187) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1122 ( .A1(DP_OP_422J2_124_3477_n1903), 
        .A2(DP_OP_422J2_124_3477_n1909), .Y(DP_OP_422J2_124_3477_n1895) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1012 ( .A1(n369), .A2(n341), .Y(
        DP_OP_422J2_124_3477_n1785) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2001 ( .A1(DP_OP_424J2_126_3477_n2078), 
        .A2(DP_OP_422J2_124_3477_n2786), .Y(DP_OP_422J2_124_3477_n2771) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1933 ( .A1(DP_OP_425J2_127_3477_n2120), 
        .A2(DP_OP_425J2_127_3477_n2740), .Y(DP_OP_423J2_125_3477_n2704) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1141 ( .A1(DP_OP_423J2_125_3477_n1939), 
        .A2(n442), .Y(DP_OP_423J2_125_3477_n1915) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1004 ( .A1(n269), .A2(n339), .Y(
        DP_OP_423J2_125_3477_n1778) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1993 ( .A1(DP_OP_423J2_125_3477_n2772), 
        .A2(DP_OP_423J2_125_3477_n2781), .Y(DP_OP_423J2_125_3477_n2764) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1451 ( .A1(DP_OP_424J2_126_3477_n2342), 
        .A2(DP_OP_423J2_125_3477_n2254), .Y(DP_OP_423J2_125_3477_n2225) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1319 ( .A1(DP_OP_423J2_125_3477_n2117), 
        .A2(DP_OP_423J2_125_3477_n2122), .Y(DP_OP_423J2_125_3477_n2093) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1671 ( .A1(DP_OP_423J2_125_3477_n2469), 
        .A2(DP_OP_423J2_125_3477_n2474), .Y(DP_OP_423J2_125_3477_n2445) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1729 ( .A1(DP_OP_425J2_127_3477_n2340), 
        .A2(DP_OP_423J2_125_3477_n2520), .Y(DP_OP_423J2_125_3477_n2503) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2081 ( .A1(DP_OP_423J2_125_3477_n2860), 
        .A2(DP_OP_423J2_125_3477_n2869), .Y(DP_OP_423J2_125_3477_n2852) );
  XNOR2X1_HVT DP_OP_424J2_126_3477_U627 ( .A1(DP_OP_424J2_126_3477_n2002), 
        .A2(DP_OP_424J2_126_3477_n2352), .Y(DP_OP_424J2_126_3477_n1062) );
  OR2X1_HVT DP_OP_425J2_127_3477_U984 ( .A1(n381), .A2(n339), .Y(
        DP_OP_425J2_127_3477_n1773) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1113 ( .A1(DP_OP_424J2_126_3477_n1988), 
        .A2(DP_OP_423J2_125_3477_n1904), .Y(DP_OP_423J2_125_3477_n1887) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1006 ( .A1(n291), .A2(n343), .Y(
        DP_OP_425J2_127_3477_n1779) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1323 ( .A1(DP_OP_424J2_126_3477_n2120), 
        .A2(DP_OP_424J2_126_3477_n2127), .Y(DP_OP_424J2_126_3477_n2096) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1675 ( .A1(DP_OP_425J2_127_3477_n2296), 
        .A2(DP_OP_425J2_127_3477_n2476), .Y(DP_OP_424J2_126_3477_n2445) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1455 ( .A1(DP_OP_422J2_124_3477_n2603), 
        .A2(DP_OP_423J2_125_3477_n2254), .Y(DP_OP_424J2_126_3477_n2228) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1771 ( .A1(DP_OP_424J2_126_3477_n2557), 
        .A2(DP_OP_424J2_126_3477_n2565), .Y(DP_OP_424J2_126_3477_n2541) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1683 ( .A1(DP_OP_425J2_127_3477_n2296), 
        .A2(DP_OP_422J2_124_3477_n2479), .Y(DP_OP_424J2_126_3477_n2453) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1148 ( .A1(DP_OP_425J2_127_3477_n2778), 
        .A2(n442), .Y(DP_OP_424J2_126_3477_n1921) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1412 ( .A1(DP_OP_423J2_125_3477_n2116), 
        .A2(n443), .Y(DP_OP_424J2_126_3477_n2185) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1940 ( .A1(DP_OP_424J2_126_3477_n2734), 
        .A2(DP_OP_424J2_126_3477_n2740), .Y(DP_OP_424J2_126_3477_n2710) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1991 ( .A1(DP_OP_424J2_126_3477_n2777), 
        .A2(DP_OP_424J2_126_3477_n2785), .Y(DP_OP_424J2_126_3477_n2761) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1903 ( .A1(DP_OP_424J2_126_3477_n2689), 
        .A2(DP_OP_424J2_126_3477_n2697), .Y(DP_OP_424J2_126_3477_n2673) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1155 ( .A1(DP_OP_425J2_127_3477_n2777), 
        .A2(DP_OP_424J2_126_3477_n1952), .Y(DP_OP_424J2_126_3477_n1928) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1002 ( .A1(n264), .A2(n339), .Y(
        DP_OP_423J2_125_3477_n1776) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1588 ( .A1(DP_OP_424J2_126_3477_n2382), 
        .A2(DP_OP_424J2_126_3477_n2388), .Y(DP_OP_424J2_126_3477_n2358) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1317 ( .A1(DP_OP_423J2_125_3477_n2115), 
        .A2(DP_OP_423J2_125_3477_n2122), .Y(DP_OP_423J2_125_3477_n2091) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1449 ( .A1(DP_OP_423J2_125_3477_n2247), 
        .A2(DP_OP_423J2_125_3477_n2254), .Y(DP_OP_423J2_125_3477_n2223) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1669 ( .A1(DP_OP_423J2_125_3477_n2467), 
        .A2(DP_OP_423J2_125_3477_n2474), .Y(DP_OP_423J2_125_3477_n2443) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1581 ( .A1(DP_OP_422J2_124_3477_n2339), 
        .A2(DP_OP_423J2_125_3477_n2386), .Y(DP_OP_423J2_125_3477_n2355) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U992 ( .A1(n383), .A2(n339), .Y(
        DP_OP_424J2_126_3477_n167) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U991 ( .A1(n408), .A2(n343), .Y(
        DP_OP_424J2_126_3477_n165) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U990 ( .A1(n425), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_424J2_126_3477_n163) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U989 ( .A1(n396), .A2(n340), .Y(
        DP_OP_424J2_126_3477_n161) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2079 ( .A1(DP_OP_424J2_126_3477_n2865), 
        .A2(DP_OP_424J2_126_3477_n2873), .Y(DP_OP_424J2_126_3477_n2849) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1405 ( .A1(DP_OP_422J2_124_3477_n2559), 
        .A2(n443), .Y(DP_OP_423J2_125_3477_n2179) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1404 ( .A1(DP_OP_425J2_127_3477_n2424), 
        .A2(DP_OP_425J2_127_3477_n2215), .Y(DP_OP_423J2_125_3477_n2178) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1005 ( .A1(n284), .A2(n340), .Y(
        DP_OP_425J2_127_3477_n1778) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1003 ( .A1(n287), .A2(n342), .Y(
        DP_OP_425J2_127_3477_n1776) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1325 ( .A1(DP_OP_423J2_125_3477_n2029), 
        .A2(DP_OP_424J2_126_3477_n2127), .Y(DP_OP_424J2_126_3477_n2098) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2087 ( .A1(DP_OP_424J2_126_3477_n2865), 
        .A2(DP_OP_424J2_126_3477_n2874), .Y(DP_OP_424J2_126_3477_n2857) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2079 ( .A1(DP_OP_425J2_127_3477_n2865), 
        .A2(DP_OP_422J2_124_3477_n2873), .Y(DP_OP_425J2_127_3477_n2849) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1677 ( .A1(DP_OP_424J2_126_3477_n2471), 
        .A2(DP_OP_423J2_125_3477_n2474), .Y(DP_OP_424J2_126_3477_n2447) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1003 ( .A1(n274), .A2(n339), .Y(
        DP_OP_423J2_125_3477_n1777) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1010 ( .A1(n367), .A2(n341), .Y(
        DP_OP_424J2_126_3477_n1783) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1772 ( .A1(DP_OP_422J2_124_3477_n2076), 
        .A2(DP_OP_424J2_126_3477_n2565), .Y(DP_OP_424J2_126_3477_n2542) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1684 ( .A1(DP_OP_422J2_124_3477_n2164), 
        .A2(DP_OP_422J2_124_3477_n2479), .Y(DP_OP_424J2_126_3477_n2454) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1898 ( .A1(DP_OP_423J2_125_3477_n2688), 
        .A2(DP_OP_423J2_125_3477_n2695), .Y(DP_OP_423J2_125_3477_n2672) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1986 ( .A1(DP_OP_425J2_127_3477_n2077), 
        .A2(DP_OP_422J2_124_3477_n2785), .Y(DP_OP_423J2_125_3477_n2757) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1939 ( .A1(DP_OP_424J2_126_3477_n2733), 
        .A2(DP_OP_424J2_126_3477_n2740), .Y(DP_OP_424J2_126_3477_n2709) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1147 ( .A1(DP_OP_425J2_127_3477_n2777), 
        .A2(DP_OP_422J2_124_3477_n1951), .Y(DP_OP_424J2_126_3477_n1920) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1411 ( .A1(DP_OP_423J2_125_3477_n2115), 
        .A2(n443), .Y(DP_OP_424J2_126_3477_n2184) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1143 ( .A1(DP_OP_425J2_127_3477_n2691), 
        .A2(DP_OP_422J2_124_3477_n1951), .Y(DP_OP_423J2_125_3477_n1917) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1678 ( .A1(DP_OP_423J2_125_3477_n2468), 
        .A2(DP_OP_423J2_125_3477_n2475), .Y(DP_OP_423J2_125_3477_n2452) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2074 ( .A1(DP_OP_423J2_125_3477_n2861), 
        .A2(DP_OP_423J2_125_3477_n2868), .Y(DP_OP_423J2_125_3477_n2845) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1007 ( .A1(n387), .A2(n342), .Y(
        DP_OP_425J2_127_3477_n1780) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1583 ( .A1(DP_OP_422J2_124_3477_n2341), 
        .A2(DP_OP_423J2_125_3477_n2386), .Y(DP_OP_423J2_125_3477_n2357) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1587 ( .A1(DP_OP_424J2_126_3477_n2381), 
        .A2(DP_OP_424J2_126_3477_n2388), .Y(DP_OP_424J2_126_3477_n2357) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1150 ( .A1(DP_OP_425J2_127_3477_n2690), 
        .A2(DP_OP_423J2_125_3477_n1947), .Y(DP_OP_423J2_125_3477_n1924) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1769 ( .A1(DP_OP_423J2_125_3477_n2559), 
        .A2(DP_OP_422J2_124_3477_n2567), .Y(DP_OP_423J2_125_3477_n2543) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1152 ( .A1(DP_OP_424J2_126_3477_n1949), 
        .A2(n442), .Y(DP_OP_424J2_126_3477_n1925) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1416 ( .A1(DP_OP_422J2_124_3477_n2652), 
        .A2(n443), .Y(DP_OP_424J2_126_3477_n2189) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1938 ( .A1(DP_OP_423J2_125_3477_n2733), 
        .A2(DP_OP_422J2_124_3477_n2740), .Y(DP_OP_423J2_125_3477_n2709) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1158 ( .A1(DP_OP_425J2_127_3477_n2780), 
        .A2(DP_OP_424J2_126_3477_n1952), .Y(DP_OP_424J2_126_3477_n1931) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1738 ( .A1(DP_OP_423J2_125_3477_n2602), 
        .A2(DP_OP_424J2_126_3477_n2522), .Y(DP_OP_424J2_126_3477_n2508) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1679 ( .A1(DP_OP_423J2_125_3477_n2469), 
        .A2(DP_OP_423J2_125_3477_n2475), .Y(DP_OP_423J2_125_3477_n2453) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1013 ( .A1(n394), .A2(n341), .Y(
        DP_OP_424J2_126_3477_n1786) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2075 ( .A1(DP_OP_425J2_127_3477_n1990), 
        .A2(DP_OP_423J2_125_3477_n2868), .Y(DP_OP_423J2_125_3477_n2846) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2002 ( .A1(DP_OP_425J2_127_3477_n1991), 
        .A2(DP_OP_422J2_124_3477_n2786), .Y(DP_OP_424J2_126_3477_n2772) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1687 ( .A1(DP_OP_425J2_127_3477_n2300), 
        .A2(DP_OP_425J2_127_3477_n2477), .Y(DP_OP_424J2_126_3477_n2457) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1906 ( .A1(DP_OP_423J2_125_3477_n2775), 
        .A2(DP_OP_424J2_126_3477_n2697), .Y(DP_OP_424J2_126_3477_n2676) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2083 ( .A1(DP_OP_424J2_126_3477_n2869), 
        .A2(DP_OP_424J2_126_3477_n2873), .Y(DP_OP_424J2_126_3477_n2853) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1767 ( .A1(DP_OP_422J2_124_3477_n2165), 
        .A2(DP_OP_425J2_127_3477_n2565), .Y(DP_OP_423J2_125_3477_n2541) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1995 ( .A1(DP_OP_425J2_127_3477_n1992), 
        .A2(DP_OP_424J2_126_3477_n2785), .Y(DP_OP_424J2_126_3477_n2765) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1681 ( .A1(DP_OP_423J2_125_3477_n2471), 
        .A2(DP_OP_423J2_125_3477_n2475), .Y(DP_OP_423J2_125_3477_n2455) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1775 ( .A1(DP_OP_424J2_126_3477_n2561), 
        .A2(DP_OP_424J2_126_3477_n2565), .Y(DP_OP_424J2_126_3477_n2545) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1328 ( .A1(DP_OP_424J2_126_3477_n2125), 
        .A2(DP_OP_424J2_126_3477_n2127), .Y(DP_OP_424J2_126_3477_n2101) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1408 ( .A1(DP_OP_422J2_124_3477_n2562), 
        .A2(DP_OP_425J2_127_3477_n2215), .Y(DP_OP_423J2_125_3477_n2182) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1936 ( .A1(DP_OP_423J2_125_3477_n2731), 
        .A2(DP_OP_422J2_124_3477_n2740), .Y(DP_OP_423J2_125_3477_n2707) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1122 ( .A1(DP_OP_424J2_126_3477_n1903), 
        .A2(DP_OP_424J2_126_3477_n1909), .Y(DP_OP_424J2_126_3477_n1895) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1460 ( .A1(DP_OP_422J2_124_3477_n2608), 
        .A2(DP_OP_422J2_124_3477_n2258), .Y(DP_OP_424J2_126_3477_n2233) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1680 ( .A1(DP_OP_424J2_126_3477_n2474), 
        .A2(DP_OP_425J2_127_3477_n2476), .Y(DP_OP_424J2_126_3477_n2450) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1586 ( .A1(DP_OP_422J2_124_3477_n2344), 
        .A2(DP_OP_423J2_125_3477_n2386), .Y(DP_OP_423J2_125_3477_n2360) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2090 ( .A1(DP_OP_425J2_127_3477_n1903), 
        .A2(DP_OP_424J2_126_3477_n2874), .Y(DP_OP_424J2_126_3477_n2860) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1674 ( .A1(DP_OP_423J2_125_3477_n2472), 
        .A2(DP_OP_423J2_125_3477_n2474), .Y(DP_OP_423J2_125_3477_n2448) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1996 ( .A1(DP_OP_423J2_125_3477_n2775), 
        .A2(DP_OP_423J2_125_3477_n2781), .Y(DP_OP_423J2_125_3477_n2767) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1454 ( .A1(DP_OP_425J2_127_3477_n2386), 
        .A2(DP_OP_423J2_125_3477_n2254), .Y(DP_OP_423J2_125_3477_n2228) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1116 ( .A1(DP_OP_423J2_125_3477_n1898), 
        .A2(DP_OP_423J2_125_3477_n1904), .Y(DP_OP_423J2_125_3477_n1890) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2084 ( .A1(DP_OP_422J2_124_3477_n1859), 
        .A2(DP_OP_423J2_125_3477_n2869), .Y(DP_OP_423J2_125_3477_n2855) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1944 ( .A1(DP_OP_424J2_126_3477_n2738), 
        .A2(DP_OP_424J2_126_3477_n2740), .Y(DP_OP_424J2_126_3477_n2714) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1157 ( .A1(DP_OP_423J2_125_3477_n1853), 
        .A2(DP_OP_424J2_126_3477_n1952), .Y(DP_OP_424J2_126_3477_n1930) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1732 ( .A1(DP_OP_424J2_126_3477_n2428), 
        .A2(DP_OP_423J2_125_3477_n2520), .Y(DP_OP_423J2_125_3477_n2506) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1322 ( .A1(DP_OP_425J2_127_3477_n2518), 
        .A2(DP_OP_423J2_125_3477_n2122), .Y(DP_OP_423J2_125_3477_n2096) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1997 ( .A1(DP_OP_423J2_125_3477_n2776), 
        .A2(DP_OP_423J2_125_3477_n2781), .Y(DP_OP_423J2_125_3477_n2768) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1935 ( .A1(DP_OP_423J2_125_3477_n2730), 
        .A2(DP_OP_425J2_127_3477_n2740), .Y(DP_OP_423J2_125_3477_n2706) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1766 ( .A1(DP_OP_422J2_124_3477_n2164), 
        .A2(DP_OP_422J2_124_3477_n2567), .Y(DP_OP_423J2_125_3477_n2540) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1407 ( .A1(DP_OP_423J2_125_3477_n2205), 
        .A2(DP_OP_425J2_127_3477_n2215), .Y(DP_OP_423J2_125_3477_n2181) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2086 ( .A1(DP_OP_423J2_125_3477_n2865), 
        .A2(DP_OP_423J2_125_3477_n2869), .Y(DP_OP_423J2_125_3477_n2857) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1118 ( .A1(DP_OP_425J2_127_3477_n2738), 
        .A2(DP_OP_423J2_125_3477_n1904), .Y(DP_OP_423J2_125_3477_n1892) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1998 ( .A1(DP_OP_423J2_125_3477_n2777), 
        .A2(DP_OP_423J2_125_3477_n2781), .Y(DP_OP_423J2_125_3477_n2769) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1734 ( .A1(DP_OP_423J2_125_3477_n2516), 
        .A2(DP_OP_423J2_125_3477_n2520), .Y(DP_OP_423J2_125_3477_n2508) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1679 ( .A1(DP_OP_425J2_127_3477_n2300), 
        .A2(DP_OP_425J2_127_3477_n2476), .Y(DP_OP_424J2_126_3477_n2449) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1453 ( .A1(DP_OP_423J2_125_3477_n2251), 
        .A2(DP_OP_423J2_125_3477_n2254), .Y(DP_OP_423J2_125_3477_n2227) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2083 ( .A1(DP_OP_425J2_127_3477_n1990), 
        .A2(DP_OP_423J2_125_3477_n2869), .Y(DP_OP_423J2_125_3477_n2854) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1995 ( .A1(DP_OP_425J2_127_3477_n2078), 
        .A2(DP_OP_423J2_125_3477_n2781), .Y(DP_OP_423J2_125_3477_n2766) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1585 ( .A1(DP_OP_422J2_124_3477_n2343), 
        .A2(DP_OP_423J2_125_3477_n2386), .Y(DP_OP_423J2_125_3477_n2359) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1731 ( .A1(DP_OP_425J2_127_3477_n2342), 
        .A2(DP_OP_423J2_125_3477_n2520), .Y(DP_OP_423J2_125_3477_n2505) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1121 ( .A1(DP_OP_425J2_127_3477_n2823), 
        .A2(DP_OP_424J2_126_3477_n1909), .Y(DP_OP_424J2_126_3477_n1894) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1321 ( .A1(DP_OP_422J2_124_3477_n2651), 
        .A2(DP_OP_423J2_125_3477_n2122), .Y(DP_OP_423J2_125_3477_n2095) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1774 ( .A1(DP_OP_422J2_124_3477_n2078), 
        .A2(DP_OP_424J2_126_3477_n2565), .Y(DP_OP_424J2_126_3477_n2544) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2089 ( .A1(DP_OP_424J2_126_3477_n2867), 
        .A2(DP_OP_424J2_126_3477_n2874), .Y(DP_OP_424J2_126_3477_n2859) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1459 ( .A1(DP_OP_422J2_124_3477_n2607), 
        .A2(DP_OP_423J2_125_3477_n2254), .Y(DP_OP_424J2_126_3477_n2232) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1115 ( .A1(DP_OP_423J2_125_3477_n1897), 
        .A2(DP_OP_423J2_125_3477_n1904), .Y(DP_OP_423J2_125_3477_n1889) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1737 ( .A1(DP_OP_423J2_125_3477_n2601), 
        .A2(DP_OP_424J2_126_3477_n2522), .Y(DP_OP_424J2_126_3477_n2507) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1943 ( .A1(DP_OP_424J2_126_3477_n2737), 
        .A2(DP_OP_424J2_126_3477_n2740), .Y(DP_OP_424J2_126_3477_n2713) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1900 ( .A1(DP_OP_423J2_125_3477_n2690), 
        .A2(DP_OP_423J2_125_3477_n2695), .Y(DP_OP_423J2_125_3477_n2674) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1988 ( .A1(DP_OP_423J2_125_3477_n2775), 
        .A2(DP_OP_422J2_124_3477_n2785), .Y(DP_OP_423J2_125_3477_n2759) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2076 ( .A1(DP_OP_425J2_127_3477_n1991), 
        .A2(DP_OP_423J2_125_3477_n2868), .Y(DP_OP_423J2_125_3477_n2847) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1994 ( .A1(DP_OP_425J2_127_3477_n1991), 
        .A2(DP_OP_424J2_126_3477_n2785), .Y(DP_OP_424J2_126_3477_n2764) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1152 ( .A1(DP_OP_425J2_127_3477_n2692), 
        .A2(DP_OP_423J2_125_3477_n1947), .Y(DP_OP_423J2_125_3477_n1926) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1680 ( .A1(DP_OP_423J2_125_3477_n2470), 
        .A2(DP_OP_423J2_125_3477_n2475), .Y(DP_OP_423J2_125_3477_n2454) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1673 ( .A1(DP_OP_423J2_125_3477_n2471), 
        .A2(DP_OP_423J2_125_3477_n2474), .Y(DP_OP_423J2_125_3477_n2447) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2001 ( .A1(DP_OP_425J2_127_3477_n1990), 
        .A2(DP_OP_423J2_125_3477_n2781), .Y(DP_OP_424J2_126_3477_n2771) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1012 ( .A1(n371), .A2(n340), .Y(
        DP_OP_424J2_126_3477_n1785) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1327 ( .A1(DP_OP_424J2_126_3477_n2124), 
        .A2(DP_OP_424J2_126_3477_n2127), .Y(DP_OP_424J2_126_3477_n2100) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1937 ( .A1(DP_OP_423J2_125_3477_n2732), 
        .A2(DP_OP_422J2_124_3477_n2740), .Y(DP_OP_423J2_125_3477_n2708) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2082 ( .A1(DP_OP_425J2_127_3477_n1903), 
        .A2(DP_OP_424J2_126_3477_n2873), .Y(DP_OP_424J2_126_3477_n2852) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1686 ( .A1(DP_OP_424J2_126_3477_n2472), 
        .A2(DP_OP_423J2_125_3477_n2475), .Y(DP_OP_424J2_126_3477_n2456) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1768 ( .A1(DP_OP_423J2_125_3477_n2558), 
        .A2(DP_OP_422J2_124_3477_n2567), .Y(DP_OP_423J2_125_3477_n2542) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1145 ( .A1(DP_OP_423J2_125_3477_n1943), 
        .A2(DP_OP_425J2_127_3477_n1951), .Y(DP_OP_423J2_125_3477_n1919) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1907 ( .A1(DP_OP_424J2_126_3477_n2693), 
        .A2(DP_OP_424J2_126_3477_n2697), .Y(DP_OP_424J2_126_3477_n2677) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1409 ( .A1(DP_OP_425J2_127_3477_n2429), 
        .A2(n443), .Y(DP_OP_423J2_125_3477_n2183) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1410 ( .A1(DP_OP_425J2_127_3477_n2430), 
        .A2(n443), .Y(DP_OP_423J2_125_3477_n2184) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1008 ( .A1(n384), .A2(n342), .Y(
        DP_OP_423J2_125_3477_n1782) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1592 ( .A1(DP_OP_424J2_126_3477_n2386), 
        .A2(DP_OP_424J2_126_3477_n2388), .Y(DP_OP_424J2_126_3477_n2362) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1146 ( .A1(DP_OP_425J2_127_3477_n2694), 
        .A2(n442), .Y(DP_OP_423J2_125_3477_n1920) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1151 ( .A1(DP_OP_424J2_126_3477_n1948), 
        .A2(DP_OP_425J2_127_3477_n1951), .Y(DP_OP_424J2_126_3477_n1924) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1415 ( .A1(DP_OP_424J2_126_3477_n2212), 
        .A2(DP_OP_422J2_124_3477_n2214), .Y(DP_OP_424J2_126_3477_n2188) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1153 ( .A1(DP_OP_423J2_125_3477_n1943), 
        .A2(DP_OP_423J2_125_3477_n1947), .Y(DP_OP_423J2_125_3477_n1927) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2077 ( .A1(DP_OP_423J2_125_3477_n2864), 
        .A2(DP_OP_423J2_125_3477_n2868), .Y(DP_OP_423J2_125_3477_n2848) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1584 ( .A1(DP_OP_422J2_124_3477_n2342), 
        .A2(DP_OP_423J2_125_3477_n2386), .Y(DP_OP_423J2_125_3477_n2358) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1591 ( .A1(DP_OP_424J2_126_3477_n2385), 
        .A2(DP_OP_424J2_126_3477_n2388), .Y(DP_OP_424J2_126_3477_n2361) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1989 ( .A1(DP_OP_423J2_125_3477_n2776), 
        .A2(DP_OP_422J2_124_3477_n2785), .Y(DP_OP_423J2_125_3477_n2760) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1899 ( .A1(DP_OP_425J2_127_3477_n2166), 
        .A2(DP_OP_423J2_125_3477_n2695), .Y(DP_OP_423J2_125_3477_n2673) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1901 ( .A1(DP_OP_425J2_127_3477_n2168), 
        .A2(DP_OP_423J2_125_3477_n2695), .Y(DP_OP_423J2_125_3477_n2675) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1987 ( .A1(DP_OP_424J2_126_3477_n2691), 
        .A2(DP_OP_424J2_126_3477_n2785), .Y(DP_OP_423J2_125_3477_n2758) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1159 ( .A1(DP_OP_424J2_126_3477_n1948), 
        .A2(DP_OP_424J2_126_3477_n1952), .Y(DP_OP_424J2_126_3477_n1932) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2080 ( .A1(DP_OP_425J2_127_3477_n1901), 
        .A2(DP_OP_424J2_126_3477_n2873), .Y(DP_OP_424J2_126_3477_n2850) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1739 ( .A1(DP_OP_424J2_126_3477_n2517), 
        .A2(DP_OP_424J2_126_3477_n2522), .Y(DP_OP_424J2_126_3477_n2509) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1736 ( .A1(DP_OP_423J2_125_3477_n2600), 
        .A2(DP_OP_424J2_126_3477_n2522), .Y(DP_OP_424J2_126_3477_n2506) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1678 ( .A1(DP_OP_424J2_126_3477_n2472), 
        .A2(DP_OP_423J2_125_3477_n2474), .Y(DP_OP_424J2_126_3477_n2448) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1942 ( .A1(DP_OP_424J2_126_3477_n2736), 
        .A2(DP_OP_424J2_126_3477_n2740), .Y(DP_OP_424J2_126_3477_n2712) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1685 ( .A1(DP_OP_424J2_126_3477_n2471), 
        .A2(DP_OP_422J2_124_3477_n2479), .Y(DP_OP_424J2_126_3477_n2455) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1151 ( .A1(DP_OP_425J2_127_3477_n2691), 
        .A2(DP_OP_423J2_125_3477_n1947), .Y(DP_OP_423J2_125_3477_n1925) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1414 ( .A1(DP_OP_424J2_126_3477_n2211), 
        .A2(n443), .Y(DP_OP_424J2_126_3477_n2187) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2081 ( .A1(DP_OP_424J2_126_3477_n2867), 
        .A2(DP_OP_424J2_126_3477_n2873), .Y(DP_OP_424J2_126_3477_n2851) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1144 ( .A1(DP_OP_425J2_127_3477_n2692), 
        .A2(n442), .Y(DP_OP_423J2_125_3477_n1918) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1150 ( .A1(DP_OP_425J2_127_3477_n2780), 
        .A2(n442), .Y(DP_OP_424J2_126_3477_n1923) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1590 ( .A1(DP_OP_424J2_126_3477_n2384), 
        .A2(DP_OP_424J2_126_3477_n2388), .Y(DP_OP_424J2_126_3477_n2360) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1905 ( .A1(DP_OP_424J2_126_3477_n2691), 
        .A2(DP_OP_424J2_126_3477_n2697), .Y(DP_OP_424J2_126_3477_n2675) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1670 ( .A1(DP_OP_423J2_125_3477_n2468), 
        .A2(DP_OP_423J2_125_3477_n2474), .Y(DP_OP_423J2_125_3477_n2444) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2000 ( .A1(DP_OP_425J2_127_3477_n1989), 
        .A2(DP_OP_425J2_127_3477_n2786), .Y(DP_OP_424J2_126_3477_n2770) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1326 ( .A1(DP_OP_422J2_124_3477_n2736), 
        .A2(DP_OP_424J2_126_3477_n2127), .Y(DP_OP_424J2_126_3477_n2099) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U982 ( .A1(n316), .A2(n343), .Y(
        DP_OP_423J2_125_3477_n154) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1450 ( .A1(DP_OP_425J2_127_3477_n2382), 
        .A2(DP_OP_423J2_125_3477_n2254), .Y(DP_OP_423J2_125_3477_n2224) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1773 ( .A1(DP_OP_424J2_126_3477_n2559), 
        .A2(DP_OP_424J2_126_3477_n2565), .Y(DP_OP_424J2_126_3477_n2543) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1318 ( .A1(DP_OP_423J2_125_3477_n2116), 
        .A2(DP_OP_423J2_125_3477_n2122), .Y(DP_OP_423J2_125_3477_n2092) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1993 ( .A1(DP_OP_425J2_127_3477_n1990), 
        .A2(DP_OP_424J2_126_3477_n2785), .Y(DP_OP_424J2_126_3477_n2763) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U981 ( .A1(n323), .A2(n340), .Y(
        DP_OP_423J2_125_3477_n152) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1458 ( .A1(DP_OP_422J2_124_3477_n2606), 
        .A2(DP_OP_423J2_125_3477_n2254), .Y(DP_OP_424J2_126_3477_n2231) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1149 ( .A1(DP_OP_423J2_125_3477_n1939), 
        .A2(DP_OP_423J2_125_3477_n1947), .Y(DP_OP_423J2_125_3477_n1923) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2088 ( .A1(DP_OP_425J2_127_3477_n1901), 
        .A2(DP_OP_424J2_126_3477_n2874), .Y(DP_OP_424J2_126_3477_n2858) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U980 ( .A1(n326), .A2(n341), .Y(
        DP_OP_423J2_125_3477_n150) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1897 ( .A1(DP_OP_425J2_127_3477_n2164), 
        .A2(DP_OP_423J2_125_3477_n2695), .Y(DP_OP_423J2_125_3477_n2671) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1120 ( .A1(DP_OP_424J2_126_3477_n1901), 
        .A2(DP_OP_424J2_126_3477_n1909), .Y(DP_OP_424J2_126_3477_n1893) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1985 ( .A1(DP_OP_423J2_125_3477_n2772), 
        .A2(DP_OP_424J2_126_3477_n2785), .Y(DP_OP_423J2_125_3477_n2756) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1582 ( .A1(DP_OP_422J2_124_3477_n2340), 
        .A2(DP_OP_423J2_125_3477_n2386), .Y(DP_OP_423J2_125_3477_n2356) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1677 ( .A1(DP_OP_423J2_125_3477_n2467), 
        .A2(DP_OP_423J2_125_3477_n2475), .Y(DP_OP_423J2_125_3477_n2451) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2073 ( .A1(DP_OP_423J2_125_3477_n2860), 
        .A2(DP_OP_423J2_125_3477_n2868), .Y(DP_OP_423J2_125_3477_n2844) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1142 ( .A1(DP_OP_425J2_127_3477_n2690), 
        .A2(n442), .Y(DP_OP_423J2_125_3477_n1916) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1406 ( .A1(DP_OP_423J2_125_3477_n2204), 
        .A2(n443), .Y(DP_OP_423J2_125_3477_n2180) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1676 ( .A1(DP_OP_425J2_127_3477_n2297), 
        .A2(DP_OP_423J2_125_3477_n2474), .Y(DP_OP_424J2_126_3477_n2446) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1934 ( .A1(DP_OP_423J2_125_3477_n2729), 
        .A2(DP_OP_422J2_124_3477_n2740), .Y(DP_OP_423J2_125_3477_n2705) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1456 ( .A1(DP_OP_422J2_124_3477_n2604), 
        .A2(DP_OP_425J2_127_3477_n2259), .Y(DP_OP_424J2_126_3477_n2229) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1765 ( .A1(DP_OP_425J2_127_3477_n2296), 
        .A2(DP_OP_424J2_126_3477_n2565), .Y(DP_OP_423J2_125_3477_n2539) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1324 ( .A1(DP_OP_423J2_125_3477_n2028), 
        .A2(DP_OP_424J2_126_3477_n2127), .Y(DP_OP_424J2_126_3477_n2097) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1009 ( .A1(n293), .A2(n343), .Y(
        DP_OP_423J2_125_3477_n1783) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1154 ( .A1(DP_OP_425J2_127_3477_n2694), 
        .A2(DP_OP_423J2_125_3477_n1947), .Y(DP_OP_423J2_125_3477_n1928) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2092 ( .A1(DP_OP_425J2_127_3477_n1905), 
        .A2(DP_OP_424J2_126_3477_n2874), .Y(DP_OP_424J2_126_3477_n2862) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1740 ( .A1(DP_OP_423J2_125_3477_n2604), 
        .A2(DP_OP_424J2_126_3477_n2522), .Y(DP_OP_424J2_126_3477_n2510) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2004 ( .A1(DP_OP_422J2_124_3477_n1861), 
        .A2(DP_OP_423J2_125_3477_n2781), .Y(DP_OP_424J2_126_3477_n2774) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1015 ( .A1(n278), .A2(n339), .Y(
        DP_OP_424J2_126_3477_n1788) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1124 ( .A1(DP_OP_425J2_127_3477_n2826), 
        .A2(DP_OP_424J2_126_3477_n1909), .Y(DP_OP_424J2_126_3477_n1897) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2078 ( .A1(DP_OP_423J2_125_3477_n2865), 
        .A2(DP_OP_423J2_125_3477_n2868), .Y(DP_OP_423J2_125_3477_n2849) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1990 ( .A1(DP_OP_423J2_125_3477_n2777), 
        .A2(DP_OP_422J2_124_3477_n2785), .Y(DP_OP_423J2_125_3477_n2761) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1682 ( .A1(DP_OP_423J2_125_3477_n2472), 
        .A2(DP_OP_423J2_125_3477_n2475), .Y(DP_OP_423J2_125_3477_n2456) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1902 ( .A1(DP_OP_425J2_127_3477_n2169), 
        .A2(DP_OP_423J2_125_3477_n2695), .Y(DP_OP_423J2_125_3477_n2676) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1770 ( .A1(DP_OP_422J2_124_3477_n2168), 
        .A2(DP_OP_424J2_126_3477_n2565), .Y(DP_OP_423J2_125_3477_n2544) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1005 ( .A1(n273), .A2(n340), .Y(
        DP_OP_423J2_125_3477_n1779) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1452 ( .A1(DP_OP_422J2_124_3477_n2518), 
        .A2(DP_OP_423J2_125_3477_n2254), .Y(DP_OP_423J2_125_3477_n2226) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2082 ( .A1(DP_OP_423J2_125_3477_n2861), 
        .A2(DP_OP_423J2_125_3477_n2869), .Y(DP_OP_423J2_125_3477_n2853) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2085 ( .A1(DP_OP_423J2_125_3477_n2864), 
        .A2(DP_OP_423J2_125_3477_n2869), .Y(DP_OP_423J2_125_3477_n2856) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1733 ( .A1(DP_OP_423J2_125_3477_n2515), 
        .A2(DP_OP_423J2_125_3477_n2520), .Y(DP_OP_423J2_125_3477_n2507) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1908 ( .A1(DP_OP_422J2_124_3477_n1949), 
        .A2(DP_OP_424J2_126_3477_n2697), .Y(DP_OP_424J2_126_3477_n2678) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1160 ( .A1(DP_OP_424J2_126_3477_n1949), 
        .A2(DP_OP_424J2_126_3477_n1952), .Y(DP_OP_424J2_126_3477_n1933) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1114 ( .A1(DP_OP_423J2_125_3477_n1896), 
        .A2(DP_OP_423J2_125_3477_n1904), .Y(DP_OP_423J2_125_3477_n1888) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1672 ( .A1(DP_OP_423J2_125_3477_n2470), 
        .A2(DP_OP_423J2_125_3477_n2474), .Y(DP_OP_423J2_125_3477_n2446) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1730 ( .A1(DP_OP_425J2_127_3477_n2341), 
        .A2(DP_OP_423J2_125_3477_n2520), .Y(DP_OP_423J2_125_3477_n2504) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1994 ( .A1(DP_OP_425J2_127_3477_n2077), 
        .A2(DP_OP_423J2_125_3477_n2781), .Y(DP_OP_423J2_125_3477_n2765) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1117 ( .A1(DP_OP_423J2_125_3477_n1899), 
        .A2(DP_OP_423J2_125_3477_n1904), .Y(DP_OP_423J2_125_3477_n1891) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1688 ( .A1(DP_OP_424J2_126_3477_n2474), 
        .A2(DP_OP_423J2_125_3477_n2475), .Y(DP_OP_424J2_126_3477_n2458) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2084 ( .A1(DP_OP_425J2_127_3477_n1905), 
        .A2(DP_OP_424J2_126_3477_n2873), .Y(DP_OP_424J2_126_3477_n2854) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1320 ( .A1(DP_OP_422J2_124_3477_n2650), 
        .A2(DP_OP_423J2_125_3477_n2122), .Y(DP_OP_423J2_125_3477_n2094) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1996 ( .A1(DP_OP_423J2_125_3477_n2865), 
        .A2(DP_OP_424J2_126_3477_n2785), .Y(DP_OP_424J2_126_3477_n2766) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1776 ( .A1(DP_OP_425J2_127_3477_n2213), 
        .A2(DP_OP_424J2_126_3477_n2565), .Y(DP_OP_424J2_126_3477_n2546) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2003 ( .A1(DP_OP_423J2_125_3477_n2864), 
        .A2(DP_OP_425J2_127_3477_n2786), .Y(DP_OP_424J2_126_3477_n2773) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1123 ( .A1(DP_OP_424J2_126_3477_n1904), 
        .A2(DP_OP_424J2_126_3477_n1909), .Y(DP_OP_424J2_126_3477_n1896) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2091 ( .A1(DP_OP_424J2_126_3477_n2869), 
        .A2(DP_OP_424J2_126_3477_n2874), .Y(DP_OP_424J2_126_3477_n2861) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1411 ( .A1(DP_OP_423J2_125_3477_n2643), 
        .A2(DP_OP_425J2_127_3477_n2215), .Y(DP_OP_425J2_127_3477_n2184) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1939 ( .A1(DP_OP_424J2_126_3477_n1988), 
        .A2(DP_OP_425J2_127_3477_n2740), .Y(DP_OP_425J2_127_3477_n2709) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1323 ( .A1(DP_OP_425J2_127_3477_n2120), 
        .A2(DP_OP_425J2_127_3477_n2127), .Y(DP_OP_425J2_127_3477_n2096) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1676 ( .A1(DP_OP_423J2_125_3477_n2160), 
        .A2(DP_OP_425J2_127_3477_n2476), .Y(DP_OP_425J2_127_3477_n2446) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1324 ( .A1(DP_OP_423J2_125_3477_n2729), 
        .A2(DP_OP_425J2_127_3477_n2127), .Y(DP_OP_425J2_127_3477_n2097) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1999 ( .A1(DP_OP_425J2_127_3477_n2777), 
        .A2(DP_OP_425J2_127_3477_n2786), .Y(DP_OP_425J2_127_3477_n2769) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1149 ( .A1(DP_OP_423J2_125_3477_n2906), 
        .A2(DP_OP_425J2_127_3477_n1951), .Y(DP_OP_425J2_127_3477_n1922) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1010 ( .A1(n268), .A2(n340), .Y(
        DP_OP_425J2_127_3477_n1783) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U999 ( .A1(n283), .A2(n341), .Y(
        DP_OP_423J2_125_3477_n1773) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2080 ( .A1(DP_OP_424J2_126_3477_n1857), 
        .A2(DP_OP_423J2_125_3477_n2868), .Y(DP_OP_425J2_127_3477_n2850) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1455 ( .A1(DP_OP_425J2_127_3477_n2252), 
        .A2(DP_OP_425J2_127_3477_n2259), .Y(DP_OP_425J2_127_3477_n2228) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1771 ( .A1(DP_OP_425J2_127_3477_n2557), 
        .A2(DP_OP_425J2_127_3477_n2565), .Y(DP_OP_425J2_127_3477_n2541) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2087 ( .A1(DP_OP_425J2_127_3477_n2865), 
        .A2(DP_OP_425J2_127_3477_n2874), .Y(DP_OP_425J2_127_3477_n2857) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1735 ( .A1(DP_OP_422J2_124_3477_n2647), 
        .A2(DP_OP_423J2_125_3477_n2520), .Y(DP_OP_425J2_127_3477_n2505) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1325 ( .A1(DP_OP_425J2_127_3477_n2122), 
        .A2(DP_OP_425J2_127_3477_n2127), .Y(DP_OP_425J2_127_3477_n2098) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1148 ( .A1(DP_OP_425J2_127_3477_n1945), 
        .A2(DP_OP_425J2_127_3477_n1951), .Y(DP_OP_425J2_127_3477_n1921) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1940 ( .A1(DP_OP_425J2_127_3477_n2734), 
        .A2(DP_OP_425J2_127_3477_n2740), .Y(DP_OP_425J2_127_3477_n2710) );
  XNOR2X1_HVT DP_OP_425J2_127_3477_U627 ( .A1(DP_OP_425J2_127_3477_n2703), 
        .A2(DP_OP_425J2_127_3477_n2352), .Y(DP_OP_425J2_127_3477_n1062) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1456 ( .A1(DP_OP_422J2_124_3477_n2120), 
        .A2(DP_OP_425J2_127_3477_n2259), .Y(DP_OP_425J2_127_3477_n2229) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1683 ( .A1(DP_OP_425J2_127_3477_n2469), 
        .A2(DP_OP_425J2_127_3477_n2477), .Y(DP_OP_425J2_127_3477_n2453) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1991 ( .A1(DP_OP_425J2_127_3477_n2777), 
        .A2(DP_OP_425J2_127_3477_n2785), .Y(DP_OP_425J2_127_3477_n2761) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2000 ( .A1(DP_OP_425J2_127_3477_n2778), 
        .A2(DP_OP_425J2_127_3477_n2786), .Y(DP_OP_425J2_127_3477_n2770) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1992 ( .A1(DP_OP_423J2_125_3477_n2861), 
        .A2(DP_OP_424J2_126_3477_n2785), .Y(DP_OP_424J2_126_3477_n2762) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1678 ( .A1(DP_OP_425J2_127_3477_n2472), 
        .A2(DP_OP_425J2_127_3477_n2476), .Y(DP_OP_425J2_127_3477_n2448) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1941 ( .A1(DP_OP_424J2_126_3477_n2735), 
        .A2(DP_OP_424J2_126_3477_n2740), .Y(DP_OP_424J2_126_3477_n2711) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1992 ( .A1(DP_OP_425J2_127_3477_n2778), 
        .A2(DP_OP_425J2_127_3477_n2785), .Y(DP_OP_425J2_127_3477_n2762) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1458 ( .A1(DP_OP_425J2_127_3477_n2255), 
        .A2(DP_OP_425J2_127_3477_n2259), .Y(DP_OP_425J2_127_3477_n2231) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1684 ( .A1(DP_OP_423J2_125_3477_n2160), 
        .A2(DP_OP_425J2_127_3477_n2477), .Y(DP_OP_425J2_127_3477_n2454) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1903 ( .A1(DP_OP_423J2_125_3477_n1939), 
        .A2(DP_OP_422J2_124_3477_n2699), .Y(DP_OP_425J2_127_3477_n2673) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1155 ( .A1(DP_OP_423J2_125_3477_n2904), 
        .A2(DP_OP_423J2_125_3477_n1947), .Y(DP_OP_425J2_127_3477_n1928) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1003 ( .A1(n404), .A2(n340), .Y(
        DP_OP_424J2_126_3477_n1776) );
  OR2X1_HVT DP_OP_423J2_125_3477_U978 ( .A1(n380), .A2(n340), .Y(
        DP_OP_423J2_125_3477_n1768) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1007 ( .A1(n276), .A2(n343), .Y(
        DP_OP_424J2_126_3477_n1780) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U979 ( .A1(n320), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_423J2_125_3477_n148) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1414 ( .A1(DP_OP_422J2_124_3477_n2078), 
        .A2(DP_OP_425J2_127_3477_n2215), .Y(DP_OP_425J2_127_3477_n2187) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1736 ( .A1(DP_OP_423J2_125_3477_n2116), 
        .A2(DP_OP_424J2_126_3477_n2522), .Y(DP_OP_425J2_127_3477_n2506) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2088 ( .A1(DP_OP_424J2_126_3477_n1857), 
        .A2(DP_OP_425J2_127_3477_n2874), .Y(DP_OP_425J2_127_3477_n2858) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1735 ( .A1(DP_OP_423J2_125_3477_n2599), 
        .A2(DP_OP_424J2_126_3477_n2522), .Y(DP_OP_424J2_126_3477_n2505) );
  OR2X1_HVT DP_OP_424J2_126_3477_U33 ( .A1(DP_OP_424J2_126_3477_n179), .A2(
        DP_OP_424J2_126_3477_n178), .Y(DP_OP_424J2_126_3477_n45) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1150 ( .A1(DP_OP_423J2_125_3477_n2907), 
        .A2(DP_OP_425J2_127_3477_n1951), .Y(DP_OP_425J2_127_3477_n1923) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1999 ( .A1(DP_OP_424J2_126_3477_n2777), 
        .A2(DP_OP_423J2_125_3477_n2781), .Y(DP_OP_424J2_126_3477_n2769) );
  OR2X1_HVT DP_OP_424J2_126_3477_U984 ( .A1(n314), .A2(n343), .Y(
        DP_OP_424J2_126_3477_n1773) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1140 ( .A1(DP_OP_425J2_127_3477_n2688), 
        .A2(n442), .Y(DP_OP_423J2_125_3477_n1914) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1457 ( .A1(DP_OP_422J2_124_3477_n2605), 
        .A2(DP_OP_425J2_127_3477_n2259), .Y(DP_OP_424J2_126_3477_n2230) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1326 ( .A1(DP_OP_423J2_125_3477_n2731), 
        .A2(DP_OP_425J2_127_3477_n2127), .Y(DP_OP_425J2_127_3477_n2099) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1942 ( .A1(DP_OP_423J2_125_3477_n1898), 
        .A2(DP_OP_425J2_127_3477_n2740), .Y(DP_OP_425J2_127_3477_n2712) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1412 ( .A1(DP_OP_425J2_127_3477_n2209), 
        .A2(DP_OP_425J2_127_3477_n2215), .Y(DP_OP_425J2_127_3477_n2185) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1149 ( .A1(DP_OP_425J2_127_3477_n2779), 
        .A2(n442), .Y(DP_OP_424J2_126_3477_n1922) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1685 ( .A1(DP_OP_423J2_125_3477_n2161), 
        .A2(DP_OP_425J2_127_3477_n2477), .Y(DP_OP_425J2_127_3477_n2455) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1993 ( .A1(DP_OP_425J2_127_3477_n2779), 
        .A2(DP_OP_425J2_127_3477_n2785), .Y(DP_OP_425J2_127_3477_n2763) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1772 ( .A1(DP_OP_425J2_127_3477_n2558), 
        .A2(DP_OP_425J2_127_3477_n2565), .Y(DP_OP_425J2_127_3477_n2542) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1156 ( .A1(DP_OP_425J2_127_3477_n2778), 
        .A2(DP_OP_424J2_126_3477_n1952), .Y(DP_OP_424J2_126_3477_n1929) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1773 ( .A1(DP_OP_425J2_127_3477_n2559), 
        .A2(DP_OP_425J2_127_3477_n2565), .Y(DP_OP_425J2_127_3477_n2543) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1147 ( .A1(DP_OP_423J2_125_3477_n2904), 
        .A2(DP_OP_425J2_127_3477_n1951), .Y(DP_OP_425J2_127_3477_n1920) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2081 ( .A1(DP_OP_424J2_126_3477_n1858), 
        .A2(DP_OP_423J2_125_3477_n2868), .Y(DP_OP_425J2_127_3477_n2851) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U998 ( .A1(n281), .A2(n341), .Y(
        DP_OP_423J2_125_3477_n1772) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1675 ( .A1(DP_OP_425J2_127_3477_n2469), 
        .A2(DP_OP_425J2_127_3477_n2476), .Y(DP_OP_425J2_127_3477_n2445) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1413 ( .A1(DP_OP_423J2_125_3477_n2645), 
        .A2(DP_OP_425J2_127_3477_n2215), .Y(DP_OP_425J2_127_3477_n2186) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1677 ( .A1(DP_OP_423J2_125_3477_n2161), 
        .A2(DP_OP_425J2_127_3477_n2476), .Y(DP_OP_425J2_127_3477_n2447) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1457 ( .A1(DP_OP_423J2_125_3477_n2601), 
        .A2(DP_OP_425J2_127_3477_n2259), .Y(DP_OP_425J2_127_3477_n2230) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1941 ( .A1(DP_OP_425J2_127_3477_n2735), 
        .A2(DP_OP_425J2_127_3477_n2740), .Y(DP_OP_425J2_127_3477_n2711) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1413 ( .A1(DP_OP_423J2_125_3477_n2117), 
        .A2(n443), .Y(DP_OP_424J2_126_3477_n2186) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1589 ( .A1(DP_OP_424J2_126_3477_n2383), 
        .A2(DP_OP_424J2_126_3477_n2388), .Y(DP_OP_424J2_126_3477_n2359) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1588 ( .A1(DP_OP_425J2_127_3477_n2382), 
        .A2(DP_OP_423J2_125_3477_n2386), .Y(DP_OP_425J2_127_3477_n2358) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1904 ( .A1(DP_OP_425J2_127_3477_n2077), 
        .A2(DP_OP_424J2_126_3477_n2697), .Y(DP_OP_424J2_126_3477_n2674) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1011 ( .A1(n272), .A2(n342), .Y(
        DP_OP_425J2_127_3477_n1784) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1281 ( .A1(DP_OP_423J2_125_3477_n2645), 
        .A2(DP_OP_422J2_124_3477_n2082), .Y(DP_OP_422J2_124_3477_n2053) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1197 ( .A1(DP_OP_422J2_124_3477_n2781), 
        .A2(DP_OP_423J2_125_3477_n1991), .Y(DP_OP_423J2_125_3477_n1971) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1542 ( .A1(DP_OP_422J2_124_3477_n2432), 
        .A2(DP_OP_425J2_127_3477_n2347), .Y(DP_OP_423J2_125_3477_n2316) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1200 ( .A1(DP_OP_422J2_124_3477_n1989), 
        .A2(DP_OP_422J2_124_3477_n1996), .Y(DP_OP_422J2_124_3477_n1973) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1282 ( .A1(DP_OP_422J2_124_3477_n2078), 
        .A2(DP_OP_422J2_124_3477_n2082), .Y(DP_OP_422J2_124_3477_n2054) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1278 ( .A1(DP_OP_423J2_125_3477_n2076), 
        .A2(n447), .Y(DP_OP_423J2_125_3477_n2052) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2029 ( .A1(DP_OP_424J2_126_3477_n2034), 
        .A2(DP_OP_423J2_125_3477_n2823), .Y(DP_OP_422J2_124_3477_n2799) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1055 ( .A1(DP_OP_423J2_125_3477_n1853), 
        .A2(DP_OP_423J2_125_3477_n1858), .Y(DP_OP_423J2_125_3477_n1829) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1060 ( .A1(DP_OP_425J2_127_3477_n1989), 
        .A2(DP_OP_422J2_124_3477_n1863), .Y(DP_OP_422J2_124_3477_n1833) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1057 ( .A1(DP_OP_424J2_126_3477_n1948), 
        .A2(DP_OP_423J2_125_3477_n1858), .Y(DP_OP_423J2_125_3477_n1831) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2024 ( .A1(DP_OP_424J2_126_3477_n2736), 
        .A2(DP_OP_423J2_125_3477_n2823), .Y(DP_OP_423J2_125_3477_n2795) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1850 ( .A1(DP_OP_423J2_125_3477_n2648), 
        .A2(DP_OP_422J2_124_3477_n2654), .Y(DP_OP_423J2_125_3477_n2624) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2039 ( .A1(DP_OP_422J2_124_3477_n1902), 
        .A2(DP_OP_424J2_126_3477_n2830), .Y(DP_OP_423J2_125_3477_n2810) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1544 ( .A1(DP_OP_422J2_124_3477_n2340), 
        .A2(DP_OP_422J2_124_3477_n2346), .Y(DP_OP_422J2_124_3477_n2316) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1541 ( .A1(DP_OP_423J2_125_3477_n2339), 
        .A2(DP_OP_425J2_127_3477_n2347), .Y(DP_OP_423J2_125_3477_n2315) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2026 ( .A1(DP_OP_422J2_124_3477_n1905), 
        .A2(DP_OP_423J2_125_3477_n2823), .Y(DP_OP_423J2_125_3477_n2797) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2040 ( .A1(DP_OP_422J2_124_3477_n1903), 
        .A2(DP_OP_424J2_126_3477_n2830), .Y(DP_OP_423J2_125_3477_n2811) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1058 ( .A1(DP_OP_423J2_125_3477_n1856), 
        .A2(DP_OP_423J2_125_3477_n1858), .Y(DP_OP_423J2_125_3477_n1832) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1196 ( .A1(DP_OP_423J2_125_3477_n1986), 
        .A2(DP_OP_423J2_125_3477_n1991), .Y(DP_OP_423J2_125_3477_n1970) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1280 ( .A1(DP_OP_422J2_124_3477_n2076), 
        .A2(DP_OP_422J2_124_3477_n2082), .Y(DP_OP_422J2_124_3477_n2052) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1056 ( .A1(DP_OP_425J2_127_3477_n2780), 
        .A2(DP_OP_423J2_125_3477_n1858), .Y(DP_OP_423J2_125_3477_n1830) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1849 ( .A1(DP_OP_423J2_125_3477_n2647), 
        .A2(DP_OP_425J2_127_3477_n2652), .Y(DP_OP_423J2_125_3477_n2623) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1199 ( .A1(DP_OP_422J2_124_3477_n1988), 
        .A2(DP_OP_422J2_124_3477_n1996), .Y(DP_OP_422J2_124_3477_n1972) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1062 ( .A1(DP_OP_422J2_124_3477_n1859), 
        .A2(DP_OP_422J2_124_3477_n1863), .Y(DP_OP_422J2_124_3477_n1835) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1277 ( .A1(DP_OP_422J2_124_3477_n2695), 
        .A2(DP_OP_425J2_127_3477_n2083), .Y(DP_OP_423J2_125_3477_n2051) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2025 ( .A1(DP_OP_424J2_126_3477_n2737), 
        .A2(DP_OP_423J2_125_3477_n2823), .Y(DP_OP_423J2_125_3477_n2796) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2047 ( .A1(DP_OP_422J2_124_3477_n2825), 
        .A2(DP_OP_422J2_124_3477_n2830), .Y(DP_OP_422J2_124_3477_n2817) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1204 ( .A1(DP_OP_424J2_126_3477_n2650), 
        .A2(DP_OP_422J2_124_3477_n1996), .Y(DP_OP_422J2_124_3477_n1977) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2043 ( .A1(DP_OP_424J2_126_3477_n2032), 
        .A2(DP_OP_422J2_124_3477_n2830), .Y(DP_OP_422J2_124_3477_n2813) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1546 ( .A1(DP_OP_422J2_124_3477_n2342), 
        .A2(DP_OP_422J2_124_3477_n2346), .Y(DP_OP_422J2_124_3477_n2318) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2048 ( .A1(DP_OP_424J2_126_3477_n2037), 
        .A2(DP_OP_422J2_124_3477_n2830), .Y(DP_OP_422J2_124_3477_n2818) );
  OR2X1_HVT DP_OP_423J2_125_3477_U33 ( .A1(DP_OP_423J2_125_3477_n174), .A2(
        DP_OP_423J2_125_3477_n173), .Y(DP_OP_423J2_125_3477_n43) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1063 ( .A1(DP_OP_425J2_127_3477_n1992), 
        .A2(DP_OP_422J2_124_3477_n1863), .Y(DP_OP_422J2_124_3477_n1836) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1274 ( .A1(DP_OP_422J2_124_3477_n2692), 
        .A2(DP_OP_425J2_127_3477_n2083), .Y(DP_OP_423J2_125_3477_n2048) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2031 ( .A1(DP_OP_422J2_124_3477_n2825), 
        .A2(DP_OP_424J2_126_3477_n2828), .Y(DP_OP_422J2_124_3477_n2801) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1538 ( .A1(DP_OP_422J2_124_3477_n2428), 
        .A2(n448), .Y(DP_OP_423J2_125_3477_n2312) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2022 ( .A1(DP_OP_424J2_126_3477_n2734), 
        .A2(DP_OP_423J2_125_3477_n2823), .Y(DP_OP_423J2_125_3477_n2793) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1846 ( .A1(DP_OP_425J2_127_3477_n2209), 
        .A2(DP_OP_425J2_127_3477_n2652), .Y(DP_OP_423J2_125_3477_n2620) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2027 ( .A1(DP_OP_424J2_126_3477_n2032), 
        .A2(DP_OP_423J2_125_3477_n2823), .Y(DP_OP_422J2_124_3477_n2797) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1193 ( .A1(DP_OP_423J2_125_3477_n1983), 
        .A2(DP_OP_423J2_125_3477_n1991), .Y(DP_OP_423J2_125_3477_n1967) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1847 ( .A1(DP_OP_423J2_125_3477_n2645), 
        .A2(DP_OP_424J2_126_3477_n2652), .Y(DP_OP_423J2_125_3477_n2621) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2032 ( .A1(DP_OP_424J2_126_3477_n2037), 
        .A2(DP_OP_423J2_125_3477_n2823), .Y(DP_OP_422J2_124_3477_n2802) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1202 ( .A1(DP_OP_422J2_124_3477_n1991), 
        .A2(DP_OP_422J2_124_3477_n1996), .Y(DP_OP_422J2_124_3477_n1975) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2045 ( .A1(DP_OP_424J2_126_3477_n2034), 
        .A2(DP_OP_422J2_124_3477_n2830), .Y(DP_OP_422J2_124_3477_n2815) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2038 ( .A1(DP_OP_424J2_126_3477_n2734), 
        .A2(DP_OP_425J2_127_3477_n2830), .Y(DP_OP_423J2_125_3477_n2809) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2023 ( .A1(DP_OP_422J2_124_3477_n1902), 
        .A2(DP_OP_423J2_125_3477_n2823), .Y(DP_OP_423J2_125_3477_n2794) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2046 ( .A1(DP_OP_424J2_126_3477_n2035), 
        .A2(DP_OP_422J2_124_3477_n2830), .Y(DP_OP_422J2_124_3477_n2816) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1203 ( .A1(DP_OP_424J2_126_3477_n2649), 
        .A2(DP_OP_422J2_124_3477_n1996), .Y(DP_OP_422J2_124_3477_n1976) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1275 ( .A1(DP_OP_423J2_125_3477_n2073), 
        .A2(DP_OP_422J2_124_3477_n2082), .Y(DP_OP_423J2_125_3477_n2049) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1855 ( .A1(DP_OP_422J2_124_3477_n2651), 
        .A2(DP_OP_422J2_124_3477_n2654), .Y(DP_OP_422J2_124_3477_n2627) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1276 ( .A1(DP_OP_423J2_125_3477_n2074), 
        .A2(DP_OP_425J2_127_3477_n2083), .Y(DP_OP_423J2_125_3477_n2050) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1195 ( .A1(DP_OP_423J2_125_3477_n1985), 
        .A2(DP_OP_423J2_125_3477_n1991), .Y(DP_OP_423J2_125_3477_n1969) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1539 ( .A1(DP_OP_422J2_124_3477_n2429), 
        .A2(n448), .Y(DP_OP_423J2_125_3477_n2313) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1540 ( .A1(DP_OP_422J2_124_3477_n2430), 
        .A2(DP_OP_422J2_124_3477_n2346), .Y(DP_OP_423J2_125_3477_n2314) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1543 ( .A1(DP_OP_422J2_124_3477_n2339), 
        .A2(DP_OP_422J2_124_3477_n2346), .Y(DP_OP_422J2_124_3477_n2315) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1547 ( .A1(DP_OP_422J2_124_3477_n2343), 
        .A2(DP_OP_422J2_124_3477_n2346), .Y(DP_OP_422J2_124_3477_n2319) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1537 ( .A1(DP_OP_422J2_124_3477_n2427), 
        .A2(DP_OP_425J2_127_3477_n2347), .Y(DP_OP_423J2_125_3477_n2311) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2021 ( .A1(DP_OP_422J2_124_3477_n1900), 
        .A2(DP_OP_423J2_125_3477_n2823), .Y(DP_OP_423J2_125_3477_n2792) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1845 ( .A1(DP_OP_423J2_125_3477_n2643), 
        .A2(DP_OP_422J2_124_3477_n2654), .Y(DP_OP_423J2_125_3477_n2619) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1053 ( .A1(DP_OP_425J2_127_3477_n2777), 
        .A2(DP_OP_423J2_125_3477_n1858), .Y(DP_OP_423J2_125_3477_n1827) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1851 ( .A1(DP_OP_422J2_124_3477_n2647), 
        .A2(DP_OP_422J2_124_3477_n2654), .Y(DP_OP_422J2_124_3477_n2623) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1283 ( .A1(DP_OP_423J2_125_3477_n2647), 
        .A2(DP_OP_422J2_124_3477_n2082), .Y(DP_OP_422J2_124_3477_n2055) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1273 ( .A1(DP_OP_424J2_126_3477_n2164), 
        .A2(n447), .Y(DP_OP_423J2_125_3477_n2047) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1059 ( .A1(DP_OP_424J2_126_3477_n2777), 
        .A2(DP_OP_422J2_124_3477_n1863), .Y(DP_OP_422J2_124_3477_n1832) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1054 ( .A1(DP_OP_423J2_125_3477_n1852), 
        .A2(DP_OP_423J2_125_3477_n1858), .Y(DP_OP_423J2_125_3477_n1828) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1284 ( .A1(DP_OP_423J2_125_3477_n2648), 
        .A2(DP_OP_422J2_124_3477_n2082), .Y(DP_OP_422J2_124_3477_n2056) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1548 ( .A1(DP_OP_422J2_124_3477_n2344), 
        .A2(DP_OP_422J2_124_3477_n2346), .Y(DP_OP_422J2_124_3477_n2320) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2028 ( .A1(DP_OP_424J2_126_3477_n2033), 
        .A2(DP_OP_423J2_125_3477_n2823), .Y(DP_OP_422J2_124_3477_n2798) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1852 ( .A1(DP_OP_422J2_124_3477_n2648), 
        .A2(DP_OP_422J2_124_3477_n2654), .Y(DP_OP_422J2_124_3477_n2624) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2041 ( .A1(DP_OP_424J2_126_3477_n2737), 
        .A2(DP_OP_422J2_124_3477_n2830), .Y(DP_OP_423J2_125_3477_n2812) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1198 ( .A1(DP_OP_425J2_127_3477_n2650), 
        .A2(DP_OP_423J2_125_3477_n1991), .Y(DP_OP_423J2_125_3477_n1972) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1061 ( .A1(DP_OP_422J2_124_3477_n1858), 
        .A2(DP_OP_422J2_124_3477_n1863), .Y(DP_OP_422J2_124_3477_n1834) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2037 ( .A1(DP_OP_422J2_124_3477_n1900), 
        .A2(DP_OP_422J2_124_3477_n2830), .Y(DP_OP_423J2_125_3477_n2808) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1545 ( .A1(DP_OP_422J2_124_3477_n2341), 
        .A2(DP_OP_422J2_124_3477_n2346), .Y(DP_OP_422J2_124_3477_n2317) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1853 ( .A1(DP_OP_422J2_124_3477_n2649), 
        .A2(DP_OP_422J2_124_3477_n2654), .Y(DP_OP_422J2_124_3477_n2625) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1279 ( .A1(DP_OP_424J2_126_3477_n2557), 
        .A2(DP_OP_422J2_124_3477_n2082), .Y(DP_OP_422J2_124_3477_n2051) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1848 ( .A1(DP_OP_423J2_125_3477_n2646), 
        .A2(DP_OP_422J2_124_3477_n2654), .Y(DP_OP_423J2_125_3477_n2622) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1194 ( .A1(DP_OP_424J2_126_3477_n2077), 
        .A2(DP_OP_423J2_125_3477_n1991), .Y(DP_OP_423J2_125_3477_n1968) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1856 ( .A1(DP_OP_422J2_124_3477_n2652), 
        .A2(DP_OP_422J2_124_3477_n2654), .Y(DP_OP_422J2_124_3477_n2628) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2042 ( .A1(DP_OP_424J2_126_3477_n2738), 
        .A2(DP_OP_422J2_124_3477_n2830), .Y(DP_OP_423J2_125_3477_n2813) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2030 ( .A1(DP_OP_424J2_126_3477_n2035), 
        .A2(DP_OP_424J2_126_3477_n2828), .Y(DP_OP_422J2_124_3477_n2800) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2044 ( .A1(DP_OP_424J2_126_3477_n2033), 
        .A2(DP_OP_422J2_124_3477_n2830), .Y(DP_OP_422J2_124_3477_n2814) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1064 ( .A1(DP_OP_422J2_124_3477_n1861), 
        .A2(DP_OP_422J2_124_3477_n1863), .Y(DP_OP_422J2_124_3477_n1837) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1201 ( .A1(DP_OP_425J2_127_3477_n2122), 
        .A2(DP_OP_422J2_124_3477_n1996), .Y(DP_OP_422J2_124_3477_n1974) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1854 ( .A1(DP_OP_422J2_124_3477_n2650), 
        .A2(DP_OP_422J2_124_3477_n2654), .Y(DP_OP_422J2_124_3477_n2626) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1855 ( .A1(DP_OP_425J2_127_3477_n2649), 
        .A2(DP_OP_425J2_127_3477_n2652), .Y(DP_OP_425J2_127_3477_n2625) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1064 ( .A1(DP_OP_425J2_127_3477_n2870), 
        .A2(DP_OP_425J2_127_3477_n1863), .Y(DP_OP_424J2_126_3477_n1837) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1548 ( .A1(DP_OP_422J2_124_3477_n2520), 
        .A2(n448), .Y(DP_OP_424J2_126_3477_n2321) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1284 ( .A1(DP_OP_422J2_124_3477_n2782), 
        .A2(n447), .Y(DP_OP_424J2_126_3477_n2057) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1856 ( .A1(DP_OP_424J2_126_3477_n2650), 
        .A2(DP_OP_424J2_126_3477_n2652), .Y(DP_OP_424J2_126_3477_n2626) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2046 ( .A1(DP_OP_424J2_126_3477_n2824), 
        .A2(DP_OP_424J2_126_3477_n2830), .Y(DP_OP_424J2_126_3477_n2816) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2032 ( .A1(DP_OP_424J2_126_3477_n2826), 
        .A2(DP_OP_424J2_126_3477_n2828), .Y(DP_OP_424J2_126_3477_n2802) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1203 ( .A1(DP_OP_422J2_124_3477_n2869), 
        .A2(DP_OP_424J2_126_3477_n1996), .Y(DP_OP_424J2_126_3477_n1976) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2047 ( .A1(DP_OP_424J2_126_3477_n2825), 
        .A2(DP_OP_424J2_126_3477_n2830), .Y(DP_OP_424J2_126_3477_n2817) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1204 ( .A1(DP_OP_422J2_124_3477_n2870), 
        .A2(DP_OP_424J2_126_3477_n1996), .Y(DP_OP_424J2_126_3477_n1977) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2048 ( .A1(DP_OP_424J2_126_3477_n2826), 
        .A2(DP_OP_424J2_126_3477_n2830), .Y(DP_OP_424J2_126_3477_n2818) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2028 ( .A1(DP_OP_424J2_126_3477_n2822), 
        .A2(DP_OP_424J2_126_3477_n2828), .Y(DP_OP_424J2_126_3477_n2798) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1544 ( .A1(DP_OP_424J2_126_3477_n2341), 
        .A2(n448), .Y(DP_OP_424J2_126_3477_n2317) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1199 ( .A1(DP_OP_424J2_126_3477_n1988), 
        .A2(DP_OP_424J2_126_3477_n1996), .Y(DP_OP_424J2_126_3477_n1972) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1852 ( .A1(DP_OP_422J2_124_3477_n1989), 
        .A2(DP_OP_424J2_126_3477_n2652), .Y(DP_OP_424J2_126_3477_n2622) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1280 ( .A1(DP_OP_424J2_126_3477_n2077), 
        .A2(n447), .Y(DP_OP_424J2_126_3477_n2053) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1282 ( .A1(DP_OP_422J2_124_3477_n2780), 
        .A2(n447), .Y(DP_OP_424J2_126_3477_n2055) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2030 ( .A1(DP_OP_424J2_126_3477_n2824), 
        .A2(DP_OP_424J2_126_3477_n2828), .Y(DP_OP_424J2_126_3477_n2800) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1062 ( .A1(DP_OP_425J2_127_3477_n2868), 
        .A2(DP_OP_423J2_125_3477_n1858), .Y(DP_OP_424J2_126_3477_n1835) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1854 ( .A1(DP_OP_423J2_125_3477_n2731), 
        .A2(DP_OP_424J2_126_3477_n2652), .Y(DP_OP_424J2_126_3477_n2624) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1546 ( .A1(DP_OP_422J2_124_3477_n2518), 
        .A2(n448), .Y(DP_OP_424J2_126_3477_n2319) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2029 ( .A1(DP_OP_424J2_126_3477_n2823), 
        .A2(DP_OP_424J2_126_3477_n2828), .Y(DP_OP_424J2_126_3477_n2799) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2044 ( .A1(DP_OP_424J2_126_3477_n2822), 
        .A2(DP_OP_424J2_126_3477_n2830), .Y(DP_OP_424J2_126_3477_n2814) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1201 ( .A1(DP_OP_423J2_125_3477_n1897), 
        .A2(DP_OP_424J2_126_3477_n1996), .Y(DP_OP_424J2_126_3477_n1974) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1283 ( .A1(DP_OP_422J2_124_3477_n2781), 
        .A2(n447), .Y(DP_OP_424J2_126_3477_n2056) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1547 ( .A1(DP_OP_424J2_126_3477_n2344), 
        .A2(n448), .Y(DP_OP_424J2_126_3477_n2320) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2045 ( .A1(DP_OP_424J2_126_3477_n2823), 
        .A2(DP_OP_424J2_126_3477_n2830), .Y(DP_OP_424J2_126_3477_n2815) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1855 ( .A1(DP_OP_424J2_126_3477_n2649), 
        .A2(DP_OP_424J2_126_3477_n2652), .Y(DP_OP_424J2_126_3477_n2625) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1063 ( .A1(DP_OP_425J2_127_3477_n2869), 
        .A2(DP_OP_423J2_125_3477_n1858), .Y(DP_OP_424J2_126_3477_n1836) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1202 ( .A1(DP_OP_423J2_125_3477_n1898), 
        .A2(DP_OP_424J2_126_3477_n1996), .Y(DP_OP_424J2_126_3477_n1975) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2031 ( .A1(DP_OP_424J2_126_3477_n2825), 
        .A2(DP_OP_424J2_126_3477_n2828), .Y(DP_OP_424J2_126_3477_n2801) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1544 ( .A1(DP_OP_425J2_127_3477_n2341), 
        .A2(DP_OP_425J2_127_3477_n2347), .Y(DP_OP_425J2_127_3477_n2317) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2044 ( .A1(DP_OP_424J2_126_3477_n1901), 
        .A2(DP_OP_425J2_127_3477_n2830), .Y(DP_OP_425J2_127_3477_n2814) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1546 ( .A1(DP_OP_424J2_126_3477_n2428), 
        .A2(DP_OP_425J2_127_3477_n2347), .Y(DP_OP_425J2_127_3477_n2319) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1282 ( .A1(DP_OP_425J2_127_3477_n2079), 
        .A2(DP_OP_425J2_127_3477_n2083), .Y(DP_OP_425J2_127_3477_n2055) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1200 ( .A1(DP_OP_425J2_127_3477_n1989), 
        .A2(DP_OP_422J2_124_3477_n1996), .Y(DP_OP_425J2_127_3477_n1973) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1853 ( .A1(DP_OP_424J2_126_3477_n2078), 
        .A2(DP_OP_425J2_127_3477_n2652), .Y(DP_OP_425J2_127_3477_n2623) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2030 ( .A1(DP_OP_424J2_126_3477_n1903), 
        .A2(DP_OP_425J2_127_3477_n2828), .Y(DP_OP_425J2_127_3477_n2800) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1201 ( .A1(DP_OP_425J2_127_3477_n1990), 
        .A2(DP_OP_424J2_126_3477_n1996), .Y(DP_OP_425J2_127_3477_n1974) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1854 ( .A1(DP_OP_422J2_124_3477_n2780), 
        .A2(DP_OP_425J2_127_3477_n2652), .Y(DP_OP_425J2_127_3477_n2624) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1062 ( .A1(DP_OP_424J2_126_3477_n2912), 
        .A2(DP_OP_425J2_127_3477_n1863), .Y(DP_OP_425J2_127_3477_n1835) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2045 ( .A1(DP_OP_425J2_127_3477_n2823), 
        .A2(DP_OP_425J2_127_3477_n2830), .Y(DP_OP_425J2_127_3477_n2815) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1202 ( .A1(DP_OP_425J2_127_3477_n1991), 
        .A2(DP_OP_424J2_126_3477_n1996), .Y(DP_OP_425J2_127_3477_n1975) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2031 ( .A1(DP_OP_424J2_126_3477_n1904), 
        .A2(DP_OP_425J2_127_3477_n2828), .Y(DP_OP_425J2_127_3477_n2801) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1063 ( .A1(DP_OP_425J2_127_3477_n1860), 
        .A2(DP_OP_425J2_127_3477_n1863), .Y(DP_OP_425J2_127_3477_n1836) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1547 ( .A1(DP_OP_423J2_125_3477_n2515), 
        .A2(DP_OP_425J2_127_3477_n2347), .Y(DP_OP_425J2_127_3477_n2320) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1283 ( .A1(DP_OP_424J2_126_3477_n2693), 
        .A2(DP_OP_425J2_127_3477_n2083), .Y(DP_OP_425J2_127_3477_n2056) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1204 ( .A1(DP_OP_422J2_124_3477_n1861), 
        .A2(DP_OP_423J2_125_3477_n1991), .Y(DP_OP_425J2_127_3477_n1977) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2047 ( .A1(DP_OP_424J2_126_3477_n1904), 
        .A2(DP_OP_425J2_127_3477_n2830), .Y(DP_OP_425J2_127_3477_n2817) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2046 ( .A1(DP_OP_424J2_126_3477_n1903), 
        .A2(DP_OP_425J2_127_3477_n2830), .Y(DP_OP_425J2_127_3477_n2816) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2032 ( .A1(DP_OP_425J2_127_3477_n2826), 
        .A2(DP_OP_425J2_127_3477_n2828), .Y(DP_OP_425J2_127_3477_n2802) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1856 ( .A1(DP_OP_425J2_127_3477_n2650), 
        .A2(DP_OP_425J2_127_3477_n2652), .Y(DP_OP_425J2_127_3477_n2626) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1203 ( .A1(DP_OP_425J2_127_3477_n1992), 
        .A2(DP_OP_423J2_125_3477_n1991), .Y(DP_OP_425J2_127_3477_n1976) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1064 ( .A1(DP_OP_425J2_127_3477_n1861), 
        .A2(DP_OP_425J2_127_3477_n1863), .Y(DP_OP_425J2_127_3477_n1837) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1548 ( .A1(DP_OP_424J2_126_3477_n2430), 
        .A2(DP_OP_425J2_127_3477_n2347), .Y(DP_OP_425J2_127_3477_n2321) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1284 ( .A1(DP_OP_423J2_125_3477_n2777), 
        .A2(DP_OP_425J2_127_3477_n2083), .Y(DP_OP_425J2_127_3477_n2057) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1061 ( .A1(DP_OP_425J2_127_3477_n1858), 
        .A2(DP_OP_425J2_127_3477_n1863), .Y(DP_OP_425J2_127_3477_n1834) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2029 ( .A1(DP_OP_425J2_127_3477_n2823), 
        .A2(DP_OP_425J2_127_3477_n2828), .Y(DP_OP_425J2_127_3477_n2799) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2043 ( .A1(DP_OP_425J2_127_3477_n2821), 
        .A2(DP_OP_425J2_127_3477_n2830), .Y(DP_OP_425J2_127_3477_n2813) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1281 ( .A1(DP_OP_425J2_127_3477_n2078), 
        .A2(DP_OP_425J2_127_3477_n2083), .Y(DP_OP_425J2_127_3477_n2054) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1545 ( .A1(DP_OP_425J2_127_3477_n2342), 
        .A2(DP_OP_425J2_127_3477_n2347), .Y(DP_OP_425J2_127_3477_n2318) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1280 ( .A1(DP_OP_425J2_127_3477_n2077), 
        .A2(DP_OP_425J2_127_3477_n2083), .Y(DP_OP_425J2_127_3477_n2053) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2027 ( .A1(DP_OP_425J2_127_3477_n2821), 
        .A2(DP_OP_425J2_127_3477_n2828), .Y(DP_OP_425J2_127_3477_n2797) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1851 ( .A1(DP_OP_423J2_125_3477_n1983), 
        .A2(DP_OP_425J2_127_3477_n2652), .Y(DP_OP_425J2_127_3477_n2621) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2048 ( .A1(DP_OP_425J2_127_3477_n2826), 
        .A2(DP_OP_425J2_127_3477_n2830), .Y(DP_OP_425J2_127_3477_n2818) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1543 ( .A1(DP_OP_425J2_127_3477_n2340), 
        .A2(DP_OP_425J2_127_3477_n2347), .Y(DP_OP_425J2_127_3477_n2316) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1198 ( .A1(DP_OP_423J2_125_3477_n2859), 
        .A2(DP_OP_422J2_124_3477_n1996), .Y(DP_OP_425J2_127_3477_n1971) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1059 ( .A1(DP_OP_424J2_126_3477_n2909), 
        .A2(DP_OP_425J2_127_3477_n1863), .Y(DP_OP_425J2_127_3477_n1832) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1279 ( .A1(DP_OP_423J2_125_3477_n2772), 
        .A2(DP_OP_425J2_127_3477_n2083), .Y(DP_OP_425J2_127_3477_n2052) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1060 ( .A1(DP_OP_424J2_126_3477_n2910), 
        .A2(DP_OP_425J2_127_3477_n1863), .Y(DP_OP_425J2_127_3477_n1833) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1852 ( .A1(DP_OP_425J2_127_3477_n2646), 
        .A2(DP_OP_425J2_127_3477_n2652), .Y(DP_OP_425J2_127_3477_n2622) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1199 ( .A1(DP_OP_423J2_125_3477_n2860), 
        .A2(DP_OP_423J2_125_3477_n1991), .Y(DP_OP_425J2_127_3477_n1972) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2028 ( .A1(DP_OP_424J2_126_3477_n1901), 
        .A2(DP_OP_425J2_127_3477_n2828), .Y(DP_OP_425J2_127_3477_n2798) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1279 ( .A1(DP_OP_423J2_125_3477_n1983), 
        .A2(DP_OP_422J2_124_3477_n2082), .Y(DP_OP_424J2_126_3477_n2052) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1851 ( .A1(DP_OP_422J2_124_3477_n1988), 
        .A2(DP_OP_424J2_126_3477_n2652), .Y(DP_OP_424J2_126_3477_n2621) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1543 ( .A1(DP_OP_423J2_125_3477_n2247), 
        .A2(n448), .Y(DP_OP_424J2_126_3477_n2316) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2027 ( .A1(DP_OP_424J2_126_3477_n2821), 
        .A2(DP_OP_424J2_126_3477_n2828), .Y(DP_OP_424J2_126_3477_n2797) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1059 ( .A1(DP_OP_425J2_127_3477_n2865), 
        .A2(DP_OP_423J2_125_3477_n1858), .Y(DP_OP_424J2_126_3477_n1832) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1281 ( .A1(DP_OP_424J2_126_3477_n2078), 
        .A2(n447), .Y(DP_OP_424J2_126_3477_n2054) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1853 ( .A1(DP_OP_423J2_125_3477_n2730), 
        .A2(DP_OP_424J2_126_3477_n2652), .Y(DP_OP_424J2_126_3477_n2623) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1061 ( .A1(DP_OP_424J2_126_3477_n1858), 
        .A2(DP_OP_423J2_125_3477_n1858), .Y(DP_OP_424J2_126_3477_n1834) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1545 ( .A1(DP_OP_424J2_126_3477_n2342), 
        .A2(n448), .Y(DP_OP_424J2_126_3477_n2318) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1200 ( .A1(DP_OP_425J2_127_3477_n2734), 
        .A2(DP_OP_424J2_126_3477_n1996), .Y(DP_OP_424J2_126_3477_n1973) );
  XOR2X1_HVT DP_OP_422J2_124_3477_U4 ( .A1(DP_OP_422J2_124_3477_n1773), .A2(
        DP_OP_422J2_124_3477_n153), .Y(DP_OP_422J2_124_3477_n3) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1060 ( .A1(DP_OP_424J2_126_3477_n1857), 
        .A2(DP_OP_422J2_124_3477_n1863), .Y(DP_OP_424J2_126_3477_n1833) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1103 ( .A1(DP_OP_425J2_127_3477_n2821), 
        .A2(DP_OP_424J2_126_3477_n1907), .Y(DP_OP_424J2_126_3477_n1876) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1608 ( .A1(DP_OP_422J2_124_3477_n2388), 
        .A2(DP_OP_422J2_124_3477_n2392), .Y(DP_OP_422J2_124_3477_n2380) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2135 ( .A1(DP_OP_425J2_127_3477_n2913), 
        .A2(DP_OP_425J2_127_3477_n2918), .Y(DP_OP_425J2_127_3477_n2905) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1944 ( .A1(DP_OP_423J2_125_3477_n2731), 
        .A2(DP_OP_422J2_124_3477_n2741), .Y(DP_OP_423J2_125_3477_n2715) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1108 ( .A1(DP_OP_422J2_124_3477_n1905), 
        .A2(DP_OP_422J2_124_3477_n1907), .Y(DP_OP_422J2_124_3477_n1881) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2136 ( .A1(DP_OP_423J2_125_3477_n1856), 
        .A2(DP_OP_422J2_124_3477_n2918), .Y(DP_OP_422J2_124_3477_n2906) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1896 ( .A1(DP_OP_422J2_124_3477_n2692), 
        .A2(DP_OP_422J2_124_3477_n2698), .Y(DP_OP_422J2_124_3477_n2668) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2130 ( .A1(DP_OP_423J2_125_3477_n2909), 
        .A2(DP_OP_423J2_125_3477_n2913), .Y(DP_OP_423J2_125_3477_n2901) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1104 ( .A1(DP_OP_425J2_127_3477_n1901), 
        .A2(DP_OP_425J2_127_3477_n1907), .Y(DP_OP_425J2_127_3477_n1877) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1604 ( .A1(DP_OP_425J2_127_3477_n2382), 
        .A2(DP_OP_424J2_126_3477_n2390), .Y(DP_OP_425J2_127_3477_n2374) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2127 ( .A1(DP_OP_423J2_125_3477_n2906), 
        .A2(DP_OP_423J2_125_3477_n2913), .Y(DP_OP_423J2_125_3477_n2898) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1952 ( .A1(DP_OP_425J2_127_3477_n2738), 
        .A2(DP_OP_425J2_127_3477_n2741), .Y(DP_OP_425J2_127_3477_n2722) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1949 ( .A1(DP_OP_425J2_127_3477_n2735), 
        .A2(DP_OP_425J2_127_3477_n2741), .Y(DP_OP_425J2_127_3477_n2719) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1602 ( .A1(DP_OP_422J2_124_3477_n2344), 
        .A2(DP_OP_423J2_125_3477_n2388), .Y(DP_OP_423J2_125_3477_n2376) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1896 ( .A1(DP_OP_425J2_127_3477_n2690), 
        .A2(DP_OP_425J2_127_3477_n2696), .Y(DP_OP_425J2_127_3477_n2666) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1952 ( .A1(DP_OP_423J2_125_3477_n2032), 
        .A2(DP_OP_422J2_124_3477_n2741), .Y(DP_OP_422J2_124_3477_n2722) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2134 ( .A1(DP_OP_424J2_126_3477_n2912), 
        .A2(DP_OP_422J2_124_3477_n2918), .Y(DP_OP_424J2_126_3477_n2904) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1892 ( .A1(DP_OP_423J2_125_3477_n2690), 
        .A2(DP_OP_425J2_127_3477_n2696), .Y(DP_OP_423J2_125_3477_n2666) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1106 ( .A1(DP_OP_425J2_127_3477_n1903), 
        .A2(DP_OP_425J2_127_3477_n1907), .Y(DP_OP_425J2_127_3477_n1879) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1898 ( .A1(DP_OP_425J2_127_3477_n2692), 
        .A2(DP_OP_425J2_127_3477_n2696), .Y(DP_OP_425J2_127_3477_n2668) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2135 ( .A1(DP_OP_422J2_124_3477_n2913), 
        .A2(DP_OP_422J2_124_3477_n2918), .Y(DP_OP_422J2_124_3477_n2905) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1940 ( .A1(DP_OP_425J2_127_3477_n2119), 
        .A2(DP_OP_424J2_126_3477_n2741), .Y(DP_OP_423J2_125_3477_n2711) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1607 ( .A1(DP_OP_422J2_124_3477_n2387), 
        .A2(DP_OP_422J2_124_3477_n2392), .Y(DP_OP_422J2_124_3477_n2379) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1947 ( .A1(DP_OP_424J2_126_3477_n1988), 
        .A2(DP_OP_425J2_127_3477_n2741), .Y(DP_OP_425J2_127_3477_n2717) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1949 ( .A1(DP_OP_424J2_126_3477_n2735), 
        .A2(DP_OP_424J2_126_3477_n2741), .Y(DP_OP_424J2_126_3477_n2719) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1097 ( .A1(DP_OP_422J2_124_3477_n2865), 
        .A2(DP_OP_424J2_126_3477_n1907), .Y(DP_OP_423J2_125_3477_n1871) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1105 ( .A1(DP_OP_425J2_127_3477_n2823), 
        .A2(DP_OP_424J2_126_3477_n1907), .Y(DP_OP_424J2_126_3477_n1878) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1606 ( .A1(DP_OP_424J2_126_3477_n2384), 
        .A2(DP_OP_424J2_126_3477_n2390), .Y(DP_OP_424J2_126_3477_n2376) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1108 ( .A1(DP_OP_425J2_127_3477_n2826), 
        .A2(DP_OP_424J2_126_3477_n1907), .Y(DP_OP_424J2_126_3477_n1881) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1948 ( .A1(DP_OP_424J2_126_3477_n2734), 
        .A2(DP_OP_424J2_126_3477_n2741), .Y(DP_OP_424J2_126_3477_n2718) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1951 ( .A1(DP_OP_424J2_126_3477_n2737), 
        .A2(DP_OP_424J2_126_3477_n2741), .Y(DP_OP_424J2_126_3477_n2721) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1603 ( .A1(DP_OP_424J2_126_3477_n2381), 
        .A2(DP_OP_424J2_126_3477_n2390), .Y(DP_OP_424J2_126_3477_n2373) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1897 ( .A1(DP_OP_424J2_126_3477_n2691), 
        .A2(DP_OP_424J2_126_3477_n2696), .Y(DP_OP_424J2_126_3477_n2667) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1898 ( .A1(DP_OP_425J2_127_3477_n2079), 
        .A2(DP_OP_424J2_126_3477_n2696), .Y(DP_OP_424J2_126_3477_n2668) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2131 ( .A1(DP_OP_424J2_126_3477_n2909), 
        .A2(DP_OP_425J2_127_3477_n2918), .Y(DP_OP_424J2_126_3477_n2901) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1605 ( .A1(DP_OP_424J2_126_3477_n2383), 
        .A2(DP_OP_424J2_126_3477_n2390), .Y(DP_OP_424J2_126_3477_n2375) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1107 ( .A1(DP_OP_424J2_126_3477_n1904), 
        .A2(DP_OP_424J2_126_3477_n1907), .Y(DP_OP_424J2_126_3477_n1880) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1605 ( .A1(DP_OP_425J2_127_3477_n2383), 
        .A2(DP_OP_423J2_125_3477_n2388), .Y(DP_OP_425J2_127_3477_n2375) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1950 ( .A1(DP_OP_422J2_124_3477_n2868), 
        .A2(DP_OP_425J2_127_3477_n2741), .Y(DP_OP_425J2_127_3477_n2720) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1602 ( .A1(DP_OP_422J2_124_3477_n2382), 
        .A2(DP_OP_422J2_124_3477_n2392), .Y(DP_OP_422J2_124_3477_n2374) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1898 ( .A1(DP_OP_422J2_124_3477_n2694), 
        .A2(DP_OP_422J2_124_3477_n2698), .Y(DP_OP_422J2_124_3477_n2670) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1106 ( .A1(DP_OP_422J2_124_3477_n1903), 
        .A2(DP_OP_422J2_124_3477_n1907), .Y(DP_OP_422J2_124_3477_n1879) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1600 ( .A1(DP_OP_422J2_124_3477_n2342), 
        .A2(DP_OP_423J2_125_3477_n2388), .Y(DP_OP_423J2_125_3477_n2374) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1899 ( .A1(DP_OP_424J2_126_3477_n2693), 
        .A2(DP_OP_424J2_126_3477_n2696), .Y(DP_OP_424J2_126_3477_n2669) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1895 ( .A1(DP_OP_424J2_126_3477_n2689), 
        .A2(DP_OP_424J2_126_3477_n2696), .Y(DP_OP_424J2_126_3477_n2665) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2133 ( .A1(DP_OP_425J2_127_3477_n2911), 
        .A2(DP_OP_425J2_127_3477_n2918), .Y(DP_OP_425J2_127_3477_n2903) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1949 ( .A1(DP_OP_422J2_124_3477_n2735), 
        .A2(DP_OP_422J2_124_3477_n2741), .Y(DP_OP_422J2_124_3477_n2719) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1596 ( .A1(DP_OP_422J2_124_3477_n2338), 
        .A2(DP_OP_423J2_125_3477_n2388), .Y(DP_OP_423J2_125_3477_n2370) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1107 ( .A1(DP_OP_424J2_126_3477_n2869), 
        .A2(DP_OP_425J2_127_3477_n1907), .Y(DP_OP_425J2_127_3477_n1880) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2133 ( .A1(DP_OP_425J2_127_3477_n1858), 
        .A2(DP_OP_422J2_124_3477_n2918), .Y(DP_OP_424J2_126_3477_n2903) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1900 ( .A1(DP_OP_422J2_124_3477_n2696), 
        .A2(DP_OP_422J2_124_3477_n2698), .Y(DP_OP_422J2_124_3477_n2672) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2132 ( .A1(DP_OP_425J2_127_3477_n2778), 
        .A2(DP_OP_422J2_124_3477_n2918), .Y(DP_OP_422J2_124_3477_n2902) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1890 ( .A1(DP_OP_423J2_125_3477_n2688), 
        .A2(DP_OP_424J2_126_3477_n2696), .Y(DP_OP_423J2_125_3477_n2664) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1098 ( .A1(DP_OP_423J2_125_3477_n1896), 
        .A2(DP_OP_424J2_126_3477_n1907), .Y(DP_OP_423J2_125_3477_n1872) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1102 ( .A1(DP_OP_425J2_127_3477_n2738), 
        .A2(DP_OP_422J2_124_3477_n1907), .Y(DP_OP_423J2_125_3477_n1876) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1604 ( .A1(DP_OP_422J2_124_3477_n2384), 
        .A2(DP_OP_422J2_124_3477_n2392), .Y(DP_OP_422J2_124_3477_n2376) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1606 ( .A1(DP_OP_422J2_124_3477_n2386), 
        .A2(DP_OP_422J2_124_3477_n2392), .Y(DP_OP_422J2_124_3477_n2378) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2128 ( .A1(DP_OP_423J2_125_3477_n2907), 
        .A2(DP_OP_423J2_125_3477_n2913), .Y(DP_OP_423J2_125_3477_n2899) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2132 ( .A1(DP_OP_425J2_127_3477_n2910), 
        .A2(DP_OP_425J2_127_3477_n2918), .Y(DP_OP_425J2_127_3477_n2902) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2134 ( .A1(DP_OP_422J2_124_3477_n2912), 
        .A2(DP_OP_422J2_124_3477_n2918), .Y(DP_OP_422J2_124_3477_n2904) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1601 ( .A1(DP_OP_422J2_124_3477_n2343), 
        .A2(DP_OP_423J2_125_3477_n2388), .Y(DP_OP_423J2_125_3477_n2375) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1951 ( .A1(DP_OP_423J2_125_3477_n2031), 
        .A2(DP_OP_422J2_124_3477_n2741), .Y(DP_OP_422J2_124_3477_n2721) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1894 ( .A1(DP_OP_425J2_127_3477_n2169), 
        .A2(DP_OP_425J2_127_3477_n2696), .Y(DP_OP_423J2_125_3477_n2668) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2136 ( .A1(DP_OP_425J2_127_3477_n1861), 
        .A2(DP_OP_422J2_124_3477_n2918), .Y(DP_OP_424J2_126_3477_n2906) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1608 ( .A1(DP_OP_424J2_126_3477_n2386), 
        .A2(DP_OP_424J2_126_3477_n2390), .Y(DP_OP_424J2_126_3477_n2378) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1950 ( .A1(DP_OP_424J2_126_3477_n2736), 
        .A2(DP_OP_424J2_126_3477_n2741), .Y(DP_OP_424J2_126_3477_n2720) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1893 ( .A1(DP_OP_425J2_127_3477_n2168), 
        .A2(DP_OP_424J2_126_3477_n2696), .Y(DP_OP_423J2_125_3477_n2667) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1599 ( .A1(DP_OP_422J2_124_3477_n2341), 
        .A2(DP_OP_423J2_125_3477_n2388), .Y(DP_OP_423J2_125_3477_n2373) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1106 ( .A1(DP_OP_424J2_126_3477_n1903), 
        .A2(DP_OP_424J2_126_3477_n1907), .Y(DP_OP_424J2_126_3477_n1879) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1945 ( .A1(DP_OP_423J2_125_3477_n2732), 
        .A2(DP_OP_424J2_126_3477_n2741), .Y(DP_OP_423J2_125_3477_n2716) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1946 ( .A1(DP_OP_423J2_125_3477_n2733), 
        .A2(DP_OP_425J2_127_3477_n2741), .Y(DP_OP_423J2_125_3477_n2717) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1899 ( .A1(DP_OP_423J2_125_3477_n1943), 
        .A2(DP_OP_425J2_127_3477_n2696), .Y(DP_OP_425J2_127_3477_n2669) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1101 ( .A1(DP_OP_423J2_125_3477_n1899), 
        .A2(DP_OP_422J2_124_3477_n1907), .Y(DP_OP_423J2_125_3477_n1875) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2136 ( .A1(DP_OP_425J2_127_3477_n2914), 
        .A2(DP_OP_425J2_127_3477_n2918), .Y(DP_OP_425J2_127_3477_n2906) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2131 ( .A1(DP_OP_425J2_127_3477_n2909), 
        .A2(DP_OP_425J2_127_3477_n2918), .Y(DP_OP_425J2_127_3477_n2901) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2131 ( .A1(DP_OP_422J2_124_3477_n2909), 
        .A2(DP_OP_422J2_124_3477_n2918), .Y(DP_OP_422J2_124_3477_n2901) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1900 ( .A1(DP_OP_425J2_127_3477_n2694), 
        .A2(DP_OP_425J2_127_3477_n2696), .Y(DP_OP_425J2_127_3477_n2670) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1105 ( .A1(DP_OP_422J2_124_3477_n1902), 
        .A2(DP_OP_422J2_124_3477_n1907), .Y(DP_OP_422J2_124_3477_n1878) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2133 ( .A1(DP_OP_423J2_125_3477_n1853), 
        .A2(DP_OP_422J2_124_3477_n2918), .Y(DP_OP_422J2_124_3477_n2903) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1103 ( .A1(DP_OP_422J2_124_3477_n1900), 
        .A2(DP_OP_422J2_124_3477_n1907), .Y(DP_OP_422J2_124_3477_n1876) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1605 ( .A1(DP_OP_422J2_124_3477_n2385), 
        .A2(DP_OP_422J2_124_3477_n2392), .Y(DP_OP_422J2_124_3477_n2377) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1896 ( .A1(DP_OP_422J2_124_3477_n1945), 
        .A2(DP_OP_424J2_126_3477_n2696), .Y(DP_OP_424J2_126_3477_n2666) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1104 ( .A1(DP_OP_424J2_126_3477_n2734), 
        .A2(DP_OP_422J2_124_3477_n1907), .Y(DP_OP_422J2_124_3477_n1877) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1943 ( .A1(DP_OP_423J2_125_3477_n2730), 
        .A2(DP_OP_425J2_127_3477_n2741), .Y(DP_OP_423J2_125_3477_n2714) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2129 ( .A1(DP_OP_423J2_125_3477_n2908), 
        .A2(DP_OP_423J2_125_3477_n2913), .Y(DP_OP_423J2_125_3477_n2900) );
  XOR2X1_HVT DP_OP_425J2_127_3477_U4 ( .A1(DP_OP_425J2_127_3477_n1773), .A2(
        DP_OP_425J2_127_3477_n153), .Y(DP_OP_425J2_127_3477_n3) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1891 ( .A1(DP_OP_425J2_127_3477_n2166), 
        .A2(DP_OP_425J2_127_3477_n2696), .Y(DP_OP_423J2_125_3477_n2665) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1099 ( .A1(DP_OP_423J2_125_3477_n1897), 
        .A2(DP_OP_425J2_127_3477_n1907), .Y(DP_OP_423J2_125_3477_n1873) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1950 ( .A1(DP_OP_422J2_124_3477_n2736), 
        .A2(DP_OP_422J2_124_3477_n2741), .Y(DP_OP_422J2_124_3477_n2720) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1897 ( .A1(DP_OP_425J2_127_3477_n2691), 
        .A2(DP_OP_425J2_127_3477_n2696), .Y(DP_OP_425J2_127_3477_n2667) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1105 ( .A1(DP_OP_424J2_126_3477_n2867), 
        .A2(DP_OP_425J2_127_3477_n1907), .Y(DP_OP_425J2_127_3477_n1878) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1947 ( .A1(DP_OP_424J2_126_3477_n2733), 
        .A2(DP_OP_424J2_126_3477_n2741), .Y(DP_OP_424J2_126_3477_n2717) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1107 ( .A1(DP_OP_422J2_124_3477_n1904), 
        .A2(DP_OP_422J2_124_3477_n1907), .Y(DP_OP_422J2_124_3477_n1880) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1608 ( .A1(DP_OP_425J2_127_3477_n2386), 
        .A2(DP_OP_422J2_124_3477_n2392), .Y(DP_OP_425J2_127_3477_n2378) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1103 ( .A1(DP_OP_424J2_126_3477_n2865), 
        .A2(DP_OP_425J2_127_3477_n1907), .Y(DP_OP_425J2_127_3477_n1876) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2135 ( .A1(DP_OP_425J2_127_3477_n1860), 
        .A2(DP_OP_423J2_125_3477_n2913), .Y(DP_OP_424J2_126_3477_n2905) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1606 ( .A1(DP_OP_425J2_127_3477_n2384), 
        .A2(DP_OP_423J2_125_3477_n2388), .Y(DP_OP_425J2_127_3477_n2376) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1900 ( .A1(DP_OP_423J2_125_3477_n2777), 
        .A2(DP_OP_424J2_126_3477_n2696), .Y(DP_OP_424J2_126_3477_n2670) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2134 ( .A1(DP_OP_425J2_127_3477_n2912), 
        .A2(DP_OP_425J2_127_3477_n2918), .Y(DP_OP_425J2_127_3477_n2904) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1100 ( .A1(DP_OP_423J2_125_3477_n1898), 
        .A2(DP_OP_425J2_127_3477_n1907), .Y(DP_OP_423J2_125_3477_n1874) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2132 ( .A1(DP_OP_424J2_126_3477_n2910), 
        .A2(DP_OP_423J2_125_3477_n2913), .Y(DP_OP_424J2_126_3477_n2902) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1951 ( .A1(DP_OP_423J2_125_3477_n1899), 
        .A2(DP_OP_425J2_127_3477_n2741), .Y(DP_OP_425J2_127_3477_n2721) );
  OR2X1_HVT DP_OP_425J2_127_3477_U33 ( .A1(DP_OP_425J2_127_3477_n179), .A2(
        DP_OP_425J2_127_3477_n178), .Y(DP_OP_425J2_127_3477_n45) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1895 ( .A1(DP_OP_425J2_127_3477_n2557), 
        .A2(DP_OP_422J2_124_3477_n2698), .Y(DP_OP_422J2_124_3477_n2667) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1104 ( .A1(DP_OP_424J2_126_3477_n1901), 
        .A2(DP_OP_424J2_126_3477_n1907), .Y(DP_OP_424J2_126_3477_n1877) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1604 ( .A1(DP_OP_424J2_126_3477_n2382), 
        .A2(DP_OP_424J2_126_3477_n2390), .Y(DP_OP_424J2_126_3477_n2374) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1889 ( .A1(DP_OP_425J2_127_3477_n2164), 
        .A2(DP_OP_424J2_126_3477_n2696), .Y(DP_OP_423J2_125_3477_n2663) );
  XOR2X1_HVT DP_OP_424J2_126_3477_U4 ( .A1(DP_OP_424J2_126_3477_n1773), .A2(
        DP_OP_424J2_126_3477_n153), .Y(DP_OP_424J2_126_3477_n3) );
  XOR2X1_HVT DP_OP_423J2_125_3477_U4 ( .A1(DP_OP_423J2_125_3477_n1768), .A2(
        DP_OP_423J2_125_3477_n148), .Y(DP_OP_423J2_125_3477_n3) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1899 ( .A1(DP_OP_422J2_124_3477_n2695), 
        .A2(DP_OP_422J2_124_3477_n2698), .Y(DP_OP_422J2_124_3477_n2671) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1598 ( .A1(DP_OP_422J2_124_3477_n2340), 
        .A2(DP_OP_423J2_125_3477_n2388), .Y(DP_OP_423J2_125_3477_n2372) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1897 ( .A1(DP_OP_425J2_127_3477_n2559), 
        .A2(DP_OP_422J2_124_3477_n2698), .Y(DP_OP_422J2_124_3477_n2669) );
  OR2X1_HVT DP_OP_422J2_124_3477_U33 ( .A1(DP_OP_422J2_124_3477_n179), .A2(
        DP_OP_422J2_124_3477_n178), .Y(DP_OP_422J2_124_3477_n45) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1597 ( .A1(DP_OP_422J2_124_3477_n2339), 
        .A2(DP_OP_423J2_125_3477_n2388), .Y(DP_OP_423J2_125_3477_n2371) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1895 ( .A1(DP_OP_423J2_125_3477_n1939), 
        .A2(DP_OP_425J2_127_3477_n2696), .Y(DP_OP_425J2_127_3477_n2665) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2126 ( .A1(DP_OP_425J2_127_3477_n1945), 
        .A2(DP_OP_423J2_125_3477_n2913), .Y(DP_OP_423J2_125_3477_n2897) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1603 ( .A1(DP_OP_422J2_124_3477_n2383), 
        .A2(DP_OP_422J2_124_3477_n2392), .Y(DP_OP_422J2_124_3477_n2375) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1948 ( .A1(DP_OP_425J2_127_3477_n2734), 
        .A2(DP_OP_425J2_127_3477_n2741), .Y(DP_OP_425J2_127_3477_n2718) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1948 ( .A1(DP_OP_422J2_124_3477_n2734), 
        .A2(DP_OP_422J2_124_3477_n2741), .Y(DP_OP_422J2_124_3477_n2718) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1108 ( .A1(DP_OP_425J2_127_3477_n1905), 
        .A2(DP_OP_425J2_127_3477_n1907), .Y(DP_OP_425J2_127_3477_n1881) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1952 ( .A1(DP_OP_424J2_126_3477_n2738), 
        .A2(DP_OP_424J2_126_3477_n2741), .Y(DP_OP_424J2_126_3477_n2722) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1607 ( .A1(DP_OP_424J2_126_3477_n2344), 
        .A2(DP_OP_423J2_125_3477_n2388), .Y(DP_OP_425J2_127_3477_n2377) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1942 ( .A1(DP_OP_423J2_125_3477_n2729), 
        .A2(DP_OP_422J2_124_3477_n2741), .Y(DP_OP_423J2_125_3477_n2713) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1607 ( .A1(DP_OP_424J2_126_3477_n2385), 
        .A2(DP_OP_424J2_126_3477_n2390), .Y(DP_OP_424J2_126_3477_n2377) );
  OR2X1_HVT DP_OP_422J2_124_3477_U162 ( .A1(DP_OP_422J2_124_3477_n1584), .A2(
        DP_OP_422J2_124_3477_n1582), .Y(DP_OP_422J2_124_3477_n126) );
  OR2X1_HVT DP_OP_423J2_125_3477_U162 ( .A1(DP_OP_423J2_125_3477_n1579), .A2(
        DP_OP_423J2_125_3477_n1577), .Y(DP_OP_423J2_125_3477_n124) );
  OR2X1_HVT DP_OP_425J2_127_3477_U162 ( .A1(DP_OP_425J2_127_3477_n1584), .A2(
        DP_OP_425J2_127_3477_n1582), .Y(DP_OP_425J2_127_3477_n126) );
  OR2X1_HVT DP_OP_424J2_126_3477_U162 ( .A1(DP_OP_424J2_126_3477_n1584), .A2(
        DP_OP_424J2_126_3477_n1582), .Y(DP_OP_424J2_126_3477_n126) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U165 ( .A1(DP_OP_424J2_126_3477_n4), .A2(
        DP_OP_424J2_126_3477_n129), .A3(DP_OP_424J2_126_3477_n130), .Y(
        DP_OP_424J2_126_3477_n128) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U165 ( .A1(DP_OP_422J2_124_3477_n4), .A2(
        DP_OP_422J2_124_3477_n129), .A3(DP_OP_422J2_124_3477_n130), .Y(
        DP_OP_422J2_124_3477_n128) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U165 ( .A1(DP_OP_425J2_127_3477_n4), .A2(
        DP_OP_425J2_127_3477_n129), .A3(DP_OP_425J2_127_3477_n130), .Y(
        DP_OP_425J2_127_3477_n128) );
  OR2X1_HVT DP_OP_423J2_125_3477_U148 ( .A1(DP_OP_423J2_125_3477_n1249), .A2(
        DP_OP_423J2_125_3477_n1247), .Y(DP_OP_423J2_125_3477_n116) );
  OR2X1_HVT DP_OP_422J2_124_3477_U148 ( .A1(DP_OP_422J2_124_3477_n1254), .A2(
        DP_OP_422J2_124_3477_n1252), .Y(DP_OP_422J2_124_3477_n118) );
  OR2X1_HVT DP_OP_424J2_126_3477_U148 ( .A1(DP_OP_424J2_126_3477_n1254), .A2(
        DP_OP_424J2_126_3477_n1252), .Y(DP_OP_424J2_126_3477_n118) );
  OR2X1_HVT DP_OP_425J2_127_3477_U148 ( .A1(DP_OP_425J2_127_3477_n1254), .A2(
        DP_OP_425J2_127_3477_n1252), .Y(DP_OP_425J2_127_3477_n118) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U151 ( .A1(DP_OP_424J2_126_3477_n123), .A2(
        DP_OP_424J2_126_3477_n121), .A3(DP_OP_424J2_126_3477_n122), .Y(
        DP_OP_424J2_126_3477_n120) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U151 ( .A1(DP_OP_422J2_124_3477_n123), .A2(
        DP_OP_422J2_124_3477_n121), .A3(DP_OP_422J2_124_3477_n122), .Y(
        DP_OP_422J2_124_3477_n120) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U151 ( .A1(DP_OP_425J2_127_3477_n123), .A2(
        DP_OP_425J2_127_3477_n121), .A3(DP_OP_425J2_127_3477_n122), .Y(
        DP_OP_425J2_127_3477_n120) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U151 ( .A1(DP_OP_423J2_125_3477_n121), .A2(
        DP_OP_423J2_125_3477_n119), .A3(DP_OP_423J2_125_3477_n120), .Y(
        DP_OP_423J2_125_3477_n118) );
  OR2X1_HVT DP_OP_423J2_125_3477_U134 ( .A1(DP_OP_423J2_125_3477_n867), .A2(
        DP_OP_423J2_125_3477_n865), .Y(DP_OP_423J2_125_3477_n108) );
  OR2X1_HVT DP_OP_425J2_127_3477_U134 ( .A1(DP_OP_425J2_127_3477_n872), .A2(
        DP_OP_425J2_127_3477_n870), .Y(DP_OP_425J2_127_3477_n110) );
  OR2X1_HVT DP_OP_422J2_124_3477_U134 ( .A1(DP_OP_422J2_124_3477_n872), .A2(
        DP_OP_422J2_124_3477_n870), .Y(DP_OP_422J2_124_3477_n110) );
  OR2X1_HVT DP_OP_424J2_126_3477_U134 ( .A1(DP_OP_424J2_126_3477_n872), .A2(
        DP_OP_424J2_126_3477_n870), .Y(DP_OP_424J2_126_3477_n110) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U137 ( .A1(DP_OP_423J2_125_3477_n113), .A2(
        DP_OP_423J2_125_3477_n111), .A3(DP_OP_423J2_125_3477_n112), .Y(
        DP_OP_423J2_125_3477_n110) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U137 ( .A1(DP_OP_425J2_127_3477_n115), .A2(
        DP_OP_425J2_127_3477_n113), .A3(DP_OP_425J2_127_3477_n114), .Y(
        DP_OP_425J2_127_3477_n112) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U137 ( .A1(DP_OP_424J2_126_3477_n115), .A2(
        DP_OP_424J2_126_3477_n113), .A3(DP_OP_424J2_126_3477_n114), .Y(
        DP_OP_424J2_126_3477_n112) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U137 ( .A1(DP_OP_422J2_124_3477_n115), .A2(
        DP_OP_422J2_124_3477_n113), .A3(DP_OP_422J2_124_3477_n114), .Y(
        DP_OP_422J2_124_3477_n112) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U71 ( .A1(DP_OP_422J2_124_3477_n186), .A2(
        DP_OP_422J2_124_3477_n191), .Y(DP_OP_422J2_124_3477_n67) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U71 ( .A1(DP_OP_424J2_126_3477_n186), .A2(
        DP_OP_424J2_126_3477_n191), .Y(DP_OP_424J2_126_3477_n67) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U79 ( .A1(DP_OP_422J2_124_3477_n79), .A2(
        DP_OP_422J2_124_3477_n83), .A3(DP_OP_422J2_124_3477_n80), .Y(
        DP_OP_422J2_124_3477_n78) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U123 ( .A1(DP_OP_423J2_125_3477_n103), .A2(
        DP_OP_423J2_125_3477_n105), .A3(DP_OP_423J2_125_3477_n104), .Y(
        DP_OP_423J2_125_3477_n102) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U123 ( .A1(DP_OP_424J2_126_3477_n105), .A2(
        DP_OP_424J2_126_3477_n107), .A3(DP_OP_424J2_126_3477_n106), .Y(
        DP_OP_424J2_126_3477_n104) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U123 ( .A1(DP_OP_425J2_127_3477_n105), .A2(
        DP_OP_425J2_127_3477_n107), .A3(DP_OP_425J2_127_3477_n106), .Y(
        DP_OP_425J2_127_3477_n104) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U93 ( .A1(DP_OP_422J2_124_3477_n93), .A2(
        DP_OP_422J2_124_3477_n87), .A3(DP_OP_422J2_124_3477_n88), .Y(
        DP_OP_422J2_124_3477_n86) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U93 ( .A1(DP_OP_424J2_126_3477_n93), .A2(
        DP_OP_424J2_126_3477_n87), .A3(DP_OP_424J2_126_3477_n88), .Y(
        DP_OP_424J2_126_3477_n86) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U123 ( .A1(DP_OP_422J2_124_3477_n105), .A2(
        DP_OP_422J2_124_3477_n107), .A3(DP_OP_422J2_124_3477_n106), .Y(
        DP_OP_422J2_124_3477_n104) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U93 ( .A1(DP_OP_423J2_125_3477_n91), .A2(
        DP_OP_423J2_125_3477_n85), .A3(DP_OP_423J2_125_3477_n86), .Y(
        DP_OP_423J2_125_3477_n84) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U79 ( .A1(DP_OP_424J2_126_3477_n79), .A2(
        DP_OP_424J2_126_3477_n83), .A3(DP_OP_424J2_126_3477_n80), .Y(
        DP_OP_424J2_126_3477_n78) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U79 ( .A1(DP_OP_423J2_125_3477_n77), .A2(
        DP_OP_423J2_125_3477_n81), .A3(DP_OP_423J2_125_3477_n78), .Y(
        DP_OP_423J2_125_3477_n76) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U79 ( .A1(DP_OP_425J2_127_3477_n79), .A2(
        DP_OP_425J2_127_3477_n83), .A3(DP_OP_425J2_127_3477_n80), .Y(
        DP_OP_425J2_127_3477_n78) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U93 ( .A1(DP_OP_425J2_127_3477_n93), .A2(
        DP_OP_425J2_127_3477_n87), .A3(DP_OP_425J2_127_3477_n88), .Y(
        DP_OP_425J2_127_3477_n86) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U40 ( .A1(DP_OP_424J2_126_3477_n52), .A2(
        DP_OP_424J2_126_3477_n56), .A3(DP_OP_424J2_126_3477_n53), .Y(
        DP_OP_424J2_126_3477_n51) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U75 ( .A1(DP_OP_422J2_124_3477_n75), .A2(
        DP_OP_422J2_124_3477_n95), .A3(DP_OP_422J2_124_3477_n76), .Y(
        DP_OP_422J2_124_3477_n74) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U75 ( .A1(DP_OP_424J2_126_3477_n75), .A2(
        DP_OP_424J2_126_3477_n95), .A3(DP_OP_424J2_126_3477_n76), .Y(
        DP_OP_424J2_126_3477_n74) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U40 ( .A1(DP_OP_425J2_127_3477_n52), .A2(
        DP_OP_425J2_127_3477_n56), .A3(DP_OP_425J2_127_3477_n53), .Y(
        DP_OP_425J2_127_3477_n51) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U40 ( .A1(DP_OP_423J2_125_3477_n50), .A2(
        DP_OP_423J2_125_3477_n54), .A3(DP_OP_423J2_125_3477_n51), .Y(
        DP_OP_423J2_125_3477_n49) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U40 ( .A1(DP_OP_422J2_124_3477_n52), .A2(
        DP_OP_422J2_124_3477_n56), .A3(DP_OP_422J2_124_3477_n53), .Y(
        DP_OP_422J2_124_3477_n51) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U75 ( .A1(DP_OP_423J2_125_3477_n73), .A2(
        DP_OP_423J2_125_3477_n93), .A3(DP_OP_423J2_125_3477_n74), .Y(
        DP_OP_423J2_125_3477_n72) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U75 ( .A1(DP_OP_425J2_127_3477_n75), .A2(
        DP_OP_425J2_127_3477_n95), .A3(DP_OP_425J2_127_3477_n76), .Y(
        DP_OP_425J2_127_3477_n74) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U64 ( .A1(DP_OP_424J2_126_3477_n67), .A2(
        DP_OP_424J2_126_3477_n73), .A3(DP_OP_424J2_126_3477_n68), .Y(
        DP_OP_424J2_126_3477_n66) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U20 ( .A1(DP_OP_422J2_124_3477_n38), .A2(
        DP_OP_422J2_124_3477_n42), .A3(DP_OP_422J2_124_3477_n39), .Y(
        DP_OP_422J2_124_3477_n37) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U64 ( .A1(DP_OP_422J2_124_3477_n67), .A2(
        DP_OP_422J2_124_3477_n73), .A3(DP_OP_422J2_124_3477_n68), .Y(
        DP_OP_422J2_124_3477_n66) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U20 ( .A1(DP_OP_424J2_126_3477_n38), .A2(
        DP_OP_424J2_126_3477_n42), .A3(DP_OP_424J2_126_3477_n39), .Y(
        DP_OP_424J2_126_3477_n37) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U64 ( .A1(DP_OP_423J2_125_3477_n65), .A2(
        DP_OP_423J2_125_3477_n71), .A3(DP_OP_423J2_125_3477_n66), .Y(
        DP_OP_423J2_125_3477_n64) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U20 ( .A1(DP_OP_423J2_125_3477_n36), .A2(
        DP_OP_423J2_125_3477_n40), .A3(DP_OP_423J2_125_3477_n37), .Y(
        DP_OP_423J2_125_3477_n35) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U20 ( .A1(DP_OP_425J2_127_3477_n38), .A2(
        DP_OP_425J2_127_3477_n42), .A3(DP_OP_425J2_127_3477_n39), .Y(
        DP_OP_425J2_127_3477_n37) );
  AO21X1_HVT DP_OP_425J2_127_3477_U18 ( .A1(DP_OP_425J2_127_3477_n74), .A2(
        DP_OP_425J2_127_3477_n36), .A3(DP_OP_425J2_127_3477_n37), .Y(
        DP_OP_425J2_127_3477_n35) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U64 ( .A1(DP_OP_425J2_127_3477_n67), .A2(
        DP_OP_425J2_127_3477_n73), .A3(DP_OP_425J2_127_3477_n68), .Y(
        DP_OP_425J2_127_3477_n66) );
  AO21X1_HVT DP_OP_424J2_126_3477_U18 ( .A1(DP_OP_424J2_126_3477_n74), .A2(
        DP_OP_424J2_126_3477_n36), .A3(DP_OP_424J2_126_3477_n37), .Y(
        DP_OP_424J2_126_3477_n35) );
  AO21X1_HVT DP_OP_422J2_124_3477_U18 ( .A1(DP_OP_422J2_124_3477_n74), .A2(
        DP_OP_422J2_124_3477_n36), .A3(DP_OP_422J2_124_3477_n37), .Y(
        DP_OP_422J2_124_3477_n35) );
  AO21X1_HVT DP_OP_423J2_125_3477_U18 ( .A1(DP_OP_423J2_125_3477_n72), .A2(
        DP_OP_423J2_125_3477_n34), .A3(DP_OP_423J2_125_3477_n35), .Y(
        DP_OP_423J2_125_3477_n33) );
  XOR2X1_HVT DP_OP_422J2_124_3477_U3 ( .A1(DP_OP_422J2_124_3477_n24), .A2(
        DP_OP_422J2_124_3477_n3), .Y(n_conv2_sum_a[31]) );
  XOR2X1_HVT DP_OP_423J2_125_3477_U3 ( .A1(DP_OP_423J2_125_3477_n22), .A2(
        DP_OP_423J2_125_3477_n3), .Y(n_conv2_sum_b[31]) );
  XOR2X1_HVT DP_OP_425J2_127_3477_U3 ( .A1(DP_OP_425J2_127_3477_n24), .A2(
        DP_OP_425J2_127_3477_n3), .Y(n_conv2_sum_d[31]) );
  XOR2X1_HVT DP_OP_424J2_126_3477_U3 ( .A1(DP_OP_424J2_126_3477_n24), .A2(
        DP_OP_424J2_126_3477_n3), .Y(n_conv2_sum_c[31]) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1075 ( .A1(DP_OP_425J2_127_3477_n2865), 
        .A2(DP_OP_424J2_126_3477_n1865), .Y(DP_OP_424J2_126_3477_n1848) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1823 ( .A1(DP_OP_422J2_124_3477_n2031), 
        .A2(DP_OP_424J2_126_3477_n2610), .Y(DP_OP_424J2_126_3477_n2593) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1163 ( .A1(DP_OP_422J2_124_3477_n2909), 
        .A2(DP_OP_424J2_126_3477_n1953), .Y(DP_OP_424J2_126_3477_n1936) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1647 ( .A1(DP_OP_422J2_124_3477_n2427), 
        .A2(DP_OP_422J2_124_3477_n2436), .Y(DP_OP_422J2_124_3477_n2419) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1559 ( .A1(DP_OP_423J2_125_3477_n2247), 
        .A2(DP_OP_424J2_126_3477_n2349), .Y(DP_OP_424J2_126_3477_n2332) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1002 ( .A1(n399), .A2(n337), .Y(
        DP_OP_422J2_124_3477_n1775) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1383 ( .A1(DP_OP_424J2_126_3477_n2164), 
        .A2(DP_OP_424J2_126_3477_n2173), .Y(DP_OP_424J2_126_3477_n2156) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1427 ( .A1(DP_OP_422J2_124_3477_n2207), 
        .A2(DP_OP_422J2_124_3477_n2216), .Y(DP_OP_422J2_124_3477_n2199) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1647 ( .A1(DP_OP_422J2_124_3477_n2207), 
        .A2(DP_OP_423J2_125_3477_n2432), .Y(DP_OP_424J2_126_3477_n2417) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1779 ( .A1(DP_OP_424J2_126_3477_n2557), 
        .A2(DP_OP_424J2_126_3477_n2566), .Y(DP_OP_424J2_126_3477_n2549) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1427 ( .A1(DP_OP_422J2_124_3477_n2647), 
        .A2(DP_OP_422J2_124_3477_n2216), .Y(DP_OP_424J2_126_3477_n2200) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1691 ( .A1(DP_OP_423J2_125_3477_n2291), 
        .A2(DP_OP_422J2_124_3477_n2480), .Y(DP_OP_422J2_124_3477_n2463) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1685 ( .A1(DP_OP_423J2_125_3477_n2467), 
        .A2(DP_OP_423J2_125_3477_n2476), .Y(DP_OP_423J2_125_3477_n2459) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1818 ( .A1(DP_OP_423J2_125_3477_n2600), 
        .A2(DP_OP_425J2_127_3477_n2610), .Y(DP_OP_423J2_125_3477_n2592) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1554 ( .A1(DP_OP_422J2_124_3477_n2428), 
        .A2(DP_OP_423J2_125_3477_n2344), .Y(DP_OP_423J2_125_3477_n2328) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1641 ( .A1(DP_OP_422J2_124_3477_n2295), 
        .A2(DP_OP_423J2_125_3477_n2432), .Y(DP_OP_423J2_125_3477_n2415) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1560 ( .A1(DP_OP_422J2_124_3477_n2340), 
        .A2(DP_OP_425J2_127_3477_n2349), .Y(DP_OP_422J2_124_3477_n2332) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1340 ( .A1(DP_OP_422J2_124_3477_n2120), 
        .A2(DP_OP_422J2_124_3477_n2128), .Y(DP_OP_422J2_124_3477_n2112) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1780 ( .A1(DP_OP_425J2_127_3477_n2558), 
        .A2(DP_OP_425J2_127_3477_n2566), .Y(DP_OP_425J2_127_3477_n2550) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1560 ( .A1(DP_OP_425J2_127_3477_n2341), 
        .A2(DP_OP_425J2_127_3477_n2349), .Y(DP_OP_425J2_127_3477_n2333) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1164 ( .A1(DP_OP_422J2_124_3477_n1945), 
        .A2(DP_OP_423J2_125_3477_n1948), .Y(DP_OP_422J2_124_3477_n1937) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1861 ( .A1(DP_OP_423J2_125_3477_n2643), 
        .A2(DP_OP_424J2_126_3477_n2654), .Y(DP_OP_423J2_125_3477_n2635) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1773 ( .A1(DP_OP_422J2_124_3477_n2163), 
        .A2(DP_OP_424J2_126_3477_n2566), .Y(DP_OP_423J2_125_3477_n2547) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1163 ( .A1(DP_OP_424J2_126_3477_n2689), 
        .A2(DP_OP_424J2_126_3477_n1953), .Y(DP_OP_422J2_124_3477_n1936) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1158 ( .A1(DP_OP_425J2_127_3477_n2690), 
        .A2(DP_OP_423J2_125_3477_n1948), .Y(DP_OP_423J2_125_3477_n1932) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U986 ( .A1(n302), .A2(
        DP_OP_424J2_126_3477_n2), .Y(DP_OP_423J2_125_3477_n162) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1243 ( .A1(DP_OP_422J2_124_3477_n2031), 
        .A2(DP_OP_422J2_124_3477_n2039), .Y(DP_OP_422J2_124_3477_n2015) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1243 ( .A1(DP_OP_422J2_124_3477_n1900), 
        .A2(DP_OP_425J2_127_3477_n2040), .Y(DP_OP_425J2_127_3477_n2016) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1243 ( .A1(DP_OP_424J2_126_3477_n2032), 
        .A2(DP_OP_424J2_126_3477_n2040), .Y(DP_OP_424J2_126_3477_n2016) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1624 ( .A1(DP_OP_422J2_124_3477_n2294), 
        .A2(DP_OP_423J2_125_3477_n2430), .Y(DP_OP_423J2_125_3477_n2398) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1647 ( .A1(DP_OP_424J2_126_3477_n2296), 
        .A2(DP_OP_425J2_127_3477_n2434), .Y(DP_OP_425J2_127_3477_n2417) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1823 ( .A1(DP_OP_424J2_126_3477_n2120), 
        .A2(DP_OP_425J2_127_3477_n2610), .Y(DP_OP_425J2_127_3477_n2593) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U991 ( .A1(n322), .A2(
        DP_OP_423J2_125_3477_n2), .Y(DP_OP_425J2_127_3477_n165) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1427 ( .A1(DP_OP_423J2_125_3477_n2643), 
        .A2(DP_OP_425J2_127_3477_n2217), .Y(DP_OP_425J2_127_3477_n2200) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U993 ( .A1(n307), .A2(
        DP_OP_425J2_127_3477_n2), .Y(DP_OP_425J2_127_3477_n169) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1163 ( .A1(DP_OP_423J2_125_3477_n2904), 
        .A2(DP_OP_425J2_127_3477_n1953), .Y(DP_OP_425J2_127_3477_n1936) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U995 ( .A1(n406), .A2(
        DP_OP_425J2_127_3477_n2), .Y(DP_OP_422J2_124_3477_n173) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1867 ( .A1(DP_OP_422J2_124_3477_n2777), 
        .A2(DP_OP_425J2_127_3477_n2654), .Y(DP_OP_425J2_127_3477_n2637) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U993 ( .A1(n411), .A2(
        DP_OP_423J2_125_3477_n2), .Y(DP_OP_422J2_124_3477_n169) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U994 ( .A1(n422), .A2(n338), .Y(
        DP_OP_422J2_124_3477_n171) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1338 ( .A1(DP_OP_425J2_127_3477_n2119), 
        .A2(DP_OP_425J2_127_3477_n2129), .Y(DP_OP_425J2_127_3477_n2111) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1932 ( .A1(DP_OP_424J2_126_3477_n2644), 
        .A2(DP_OP_425J2_127_3477_n2740), .Y(DP_OP_423J2_125_3477_n2703) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1060 ( .A1(DP_OP_423J2_125_3477_n1850), 
        .A2(DP_OP_423J2_125_3477_n1859), .Y(DP_OP_423J2_125_3477_n1834) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1720 ( .A1(DP_OP_423J2_125_3477_n2510), 
        .A2(DP_OP_423J2_125_3477_n2519), .Y(DP_OP_423J2_125_3477_n2494) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1632 ( .A1(DP_OP_422J2_124_3477_n2294), 
        .A2(DP_OP_423J2_125_3477_n2431), .Y(DP_OP_423J2_125_3477_n2406) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2116 ( .A1(DP_OP_423J2_125_3477_n2903), 
        .A2(DP_OP_425J2_127_3477_n2917), .Y(DP_OP_423J2_125_3477_n2887) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1756 ( .A1(DP_OP_423J2_125_3477_n2554), 
        .A2(DP_OP_423J2_125_3477_n2562), .Y(DP_OP_423J2_125_3477_n2530) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2028 ( .A1(DP_OP_424J2_126_3477_n2732), 
        .A2(DP_OP_423J2_125_3477_n2824), .Y(DP_OP_423J2_125_3477_n2799) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2026 ( .A1(DP_OP_425J2_127_3477_n2820), 
        .A2(DP_OP_425J2_127_3477_n2828), .Y(DP_OP_425J2_127_3477_n2796) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1289 ( .A1(DP_OP_424J2_126_3477_n2164), 
        .A2(DP_OP_423J2_125_3477_n2080), .Y(DP_OP_423J2_125_3477_n2063) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1190 ( .A1(DP_OP_423J2_125_3477_n2859), 
        .A2(DP_OP_425J2_127_3477_n1995), .Y(DP_OP_425J2_127_3477_n1963) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1207 ( .A1(DP_OP_424J2_126_3477_n2777), 
        .A2(DP_OP_425J2_127_3477_n1997), .Y(DP_OP_425J2_127_3477_n1980) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1418 ( .A1(DP_OP_423J2_125_3477_n2642), 
        .A2(DP_OP_423J2_125_3477_n2211), .Y(DP_OP_425J2_127_3477_n2191) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1228 ( .A1(DP_OP_424J2_126_3477_n2119), 
        .A2(DP_OP_423J2_125_3477_n2034), .Y(DP_OP_423J2_125_3477_n2002) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1859 ( .A1(DP_OP_422J2_124_3477_n2777), 
        .A2(DP_OP_424J2_126_3477_n2653), .Y(DP_OP_425J2_127_3477_n2629) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1119 ( .A1(DP_OP_424J2_126_3477_n2865), 
        .A2(DP_OP_423J2_125_3477_n1904), .Y(DP_OP_425J2_127_3477_n1892) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1251 ( .A1(DP_OP_422J2_124_3477_n1900), 
        .A2(DP_OP_425J2_127_3477_n2041), .Y(DP_OP_425J2_127_3477_n2024) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1245 ( .A1(DP_OP_424J2_126_3477_n2120), 
        .A2(DP_OP_424J2_126_3477_n2041), .Y(DP_OP_423J2_125_3477_n2019) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1201 ( .A1(DP_OP_423J2_125_3477_n1983), 
        .A2(DP_OP_423J2_125_3477_n1992), .Y(DP_OP_423J2_125_3477_n1975) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1911 ( .A1(DP_OP_423J2_125_3477_n1939), 
        .A2(DP_OP_422J2_124_3477_n2700), .Y(DP_OP_425J2_127_3477_n2681) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1938 ( .A1(DP_OP_425J2_127_3477_n2732), 
        .A2(DP_OP_425J2_127_3477_n2740), .Y(DP_OP_425J2_127_3477_n2708) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1594 ( .A1(DP_OP_422J2_124_3477_n2514), 
        .A2(DP_OP_422J2_124_3477_n2391), .Y(DP_OP_425J2_127_3477_n2364) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1454 ( .A1(DP_OP_424J2_126_3477_n2512), 
        .A2(DP_OP_425J2_127_3477_n2259), .Y(DP_OP_425J2_127_3477_n2227) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1198 ( .A1(DP_OP_425J2_127_3477_n2732), 
        .A2(DP_OP_424J2_126_3477_n1996), .Y(DP_OP_424J2_126_3477_n1971) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1770 ( .A1(DP_OP_423J2_125_3477_n2642), 
        .A2(DP_OP_424J2_126_3477_n2565), .Y(DP_OP_424J2_126_3477_n2540) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1770 ( .A1(DP_OP_422J2_124_3477_n2558), 
        .A2(DP_OP_422J2_124_3477_n2567), .Y(DP_OP_422J2_124_3477_n2542) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1154 ( .A1(DP_OP_422J2_124_3477_n1943), 
        .A2(DP_OP_422J2_124_3477_n1952), .Y(DP_OP_422J2_124_3477_n1927) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1462 ( .A1(DP_OP_422J2_124_3477_n2602), 
        .A2(DP_OP_424J2_126_3477_n2260), .Y(DP_OP_424J2_126_3477_n2235) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1418 ( .A1(DP_OP_422J2_124_3477_n2646), 
        .A2(DP_OP_424J2_126_3477_n2216), .Y(DP_OP_424J2_126_3477_n2191) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1726 ( .A1(DP_OP_424J2_126_3477_n2512), 
        .A2(DP_OP_424J2_126_3477_n2521), .Y(DP_OP_424J2_126_3477_n2496) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2026 ( .A1(DP_OP_424J2_126_3477_n2820), 
        .A2(DP_OP_424J2_126_3477_n2828), .Y(DP_OP_424J2_126_3477_n2796) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1119 ( .A1(DP_OP_422J2_124_3477_n1900), 
        .A2(DP_OP_422J2_124_3477_n1909), .Y(DP_OP_422J2_124_3477_n1892) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1911 ( .A1(DP_OP_425J2_127_3477_n2557), 
        .A2(DP_OP_422J2_124_3477_n2700), .Y(DP_OP_422J2_124_3477_n2683) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1119 ( .A1(DP_OP_425J2_127_3477_n2821), 
        .A2(DP_OP_424J2_126_3477_n1909), .Y(DP_OP_424J2_126_3477_n1892) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1207 ( .A1(DP_OP_424J2_126_3477_n1988), 
        .A2(DP_OP_422J2_124_3477_n1997), .Y(DP_OP_424J2_126_3477_n1980) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1251 ( .A1(DP_OP_424J2_126_3477_n2032), 
        .A2(DP_OP_424J2_126_3477_n2041), .Y(DP_OP_424J2_126_3477_n2024) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1955 ( .A1(DP_OP_424J2_126_3477_n2733), 
        .A2(DP_OP_424J2_126_3477_n2742), .Y(DP_OP_424J2_126_3477_n2725) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1198 ( .A1(DP_OP_425J2_127_3477_n2119), 
        .A2(DP_OP_422J2_124_3477_n1996), .Y(DP_OP_422J2_124_3477_n1971) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1859 ( .A1(DP_OP_425J2_127_3477_n2120), 
        .A2(DP_OP_424J2_126_3477_n2653), .Y(DP_OP_424J2_126_3477_n2629) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1551 ( .A1(DP_OP_423J2_125_3477_n2247), 
        .A2(DP_OP_423J2_125_3477_n2343), .Y(DP_OP_424J2_126_3477_n2324) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1727 ( .A1(DP_OP_423J2_125_3477_n2599), 
        .A2(DP_OP_424J2_126_3477_n2521), .Y(DP_OP_424J2_126_3477_n2497) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2042 ( .A1(DP_OP_422J2_124_3477_n2820), 
        .A2(DP_OP_422J2_124_3477_n2830), .Y(DP_OP_422J2_124_3477_n2812) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1726 ( .A1(DP_OP_422J2_124_3477_n2514), 
        .A2(DP_OP_422J2_124_3477_n2523), .Y(DP_OP_422J2_124_3477_n2498) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1295 ( .A1(DP_OP_423J2_125_3477_n2643), 
        .A2(n441), .Y(DP_OP_422J2_124_3477_n2067) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1251 ( .A1(DP_OP_422J2_124_3477_n2031), 
        .A2(DP_OP_422J2_124_3477_n2040), .Y(DP_OP_422J2_124_3477_n2023) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1595 ( .A1(DP_OP_424J2_126_3477_n2381), 
        .A2(DP_OP_424J2_126_3477_n2389), .Y(DP_OP_424J2_126_3477_n2365) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1762 ( .A1(DP_OP_422J2_124_3477_n2558), 
        .A2(DP_OP_422J2_124_3477_n2566), .Y(DP_OP_422J2_124_3477_n2534) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1322 ( .A1(DP_OP_422J2_124_3477_n2118), 
        .A2(DP_OP_423J2_125_3477_n2122), .Y(DP_OP_422J2_124_3477_n2094) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1551 ( .A1(DP_OP_422J2_124_3477_n2339), 
        .A2(DP_OP_422J2_124_3477_n2347), .Y(DP_OP_422J2_124_3477_n2323) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1120 ( .A1(DP_OP_425J2_127_3477_n1901), 
        .A2(DP_OP_424J2_126_3477_n1909), .Y(DP_OP_425J2_127_3477_n1893) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2043 ( .A1(DP_OP_424J2_126_3477_n2821), 
        .A2(DP_OP_424J2_126_3477_n2830), .Y(DP_OP_424J2_126_3477_n2813) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2130 ( .A1(DP_OP_422J2_124_3477_n2908), 
        .A2(DP_OP_422J2_124_3477_n2918), .Y(DP_OP_422J2_124_3477_n2900) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2130 ( .A1(DP_OP_425J2_127_3477_n1855), 
        .A2(DP_OP_422J2_124_3477_n2918), .Y(DP_OP_424J2_126_3477_n2900) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1002 ( .A1(n401), .A2(n341), .Y(
        DP_OP_424J2_126_3477_n1775) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1000 ( .A1(n374), .A2(n340), .Y(
        DP_OP_424J2_126_3477_n1774) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1001 ( .A1(n413), .A2(n343), .Y(
        DP_OP_422J2_124_3477_n189) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U994 ( .A1(n310), .A2(n341), .Y(
        DP_OP_425J2_127_3477_n171) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1330 ( .A1(DP_OP_424J2_126_3477_n2119), 
        .A2(DP_OP_422J2_124_3477_n2127), .Y(DP_OP_424J2_126_3477_n2103) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U987 ( .A1(n306), .A2(n342), .Y(
        DP_OP_423J2_125_3477_n164) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U993 ( .A1(n415), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_424J2_126_3477_n169) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U996 ( .A1(n290), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_423J2_125_3477_n1770) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U994 ( .A1(n295), .A2(n342), .Y(
        DP_OP_423J2_125_3477_n1769) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2125 ( .A1(DP_OP_423J2_125_3477_n2904), 
        .A2(DP_OP_423J2_125_3477_n2913), .Y(DP_OP_423J2_125_3477_n2896) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1465 ( .A1(DP_OP_423J2_125_3477_n2247), 
        .A2(DP_OP_423J2_125_3477_n2256), .Y(DP_OP_423J2_125_3477_n2239) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1902 ( .A1(DP_OP_425J2_127_3477_n2688), 
        .A2(DP_OP_422J2_124_3477_n2699), .Y(DP_OP_425J2_127_3477_n2672) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U992 ( .A1(n300), .A2(n343), .Y(
        DP_OP_423J2_125_3477_n174) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1000 ( .A1(n294), .A2(n340), .Y(
        DP_OP_425J2_127_3477_n1774) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U993 ( .A1(n397), .A2(n341), .Y(
        DP_OP_423J2_125_3477_n176) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1002 ( .A1(n289), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_425J2_127_3477_n1775) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1587 ( .A1(DP_OP_425J2_127_3477_n2381), 
        .A2(DP_OP_423J2_125_3477_n2386), .Y(DP_OP_425J2_127_3477_n2357) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1536 ( .A1(DP_OP_423J2_125_3477_n2334), 
        .A2(DP_OP_422J2_124_3477_n2346), .Y(DP_OP_423J2_125_3477_n2310) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U997 ( .A1(n312), .A2(n339), .Y(
        DP_OP_425J2_127_3477_n177) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1278 ( .A1(DP_OP_425J2_127_3477_n2075), 
        .A2(DP_OP_425J2_127_3477_n2083), .Y(DP_OP_425J2_127_3477_n2051) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1990 ( .A1(DP_OP_423J2_125_3477_n1850), 
        .A2(DP_OP_425J2_127_3477_n2785), .Y(DP_OP_425J2_127_3477_n2760) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1471 ( .A1(DP_OP_425J2_127_3477_n2252), 
        .A2(DP_OP_425J2_127_3477_n2261), .Y(DP_OP_425J2_127_3477_n2244) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1946 ( .A1(DP_OP_424J2_126_3477_n2732), 
        .A2(DP_OP_424J2_126_3477_n2741), .Y(DP_OP_424J2_126_3477_n2716) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1941 ( .A1(DP_OP_422J2_124_3477_n1988), 
        .A2(DP_OP_424J2_126_3477_n2741), .Y(DP_OP_423J2_125_3477_n2712) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1602 ( .A1(DP_OP_422J2_124_3477_n2250), 
        .A2(DP_OP_424J2_126_3477_n2390), .Y(DP_OP_424J2_126_3477_n2372) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1946 ( .A1(DP_OP_425J2_127_3477_n2732), 
        .A2(DP_OP_425J2_127_3477_n2741), .Y(DP_OP_425J2_127_3477_n2716) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1947 ( .A1(DP_OP_422J2_124_3477_n2733), 
        .A2(DP_OP_422J2_124_3477_n2741), .Y(DP_OP_422J2_124_3477_n2717) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1888 ( .A1(DP_OP_425J2_127_3477_n2163), 
        .A2(DP_OP_424J2_126_3477_n2696), .Y(DP_OP_423J2_125_3477_n2662) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1096 ( .A1(DP_OP_425J2_127_3477_n2732), 
        .A2(DP_OP_422J2_124_3477_n1907), .Y(DP_OP_423J2_125_3477_n1870) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1602 ( .A1(DP_OP_424J2_126_3477_n2339), 
        .A2(DP_OP_423J2_125_3477_n2388), .Y(DP_OP_425J2_127_3477_n2372) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1894 ( .A1(DP_OP_425J2_127_3477_n2075), 
        .A2(DP_OP_424J2_126_3477_n2696), .Y(DP_OP_424J2_126_3477_n2664) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1146 ( .A1(DP_OP_423J2_125_3477_n1850), 
        .A2(n442), .Y(DP_OP_424J2_126_3477_n1919) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1603 ( .A1(DP_OP_425J2_127_3477_n2381), 
        .A2(DP_OP_424J2_126_3477_n2390), .Y(DP_OP_425J2_127_3477_n2373) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1946 ( .A1(DP_OP_422J2_124_3477_n2732), 
        .A2(DP_OP_422J2_124_3477_n2741), .Y(DP_OP_422J2_124_3477_n2716) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U71 ( .A1(DP_OP_423J2_125_3477_n181), .A2(
        DP_OP_423J2_125_3477_n186), .Y(DP_OP_423J2_125_3477_n65) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U19 ( .A1(DP_OP_422J2_124_3477_n38), .A2(
        DP_OP_422J2_124_3477_n41), .Y(DP_OP_422J2_124_3477_n36) );
  AO221X1_HVT U3 ( .A1(1'b1), .A2(n537), .A3(n407), .A4(conv2_sum_d[28]), .A5(
        n214), .Y(n538) );
  AO221X1_HVT U4 ( .A1(1'b1), .A2(n549), .A3(n419), .A4(conv2_sum_d[20]), .A5(
        n211), .Y(n585) );
  AO221X1_HVT U5 ( .A1(1'b1), .A2(n463), .A3(n405), .A4(conv2_sum_b[28]), .A5(
        n103), .Y(n464) );
  AO221X1_HVT U6 ( .A1(1'b1), .A2(n562), .A3(n404), .A4(conv2_sum_d[12]), .A5(
        n101), .Y(n565) );
  AO221X1_HVT U7 ( .A1(1'b1), .A2(n478), .A3(n406), .A4(conv2_sum_b[20]), .A5(
        n99), .Y(n514) );
  AO221X1_HVT U8 ( .A1(1'b1), .A2(n607), .A3(tmp_big2[28]), .A4(n72), .A5(n73), 
        .Y(n608) );
  AO221X1_HVT U9 ( .A1(1'b1), .A2(n632), .A3(tmp_big2[12]), .A4(n701), .A5(n71), .Y(n635) );
  AO221X1_HVT U10 ( .A1(1'b1), .A2(n619), .A3(tmp_big2[20]), .A4(n51), .A5(n52), .Y(n649) );
  AO221X1_HVT U11 ( .A1(1'b1), .A2(n491), .A3(n403), .A4(conv2_sum_b[12]), 
        .A5(n3), .Y(n494) );
  OA221X1_HVT U12 ( .A1(n155), .A2(n464), .A3(n462), .A4(conv2_sum_b[30]), 
        .A5(n157), .Y(n158) );
  OA221X1_HVT U13 ( .A1(1'b0), .A2(DP_OP_424J2_126_3477_n60), .A3(
        DP_OP_424J2_126_3477_n59), .A4(DP_OP_424J2_126_3477_n65), .A5(n26), 
        .Y(DP_OP_424J2_126_3477_n56) );
  OA221X1_HVT U14 ( .A1(1'b0), .A2(DP_OP_425J2_127_3477_n60), .A3(
        DP_OP_425J2_127_3477_n59), .A4(DP_OP_425J2_127_3477_n65), .A5(n24), 
        .Y(DP_OP_425J2_127_3477_n56) );
  OA221X1_HVT U15 ( .A1(1'b0), .A2(DP_OP_422J2_124_3477_n60), .A3(
        DP_OP_422J2_124_3477_n59), .A4(DP_OP_422J2_124_3477_n65), .A5(n21), 
        .Y(DP_OP_422J2_124_3477_n56) );
  OA221X1_HVT U16 ( .A1(1'b0), .A2(DP_OP_423J2_125_3477_n58), .A3(
        DP_OP_423J2_125_3477_n57), .A4(DP_OP_423J2_125_3477_n63), .A5(n18), 
        .Y(DP_OP_423J2_125_3477_n54) );
  OA221X1_HVT U17 ( .A1(1'b0), .A2(DP_OP_424J2_126_3477_n99), .A3(
        DP_OP_424J2_126_3477_n98), .A4(DP_OP_424J2_126_3477_n102), .A5(n14), 
        .Y(DP_OP_424J2_126_3477_n95) );
  OA221X1_HVT U18 ( .A1(1'b0), .A2(DP_OP_425J2_127_3477_n99), .A3(
        DP_OP_425J2_127_3477_n98), .A4(DP_OP_425J2_127_3477_n102), .A5(n12), 
        .Y(DP_OP_425J2_127_3477_n95) );
  OA221X1_HVT U19 ( .A1(1'b0), .A2(DP_OP_422J2_124_3477_n99), .A3(
        DP_OP_422J2_124_3477_n98), .A4(DP_OP_422J2_124_3477_n102), .A5(n900), 
        .Y(DP_OP_422J2_124_3477_n95) );
  OA221X1_HVT U20 ( .A1(1'b0), .A2(DP_OP_423J2_125_3477_n97), .A3(
        DP_OP_423J2_125_3477_n96), .A4(DP_OP_423J2_125_3477_n100), .A5(n6), 
        .Y(DP_OP_423J2_125_3477_n93) );
  INVX0_HVT U21 ( .A(n352), .Y(n1) );
  AOI22X1_HVT U22 ( .A1(n352), .A2(conv1_sram_rdata_weight[79]), .A3(n1), .A4(
        conv2_sram_rdata_weight[79]), .Y(n450) );
  AO22X1_HVT U23 ( .A1(n439), .A2(conv2_sram_rdata_weight[98]), .A3(
        conv1_sram_rdata_weight[98]), .A4(n349), .Y(conv_weight_box[92]) );
  INVX0_HVT U25 ( .A(n480), .Y(n3) );
  INVX0_HVT U27 ( .A(DP_OP_423J2_125_3477_n102), .Y(n5010) );
  OR3X1_HVT U28 ( .A1(n5010), .A2(DP_OP_423J2_125_3477_n99), .A3(
        DP_OP_423J2_125_3477_n96), .Y(n6) );
  INVX0_HVT U30 ( .A(DP_OP_422J2_124_3477_n104), .Y(n8) );
  OR3X1_HVT U31 ( .A1(n8), .A2(DP_OP_422J2_124_3477_n101), .A3(
        DP_OP_422J2_124_3477_n98), .Y(n900) );
  INVX0_HVT U33 ( .A(DP_OP_425J2_127_3477_n104), .Y(n11) );
  OR3X1_HVT U34 ( .A1(n11), .A2(DP_OP_425J2_127_3477_n101), .A3(
        DP_OP_425J2_127_3477_n98), .Y(n12) );
  OR3X1_HVT U35 ( .A1(n13), .A2(DP_OP_424J2_126_3477_n101), .A3(
        DP_OP_424J2_126_3477_n98), .Y(n14) );
  INVX0_HVT U37 ( .A(DP_OP_424J2_126_3477_n104), .Y(n13) );
  INVX0_HVT U39 ( .A(DP_OP_423J2_125_3477_n66), .Y(n17) );
  NAND2X0_HVT U40 ( .A1(DP_OP_423J2_125_3477_n55), .A2(n17), .Y(n18) );
  INVX0_HVT U42 ( .A(DP_OP_422J2_124_3477_n68), .Y(n20) );
  NAND2X0_HVT U43 ( .A1(DP_OP_422J2_124_3477_n57), .A2(n20), .Y(n21) );
  INVX0_HVT U45 ( .A(DP_OP_425J2_127_3477_n68), .Y(n23) );
  NAND2X0_HVT U46 ( .A1(DP_OP_425J2_127_3477_n57), .A2(n23), .Y(n24) );
  INVX0_HVT U47 ( .A(DP_OP_424J2_126_3477_n68), .Y(n25) );
  NAND2X0_HVT U48 ( .A1(DP_OP_424J2_126_3477_n57), .A2(n25), .Y(n26) );
  INVX0_HVT U50 ( .A(n353), .Y(n28) );
  AOI22X1_HVT U51 ( .A1(n353), .A2(conv1_sram_rdata_weight[74]), .A3(n28), 
        .A4(conv2_sram_rdata_weight[74]), .Y(n444) );
  NAND2X0_HVT U52 ( .A1(n646), .A2(tmp_big1[6]), .Y(n29) );
  INVX0_HVT U53 ( .A(tmp_big1[6]), .Y(n30) );
  AO22X1_HVT U54 ( .A1(tmp_big2[7]), .A2(n685), .A3(tmp_big2[6]), .A4(n30), 
        .Y(n31) );
  NAND2X0_HVT U55 ( .A1(n645), .A2(tmp_big1[4]), .Y(n32) );
  OA21X1_HVT U56 ( .A1(n642), .A2(n643), .A3(n644), .Y(n33) );
  OA222X1_HVT U57 ( .A1(n32), .A2(tmp_big2[4]), .A3(tmp_big2[5]), .A4(n684), 
        .A5(n33), .A6(n641), .Y(n34) );
  OA222X1_HVT U58 ( .A1(n29), .A2(tmp_big2[6]), .A3(n31), .A4(n34), .A5(
        tmp_big2[7]), .A6(n685), .Y(n651) );
  OA22X1_HVT U59 ( .A1(conv2_sum_d[22]), .A2(n548), .A3(conv2_sum_d[23]), .A4(
        n383), .Y(n35) );
  OA22X1_HVT U60 ( .A1(conv2_sum_d[20]), .A2(n540), .A3(n426), .A4(
        conv2_sum_d[21]), .Y(n36) );
  OA21X1_HVT U61 ( .A1(n586), .A2(n545), .A3(n546), .Y(n37) );
  OA22X1_HVT U62 ( .A1(n549), .A2(n36), .A3(n585), .A4(n37), .Y(n38) );
  OR3X1_HVT U63 ( .A1(n565), .A2(n566), .A3(n564), .Y(n39) );
  OR3X1_HVT U64 ( .A1(n585), .A2(n586), .A3(n584), .Y(n40) );
  AO221X1_HVT U65 ( .A1(n588), .A2(n587), .A3(n588), .A4(n39), .A5(n40), .Y(
        n41) );
  NAND3X0_HVT U66 ( .A1(n35), .A2(n38), .A3(n41), .Y(n589) );
  INVX0_HVT U67 ( .A(n432), .Y(n42) );
  OR3X1_HVT U68 ( .A1(channel[4]), .A2(channel[1]), .A3(channel[3]), .Y(n43)
         );
  AO222X1_HVT U69 ( .A1(n42), .A2(channel[0]), .A3(n42), .A4(channel[2]), .A5(
        n42), .A6(n43), .Y(n437) );
  NAND2X0_HVT U70 ( .A1(DP_OP_423J2_125_3477_n67), .A2(
        DP_OP_423J2_125_3477_n66), .Y(n44) );
  HADDX1_HVT U71 ( .A0(DP_OP_423J2_125_3477_n71), .B0(n44), .SO(
        n_conv2_sum_b[14]) );
  NAND2X0_HVT U72 ( .A1(DP_OP_422J2_124_3477_n69), .A2(
        DP_OP_422J2_124_3477_n68), .Y(n45) );
  HADDX1_HVT U73 ( .A0(DP_OP_422J2_124_3477_n73), .B0(n45), .SO(
        n_conv2_sum_a[14]) );
  NAND2X0_HVT U74 ( .A1(DP_OP_425J2_127_3477_n69), .A2(
        DP_OP_425J2_127_3477_n68), .Y(n46) );
  HADDX1_HVT U75 ( .A0(DP_OP_425J2_127_3477_n73), .B0(n46), .SO(
        n_conv2_sum_d[14]) );
  NAND2X0_HVT U76 ( .A1(DP_OP_424J2_126_3477_n69), .A2(
        DP_OP_424J2_126_3477_n68), .Y(n47) );
  HADDX1_HVT U77 ( .A0(DP_OP_424J2_126_3477_n73), .B0(n47), .SO(
        n_conv2_sum_c[14]) );
  INVX0_HVT U78 ( .A(n350), .Y(n48) );
  AOI22X1_HVT U79 ( .A1(n350), .A2(conv1_sram_rdata_weight[62]), .A3(n48), 
        .A4(conv2_sram_rdata_weight[62]), .Y(n452) );
  AO22X1_HVT U80 ( .A1(n438), .A2(conv2_sram_rdata_weight[42]), .A3(
        conv1_sram_rdata_weight[42]), .A4(n334), .Y(DP_OP_425J2_127_3477_n3110) );
  INVX0_HVT U81 ( .A(n453), .Y(n49) );
  AOI22X1_HVT U82 ( .A1(n453), .A2(conv2_sram_rdata_weight[22]), .A3(n49), 
        .A4(conv1_sram_rdata_weight[22]), .Y(n442) );
  INVX0_HVT U84 ( .A(tmp_big1[20]), .Y(n51) );
  INVX0_HVT U85 ( .A(n611), .Y(n52) );
  NAND2X0_HVT U86 ( .A1(DP_OP_423J2_125_3477_n110), .A2(
        DP_OP_423J2_125_3477_n108), .Y(n53) );
  AND2X1_HVT U87 ( .A1(n53), .A2(DP_OP_423J2_125_3477_n109), .Y(
        DP_OP_423J2_125_3477_n105) );
  NAND2X0_HVT U88 ( .A1(DP_OP_422J2_124_3477_n112), .A2(
        DP_OP_422J2_124_3477_n110), .Y(n54) );
  AND2X1_HVT U89 ( .A1(n54), .A2(DP_OP_422J2_124_3477_n111), .Y(
        DP_OP_422J2_124_3477_n107) );
  NAND2X0_HVT U90 ( .A1(DP_OP_425J2_127_3477_n112), .A2(
        DP_OP_425J2_127_3477_n110), .Y(n55) );
  AND2X1_HVT U91 ( .A1(n55), .A2(DP_OP_425J2_127_3477_n111), .Y(
        DP_OP_425J2_127_3477_n107) );
  NAND2X0_HVT U92 ( .A1(DP_OP_424J2_126_3477_n112), .A2(
        DP_OP_424J2_126_3477_n110), .Y(n56) );
  AND2X1_HVT U93 ( .A1(n56), .A2(DP_OP_424J2_126_3477_n111), .Y(
        DP_OP_424J2_126_3477_n107) );
  INVX0_HVT U94 ( .A(DP_OP_423J2_125_3477_n57), .Y(n57) );
  NAND2X0_HVT U95 ( .A1(DP_OP_423J2_125_3477_n64), .A2(
        DP_OP_423J2_125_3477_n60), .Y(n58) );
  AO22X1_HVT U96 ( .A1(n57), .A2(DP_OP_423J2_125_3477_n58), .A3(
        DP_OP_423J2_125_3477_n63), .A4(n58), .Y(n59) );
  NAND4X0_HVT U97 ( .A1(n57), .A2(DP_OP_423J2_125_3477_n58), .A3(
        DP_OP_423J2_125_3477_n63), .A4(n58), .Y(n60) );
  NAND2X0_HVT U98 ( .A1(n59), .A2(n60), .Y(n_conv2_sum_b[16]) );
  AND2X1_HVT U99 ( .A1(DP_OP_422J2_124_3477_n62), .A2(DP_OP_422J2_124_3477_n65), .Y(n61) );
  HADDX1_HVT U100 ( .A0(n61), .B0(DP_OP_422J2_124_3477_n66), .SO(
        n_conv2_sum_a[15]) );
  INVX0_HVT U101 ( .A(DP_OP_425J2_127_3477_n59), .Y(n62) );
  NAND2X0_HVT U102 ( .A1(DP_OP_425J2_127_3477_n66), .A2(
        DP_OP_425J2_127_3477_n62), .Y(n63) );
  AO22X1_HVT U103 ( .A1(n62), .A2(DP_OP_425J2_127_3477_n60), .A3(
        DP_OP_425J2_127_3477_n65), .A4(n63), .Y(n64) );
  NAND4X0_HVT U104 ( .A1(n62), .A2(DP_OP_425J2_127_3477_n60), .A3(
        DP_OP_425J2_127_3477_n65), .A4(n63), .Y(n65) );
  NAND2X0_HVT U105 ( .A1(n64), .A2(n65), .Y(n_conv2_sum_d[16]) );
  AND2X1_HVT U106 ( .A1(DP_OP_424J2_126_3477_n62), .A2(
        DP_OP_424J2_126_3477_n65), .Y(n66) );
  HADDX1_HVT U107 ( .A0(n66), .B0(DP_OP_424J2_126_3477_n66), .SO(
        n_conv2_sum_c[15]) );
  INVX0_HVT U108 ( .A(n348), .Y(n67) );
  AOI22X1_HVT U109 ( .A1(n348), .A2(conv1_sram_rdata_weight[58]), .A3(n67), 
        .A4(conv2_sram_rdata_weight[58]), .Y(n451) );
  INVX0_HVT U110 ( .A(n438), .Y(n68) );
  AOI22X1_HVT U111 ( .A1(n438), .A2(conv2_sram_rdata_weight[70]), .A3(n68), 
        .A4(conv1_sram_rdata_weight[70]), .Y(n443) );
  AO22X1_HVT U112 ( .A1(n453), .A2(conv2_sram_rdata_weight[25]), .A3(
        conv1_sram_rdata_weight[25]), .A4(n336), .Y(conv_weight_box[23]) );
  INVX0_HVT U114 ( .A(tmp_big1[12]), .Y(n701) );
  INVX0_HVT U115 ( .A(n621), .Y(n71) );
  INVX0_HVT U116 ( .A(tmp_big1[28]), .Y(n72) );
  INVX0_HVT U117 ( .A(n596), .Y(n73) );
  NAND2X0_HVT U119 ( .A1(DP_OP_423J2_125_3477_n116), .A2(
        DP_OP_423J2_125_3477_n118), .Y(n75) );
  AND2X1_HVT U120 ( .A1(n75), .A2(DP_OP_423J2_125_3477_n117), .Y(
        DP_OP_423J2_125_3477_n113) );
  NAND2X0_HVT U121 ( .A1(DP_OP_423J2_125_3477_n49), .A2(
        DP_OP_423J2_125_3477_n43), .Y(n76) );
  AND2X1_HVT U122 ( .A1(n76), .A2(DP_OP_423J2_125_3477_n44), .Y(
        DP_OP_423J2_125_3477_n40) );
  NAND2X0_HVT U123 ( .A1(DP_OP_422J2_124_3477_n118), .A2(
        DP_OP_422J2_124_3477_n120), .Y(n77) );
  AND2X1_HVT U124 ( .A1(n77), .A2(DP_OP_422J2_124_3477_n119), .Y(
        DP_OP_422J2_124_3477_n115) );
  NAND2X0_HVT U125 ( .A1(DP_OP_422J2_124_3477_n51), .A2(
        DP_OP_422J2_124_3477_n45), .Y(n78) );
  AND2X1_HVT U126 ( .A1(n78), .A2(DP_OP_422J2_124_3477_n46), .Y(
        DP_OP_422J2_124_3477_n42) );
  NAND2X0_HVT U127 ( .A1(DP_OP_425J2_127_3477_n118), .A2(
        DP_OP_425J2_127_3477_n120), .Y(n79) );
  AND2X1_HVT U128 ( .A1(n79), .A2(DP_OP_425J2_127_3477_n119), .Y(
        DP_OP_425J2_127_3477_n115) );
  NAND2X0_HVT U129 ( .A1(DP_OP_425J2_127_3477_n51), .A2(
        DP_OP_425J2_127_3477_n45), .Y(n80) );
  AND2X1_HVT U130 ( .A1(n80), .A2(DP_OP_425J2_127_3477_n46), .Y(
        DP_OP_425J2_127_3477_n42) );
  NAND2X0_HVT U131 ( .A1(DP_OP_424J2_126_3477_n118), .A2(
        DP_OP_424J2_126_3477_n120), .Y(n81) );
  AND2X1_HVT U132 ( .A1(n81), .A2(DP_OP_424J2_126_3477_n119), .Y(
        DP_OP_424J2_126_3477_n115) );
  NAND2X0_HVT U133 ( .A1(DP_OP_424J2_126_3477_n51), .A2(
        DP_OP_424J2_126_3477_n45), .Y(n82) );
  AND2X1_HVT U134 ( .A1(n82), .A2(DP_OP_424J2_126_3477_n46), .Y(
        DP_OP_424J2_126_3477_n42) );
  AND2X1_HVT U135 ( .A1(DP_OP_423J2_125_3477_n88), .A2(
        DP_OP_423J2_125_3477_n91), .Y(n83) );
  HADDX1_HVT U136 ( .A0(n83), .B0(DP_OP_423J2_125_3477_n92), .SO(
        n_conv2_sum_b[10]) );
  AND2X1_HVT U137 ( .A1(DP_OP_423J2_125_3477_n60), .A2(
        DP_OP_423J2_125_3477_n63), .Y(n84) );
  HADDX1_HVT U138 ( .A0(n84), .B0(DP_OP_423J2_125_3477_n64), .SO(
        n_conv2_sum_b[15]) );
  AND2X1_HVT U139 ( .A1(DP_OP_422J2_124_3477_n90), .A2(
        DP_OP_422J2_124_3477_n93), .Y(n85) );
  HADDX1_HVT U140 ( .A0(n85), .B0(DP_OP_422J2_124_3477_n94), .SO(
        n_conv2_sum_a[10]) );
  INVX0_HVT U141 ( .A(DP_OP_422J2_124_3477_n59), .Y(n86) );
  NAND2X0_HVT U142 ( .A1(DP_OP_422J2_124_3477_n66), .A2(
        DP_OP_422J2_124_3477_n62), .Y(n87) );
  AO22X1_HVT U143 ( .A1(n86), .A2(DP_OP_422J2_124_3477_n60), .A3(
        DP_OP_422J2_124_3477_n65), .A4(n87), .Y(n88) );
  NAND4X0_HVT U144 ( .A1(n86), .A2(DP_OP_422J2_124_3477_n60), .A3(
        DP_OP_422J2_124_3477_n65), .A4(n87), .Y(n89) );
  NAND2X0_HVT U145 ( .A1(n88), .A2(n89), .Y(n_conv2_sum_a[16]) );
  AND2X1_HVT U146 ( .A1(DP_OP_425J2_127_3477_n90), .A2(
        DP_OP_425J2_127_3477_n93), .Y(n901) );
  HADDX1_HVT U147 ( .A0(n901), .B0(DP_OP_425J2_127_3477_n94), .SO(
        n_conv2_sum_d[10]) );
  AND2X1_HVT U148 ( .A1(DP_OP_425J2_127_3477_n62), .A2(
        DP_OP_425J2_127_3477_n65), .Y(n91) );
  HADDX1_HVT U149 ( .A0(n91), .B0(DP_OP_425J2_127_3477_n66), .SO(
        n_conv2_sum_d[15]) );
  AND2X1_HVT U150 ( .A1(DP_OP_424J2_126_3477_n90), .A2(
        DP_OP_424J2_126_3477_n93), .Y(n92) );
  HADDX1_HVT U151 ( .A0(n92), .B0(DP_OP_424J2_126_3477_n94), .SO(
        n_conv2_sum_c[10]) );
  INVX0_HVT U152 ( .A(DP_OP_424J2_126_3477_n59), .Y(n93) );
  NAND2X0_HVT U153 ( .A1(DP_OP_424J2_126_3477_n66), .A2(
        DP_OP_424J2_126_3477_n62), .Y(n94) );
  AO22X1_HVT U154 ( .A1(n93), .A2(DP_OP_424J2_126_3477_n60), .A3(
        DP_OP_424J2_126_3477_n65), .A4(n94), .Y(n95) );
  NAND4X0_HVT U155 ( .A1(n93), .A2(DP_OP_424J2_126_3477_n60), .A3(
        DP_OP_424J2_126_3477_n65), .A4(n94), .Y(n96) );
  NAND2X0_HVT U156 ( .A1(n95), .A2(n96), .Y(n_conv2_sum_c[16]) );
  INVX0_HVT U157 ( .A(n350), .Y(n97) );
  AOI22X1_HVT U158 ( .A1(n350), .A2(conv1_sram_rdata_weight[86]), .A3(n97), 
        .A4(conv2_sram_rdata_weight[86]), .Y(n445) );
  AO22X1_HVT U159 ( .A1(n438), .A2(conv2_sram_rdata_weight[41]), .A3(
        conv1_sram_rdata_weight[41]), .A4(n336), .Y(conv_weight_box[38]) );
  INVX0_HVT U161 ( .A(n467), .Y(n99) );
  INVX0_HVT U163 ( .A(n551), .Y(n101) );
  INVX0_HVT U165 ( .A(n455), .Y(n103) );
  OA22X1_HVT U166 ( .A1(tmp_big2[22]), .A2(n618), .A3(tmp_big2[23]), .A4(n674), 
        .Y(n104) );
  OA22X1_HVT U167 ( .A1(n610), .A2(tmp_big2[20]), .A3(n672), .A4(tmp_big2[21]), 
        .Y(n105) );
  OA21X1_HVT U168 ( .A1(n650), .A2(n615), .A3(n616), .Y(n106) );
  OA22X1_HVT U169 ( .A1(n619), .A2(n105), .A3(n649), .A4(n106), .Y(n107) );
  OR3X1_HVT U170 ( .A1(n649), .A2(n650), .A3(n648), .Y(n108) );
  AO221X1_HVT U171 ( .A1(n653), .A2(n651), .A3(n653), .A4(n652), .A5(n108), 
        .Y(n109) );
  NAND3X0_HVT U172 ( .A1(n104), .A2(n107), .A3(n109), .Y(n654) );
  NAND2X0_HVT U173 ( .A1(DP_OP_423J2_125_3477_n124), .A2(
        DP_OP_423J2_125_3477_n126), .Y(n110) );
  AND2X1_HVT U174 ( .A1(n110), .A2(DP_OP_423J2_125_3477_n125), .Y(
        DP_OP_423J2_125_3477_n121) );
  NAND2X0_HVT U175 ( .A1(DP_OP_422J2_124_3477_n126), .A2(
        DP_OP_422J2_124_3477_n128), .Y(n111) );
  AND2X1_HVT U176 ( .A1(n111), .A2(DP_OP_422J2_124_3477_n127), .Y(
        DP_OP_422J2_124_3477_n123) );
  NAND2X0_HVT U177 ( .A1(DP_OP_425J2_127_3477_n126), .A2(
        DP_OP_425J2_127_3477_n128), .Y(n112) );
  AND2X1_HVT U178 ( .A1(n112), .A2(DP_OP_425J2_127_3477_n127), .Y(
        DP_OP_425J2_127_3477_n123) );
  NAND2X0_HVT U179 ( .A1(DP_OP_424J2_126_3477_n126), .A2(
        DP_OP_424J2_126_3477_n128), .Y(n113) );
  AND2X1_HVT U180 ( .A1(n113), .A2(DP_OP_424J2_126_3477_n127), .Y(
        DP_OP_424J2_126_3477_n123) );
  INVX0_HVT U181 ( .A(DP_OP_423J2_125_3477_n103), .Y(n114) );
  NAND2X0_HVT U182 ( .A1(n114), .A2(DP_OP_423J2_125_3477_n104), .Y(n115) );
  HADDX1_HVT U183 ( .A0(DP_OP_423J2_125_3477_n105), .B0(n115), .SO(
        n_conv2_sum_b[7]) );
  INVX0_HVT U184 ( .A(DP_OP_423J2_125_3477_n85), .Y(n116) );
  NAND2X0_HVT U185 ( .A1(DP_OP_423J2_125_3477_n92), .A2(
        DP_OP_423J2_125_3477_n88), .Y(n117) );
  AO22X1_HVT U186 ( .A1(n116), .A2(DP_OP_423J2_125_3477_n86), .A3(
        DP_OP_423J2_125_3477_n91), .A4(n117), .Y(n118) );
  NAND4X0_HVT U187 ( .A1(n116), .A2(DP_OP_423J2_125_3477_n86), .A3(
        DP_OP_423J2_125_3477_n91), .A4(n117), .Y(n119) );
  NAND2X0_HVT U188 ( .A1(n118), .A2(n119), .Y(n_conv2_sum_b[11]) );
  OA21X1_HVT U189 ( .A1(DP_OP_423J2_125_3477_n53), .A2(
        DP_OP_423J2_125_3477_n71), .A3(DP_OP_423J2_125_3477_n54), .Y(n120) );
  INVX0_HVT U190 ( .A(DP_OP_423J2_125_3477_n50), .Y(n121) );
  NAND2X0_HVT U191 ( .A1(n121), .A2(DP_OP_423J2_125_3477_n51), .Y(n122) );
  HADDX1_HVT U192 ( .A0(n120), .B0(n122), .SO(n_conv2_sum_b[17]) );
  INVX0_HVT U193 ( .A(DP_OP_422J2_124_3477_n105), .Y(n123) );
  NAND2X0_HVT U194 ( .A1(n123), .A2(DP_OP_422J2_124_3477_n106), .Y(n124) );
  HADDX1_HVT U195 ( .A0(DP_OP_422J2_124_3477_n107), .B0(n124), .SO(
        n_conv2_sum_a[7]) );
  INVX0_HVT U196 ( .A(DP_OP_422J2_124_3477_n87), .Y(n125) );
  NAND2X0_HVT U197 ( .A1(DP_OP_422J2_124_3477_n94), .A2(
        DP_OP_422J2_124_3477_n90), .Y(n126) );
  AO22X1_HVT U198 ( .A1(n125), .A2(DP_OP_422J2_124_3477_n88), .A3(
        DP_OP_422J2_124_3477_n93), .A4(n126), .Y(n127) );
  NAND4X0_HVT U199 ( .A1(n125), .A2(DP_OP_422J2_124_3477_n88), .A3(
        DP_OP_422J2_124_3477_n93), .A4(n126), .Y(n129) );
  NAND2X0_HVT U200 ( .A1(n127), .A2(n129), .Y(n_conv2_sum_a[11]) );
  OA21X1_HVT U201 ( .A1(DP_OP_422J2_124_3477_n55), .A2(
        DP_OP_422J2_124_3477_n73), .A3(DP_OP_422J2_124_3477_n56), .Y(n130) );
  INVX0_HVT U202 ( .A(DP_OP_422J2_124_3477_n52), .Y(n131) );
  NAND2X0_HVT U203 ( .A1(n131), .A2(DP_OP_422J2_124_3477_n53), .Y(n132) );
  HADDX1_HVT U204 ( .A0(n130), .B0(n132), .SO(n_conv2_sum_a[17]) );
  INVX0_HVT U205 ( .A(DP_OP_425J2_127_3477_n105), .Y(n133) );
  NAND2X0_HVT U206 ( .A1(n133), .A2(DP_OP_425J2_127_3477_n106), .Y(n134) );
  HADDX1_HVT U207 ( .A0(DP_OP_425J2_127_3477_n107), .B0(n134), .SO(
        n_conv2_sum_d[7]) );
  INVX0_HVT U208 ( .A(DP_OP_425J2_127_3477_n87), .Y(n135) );
  NAND2X0_HVT U209 ( .A1(DP_OP_425J2_127_3477_n94), .A2(
        DP_OP_425J2_127_3477_n90), .Y(n136) );
  AO22X1_HVT U210 ( .A1(n135), .A2(DP_OP_425J2_127_3477_n88), .A3(
        DP_OP_425J2_127_3477_n93), .A4(n136), .Y(n137) );
  NAND4X0_HVT U211 ( .A1(n135), .A2(DP_OP_425J2_127_3477_n88), .A3(
        DP_OP_425J2_127_3477_n93), .A4(n136), .Y(n138) );
  NAND2X0_HVT U212 ( .A1(n137), .A2(n138), .Y(n_conv2_sum_d[11]) );
  OA21X1_HVT U213 ( .A1(DP_OP_425J2_127_3477_n55), .A2(
        DP_OP_425J2_127_3477_n73), .A3(DP_OP_425J2_127_3477_n56), .Y(n139) );
  INVX0_HVT U214 ( .A(DP_OP_425J2_127_3477_n52), .Y(n140) );
  NAND2X0_HVT U215 ( .A1(n140), .A2(DP_OP_425J2_127_3477_n53), .Y(n141) );
  HADDX1_HVT U216 ( .A0(n139), .B0(n141), .SO(n_conv2_sum_d[17]) );
  INVX0_HVT U217 ( .A(DP_OP_424J2_126_3477_n105), .Y(n142) );
  NAND2X0_HVT U218 ( .A1(n142), .A2(DP_OP_424J2_126_3477_n106), .Y(n143) );
  HADDX1_HVT U219 ( .A0(DP_OP_424J2_126_3477_n107), .B0(n143), .SO(
        n_conv2_sum_c[7]) );
  INVX0_HVT U220 ( .A(DP_OP_424J2_126_3477_n87), .Y(n144) );
  NAND2X0_HVT U221 ( .A1(DP_OP_424J2_126_3477_n94), .A2(
        DP_OP_424J2_126_3477_n90), .Y(n145) );
  AO22X1_HVT U222 ( .A1(n144), .A2(DP_OP_424J2_126_3477_n88), .A3(
        DP_OP_424J2_126_3477_n93), .A4(n145), .Y(n146) );
  NAND4X0_HVT U223 ( .A1(n144), .A2(DP_OP_424J2_126_3477_n88), .A3(
        DP_OP_424J2_126_3477_n93), .A4(n145), .Y(n147) );
  NAND2X0_HVT U224 ( .A1(n146), .A2(n147), .Y(n_conv2_sum_c[11]) );
  OA21X1_HVT U225 ( .A1(DP_OP_424J2_126_3477_n55), .A2(
        DP_OP_424J2_126_3477_n73), .A3(DP_OP_424J2_126_3477_n56), .Y(n148) );
  INVX0_HVT U226 ( .A(DP_OP_424J2_126_3477_n52), .Y(n149) );
  NAND2X0_HVT U227 ( .A1(n149), .A2(DP_OP_424J2_126_3477_n53), .Y(n150) );
  HADDX1_HVT U228 ( .A0(n148), .B0(n150), .SO(n_conv2_sum_c[17]) );
  INVX0_HVT U229 ( .A(n332), .Y(n151) );
  AOI22X1_HVT U230 ( .A1(n332), .A2(conv1_sram_rdata_weight[46]), .A3(n151), 
        .A4(conv2_sram_rdata_weight[46]), .Y(n447) );
  INVX0_HVT U231 ( .A(n351), .Y(n152) );
  AOI22X1_HVT U232 ( .A1(n351), .A2(conv1_sram_rdata_weight[13]), .A3(n152), 
        .A4(conv2_sram_rdata_weight[13]), .Y(n449) );
  INVX0_HVT U233 ( .A(n350), .Y(n153) );
  AOI22X1_HVT U234 ( .A1(n350), .A2(conv1_sram_rdata_weight[44]), .A3(n153), 
        .A4(conv2_sram_rdata_weight[44]), .Y(n441) );
  NAND3X0_HVT U235 ( .A1(n522), .A2(n524), .A3(n523), .Y(n154) );
  OA21X1_HVT U236 ( .A1(n465), .A2(n459), .A3(n460), .Y(n155) );
  OA22X1_HVT U237 ( .A1(n420), .A2(conv2_sum_b[29]), .A3(n454), .A4(
        conv2_sum_b[28]), .Y(n156) );
  OA22X1_HVT U238 ( .A1(conv2_sum_a[31]), .A2(n380), .A3(n463), .A4(n156), .Y(
        n157) );
  OA221X1_HVT U239 ( .A1(n154), .A2(conv2_sum_b[24]), .A3(n154), .A4(n418), 
        .A5(n158), .Y(N5) );
  INVX0_HVT U240 ( .A(DP_OP_423J2_125_3477_n119), .Y(n159) );
  NAND2X0_HVT U241 ( .A1(n159), .A2(DP_OP_423J2_125_3477_n120), .Y(n160) );
  HADDX1_HVT U242 ( .A0(DP_OP_423J2_125_3477_n121), .B0(n160), .SO(
        n_conv2_sum_b[3]) );
  INVX0_HVT U243 ( .A(DP_OP_423J2_125_3477_n111), .Y(n161) );
  NAND2X0_HVT U244 ( .A1(n161), .A2(DP_OP_423J2_125_3477_n112), .Y(n162) );
  HADDX1_HVT U245 ( .A0(DP_OP_423J2_125_3477_n113), .B0(n162), .SO(
        n_conv2_sum_b[5]) );
  INVX0_HVT U246 ( .A(DP_OP_423J2_125_3477_n99), .Y(n163) );
  NAND2X0_HVT U247 ( .A1(n163), .A2(DP_OP_423J2_125_3477_n100), .Y(n164) );
  HADDX1_HVT U248 ( .A0(DP_OP_423J2_125_3477_n101), .B0(n164), .SO(
        n_conv2_sum_b[8]) );
  INVX0_HVT U249 ( .A(DP_OP_423J2_125_3477_n80), .Y(n165) );
  NAND2X0_HVT U250 ( .A1(n165), .A2(DP_OP_423J2_125_3477_n81), .Y(n166) );
  HADDX1_HVT U251 ( .A0(DP_OP_423J2_125_3477_n82), .B0(n166), .SO(
        n_conv2_sum_b[12]) );
  INVX0_HVT U252 ( .A(DP_OP_423J2_125_3477_n71), .Y(n167) );
  AOI21X1_HVT U253 ( .A1(DP_OP_423J2_125_3477_n48), .A2(n167), .A3(
        DP_OP_423J2_125_3477_n49), .Y(n168) );
  NAND2X0_HVT U254 ( .A1(DP_OP_423J2_125_3477_n43), .A2(
        DP_OP_423J2_125_3477_n44), .Y(n169) );
  HADDX1_HVT U255 ( .A0(n168), .B0(n169), .SO(n_conv2_sum_b[18]) );
  INVX0_HVT U256 ( .A(DP_OP_422J2_124_3477_n129), .Y(n170) );
  AND2X1_HVT U257 ( .A1(n170), .A2(DP_OP_422J2_124_3477_n130), .Y(n171) );
  HADDX1_HVT U258 ( .A0(n171), .B0(DP_OP_422J2_124_3477_n131), .SO(
        n_conv2_sum_a[1]) );
  INVX0_HVT U259 ( .A(DP_OP_422J2_124_3477_n121), .Y(n172) );
  NAND2X0_HVT U260 ( .A1(n172), .A2(DP_OP_422J2_124_3477_n122), .Y(n173) );
  HADDX1_HVT U261 ( .A0(DP_OP_422J2_124_3477_n123), .B0(n173), .SO(
        n_conv2_sum_a[3]) );
  INVX0_HVT U262 ( .A(DP_OP_422J2_124_3477_n113), .Y(n174) );
  NAND2X0_HVT U263 ( .A1(n174), .A2(DP_OP_422J2_124_3477_n114), .Y(n175) );
  HADDX1_HVT U264 ( .A0(DP_OP_422J2_124_3477_n115), .B0(n175), .SO(
        n_conv2_sum_a[5]) );
  INVX0_HVT U265 ( .A(DP_OP_422J2_124_3477_n101), .Y(n176) );
  NAND2X0_HVT U266 ( .A1(n176), .A2(DP_OP_422J2_124_3477_n102), .Y(n177) );
  HADDX1_HVT U267 ( .A0(DP_OP_422J2_124_3477_n103), .B0(n177), .SO(
        n_conv2_sum_a[8]) );
  INVX0_HVT U268 ( .A(DP_OP_422J2_124_3477_n82), .Y(n178) );
  NAND2X0_HVT U269 ( .A1(n178), .A2(DP_OP_422J2_124_3477_n83), .Y(n179) );
  HADDX1_HVT U270 ( .A0(DP_OP_422J2_124_3477_n84), .B0(n179), .SO(
        n_conv2_sum_a[12]) );
  INVX0_HVT U271 ( .A(DP_OP_422J2_124_3477_n73), .Y(n180) );
  AOI21X1_HVT U272 ( .A1(DP_OP_422J2_124_3477_n50), .A2(n180), .A3(
        DP_OP_422J2_124_3477_n51), .Y(n181) );
  NAND2X0_HVT U273 ( .A1(DP_OP_422J2_124_3477_n45), .A2(
        DP_OP_422J2_124_3477_n46), .Y(n182) );
  HADDX1_HVT U274 ( .A0(n181), .B0(n182), .SO(n_conv2_sum_a[18]) );
  INVX0_HVT U275 ( .A(DP_OP_425J2_127_3477_n129), .Y(n183) );
  AND2X1_HVT U276 ( .A1(n183), .A2(DP_OP_425J2_127_3477_n130), .Y(n184) );
  HADDX1_HVT U277 ( .A0(n184), .B0(DP_OP_425J2_127_3477_n131), .SO(
        n_conv2_sum_d[1]) );
  INVX0_HVT U278 ( .A(DP_OP_425J2_127_3477_n121), .Y(n185) );
  NAND2X0_HVT U279 ( .A1(n185), .A2(DP_OP_425J2_127_3477_n122), .Y(n186) );
  HADDX1_HVT U280 ( .A0(DP_OP_425J2_127_3477_n123), .B0(n186), .SO(
        n_conv2_sum_d[3]) );
  INVX0_HVT U281 ( .A(DP_OP_425J2_127_3477_n113), .Y(n187) );
  NAND2X0_HVT U282 ( .A1(n187), .A2(DP_OP_425J2_127_3477_n114), .Y(n188) );
  HADDX1_HVT U283 ( .A0(DP_OP_425J2_127_3477_n115), .B0(n188), .SO(
        n_conv2_sum_d[5]) );
  INVX0_HVT U284 ( .A(DP_OP_425J2_127_3477_n101), .Y(n189) );
  NAND2X0_HVT U285 ( .A1(n189), .A2(DP_OP_425J2_127_3477_n102), .Y(n190) );
  HADDX1_HVT U286 ( .A0(DP_OP_425J2_127_3477_n103), .B0(n190), .SO(
        n_conv2_sum_d[8]) );
  INVX0_HVT U287 ( .A(DP_OP_425J2_127_3477_n82), .Y(n191) );
  NAND2X0_HVT U288 ( .A1(n191), .A2(DP_OP_425J2_127_3477_n83), .Y(n192) );
  HADDX1_HVT U289 ( .A0(DP_OP_425J2_127_3477_n84), .B0(n192), .SO(
        n_conv2_sum_d[12]) );
  INVX0_HVT U290 ( .A(DP_OP_425J2_127_3477_n73), .Y(n193) );
  AOI21X1_HVT U291 ( .A1(DP_OP_425J2_127_3477_n50), .A2(n193), .A3(
        DP_OP_425J2_127_3477_n51), .Y(n194) );
  NAND2X0_HVT U292 ( .A1(DP_OP_425J2_127_3477_n45), .A2(
        DP_OP_425J2_127_3477_n46), .Y(n195) );
  HADDX1_HVT U293 ( .A0(n194), .B0(n195), .SO(n_conv2_sum_d[18]) );
  INVX0_HVT U294 ( .A(DP_OP_424J2_126_3477_n129), .Y(n196) );
  AND2X1_HVT U295 ( .A1(n196), .A2(DP_OP_424J2_126_3477_n130), .Y(n197) );
  HADDX1_HVT U296 ( .A0(n197), .B0(DP_OP_424J2_126_3477_n131), .SO(
        n_conv2_sum_c[1]) );
  INVX0_HVT U297 ( .A(DP_OP_424J2_126_3477_n121), .Y(n198) );
  NAND2X0_HVT U298 ( .A1(n198), .A2(DP_OP_424J2_126_3477_n122), .Y(n199) );
  HADDX1_HVT U299 ( .A0(DP_OP_424J2_126_3477_n123), .B0(n199), .SO(
        n_conv2_sum_c[3]) );
  INVX0_HVT U300 ( .A(DP_OP_424J2_126_3477_n113), .Y(n200) );
  NAND2X0_HVT U301 ( .A1(n200), .A2(DP_OP_424J2_126_3477_n114), .Y(n201) );
  HADDX1_HVT U302 ( .A0(DP_OP_424J2_126_3477_n115), .B0(n201), .SO(
        n_conv2_sum_c[5]) );
  INVX0_HVT U303 ( .A(DP_OP_424J2_126_3477_n101), .Y(n202) );
  NAND2X0_HVT U304 ( .A1(n202), .A2(DP_OP_424J2_126_3477_n102), .Y(n203) );
  HADDX1_HVT U305 ( .A0(DP_OP_424J2_126_3477_n103), .B0(n203), .SO(
        n_conv2_sum_c[8]) );
  INVX0_HVT U306 ( .A(DP_OP_424J2_126_3477_n82), .Y(n204) );
  NAND2X0_HVT U307 ( .A1(n204), .A2(DP_OP_424J2_126_3477_n83), .Y(n205) );
  HADDX1_HVT U308 ( .A0(DP_OP_424J2_126_3477_n84), .B0(n205), .SO(
        n_conv2_sum_c[12]) );
  INVX0_HVT U309 ( .A(DP_OP_424J2_126_3477_n73), .Y(n206) );
  AOI21X1_HVT U310 ( .A1(DP_OP_424J2_126_3477_n50), .A2(n206), .A3(
        DP_OP_424J2_126_3477_n51), .Y(n207) );
  NAND2X0_HVT U311 ( .A1(DP_OP_424J2_126_3477_n45), .A2(
        DP_OP_424J2_126_3477_n46), .Y(n208) );
  HADDX1_HVT U312 ( .A0(n207), .B0(n208), .SO(n_conv2_sum_c[18]) );
  INVX0_HVT U313 ( .A(n332), .Y(n209) );
  AOI22X1_HVT U314 ( .A1(n332), .A2(conv1_sram_rdata_weight[94]), .A3(n209), 
        .A4(conv2_sram_rdata_weight[94]), .Y(n448) );
  INVX0_HVT U316 ( .A(n541), .Y(n211) );
  INVX0_HVT U317 ( .A(n352), .Y(n212) );
  AOI22X1_HVT U318 ( .A1(n352), .A2(conv1_sram_rdata_weight[53]), .A3(n212), 
        .A4(conv2_sram_rdata_weight[53]), .Y(n440) );
  INVX0_HVT U319 ( .A(n350), .Y(n213) );
  AOI22X1_HVT U320 ( .A1(n350), .A2(conv1_sram_rdata_weight[84]), .A3(n213), 
        .A4(conv2_sram_rdata_weight[84]), .Y(n446) );
  INVX0_HVT U321 ( .A(n526), .Y(n214) );
  AND2X1_HVT U323 ( .A1(DP_OP_423J2_125_3477_n125), .A2(
        DP_OP_423J2_125_3477_n124), .Y(n216) );
  HADDX1_HVT U324 ( .A0(n216), .B0(DP_OP_423J2_125_3477_n126), .SO(
        n_conv2_sum_b[2]) );
  AND2X1_HVT U325 ( .A1(DP_OP_423J2_125_3477_n117), .A2(
        DP_OP_423J2_125_3477_n116), .Y(n217) );
  HADDX1_HVT U326 ( .A0(n217), .B0(DP_OP_423J2_125_3477_n118), .SO(
        n_conv2_sum_b[4]) );
  AND2X1_HVT U327 ( .A1(DP_OP_423J2_125_3477_n109), .A2(
        DP_OP_423J2_125_3477_n108), .Y(n218) );
  HADDX1_HVT U328 ( .A0(n218), .B0(DP_OP_423J2_125_3477_n110), .SO(
        n_conv2_sum_b[6]) );
  OA21X1_HVT U329 ( .A1(DP_OP_423J2_125_3477_n99), .A2(
        DP_OP_423J2_125_3477_n101), .A3(DP_OP_423J2_125_3477_n100), .Y(n219)
         );
  INVX0_HVT U330 ( .A(DP_OP_423J2_125_3477_n96), .Y(n220) );
  NAND2X0_HVT U331 ( .A1(n220), .A2(DP_OP_423J2_125_3477_n97), .Y(n221) );
  HADDX1_HVT U332 ( .A0(n219), .B0(n221), .SO(n_conv2_sum_b[9]) );
  OA21X1_HVT U333 ( .A1(DP_OP_423J2_125_3477_n80), .A2(
        DP_OP_423J2_125_3477_n82), .A3(DP_OP_423J2_125_3477_n81), .Y(n222) );
  INVX0_HVT U334 ( .A(DP_OP_423J2_125_3477_n77), .Y(n223) );
  NAND2X0_HVT U335 ( .A1(n223), .A2(DP_OP_423J2_125_3477_n78), .Y(n224) );
  HADDX1_HVT U336 ( .A0(n222), .B0(n224), .SO(n_conv2_sum_b[13]) );
  OA21X1_HVT U337 ( .A1(DP_OP_423J2_125_3477_n39), .A2(
        DP_OP_423J2_125_3477_n71), .A3(DP_OP_423J2_125_3477_n40), .Y(n225) );
  INVX0_HVT U338 ( .A(DP_OP_423J2_125_3477_n36), .Y(n226) );
  NAND2X0_HVT U339 ( .A1(n226), .A2(DP_OP_423J2_125_3477_n37), .Y(n227) );
  HADDX1_HVT U340 ( .A0(n225), .B0(n227), .SO(n_conv2_sum_b[19]) );
  AND2X1_HVT U341 ( .A1(DP_OP_422J2_124_3477_n127), .A2(
        DP_OP_422J2_124_3477_n126), .Y(n228) );
  HADDX1_HVT U342 ( .A0(n228), .B0(DP_OP_422J2_124_3477_n128), .SO(
        n_conv2_sum_a[2]) );
  AND2X1_HVT U343 ( .A1(DP_OP_422J2_124_3477_n119), .A2(
        DP_OP_422J2_124_3477_n118), .Y(n229) );
  HADDX1_HVT U344 ( .A0(n229), .B0(DP_OP_422J2_124_3477_n120), .SO(
        n_conv2_sum_a[4]) );
  AND2X1_HVT U345 ( .A1(DP_OP_422J2_124_3477_n111), .A2(
        DP_OP_422J2_124_3477_n110), .Y(n230) );
  HADDX1_HVT U346 ( .A0(n230), .B0(DP_OP_422J2_124_3477_n112), .SO(
        n_conv2_sum_a[6]) );
  OA21X1_HVT U347 ( .A1(DP_OP_422J2_124_3477_n101), .A2(
        DP_OP_422J2_124_3477_n103), .A3(DP_OP_422J2_124_3477_n102), .Y(n231)
         );
  INVX0_HVT U348 ( .A(DP_OP_422J2_124_3477_n98), .Y(n232) );
  NAND2X0_HVT U349 ( .A1(n232), .A2(DP_OP_422J2_124_3477_n99), .Y(n233) );
  HADDX1_HVT U350 ( .A0(n231), .B0(n233), .SO(n_conv2_sum_a[9]) );
  OA21X1_HVT U351 ( .A1(DP_OP_422J2_124_3477_n82), .A2(
        DP_OP_422J2_124_3477_n84), .A3(DP_OP_422J2_124_3477_n83), .Y(n234) );
  INVX0_HVT U352 ( .A(DP_OP_422J2_124_3477_n79), .Y(n235) );
  NAND2X0_HVT U353 ( .A1(n235), .A2(DP_OP_422J2_124_3477_n80), .Y(n236) );
  HADDX1_HVT U354 ( .A0(n234), .B0(n236), .SO(n_conv2_sum_a[13]) );
  OA21X1_HVT U355 ( .A1(DP_OP_422J2_124_3477_n41), .A2(
        DP_OP_422J2_124_3477_n73), .A3(DP_OP_422J2_124_3477_n42), .Y(n237) );
  INVX0_HVT U356 ( .A(DP_OP_422J2_124_3477_n38), .Y(n238) );
  NAND2X0_HVT U357 ( .A1(n238), .A2(DP_OP_422J2_124_3477_n39), .Y(n239) );
  HADDX1_HVT U358 ( .A0(n237), .B0(n239), .SO(n_conv2_sum_a[19]) );
  AND2X1_HVT U359 ( .A1(DP_OP_425J2_127_3477_n127), .A2(
        DP_OP_425J2_127_3477_n126), .Y(n240) );
  HADDX1_HVT U360 ( .A0(n240), .B0(DP_OP_425J2_127_3477_n128), .SO(
        n_conv2_sum_d[2]) );
  AND2X1_HVT U361 ( .A1(DP_OP_425J2_127_3477_n119), .A2(
        DP_OP_425J2_127_3477_n118), .Y(n241) );
  HADDX1_HVT U362 ( .A0(n241), .B0(DP_OP_425J2_127_3477_n120), .SO(
        n_conv2_sum_d[4]) );
  AND2X1_HVT U363 ( .A1(DP_OP_425J2_127_3477_n111), .A2(
        DP_OP_425J2_127_3477_n110), .Y(n242) );
  HADDX1_HVT U364 ( .A0(n242), .B0(DP_OP_425J2_127_3477_n112), .SO(
        n_conv2_sum_d[6]) );
  OA21X1_HVT U365 ( .A1(DP_OP_425J2_127_3477_n101), .A2(
        DP_OP_425J2_127_3477_n103), .A3(DP_OP_425J2_127_3477_n102), .Y(n243)
         );
  INVX0_HVT U366 ( .A(DP_OP_425J2_127_3477_n98), .Y(n244) );
  NAND2X0_HVT U367 ( .A1(n244), .A2(DP_OP_425J2_127_3477_n99), .Y(n245) );
  HADDX1_HVT U368 ( .A0(n243), .B0(n245), .SO(n_conv2_sum_d[9]) );
  OA21X1_HVT U369 ( .A1(DP_OP_425J2_127_3477_n82), .A2(
        DP_OP_425J2_127_3477_n84), .A3(DP_OP_425J2_127_3477_n83), .Y(n246) );
  INVX0_HVT U370 ( .A(DP_OP_425J2_127_3477_n79), .Y(n247) );
  NAND2X0_HVT U371 ( .A1(n247), .A2(DP_OP_425J2_127_3477_n80), .Y(n248) );
  HADDX1_HVT U372 ( .A0(n246), .B0(n248), .SO(n_conv2_sum_d[13]) );
  OA21X1_HVT U373 ( .A1(DP_OP_425J2_127_3477_n41), .A2(
        DP_OP_425J2_127_3477_n73), .A3(DP_OP_425J2_127_3477_n42), .Y(n249) );
  INVX0_HVT U374 ( .A(DP_OP_425J2_127_3477_n38), .Y(n250) );
  NAND2X0_HVT U375 ( .A1(n250), .A2(DP_OP_425J2_127_3477_n39), .Y(n251) );
  HADDX1_HVT U376 ( .A0(n249), .B0(n251), .SO(n_conv2_sum_d[19]) );
  AND2X1_HVT U377 ( .A1(DP_OP_424J2_126_3477_n127), .A2(
        DP_OP_424J2_126_3477_n126), .Y(n252) );
  HADDX1_HVT U378 ( .A0(n252), .B0(DP_OP_424J2_126_3477_n128), .SO(
        n_conv2_sum_c[2]) );
  AND2X1_HVT U379 ( .A1(DP_OP_424J2_126_3477_n119), .A2(
        DP_OP_424J2_126_3477_n118), .Y(n253) );
  HADDX1_HVT U380 ( .A0(n253), .B0(DP_OP_424J2_126_3477_n120), .SO(
        n_conv2_sum_c[4]) );
  AND2X1_HVT U381 ( .A1(DP_OP_424J2_126_3477_n111), .A2(
        DP_OP_424J2_126_3477_n110), .Y(n254) );
  HADDX1_HVT U382 ( .A0(n254), .B0(DP_OP_424J2_126_3477_n112), .SO(
        n_conv2_sum_c[6]) );
  OA21X1_HVT U383 ( .A1(DP_OP_424J2_126_3477_n101), .A2(
        DP_OP_424J2_126_3477_n103), .A3(DP_OP_424J2_126_3477_n102), .Y(n255)
         );
  INVX0_HVT U384 ( .A(DP_OP_424J2_126_3477_n98), .Y(n256) );
  NAND2X0_HVT U385 ( .A1(n256), .A2(DP_OP_424J2_126_3477_n99), .Y(n257) );
  HADDX1_HVT U386 ( .A0(n255), .B0(n257), .SO(n_conv2_sum_c[9]) );
  OA21X1_HVT U387 ( .A1(DP_OP_424J2_126_3477_n82), .A2(
        DP_OP_424J2_126_3477_n84), .A3(DP_OP_424J2_126_3477_n83), .Y(n258) );
  INVX0_HVT U388 ( .A(DP_OP_424J2_126_3477_n79), .Y(n259) );
  NAND2X0_HVT U389 ( .A1(n259), .A2(DP_OP_424J2_126_3477_n80), .Y(n260) );
  HADDX1_HVT U390 ( .A0(n258), .B0(n260), .SO(n_conv2_sum_c[13]) );
  OA21X1_HVT U391 ( .A1(DP_OP_424J2_126_3477_n41), .A2(
        DP_OP_424J2_126_3477_n73), .A3(DP_OP_424J2_126_3477_n42), .Y(n261) );
  INVX0_HVT U392 ( .A(DP_OP_424J2_126_3477_n38), .Y(n262) );
  NAND2X0_HVT U393 ( .A1(n262), .A2(DP_OP_424J2_126_3477_n39), .Y(n263) );
  HADDX1_HVT U394 ( .A0(n261), .B0(n263), .SO(n_conv2_sum_c[19]) );
  AND2X1_HVT U395 ( .A1(mode[1]), .A2(n687), .Y(n453) );
  INVX1_HVT U396 ( .A(tmp_big1[26]), .Y(n677) );
  INVX1_HVT U397 ( .A(tmp_big2[8]), .Y(n663) );
  INVX1_HVT U398 ( .A(n443), .Y(conv_weight_box[66]) );
  NAND2X0_HVT U399 ( .A1(n436), .A2(n435), .Y(DP_OP_425J2_127_3477_n3255) );
  INVX1_HVT U400 ( .A(n442), .Y(conv_weight_box[20]) );
  INVX1_HVT U401 ( .A(n437), .Y(n341) );
  INVX1_HVT U402 ( .A(n437), .Y(n340) );
  INVX1_HVT U403 ( .A(n437), .Y(n342) );
  INVX1_HVT U404 ( .A(n437), .Y(n343) );
  INVX1_HVT U405 ( .A(n437), .Y(n339) );
  AO22X1_HVT U406 ( .A1(n334), .A2(conv1_sram_rdata_weight[33]), .A3(n438), 
        .A4(conv2_sram_rdata_weight[33]), .Y(n428) );
  INVX1_HVT U407 ( .A(n447), .Y(conv_weight_box[42]) );
  INVX1_HVT U408 ( .A(n448), .Y(conv_weight_box[89]) );
  AO22X1_HVT U409 ( .A1(n332), .A2(conv1_sram_rdata_weight[96]), .A3(n438), 
        .A4(conv2_sram_rdata_weight[96]), .Y(n430) );
  AO22X1_HVT U410 ( .A1(n333), .A2(conv1_sram_rdata_weight[14]), .A3(n438), 
        .A4(conv2_sram_rdata_weight[14]), .Y(n431) );
  INVX1_HVT U411 ( .A(n437), .Y(DP_OP_425J2_127_3477_n2) );
  INVX1_HVT U412 ( .A(n451), .Y(conv_weight_box[54]) );
  INVX1_HVT U413 ( .A(n437), .Y(DP_OP_424J2_126_3477_n2) );
  INVX1_HVT U414 ( .A(n437), .Y(DP_OP_423J2_125_3477_n2) );
  INVX1_HVT U415 ( .A(n438), .Y(n333) );
  INVX1_HVT U416 ( .A(n438), .Y(n332) );
  INVX1_HVT U417 ( .A(srstn), .Y(n330) );
  INVX0_HVT U418 ( .A(DP_OP_424J2_126_3477_n95), .Y(DP_OP_424J2_126_3477_n94)
         );
  INVX0_HVT U419 ( .A(DP_OP_425J2_127_3477_n95), .Y(DP_OP_425J2_127_3477_n94)
         );
  INVX0_HVT U420 ( .A(DP_OP_422J2_124_3477_n95), .Y(DP_OP_422J2_124_3477_n94)
         );
  INVX0_HVT U421 ( .A(DP_OP_423J2_125_3477_n93), .Y(DP_OP_423J2_125_3477_n92)
         );
  INVX0_HVT U422 ( .A(DP_OP_425J2_127_3477_n104), .Y(DP_OP_425J2_127_3477_n103) );
  INVX0_HVT U423 ( .A(DP_OP_424J2_126_3477_n104), .Y(DP_OP_424J2_126_3477_n103) );
  INVX0_HVT U424 ( .A(DP_OP_425J2_127_3477_n92), .Y(DP_OP_425J2_127_3477_n90)
         );
  INVX0_HVT U425 ( .A(DP_OP_422J2_124_3477_n104), .Y(DP_OP_422J2_124_3477_n103) );
  INVX0_HVT U426 ( .A(DP_OP_423J2_125_3477_n102), .Y(DP_OP_423J2_125_3477_n101) );
  INVX0_HVT U427 ( .A(DP_OP_424J2_126_3477_n92), .Y(DP_OP_424J2_126_3477_n90)
         );
  INVX0_HVT U428 ( .A(DP_OP_422J2_124_3477_n92), .Y(DP_OP_422J2_124_3477_n90)
         );
  INVX0_HVT U429 ( .A(DP_OP_423J2_125_3477_n90), .Y(DP_OP_423J2_125_3477_n88)
         );
  INVX0_HVT U430 ( .A(DP_OP_422J2_124_3477_n64), .Y(DP_OP_422J2_124_3477_n62)
         );
  INVX0_HVT U431 ( .A(DP_OP_425J2_127_3477_n64), .Y(DP_OP_425J2_127_3477_n62)
         );
  INVX0_HVT U432 ( .A(DP_OP_423J2_125_3477_n62), .Y(DP_OP_423J2_125_3477_n60)
         );
  INVX0_HVT U433 ( .A(DP_OP_424J2_126_3477_n64), .Y(DP_OP_424J2_126_3477_n62)
         );
  MUX21X1_HVT U434 ( .A1(tmp_big2[18]), .A2(tmp_big1[18]), .S0(n355), .Y(
        data_out[18]) );
  MUX21X1_HVT U435 ( .A1(tmp_big2[19]), .A2(tmp_big1[19]), .S0(n356), .Y(
        data_out[19]) );
  INVX1_HVT U436 ( .A(N9), .Y(n355) );
  INVX1_HVT U437 ( .A(N9), .Y(n354) );
  INVX1_HVT U438 ( .A(N9), .Y(n356) );
  INVX1_HVT U439 ( .A(N9), .Y(n357) );
  INVX0_HVT U440 ( .A(DP_OP_425J2_127_3477_n131), .Y(DP_OP_425J2_127_3477_n4)
         );
  NOR2X1_HVT U441 ( .A1(n609), .A2(n608), .Y(n655) );
  INVX0_HVT U442 ( .A(DP_OP_422J2_124_3477_n131), .Y(DP_OP_422J2_124_3477_n4)
         );
  INVX0_HVT U443 ( .A(DP_OP_424J2_126_3477_n131), .Y(DP_OP_424J2_126_3477_n4)
         );
  INVX0_HVT U444 ( .A(tmp_big1[4]), .Y(n683) );
  INVX0_HVT U445 ( .A(tmp_big1[2]), .Y(n680) );
  INVX0_HVT U446 ( .A(tmp_big1[10]), .Y(n664) );
  INVX0_HVT U447 ( .A(tmp_big1[22]), .Y(n673) );
  INVX0_HVT U448 ( .A(tmp_big2[16]), .Y(n660) );
  INVX0_HVT U449 ( .A(tmp_big1[18]), .Y(n670) );
  INVX1_HVT U450 ( .A(N5), .Y(n365) );
  INVX1_HVT U451 ( .A(N7), .Y(n361) );
  INVX1_HVT U452 ( .A(N7), .Y(n360) );
  INVX1_HVT U453 ( .A(N7), .Y(n358) );
  INVX1_HVT U454 ( .A(N5), .Y(n364) );
  INVX1_HVT U455 ( .A(N5), .Y(n362) );
  INVX1_HVT U456 ( .A(N5), .Y(n363) );
  INVX1_HVT U457 ( .A(N7), .Y(n359) );
  AO22X1_HVT U458 ( .A1(n333), .A2(conv1_sram_rdata_weight[0]), .A3(n438), 
        .A4(conv2_sram_rdata_weight[0]), .Y(n429) );
  MUX21X1_HVT U459 ( .A1(conv2_sram_rdata_weight[6]), .A2(
        conv1_sram_rdata_weight[6]), .S0(n333), .Y(conv_weight_box[5]) );
  MUX21X1_HVT U460 ( .A1(conv2_sram_rdata_weight[82]), .A2(
        conv1_sram_rdata_weight[82]), .S0(n333), .Y(conv_weight_box[78]) );
  NAND2X0_HVT U461 ( .A1(n434), .A2(n433), .Y(conv_weight_box[77]) );
  MUX21X1_HVT U462 ( .A1(conv2_sram_rdata_weight[78]), .A2(
        conv1_sram_rdata_weight[78]), .S0(n334), .Y(conv_weight_box[74]) );
  MUX21X1_HVT U463 ( .A1(conv2_sram_rdata_weight[54]), .A2(
        conv1_sram_rdata_weight[54]), .S0(n334), .Y(conv_weight_box[50]) );
  MUX21X1_HVT U464 ( .A1(conv2_sram_rdata_weight[27]), .A2(
        conv1_sram_rdata_weight[27]), .S0(n333), .Y(conv_weight_box[25]) );
  MUX21X1_HVT U465 ( .A1(conv2_sram_rdata_weight[31]), .A2(
        conv1_sram_rdata_weight[31]), .S0(n332), .Y(conv_weight_box[29]) );
  MUX21X1_HVT U466 ( .A1(conv2_sram_rdata_weight[24]), .A2(
        conv1_sram_rdata_weight[24]), .S0(n332), .Y(conv_weight_box[22]) );
  MUX21X1_HVT U467 ( .A1(conv2_sram_rdata_weight[8]), .A2(
        conv1_sram_rdata_weight[8]), .S0(n333), .Y(conv_weight_box[7]) );
  MUX21X1_HVT U468 ( .A1(conv2_sram_rdata_weight[12]), .A2(
        conv1_sram_rdata_weight[12]), .S0(n334), .Y(conv_weight_box[11]) );
  MUX21X1_HVT U469 ( .A1(conv2_sram_rdata_weight[72]), .A2(
        conv1_sram_rdata_weight[72]), .S0(n333), .Y(conv_weight_box[68]) );
  MUX21X1_HVT U470 ( .A1(conv2_sram_rdata_weight[36]), .A2(
        conv1_sram_rdata_weight[36]), .S0(n335), .Y(conv_weight_box[33]) );
  MUX21X1_HVT U471 ( .A1(conv2_sram_rdata_weight[40]), .A2(
        conv1_sram_rdata_weight[40]), .S0(n336), .Y(conv_weight_box[37]) );
  INVX1_HVT U472 ( .A(n441), .Y(conv_weight_box[40]) );
  MUX21X1_HVT U473 ( .A1(conv2_sram_rdata_weight[43]), .A2(
        conv1_sram_rdata_weight[43]), .S0(n335), .Y(conv_weight_box[39]) );
  MUX21X1_HVT U474 ( .A1(conv2_sram_rdata_weight[15]), .A2(
        conv1_sram_rdata_weight[15]), .S0(n353), .Y(conv_weight_box[13]) );
  MUX21X1_HVT U475 ( .A1(conv1_sram_rdata_weight[76]), .A2(
        conv2_sram_rdata_weight[76]), .S0(n453), .Y(conv_weight_box[72]) );
  MUX21X1_HVT U476 ( .A1(conv2_sram_rdata_weight[19]), .A2(
        conv1_sram_rdata_weight[19]), .S0(n334), .Y(conv_weight_box[17]) );
  MUX21X1_HVT U477 ( .A1(conv2_sram_rdata_weight[55]), .A2(
        conv1_sram_rdata_weight[55]), .S0(n334), .Y(conv_weight_box[51]) );
  INVX1_HVT U478 ( .A(n444), .Y(conv_weight_box[70]) );
  MUX21X1_HVT U479 ( .A1(conv2_sram_rdata_weight[28]), .A2(
        conv1_sram_rdata_weight[28]), .S0(n335), .Y(conv_weight_box[26]) );
  MUX21X1_HVT U480 ( .A1(conv2_sram_rdata_weight[7]), .A2(
        conv1_sram_rdata_weight[7]), .S0(n336), .Y(conv_weight_box[6]) );
  INVX1_HVT U481 ( .A(n445), .Y(conv_weight_box[82]) );
  INVX1_HVT U482 ( .A(n446), .Y(conv_weight_box[80]) );
  INVX1_HVT U483 ( .A(n452), .Y(conv_weight_box[58]) );
  MUX21X1_HVT U484 ( .A1(conv2_sram_rdata_weight[11]), .A2(
        conv1_sram_rdata_weight[11]), .S0(n335), .Y(conv_weight_box[10]) );
  MUX21X1_HVT U485 ( .A1(conv2_sram_rdata_weight[63]), .A2(
        conv1_sram_rdata_weight[63]), .S0(n335), .Y(conv_weight_box[59]) );
  MUX21X1_HVT U486 ( .A1(conv2_sram_rdata_weight[87]), .A2(
        conv1_sram_rdata_weight[87]), .S0(n335), .Y(conv_weight_box[83]) );
  MUX21X1_HVT U487 ( .A1(conv2_sram_rdata_weight[26]), .A2(
        conv1_sram_rdata_weight[26]), .S0(n336), .Y(conv_weight_box[24]) );
  MUX21X1_HVT U488 ( .A1(conv2_sram_rdata_weight[51]), .A2(
        conv1_sram_rdata_weight[51]), .S0(n336), .Y(conv_weight_box[47]) );
  INVX1_HVT U489 ( .A(n438), .Y(n334) );
  MUX21X1_HVT U490 ( .A1(conv2_sram_rdata_weight[95]), .A2(
        conv1_sram_rdata_weight[95]), .S0(n336), .Y(conv_weight_box[90]) );
  MUX21X1_HVT U491 ( .A1(conv2_sram_rdata_weight[99]), .A2(
        conv1_sram_rdata_weight[99]), .S0(n336), .Y(conv_weight_box[93]) );
  INVX1_HVT U492 ( .A(n450), .Y(conv_weight_box[75]) );
  MUX21X1_HVT U493 ( .A1(conv2_sram_rdata_weight[49]), .A2(
        conv1_sram_rdata_weight[49]), .S0(n333), .Y(conv_weight_box[45]) );
  MUX21X1_HVT U494 ( .A1(conv2_sram_rdata_weight[45]), .A2(
        conv1_sram_rdata_weight[45]), .S0(n353), .Y(conv_weight_box[41]) );
  INVX1_HVT U495 ( .A(n440), .Y(conv_weight_box[49]) );
  MUX21X1_HVT U496 ( .A1(conv2_sram_rdata_weight[57]), .A2(
        conv1_sram_rdata_weight[57]), .S0(n353), .Y(conv_weight_box[53]) );
  MUX21X1_HVT U497 ( .A1(conv2_sram_rdata_weight[5]), .A2(
        conv1_sram_rdata_weight[5]), .S0(n335), .Y(conv_weight_box[4]) );
  MUX21X1_HVT U498 ( .A1(conv2_sram_rdata_weight[9]), .A2(
        conv1_sram_rdata_weight[9]), .S0(n352), .Y(conv_weight_box[8]) );
  INVX1_HVT U499 ( .A(n449), .Y(conv_weight_box[12]) );
  MUX21X1_HVT U500 ( .A1(conv2_sram_rdata_weight[73]), .A2(
        conv1_sram_rdata_weight[73]), .S0(n352), .Y(conv_weight_box[69]) );
  MUX21X1_HVT U501 ( .A1(conv2_sram_rdata_weight[93]), .A2(
        conv1_sram_rdata_weight[93]), .S0(n332), .Y(conv_weight_box[88]) );
  INVX1_HVT U502 ( .A(n453), .Y(n336) );
  INVX1_HVT U503 ( .A(n453), .Y(n335) );
  INVX1_HVT U504 ( .A(n453), .Y(n353) );
  INVX1_HVT U505 ( .A(n439), .Y(n349) );
  INVX1_HVT U506 ( .A(n453), .Y(n351) );
  INVX1_HVT U507 ( .A(n439), .Y(n350) );
  INVX1_HVT U508 ( .A(n439), .Y(n348) );
  INVX0_HVT U509 ( .A(n432), .Y(n438) );
  INVX1_HVT U510 ( .A(n453), .Y(n352) );
  NOR2X1_HVT U511 ( .A1(n539), .A2(n538), .Y(n590) );
  NOR2X1_HVT U512 ( .A1(n465), .A2(n464), .Y(n523) );
  INVX1_HVT U513 ( .A(srstn), .Y(n331) );
  NAND2X0_HVT U514 ( .A1(mode[1]), .A2(n687), .Y(n432) );
  AND2X1_HVT U515 ( .A1(n687), .A2(mode[1]), .Y(n439) );
  INVX1_HVT U516 ( .A(mode[0]), .Y(n687) );
  INVX2_HVT U517 ( .A(srstn), .Y(n346) );
  INVX1_HVT U518 ( .A(srstn), .Y(n347) );
  INVX2_HVT U519 ( .A(srstn), .Y(n345) );
  INVX2_HVT U520 ( .A(srstn), .Y(n344) );
  INVX1_HVT U521 ( .A(n437), .Y(n337) );
  INVX1_HVT U522 ( .A(n437), .Y(n338) );
  INVX1_HVT U523 ( .A(n437), .Y(DP_OP_422J2_124_3477_n2) );
  MUX21X1_HVT U524 ( .A1(conv2_sram_rdata_weight[48]), .A2(
        conv1_sram_rdata_weight[48]), .S0(n349), .Y(conv_weight_box[44]) );
  MUX21X1_HVT U525 ( .A1(conv2_sram_rdata_weight[35]), .A2(
        conv1_sram_rdata_weight[35]), .S0(n349), .Y(conv_weight_box[32]) );
  MUX21X1_HVT U526 ( .A1(conv2_sram_rdata_weight[2]), .A2(
        conv1_sram_rdata_weight[2]), .S0(n348), .Y(conv_weight_box[1]) );
  MUX21X1_HVT U527 ( .A1(conv2_sram_rdata_weight[64]), .A2(
        conv1_sram_rdata_weight[64]), .S0(n349), .Y(conv_weight_box[60]) );
  MUX21X1_HVT U528 ( .A1(conv2_sram_rdata_weight[10]), .A2(
        conv1_sram_rdata_weight[10]), .S0(n349), .Y(conv_weight_box[9]) );
  MUX21X1_HVT U529 ( .A1(conv2_sram_rdata_weight[4]), .A2(
        conv1_sram_rdata_weight[4]), .S0(n348), .Y(conv_weight_box[3]) );
  MUX21X1_HVT U530 ( .A1(conv2_sram_rdata_weight[68]), .A2(
        conv1_sram_rdata_weight[68]), .S0(n350), .Y(conv_weight_box[64]) );
  MUX21X1_HVT U531 ( .A1(conv2_sram_rdata_weight[52]), .A2(
        conv1_sram_rdata_weight[52]), .S0(n348), .Y(conv_weight_box[48]) );
  MUX21X1_HVT U532 ( .A1(conv2_sram_rdata_weight[92]), .A2(
        conv1_sram_rdata_weight[92]), .S0(n349), .Y(conv_weight_box[87]) );
  MUX21X1_HVT U533 ( .A1(conv2_sram_rdata_weight[88]), .A2(
        conv1_sram_rdata_weight[88]), .S0(n348), .Y(conv_weight_box[84]) );
  MUX21X1_HVT U534 ( .A1(conv2_sram_rdata_weight[39]), .A2(
        conv1_sram_rdata_weight[39]), .S0(n349), .Y(conv_weight_box[36]) );
  MUX21X1_HVT U535 ( .A1(conv2_sram_rdata_weight[20]), .A2(
        conv1_sram_rdata_weight[20]), .S0(n350), .Y(conv_weight_box[18]) );
  MUX21X1_HVT U536 ( .A1(conv2_sram_rdata_weight[56]), .A2(
        conv1_sram_rdata_weight[56]), .S0(n349), .Y(conv_weight_box[52]) );
  MUX21X1_HVT U537 ( .A1(conv2_sram_rdata_weight[80]), .A2(
        conv1_sram_rdata_weight[80]), .S0(n348), .Y(conv_weight_box[76]) );
  MUX21X1_HVT U538 ( .A1(conv2_sram_rdata_weight[47]), .A2(
        conv1_sram_rdata_weight[47]), .S0(n353), .Y(conv_weight_box[43]) );
  MUX21X1_HVT U539 ( .A1(conv2_sram_rdata_weight[23]), .A2(
        conv1_sram_rdata_weight[23]), .S0(n351), .Y(conv_weight_box[21]) );
  MUX21X1_HVT U540 ( .A1(conv2_sram_rdata_weight[59]), .A2(
        conv1_sram_rdata_weight[59]), .S0(n352), .Y(conv_weight_box[55]) );
  MUX21X1_HVT U541 ( .A1(conv2_sram_rdata_weight[75]), .A2(
        conv1_sram_rdata_weight[75]), .S0(n351), .Y(conv_weight_box[71]) );
  MUX21X1_HVT U542 ( .A1(conv2_sram_rdata_weight[67]), .A2(
        conv1_sram_rdata_weight[67]), .S0(n351), .Y(conv_weight_box[63]) );
  MUX21X1_HVT U543 ( .A1(conv2_sram_rdata_weight[3]), .A2(
        conv1_sram_rdata_weight[3]), .S0(n353), .Y(conv_weight_box[2]) );
  MUX21X1_HVT U544 ( .A1(conv2_sram_rdata_weight[66]), .A2(
        conv1_sram_rdata_weight[66]), .S0(n352), .Y(conv_weight_box[62]) );
  MUX21X1_HVT U545 ( .A1(conv2_sram_rdata_weight[71]), .A2(
        conv1_sram_rdata_weight[71]), .S0(n432), .Y(conv_weight_box[67]) );
  MUX21X1_HVT U546 ( .A1(conv2_sram_rdata_weight[83]), .A2(
        conv1_sram_rdata_weight[83]), .S0(n332), .Y(conv_weight_box[79]) );
  MUX21X1_HVT U547 ( .A1(conv2_sram_rdata_weight[30]), .A2(
        conv1_sram_rdata_weight[30]), .S0(n351), .Y(conv_weight_box[28]) );
  MUX21X1_HVT U548 ( .A1(conv2_sram_rdata_weight[89]), .A2(
        conv1_sram_rdata_weight[89]), .S0(n351), .Y(conv_weight_box[85]) );
  MUX21X1_HVT U549 ( .A1(conv2_sram_rdata_weight[32]), .A2(
        conv1_sram_rdata_weight[32]), .S0(n352), .Y(conv_weight_box[30]) );
  MUX21X1_HVT U550 ( .A1(conv2_sram_rdata_weight[61]), .A2(
        conv1_sram_rdata_weight[61]), .S0(n351), .Y(conv_weight_box[57]) );
  MUX21X1_HVT U551 ( .A1(conv2_sram_rdata_weight[1]), .A2(
        conv1_sram_rdata_weight[1]), .S0(n352), .Y(conv_weight_box[0]) );
  AND2X1_HVT U552 ( .A1(n659), .A2(n658), .Y(N9) );
  AND2X1_HVT U553 ( .A1(n594), .A2(n593), .Y(N7) );
  INVX1_HVT U554 ( .A(DP_OP_423J2_125_3477_n65), .Y(DP_OP_423J2_125_3477_n67)
         );
  INVX1_HVT U555 ( .A(DP_OP_423J2_125_3477_n148), .Y(DP_OP_423J2_125_3477_n149) );
  INVX1_HVT U556 ( .A(DP_OP_423J2_125_3477_n150), .Y(DP_OP_423J2_125_3477_n151) );
  INVX1_HVT U557 ( .A(DP_OP_423J2_125_3477_n152), .Y(DP_OP_423J2_125_3477_n153) );
  INVX1_HVT U558 ( .A(DP_OP_423J2_125_3477_n154), .Y(DP_OP_423J2_125_3477_n155) );
  INVX1_HVT U559 ( .A(DP_OP_423J2_125_3477_n156), .Y(DP_OP_423J2_125_3477_n157) );
  INVX1_HVT U560 ( .A(DP_OP_423J2_125_3477_n1574), .Y(
        DP_OP_423J2_125_3477_n1575) );
  INVX1_HVT U561 ( .A(DP_OP_423J2_125_3477_n158), .Y(DP_OP_423J2_125_3477_n159) );
  INVX1_HVT U562 ( .A(DP_OP_423J2_125_3477_n160), .Y(DP_OP_423J2_125_3477_n161) );
  INVX1_HVT U563 ( .A(DP_OP_423J2_125_3477_n162), .Y(DP_OP_423J2_125_3477_n163) );
  INVX1_HVT U564 ( .A(DP_OP_423J2_125_3477_n164), .Y(DP_OP_423J2_125_3477_n165) );
  INVX1_HVT U565 ( .A(DP_OP_423J2_125_3477_n166), .Y(DP_OP_423J2_125_3477_n167) );
  INVX1_HVT U566 ( .A(DP_OP_423J2_125_3477_n168), .Y(DP_OP_423J2_125_3477_n169) );
  INVX1_HVT U567 ( .A(DP_OP_423J2_125_3477_n170), .Y(DP_OP_423J2_125_3477_n171) );
  INVX1_HVT U568 ( .A(DP_OP_423J2_125_3477_n172), .Y(DP_OP_423J2_125_3477_n173) );
  INVX1_HVT U569 ( .A(DP_OP_423J2_125_3477_n174), .Y(DP_OP_423J2_125_3477_n175) );
  INVX1_HVT U570 ( .A(DP_OP_423J2_125_3477_n176), .Y(DP_OP_423J2_125_3477_n177) );
  INVX1_HVT U571 ( .A(src_window[63]), .Y(DP_OP_423J2_125_3477_n1849) );
  INVX1_HVT U572 ( .A(DP_OP_423J2_125_3477_n184), .Y(DP_OP_423J2_125_3477_n185) );
  INVX1_HVT U573 ( .A(src_window[62]), .Y(DP_OP_423J2_125_3477_n1850) );
  INVX1_HVT U574 ( .A(src_window[60]), .Y(DP_OP_423J2_125_3477_n1852) );
  INVX1_HVT U575 ( .A(src_window[59]), .Y(DP_OP_423J2_125_3477_n1853) );
  INVX1_HVT U576 ( .A(src_window[56]), .Y(DP_OP_423J2_125_3477_n1856) );
  INVX1_HVT U577 ( .A(conv_weight_box[5]), .Y(DP_OP_423J2_125_3477_n1858) );
  INVX1_HVT U578 ( .A(conv_weight_box[4]), .Y(DP_OP_423J2_125_3477_n1859) );
  INVX1_HVT U579 ( .A(conv_weight_box[3]), .Y(DP_OP_423J2_125_3477_n1860) );
  INVX1_HVT U580 ( .A(src_window[79]), .Y(DP_OP_423J2_125_3477_n1893) );
  INVX1_HVT U581 ( .A(src_window[76]), .Y(DP_OP_423J2_125_3477_n1896) );
  INVX1_HVT U582 ( .A(src_window[75]), .Y(DP_OP_423J2_125_3477_n1897) );
  INVX1_HVT U583 ( .A(src_window[74]), .Y(DP_OP_423J2_125_3477_n1898) );
  INVX1_HVT U584 ( .A(src_window[73]), .Y(DP_OP_423J2_125_3477_n1899) );
  INVX1_HVT U585 ( .A(conv_weight_box[13]), .Y(DP_OP_423J2_125_3477_n1901) );
  INVX1_HVT U586 ( .A(conv_weight_box[11]), .Y(DP_OP_423J2_125_3477_n1904) );
  INVX1_HVT U587 ( .A(src_window[103]), .Y(DP_OP_423J2_125_3477_n1937) );
  INVX1_HVT U588 ( .A(src_window[101]), .Y(DP_OP_423J2_125_3477_n1939) );
  INVX1_HVT U589 ( .A(src_window[97]), .Y(DP_OP_423J2_125_3477_n1943) );
  INVX1_HVT U590 ( .A(conv_weight_box[19]), .Y(DP_OP_423J2_125_3477_n1947) );
  INVX1_HVT U591 ( .A(conv_weight_box[18]), .Y(DP_OP_423J2_125_3477_n1948) );
  INVX1_HVT U592 ( .A(src_window[117]), .Y(DP_OP_423J2_125_3477_n1983) );
  INVX1_HVT U593 ( .A(src_window[115]), .Y(DP_OP_423J2_125_3477_n1985) );
  INVX1_HVT U594 ( .A(src_window[114]), .Y(DP_OP_423J2_125_3477_n1986) );
  INVX1_HVT U595 ( .A(conv_weight_box[29]), .Y(DP_OP_423J2_125_3477_n1989) );
  INVX1_HVT U596 ( .A(conv_weight_box[27]), .Y(DP_OP_423J2_125_3477_n1991) );
  INVX1_HVT U597 ( .A(conv_weight_box[26]), .Y(DP_OP_423J2_125_3477_n1992) );
  INVX1_HVT U598 ( .A(src_window[132]), .Y(DP_OP_423J2_125_3477_n2028) );
  INVX1_HVT U599 ( .A(src_window[131]), .Y(DP_OP_423J2_125_3477_n2029) );
  INVX1_HVT U600 ( .A(src_window[130]), .Y(DP_OP_423J2_125_3477_n2030) );
  INVX1_HVT U601 ( .A(src_window[129]), .Y(DP_OP_423J2_125_3477_n2031) );
  INVX1_HVT U602 ( .A(src_window[128]), .Y(DP_OP_423J2_125_3477_n2032) );
  INVX1_HVT U603 ( .A(conv_weight_box[36]), .Y(DP_OP_423J2_125_3477_n2033) );
  INVX1_HVT U604 ( .A(conv_weight_box[35]), .Y(DP_OP_423J2_125_3477_n2034) );
  INVX1_HVT U605 ( .A(src_window[155]), .Y(DP_OP_423J2_125_3477_n2073) );
  INVX1_HVT U606 ( .A(src_window[154]), .Y(DP_OP_423J2_125_3477_n2074) );
  INVX1_HVT U607 ( .A(src_window[152]), .Y(DP_OP_423J2_125_3477_n2076) );
  INVX1_HVT U608 ( .A(conv_weight_box[43]), .Y(DP_OP_423J2_125_3477_n2077) );
  INVX1_HVT U609 ( .A(conv_weight_box[40]), .Y(DP_OP_423J2_125_3477_n2080) );
  INVX1_HVT U610 ( .A(src_window[174]), .Y(DP_OP_423J2_125_3477_n2114) );
  INVX1_HVT U611 ( .A(src_window[173]), .Y(DP_OP_423J2_125_3477_n2115) );
  INVX1_HVT U612 ( .A(src_window[172]), .Y(DP_OP_423J2_125_3477_n2116) );
  INVX1_HVT U613 ( .A(src_window[171]), .Y(DP_OP_423J2_125_3477_n2117) );
  INVX1_HVT U614 ( .A(conv_weight_box[50]), .Y(DP_OP_423J2_125_3477_n2122) );
  INVX1_HVT U615 ( .A(src_window[199]), .Y(DP_OP_423J2_125_3477_n2157) );
  INVX1_HVT U616 ( .A(src_window[198]), .Y(DP_OP_423J2_125_3477_n2158) );
  INVX1_HVT U617 ( .A(src_window[196]), .Y(DP_OP_423J2_125_3477_n2160) );
  INVX1_HVT U618 ( .A(src_window[195]), .Y(DP_OP_423J2_125_3477_n2161) );
  INVX1_HVT U619 ( .A(src_window[193]), .Y(DP_OP_423J2_125_3477_n2163) );
  INVX1_HVT U620 ( .A(src_window[192]), .Y(DP_OP_423J2_125_3477_n2164) );
  INVX1_HVT U621 ( .A(conv_weight_box[59]), .Y(DP_OP_423J2_125_3477_n2165) );
  INVX1_HVT U622 ( .A(conv_weight_box[57]), .Y(DP_OP_423J2_125_3477_n2167) );
  INVX1_HVT U623 ( .A(conv_weight_box[56]), .Y(DP_OP_423J2_125_3477_n2168) );
  INVX1_HVT U624 ( .A(src_window[212]), .Y(DP_OP_423J2_125_3477_n2204) );
  INVX1_HVT U625 ( .A(src_window[211]), .Y(DP_OP_423J2_125_3477_n2205) );
  INVX1_HVT U626 ( .A(conv_weight_box[67]), .Y(DP_OP_423J2_125_3477_n2209) );
  INVX1_HVT U627 ( .A(conv_weight_box[65]), .Y(DP_OP_423J2_125_3477_n2211) );
  INVX1_HVT U628 ( .A(conv_weight_box[64]), .Y(DP_OP_423J2_125_3477_n2212) );
  INVX1_HVT U629 ( .A(src_window[229]), .Y(DP_OP_423J2_125_3477_n2247) );
  INVX1_HVT U630 ( .A(src_window[225]), .Y(DP_OP_423J2_125_3477_n2251) );
  INVX1_HVT U631 ( .A(conv_weight_box[74]), .Y(DP_OP_423J2_125_3477_n2254) );
  INVX1_HVT U632 ( .A(conv_weight_box[72]), .Y(DP_OP_423J2_125_3477_n2256) );
  INVX1_HVT U633 ( .A(src_window[253]), .Y(DP_OP_423J2_125_3477_n2291) );
  INVX1_HVT U634 ( .A(src_window[250]), .Y(DP_OP_423J2_125_3477_n2294) );
  INVX1_HVT U635 ( .A(src_window[249]), .Y(DP_OP_423J2_125_3477_n2295) );
  INVX1_HVT U636 ( .A(conv_weight_box[82]), .Y(DP_OP_423J2_125_3477_n2298) );
  INVX1_HVT U637 ( .A(conv_weight_box[81]), .Y(DP_OP_423J2_125_3477_n2299) );
  INVX1_HVT U638 ( .A(src_window[271]), .Y(DP_OP_423J2_125_3477_n2333) );
  INVX1_HVT U639 ( .A(src_window[270]), .Y(DP_OP_423J2_125_3477_n2334) );
  INVX1_HVT U640 ( .A(src_window[265]), .Y(DP_OP_423J2_125_3477_n2339) );
  INVX1_HVT U641 ( .A(conv_weight_box[90]), .Y(DP_OP_423J2_125_3477_n2341) );
  INVX1_HVT U642 ( .A(conv_weight_box[88]), .Y(DP_OP_423J2_125_3477_n2343) );
  INVX1_HVT U643 ( .A(conv_weight_box[87]), .Y(DP_OP_423J2_125_3477_n2344) );
  INVX1_HVT U644 ( .A(src_window[279]), .Y(DP_OP_423J2_125_3477_n2377) );
  INVX1_HVT U645 ( .A(conv_weight_box[92]), .Y(DP_OP_423J2_125_3477_n2386) );
  INVX1_HVT U646 ( .A(conv_weight_box[91]), .Y(DP_OP_423J2_125_3477_n2387) );
  INVX1_HVT U647 ( .A(n430), .Y(DP_OP_423J2_125_3477_n2388) );
  INVX1_HVT U648 ( .A(src_window[263]), .Y(DP_OP_423J2_125_3477_n2421) );
  INVX1_HVT U649 ( .A(src_window[260]), .Y(DP_OP_423J2_125_3477_n2424) );
  INVX1_HVT U650 ( .A(src_window[259]), .Y(DP_OP_423J2_125_3477_n2425) );
  INVX1_HVT U651 ( .A(src_window[256]), .Y(DP_OP_423J2_125_3477_n2428) );
  INVX1_HVT U652 ( .A(DP_OP_425J2_127_3477_n3255), .Y(
        DP_OP_423J2_125_3477_n2429) );
  INVX1_HVT U653 ( .A(conv_weight_box[86]), .Y(DP_OP_423J2_125_3477_n2430) );
  INVX1_HVT U654 ( .A(conv_weight_box[85]), .Y(DP_OP_423J2_125_3477_n2431) );
  INVX1_HVT U655 ( .A(conv_weight_box[84]), .Y(DP_OP_423J2_125_3477_n2432) );
  INVX1_HVT U656 ( .A(src_window[247]), .Y(DP_OP_423J2_125_3477_n2465) );
  INVX1_HVT U657 ( .A(src_window[246]), .Y(DP_OP_423J2_125_3477_n2466) );
  INVX1_HVT U658 ( .A(src_window[245]), .Y(DP_OP_423J2_125_3477_n2467) );
  INVX1_HVT U659 ( .A(src_window[244]), .Y(DP_OP_423J2_125_3477_n2468) );
  INVX1_HVT U660 ( .A(src_window[243]), .Y(DP_OP_423J2_125_3477_n2469) );
  INVX1_HVT U661 ( .A(src_window[242]), .Y(DP_OP_423J2_125_3477_n2470) );
  INVX1_HVT U662 ( .A(src_window[241]), .Y(DP_OP_423J2_125_3477_n2471) );
  INVX1_HVT U663 ( .A(src_window[240]), .Y(DP_OP_423J2_125_3477_n2472) );
  INVX1_HVT U664 ( .A(conv_weight_box[78]), .Y(DP_OP_423J2_125_3477_n2474) );
  INVX1_HVT U665 ( .A(conv_weight_box[77]), .Y(DP_OP_423J2_125_3477_n2475) );
  INVX1_HVT U666 ( .A(conv_weight_box[76]), .Y(DP_OP_423J2_125_3477_n2476) );
  INVX1_HVT U667 ( .A(src_window[223]), .Y(DP_OP_423J2_125_3477_n2509) );
  INVX1_HVT U668 ( .A(src_window[222]), .Y(DP_OP_423J2_125_3477_n2510) );
  INVX1_HVT U669 ( .A(src_window[217]), .Y(DP_OP_423J2_125_3477_n2515) );
  INVX1_HVT U670 ( .A(src_window[216]), .Y(DP_OP_423J2_125_3477_n2516) );
  INVX1_HVT U671 ( .A(conv_weight_box[71]), .Y(DP_OP_423J2_125_3477_n2517) );
  INVX1_HVT U672 ( .A(conv_weight_box[69]), .Y(DP_OP_423J2_125_3477_n2519) );
  INVX1_HVT U673 ( .A(conv_weight_box[68]), .Y(DP_OP_423J2_125_3477_n2520) );
  INVX1_HVT U674 ( .A(src_window[207]), .Y(DP_OP_423J2_125_3477_n2553) );
  INVX1_HVT U675 ( .A(src_window[206]), .Y(DP_OP_423J2_125_3477_n2554) );
  INVX1_HVT U676 ( .A(src_window[202]), .Y(DP_OP_423J2_125_3477_n2558) );
  INVX1_HVT U677 ( .A(src_window[201]), .Y(DP_OP_423J2_125_3477_n2559) );
  INVX1_HVT U678 ( .A(conv_weight_box[63]), .Y(DP_OP_423J2_125_3477_n2561) );
  INVX1_HVT U679 ( .A(conv_weight_box[62]), .Y(DP_OP_423J2_125_3477_n2562) );
  INVX1_HVT U680 ( .A(src_window[181]), .Y(DP_OP_423J2_125_3477_n2599) );
  INVX1_HVT U681 ( .A(src_window[180]), .Y(DP_OP_423J2_125_3477_n2600) );
  INVX1_HVT U682 ( .A(src_window[179]), .Y(DP_OP_423J2_125_3477_n2601) );
  INVX1_HVT U683 ( .A(src_window[178]), .Y(DP_OP_423J2_125_3477_n2602) );
  INVX1_HVT U684 ( .A(src_window[177]), .Y(DP_OP_423J2_125_3477_n2603) );
  INVX1_HVT U685 ( .A(src_window[176]), .Y(DP_OP_423J2_125_3477_n2604) );
  INVX1_HVT U686 ( .A(conv_weight_box[55]), .Y(DP_OP_423J2_125_3477_n2605) );
  INVX1_HVT U687 ( .A(conv_weight_box[53]), .Y(DP_OP_423J2_125_3477_n2607) );
  INVX1_HVT U688 ( .A(src_window[166]), .Y(DP_OP_423J2_125_3477_n2642) );
  INVX1_HVT U689 ( .A(src_window[165]), .Y(DP_OP_423J2_125_3477_n2643) );
  INVX1_HVT U690 ( .A(src_window[163]), .Y(DP_OP_423J2_125_3477_n2645) );
  INVX1_HVT U691 ( .A(src_window[162]), .Y(DP_OP_423J2_125_3477_n2646) );
  INVX1_HVT U692 ( .A(src_window[161]), .Y(DP_OP_423J2_125_3477_n2647) );
  INVX1_HVT U693 ( .A(src_window[160]), .Y(DP_OP_423J2_125_3477_n2648) );
  INVX1_HVT U694 ( .A(conv_weight_box[47]), .Y(DP_OP_423J2_125_3477_n2649) );
  INVX1_HVT U695 ( .A(conv_weight_box[45]), .Y(DP_OP_423J2_125_3477_n2651) );
  INVX1_HVT U696 ( .A(src_window[148]), .Y(DP_OP_423J2_125_3477_n2688) );
  INVX1_HVT U697 ( .A(src_window[146]), .Y(DP_OP_423J2_125_3477_n2690) );
  INVX1_HVT U698 ( .A(conv_weight_box[39]), .Y(DP_OP_423J2_125_3477_n2693) );
  INVX1_HVT U699 ( .A(conv_weight_box[38]), .Y(DP_OP_423J2_125_3477_n2695) );
  INVX1_HVT U700 ( .A(conv_weight_box[37]), .Y(DP_OP_423J2_125_3477_n2696) );
  INVX1_HVT U701 ( .A(src_window[127]), .Y(DP_OP_423J2_125_3477_n2726) );
  INVX1_HVT U702 ( .A(src_window[124]), .Y(DP_OP_423J2_125_3477_n2729) );
  INVX1_HVT U703 ( .A(src_window[123]), .Y(DP_OP_423J2_125_3477_n2730) );
  INVX1_HVT U704 ( .A(src_window[122]), .Y(DP_OP_423J2_125_3477_n2731) );
  INVX1_HVT U705 ( .A(src_window[121]), .Y(DP_OP_423J2_125_3477_n2732) );
  INVX1_HVT U706 ( .A(src_window[120]), .Y(DP_OP_423J2_125_3477_n2733) );
  INVX1_HVT U707 ( .A(conv_weight_box[32]), .Y(DP_OP_423J2_125_3477_n2734) );
  INVX1_HVT U708 ( .A(conv_weight_box[30]), .Y(DP_OP_423J2_125_3477_n2737) );
  INVX1_HVT U709 ( .A(src_window[111]), .Y(DP_OP_423J2_125_3477_n2770) );
  INVX1_HVT U710 ( .A(src_window[109]), .Y(DP_OP_423J2_125_3477_n2772) );
  INVX1_HVT U711 ( .A(src_window[106]), .Y(DP_OP_423J2_125_3477_n2775) );
  INVX1_HVT U712 ( .A(src_window[105]), .Y(DP_OP_423J2_125_3477_n2776) );
  INVX1_HVT U713 ( .A(src_window[104]), .Y(DP_OP_423J2_125_3477_n2777) );
  INVX1_HVT U714 ( .A(conv_weight_box[25]), .Y(DP_OP_423J2_125_3477_n2778) );
  INVX1_HVT U715 ( .A(conv_weight_box[24]), .Y(DP_OP_423J2_125_3477_n2779) );
  INVX1_HVT U716 ( .A(conv_weight_box[22]), .Y(DP_OP_423J2_125_3477_n2781) );
  INVX1_HVT U717 ( .A(conv_weight_box[16]), .Y(DP_OP_423J2_125_3477_n2823) );
  INVX1_HVT U718 ( .A(conv_weight_box[15]), .Y(DP_OP_423J2_125_3477_n2824) );
  INVX1_HVT U719 ( .A(src_window[70]), .Y(DP_OP_423J2_125_3477_n2859) );
  INVX1_HVT U720 ( .A(src_window[69]), .Y(DP_OP_423J2_125_3477_n2860) );
  INVX1_HVT U721 ( .A(src_window[68]), .Y(DP_OP_423J2_125_3477_n2861) );
  INVX1_HVT U722 ( .A(src_window[65]), .Y(DP_OP_423J2_125_3477_n2864) );
  INVX1_HVT U723 ( .A(src_window[64]), .Y(DP_OP_423J2_125_3477_n2865) );
  INVX1_HVT U724 ( .A(conv_weight_box[10]), .Y(DP_OP_423J2_125_3477_n2866) );
  INVX1_HVT U725 ( .A(conv_weight_box[9]), .Y(DP_OP_423J2_125_3477_n2867) );
  INVX1_HVT U726 ( .A(conv_weight_box[8]), .Y(DP_OP_423J2_125_3477_n2868) );
  INVX1_HVT U727 ( .A(conv_weight_box[7]), .Y(DP_OP_423J2_125_3477_n2869) );
  INVX1_HVT U728 ( .A(src_window[55]), .Y(DP_OP_423J2_125_3477_n2902) );
  INVX1_HVT U729 ( .A(src_window[54]), .Y(DP_OP_423J2_125_3477_n2903) );
  INVX1_HVT U730 ( .A(src_window[53]), .Y(DP_OP_423J2_125_3477_n2904) );
  INVX1_HVT U731 ( .A(src_window[51]), .Y(DP_OP_423J2_125_3477_n2906) );
  INVX1_HVT U732 ( .A(src_window[50]), .Y(DP_OP_423J2_125_3477_n2907) );
  INVX1_HVT U733 ( .A(src_window[49]), .Y(DP_OP_423J2_125_3477_n2908) );
  INVX1_HVT U734 ( .A(src_window[48]), .Y(DP_OP_423J2_125_3477_n2909) );
  INVX1_HVT U735 ( .A(conv_weight_box[2]), .Y(DP_OP_423J2_125_3477_n2910) );
  INVX1_HVT U736 ( .A(conv_weight_box[1]), .Y(DP_OP_423J2_125_3477_n2911) );
  INVX1_HVT U737 ( .A(n429), .Y(DP_OP_423J2_125_3477_n2913) );
  INVX1_HVT U738 ( .A(DP_OP_423J2_125_3477_n356), .Y(DP_OP_423J2_125_3477_n357) );
  INVX1_HVT U739 ( .A(DP_OP_423J2_125_3477_n666), .Y(DP_OP_423J2_125_3477_n667) );
  INVX1_HVT U740 ( .A(DP_OP_423J2_125_3477_n72), .Y(DP_OP_423J2_125_3477_n71)
         );
  INVX1_HVT U741 ( .A(DP_OP_422J2_124_3477_n67), .Y(DP_OP_422J2_124_3477_n69)
         );
  INVX1_HVT U742 ( .A(DP_OP_422J2_124_3477_n153), .Y(DP_OP_422J2_124_3477_n154) );
  INVX1_HVT U743 ( .A(DP_OP_422J2_124_3477_n155), .Y(DP_OP_422J2_124_3477_n156) );
  INVX1_HVT U744 ( .A(DP_OP_422J2_124_3477_n157), .Y(DP_OP_422J2_124_3477_n158) );
  INVX1_HVT U745 ( .A(DP_OP_422J2_124_3477_n1579), .Y(
        DP_OP_422J2_124_3477_n1580) );
  INVX1_HVT U746 ( .A(DP_OP_422J2_124_3477_n159), .Y(DP_OP_422J2_124_3477_n160) );
  INVX1_HVT U747 ( .A(DP_OP_422J2_124_3477_n161), .Y(DP_OP_422J2_124_3477_n162) );
  INVX1_HVT U748 ( .A(DP_OP_422J2_124_3477_n163), .Y(DP_OP_422J2_124_3477_n164) );
  INVX1_HVT U749 ( .A(DP_OP_422J2_124_3477_n165), .Y(DP_OP_422J2_124_3477_n166) );
  INVX1_HVT U750 ( .A(DP_OP_422J2_124_3477_n167), .Y(DP_OP_422J2_124_3477_n168) );
  INVX1_HVT U751 ( .A(DP_OP_422J2_124_3477_n169), .Y(DP_OP_422J2_124_3477_n170) );
  INVX1_HVT U752 ( .A(DP_OP_422J2_124_3477_n171), .Y(DP_OP_422J2_124_3477_n172) );
  INVX1_HVT U753 ( .A(DP_OP_422J2_124_3477_n173), .Y(DP_OP_422J2_124_3477_n174) );
  INVX1_HVT U754 ( .A(DP_OP_422J2_124_3477_n175), .Y(DP_OP_422J2_124_3477_n176) );
  INVX1_HVT U755 ( .A(DP_OP_422J2_124_3477_n177), .Y(DP_OP_422J2_124_3477_n178) );
  INVX1_HVT U756 ( .A(DP_OP_422J2_124_3477_n179), .Y(DP_OP_422J2_124_3477_n180) );
  INVX1_HVT U757 ( .A(DP_OP_422J2_124_3477_n181), .Y(DP_OP_422J2_124_3477_n182) );
  INVX1_HVT U758 ( .A(src_window[71]), .Y(DP_OP_422J2_124_3477_n1854) );
  INVX1_HVT U759 ( .A(src_window[70]), .Y(DP_OP_422J2_124_3477_n1855) );
  INVX1_HVT U760 ( .A(src_window[67]), .Y(DP_OP_422J2_124_3477_n1858) );
  INVX1_HVT U761 ( .A(src_window[66]), .Y(DP_OP_422J2_124_3477_n1859) );
  INVX1_HVT U762 ( .A(src_window[64]), .Y(DP_OP_422J2_124_3477_n1861) );
  INVX1_HVT U763 ( .A(conv_weight_box[6]), .Y(DP_OP_422J2_124_3477_n1862) );
  INVX1_HVT U764 ( .A(conv_weight_box[5]), .Y(DP_OP_422J2_124_3477_n1863) );
  INVX1_HVT U765 ( .A(conv_weight_box[4]), .Y(DP_OP_422J2_124_3477_n1864) );
  INVX1_HVT U766 ( .A(conv_weight_box[3]), .Y(DP_OP_422J2_124_3477_n1865) );
  INVX1_HVT U767 ( .A(src_window[87]), .Y(DP_OP_422J2_124_3477_n1898) );
  INVX1_HVT U768 ( .A(src_window[86]), .Y(DP_OP_422J2_124_3477_n1899) );
  INVX1_HVT U769 ( .A(DP_OP_422J2_124_3477_n189), .Y(DP_OP_422J2_124_3477_n190) );
  INVX1_HVT U770 ( .A(src_window[85]), .Y(DP_OP_422J2_124_3477_n1900) );
  INVX1_HVT U771 ( .A(src_window[83]), .Y(DP_OP_422J2_124_3477_n1902) );
  INVX1_HVT U772 ( .A(src_window[82]), .Y(DP_OP_422J2_124_3477_n1903) );
  INVX1_HVT U773 ( .A(src_window[81]), .Y(DP_OP_422J2_124_3477_n1904) );
  INVX1_HVT U774 ( .A(src_window[80]), .Y(DP_OP_422J2_124_3477_n1905) );
  INVX1_HVT U775 ( .A(conv_weight_box[13]), .Y(DP_OP_422J2_124_3477_n1906) );
  INVX1_HVT U776 ( .A(n431), .Y(DP_OP_422J2_124_3477_n1907) );
  INVX1_HVT U777 ( .A(conv_weight_box[12]), .Y(DP_OP_422J2_124_3477_n1908) );
  INVX1_HVT U778 ( .A(conv_weight_box[11]), .Y(DP_OP_422J2_124_3477_n1909) );
  INVX1_HVT U779 ( .A(src_window[110]), .Y(DP_OP_422J2_124_3477_n1943) );
  INVX1_HVT U780 ( .A(src_window[108]), .Y(DP_OP_422J2_124_3477_n1945) );
  INVX1_HVT U781 ( .A(src_window[104]), .Y(DP_OP_422J2_124_3477_n1949) );
  INVX1_HVT U782 ( .A(conv_weight_box[21]), .Y(DP_OP_422J2_124_3477_n1950) );
  INVX1_HVT U783 ( .A(conv_weight_box[20]), .Y(DP_OP_422J2_124_3477_n1951) );
  INVX1_HVT U784 ( .A(conv_weight_box[19]), .Y(DP_OP_422J2_124_3477_n1952) );
  INVX1_HVT U785 ( .A(src_window[125]), .Y(DP_OP_422J2_124_3477_n1988) );
  INVX1_HVT U786 ( .A(src_window[124]), .Y(DP_OP_422J2_124_3477_n1989) );
  INVX1_HVT U787 ( .A(src_window[122]), .Y(DP_OP_422J2_124_3477_n1991) );
  INVX1_HVT U788 ( .A(conv_weight_box[29]), .Y(DP_OP_422J2_124_3477_n1994) );
  INVX1_HVT U789 ( .A(conv_weight_box[28]), .Y(DP_OP_422J2_124_3477_n1995) );
  INVX1_HVT U790 ( .A(conv_weight_box[27]), .Y(DP_OP_422J2_124_3477_n1996) );
  INVX1_HVT U791 ( .A(conv_weight_box[26]), .Y(DP_OP_422J2_124_3477_n1997) );
  INVX1_HVT U792 ( .A(src_window[143]), .Y(DP_OP_422J2_124_3477_n2029) );
  INVX1_HVT U793 ( .A(src_window[141]), .Y(DP_OP_422J2_124_3477_n2031) );
  INVX1_HVT U794 ( .A(src_window[140]), .Y(DP_OP_422J2_124_3477_n2032) );
  INVX1_HVT U795 ( .A(src_window[139]), .Y(DP_OP_422J2_124_3477_n2033) );
  INVX1_HVT U796 ( .A(src_window[137]), .Y(DP_OP_422J2_124_3477_n2035) );
  INVX1_HVT U797 ( .A(src_window[136]), .Y(DP_OP_422J2_124_3477_n2036) );
  INVX1_HVT U798 ( .A(conv_weight_box[36]), .Y(DP_OP_422J2_124_3477_n2037) );
  INVX1_HVT U799 ( .A(conv_weight_box[34]), .Y(DP_OP_422J2_124_3477_n2039) );
  INVX1_HVT U800 ( .A(conv_weight_box[33]), .Y(DP_OP_422J2_124_3477_n2040) );
  INVX1_HVT U801 ( .A(src_window[167]), .Y(DP_OP_422J2_124_3477_n2073) );
  INVX1_HVT U802 ( .A(src_window[166]), .Y(DP_OP_422J2_124_3477_n2074) );
  INVX1_HVT U803 ( .A(src_window[164]), .Y(DP_OP_422J2_124_3477_n2076) );
  INVX1_HVT U804 ( .A(src_window[162]), .Y(DP_OP_422J2_124_3477_n2078) );
  INVX1_HVT U805 ( .A(conv_weight_box[43]), .Y(DP_OP_422J2_124_3477_n2081) );
  INVX1_HVT U806 ( .A(conv_weight_box[42]), .Y(DP_OP_422J2_124_3477_n2082) );
  INVX1_HVT U807 ( .A(conv_weight_box[41]), .Y(DP_OP_422J2_124_3477_n2083) );
  INVX1_HVT U808 ( .A(src_window[183]), .Y(DP_OP_422J2_124_3477_n2117) );
  INVX1_HVT U809 ( .A(src_window[182]), .Y(DP_OP_422J2_124_3477_n2118) );
  INVX1_HVT U810 ( .A(src_window[180]), .Y(DP_OP_422J2_124_3477_n2120) );
  INVX1_HVT U811 ( .A(src_window[179]), .Y(DP_OP_422J2_124_3477_n2121) );
  INVX1_HVT U812 ( .A(src_window[176]), .Y(DP_OP_422J2_124_3477_n2124) );
  INVX1_HVT U813 ( .A(conv_weight_box[51]), .Y(DP_OP_422J2_124_3477_n2125) );
  INVX1_HVT U814 ( .A(conv_weight_box[49]), .Y(DP_OP_422J2_124_3477_n2127) );
  INVX1_HVT U815 ( .A(conv_weight_box[48]), .Y(DP_OP_422J2_124_3477_n2128) );
  INVX1_HVT U816 ( .A(src_window[206]), .Y(DP_OP_422J2_124_3477_n2162) );
  INVX1_HVT U817 ( .A(src_window[205]), .Y(DP_OP_422J2_124_3477_n2163) );
  INVX1_HVT U818 ( .A(src_window[204]), .Y(DP_OP_422J2_124_3477_n2164) );
  INVX1_HVT U819 ( .A(src_window[203]), .Y(DP_OP_422J2_124_3477_n2165) );
  INVX1_HVT U820 ( .A(src_window[200]), .Y(DP_OP_422J2_124_3477_n2168) );
  INVX1_HVT U821 ( .A(conv_weight_box[59]), .Y(DP_OP_422J2_124_3477_n2169) );
  INVX1_HVT U822 ( .A(conv_weight_box[58]), .Y(DP_OP_422J2_124_3477_n2170) );
  INVX1_HVT U823 ( .A(conv_weight_box[57]), .Y(DP_OP_422J2_124_3477_n2171) );
  INVX1_HVT U824 ( .A(src_window[221]), .Y(DP_OP_422J2_124_3477_n2207) );
  INVX1_HVT U825 ( .A(src_window[220]), .Y(DP_OP_422J2_124_3477_n2208) );
  INVX1_HVT U826 ( .A(src_window[219]), .Y(DP_OP_422J2_124_3477_n2209) );
  INVX1_HVT U827 ( .A(src_window[218]), .Y(DP_OP_422J2_124_3477_n2210) );
  INVX1_HVT U828 ( .A(src_window[217]), .Y(DP_OP_422J2_124_3477_n2211) );
  INVX1_HVT U829 ( .A(conv_weight_box[67]), .Y(DP_OP_422J2_124_3477_n2213) );
  INVX1_HVT U830 ( .A(conv_weight_box[66]), .Y(DP_OP_422J2_124_3477_n2214) );
  INVX1_HVT U831 ( .A(conv_weight_box[65]), .Y(DP_OP_422J2_124_3477_n2215) );
  INVX1_HVT U832 ( .A(conv_weight_box[64]), .Y(DP_OP_422J2_124_3477_n2216) );
  INVX1_HVT U833 ( .A(src_window[239]), .Y(DP_OP_422J2_124_3477_n2249) );
  INVX1_HVT U834 ( .A(src_window[238]), .Y(DP_OP_422J2_124_3477_n2250) );
  INVX1_HVT U835 ( .A(conv_weight_box[75]), .Y(DP_OP_422J2_124_3477_n2257) );
  INVX1_HVT U836 ( .A(conv_weight_box[74]), .Y(DP_OP_422J2_124_3477_n2258) );
  INVX1_HVT U837 ( .A(conv_weight_box[73]), .Y(DP_OP_422J2_124_3477_n2259) );
  INVX1_HVT U838 ( .A(conv_weight_box[72]), .Y(DP_OP_422J2_124_3477_n2260) );
  INVX1_HVT U839 ( .A(src_window[262]), .Y(DP_OP_422J2_124_3477_n2294) );
  INVX1_HVT U840 ( .A(src_window[261]), .Y(DP_OP_422J2_124_3477_n2295) );
  INVX1_HVT U841 ( .A(src_window[258]), .Y(DP_OP_422J2_124_3477_n2298) );
  INVX1_HVT U842 ( .A(src_window[257]), .Y(DP_OP_422J2_124_3477_n2299) );
  INVX1_HVT U843 ( .A(conv_weight_box[83]), .Y(DP_OP_422J2_124_3477_n2301) );
  INVX1_HVT U844 ( .A(conv_weight_box[82]), .Y(DP_OP_422J2_124_3477_n2302) );
  INVX1_HVT U845 ( .A(conv_weight_box[80]), .Y(DP_OP_422J2_124_3477_n2304) );
  INVX1_HVT U846 ( .A(src_window[278]), .Y(DP_OP_422J2_124_3477_n2338) );
  INVX1_HVT U847 ( .A(src_window[277]), .Y(DP_OP_422J2_124_3477_n2339) );
  INVX1_HVT U848 ( .A(src_window[276]), .Y(DP_OP_422J2_124_3477_n2340) );
  INVX1_HVT U849 ( .A(src_window[275]), .Y(DP_OP_422J2_124_3477_n2341) );
  INVX1_HVT U850 ( .A(src_window[274]), .Y(DP_OP_422J2_124_3477_n2342) );
  INVX1_HVT U851 ( .A(src_window[273]), .Y(DP_OP_422J2_124_3477_n2343) );
  INVX1_HVT U852 ( .A(src_window[272]), .Y(DP_OP_422J2_124_3477_n2344) );
  INVX1_HVT U853 ( .A(conv_weight_box[90]), .Y(DP_OP_422J2_124_3477_n2345) );
  INVX1_HVT U854 ( .A(conv_weight_box[89]), .Y(DP_OP_422J2_124_3477_n2346) );
  INVX1_HVT U855 ( .A(conv_weight_box[88]), .Y(DP_OP_422J2_124_3477_n2347) );
  INVX1_HVT U856 ( .A(src_window[287]), .Y(DP_OP_422J2_124_3477_n2381) );
  INVX1_HVT U857 ( .A(src_window[286]), .Y(DP_OP_422J2_124_3477_n2382) );
  INVX1_HVT U858 ( .A(src_window[285]), .Y(DP_OP_422J2_124_3477_n2383) );
  INVX1_HVT U859 ( .A(src_window[284]), .Y(DP_OP_422J2_124_3477_n2384) );
  INVX1_HVT U860 ( .A(src_window[283]), .Y(DP_OP_422J2_124_3477_n2385) );
  INVX1_HVT U861 ( .A(src_window[282]), .Y(DP_OP_422J2_124_3477_n2386) );
  INVX1_HVT U862 ( .A(src_window[281]), .Y(DP_OP_422J2_124_3477_n2387) );
  INVX1_HVT U863 ( .A(src_window[280]), .Y(DP_OP_422J2_124_3477_n2388) );
  INVX1_HVT U864 ( .A(conv_weight_box[93]), .Y(DP_OP_422J2_124_3477_n2389) );
  INVX1_HVT U865 ( .A(conv_weight_box[92]), .Y(DP_OP_422J2_124_3477_n2390) );
  INVX1_HVT U866 ( .A(conv_weight_box[91]), .Y(DP_OP_422J2_124_3477_n2391) );
  INVX1_HVT U867 ( .A(n430), .Y(DP_OP_422J2_124_3477_n2392) );
  INVX1_HVT U868 ( .A(src_window[269]), .Y(DP_OP_422J2_124_3477_n2427) );
  INVX1_HVT U869 ( .A(src_window[268]), .Y(DP_OP_422J2_124_3477_n2428) );
  INVX1_HVT U870 ( .A(src_window[267]), .Y(DP_OP_422J2_124_3477_n2429) );
  INVX1_HVT U871 ( .A(src_window[266]), .Y(DP_OP_422J2_124_3477_n2430) );
  INVX1_HVT U872 ( .A(src_window[264]), .Y(DP_OP_422J2_124_3477_n2432) );
  INVX1_HVT U873 ( .A(DP_OP_425J2_127_3477_n3255), .Y(
        DP_OP_422J2_124_3477_n2433) );
  INVX1_HVT U874 ( .A(conv_weight_box[86]), .Y(DP_OP_422J2_124_3477_n2434) );
  INVX1_HVT U875 ( .A(conv_weight_box[85]), .Y(DP_OP_422J2_124_3477_n2435) );
  INVX1_HVT U876 ( .A(conv_weight_box[84]), .Y(DP_OP_422J2_124_3477_n2436) );
  INVX1_HVT U877 ( .A(src_window[255]), .Y(DP_OP_422J2_124_3477_n2469) );
  INVX1_HVT U878 ( .A(src_window[254]), .Y(DP_OP_422J2_124_3477_n2470) );
  INVX1_HVT U879 ( .A(src_window[252]), .Y(DP_OP_422J2_124_3477_n2472) );
  INVX1_HVT U880 ( .A(src_window[251]), .Y(DP_OP_422J2_124_3477_n2473) );
  INVX1_HVT U881 ( .A(src_window[248]), .Y(DP_OP_422J2_124_3477_n2476) );
  INVX1_HVT U882 ( .A(conv_weight_box[79]), .Y(DP_OP_422J2_124_3477_n2477) );
  INVX1_HVT U883 ( .A(conv_weight_box[78]), .Y(DP_OP_422J2_124_3477_n2478) );
  INVX1_HVT U884 ( .A(conv_weight_box[77]), .Y(DP_OP_422J2_124_3477_n2479) );
  INVX1_HVT U885 ( .A(conv_weight_box[76]), .Y(DP_OP_422J2_124_3477_n2480) );
  INVX1_HVT U886 ( .A(src_window[231]), .Y(DP_OP_422J2_124_3477_n2513) );
  INVX1_HVT U887 ( .A(src_window[230]), .Y(DP_OP_422J2_124_3477_n2514) );
  INVX1_HVT U888 ( .A(src_window[226]), .Y(DP_OP_422J2_124_3477_n2518) );
  INVX1_HVT U889 ( .A(src_window[224]), .Y(DP_OP_422J2_124_3477_n2520) );
  INVX1_HVT U890 ( .A(conv_weight_box[71]), .Y(DP_OP_422J2_124_3477_n2521) );
  INVX1_HVT U891 ( .A(conv_weight_box[70]), .Y(DP_OP_422J2_124_3477_n2522) );
  INVX1_HVT U892 ( .A(conv_weight_box[69]), .Y(DP_OP_422J2_124_3477_n2523) );
  INVX1_HVT U893 ( .A(conv_weight_box[68]), .Y(DP_OP_422J2_124_3477_n2524) );
  INVX1_HVT U894 ( .A(src_window[215]), .Y(DP_OP_422J2_124_3477_n2557) );
  INVX1_HVT U895 ( .A(src_window[214]), .Y(DP_OP_422J2_124_3477_n2558) );
  INVX1_HVT U896 ( .A(src_window[213]), .Y(DP_OP_422J2_124_3477_n2559) );
  INVX1_HVT U897 ( .A(src_window[212]), .Y(DP_OP_422J2_124_3477_n2560) );
  INVX1_HVT U898 ( .A(src_window[210]), .Y(DP_OP_422J2_124_3477_n2562) );
  INVX1_HVT U899 ( .A(src_window[209]), .Y(DP_OP_422J2_124_3477_n2563) );
  INVX1_HVT U900 ( .A(src_window[208]), .Y(DP_OP_422J2_124_3477_n2564) );
  INVX1_HVT U901 ( .A(conv_weight_box[62]), .Y(DP_OP_422J2_124_3477_n2566) );
  INVX1_HVT U902 ( .A(conv_weight_box[61]), .Y(DP_OP_422J2_124_3477_n2567) );
  INVX1_HVT U903 ( .A(conv_weight_box[60]), .Y(DP_OP_422J2_124_3477_n2568) );
  INVX1_HVT U904 ( .A(src_window[191]), .Y(DP_OP_422J2_124_3477_n2601) );
  INVX1_HVT U905 ( .A(src_window[190]), .Y(DP_OP_422J2_124_3477_n2602) );
  INVX1_HVT U906 ( .A(src_window[189]), .Y(DP_OP_422J2_124_3477_n2603) );
  INVX1_HVT U907 ( .A(src_window[188]), .Y(DP_OP_422J2_124_3477_n2604) );
  INVX1_HVT U908 ( .A(src_window[187]), .Y(DP_OP_422J2_124_3477_n2605) );
  INVX1_HVT U909 ( .A(src_window[186]), .Y(DP_OP_422J2_124_3477_n2606) );
  INVX1_HVT U910 ( .A(src_window[185]), .Y(DP_OP_422J2_124_3477_n2607) );
  INVX1_HVT U911 ( .A(src_window[184]), .Y(DP_OP_422J2_124_3477_n2608) );
  INVX1_HVT U912 ( .A(conv_weight_box[55]), .Y(DP_OP_422J2_124_3477_n2609) );
  INVX1_HVT U913 ( .A(conv_weight_box[54]), .Y(DP_OP_422J2_124_3477_n2610) );
  INVX1_HVT U914 ( .A(conv_weight_box[53]), .Y(DP_OP_422J2_124_3477_n2611) );
  INVX1_HVT U915 ( .A(conv_weight_box[52]), .Y(DP_OP_422J2_124_3477_n2612) );
  INVX1_HVT U916 ( .A(src_window[175]), .Y(DP_OP_422J2_124_3477_n2645) );
  INVX1_HVT U917 ( .A(src_window[174]), .Y(DP_OP_422J2_124_3477_n2646) );
  INVX1_HVT U918 ( .A(src_window[173]), .Y(DP_OP_422J2_124_3477_n2647) );
  INVX1_HVT U919 ( .A(src_window[172]), .Y(DP_OP_422J2_124_3477_n2648) );
  INVX1_HVT U920 ( .A(src_window[171]), .Y(DP_OP_422J2_124_3477_n2649) );
  INVX1_HVT U921 ( .A(src_window[170]), .Y(DP_OP_422J2_124_3477_n2650) );
  INVX1_HVT U922 ( .A(src_window[169]), .Y(DP_OP_422J2_124_3477_n2651) );
  INVX1_HVT U923 ( .A(src_window[168]), .Y(DP_OP_422J2_124_3477_n2652) );
  INVX1_HVT U924 ( .A(conv_weight_box[47]), .Y(DP_OP_422J2_124_3477_n2653) );
  INVX1_HVT U925 ( .A(conv_weight_box[46]), .Y(DP_OP_422J2_124_3477_n2654) );
  INVX1_HVT U926 ( .A(conv_weight_box[45]), .Y(DP_OP_422J2_124_3477_n2655) );
  INVX1_HVT U927 ( .A(conv_weight_box[44]), .Y(DP_OP_422J2_124_3477_n2656) );
  INVX1_HVT U928 ( .A(src_window[159]), .Y(DP_OP_422J2_124_3477_n2689) );
  INVX1_HVT U929 ( .A(src_window[158]), .Y(DP_OP_422J2_124_3477_n2690) );
  INVX1_HVT U930 ( .A(src_window[156]), .Y(DP_OP_422J2_124_3477_n2692) );
  INVX1_HVT U931 ( .A(src_window[154]), .Y(DP_OP_422J2_124_3477_n2694) );
  INVX1_HVT U932 ( .A(src_window[153]), .Y(DP_OP_422J2_124_3477_n2695) );
  INVX1_HVT U933 ( .A(src_window[152]), .Y(DP_OP_422J2_124_3477_n2696) );
  INVX1_HVT U934 ( .A(conv_weight_box[39]), .Y(DP_OP_422J2_124_3477_n2697) );
  INVX1_HVT U935 ( .A(DP_OP_425J2_127_3477_n3110), .Y(
        DP_OP_422J2_124_3477_n2698) );
  INVX1_HVT U936 ( .A(conv_weight_box[38]), .Y(DP_OP_422J2_124_3477_n2699) );
  INVX1_HVT U937 ( .A(conv_weight_box[37]), .Y(DP_OP_422J2_124_3477_n2700) );
  INVX1_HVT U938 ( .A(src_window[135]), .Y(DP_OP_422J2_124_3477_n2731) );
  INVX1_HVT U939 ( .A(src_window[134]), .Y(DP_OP_422J2_124_3477_n2732) );
  INVX1_HVT U940 ( .A(src_window[133]), .Y(DP_OP_422J2_124_3477_n2733) );
  INVX1_HVT U941 ( .A(src_window[132]), .Y(DP_OP_422J2_124_3477_n2734) );
  INVX1_HVT U942 ( .A(src_window[131]), .Y(DP_OP_422J2_124_3477_n2735) );
  INVX1_HVT U943 ( .A(src_window[130]), .Y(DP_OP_422J2_124_3477_n2736) );
  INVX1_HVT U944 ( .A(conv_weight_box[32]), .Y(DP_OP_422J2_124_3477_n2739) );
  INVX1_HVT U945 ( .A(conv_weight_box[31]), .Y(DP_OP_422J2_124_3477_n2740) );
  INVX1_HVT U946 ( .A(n428), .Y(DP_OP_422J2_124_3477_n2741) );
  INVX1_HVT U947 ( .A(conv_weight_box[30]), .Y(DP_OP_422J2_124_3477_n2742) );
  INVX1_HVT U948 ( .A(src_window[118]), .Y(DP_OP_422J2_124_3477_n2776) );
  INVX1_HVT U949 ( .A(src_window[117]), .Y(DP_OP_422J2_124_3477_n2777) );
  INVX1_HVT U950 ( .A(src_window[114]), .Y(DP_OP_422J2_124_3477_n2780) );
  INVX1_HVT U951 ( .A(src_window[113]), .Y(DP_OP_422J2_124_3477_n2781) );
  INVX1_HVT U952 ( .A(src_window[112]), .Y(DP_OP_422J2_124_3477_n2782) );
  INVX1_HVT U953 ( .A(conv_weight_box[24]), .Y(DP_OP_422J2_124_3477_n2784) );
  INVX1_HVT U954 ( .A(conv_weight_box[23]), .Y(DP_OP_422J2_124_3477_n2785) );
  INVX1_HVT U955 ( .A(conv_weight_box[22]), .Y(DP_OP_422J2_124_3477_n2786) );
  INVX1_HVT U956 ( .A(src_window[95]), .Y(DP_OP_422J2_124_3477_n2819) );
  INVX1_HVT U957 ( .A(src_window[94]), .Y(DP_OP_422J2_124_3477_n2820) );
  INVX1_HVT U958 ( .A(src_window[89]), .Y(DP_OP_422J2_124_3477_n2825) );
  INVX1_HVT U959 ( .A(conv_weight_box[17]), .Y(DP_OP_422J2_124_3477_n2827) );
  INVX1_HVT U960 ( .A(conv_weight_box[14]), .Y(DP_OP_422J2_124_3477_n2830) );
  INVX1_HVT U961 ( .A(src_window[78]), .Y(DP_OP_422J2_124_3477_n2864) );
  INVX1_HVT U962 ( .A(src_window[77]), .Y(DP_OP_422J2_124_3477_n2865) );
  INVX1_HVT U963 ( .A(src_window[74]), .Y(DP_OP_422J2_124_3477_n2868) );
  INVX1_HVT U964 ( .A(src_window[73]), .Y(DP_OP_422J2_124_3477_n2869) );
  INVX1_HVT U965 ( .A(src_window[72]), .Y(DP_OP_422J2_124_3477_n2870) );
  INVX1_HVT U966 ( .A(conv_weight_box[10]), .Y(DP_OP_422J2_124_3477_n2871) );
  INVX1_HVT U967 ( .A(conv_weight_box[9]), .Y(DP_OP_422J2_124_3477_n2872) );
  INVX1_HVT U968 ( .A(conv_weight_box[8]), .Y(DP_OP_422J2_124_3477_n2873) );
  INVX1_HVT U969 ( .A(src_window[62]), .Y(DP_OP_422J2_124_3477_n2908) );
  INVX1_HVT U970 ( .A(src_window[61]), .Y(DP_OP_422J2_124_3477_n2909) );
  INVX1_HVT U971 ( .A(src_window[58]), .Y(DP_OP_422J2_124_3477_n2912) );
  INVX1_HVT U972 ( .A(src_window[57]), .Y(DP_OP_422J2_124_3477_n2913) );
  INVX1_HVT U973 ( .A(conv_weight_box[1]), .Y(DP_OP_422J2_124_3477_n2916) );
  INVX1_HVT U974 ( .A(conv_weight_box[0]), .Y(DP_OP_422J2_124_3477_n2917) );
  INVX1_HVT U975 ( .A(n429), .Y(DP_OP_422J2_124_3477_n2918) );
  INVX1_HVT U976 ( .A(DP_OP_422J2_124_3477_n361), .Y(DP_OP_422J2_124_3477_n362) );
  INVX1_HVT U977 ( .A(DP_OP_422J2_124_3477_n671), .Y(DP_OP_422J2_124_3477_n672) );
  INVX1_HVT U978 ( .A(DP_OP_422J2_124_3477_n74), .Y(DP_OP_422J2_124_3477_n73)
         );
  INVX1_HVT U979 ( .A(DP_OP_424J2_126_3477_n67), .Y(DP_OP_424J2_126_3477_n69)
         );
  INVX1_HVT U980 ( .A(DP_OP_424J2_126_3477_n153), .Y(DP_OP_424J2_126_3477_n154) );
  INVX1_HVT U981 ( .A(DP_OP_424J2_126_3477_n155), .Y(DP_OP_424J2_126_3477_n156) );
  INVX1_HVT U982 ( .A(DP_OP_424J2_126_3477_n157), .Y(DP_OP_424J2_126_3477_n158) );
  INVX1_HVT U983 ( .A(DP_OP_424J2_126_3477_n1579), .Y(
        DP_OP_424J2_126_3477_n1580) );
  INVX1_HVT U984 ( .A(DP_OP_424J2_126_3477_n159), .Y(DP_OP_424J2_126_3477_n160) );
  INVX1_HVT U985 ( .A(DP_OP_424J2_126_3477_n161), .Y(DP_OP_424J2_126_3477_n162) );
  INVX1_HVT U986 ( .A(DP_OP_424J2_126_3477_n163), .Y(DP_OP_424J2_126_3477_n164) );
  INVX1_HVT U987 ( .A(DP_OP_424J2_126_3477_n165), .Y(DP_OP_424J2_126_3477_n166) );
  INVX1_HVT U988 ( .A(DP_OP_424J2_126_3477_n167), .Y(DP_OP_424J2_126_3477_n168) );
  INVX1_HVT U989 ( .A(DP_OP_424J2_126_3477_n169), .Y(DP_OP_424J2_126_3477_n170) );
  INVX1_HVT U990 ( .A(DP_OP_424J2_126_3477_n171), .Y(DP_OP_424J2_126_3477_n172) );
  INVX1_HVT U991 ( .A(DP_OP_424J2_126_3477_n173), .Y(DP_OP_424J2_126_3477_n174) );
  INVX1_HVT U992 ( .A(DP_OP_424J2_126_3477_n175), .Y(DP_OP_424J2_126_3477_n176) );
  INVX1_HVT U993 ( .A(DP_OP_424J2_126_3477_n177), .Y(DP_OP_424J2_126_3477_n178) );
  INVX1_HVT U994 ( .A(DP_OP_424J2_126_3477_n179), .Y(DP_OP_424J2_126_3477_n180) );
  INVX1_HVT U995 ( .A(DP_OP_424J2_126_3477_n181), .Y(DP_OP_424J2_126_3477_n182) );
  INVX1_HVT U996 ( .A(src_window[23]), .Y(DP_OP_424J2_126_3477_n1854) );
  INVX1_HVT U997 ( .A(src_window[20]), .Y(DP_OP_424J2_126_3477_n1857) );
  INVX1_HVT U998 ( .A(src_window[19]), .Y(DP_OP_424J2_126_3477_n1858) );
  INVX1_HVT U999 ( .A(conv_weight_box[6]), .Y(DP_OP_424J2_126_3477_n1862) );
  INVX1_HVT U1000 ( .A(conv_weight_box[3]), .Y(DP_OP_424J2_126_3477_n1865) );
  INVX1_HVT U1001 ( .A(src_window[39]), .Y(DP_OP_424J2_126_3477_n1898) );
  INVX1_HVT U1002 ( .A(DP_OP_424J2_126_3477_n189), .Y(
        DP_OP_424J2_126_3477_n190) );
  INVX1_HVT U1003 ( .A(src_window[36]), .Y(DP_OP_424J2_126_3477_n1901) );
  INVX1_HVT U1004 ( .A(src_window[34]), .Y(DP_OP_424J2_126_3477_n1903) );
  INVX1_HVT U1005 ( .A(src_window[33]), .Y(DP_OP_424J2_126_3477_n1904) );
  INVX1_HVT U1006 ( .A(conv_weight_box[13]), .Y(DP_OP_424J2_126_3477_n1906) );
  INVX1_HVT U1007 ( .A(n431), .Y(DP_OP_424J2_126_3477_n1907) );
  INVX1_HVT U1008 ( .A(conv_weight_box[12]), .Y(DP_OP_424J2_126_3477_n1908) );
  INVX1_HVT U1009 ( .A(conv_weight_box[11]), .Y(DP_OP_424J2_126_3477_n1909) );
  INVX1_HVT U1010 ( .A(src_window[63]), .Y(DP_OP_424J2_126_3477_n1942) );
  INVX1_HVT U1011 ( .A(src_window[57]), .Y(DP_OP_424J2_126_3477_n1948) );
  INVX1_HVT U1012 ( .A(src_window[56]), .Y(DP_OP_424J2_126_3477_n1949) );
  INVX1_HVT U1013 ( .A(conv_weight_box[21]), .Y(DP_OP_424J2_126_3477_n1950) );
  INVX1_HVT U1014 ( .A(conv_weight_box[19]), .Y(DP_OP_424J2_126_3477_n1952) );
  INVX1_HVT U1015 ( .A(conv_weight_box[18]), .Y(DP_OP_424J2_126_3477_n1953) );
  INVX1_HVT U1016 ( .A(src_window[79]), .Y(DP_OP_424J2_126_3477_n1986) );
  INVX1_HVT U1017 ( .A(src_window[77]), .Y(DP_OP_424J2_126_3477_n1988) );
  INVX1_HVT U1018 ( .A(conv_weight_box[29]), .Y(DP_OP_424J2_126_3477_n1994) );
  INVX1_HVT U1019 ( .A(conv_weight_box[28]), .Y(DP_OP_424J2_126_3477_n1995) );
  INVX1_HVT U1020 ( .A(conv_weight_box[27]), .Y(DP_OP_424J2_126_3477_n1996) );
  INVX1_HVT U1021 ( .A(src_window[93]), .Y(DP_OP_424J2_126_3477_n2032) );
  INVX1_HVT U1022 ( .A(src_window[92]), .Y(DP_OP_424J2_126_3477_n2033) );
  INVX1_HVT U1023 ( .A(src_window[91]), .Y(DP_OP_424J2_126_3477_n2034) );
  INVX1_HVT U1024 ( .A(src_window[90]), .Y(DP_OP_424J2_126_3477_n2035) );
  INVX1_HVT U1025 ( .A(src_window[88]), .Y(DP_OP_424J2_126_3477_n2037) );
  INVX1_HVT U1026 ( .A(conv_weight_box[36]), .Y(DP_OP_424J2_126_3477_n2038) );
  INVX1_HVT U1027 ( .A(conv_weight_box[35]), .Y(DP_OP_424J2_126_3477_n2039) );
  INVX1_HVT U1028 ( .A(conv_weight_box[34]), .Y(DP_OP_424J2_126_3477_n2040) );
  INVX1_HVT U1029 ( .A(conv_weight_box[33]), .Y(DP_OP_424J2_126_3477_n2041) );
  INVX1_HVT U1030 ( .A(src_window[119]), .Y(DP_OP_424J2_126_3477_n2074) );
  INVX1_HVT U1031 ( .A(src_window[116]), .Y(DP_OP_424J2_126_3477_n2077) );
  INVX1_HVT U1032 ( .A(src_window[115]), .Y(DP_OP_424J2_126_3477_n2078) );
  INVX1_HVT U1033 ( .A(conv_weight_box[43]), .Y(DP_OP_424J2_126_3477_n2082) );
  INVX1_HVT U1034 ( .A(conv_weight_box[41]), .Y(DP_OP_424J2_126_3477_n2084) );
  INVX1_HVT U1035 ( .A(conv_weight_box[40]), .Y(DP_OP_424J2_126_3477_n2085) );
  INVX1_HVT U1036 ( .A(src_window[135]), .Y(DP_OP_424J2_126_3477_n2118) );
  INVX1_HVT U1037 ( .A(src_window[134]), .Y(DP_OP_424J2_126_3477_n2119) );
  INVX1_HVT U1038 ( .A(src_window[133]), .Y(DP_OP_424J2_126_3477_n2120) );
  INVX1_HVT U1039 ( .A(src_window[129]), .Y(DP_OP_424J2_126_3477_n2124) );
  INVX1_HVT U1040 ( .A(src_window[128]), .Y(DP_OP_424J2_126_3477_n2125) );
  INVX1_HVT U1041 ( .A(conv_weight_box[51]), .Y(DP_OP_424J2_126_3477_n2126) );
  INVX1_HVT U1042 ( .A(conv_weight_box[50]), .Y(DP_OP_424J2_126_3477_n2127) );
  INVX1_HVT U1043 ( .A(conv_weight_box[48]), .Y(DP_OP_424J2_126_3477_n2129) );
  INVX1_HVT U1044 ( .A(src_window[158]), .Y(DP_OP_424J2_126_3477_n2163) );
  INVX1_HVT U1045 ( .A(src_window[157]), .Y(DP_OP_424J2_126_3477_n2164) );
  INVX1_HVT U1046 ( .A(src_window[153]), .Y(DP_OP_424J2_126_3477_n2168) );
  INVX1_HVT U1047 ( .A(conv_weight_box[59]), .Y(DP_OP_424J2_126_3477_n2170) );
  INVX1_HVT U1048 ( .A(conv_weight_box[58]), .Y(DP_OP_424J2_126_3477_n2171) );
  INVX1_HVT U1049 ( .A(conv_weight_box[56]), .Y(DP_OP_424J2_126_3477_n2173) );
  INVX1_HVT U1050 ( .A(src_window[170]), .Y(DP_OP_424J2_126_3477_n2211) );
  INVX1_HVT U1051 ( .A(src_window[169]), .Y(DP_OP_424J2_126_3477_n2212) );
  INVX1_HVT U1052 ( .A(conv_weight_box[65]), .Y(DP_OP_424J2_126_3477_n2216) );
  INVX1_HVT U1053 ( .A(conv_weight_box[75]), .Y(DP_OP_424J2_126_3477_n2258) );
  INVX1_HVT U1054 ( .A(conv_weight_box[73]), .Y(DP_OP_424J2_126_3477_n2260) );
  INVX1_HVT U1055 ( .A(src_window[213]), .Y(DP_OP_424J2_126_3477_n2296) );
  INVX1_HVT U1056 ( .A(conv_weight_box[83]), .Y(DP_OP_424J2_126_3477_n2302) );
  INVX1_HVT U1057 ( .A(conv_weight_box[81]), .Y(DP_OP_424J2_126_3477_n2304) );
  INVX1_HVT U1058 ( .A(src_window[231]), .Y(DP_OP_424J2_126_3477_n2338) );
  INVX1_HVT U1059 ( .A(src_window[230]), .Y(DP_OP_424J2_126_3477_n2339) );
  INVX1_HVT U1060 ( .A(src_window[228]), .Y(DP_OP_424J2_126_3477_n2341) );
  INVX1_HVT U1061 ( .A(src_window[227]), .Y(DP_OP_424J2_126_3477_n2342) );
  INVX1_HVT U1062 ( .A(src_window[225]), .Y(DP_OP_424J2_126_3477_n2344) );
  INVX1_HVT U1063 ( .A(conv_weight_box[87]), .Y(DP_OP_424J2_126_3477_n2349) );
  INVX1_HVT U1064 ( .A(src_window[237]), .Y(DP_OP_424J2_126_3477_n2381) );
  INVX1_HVT U1065 ( .A(src_window[236]), .Y(DP_OP_424J2_126_3477_n2382) );
  INVX1_HVT U1066 ( .A(src_window[235]), .Y(DP_OP_424J2_126_3477_n2383) );
  INVX1_HVT U1067 ( .A(src_window[234]), .Y(DP_OP_424J2_126_3477_n2384) );
  INVX1_HVT U1068 ( .A(src_window[233]), .Y(DP_OP_424J2_126_3477_n2385) );
  INVX1_HVT U1069 ( .A(src_window[232]), .Y(DP_OP_424J2_126_3477_n2386) );
  INVX1_HVT U1070 ( .A(conv_weight_box[93]), .Y(DP_OP_424J2_126_3477_n2387) );
  INVX1_HVT U1071 ( .A(conv_weight_box[92]), .Y(DP_OP_424J2_126_3477_n2388) );
  INVX1_HVT U1072 ( .A(conv_weight_box[91]), .Y(DP_OP_424J2_126_3477_n2389) );
  INVX1_HVT U1073 ( .A(n430), .Y(DP_OP_424J2_126_3477_n2390) );
  INVX1_HVT U1074 ( .A(src_window[223]), .Y(DP_OP_424J2_126_3477_n2423) );
  INVX1_HVT U1075 ( .A(src_window[218]), .Y(DP_OP_424J2_126_3477_n2428) );
  INVX1_HVT U1076 ( .A(src_window[216]), .Y(DP_OP_424J2_126_3477_n2430) );
  INVX1_HVT U1077 ( .A(conv_weight_box[86]), .Y(DP_OP_424J2_126_3477_n2432) );
  INVX1_HVT U1078 ( .A(src_window[203]), .Y(DP_OP_424J2_126_3477_n2471) );
  INVX1_HVT U1079 ( .A(src_window[202]), .Y(DP_OP_424J2_126_3477_n2472) );
  INVX1_HVT U1080 ( .A(src_window[200]), .Y(DP_OP_424J2_126_3477_n2474) );
  INVX1_HVT U1081 ( .A(conv_weight_box[79]), .Y(DP_OP_424J2_126_3477_n2475) );
  INVX1_HVT U1082 ( .A(conv_weight_box[76]), .Y(DP_OP_424J2_126_3477_n2478) );
  INVX1_HVT U1083 ( .A(src_window[182]), .Y(DP_OP_424J2_126_3477_n2512) );
  INVX1_HVT U1084 ( .A(src_window[177]), .Y(DP_OP_424J2_126_3477_n2517) );
  INVX1_HVT U1085 ( .A(conv_weight_box[70]), .Y(DP_OP_424J2_126_3477_n2520) );
  INVX1_HVT U1086 ( .A(conv_weight_box[69]), .Y(DP_OP_424J2_126_3477_n2521) );
  INVX1_HVT U1087 ( .A(conv_weight_box[68]), .Y(DP_OP_424J2_126_3477_n2522) );
  INVX1_HVT U1088 ( .A(src_window[167]), .Y(DP_OP_424J2_126_3477_n2555) );
  INVX1_HVT U1089 ( .A(src_window[165]), .Y(DP_OP_424J2_126_3477_n2557) );
  INVX1_HVT U1090 ( .A(src_window[163]), .Y(DP_OP_424J2_126_3477_n2559) );
  INVX1_HVT U1091 ( .A(src_window[161]), .Y(DP_OP_424J2_126_3477_n2561) );
  INVX1_HVT U1092 ( .A(conv_weight_box[63]), .Y(DP_OP_424J2_126_3477_n2563) );
  INVX1_HVT U1093 ( .A(conv_weight_box[61]), .Y(DP_OP_424J2_126_3477_n2565) );
  INVX1_HVT U1094 ( .A(conv_weight_box[60]), .Y(DP_OP_424J2_126_3477_n2566) );
  INVX1_HVT U1095 ( .A(src_window[142]), .Y(DP_OP_424J2_126_3477_n2600) );
  INVX1_HVT U1096 ( .A(src_window[138]), .Y(DP_OP_424J2_126_3477_n2604) );
  INVX1_HVT U1097 ( .A(conv_weight_box[55]), .Y(DP_OP_424J2_126_3477_n2607) );
  INVX1_HVT U1098 ( .A(conv_weight_box[54]), .Y(DP_OP_424J2_126_3477_n2608) );
  INVX1_HVT U1099 ( .A(conv_weight_box[53]), .Y(DP_OP_424J2_126_3477_n2609) );
  INVX1_HVT U1100 ( .A(conv_weight_box[52]), .Y(DP_OP_424J2_126_3477_n2610) );
  INVX1_HVT U1101 ( .A(src_window[126]), .Y(DP_OP_424J2_126_3477_n2644) );
  INVX1_HVT U1102 ( .A(src_window[121]), .Y(DP_OP_424J2_126_3477_n2649) );
  INVX1_HVT U1103 ( .A(src_window[120]), .Y(DP_OP_424J2_126_3477_n2650) );
  INVX1_HVT U1104 ( .A(conv_weight_box[47]), .Y(DP_OP_424J2_126_3477_n2651) );
  INVX1_HVT U1105 ( .A(conv_weight_box[46]), .Y(DP_OP_424J2_126_3477_n2652) );
  INVX1_HVT U1106 ( .A(conv_weight_box[45]), .Y(DP_OP_424J2_126_3477_n2653) );
  INVX1_HVT U1107 ( .A(conv_weight_box[44]), .Y(DP_OP_424J2_126_3477_n2654) );
  INVX1_HVT U1108 ( .A(src_window[109]), .Y(DP_OP_424J2_126_3477_n2689) );
  INVX1_HVT U1109 ( .A(src_window[107]), .Y(DP_OP_424J2_126_3477_n2691) );
  INVX1_HVT U1110 ( .A(src_window[105]), .Y(DP_OP_424J2_126_3477_n2693) );
  INVX1_HVT U1111 ( .A(conv_weight_box[39]), .Y(DP_OP_424J2_126_3477_n2695) );
  INVX1_HVT U1112 ( .A(DP_OP_425J2_127_3477_n3110), .Y(
        DP_OP_424J2_126_3477_n2696) );
  INVX1_HVT U1113 ( .A(conv_weight_box[38]), .Y(DP_OP_424J2_126_3477_n2697) );
  INVX1_HVT U1114 ( .A(conv_weight_box[37]), .Y(DP_OP_424J2_126_3477_n2698) );
  INVX1_HVT U1115 ( .A(src_window[87]), .Y(DP_OP_424J2_126_3477_n2731) );
  INVX1_HVT U1116 ( .A(src_window[86]), .Y(DP_OP_424J2_126_3477_n2732) );
  INVX1_HVT U1117 ( .A(src_window[85]), .Y(DP_OP_424J2_126_3477_n2733) );
  INVX1_HVT U1118 ( .A(src_window[84]), .Y(DP_OP_424J2_126_3477_n2734) );
  INVX1_HVT U1119 ( .A(src_window[83]), .Y(DP_OP_424J2_126_3477_n2735) );
  INVX1_HVT U1120 ( .A(src_window[82]), .Y(DP_OP_424J2_126_3477_n2736) );
  INVX1_HVT U1121 ( .A(src_window[81]), .Y(DP_OP_424J2_126_3477_n2737) );
  INVX1_HVT U1122 ( .A(src_window[80]), .Y(DP_OP_424J2_126_3477_n2738) );
  INVX1_HVT U1123 ( .A(conv_weight_box[31]), .Y(DP_OP_424J2_126_3477_n2740) );
  INVX1_HVT U1124 ( .A(n428), .Y(DP_OP_424J2_126_3477_n2741) );
  INVX1_HVT U1125 ( .A(conv_weight_box[30]), .Y(DP_OP_424J2_126_3477_n2742) );
  INVX1_HVT U1126 ( .A(src_window[71]), .Y(DP_OP_424J2_126_3477_n2775) );
  INVX1_HVT U1127 ( .A(src_window[69]), .Y(DP_OP_424J2_126_3477_n2777) );
  INVX1_HVT U1128 ( .A(conv_weight_box[25]), .Y(DP_OP_424J2_126_3477_n2783) );
  INVX1_HVT U1129 ( .A(conv_weight_box[24]), .Y(DP_OP_424J2_126_3477_n2784) );
  INVX1_HVT U1130 ( .A(conv_weight_box[23]), .Y(DP_OP_424J2_126_3477_n2785) );
  INVX1_HVT U1131 ( .A(src_window[47]), .Y(DP_OP_424J2_126_3477_n2819) );
  INVX1_HVT U1132 ( .A(src_window[46]), .Y(DP_OP_424J2_126_3477_n2820) );
  INVX1_HVT U1133 ( .A(src_window[45]), .Y(DP_OP_424J2_126_3477_n2821) );
  INVX1_HVT U1134 ( .A(src_window[44]), .Y(DP_OP_424J2_126_3477_n2822) );
  INVX1_HVT U1135 ( .A(src_window[43]), .Y(DP_OP_424J2_126_3477_n2823) );
  INVX1_HVT U1136 ( .A(src_window[42]), .Y(DP_OP_424J2_126_3477_n2824) );
  INVX1_HVT U1137 ( .A(src_window[41]), .Y(DP_OP_424J2_126_3477_n2825) );
  INVX1_HVT U1138 ( .A(src_window[40]), .Y(DP_OP_424J2_126_3477_n2826) );
  INVX1_HVT U1139 ( .A(conv_weight_box[17]), .Y(DP_OP_424J2_126_3477_n2827) );
  INVX1_HVT U1140 ( .A(conv_weight_box[16]), .Y(DP_OP_424J2_126_3477_n2828) );
  INVX1_HVT U1141 ( .A(conv_weight_box[15]), .Y(DP_OP_424J2_126_3477_n2829) );
  INVX1_HVT U1142 ( .A(conv_weight_box[14]), .Y(DP_OP_424J2_126_3477_n2830) );
  INVX1_HVT U1143 ( .A(src_window[31]), .Y(DP_OP_424J2_126_3477_n2863) );
  INVX1_HVT U1144 ( .A(src_window[30]), .Y(DP_OP_424J2_126_3477_n2864) );
  INVX1_HVT U1145 ( .A(src_window[29]), .Y(DP_OP_424J2_126_3477_n2865) );
  INVX1_HVT U1146 ( .A(src_window[27]), .Y(DP_OP_424J2_126_3477_n2867) );
  INVX1_HVT U1147 ( .A(src_window[25]), .Y(DP_OP_424J2_126_3477_n2869) );
  INVX1_HVT U1148 ( .A(conv_weight_box[8]), .Y(DP_OP_424J2_126_3477_n2873) );
  INVX1_HVT U1149 ( .A(conv_weight_box[7]), .Y(DP_OP_424J2_126_3477_n2874) );
  INVX1_HVT U1150 ( .A(src_window[13]), .Y(DP_OP_424J2_126_3477_n2909) );
  INVX1_HVT U1151 ( .A(src_window[12]), .Y(DP_OP_424J2_126_3477_n2910) );
  INVX1_HVT U1152 ( .A(src_window[10]), .Y(DP_OP_424J2_126_3477_n2912) );
  INVX1_HVT U1153 ( .A(conv_weight_box[2]), .Y(DP_OP_424J2_126_3477_n2915) );
  INVX1_HVT U1154 ( .A(conv_weight_box[0]), .Y(DP_OP_424J2_126_3477_n2917) );
  INVX1_HVT U1155 ( .A(DP_OP_424J2_126_3477_n361), .Y(
        DP_OP_424J2_126_3477_n362) );
  INVX1_HVT U1156 ( .A(DP_OP_424J2_126_3477_n671), .Y(
        DP_OP_424J2_126_3477_n672) );
  INVX1_HVT U1157 ( .A(DP_OP_424J2_126_3477_n74), .Y(DP_OP_424J2_126_3477_n73)
         );
  INVX1_HVT U1158 ( .A(DP_OP_425J2_127_3477_n67), .Y(DP_OP_425J2_127_3477_n69)
         );
  INVX1_HVT U1159 ( .A(DP_OP_425J2_127_3477_n153), .Y(
        DP_OP_425J2_127_3477_n154) );
  INVX1_HVT U1160 ( .A(DP_OP_425J2_127_3477_n155), .Y(
        DP_OP_425J2_127_3477_n156) );
  INVX1_HVT U1161 ( .A(DP_OP_425J2_127_3477_n157), .Y(
        DP_OP_425J2_127_3477_n158) );
  INVX1_HVT U1162 ( .A(DP_OP_425J2_127_3477_n1579), .Y(
        DP_OP_425J2_127_3477_n1580) );
  INVX1_HVT U1163 ( .A(DP_OP_425J2_127_3477_n159), .Y(
        DP_OP_425J2_127_3477_n160) );
  INVX1_HVT U1164 ( .A(DP_OP_425J2_127_3477_n161), .Y(
        DP_OP_425J2_127_3477_n162) );
  INVX1_HVT U1165 ( .A(DP_OP_425J2_127_3477_n163), .Y(
        DP_OP_425J2_127_3477_n164) );
  INVX1_HVT U1166 ( .A(DP_OP_425J2_127_3477_n165), .Y(
        DP_OP_425J2_127_3477_n166) );
  INVX1_HVT U1167 ( .A(DP_OP_425J2_127_3477_n167), .Y(
        DP_OP_425J2_127_3477_n168) );
  INVX1_HVT U1168 ( .A(DP_OP_425J2_127_3477_n169), .Y(
        DP_OP_425J2_127_3477_n170) );
  INVX1_HVT U1169 ( .A(DP_OP_425J2_127_3477_n171), .Y(
        DP_OP_425J2_127_3477_n172) );
  INVX1_HVT U1170 ( .A(DP_OP_425J2_127_3477_n173), .Y(
        DP_OP_425J2_127_3477_n174) );
  INVX1_HVT U1171 ( .A(DP_OP_425J2_127_3477_n175), .Y(
        DP_OP_425J2_127_3477_n176) );
  INVX1_HVT U1172 ( .A(DP_OP_425J2_127_3477_n177), .Y(
        DP_OP_425J2_127_3477_n178) );
  INVX1_HVT U1173 ( .A(DP_OP_425J2_127_3477_n179), .Y(
        DP_OP_425J2_127_3477_n180) );
  INVX1_HVT U1174 ( .A(DP_OP_425J2_127_3477_n181), .Y(
        DP_OP_425J2_127_3477_n182) );
  INVX1_HVT U1175 ( .A(src_window[15]), .Y(DP_OP_425J2_127_3477_n1854) );
  INVX1_HVT U1176 ( .A(src_window[14]), .Y(DP_OP_425J2_127_3477_n1855) );
  INVX1_HVT U1177 ( .A(src_window[11]), .Y(DP_OP_425J2_127_3477_n1858) );
  INVX1_HVT U1178 ( .A(src_window[9]), .Y(DP_OP_425J2_127_3477_n1860) );
  INVX1_HVT U1179 ( .A(src_window[8]), .Y(DP_OP_425J2_127_3477_n1861) );
  INVX1_HVT U1180 ( .A(conv_weight_box[6]), .Y(DP_OP_425J2_127_3477_n1862) );
  INVX1_HVT U1181 ( .A(conv_weight_box[5]), .Y(DP_OP_425J2_127_3477_n1863) );
  INVX1_HVT U1182 ( .A(conv_weight_box[4]), .Y(DP_OP_425J2_127_3477_n1864) );
  INVX1_HVT U1183 ( .A(DP_OP_425J2_127_3477_n189), .Y(
        DP_OP_425J2_127_3477_n190) );
  INVX1_HVT U1184 ( .A(src_window[28]), .Y(DP_OP_425J2_127_3477_n1901) );
  INVX1_HVT U1185 ( .A(src_window[26]), .Y(DP_OP_425J2_127_3477_n1903) );
  INVX1_HVT U1186 ( .A(src_window[24]), .Y(DP_OP_425J2_127_3477_n1905) );
  INVX1_HVT U1187 ( .A(n431), .Y(DP_OP_425J2_127_3477_n1907) );
  INVX1_HVT U1188 ( .A(src_window[52]), .Y(DP_OP_425J2_127_3477_n1945) );
  INVX1_HVT U1189 ( .A(conv_weight_box[21]), .Y(DP_OP_425J2_127_3477_n1950) );
  INVX1_HVT U1190 ( .A(conv_weight_box[20]), .Y(DP_OP_425J2_127_3477_n1951) );
  INVX1_HVT U1191 ( .A(conv_weight_box[18]), .Y(DP_OP_425J2_127_3477_n1953) );
  INVX1_HVT U1192 ( .A(src_window[68]), .Y(DP_OP_425J2_127_3477_n1989) );
  INVX1_HVT U1193 ( .A(src_window[67]), .Y(DP_OP_425J2_127_3477_n1990) );
  INVX1_HVT U1194 ( .A(src_window[66]), .Y(DP_OP_425J2_127_3477_n1991) );
  INVX1_HVT U1195 ( .A(src_window[65]), .Y(DP_OP_425J2_127_3477_n1992) );
  INVX1_HVT U1196 ( .A(conv_weight_box[28]), .Y(DP_OP_425J2_127_3477_n1995) );
  INVX1_HVT U1197 ( .A(conv_weight_box[26]), .Y(DP_OP_425J2_127_3477_n1997) );
  INVX1_HVT U1198 ( .A(src_window[84]), .Y(DP_OP_425J2_127_3477_n2033) );
  INVX1_HVT U1199 ( .A(conv_weight_box[35]), .Y(DP_OP_425J2_127_3477_n2039) );
  INVX1_HVT U1200 ( .A(conv_weight_box[34]), .Y(DP_OP_425J2_127_3477_n2040) );
  INVX1_HVT U1201 ( .A(conv_weight_box[33]), .Y(DP_OP_425J2_127_3477_n2041) );
  INVX1_HVT U1202 ( .A(src_window[111]), .Y(DP_OP_425J2_127_3477_n2074) );
  INVX1_HVT U1203 ( .A(src_window[110]), .Y(DP_OP_425J2_127_3477_n2075) );
  INVX1_HVT U1204 ( .A(src_window[108]), .Y(DP_OP_425J2_127_3477_n2077) );
  INVX1_HVT U1205 ( .A(src_window[107]), .Y(DP_OP_425J2_127_3477_n2078) );
  INVX1_HVT U1206 ( .A(src_window[106]), .Y(DP_OP_425J2_127_3477_n2079) );
  INVX1_HVT U1207 ( .A(conv_weight_box[42]), .Y(DP_OP_425J2_127_3477_n2083) );
  INVX1_HVT U1208 ( .A(conv_weight_box[41]), .Y(DP_OP_425J2_127_3477_n2084) );
  INVX1_HVT U1209 ( .A(src_window[127]), .Y(DP_OP_425J2_127_3477_n2118) );
  INVX1_HVT U1210 ( .A(src_window[126]), .Y(DP_OP_425J2_127_3477_n2119) );
  INVX1_HVT U1211 ( .A(src_window[125]), .Y(DP_OP_425J2_127_3477_n2120) );
  INVX1_HVT U1212 ( .A(src_window[123]), .Y(DP_OP_425J2_127_3477_n2122) );
  INVX1_HVT U1213 ( .A(conv_weight_box[51]), .Y(DP_OP_425J2_127_3477_n2126) );
  INVX1_HVT U1214 ( .A(conv_weight_box[50]), .Y(DP_OP_425J2_127_3477_n2127) );
  INVX1_HVT U1215 ( .A(conv_weight_box[49]), .Y(DP_OP_425J2_127_3477_n2128) );
  INVX1_HVT U1216 ( .A(conv_weight_box[48]), .Y(DP_OP_425J2_127_3477_n2129) );
  INVX1_HVT U1217 ( .A(src_window[151]), .Y(DP_OP_425J2_127_3477_n2162) );
  INVX1_HVT U1218 ( .A(src_window[150]), .Y(DP_OP_425J2_127_3477_n2163) );
  INVX1_HVT U1219 ( .A(src_window[149]), .Y(DP_OP_425J2_127_3477_n2164) );
  INVX1_HVT U1220 ( .A(src_window[147]), .Y(DP_OP_425J2_127_3477_n2166) );
  INVX1_HVT U1221 ( .A(src_window[145]), .Y(DP_OP_425J2_127_3477_n2168) );
  INVX1_HVT U1222 ( .A(src_window[144]), .Y(DP_OP_425J2_127_3477_n2169) );
  INVX1_HVT U1223 ( .A(conv_weight_box[57]), .Y(DP_OP_425J2_127_3477_n2172) );
  INVX1_HVT U1224 ( .A(conv_weight_box[56]), .Y(DP_OP_425J2_127_3477_n2173) );
  INVX1_HVT U1225 ( .A(src_window[164]), .Y(DP_OP_425J2_127_3477_n2209) );
  INVX1_HVT U1226 ( .A(src_window[160]), .Y(DP_OP_425J2_127_3477_n2213) );
  INVX1_HVT U1227 ( .A(conv_weight_box[67]), .Y(DP_OP_425J2_127_3477_n2214) );
  INVX1_HVT U1228 ( .A(conv_weight_box[66]), .Y(DP_OP_425J2_127_3477_n2215) );
  INVX1_HVT U1229 ( .A(conv_weight_box[64]), .Y(DP_OP_425J2_127_3477_n2217) );
  INVX1_HVT U1230 ( .A(src_window[183]), .Y(DP_OP_425J2_127_3477_n2250) );
  INVX1_HVT U1231 ( .A(src_window[181]), .Y(DP_OP_425J2_127_3477_n2252) );
  INVX1_HVT U1232 ( .A(src_window[178]), .Y(DP_OP_425J2_127_3477_n2255) );
  INVX1_HVT U1233 ( .A(conv_weight_box[74]), .Y(DP_OP_425J2_127_3477_n2259) );
  INVX1_HVT U1234 ( .A(conv_weight_box[73]), .Y(DP_OP_425J2_127_3477_n2260) );
  INVX1_HVT U1235 ( .A(conv_weight_box[72]), .Y(DP_OP_425J2_127_3477_n2261) );
  INVX1_HVT U1236 ( .A(src_window[207]), .Y(DP_OP_425J2_127_3477_n2294) );
  INVX1_HVT U1237 ( .A(src_window[205]), .Y(DP_OP_425J2_127_3477_n2296) );
  INVX1_HVT U1238 ( .A(src_window[204]), .Y(DP_OP_425J2_127_3477_n2297) );
  INVX1_HVT U1239 ( .A(src_window[201]), .Y(DP_OP_425J2_127_3477_n2300) );
  INVX1_HVT U1240 ( .A(conv_weight_box[83]), .Y(DP_OP_425J2_127_3477_n2302) );
  INVX1_HVT U1241 ( .A(conv_weight_box[81]), .Y(DP_OP_425J2_127_3477_n2304) );
  INVX1_HVT U1242 ( .A(conv_weight_box[80]), .Y(DP_OP_425J2_127_3477_n2305) );
  INVX1_HVT U1243 ( .A(src_window[222]), .Y(DP_OP_425J2_127_3477_n2339) );
  INVX1_HVT U1244 ( .A(src_window[221]), .Y(DP_OP_425J2_127_3477_n2340) );
  INVX1_HVT U1245 ( .A(src_window[220]), .Y(DP_OP_425J2_127_3477_n2341) );
  INVX1_HVT U1246 ( .A(src_window[219]), .Y(DP_OP_425J2_127_3477_n2342) );
  INVX1_HVT U1247 ( .A(conv_weight_box[90]), .Y(DP_OP_425J2_127_3477_n2346) );
  INVX1_HVT U1248 ( .A(conv_weight_box[89]), .Y(DP_OP_425J2_127_3477_n2347) );
  INVX1_HVT U1249 ( .A(conv_weight_box[88]), .Y(DP_OP_425J2_127_3477_n2348) );
  INVX1_HVT U1250 ( .A(conv_weight_box[87]), .Y(DP_OP_425J2_127_3477_n2349) );
  INVX1_HVT U1251 ( .A(src_window[229]), .Y(DP_OP_425J2_127_3477_n2381) );
  INVX1_HVT U1252 ( .A(src_window[228]), .Y(DP_OP_425J2_127_3477_n2382) );
  INVX1_HVT U1253 ( .A(src_window[227]), .Y(DP_OP_425J2_127_3477_n2383) );
  INVX1_HVT U1254 ( .A(src_window[226]), .Y(DP_OP_425J2_127_3477_n2384) );
  INVX1_HVT U1255 ( .A(src_window[224]), .Y(DP_OP_425J2_127_3477_n2386) );
  INVX1_HVT U1256 ( .A(conv_weight_box[93]), .Y(DP_OP_425J2_127_3477_n2387) );
  INVX1_HVT U1257 ( .A(src_window[215]), .Y(DP_OP_425J2_127_3477_n2423) );
  INVX1_HVT U1258 ( .A(src_window[214]), .Y(DP_OP_425J2_127_3477_n2424) );
  INVX1_HVT U1259 ( .A(src_window[211]), .Y(DP_OP_425J2_127_3477_n2427) );
  INVX1_HVT U1260 ( .A(src_window[210]), .Y(DP_OP_425J2_127_3477_n2428) );
  INVX1_HVT U1261 ( .A(src_window[209]), .Y(DP_OP_425J2_127_3477_n2429) );
  INVX1_HVT U1262 ( .A(src_window[208]), .Y(DP_OP_425J2_127_3477_n2430) );
  INVX1_HVT U1263 ( .A(DP_OP_425J2_127_3477_n3255), .Y(
        DP_OP_425J2_127_3477_n2431) );
  INVX1_HVT U1264 ( .A(conv_weight_box[85]), .Y(DP_OP_425J2_127_3477_n2433) );
  INVX1_HVT U1265 ( .A(conv_weight_box[84]), .Y(DP_OP_425J2_127_3477_n2434) );
  INVX1_HVT U1266 ( .A(src_window[197]), .Y(DP_OP_425J2_127_3477_n2469) );
  INVX1_HVT U1267 ( .A(src_window[194]), .Y(DP_OP_425J2_127_3477_n2472) );
  INVX1_HVT U1268 ( .A(conv_weight_box[79]), .Y(DP_OP_425J2_127_3477_n2475) );
  INVX1_HVT U1269 ( .A(conv_weight_box[78]), .Y(DP_OP_425J2_127_3477_n2476) );
  INVX1_HVT U1270 ( .A(conv_weight_box[77]), .Y(DP_OP_425J2_127_3477_n2477) );
  INVX1_HVT U1271 ( .A(src_window[175]), .Y(DP_OP_425J2_127_3477_n2511) );
  INVX1_HVT U1272 ( .A(src_window[168]), .Y(DP_OP_425J2_127_3477_n2518) );
  INVX1_HVT U1273 ( .A(conv_weight_box[71]), .Y(DP_OP_425J2_127_3477_n2519) );
  INVX1_HVT U1274 ( .A(src_window[159]), .Y(DP_OP_425J2_127_3477_n2555) );
  INVX1_HVT U1275 ( .A(src_window[157]), .Y(DP_OP_425J2_127_3477_n2557) );
  INVX1_HVT U1276 ( .A(src_window[156]), .Y(DP_OP_425J2_127_3477_n2558) );
  INVX1_HVT U1277 ( .A(src_window[155]), .Y(DP_OP_425J2_127_3477_n2559) );
  INVX1_HVT U1278 ( .A(conv_weight_box[63]), .Y(DP_OP_425J2_127_3477_n2563) );
  INVX1_HVT U1279 ( .A(conv_weight_box[62]), .Y(DP_OP_425J2_127_3477_n2564) );
  INVX1_HVT U1280 ( .A(conv_weight_box[61]), .Y(DP_OP_425J2_127_3477_n2565) );
  INVX1_HVT U1281 ( .A(conv_weight_box[60]), .Y(DP_OP_425J2_127_3477_n2566) );
  INVX1_HVT U1282 ( .A(conv_weight_box[52]), .Y(DP_OP_425J2_127_3477_n2610) );
  INVX1_HVT U1283 ( .A(src_window[119]), .Y(DP_OP_425J2_127_3477_n2643) );
  INVX1_HVT U1284 ( .A(src_window[118]), .Y(DP_OP_425J2_127_3477_n2644) );
  INVX1_HVT U1285 ( .A(src_window[116]), .Y(DP_OP_425J2_127_3477_n2646) );
  INVX1_HVT U1286 ( .A(src_window[113]), .Y(DP_OP_425J2_127_3477_n2649) );
  INVX1_HVT U1287 ( .A(src_window[112]), .Y(DP_OP_425J2_127_3477_n2650) );
  INVX1_HVT U1288 ( .A(conv_weight_box[46]), .Y(DP_OP_425J2_127_3477_n2652) );
  INVX1_HVT U1289 ( .A(conv_weight_box[44]), .Y(DP_OP_425J2_127_3477_n2654) );
  INVX1_HVT U1290 ( .A(src_window[102]), .Y(DP_OP_425J2_127_3477_n2688) );
  INVX1_HVT U1291 ( .A(src_window[100]), .Y(DP_OP_425J2_127_3477_n2690) );
  INVX1_HVT U1292 ( .A(src_window[99]), .Y(DP_OP_425J2_127_3477_n2691) );
  INVX1_HVT U1293 ( .A(src_window[98]), .Y(DP_OP_425J2_127_3477_n2692) );
  INVX1_HVT U1294 ( .A(src_window[96]), .Y(DP_OP_425J2_127_3477_n2694) );
  INVX1_HVT U1295 ( .A(DP_OP_425J2_127_3477_n3110), .Y(
        DP_OP_425J2_127_3477_n2696) );
  INVX1_HVT U1296 ( .A(src_window[78]), .Y(DP_OP_425J2_127_3477_n2732) );
  INVX1_HVT U1297 ( .A(src_window[76]), .Y(DP_OP_425J2_127_3477_n2734) );
  INVX1_HVT U1298 ( .A(src_window[75]), .Y(DP_OP_425J2_127_3477_n2735) );
  INVX1_HVT U1299 ( .A(src_window[72]), .Y(DP_OP_425J2_127_3477_n2738) );
  INVX1_HVT U1300 ( .A(conv_weight_box[32]), .Y(DP_OP_425J2_127_3477_n2739) );
  INVX1_HVT U1301 ( .A(conv_weight_box[31]), .Y(DP_OP_425J2_127_3477_n2740) );
  INVX1_HVT U1302 ( .A(n428), .Y(DP_OP_425J2_127_3477_n2741) );
  INVX1_HVT U1303 ( .A(src_window[61]), .Y(DP_OP_425J2_127_3477_n2777) );
  INVX1_HVT U1304 ( .A(src_window[60]), .Y(DP_OP_425J2_127_3477_n2778) );
  INVX1_HVT U1305 ( .A(src_window[59]), .Y(DP_OP_425J2_127_3477_n2779) );
  INVX1_HVT U1306 ( .A(src_window[58]), .Y(DP_OP_425J2_127_3477_n2780) );
  INVX1_HVT U1307 ( .A(conv_weight_box[25]), .Y(DP_OP_425J2_127_3477_n2783) );
  INVX1_HVT U1308 ( .A(conv_weight_box[23]), .Y(DP_OP_425J2_127_3477_n2785) );
  INVX1_HVT U1309 ( .A(conv_weight_box[22]), .Y(DP_OP_425J2_127_3477_n2786) );
  INVX1_HVT U1310 ( .A(src_window[38]), .Y(DP_OP_425J2_127_3477_n2820) );
  INVX1_HVT U1311 ( .A(src_window[37]), .Y(DP_OP_425J2_127_3477_n2821) );
  INVX1_HVT U1312 ( .A(src_window[35]), .Y(DP_OP_425J2_127_3477_n2823) );
  INVX1_HVT U1313 ( .A(src_window[32]), .Y(DP_OP_425J2_127_3477_n2826) );
  INVX1_HVT U1314 ( .A(conv_weight_box[17]), .Y(DP_OP_425J2_127_3477_n2827) );
  INVX1_HVT U1315 ( .A(conv_weight_box[16]), .Y(DP_OP_425J2_127_3477_n2828) );
  INVX1_HVT U1316 ( .A(conv_weight_box[15]), .Y(DP_OP_425J2_127_3477_n2829) );
  INVX1_HVT U1317 ( .A(conv_weight_box[14]), .Y(DP_OP_425J2_127_3477_n2830) );
  INVX1_HVT U1318 ( .A(src_window[22]), .Y(DP_OP_425J2_127_3477_n2864) );
  INVX1_HVT U1319 ( .A(src_window[21]), .Y(DP_OP_425J2_127_3477_n2865) );
  INVX1_HVT U1320 ( .A(src_window[18]), .Y(DP_OP_425J2_127_3477_n2868) );
  INVX1_HVT U1321 ( .A(src_window[17]), .Y(DP_OP_425J2_127_3477_n2869) );
  INVX1_HVT U1322 ( .A(src_window[16]), .Y(DP_OP_425J2_127_3477_n2870) );
  INVX1_HVT U1323 ( .A(conv_weight_box[10]), .Y(DP_OP_425J2_127_3477_n2871) );
  INVX1_HVT U1324 ( .A(conv_weight_box[9]), .Y(DP_OP_425J2_127_3477_n2872) );
  INVX1_HVT U1325 ( .A(conv_weight_box[7]), .Y(DP_OP_425J2_127_3477_n2874) );
  INVX1_HVT U1326 ( .A(src_window[7]), .Y(DP_OP_425J2_127_3477_n2907) );
  INVX1_HVT U1327 ( .A(src_window[6]), .Y(DP_OP_425J2_127_3477_n2908) );
  INVX1_HVT U1328 ( .A(src_window[5]), .Y(DP_OP_425J2_127_3477_n2909) );
  INVX1_HVT U1329 ( .A(src_window[4]), .Y(DP_OP_425J2_127_3477_n2910) );
  INVX1_HVT U1330 ( .A(src_window[3]), .Y(DP_OP_425J2_127_3477_n2911) );
  INVX1_HVT U1331 ( .A(src_window[2]), .Y(DP_OP_425J2_127_3477_n2912) );
  INVX1_HVT U1332 ( .A(src_window[1]), .Y(DP_OP_425J2_127_3477_n2913) );
  INVX1_HVT U1333 ( .A(src_window[0]), .Y(DP_OP_425J2_127_3477_n2914) );
  INVX1_HVT U1334 ( .A(conv_weight_box[2]), .Y(DP_OP_425J2_127_3477_n2915) );
  INVX1_HVT U1335 ( .A(conv_weight_box[1]), .Y(DP_OP_425J2_127_3477_n2916) );
  INVX1_HVT U1336 ( .A(conv_weight_box[0]), .Y(DP_OP_425J2_127_3477_n2917) );
  INVX1_HVT U1337 ( .A(n429), .Y(DP_OP_425J2_127_3477_n2918) );
  INVX1_HVT U1338 ( .A(DP_OP_425J2_127_3477_n361), .Y(
        DP_OP_425J2_127_3477_n362) );
  INVX1_HVT U1339 ( .A(DP_OP_425J2_127_3477_n671), .Y(
        DP_OP_425J2_127_3477_n672) );
  INVX1_HVT U1340 ( .A(DP_OP_425J2_127_3477_n74), .Y(DP_OP_425J2_127_3477_n73)
         );
  MUX21X1_HVT U1341 ( .A1(tmp_big2[20]), .A2(tmp_big1[20]), .S0(n357), .Y(
        data_out[20]) );
  MUX21X1_HVT U1342 ( .A1(tmp_big2[21]), .A2(tmp_big1[21]), .S0(n354), .Y(
        data_out[21]) );
  MUX21X1_HVT U1343 ( .A1(tmp_big2[22]), .A2(tmp_big1[22]), .S0(n355), .Y(
        data_out[22]) );
  MUX21X1_HVT U1344 ( .A1(tmp_big2[23]), .A2(tmp_big1[23]), .S0(n356), .Y(
        data_out[23]) );
  MUX21X1_HVT U1345 ( .A1(tmp_big2[24]), .A2(tmp_big1[24]), .S0(n357), .Y(
        data_out[24]) );
  MUX21X1_HVT U1346 ( .A1(tmp_big2[25]), .A2(tmp_big1[25]), .S0(n354), .Y(
        data_out[25]) );
  MUX21X1_HVT U1347 ( .A1(tmp_big2[26]), .A2(tmp_big1[26]), .S0(n355), .Y(
        data_out[26]) );
  MUX21X1_HVT U1348 ( .A1(tmp_big2[27]), .A2(tmp_big1[27]), .S0(n356), .Y(
        data_out[27]) );
  MUX21X1_HVT U1349 ( .A1(tmp_big2[28]), .A2(tmp_big1[28]), .S0(n357), .Y(
        data_out[28]) );
  MUX21X1_HVT U1350 ( .A1(tmp_big2[29]), .A2(tmp_big1[29]), .S0(n354), .Y(
        data_out[29]) );
  MUX21X1_HVT U1351 ( .A1(tmp_big2[30]), .A2(tmp_big1[30]), .S0(n355), .Y(
        data_out[30]) );
  MUX21X1_HVT U1352 ( .A1(tmp_big2[31]), .A2(tmp_big1[31]), .S0(n356), .Y(
        data_out[31]) );
  MUX21X1_HVT U1353 ( .A1(tmp_big2[6]), .A2(tmp_big1[6]), .S0(n357), .Y(
        data_out[6]) );
  MUX21X1_HVT U1354 ( .A1(conv2_sum_b[31]), .A2(conv2_sum_a[31]), .S0(n362), 
        .Y(tmp_big1[31]) );
  MUX21X1_HVT U1355 ( .A1(tmp_big2[5]), .A2(tmp_big1[5]), .S0(n354), .Y(
        data_out[5]) );
  MUX21X1_HVT U1356 ( .A1(tmp_big2[7]), .A2(tmp_big1[7]), .S0(n356), .Y(
        data_out[7]) );
  MUX21X1_HVT U1357 ( .A1(tmp_big2[8]), .A2(tmp_big1[8]), .S0(n356), .Y(
        data_out[8]) );
  MUX21X1_HVT U1358 ( .A1(tmp_big2[9]), .A2(tmp_big1[9]), .S0(n354), .Y(
        data_out[9]) );
  MUX21X1_HVT U1359 ( .A1(tmp_big2[12]), .A2(tmp_big1[12]), .S0(n355), .Y(
        data_out[12]) );
  MUX21X1_HVT U1360 ( .A1(tmp_big2[13]), .A2(tmp_big1[13]), .S0(n354), .Y(
        data_out[13]) );
  MUX21X1_HVT U1361 ( .A1(tmp_big2[10]), .A2(tmp_big1[10]), .S0(n356), .Y(
        data_out[10]) );
  MUX21X1_HVT U1362 ( .A1(tmp_big2[11]), .A2(tmp_big1[11]), .S0(n355), .Y(
        data_out[11]) );
  MUX21X1_HVT U1363 ( .A1(conv2_sum_b[7]), .A2(conv2_sum_a[7]), .S0(n365), .Y(
        tmp_big1[7]) );
  MUX21X1_HVT U1364 ( .A1(conv2_sum_d[7]), .A2(conv2_sum_c[7]), .S0(n361), .Y(
        tmp_big2[7]) );
  MUX21X1_HVT U1365 ( .A1(conv2_sum_b[6]), .A2(conv2_sum_a[6]), .S0(n365), .Y(
        tmp_big1[6]) );
  MUX21X1_HVT U1366 ( .A1(conv2_sum_d[6]), .A2(conv2_sum_c[6]), .S0(n361), .Y(
        tmp_big2[6]) );
  MUX21X1_HVT U1367 ( .A1(conv2_sum_b[4]), .A2(conv2_sum_a[4]), .S0(n362), .Y(
        tmp_big1[4]) );
  MUX21X1_HVT U1368 ( .A1(conv2_sum_d[4]), .A2(conv2_sum_c[4]), .S0(n358), .Y(
        tmp_big2[4]) );
  MUX21X1_HVT U1369 ( .A1(conv2_sum_b[5]), .A2(conv2_sum_a[5]), .S0(n362), .Y(
        tmp_big1[5]) );
  MUX21X1_HVT U1370 ( .A1(conv2_sum_d[5]), .A2(conv2_sum_c[5]), .S0(n361), .Y(
        tmp_big2[5]) );
  MUX21X1_HVT U1371 ( .A1(conv2_sum_b[1]), .A2(conv2_sum_a[1]), .S0(n365), .Y(
        tmp_big1[1]) );
  MUX21X1_HVT U1372 ( .A1(conv2_sum_d[1]), .A2(conv2_sum_c[1]), .S0(n358), .Y(
        tmp_big2[1]) );
  MUX21X1_HVT U1373 ( .A1(conv2_sum_d[0]), .A2(conv2_sum_c[0]), .S0(n358), .Y(
        tmp_big2[0]) );
  MUX21X1_HVT U1374 ( .A1(conv2_sum_b[0]), .A2(conv2_sum_a[0]), .S0(n365), .Y(
        tmp_big1[0]) );
  MUX21X1_HVT U1375 ( .A1(conv2_sum_b[2]), .A2(conv2_sum_a[2]), .S0(n362), .Y(
        tmp_big1[2]) );
  MUX21X1_HVT U1376 ( .A1(conv2_sum_d[2]), .A2(conv2_sum_c[2]), .S0(n359), .Y(
        tmp_big2[2]) );
  MUX21X1_HVT U1377 ( .A1(conv2_sum_b[3]), .A2(conv2_sum_a[3]), .S0(n363), .Y(
        tmp_big1[3]) );
  MUX21X1_HVT U1378 ( .A1(conv2_sum_d[3]), .A2(conv2_sum_c[3]), .S0(n360), .Y(
        tmp_big2[3]) );
  MUX21X1_HVT U1379 ( .A1(conv2_sum_b[29]), .A2(conv2_sum_a[29]), .S0(n364), 
        .Y(tmp_big1[29]) );
  MUX21X1_HVT U1380 ( .A1(conv2_sum_d[29]), .A2(conv2_sum_c[29]), .S0(n358), 
        .Y(tmp_big2[29]) );
  MUX21X1_HVT U1381 ( .A1(conv2_sum_d[31]), .A2(conv2_sum_c[31]), .S0(n360), 
        .Y(tmp_big2[31]) );
  MUX21X1_HVT U1382 ( .A1(conv2_sum_b[28]), .A2(conv2_sum_a[28]), .S0(n365), 
        .Y(tmp_big1[28]) );
  MUX21X1_HVT U1383 ( .A1(conv2_sum_d[28]), .A2(conv2_sum_c[28]), .S0(n361), 
        .Y(tmp_big2[28]) );
  MUX21X1_HVT U1384 ( .A1(conv2_sum_b[24]), .A2(conv2_sum_a[24]), .S0(n365), 
        .Y(tmp_big1[24]) );
  MUX21X1_HVT U1385 ( .A1(conv2_sum_d[25]), .A2(conv2_sum_c[25]), .S0(n358), 
        .Y(tmp_big2[25]) );
  MUX21X1_HVT U1386 ( .A1(conv2_sum_b[30]), .A2(conv2_sum_a[30]), .S0(n364), 
        .Y(tmp_big1[30]) );
  MUX21X1_HVT U1387 ( .A1(conv2_sum_d[30]), .A2(conv2_sum_c[30]), .S0(n361), 
        .Y(tmp_big2[30]) );
  INVX1_HVT U1388 ( .A(tmp_big1[7]), .Y(n685) );
  INVX1_HVT U1389 ( .A(tmp_big1[5]), .Y(n684) );
  INVX1_HVT U1390 ( .A(tmp_big2[1]), .Y(n661) );
  INVX1_HVT U1391 ( .A(tmp_big1[3]), .Y(n682) );
  INVX1_HVT U1392 ( .A(tmp_big1[13]), .Y(n666) );
  INVX1_HVT U1393 ( .A(tmp_big1[15]), .Y(n668) );
  INVX1_HVT U1394 ( .A(tmp_big1[14]), .Y(n667) );
  INVX1_HVT U1395 ( .A(tmp_big1[9]), .Y(n686) );
  INVX1_HVT U1396 ( .A(tmp_big1[11]), .Y(n665) );
  INVX1_HVT U1397 ( .A(tmp_big1[21]), .Y(n672) );
  INVX1_HVT U1398 ( .A(tmp_big1[23]), .Y(n674) );
  INVX1_HVT U1399 ( .A(tmp_big1[17]), .Y(n669) );
  INVX1_HVT U1400 ( .A(tmp_big1[19]), .Y(n671) );
  INVX1_HVT U1401 ( .A(tmp_big1[24]), .Y(n675) );
  INVX1_HVT U1402 ( .A(tmp_big1[29]), .Y(n679) );
  INVX1_HVT U1403 ( .A(tmp_big2[31]), .Y(n662) );
  INVX1_HVT U1404 ( .A(tmp_big1[30]), .Y(n681) );
  INVX1_HVT U1405 ( .A(tmp_big1[25]), .Y(n676) );
  INVX1_HVT U1406 ( .A(tmp_big1[27]), .Y(n678) );
  NAND2X0_HVT U1407 ( .A1(n353), .A2(conv1_sram_rdata_weight[81]), .Y(n433) );
  NAND2X0_HVT U1408 ( .A1(n438), .A2(conv2_sram_rdata_weight[81]), .Y(n434) );
  NAND2X0_HVT U1409 ( .A1(n352), .A2(conv1_sram_rdata_weight[91]), .Y(n435) );
  NAND2X0_HVT U1410 ( .A1(n438), .A2(conv2_sram_rdata_weight[91]), .Y(n436) );
  AO22X1_HVT U1411 ( .A1(conv2_sum_b[30]), .A2(n409), .A3(conv2_sum_a[31]), 
        .A4(n380), .Y(n463) );
  NAND2X0_HVT U1412 ( .A1(conv2_sum_b[29]), .A2(n420), .Y(n455) );
  NAND2X0_HVT U1413 ( .A1(conv2_sum_a[28]), .A2(n455), .Y(n454) );
  NAND2X0_HVT U1414 ( .A1(conv2_sum_b[27]), .A2(n376), .Y(n456) );
  NAND2X0_HVT U1415 ( .A1(conv2_sum_a[26]), .A2(n456), .Y(n457) );
  OA22X1_HVT U1416 ( .A1(conv2_sum_b[27]), .A2(n376), .A3(conv2_sum_b[26]), 
        .A4(n457), .Y(n460) );
  NAND2X0_HVT U1417 ( .A1(conv2_sum_b[25]), .A2(n421), .Y(n524) );
  NAND2X0_HVT U1418 ( .A1(conv2_sum_a[24]), .A2(n524), .Y(n458) );
  OA22X1_HVT U1419 ( .A1(n421), .A2(conv2_sum_b[25]), .A3(n458), .A4(
        conv2_sum_b[24]), .Y(n459) );
  AO22X1_HVT U1420 ( .A1(conv2_sum_b[26]), .A2(n410), .A3(conv2_sum_b[27]), 
        .A4(n376), .Y(n465) );
  NAND2X0_HVT U1421 ( .A1(conv2_sum_a[31]), .A2(n380), .Y(n461) );
  NAND2X0_HVT U1422 ( .A1(conv2_sum_a[30]), .A2(n461), .Y(n462) );
  AO22X1_HVT U1423 ( .A1(conv2_sum_b[22]), .A2(n411), .A3(conv2_sum_b[23]), 
        .A4(n382), .Y(n478) );
  NAND2X0_HVT U1424 ( .A1(conv2_sum_b[21]), .A2(n422), .Y(n467) );
  NAND2X0_HVT U1425 ( .A1(conv2_sum_a[20]), .A2(n467), .Y(n466) );
  OA22X1_HVT U1426 ( .A1(n422), .A2(conv2_sum_b[21]), .A3(n466), .A4(
        conv2_sum_b[20]), .Y(n477) );
  NAND2X0_HVT U1427 ( .A1(conv2_sum_b[19]), .A2(n377), .Y(n468) );
  NAND2X0_HVT U1428 ( .A1(conv2_sum_a[18]), .A2(n468), .Y(n469) );
  OA22X1_HVT U1429 ( .A1(conv2_sum_b[19]), .A2(n377), .A3(conv2_sum_b[18]), 
        .A4(n469), .Y(n472) );
  NAND2X0_HVT U1430 ( .A1(conv2_sum_b[17]), .A2(n423), .Y(n512) );
  NAND2X0_HVT U1431 ( .A1(conv2_sum_a[16]), .A2(n512), .Y(n470) );
  OA22X1_HVT U1432 ( .A1(n423), .A2(conv2_sum_b[17]), .A3(n470), .A4(
        conv2_sum_b[16]), .Y(n471) );
  AO22X1_HVT U1433 ( .A1(conv2_sum_b[18]), .A2(n412), .A3(conv2_sum_b[19]), 
        .A4(n377), .Y(n515) );
  AO22X1_HVT U1434 ( .A1(n472), .A2(n471), .A3(n472), .A4(n515), .Y(n476) );
  NAND2X0_HVT U1435 ( .A1(conv2_sum_b[23]), .A2(n382), .Y(n473) );
  NAND2X0_HVT U1436 ( .A1(conv2_sum_a[22]), .A2(n473), .Y(n474) );
  OA22X1_HVT U1437 ( .A1(n382), .A2(conv2_sum_b[23]), .A3(n474), .A4(
        conv2_sum_b[22]), .Y(n475) );
  AO22X1_HVT U1438 ( .A1(conv2_sum_b[14]), .A2(n413), .A3(conv2_sum_b[15]), 
        .A4(n372), .Y(n491) );
  NAND2X0_HVT U1439 ( .A1(conv2_sum_b[13]), .A2(n399), .Y(n480) );
  NAND2X0_HVT U1440 ( .A1(conv2_sum_a[12]), .A2(n480), .Y(n479) );
  OA22X1_HVT U1441 ( .A1(n399), .A2(conv2_sum_b[13]), .A3(n479), .A4(
        conv2_sum_b[12]), .Y(n490) );
  NAND2X0_HVT U1442 ( .A1(conv2_sum_b[11]), .A2(n368), .Y(n481) );
  NAND2X0_HVT U1443 ( .A1(conv2_sum_a[10]), .A2(n481), .Y(n482) );
  OA22X1_HVT U1444 ( .A1(conv2_sum_b[11]), .A2(n368), .A3(conv2_sum_b[10]), 
        .A4(n482), .Y(n485) );
  NAND2X0_HVT U1445 ( .A1(conv2_sum_b[9]), .A2(n400), .Y(n492) );
  NAND2X0_HVT U1446 ( .A1(conv2_sum_a[8]), .A2(n492), .Y(n483) );
  OA22X1_HVT U1447 ( .A1(n400), .A2(conv2_sum_b[9]), .A3(n483), .A4(
        conv2_sum_b[8]), .Y(n484) );
  AO22X1_HVT U1448 ( .A1(conv2_sum_b[10]), .A2(n390), .A3(conv2_sum_b[11]), 
        .A4(n368), .Y(n495) );
  AO22X1_HVT U1449 ( .A1(n485), .A2(n484), .A3(n485), .A4(n495), .Y(n489) );
  NAND2X0_HVT U1450 ( .A1(conv2_sum_b[15]), .A2(n372), .Y(n486) );
  NAND2X0_HVT U1451 ( .A1(conv2_sum_a[14]), .A2(n486), .Y(n487) );
  OA22X1_HVT U1452 ( .A1(n372), .A2(conv2_sum_b[15]), .A3(n487), .A4(
        conv2_sum_b[14]), .Y(n488) );
  OAI21X1_HVT U1453 ( .A1(conv2_sum_a[8]), .A2(n386), .A3(n492), .Y(n493) );
  OR3X1_HVT U1454 ( .A1(n495), .A2(n494), .A3(n493), .Y(n518) );
  NAND2X0_HVT U1455 ( .A1(conv2_sum_b[3]), .A2(n369), .Y(n496) );
  NAND2X0_HVT U1456 ( .A1(conv2_sum_a[2]), .A2(n496), .Y(n497) );
  OA22X1_HVT U1457 ( .A1(conv2_sum_b[3]), .A2(n369), .A3(conv2_sum_b[2]), .A4(
        n497), .Y(n503) );
  AO22X1_HVT U1458 ( .A1(conv2_sum_b[2]), .A2(n391), .A3(conv2_sum_b[3]), .A4(
        n369), .Y(n502) );
  NAND2X0_HVT U1459 ( .A1(n384), .A2(conv2_sum_a[1]), .Y(n498) );
  NAND2X0_HVT U1460 ( .A1(conv2_sum_b[0]), .A2(n498), .Y(n499) );
  OAI22X1_HVT U1461 ( .A1(conv2_sum_a[0]), .A2(n499), .A3(n384), .A4(
        conv2_sum_a[1]), .Y(n501) );
  AO22X1_HVT U1462 ( .A1(conv2_sum_b[5]), .A2(n366), .A3(conv2_sum_b[4]), .A4(
        n388), .Y(n5001) );
  AO221X1_HVT U1463 ( .A1(n503), .A2(n502), .A3(n503), .A4(n501), .A5(n5001), 
        .Y(n511) );
  AO22X1_HVT U1464 ( .A1(conv2_sum_b[6]), .A2(n392), .A3(conv2_sum_b[7]), .A4(
        n373), .Y(n510) );
  NAND2X0_HVT U1465 ( .A1(conv2_sum_b[5]), .A2(n366), .Y(n504) );
  NAND2X0_HVT U1466 ( .A1(conv2_sum_a[4]), .A2(n504), .Y(n505) );
  OA22X1_HVT U1467 ( .A1(n505), .A2(conv2_sum_b[4]), .A3(n366), .A4(
        conv2_sum_b[5]), .Y(n509) );
  NAND2X0_HVT U1468 ( .A1(conv2_sum_b[7]), .A2(n373), .Y(n506) );
  NAND2X0_HVT U1469 ( .A1(conv2_sum_a[6]), .A2(n506), .Y(n507) );
  OA22X1_HVT U1470 ( .A1(n373), .A2(conv2_sum_b[7]), .A3(n507), .A4(
        conv2_sum_b[6]), .Y(n508) );
  OA221X1_HVT U1471 ( .A1(n511), .A2(n510), .A3(n509), .A4(n510), .A5(n508), 
        .Y(n517) );
  OAI21X1_HVT U1472 ( .A1(conv2_sum_a[16]), .A2(n397), .A3(n512), .Y(n513) );
  OR3X1_HVT U1473 ( .A1(n515), .A2(n514), .A3(n513), .Y(n516) );
  AO221X1_HVT U1474 ( .A1(n519), .A2(n518), .A3(n519), .A4(n517), .A5(n516), 
        .Y(n520) );
  NAND2X0_HVT U1475 ( .A1(n521), .A2(n520), .Y(n522) );
  OA221X1_HVT U1476 ( .A1(n476), .A2(n514), .A3(n477), .A4(n478), .A5(n475), 
        .Y(n521) );
  OA221X1_HVT U1477 ( .A1(n489), .A2(n494), .A3(n490), .A4(n491), .A5(n488), 
        .Y(n519) );
  AO22X1_HVT U1478 ( .A1(conv2_sum_d[30]), .A2(n414), .A3(conv2_sum_c[31]), 
        .A4(n381), .Y(n537) );
  NAND2X0_HVT U1479 ( .A1(conv2_sum_d[29]), .A2(n424), .Y(n526) );
  NAND2X0_HVT U1480 ( .A1(conv2_sum_c[28]), .A2(n526), .Y(n525) );
  OA22X1_HVT U1481 ( .A1(n424), .A2(conv2_sum_d[29]), .A3(n525), .A4(
        conv2_sum_d[28]), .Y(n536) );
  NAND2X0_HVT U1482 ( .A1(conv2_sum_d[27]), .A2(n378), .Y(n527) );
  NAND2X0_HVT U1483 ( .A1(conv2_sum_c[26]), .A2(n527), .Y(n528) );
  OA22X1_HVT U1484 ( .A1(conv2_sum_d[27]), .A2(n378), .A3(conv2_sum_d[26]), 
        .A4(n528), .Y(n531) );
  NAND2X0_HVT U1485 ( .A1(conv2_sum_d[25]), .A2(n425), .Y(n591) );
  NAND2X0_HVT U1486 ( .A1(conv2_sum_c[24]), .A2(n591), .Y(n529) );
  OA22X1_HVT U1487 ( .A1(n425), .A2(conv2_sum_d[25]), .A3(n529), .A4(
        conv2_sum_d[24]), .Y(n530) );
  AO22X1_HVT U1488 ( .A1(conv2_sum_d[26]), .A2(n396), .A3(conv2_sum_d[27]), 
        .A4(n378), .Y(n539) );
  AO22X1_HVT U1489 ( .A1(n531), .A2(n530), .A3(n531), .A4(n539), .Y(n535) );
  NAND2X0_HVT U1490 ( .A1(conv2_sum_c[31]), .A2(n381), .Y(n532) );
  NAND2X0_HVT U1491 ( .A1(conv2_sum_c[30]), .A2(n532), .Y(n533) );
  OA22X1_HVT U1492 ( .A1(n381), .A2(conv2_sum_c[31]), .A3(n533), .A4(
        conv2_sum_d[30]), .Y(n534) );
  NAND2X0_HVT U1493 ( .A1(conv2_sum_d[24]), .A2(n408), .Y(n592) );
  AO22X1_HVT U1494 ( .A1(conv2_sum_d[22]), .A2(n415), .A3(conv2_sum_d[23]), 
        .A4(n383), .Y(n549) );
  NAND2X0_HVT U1495 ( .A1(conv2_sum_d[21]), .A2(n426), .Y(n541) );
  NAND2X0_HVT U1496 ( .A1(conv2_sum_c[20]), .A2(n541), .Y(n540) );
  NAND2X0_HVT U1497 ( .A1(conv2_sum_d[19]), .A2(n379), .Y(n542) );
  NAND2X0_HVT U1498 ( .A1(conv2_sum_c[18]), .A2(n542), .Y(n543) );
  OA22X1_HVT U1499 ( .A1(conv2_sum_d[19]), .A2(n379), .A3(conv2_sum_d[18]), 
        .A4(n543), .Y(n546) );
  NAND2X0_HVT U1500 ( .A1(conv2_sum_d[17]), .A2(n427), .Y(n583) );
  NAND2X0_HVT U1501 ( .A1(conv2_sum_c[16]), .A2(n583), .Y(n544) );
  OA22X1_HVT U1502 ( .A1(n427), .A2(conv2_sum_d[17]), .A3(n544), .A4(
        conv2_sum_d[16]), .Y(n545) );
  AO22X1_HVT U1503 ( .A1(conv2_sum_d[18]), .A2(n416), .A3(conv2_sum_d[19]), 
        .A4(n379), .Y(n586) );
  NAND2X0_HVT U1504 ( .A1(conv2_sum_d[23]), .A2(n383), .Y(n547) );
  NAND2X0_HVT U1505 ( .A1(conv2_sum_c[22]), .A2(n547), .Y(n548) );
  AO22X1_HVT U1506 ( .A1(conv2_sum_d[14]), .A2(n417), .A3(conv2_sum_d[15]), 
        .A4(n374), .Y(n562) );
  NAND2X0_HVT U1507 ( .A1(conv2_sum_d[13]), .A2(n401), .Y(n551) );
  NAND2X0_HVT U1508 ( .A1(conv2_sum_c[12]), .A2(n551), .Y(n550) );
  OA22X1_HVT U1509 ( .A1(n401), .A2(conv2_sum_d[13]), .A3(n550), .A4(
        conv2_sum_d[12]), .Y(n561) );
  NAND2X0_HVT U1510 ( .A1(conv2_sum_d[11]), .A2(n370), .Y(n552) );
  NAND2X0_HVT U1511 ( .A1(conv2_sum_c[10]), .A2(n552), .Y(n553) );
  OA22X1_HVT U1512 ( .A1(conv2_sum_d[11]), .A2(n370), .A3(conv2_sum_d[10]), 
        .A4(n553), .Y(n556) );
  NAND2X0_HVT U1513 ( .A1(conv2_sum_d[9]), .A2(n402), .Y(n563) );
  NAND2X0_HVT U1514 ( .A1(conv2_sum_c[8]), .A2(n563), .Y(n554) );
  OA22X1_HVT U1515 ( .A1(n402), .A2(conv2_sum_d[9]), .A3(n554), .A4(
        conv2_sum_d[8]), .Y(n555) );
  AO22X1_HVT U1516 ( .A1(conv2_sum_d[10]), .A2(n393), .A3(conv2_sum_d[11]), 
        .A4(n370), .Y(n566) );
  AO22X1_HVT U1517 ( .A1(n556), .A2(n555), .A3(n556), .A4(n566), .Y(n560) );
  NAND2X0_HVT U1518 ( .A1(conv2_sum_d[15]), .A2(n374), .Y(n557) );
  NAND2X0_HVT U1519 ( .A1(conv2_sum_c[14]), .A2(n557), .Y(n558) );
  OA22X1_HVT U1520 ( .A1(n374), .A2(conv2_sum_d[15]), .A3(n558), .A4(
        conv2_sum_d[14]), .Y(n559) );
  OAI21X1_HVT U1521 ( .A1(conv2_sum_c[8]), .A2(n387), .A3(n563), .Y(n564) );
  NAND2X0_HVT U1522 ( .A1(conv2_sum_d[3]), .A2(n371), .Y(n567) );
  NAND2X0_HVT U1523 ( .A1(conv2_sum_c[2]), .A2(n567), .Y(n568) );
  OA22X1_HVT U1524 ( .A1(conv2_sum_d[3]), .A2(n371), .A3(conv2_sum_d[2]), .A4(
        n568), .Y(n574) );
  AO22X1_HVT U1525 ( .A1(conv2_sum_d[2]), .A2(n394), .A3(conv2_sum_d[3]), .A4(
        n371), .Y(n573) );
  NAND2X0_HVT U1526 ( .A1(n385), .A2(conv2_sum_c[1]), .Y(n569) );
  NAND2X0_HVT U1527 ( .A1(conv2_sum_d[0]), .A2(n569), .Y(n570) );
  OAI22X1_HVT U1528 ( .A1(conv2_sum_c[0]), .A2(n570), .A3(n385), .A4(
        conv2_sum_c[1]), .Y(n572) );
  AO22X1_HVT U1529 ( .A1(conv2_sum_d[5]), .A2(n367), .A3(conv2_sum_d[4]), .A4(
        n389), .Y(n571) );
  AO221X1_HVT U1530 ( .A1(n574), .A2(n573), .A3(n574), .A4(n572), .A5(n571), 
        .Y(n582) );
  AO22X1_HVT U1531 ( .A1(conv2_sum_d[6]), .A2(n395), .A3(conv2_sum_d[7]), .A4(
        n375), .Y(n581) );
  NAND2X0_HVT U1532 ( .A1(conv2_sum_d[5]), .A2(n367), .Y(n575) );
  NAND2X0_HVT U1533 ( .A1(conv2_sum_c[4]), .A2(n575), .Y(n576) );
  OA22X1_HVT U1534 ( .A1(n576), .A2(conv2_sum_d[4]), .A3(n367), .A4(
        conv2_sum_d[5]), .Y(n580) );
  NAND2X0_HVT U1535 ( .A1(conv2_sum_d[7]), .A2(n375), .Y(n577) );
  NAND2X0_HVT U1536 ( .A1(conv2_sum_c[6]), .A2(n577), .Y(n578) );
  OA22X1_HVT U1537 ( .A1(n375), .A2(conv2_sum_d[7]), .A3(n578), .A4(
        conv2_sum_d[6]), .Y(n579) );
  OA221X1_HVT U1538 ( .A1(n582), .A2(n581), .A3(n580), .A4(n581), .A5(n579), 
        .Y(n587) );
  OAI21X1_HVT U1539 ( .A1(conv2_sum_c[16]), .A2(n398), .A3(n583), .Y(n584) );
  NAND4X0_HVT U1540 ( .A1(n592), .A2(n591), .A3(n590), .A4(n589), .Y(n593) );
  OA221X1_HVT U1541 ( .A1(n535), .A2(n538), .A3(n536), .A4(n537), .A5(n534), 
        .Y(n594) );
  OA221X1_HVT U1542 ( .A1(n560), .A2(n565), .A3(n561), .A4(n562), .A5(n559), 
        .Y(n588) );
  AO22X1_HVT U1543 ( .A1(tmp_big2[30]), .A2(n681), .A3(tmp_big1[31]), .A4(n662), .Y(n607) );
  NAND2X0_HVT U1544 ( .A1(tmp_big2[29]), .A2(n679), .Y(n596) );
  NAND2X0_HVT U1545 ( .A1(tmp_big1[28]), .A2(n596), .Y(n595) );
  OA22X1_HVT U1546 ( .A1(n679), .A2(tmp_big2[29]), .A3(n595), .A4(tmp_big2[28]), .Y(n606) );
  NAND2X0_HVT U1547 ( .A1(tmp_big2[27]), .A2(n678), .Y(n597) );
  NAND2X0_HVT U1548 ( .A1(tmp_big1[26]), .A2(n597), .Y(n598) );
  OA22X1_HVT U1549 ( .A1(tmp_big2[27]), .A2(n678), .A3(tmp_big2[26]), .A4(n598), .Y(n601) );
  NAND2X0_HVT U1550 ( .A1(tmp_big2[25]), .A2(n676), .Y(n656) );
  NAND2X0_HVT U1551 ( .A1(tmp_big1[24]), .A2(n656), .Y(n599) );
  OA22X1_HVT U1552 ( .A1(n676), .A2(tmp_big2[25]), .A3(n599), .A4(tmp_big2[24]), .Y(n600) );
  AO22X1_HVT U1553 ( .A1(tmp_big2[26]), .A2(n677), .A3(tmp_big2[27]), .A4(n678), .Y(n609) );
  AO22X1_HVT U1554 ( .A1(n601), .A2(n600), .A3(n601), .A4(n609), .Y(n605) );
  NAND2X0_HVT U1555 ( .A1(tmp_big1[31]), .A2(n662), .Y(n602) );
  NAND2X0_HVT U1556 ( .A1(tmp_big1[30]), .A2(n602), .Y(n603) );
  OA22X1_HVT U1557 ( .A1(n662), .A2(tmp_big1[31]), .A3(n603), .A4(tmp_big2[30]), .Y(n604) );
  NAND2X0_HVT U1558 ( .A1(tmp_big2[24]), .A2(n675), .Y(n657) );
  AO22X1_HVT U1559 ( .A1(tmp_big2[22]), .A2(n673), .A3(tmp_big2[23]), .A4(n674), .Y(n619) );
  NAND2X0_HVT U1560 ( .A1(tmp_big2[21]), .A2(n672), .Y(n611) );
  NAND2X0_HVT U1561 ( .A1(tmp_big1[20]), .A2(n611), .Y(n610) );
  NAND2X0_HVT U1562 ( .A1(tmp_big2[19]), .A2(n671), .Y(n612) );
  NAND2X0_HVT U1563 ( .A1(tmp_big1[18]), .A2(n612), .Y(n613) );
  OA22X1_HVT U1564 ( .A1(tmp_big2[19]), .A2(n671), .A3(tmp_big2[18]), .A4(n613), .Y(n616) );
  NAND2X0_HVT U1565 ( .A1(tmp_big2[17]), .A2(n669), .Y(n647) );
  NAND2X0_HVT U1566 ( .A1(tmp_big1[16]), .A2(n647), .Y(n614) );
  OA22X1_HVT U1567 ( .A1(n669), .A2(tmp_big2[17]), .A3(n614), .A4(tmp_big2[16]), .Y(n615) );
  AO22X1_HVT U1568 ( .A1(tmp_big2[18]), .A2(n670), .A3(tmp_big2[19]), .A4(n671), .Y(n650) );
  NAND2X0_HVT U1569 ( .A1(tmp_big2[23]), .A2(n674), .Y(n617) );
  NAND2X0_HVT U1570 ( .A1(tmp_big1[22]), .A2(n617), .Y(n618) );
  AO22X1_HVT U1571 ( .A1(tmp_big2[14]), .A2(n667), .A3(tmp_big2[15]), .A4(n668), .Y(n632) );
  NAND2X0_HVT U1572 ( .A1(tmp_big2[13]), .A2(n666), .Y(n621) );
  NAND2X0_HVT U1573 ( .A1(tmp_big1[12]), .A2(n621), .Y(n620) );
  OA22X1_HVT U1574 ( .A1(n666), .A2(tmp_big2[13]), .A3(n620), .A4(tmp_big2[12]), .Y(n631) );
  NAND2X0_HVT U1575 ( .A1(tmp_big2[11]), .A2(n665), .Y(n622) );
  NAND2X0_HVT U1576 ( .A1(tmp_big1[10]), .A2(n622), .Y(n623) );
  OA22X1_HVT U1577 ( .A1(tmp_big2[11]), .A2(n665), .A3(tmp_big2[10]), .A4(n623), .Y(n626) );
  NAND2X0_HVT U1578 ( .A1(tmp_big2[9]), .A2(n686), .Y(n633) );
  NAND2X0_HVT U1579 ( .A1(tmp_big1[8]), .A2(n633), .Y(n624) );
  OA22X1_HVT U1580 ( .A1(n686), .A2(tmp_big2[9]), .A3(n624), .A4(tmp_big2[8]), 
        .Y(n625) );
  AO22X1_HVT U1581 ( .A1(tmp_big2[10]), .A2(n664), .A3(tmp_big2[11]), .A4(n665), .Y(n636) );
  AO22X1_HVT U1582 ( .A1(n626), .A2(n625), .A3(n626), .A4(n636), .Y(n630) );
  NAND2X0_HVT U1583 ( .A1(tmp_big2[15]), .A2(n668), .Y(n627) );
  NAND2X0_HVT U1584 ( .A1(tmp_big1[14]), .A2(n627), .Y(n628) );
  OA22X1_HVT U1585 ( .A1(n668), .A2(tmp_big2[15]), .A3(n628), .A4(tmp_big2[14]), .Y(n629) );
  OAI21X1_HVT U1586 ( .A1(tmp_big1[8]), .A2(n663), .A3(n633), .Y(n634) );
  OR3X1_HVT U1587 ( .A1(n636), .A2(n635), .A3(n634), .Y(n652) );
  NAND2X0_HVT U1588 ( .A1(tmp_big2[3]), .A2(n682), .Y(n637) );
  NAND2X0_HVT U1589 ( .A1(tmp_big1[2]), .A2(n637), .Y(n638) );
  OA22X1_HVT U1590 ( .A1(tmp_big2[3]), .A2(n682), .A3(tmp_big2[2]), .A4(n638), 
        .Y(n644) );
  AO22X1_HVT U1591 ( .A1(tmp_big2[2]), .A2(n680), .A3(tmp_big2[3]), .A4(n682), 
        .Y(n643) );
  NAND2X0_HVT U1592 ( .A1(n661), .A2(tmp_big1[1]), .Y(n639) );
  NAND2X0_HVT U1593 ( .A1(tmp_big2[0]), .A2(n639), .Y(n640) );
  OAI22X1_HVT U1594 ( .A1(tmp_big1[0]), .A2(n640), .A3(n661), .A4(tmp_big1[1]), 
        .Y(n642) );
  AO22X1_HVT U1595 ( .A1(tmp_big2[5]), .A2(n684), .A3(tmp_big2[4]), .A4(n683), 
        .Y(n641) );
  NAND2X0_HVT U1596 ( .A1(tmp_big2[5]), .A2(n684), .Y(n645) );
  NAND2X0_HVT U1597 ( .A1(tmp_big2[7]), .A2(n685), .Y(n646) );
  OAI21X1_HVT U1598 ( .A1(tmp_big1[16]), .A2(n660), .A3(n647), .Y(n648) );
  NAND4X0_HVT U1599 ( .A1(n657), .A2(n656), .A3(n655), .A4(n654), .Y(n658) );
  OA221X1_HVT U1600 ( .A1(n605), .A2(n608), .A3(n606), .A4(n607), .A5(n604), 
        .Y(n659) );
  OA221X1_HVT U1601 ( .A1(n630), .A2(n635), .A3(n631), .A4(n632), .A5(n629), 
        .Y(n653) );
  MUX21X1_HVT U1602 ( .A1(conv2_sram_rdata_weight[97]), .A2(
        conv1_sram_rdata_weight[97]), .S0(n353), .Y(conv_weight_box[91]) );
  MUX21X1_HVT U1603 ( .A1(conv2_sram_rdata_weight[90]), .A2(
        conv1_sram_rdata_weight[90]), .S0(n348), .Y(conv_weight_box[86]) );
  MUX21X1_HVT U1604 ( .A1(conv2_sram_rdata_weight[85]), .A2(
        conv1_sram_rdata_weight[85]), .S0(n432), .Y(conv_weight_box[81]) );
  MUX21X1_HVT U1605 ( .A1(conv2_sram_rdata_weight[77]), .A2(
        conv1_sram_rdata_weight[77]), .S0(n432), .Y(conv_weight_box[73]) );
  MUX21X1_HVT U1606 ( .A1(conv2_sram_rdata_weight[69]), .A2(
        conv1_sram_rdata_weight[69]), .S0(n353), .Y(conv_weight_box[65]) );
  MUX21X1_HVT U1607 ( .A1(conv2_sram_rdata_weight[65]), .A2(
        conv1_sram_rdata_weight[65]), .S0(n336), .Y(conv_weight_box[61]) );
  MUX21X1_HVT U1608 ( .A1(conv2_sram_rdata_weight[60]), .A2(
        conv1_sram_rdata_weight[60]), .S0(n348), .Y(conv_weight_box[56]) );
  MUX21X1_HVT U1609 ( .A1(conv2_sram_rdata_weight[50]), .A2(
        conv1_sram_rdata_weight[50]), .S0(n332), .Y(conv_weight_box[46]) );
  MUX21X1_HVT U1610 ( .A1(conv2_sram_rdata_weight[38]), .A2(
        conv1_sram_rdata_weight[38]), .S0(n351), .Y(conv_weight_box[35]) );
  MUX21X1_HVT U1611 ( .A1(conv2_sram_rdata_weight[37]), .A2(
        conv1_sram_rdata_weight[37]), .S0(n350), .Y(conv_weight_box[34]) );
  MUX21X1_HVT U1612 ( .A1(conv2_sram_rdata_weight[34]), .A2(
        conv1_sram_rdata_weight[34]), .S0(n335), .Y(conv_weight_box[31]) );
  MUX21X1_HVT U1613 ( .A1(conv2_sram_rdata_weight[29]), .A2(
        conv1_sram_rdata_weight[29]), .S0(n334), .Y(conv_weight_box[27]) );
  MUX21X1_HVT U1614 ( .A1(conv2_sram_rdata_weight[21]), .A2(
        conv1_sram_rdata_weight[21]), .S0(n333), .Y(conv_weight_box[19]) );
  MUX21X1_HVT U1615 ( .A1(conv2_sram_rdata_weight[18]), .A2(
        conv1_sram_rdata_weight[18]), .S0(n334), .Y(conv_weight_box[16]) );
  MUX21X1_HVT U1616 ( .A1(conv2_sram_rdata_weight[17]), .A2(
        conv1_sram_rdata_weight[17]), .S0(n432), .Y(conv_weight_box[15]) );
  MUX21X1_HVT U1617 ( .A1(conv2_sram_rdata_weight[16]), .A2(
        conv1_sram_rdata_weight[16]), .S0(n332), .Y(conv_weight_box[14]) );
  MUX21X1_HVT U1618 ( .A1(conv2_sum_b[27]), .A2(conv2_sum_a[27]), .S0(n363), 
        .Y(tmp_big1[27]) );
  MUX21X1_HVT U1619 ( .A1(conv2_sum_b[26]), .A2(conv2_sum_a[26]), .S0(n363), 
        .Y(tmp_big1[26]) );
  MUX21X1_HVT U1620 ( .A1(conv2_sum_b[25]), .A2(conv2_sum_a[25]), .S0(n365), 
        .Y(tmp_big1[25]) );
  MUX21X1_HVT U1621 ( .A1(conv2_sum_b[23]), .A2(conv2_sum_a[23]), .S0(n364), 
        .Y(tmp_big1[23]) );
  MUX21X1_HVT U1622 ( .A1(conv2_sum_b[22]), .A2(conv2_sum_a[22]), .S0(n362), 
        .Y(tmp_big1[22]) );
  MUX21X1_HVT U1623 ( .A1(conv2_sum_b[21]), .A2(conv2_sum_a[21]), .S0(n364), 
        .Y(tmp_big1[21]) );
  MUX21X1_HVT U1624 ( .A1(conv2_sum_b[20]), .A2(conv2_sum_a[20]), .S0(n362), 
        .Y(tmp_big1[20]) );
  MUX21X1_HVT U1625 ( .A1(conv2_sum_b[19]), .A2(conv2_sum_a[19]), .S0(n364), 
        .Y(tmp_big1[19]) );
  MUX21X1_HVT U1626 ( .A1(conv2_sum_b[18]), .A2(conv2_sum_a[18]), .S0(n363), 
        .Y(tmp_big1[18]) );
  MUX21X1_HVT U1627 ( .A1(conv2_sum_b[17]), .A2(conv2_sum_a[17]), .S0(n363), 
        .Y(tmp_big1[17]) );
  MUX21X1_HVT U1628 ( .A1(conv2_sum_b[16]), .A2(conv2_sum_a[16]), .S0(n362), 
        .Y(tmp_big1[16]) );
  MUX21X1_HVT U1629 ( .A1(conv2_sum_b[15]), .A2(conv2_sum_a[15]), .S0(n364), 
        .Y(tmp_big1[15]) );
  MUX21X1_HVT U1630 ( .A1(conv2_sum_b[14]), .A2(conv2_sum_a[14]), .S0(n365), 
        .Y(tmp_big1[14]) );
  MUX21X1_HVT U1631 ( .A1(conv2_sum_b[13]), .A2(conv2_sum_a[13]), .S0(n363), 
        .Y(tmp_big1[13]) );
  MUX21X1_HVT U1632 ( .A1(conv2_sum_b[12]), .A2(conv2_sum_a[12]), .S0(n363), 
        .Y(tmp_big1[12]) );
  MUX21X1_HVT U1633 ( .A1(conv2_sum_b[11]), .A2(conv2_sum_a[11]), .S0(n364), 
        .Y(tmp_big1[11]) );
  MUX21X1_HVT U1634 ( .A1(conv2_sum_b[10]), .A2(conv2_sum_a[10]), .S0(n364), 
        .Y(tmp_big1[10]) );
  MUX21X1_HVT U1635 ( .A1(conv2_sum_b[9]), .A2(conv2_sum_a[9]), .S0(n362), .Y(
        tmp_big1[9]) );
  MUX21X1_HVT U1636 ( .A1(conv2_sum_b[8]), .A2(conv2_sum_a[8]), .S0(n363), .Y(
        tmp_big1[8]) );
  MUX21X1_HVT U1637 ( .A1(conv2_sum_d[27]), .A2(conv2_sum_c[27]), .S0(n359), 
        .Y(tmp_big2[27]) );
  MUX21X1_HVT U1638 ( .A1(conv2_sum_d[26]), .A2(conv2_sum_c[26]), .S0(n359), 
        .Y(tmp_big2[26]) );
  MUX21X1_HVT U1639 ( .A1(conv2_sum_d[24]), .A2(conv2_sum_c[24]), .S0(n360), 
        .Y(tmp_big2[24]) );
  MUX21X1_HVT U1640 ( .A1(conv2_sum_d[23]), .A2(conv2_sum_c[23]), .S0(n360), 
        .Y(tmp_big2[23]) );
  MUX21X1_HVT U1641 ( .A1(conv2_sum_d[22]), .A2(conv2_sum_c[22]), .S0(n358), 
        .Y(tmp_big2[22]) );
  MUX21X1_HVT U1642 ( .A1(conv2_sum_d[21]), .A2(conv2_sum_c[21]), .S0(n358), 
        .Y(tmp_big2[21]) );
  MUX21X1_HVT U1643 ( .A1(conv2_sum_d[20]), .A2(conv2_sum_c[20]), .S0(n361), 
        .Y(tmp_big2[20]) );
  MUX21X1_HVT U1644 ( .A1(conv2_sum_d[19]), .A2(conv2_sum_c[19]), .S0(n360), 
        .Y(tmp_big2[19]) );
  MUX21X1_HVT U1645 ( .A1(conv2_sum_d[18]), .A2(conv2_sum_c[18]), .S0(n360), 
        .Y(tmp_big2[18]) );
  MUX21X1_HVT U1646 ( .A1(conv2_sum_d[17]), .A2(conv2_sum_c[17]), .S0(n359), 
        .Y(tmp_big2[17]) );
  MUX21X1_HVT U1647 ( .A1(conv2_sum_d[16]), .A2(conv2_sum_c[16]), .S0(n359), 
        .Y(tmp_big2[16]) );
  MUX21X1_HVT U1648 ( .A1(conv2_sum_d[15]), .A2(conv2_sum_c[15]), .S0(n358), 
        .Y(tmp_big2[15]) );
  MUX21X1_HVT U1649 ( .A1(conv2_sum_d[14]), .A2(conv2_sum_c[14]), .S0(n360), 
        .Y(tmp_big2[14]) );
  MUX21X1_HVT U1650 ( .A1(conv2_sum_d[13]), .A2(conv2_sum_c[13]), .S0(n359), 
        .Y(tmp_big2[13]) );
  MUX21X1_HVT U1651 ( .A1(conv2_sum_d[12]), .A2(conv2_sum_c[12]), .S0(n359), 
        .Y(tmp_big2[12]) );
  MUX21X1_HVT U1652 ( .A1(conv2_sum_d[11]), .A2(conv2_sum_c[11]), .S0(n361), 
        .Y(tmp_big2[11]) );
  MUX21X1_HVT U1653 ( .A1(conv2_sum_d[10]), .A2(conv2_sum_c[10]), .S0(n361), 
        .Y(tmp_big2[10]) );
  MUX21X1_HVT U1654 ( .A1(conv2_sum_d[9]), .A2(conv2_sum_c[9]), .S0(n359), .Y(
        tmp_big2[9]) );
  MUX21X1_HVT U1655 ( .A1(conv2_sum_d[8]), .A2(conv2_sum_c[8]), .S0(n360), .Y(
        tmp_big2[8]) );
  MUX21X1_HVT U1656 ( .A1(tmp_big2[0]), .A2(tmp_big1[0]), .S0(n357), .Y(
        data_out[0]) );
  MUX21X1_HVT U1657 ( .A1(tmp_big2[1]), .A2(tmp_big1[1]), .S0(n356), .Y(
        data_out[1]) );
  MUX21X1_HVT U1658 ( .A1(tmp_big2[2]), .A2(tmp_big1[2]), .S0(n355), .Y(
        data_out[2]) );
  MUX21X1_HVT U1659 ( .A1(tmp_big2[3]), .A2(tmp_big1[3]), .S0(n357), .Y(
        data_out[3]) );
  MUX21X1_HVT U1660 ( .A1(tmp_big2[4]), .A2(tmp_big1[4]), .S0(n354), .Y(
        data_out[4]) );
  MUX21X1_HVT U1661 ( .A1(tmp_big2[14]), .A2(tmp_big1[14]), .S0(n357), .Y(
        data_out[14]) );
  MUX21X1_HVT U1662 ( .A1(tmp_big2[15]), .A2(tmp_big1[15]), .S0(n355), .Y(
        data_out[15]) );
  MUX21X1_HVT U1663 ( .A1(tmp_big2[16]), .A2(tmp_big1[16]), .S0(n354), .Y(
        data_out[16]) );
  MUX21X1_HVT U1664 ( .A1(tmp_big2[17]), .A2(tmp_big1[17]), .S0(n357), .Y(
        data_out[17]) );
endmodule


module quantize ( clk, srstn, bias_data, mode, quantized_data, ori_data_31_, 
        ori_data_30_, ori_data_29_, ori_data_28_, ori_data_27_, ori_data_26_, 
        ori_data_25_, ori_data_24_, ori_data_23_, ori_data_22_, ori_data_21_, 
        ori_data_20_, ori_data_19_, ori_data_18_, ori_data_17_, ori_data_16_, 
        ori_data_15_, ori_data_14_, ori_data_13_, ori_data_12_, ori_data_11_, 
        ori_data_10_, ori_data_9_, ori_data_8_, ori_data_7_, ori_data_6_, 
        ori_data_5_ );
  input [3:0] bias_data;
  input [1:0] mode;
  output [7:0] quantized_data;
  input clk, srstn, ori_data_31_, ori_data_30_, ori_data_29_, ori_data_28_,
         ori_data_27_, ori_data_26_, ori_data_25_, ori_data_24_, ori_data_23_,
         ori_data_22_, ori_data_21_, ori_data_20_, ori_data_19_, ori_data_18_,
         ori_data_17_, ori_data_16_, ori_data_15_, ori_data_14_, ori_data_13_,
         ori_data_12_, ori_data_11_, ori_data_10_, ori_data_9_, ori_data_8_,
         ori_data_7_, ori_data_6_, ori_data_5_;
  wire   N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N59, N60, N61, N113, N114, N115, N116, N117, N118, N119,
         N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130,
         N131, n13, DP_OP_26J5_124_4249_n311, DP_OP_26J5_124_4249_n310,
         DP_OP_26J5_124_4249_n309, DP_OP_26J5_124_4249_n308,
         DP_OP_26J5_124_4249_n306, DP_OP_26J5_124_4249_n304,
         DP_OP_26J5_124_4249_n299, DP_OP_26J5_124_4249_n298,
         DP_OP_26J5_124_4249_n297, DP_OP_26J5_124_4249_n296,
         DP_OP_26J5_124_4249_n295, DP_OP_26J5_124_4249_n294,
         DP_OP_26J5_124_4249_n293, DP_OP_26J5_124_4249_n287,
         DP_OP_26J5_124_4249_n286, DP_OP_26J5_124_4249_n285,
         DP_OP_26J5_124_4249_n284, DP_OP_26J5_124_4249_n283,
         DP_OP_26J5_124_4249_n282, DP_OP_26J5_124_4249_n281,
         DP_OP_26J5_124_4249_n280, DP_OP_26J5_124_4249_n275,
         DP_OP_26J5_124_4249_n272, DP_OP_26J5_124_4249_n271,
         DP_OP_26J5_124_4249_n270, DP_OP_26J5_124_4249_n269,
         DP_OP_26J5_124_4249_n264, DP_OP_26J5_124_4249_n263,
         DP_OP_26J5_124_4249_n262, DP_OP_26J5_124_4249_n252,
         DP_OP_26J5_124_4249_n246, DP_OP_26J5_124_4249_n245,
         DP_OP_26J5_124_4249_n244, DP_OP_26J5_124_4249_n243,
         DP_OP_26J5_124_4249_n234, DP_OP_26J5_124_4249_n233,
         DP_OP_26J5_124_4249_n232, DP_OP_26J5_124_4249_n231,
         DP_OP_26J5_124_4249_n230, DP_OP_26J5_124_4249_n225,
         DP_OP_26J5_124_4249_n224, DP_OP_26J5_124_4249_n223,
         DP_OP_26J5_124_4249_n222, DP_OP_26J5_124_4249_n221,
         DP_OP_26J5_124_4249_n212, DP_OP_26J5_124_4249_n210,
         DP_OP_26J5_124_4249_n209, DP_OP_26J5_124_4249_n208,
         DP_OP_26J5_124_4249_n206, DP_OP_26J5_124_4249_n205,
         DP_OP_26J5_124_4249_n204, DP_OP_26J5_124_4249_n199,
         DP_OP_26J5_124_4249_n198, DP_OP_26J5_124_4249_n196,
         DP_OP_26J5_124_4249_n186, DP_OP_26J5_124_4249_n185,
         DP_OP_26J5_124_4249_n183, DP_OP_26J5_124_4249_n181,
         DP_OP_26J5_124_4249_n180, DP_OP_26J5_124_4249_n179,
         DP_OP_26J5_124_4249_n178, DP_OP_26J5_124_4249_n176,
         DP_OP_26J5_124_4249_n175, DP_OP_26J5_124_4249_n174,
         DP_OP_26J5_124_4249_n173, DP_OP_26J5_124_4249_n172,
         DP_OP_26J5_124_4249_n171, DP_OP_26J5_124_4249_n170,
         DP_OP_26J5_124_4249_n169, DP_OP_26J5_124_4249_n168,
         DP_OP_26J5_124_4249_n167, DP_OP_26J5_124_4249_n166,
         DP_OP_26J5_124_4249_n165, DP_OP_26J5_124_4249_n157,
         DP_OP_26J5_124_4249_n156, DP_OP_26J5_124_4249_n155,
         DP_OP_26J5_124_4249_n154, DP_OP_26J5_124_4249_n153,
         DP_OP_26J5_124_4249_n152, DP_OP_26J5_124_4249_n148,
         DP_OP_26J5_124_4249_n147, DP_OP_26J5_124_4249_n146,
         DP_OP_26J5_124_4249_n144, DP_OP_26J5_124_4249_n142,
         DP_OP_26J5_124_4249_n132, DP_OP_26J5_124_4249_n131,
         DP_OP_26J5_124_4249_n130, DP_OP_26J5_124_4249_n129,
         DP_OP_26J5_124_4249_n128, DP_OP_26J5_124_4249_n127,
         DP_OP_26J5_124_4249_n121, DP_OP_26J5_124_4249_n120,
         DP_OP_26J5_124_4249_n119, DP_OP_26J5_124_4249_n118,
         DP_OP_26J5_124_4249_n117, DP_OP_26J5_124_4249_n116,
         DP_OP_26J5_124_4249_n115, DP_OP_26J5_124_4249_n114,
         DP_OP_26J5_124_4249_n109, DP_OP_26J5_124_4249_n106,
         DP_OP_26J5_124_4249_n105, DP_OP_26J5_124_4249_n104,
         DP_OP_26J5_124_4249_n103, DP_OP_26J5_124_4249_n98,
         DP_OP_26J5_124_4249_n97, DP_OP_26J5_124_4249_n96,
         DP_OP_26J5_124_4249_n87, DP_OP_26J5_124_4249_n86,
         DP_OP_26J5_124_4249_n85, DP_OP_26J5_124_4249_n84,
         DP_OP_26J5_124_4249_n83, DP_OP_26J5_124_4249_n82,
         DP_OP_26J5_124_4249_n81, DP_OP_26J5_124_4249_n80,
         DP_OP_26J5_124_4249_n79, DP_OP_26J5_124_4249_n78,
         DP_OP_26J5_124_4249_n77, DP_OP_26J5_124_4249_n68,
         DP_OP_26J5_124_4249_n67, DP_OP_26J5_124_4249_n66,
         DP_OP_26J5_124_4249_n65, DP_OP_26J5_124_4249_n64,
         DP_OP_26J5_124_4249_n59, DP_OP_26J5_124_4249_n58,
         DP_OP_26J5_124_4249_n57, DP_OP_26J5_124_4249_n56,
         DP_OP_26J5_124_4249_n55, DP_OP_26J5_124_4249_n46,
         DP_OP_26J5_124_4249_n45, DP_OP_26J5_124_4249_n44,
         DP_OP_26J5_124_4249_n43, DP_OP_26J5_124_4249_n42,
         DP_OP_26J5_124_4249_n40, DP_OP_26J5_124_4249_n39,
         DP_OP_26J5_124_4249_n38, DP_OP_26J5_124_4249_n33,
         DP_OP_26J5_124_4249_n32, DP_OP_26J5_124_4249_n31,
         DP_OP_26J5_124_4249_n30, DP_OP_26J5_124_4249_n29,
         DP_OP_26J5_124_4249_n27, DP_OP_26J5_124_4249_n26,
         DP_OP_26J5_124_4249_n25, DP_OP_26J5_124_4249_n24,
         DP_OP_26J5_124_4249_n23, DP_OP_26J5_124_4249_n22,
         DP_OP_26J5_124_4249_n21, DP_OP_26J5_124_4249_n20,
         DP_OP_26J5_124_4249_n19, DP_OP_26J5_124_4249_n18,
         DP_OP_26J5_124_4249_n17, DP_OP_26J5_124_4249_n16,
         DP_OP_26J5_124_4249_n7, DP_OP_26J5_124_4249_n6,
         DP_OP_26J5_124_4249_n5, DP_OP_26J5_124_4249_n4,
         DP_OP_26J5_124_4249_n3, DP_OP_26J5_124_4249_n2,
         DP_OP_26J5_124_4249_n1, n1, n2, n3, n4, n5, n6, n7, n9, n10, n11, n12,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n29, n30, n31, n32, n33, n34, n35, n37, n38, n39, n40, n41, n42, n430,
         n440, n450, n460, n470, n480, n490, n500, n510, n520, n530, n540,
         n550, n560, n570, n580, n590, n600, n610, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n1130, n1140;
  wire   [7:0] n_quantized_data;

  DFFSSRX1_HVT quantized_data_reg_7_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[7]), .CLK(clk), .Q(quantized_data[7]) );
  DFFSSRX1_HVT quantized_data_reg_6_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[6]), .CLK(clk), .Q(quantized_data[6]) );
  DFFSSRX1_HVT quantized_data_reg_5_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[5]), .CLK(clk), .Q(quantized_data[5]) );
  DFFSSRX1_HVT quantized_data_reg_4_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[4]), .CLK(clk), .Q(quantized_data[4]) );
  DFFSSRX1_HVT quantized_data_reg_3_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[3]), .CLK(clk), .Q(quantized_data[3]) );
  DFFSSRX1_HVT quantized_data_reg_2_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[2]), .CLK(clk), .Q(quantized_data[2]) );
  DFFSSRX1_HVT quantized_data_reg_1_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[1]), .CLK(clk), .Q(quantized_data[1]) );
  DFFSSRX1_HVT quantized_data_reg_0_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[0]), .CLK(clk), .Q(quantized_data[0]) );
  XOR2X1_HVT DP_OP_26J5_124_4249_U253 ( .A1(DP_OP_26J5_124_4249_n245), .A2(
        DP_OP_26J5_124_4249_n157), .Y(N43) );
  XNOR2X1_HVT DP_OP_26J5_124_4249_U82 ( .A1(DP_OP_26J5_124_4249_n87), .A2(
        DP_OP_26J5_124_4249_n7), .Y(N113) );
  OAI21X1_HVT DP_OP_26J5_124_4249_U337 ( .A1(DP_OP_26J5_124_4249_n299), .A2(
        DP_OP_26J5_124_4249_n297), .A3(DP_OP_26J5_124_4249_n298), .Y(
        DP_OP_26J5_124_4249_n296) );
  OAI21X1_HVT DP_OP_26J5_124_4249_U94 ( .A1(DP_OP_26J5_124_4249_n96), .A2(
        DP_OP_26J5_124_4249_n98), .A3(DP_OP_26J5_124_4249_n97), .Y(
        DP_OP_26J5_124_4249_n87) );
  XNOR2X1_HVT DP_OP_26J5_124_4249_U223 ( .A1(DP_OP_26J5_124_4249_n223), .A2(
        DP_OP_26J5_124_4249_n155), .Y(N45) );
  XNOR2X1_HVT DP_OP_26J5_124_4249_U193 ( .A1(DP_OP_26J5_124_4249_n199), .A2(
        DP_OP_26J5_124_4249_n153), .Y(N47) );
  XNOR2X1_HVT DP_OP_26J5_124_4249_U239 ( .A1(DP_OP_26J5_124_4249_n234), .A2(
        DP_OP_26J5_124_4249_n156), .Y(N44) );
  OAI21X1_HVT DP_OP_26J5_124_4249_U254 ( .A1(DP_OP_26J5_124_4249_n243), .A2(
        DP_OP_26J5_124_4249_n245), .A3(DP_OP_26J5_124_4249_n244), .Y(
        DP_OP_26J5_124_4249_n234) );
  XOR2X1_HVT DP_OP_26J5_124_4249_U181 ( .A1(DP_OP_26J5_124_4249_n186), .A2(
        DP_OP_26J5_124_4249_n152), .Y(N48) );
  OAI21X1_HVT DP_OP_26J5_124_4249_U210 ( .A1(DP_OP_26J5_124_4249_n204), .A2(
        DP_OP_26J5_124_4249_n245), .A3(DP_OP_26J5_124_4249_n205), .Y(
        DP_OP_26J5_124_4249_n199) );
  XOR2X1_HVT DP_OP_26J5_124_4249_U209 ( .A1(DP_OP_26J5_124_4249_n210), .A2(
        DP_OP_26J5_124_4249_n154), .Y(N46) );
  OAI21X1_HVT DP_OP_26J5_124_4249_U240 ( .A1(DP_OP_26J5_124_4249_n224), .A2(
        DP_OP_26J5_124_4249_n245), .A3(DP_OP_26J5_124_4249_n225), .Y(
        DP_OP_26J5_124_4249_n223) );
  OAI21X1_HVT DP_OP_26J5_124_4249_U248 ( .A1(DP_OP_26J5_124_4249_n244), .A2(
        DP_OP_26J5_124_4249_n232), .A3(DP_OP_26J5_124_4249_n233), .Y(
        DP_OP_26J5_124_4249_n231) );
  OAI21X1_HVT DP_OP_26J5_124_4249_U299 ( .A1(DP_OP_26J5_124_4249_n281), .A2(
        DP_OP_26J5_124_4249_n271), .A3(DP_OP_26J5_124_4249_n272), .Y(
        DP_OP_26J5_124_4249_n270) );
  OAI21X1_HVT DP_OP_26J5_124_4249_U320 ( .A1(DP_OP_26J5_124_4249_n294), .A2(
        DP_OP_26J5_124_4249_n286), .A3(DP_OP_26J5_124_4249_n287), .Y(
        DP_OP_26J5_124_4249_n285) );
  XOR2X1_HVT DP_OP_26J5_124_4249_U24 ( .A1(DP_OP_26J5_124_4249_n44), .A2(
        DP_OP_26J5_124_4249_n3), .Y(N117) );
  XNOR2X1_HVT DP_OP_26J5_124_4249_U54 ( .A1(DP_OP_26J5_124_4249_n68), .A2(
        DP_OP_26J5_124_4249_n5), .Y(N115) );
  OAI21X1_HVT DP_OP_26J5_124_4249_U69 ( .A1(DP_OP_26J5_124_4249_n77), .A2(
        DP_OP_26J5_124_4249_n79), .A3(DP_OP_26J5_124_4249_n78), .Y(
        DP_OP_26J5_124_4249_n68) );
  XNOR2X1_HVT DP_OP_26J5_124_4249_U16 ( .A1(DP_OP_26J5_124_4249_n33), .A2(
        DP_OP_26J5_124_4249_n2), .Y(N118) );
  OAI21X1_HVT DP_OP_26J5_124_4249_U25 ( .A1(DP_OP_26J5_124_4249_n38), .A2(
        DP_OP_26J5_124_4249_n79), .A3(DP_OP_26J5_124_4249_n39), .Y(
        DP_OP_26J5_124_4249_n33) );
  XNOR2X1_HVT DP_OP_26J5_124_4249_U38 ( .A1(DP_OP_26J5_124_4249_n57), .A2(
        DP_OP_26J5_124_4249_n4), .Y(N116) );
  OAI21X1_HVT DP_OP_26J5_124_4249_U55 ( .A1(DP_OP_26J5_124_4249_n58), .A2(
        DP_OP_26J5_124_4249_n79), .A3(DP_OP_26J5_124_4249_n59), .Y(
        DP_OP_26J5_124_4249_n57) );
  XOR2X1_HVT DP_OP_26J5_124_4249_U68 ( .A1(DP_OP_26J5_124_4249_n79), .A2(
        DP_OP_26J5_124_4249_n6), .Y(N114) );
  OAI21X1_HVT DP_OP_26J5_124_4249_U63 ( .A1(DP_OP_26J5_124_4249_n78), .A2(
        DP_OP_26J5_124_4249_n66), .A3(DP_OP_26J5_124_4249_n67), .Y(
        DP_OP_26J5_124_4249_n65) );
  OAI21X1_HVT DP_OP_26J5_124_4249_U88 ( .A1(DP_OP_26J5_124_4249_n97), .A2(
        DP_OP_26J5_124_4249_n85), .A3(DP_OP_26J5_124_4249_n86), .Y(
        DP_OP_26J5_124_4249_n84) );
  OAI21X1_HVT DP_OP_26J5_124_4249_U114 ( .A1(DP_OP_26J5_124_4249_n115), .A2(
        DP_OP_26J5_124_4249_n105), .A3(DP_OP_26J5_124_4249_n106), .Y(
        DP_OP_26J5_124_4249_n104) );
  OAI21X1_HVT DP_OP_26J5_124_4249_U135 ( .A1(DP_OP_26J5_124_4249_n128), .A2(
        DP_OP_26J5_124_4249_n120), .A3(DP_OP_26J5_124_4249_n121), .Y(
        DP_OP_26J5_124_4249_n119) );
  NOR2X0_HVT DP_OP_26J5_124_4249_U343 ( .A1(bias_data[0]), .A2(ori_data_5_), 
        .Y(DP_OP_26J5_124_4249_n299) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U341 ( .A1(ori_data_6_), .A2(bias_data[1]), 
        .Y(DP_OP_26J5_124_4249_n298) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U334 ( .A1(ori_data_7_), .A2(bias_data[2]), 
        .Y(DP_OP_26J5_124_4249_n294) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U324 ( .A1(ori_data_8_), .A2(n65), .Y(
        DP_OP_26J5_124_4249_n287) );
  NOR2X0_HVT DP_OP_26J5_124_4249_U323 ( .A1(n68), .A2(ori_data_8_), .Y(
        DP_OP_26J5_124_4249_n286) );
  NOR2X0_HVT DP_OP_26J5_124_4249_U319 ( .A1(DP_OP_26J5_124_4249_n286), .A2(
        DP_OP_26J5_124_4249_n293), .Y(DP_OP_26J5_124_4249_n284) );
  AOI21X1_HVT DP_OP_26J5_124_4249_U318 ( .A1(DP_OP_26J5_124_4249_n296), .A2(
        DP_OP_26J5_124_4249_n284), .A3(DP_OP_26J5_124_4249_n285), .Y(
        DP_OP_26J5_124_4249_n283) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U315 ( .A1(ori_data_9_), .A2(n68), .Y(
        DP_OP_26J5_124_4249_n281) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U303 ( .A1(ori_data_10_), .A2(n68), .Y(
        DP_OP_26J5_124_4249_n272) );
  NOR2X0_HVT DP_OP_26J5_124_4249_U302 ( .A1(n68), .A2(ori_data_10_), .Y(
        DP_OP_26J5_124_4249_n271) );
  NOR2X0_HVT DP_OP_26J5_124_4249_U298 ( .A1(DP_OP_26J5_124_4249_n271), .A2(
        DP_OP_26J5_124_4249_n280), .Y(DP_OP_26J5_124_4249_n269) );
  AOI21X1_HVT DP_OP_26J5_124_4249_U293 ( .A1(DP_OP_26J5_124_4249_n282), .A2(
        DP_OP_26J5_124_4249_n269), .A3(DP_OP_26J5_124_4249_n270), .Y(
        DP_OP_26J5_124_4249_n264) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U291 ( .A1(ori_data_11_), .A2(n68), .Y(
        DP_OP_26J5_124_4249_n263) );
  NOR2X0_HVT DP_OP_26J5_124_4249_U290 ( .A1(n68), .A2(ori_data_11_), .Y(
        DP_OP_26J5_124_4249_n262) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U277 ( .A1(ori_data_12_), .A2(n65), .Y(
        DP_OP_26J5_124_4249_n252) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U266 ( .A1(ori_data_13_), .A2(n68), .Y(
        DP_OP_26J5_124_4249_n244) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U263 ( .A1(DP_OP_26J5_124_4249_n306), .A2(
        DP_OP_26J5_124_4249_n244), .Y(DP_OP_26J5_124_4249_n157) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U252 ( .A1(ori_data_14_), .A2(n590), .Y(
        DP_OP_26J5_124_4249_n233) );
  NOR2X0_HVT DP_OP_26J5_124_4249_U251 ( .A1(n68), .A2(ori_data_14_), .Y(
        DP_OP_26J5_124_4249_n232) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U249 ( .A1(DP_OP_26J5_124_4249_n142), .A2(
        DP_OP_26J5_124_4249_n233), .Y(DP_OP_26J5_124_4249_n156) );
  NOR2X0_HVT DP_OP_26J5_124_4249_U247 ( .A1(DP_OP_26J5_124_4249_n232), .A2(
        DP_OP_26J5_124_4249_n243), .Y(DP_OP_26J5_124_4249_n230) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U238 ( .A1(ori_data_15_), .A2(n68), .Y(
        DP_OP_26J5_124_4249_n222) );
  NOR2X0_HVT DP_OP_26J5_124_4249_U237 ( .A1(n65), .A2(ori_data_15_), .Y(
        DP_OP_26J5_124_4249_n221) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U235 ( .A1(DP_OP_26J5_124_4249_n304), .A2(
        DP_OP_26J5_124_4249_n222), .Y(DP_OP_26J5_124_4249_n155) );
  AOI21X1_HVT DP_OP_26J5_124_4249_U224 ( .A1(DP_OP_26J5_124_4249_n223), .A2(
        DP_OP_26J5_124_4249_n304), .A3(DP_OP_26J5_124_4249_n212), .Y(
        DP_OP_26J5_124_4249_n210) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U222 ( .A1(ori_data_16_), .A2(n65), .Y(
        DP_OP_26J5_124_4249_n209) );
  NOR2X0_HVT DP_OP_26J5_124_4249_U221 ( .A1(n68), .A2(ori_data_16_), .Y(
        DP_OP_26J5_124_4249_n208) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U219 ( .A1(DP_OP_26J5_124_4249_n45), .A2(
        DP_OP_26J5_124_4249_n209), .Y(DP_OP_26J5_124_4249_n154) );
  NOR2X0_HVT DP_OP_26J5_124_4249_U217 ( .A1(DP_OP_26J5_124_4249_n208), .A2(
        DP_OP_26J5_124_4249_n221), .Y(DP_OP_26J5_124_4249_n206) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U215 ( .A1(DP_OP_26J5_124_4249_n230), .A2(
        DP_OP_26J5_124_4249_n206), .Y(DP_OP_26J5_124_4249_n204) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U208 ( .A1(ori_data_17_), .A2(n66), .Y(
        DP_OP_26J5_124_4249_n198) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U205 ( .A1(n70), .A2(
        DP_OP_26J5_124_4249_n198), .Y(DP_OP_26J5_124_4249_n153) );
  AOI21X1_HVT DP_OP_26J5_124_4249_U194 ( .A1(DP_OP_26J5_124_4249_n199), .A2(
        n70), .A3(DP_OP_26J5_124_4249_n196), .Y(DP_OP_26J5_124_4249_n186) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U192 ( .A1(ori_data_18_), .A2(n67), .Y(
        DP_OP_26J5_124_4249_n185) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U189 ( .A1(n73), .A2(
        DP_OP_26J5_124_4249_n185), .Y(DP_OP_26J5_124_4249_n152) );
  AOI21X1_HVT DP_OP_26J5_124_4249_U186 ( .A1(n73), .A2(
        DP_OP_26J5_124_4249_n196), .A3(DP_OP_26J5_124_4249_n183), .Y(
        DP_OP_26J5_124_4249_n181) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U185 ( .A1(n70), .A2(n73), .Y(
        DP_OP_26J5_124_4249_n180) );
  NOR2X0_HVT DP_OP_26J5_124_4249_U183 ( .A1(DP_OP_26J5_124_4249_n180), .A2(
        DP_OP_26J5_124_4249_n204), .Y(DP_OP_26J5_124_4249_n178) );
  FADDX1_HVT DP_OP_26J5_124_4249_U179 ( .A(n600), .B(ori_data_19_), .CI(n72), 
        .CO(DP_OP_26J5_124_4249_n176), .S(N49) );
  FADDX1_HVT DP_OP_26J5_124_4249_U178 ( .A(n65), .B(ori_data_20_), .CI(
        DP_OP_26J5_124_4249_n176), .CO(DP_OP_26J5_124_4249_n175), .S(N50) );
  FADDX1_HVT DP_OP_26J5_124_4249_U177 ( .A(n67), .B(ori_data_21_), .CI(
        DP_OP_26J5_124_4249_n175), .CO(DP_OP_26J5_124_4249_n174), .S(N51) );
  FADDX1_HVT DP_OP_26J5_124_4249_U176 ( .A(n63), .B(ori_data_22_), .CI(
        DP_OP_26J5_124_4249_n174), .CO(DP_OP_26J5_124_4249_n173), .S(N52) );
  FADDX1_HVT DP_OP_26J5_124_4249_U175 ( .A(bias_data[3]), .B(ori_data_23_), 
        .CI(DP_OP_26J5_124_4249_n173), .CO(DP_OP_26J5_124_4249_n172), .S(N53)
         );
  FADDX1_HVT DP_OP_26J5_124_4249_U174 ( .A(n66), .B(ori_data_24_), .CI(
        DP_OP_26J5_124_4249_n172), .CO(DP_OP_26J5_124_4249_n171), .S(N54) );
  FADDX1_HVT DP_OP_26J5_124_4249_U173 ( .A(n65), .B(ori_data_25_), .CI(
        DP_OP_26J5_124_4249_n171), .CO(DP_OP_26J5_124_4249_n170), .S(N55) );
  FADDX1_HVT DP_OP_26J5_124_4249_U172 ( .A(n67), .B(ori_data_26_), .CI(
        DP_OP_26J5_124_4249_n170), .CO(DP_OP_26J5_124_4249_n169), .S(N56) );
  FADDX1_HVT DP_OP_26J5_124_4249_U171 ( .A(n66), .B(ori_data_27_), .CI(
        DP_OP_26J5_124_4249_n169), .CO(DP_OP_26J5_124_4249_n168), .S(N57) );
  FADDX1_HVT DP_OP_26J5_124_4249_U170 ( .A(n600), .B(ori_data_28_), .CI(
        DP_OP_26J5_124_4249_n168), .CO(DP_OP_26J5_124_4249_n167), .S(N58) );
  FADDX1_HVT DP_OP_26J5_124_4249_U169 ( .A(n67), .B(ori_data_29_), .CI(
        DP_OP_26J5_124_4249_n167), .CO(DP_OP_26J5_124_4249_n166), .S(N59) );
  FADDX1_HVT DP_OP_26J5_124_4249_U168 ( .A(n66), .B(ori_data_30_), .CI(
        DP_OP_26J5_124_4249_n166), .CO(DP_OP_26J5_124_4249_n165), .S(N60) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U157 ( .A1(ori_data_5_), .A2(ori_data_6_), 
        .Y(DP_OP_26J5_124_4249_n132) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U149 ( .A1(ori_data_8_), .A2(bias_data[0]), 
        .Y(DP_OP_26J5_124_4249_n128) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U139 ( .A1(ori_data_9_), .A2(bias_data[1]), 
        .Y(DP_OP_26J5_124_4249_n121) );
  NOR2X0_HVT DP_OP_26J5_124_4249_U134 ( .A1(DP_OP_26J5_124_4249_n120), .A2(
        DP_OP_26J5_124_4249_n127), .Y(DP_OP_26J5_124_4249_n118) );
  AOI21X1_HVT DP_OP_26J5_124_4249_U133 ( .A1(DP_OP_26J5_124_4249_n118), .A2(
        DP_OP_26J5_124_4249_n130), .A3(DP_OP_26J5_124_4249_n119), .Y(
        DP_OP_26J5_124_4249_n117) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U130 ( .A1(ori_data_10_), .A2(bias_data[2]), 
        .Y(DP_OP_26J5_124_4249_n115) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U118 ( .A1(ori_data_11_), .A2(n63), .Y(
        DP_OP_26J5_124_4249_n106) );
  NOR2X0_HVT DP_OP_26J5_124_4249_U113 ( .A1(DP_OP_26J5_124_4249_n105), .A2(
        DP_OP_26J5_124_4249_n114), .Y(DP_OP_26J5_124_4249_n103) );
  AOI21X1_HVT DP_OP_26J5_124_4249_U108 ( .A1(DP_OP_26J5_124_4249_n116), .A2(
        DP_OP_26J5_124_4249_n103), .A3(DP_OP_26J5_124_4249_n104), .Y(
        DP_OP_26J5_124_4249_n98) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U106 ( .A1(ori_data_12_), .A2(n63), .Y(
        DP_OP_26J5_124_4249_n97) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U92 ( .A1(ori_data_13_), .A2(n610), .Y(
        DP_OP_26J5_124_4249_n86) );
  NOR2X0_HVT DP_OP_26J5_124_4249_U91 ( .A1(n63), .A2(ori_data_13_), .Y(
        DP_OP_26J5_124_4249_n85) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U89 ( .A1(DP_OP_26J5_124_4249_n306), .A2(
        DP_OP_26J5_124_4249_n86), .Y(DP_OP_26J5_124_4249_n7) );
  NOR2X0_HVT DP_OP_26J5_124_4249_U87 ( .A1(DP_OP_26J5_124_4249_n85), .A2(
        DP_OP_26J5_124_4249_n96), .Y(DP_OP_26J5_124_4249_n83) );
  AOI21X1_HVT DP_OP_26J5_124_4249_U86 ( .A1(DP_OP_26J5_124_4249_n104), .A2(
        DP_OP_26J5_124_4249_n83), .A3(DP_OP_26J5_124_4249_n84), .Y(
        DP_OP_26J5_124_4249_n82) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U85 ( .A1(DP_OP_26J5_124_4249_n103), .A2(
        DP_OP_26J5_124_4249_n83), .Y(DP_OP_26J5_124_4249_n81) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U81 ( .A1(ori_data_14_), .A2(n63), .Y(
        DP_OP_26J5_124_4249_n78) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U78 ( .A1(DP_OP_26J5_124_4249_n142), .A2(
        DP_OP_26J5_124_4249_n78), .Y(DP_OP_26J5_124_4249_n6) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U67 ( .A1(ori_data_15_), .A2(n64), .Y(
        DP_OP_26J5_124_4249_n67) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U64 ( .A1(DP_OP_26J5_124_4249_n304), .A2(
        DP_OP_26J5_124_4249_n67), .Y(DP_OP_26J5_124_4249_n5) );
  NOR2X0_HVT DP_OP_26J5_124_4249_U62 ( .A1(DP_OP_26J5_124_4249_n66), .A2(
        DP_OP_26J5_124_4249_n77), .Y(DP_OP_26J5_124_4249_n64) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U53 ( .A1(ori_data_16_), .A2(n63), .Y(
        DP_OP_26J5_124_4249_n56) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U50 ( .A1(DP_OP_26J5_124_4249_n45), .A2(
        DP_OP_26J5_124_4249_n56), .Y(DP_OP_26J5_124_4249_n4) );
  AOI21X1_HVT DP_OP_26J5_124_4249_U39 ( .A1(DP_OP_26J5_124_4249_n57), .A2(
        DP_OP_26J5_124_4249_n45), .A3(DP_OP_26J5_124_4249_n46), .Y(
        DP_OP_26J5_124_4249_n44) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U37 ( .A1(ori_data_17_), .A2(n64), .Y(
        DP_OP_26J5_124_4249_n43) );
  NOR2X0_HVT DP_OP_26J5_124_4249_U36 ( .A1(n63), .A2(ori_data_17_), .Y(
        DP_OP_26J5_124_4249_n42) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U34 ( .A1(n70), .A2(DP_OP_26J5_124_4249_n43), 
        .Y(DP_OP_26J5_124_4249_n3) );
  NOR2X0_HVT DP_OP_26J5_124_4249_U32 ( .A1(DP_OP_26J5_124_4249_n42), .A2(
        DP_OP_26J5_124_4249_n55), .Y(DP_OP_26J5_124_4249_n40) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U30 ( .A1(DP_OP_26J5_124_4249_n64), .A2(
        DP_OP_26J5_124_4249_n40), .Y(DP_OP_26J5_124_4249_n38) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U23 ( .A1(ori_data_18_), .A2(n64), .Y(
        DP_OP_26J5_124_4249_n32) );
  NOR2X0_HVT DP_OP_26J5_124_4249_U22 ( .A1(n64), .A2(ori_data_18_), .Y(
        DP_OP_26J5_124_4249_n31) );
  NAND2X0_HVT DP_OP_26J5_124_4249_U20 ( .A1(n73), .A2(DP_OP_26J5_124_4249_n32), 
        .Y(DP_OP_26J5_124_4249_n2) );
  FADDX1_HVT DP_OP_26J5_124_4249_U14 ( .A(n590), .B(ori_data_19_), .CI(n71), 
        .CO(DP_OP_26J5_124_4249_n27), .S(N119) );
  FADDX1_HVT DP_OP_26J5_124_4249_U13 ( .A(n610), .B(ori_data_20_), .CI(
        DP_OP_26J5_124_4249_n27), .CO(DP_OP_26J5_124_4249_n26), .S(N120) );
  FADDX1_HVT DP_OP_26J5_124_4249_U12 ( .A(n64), .B(ori_data_21_), .CI(
        DP_OP_26J5_124_4249_n26), .CO(DP_OP_26J5_124_4249_n25), .S(N121) );
  FADDX1_HVT DP_OP_26J5_124_4249_U11 ( .A(n590), .B(ori_data_22_), .CI(
        DP_OP_26J5_124_4249_n25), .CO(DP_OP_26J5_124_4249_n24), .S(N122) );
  FADDX1_HVT DP_OP_26J5_124_4249_U10 ( .A(n590), .B(ori_data_23_), .CI(
        DP_OP_26J5_124_4249_n24), .CO(DP_OP_26J5_124_4249_n23), .S(N123) );
  FADDX1_HVT DP_OP_26J5_124_4249_U9 ( .A(n610), .B(ori_data_24_), .CI(
        DP_OP_26J5_124_4249_n23), .CO(DP_OP_26J5_124_4249_n22), .S(N124) );
  FADDX1_HVT DP_OP_26J5_124_4249_U8 ( .A(n64), .B(ori_data_25_), .CI(
        DP_OP_26J5_124_4249_n22), .CO(DP_OP_26J5_124_4249_n21), .S(N125) );
  FADDX1_HVT DP_OP_26J5_124_4249_U7 ( .A(n610), .B(ori_data_26_), .CI(
        DP_OP_26J5_124_4249_n21), .CO(DP_OP_26J5_124_4249_n20), .S(N126) );
  FADDX1_HVT DP_OP_26J5_124_4249_U6 ( .A(n62), .B(ori_data_27_), .CI(
        DP_OP_26J5_124_4249_n20), .CO(DP_OP_26J5_124_4249_n19), .S(N127) );
  FADDX1_HVT DP_OP_26J5_124_4249_U5 ( .A(n600), .B(ori_data_28_), .CI(
        DP_OP_26J5_124_4249_n19), .CO(DP_OP_26J5_124_4249_n18), .S(N128) );
  FADDX1_HVT DP_OP_26J5_124_4249_U4 ( .A(n62), .B(ori_data_29_), .CI(
        DP_OP_26J5_124_4249_n18), .CO(DP_OP_26J5_124_4249_n17), .S(N129) );
  FADDX1_HVT DP_OP_26J5_124_4249_U3 ( .A(n62), .B(ori_data_30_), .CI(
        DP_OP_26J5_124_4249_n17), .CO(DP_OP_26J5_124_4249_n16), .S(N130) );
  XNOR2X1_HVT DP_OP_26J5_124_4249_U2 ( .A1(ori_data_31_), .A2(bias_data[3]), 
        .Y(DP_OP_26J5_124_4249_n1) );
  NOR2X1_HVT DP_OP_26J5_124_4249_U129 ( .A1(bias_data[2]), .A2(ori_data_10_), 
        .Y(DP_OP_26J5_124_4249_n114) );
  NOR2X1_HVT DP_OP_26J5_124_4249_U333 ( .A1(bias_data[2]), .A2(ori_data_7_), 
        .Y(DP_OP_26J5_124_4249_n293) );
  NOR2X1_HVT DP_OP_26J5_124_4249_U117 ( .A1(n63), .A2(ori_data_11_), .Y(
        DP_OP_26J5_124_4249_n105) );
  NOR2X1_HVT DP_OP_26J5_124_4249_U138 ( .A1(bias_data[1]), .A2(ori_data_9_), 
        .Y(DP_OP_26J5_124_4249_n120) );
  NOR2X1_HVT DP_OP_26J5_124_4249_U148 ( .A1(bias_data[0]), .A2(ori_data_8_), 
        .Y(DP_OP_26J5_124_4249_n127) );
  NOR2X1_HVT DP_OP_26J5_124_4249_U18 ( .A1(DP_OP_26J5_124_4249_n31), .A2(
        DP_OP_26J5_124_4249_n38), .Y(DP_OP_26J5_124_4249_n29) );
  OAI21X1_HVT DP_OP_26J5_124_4249_U19 ( .A1(DP_OP_26J5_124_4249_n31), .A2(
        DP_OP_26J5_124_4249_n39), .A3(DP_OP_26J5_124_4249_n32), .Y(
        DP_OP_26J5_124_4249_n30) );
  OAI21X1_HVT DP_OP_26J5_124_4249_U84 ( .A1(DP_OP_26J5_124_4249_n81), .A2(
        DP_OP_26J5_124_4249_n117), .A3(DP_OP_26J5_124_4249_n82), .Y(
        DP_OP_26J5_124_4249_n80) );
  OAI21X1_HVT DP_OP_26J5_124_4249_U184 ( .A1(DP_OP_26J5_124_4249_n180), .A2(
        DP_OP_26J5_124_4249_n205), .A3(DP_OP_26J5_124_4249_n181), .Y(
        DP_OP_26J5_124_4249_n179) );
  XOR2X1_HVT DP_OP_26J5_124_4249_U1 ( .A1(DP_OP_26J5_124_4249_n16), .A2(n570), 
        .Y(N131) );
  XOR2X1_HVT DP_OP_26J5_124_4249_U166 ( .A1(DP_OP_26J5_124_4249_n165), .A2(
        n580), .Y(N61) );
  NOR2X1_HVT DP_OP_26J5_124_4249_U340 ( .A1(bias_data[1]), .A2(ori_data_6_), 
        .Y(DP_OP_26J5_124_4249_n297) );
  NOR2X1_HVT DP_OP_26J5_124_4249_U265 ( .A1(n600), .A2(ori_data_13_), .Y(
        DP_OP_26J5_124_4249_n243) );
  NOR2X1_HVT DP_OP_26J5_124_4249_U52 ( .A1(n63), .A2(ori_data_16_), .Y(
        DP_OP_26J5_124_4249_n55) );
  NOR2X1_HVT DP_OP_26J5_124_4249_U66 ( .A1(n63), .A2(ori_data_15_), .Y(
        DP_OP_26J5_124_4249_n66) );
  NOR2X1_HVT DP_OP_26J5_124_4249_U105 ( .A1(n63), .A2(ori_data_12_), .Y(
        DP_OP_26J5_124_4249_n96) );
  NOR2X1_HVT DP_OP_26J5_124_4249_U80 ( .A1(n64), .A2(ori_data_14_), .Y(
        DP_OP_26J5_124_4249_n77) );
  NOR2X1_HVT DP_OP_26J5_124_4249_U314 ( .A1(n65), .A2(ori_data_9_), .Y(
        DP_OP_26J5_124_4249_n280) );
  NOR2X0_HVT DP_OP_26J5_124_4249_U152 ( .A1(DP_OP_26J5_124_4249_n131), .A2(
        DP_OP_26J5_124_4249_n132), .Y(DP_OP_26J5_124_4249_n130) );
  OA221X1_HVT U3 ( .A1(1'b0), .A2(DP_OP_26J5_124_4249_n43), .A3(
        DP_OP_26J5_124_4249_n42), .A4(DP_OP_26J5_124_4249_n56), .A5(n35), .Y(
        DP_OP_26J5_124_4249_n39) );
  OA221X1_HVT U4 ( .A1(1'b0), .A2(DP_OP_26J5_124_4249_n209), .A3(
        DP_OP_26J5_124_4249_n208), .A4(DP_OP_26J5_124_4249_n222), .A5(n29), 
        .Y(DP_OP_26J5_124_4249_n205) );
  INVX0_HVT U5 ( .A(DP_OP_26J5_124_4249_n262), .Y(n1) );
  OA21X1_HVT U6 ( .A1(ori_data_12_), .A2(n68), .A3(n1), .Y(n2) );
  INVX0_HVT U7 ( .A(DP_OP_26J5_124_4249_n283), .Y(n3) );
  NAND3X0_HVT U8 ( .A1(DP_OP_26J5_124_4249_n269), .A2(n2), .A3(n3), .Y(n4) );
  NAND2X0_HVT U9 ( .A1(n2), .A2(DP_OP_26J5_124_4249_n270), .Y(n5) );
  OR2X1_HVT U10 ( .A1(ori_data_12_), .A2(n68), .Y(n6) );
  INVX0_HVT U11 ( .A(DP_OP_26J5_124_4249_n263), .Y(n7) );
  NAND2X0_HVT U12 ( .A1(n6), .A2(n7), .Y(n9) );
  NAND4X0_HVT U13 ( .A1(DP_OP_26J5_124_4249_n252), .A2(n4), .A3(n5), .A4(n9), 
        .Y(DP_OP_26J5_124_4249_n246) );
  INVX0_HVT U14 ( .A(DP_OP_26J5_124_4249_n297), .Y(n10) );
  NAND2X0_HVT U15 ( .A1(n10), .A2(DP_OP_26J5_124_4249_n298), .Y(n11) );
  HADDX1_HVT U16 ( .A0(DP_OP_26J5_124_4249_n299), .B0(n11), .SO(n12) );
  HADDX1_HVT U17 ( .A0(ori_data_6_), .B0(ori_data_5_), .SO(n14) );
  AOI22X1_HVT U18 ( .A1(n104), .A2(n12), .A3(n14), .A4(n105), .Y(n15) );
  NAND2X0_HVT U19 ( .A1(n106), .A2(n15), .Y(n_quantized_data[0]) );
  OA21X1_HVT U20 ( .A1(DP_OP_26J5_124_4249_n293), .A2(DP_OP_26J5_124_4249_n295), .A3(DP_OP_26J5_124_4249_n294), .Y(n16) );
  NAND2X0_HVT U21 ( .A1(DP_OP_26J5_124_4249_n311), .A2(
        DP_OP_26J5_124_4249_n287), .Y(n17) );
  HADDX1_HVT U22 ( .A0(n16), .B0(n17), .SO(n18) );
  NAND2X0_HVT U23 ( .A1(DP_OP_26J5_124_4249_n148), .A2(
        DP_OP_26J5_124_4249_n128), .Y(n19) );
  HADDX1_HVT U24 ( .A0(DP_OP_26J5_124_4249_n129), .B0(n19), .SO(n20) );
  AOI22X1_HVT U25 ( .A1(n104), .A2(n18), .A3(n105), .A4(n20), .Y(n21) );
  NAND2X0_HVT U26 ( .A1(n106), .A2(n21), .Y(n_quantized_data[2]) );
  AND2X1_HVT U27 ( .A1(DP_OP_26J5_124_4249_n310), .A2(DP_OP_26J5_124_4249_n281), .Y(n22) );
  HADDX1_HVT U28 ( .A0(n22), .B0(DP_OP_26J5_124_4249_n282), .SO(n23) );
  OA21X1_HVT U29 ( .A1(DP_OP_26J5_124_4249_n127), .A2(DP_OP_26J5_124_4249_n129), .A3(DP_OP_26J5_124_4249_n128), .Y(n24) );
  NAND2X0_HVT U30 ( .A1(DP_OP_26J5_124_4249_n147), .A2(
        DP_OP_26J5_124_4249_n121), .Y(n25) );
  HADDX1_HVT U31 ( .A0(n24), .B0(n25), .SO(n26) );
  AOI22X1_HVT U32 ( .A1(n104), .A2(n23), .A3(n105), .A4(n26), .Y(n27) );
  NAND2X0_HVT U33 ( .A1(n106), .A2(n27), .Y(n_quantized_data[3]) );
  NAND2X0_HVT U35 ( .A1(DP_OP_26J5_124_4249_n206), .A2(
        DP_OP_26J5_124_4249_n231), .Y(n29) );
  INVX0_HVT U36 ( .A(DP_OP_26J5_124_4249_n293), .Y(n30) );
  NAND2X0_HVT U37 ( .A1(n30), .A2(DP_OP_26J5_124_4249_n294), .Y(n31) );
  HADDX1_HVT U38 ( .A0(DP_OP_26J5_124_4249_n295), .B0(n31), .SO(n32) );
  HADDX1_HVT U39 ( .A0(DP_OP_26J5_124_4249_n132), .B0(DP_OP_26J5_124_4249_n131), .SO(n33) );
  AOI22X1_HVT U40 ( .A1(n104), .A2(n32), .A3(n33), .A4(n105), .Y(n34) );
  NAND2X0_HVT U41 ( .A1(n106), .A2(n34), .Y(n_quantized_data[1]) );
  NAND2X0_HVT U42 ( .A1(DP_OP_26J5_124_4249_n40), .A2(DP_OP_26J5_124_4249_n65), 
        .Y(n35) );
  AO21X1_HVT U44 ( .A1(DP_OP_26J5_124_4249_n282), .A2(DP_OP_26J5_124_4249_n310), .A3(DP_OP_26J5_124_4249_n275), .Y(n37) );
  NAND2X0_HVT U45 ( .A1(DP_OP_26J5_124_4249_n309), .A2(
        DP_OP_26J5_124_4249_n272), .Y(n38) );
  HADDX1_HVT U46 ( .A0(n37), .B0(n38), .SO(n39) );
  INVX0_HVT U47 ( .A(n104), .Y(n40) );
  NAND2X0_HVT U48 ( .A1(DP_OP_26J5_124_4249_n146), .A2(
        DP_OP_26J5_124_4249_n115), .Y(n41) );
  HADDX1_HVT U49 ( .A0(DP_OP_26J5_124_4249_n116), .B0(n41), .SO(n42) );
  INVX0_HVT U50 ( .A(n105), .Y(n430) );
  OA22X1_HVT U51 ( .A1(n39), .A2(n40), .A3(n42), .A4(n430), .Y(n440) );
  NAND2X0_HVT U52 ( .A1(n106), .A2(n440), .Y(n_quantized_data[4]) );
  NAND2X0_HVT U53 ( .A1(DP_OP_26J5_124_4249_n308), .A2(
        DP_OP_26J5_124_4249_n263), .Y(n450) );
  HADDX1_HVT U54 ( .A0(DP_OP_26J5_124_4249_n264), .B0(n450), .SO(n460) );
  AOI21X1_HVT U55 ( .A1(DP_OP_26J5_124_4249_n116), .A2(
        DP_OP_26J5_124_4249_n146), .A3(DP_OP_26J5_124_4249_n109), .Y(n470) );
  NAND2X0_HVT U56 ( .A1(DP_OP_26J5_124_4249_n106), .A2(
        DP_OP_26J5_124_4249_n308), .Y(n480) );
  HADDX1_HVT U57 ( .A0(n470), .B0(n480), .SO(n490) );
  AOI22X1_HVT U58 ( .A1(n104), .A2(n460), .A3(n105), .A4(n490), .Y(n500) );
  NAND2X0_HVT U59 ( .A1(n106), .A2(n500), .Y(n_quantized_data[5]) );
  OA21X1_HVT U60 ( .A1(DP_OP_26J5_124_4249_n262), .A2(DP_OP_26J5_124_4249_n264), .A3(DP_OP_26J5_124_4249_n263), .Y(n510) );
  NAND2X0_HVT U61 ( .A1(DP_OP_26J5_124_4249_n144), .A2(
        DP_OP_26J5_124_4249_n252), .Y(n520) );
  HADDX1_HVT U62 ( .A0(n510), .B0(n520), .SO(n530) );
  NAND2X0_HVT U63 ( .A1(DP_OP_26J5_124_4249_n97), .A2(DP_OP_26J5_124_4249_n144), .Y(n540) );
  HADDX1_HVT U64 ( .A0(DP_OP_26J5_124_4249_n98), .B0(n540), .SO(n550) );
  AOI22X1_HVT U65 ( .A1(n104), .A2(n530), .A3(n105), .A4(n550), .Y(n560) );
  NAND2X0_HVT U66 ( .A1(n106), .A2(n560), .Y(n_quantized_data[6]) );
  INVX0_HVT U67 ( .A(DP_OP_26J5_124_4249_n117), .Y(DP_OP_26J5_124_4249_n116)
         );
  INVX0_HVT U68 ( .A(DP_OP_26J5_124_4249_n283), .Y(DP_OP_26J5_124_4249_n282)
         );
  INVX0_HVT U69 ( .A(DP_OP_26J5_124_4249_n296), .Y(DP_OP_26J5_124_4249_n295)
         );
  INVX0_HVT U70 ( .A(DP_OP_26J5_124_4249_n130), .Y(DP_OP_26J5_124_4249_n129)
         );
  INVX0_HVT U71 ( .A(DP_OP_26J5_124_4249_n114), .Y(DP_OP_26J5_124_4249_n146)
         );
  INVX0_HVT U72 ( .A(DP_OP_26J5_124_4249_n280), .Y(DP_OP_26J5_124_4249_n310)
         );
  INVX1_HVT U73 ( .A(n69), .Y(n63) );
  OR2X1_HVT U74 ( .A1(n1140), .A2(n112), .Y(n106) );
  INVX0_HVT U75 ( .A(DP_OP_26J5_124_4249_n80), .Y(DP_OP_26J5_124_4249_n79) );
  INVX0_HVT U76 ( .A(DP_OP_26J5_124_4249_n246), .Y(DP_OP_26J5_124_4249_n245)
         );
  INVX0_HVT U77 ( .A(DP_OP_26J5_124_4249_n230), .Y(DP_OP_26J5_124_4249_n224)
         );
  INVX1_HVT U78 ( .A(DP_OP_26J5_124_4249_n1), .Y(n580) );
  INVX0_HVT U79 ( .A(DP_OP_26J5_124_4249_n231), .Y(DP_OP_26J5_124_4249_n225)
         );
  INVX0_HVT U80 ( .A(DP_OP_26J5_124_4249_n65), .Y(DP_OP_26J5_124_4249_n59) );
  INVX0_HVT U81 ( .A(DP_OP_26J5_124_4249_n64), .Y(DP_OP_26J5_124_4249_n58) );
  INVX1_HVT U82 ( .A(DP_OP_26J5_124_4249_n1), .Y(n570) );
  INVX0_HVT U83 ( .A(DP_OP_26J5_124_4249_n222), .Y(DP_OP_26J5_124_4249_n212)
         );
  INVX0_HVT U84 ( .A(DP_OP_26J5_124_4249_n271), .Y(DP_OP_26J5_124_4249_n309)
         );
  INVX0_HVT U85 ( .A(DP_OP_26J5_124_4249_n56), .Y(DP_OP_26J5_124_4249_n46) );
  INVX0_HVT U86 ( .A(DP_OP_26J5_124_4249_n221), .Y(DP_OP_26J5_124_4249_n304)
         );
  INVX0_HVT U87 ( .A(DP_OP_26J5_124_4249_n55), .Y(DP_OP_26J5_124_4249_n45) );
  INVX0_HVT U88 ( .A(DP_OP_26J5_124_4249_n243), .Y(DP_OP_26J5_124_4249_n306)
         );
  INVX0_HVT U89 ( .A(DP_OP_26J5_124_4249_n281), .Y(DP_OP_26J5_124_4249_n275)
         );
  INVX0_HVT U90 ( .A(DP_OP_26J5_124_4249_n77), .Y(DP_OP_26J5_124_4249_n142) );
  INVX0_HVT U91 ( .A(DP_OP_26J5_124_4249_n120), .Y(DP_OP_26J5_124_4249_n147)
         );
  INVX0_HVT U92 ( .A(DP_OP_26J5_124_4249_n96), .Y(DP_OP_26J5_124_4249_n144) );
  INVX0_HVT U93 ( .A(DP_OP_26J5_124_4249_n115), .Y(DP_OP_26J5_124_4249_n109)
         );
  INVX0_HVT U94 ( .A(DP_OP_26J5_124_4249_n262), .Y(DP_OP_26J5_124_4249_n308)
         );
  INVX0_HVT U95 ( .A(DP_OP_26J5_124_4249_n185), .Y(DP_OP_26J5_124_4249_n183)
         );
  INVX0_HVT U96 ( .A(DP_OP_26J5_124_4249_n127), .Y(DP_OP_26J5_124_4249_n148)
         );
  INVX0_HVT U97 ( .A(DP_OP_26J5_124_4249_n286), .Y(DP_OP_26J5_124_4249_n311)
         );
  INVX1_HVT U98 ( .A(n69), .Y(n590) );
  INVX1_HVT U99 ( .A(n69), .Y(n600) );
  INVX1_HVT U100 ( .A(n69), .Y(n64) );
  INVX1_HVT U101 ( .A(n69), .Y(n610) );
  INVX0_HVT U102 ( .A(n96), .Y(n103) );
  INVX0_HVT U103 ( .A(mode[0]), .Y(n81) );
  INVX1_HVT U104 ( .A(bias_data[3]), .Y(n69) );
  INVX0_HVT U105 ( .A(srstn), .Y(n13) );
  INVX1_HVT U106 ( .A(n69), .Y(n62) );
  INVX1_HVT U107 ( .A(n69), .Y(n68) );
  INVX1_HVT U108 ( .A(n69), .Y(n67) );
  INVX1_HVT U109 ( .A(n69), .Y(n66) );
  INVX1_HVT U110 ( .A(n69), .Y(n65) );
  INVX1_HVT U111 ( .A(ori_data_7_), .Y(DP_OP_26J5_124_4249_n131) );
  INVX1_HVT U112 ( .A(DP_OP_26J5_124_4249_n198), .Y(DP_OP_26J5_124_4249_n196)
         );
  OR2X1_HVT U113 ( .A1(n66), .A2(ori_data_17_), .Y(n70) );
  AO21X1_HVT U114 ( .A1(DP_OP_26J5_124_4249_n80), .A2(DP_OP_26J5_124_4249_n29), 
        .A3(DP_OP_26J5_124_4249_n30), .Y(n71) );
  AO21X1_HVT U115 ( .A1(DP_OP_26J5_124_4249_n246), .A2(
        DP_OP_26J5_124_4249_n178), .A3(DP_OP_26J5_124_4249_n179), .Y(n72) );
  OR2X1_HVT U116 ( .A1(n67), .A2(ori_data_18_), .Y(n73) );
  AND2X1_HVT U117 ( .A1(n81), .A2(mode[1]), .Y(n96) );
  INVX1_HVT U118 ( .A(N43), .Y(n109) );
  INVX1_HVT U119 ( .A(N113), .Y(n107) );
  OR4X1_HVT U120 ( .A1(N50), .A2(N46), .A3(n84), .A4(N51), .Y(n85) );
  OR4X1_HVT U121 ( .A1(N43), .A2(N44), .A3(N47), .A4(N45), .Y(n83) );
  OR3X1_HVT U122 ( .A1(N114), .A2(N113), .A3(N116), .Y(n75) );
  OR3X1_HVT U123 ( .A1(N118), .A2(N115), .A3(N119), .Y(n74) );
  OR3X1_HVT U124 ( .A1(n75), .A2(n74), .A3(N117), .Y(n76) );
  OR3X1_HVT U125 ( .A1(N120), .A2(n76), .A3(N121), .Y(n77) );
  OR3X1_HVT U126 ( .A1(N122), .A2(n77), .A3(N123), .Y(n78) );
  OR3X1_HVT U127 ( .A1(N124), .A2(n78), .A3(N125), .Y(n79) );
  OR3X1_HVT U128 ( .A1(N126), .A2(n79), .A3(N127), .Y(n80) );
  NOR4X1_HVT U129 ( .A1(N129), .A2(N128), .A3(n80), .A4(N130), .Y(n82) );
  OA21X1_HVT U130 ( .A1(N131), .A2(n82), .A3(n103), .Y(n1140) );
  OR3X1_HVT U131 ( .A1(N49), .A2(N48), .A3(n83), .Y(n84) );
  OR3X1_HVT U132 ( .A1(N52), .A2(n85), .A3(N53), .Y(n86) );
  OR3X1_HVT U133 ( .A1(N54), .A2(n86), .A3(N55), .Y(n87) );
  OR3X1_HVT U134 ( .A1(N56), .A2(n87), .A3(N57), .Y(n88) );
  NOR4X1_HVT U135 ( .A1(N59), .A2(N58), .A3(n88), .A4(N60), .Y(n89) );
  OA21X1_HVT U136 ( .A1(N61), .A2(n89), .A3(n96), .Y(n112) );
  AND4X1_HVT U137 ( .A1(N47), .A2(N45), .A3(N44), .A4(N43), .Y(n90) );
  AND3X1_HVT U138 ( .A1(N48), .A2(N49), .A3(n90), .Y(n91) );
  AND4X1_HVT U139 ( .A1(N51), .A2(n91), .A3(N50), .A4(N46), .Y(n92) );
  AND4X1_HVT U140 ( .A1(N54), .A2(N53), .A3(N52), .A4(n92), .Y(n93) );
  AND4X1_HVT U141 ( .A1(N57), .A2(N56), .A3(N55), .A4(n93), .Y(n94) );
  NAND4X0_HVT U142 ( .A1(N60), .A2(N59), .A3(N58), .A4(n94), .Y(n95) );
  NAND2X0_HVT U143 ( .A1(n95), .A2(N61), .Y(n110) );
  AND2X1_HVT U144 ( .A1(n110), .A2(n96), .Y(n104) );
  AND3X1_HVT U145 ( .A1(N116), .A2(N114), .A3(N113), .Y(n97) );
  AND4X1_HVT U146 ( .A1(n97), .A2(N119), .A3(N118), .A4(N115), .Y(n98) );
  AND4X1_HVT U147 ( .A1(N121), .A2(N120), .A3(N117), .A4(n98), .Y(n99) );
  AND4X1_HVT U148 ( .A1(N124), .A2(N123), .A3(N122), .A4(n99), .Y(n100) );
  AND4X1_HVT U149 ( .A1(N127), .A2(N126), .A3(N125), .A4(n100), .Y(n101) );
  NAND4X0_HVT U150 ( .A1(N130), .A2(N129), .A3(N128), .A4(n101), .Y(n102) );
  NAND2X0_HVT U151 ( .A1(n102), .A2(N131), .Y(n108) );
  AND2X1_HVT U152 ( .A1(n108), .A2(n103), .Y(n105) );
  NAND2X0_HVT U153 ( .A1(n108), .A2(n107), .Y(n1130) );
  NAND2X0_HVT U154 ( .A1(n110), .A2(n109), .Y(n111) );
  AO22X1_HVT U155 ( .A1(n1140), .A2(n1130), .A3(n112), .A4(n111), .Y(
        n_quantized_data[7]) );
endmodule


module conv_top ( clk, srstn, conv_start, sram_rdata_a0, sram_rdata_a1, 
        sram_rdata_a2, sram_rdata_a3, sram_rdata_a4, sram_rdata_a5, 
        sram_rdata_a6, sram_rdata_a7, sram_rdata_a8, sram_rdata_b0, 
        sram_rdata_b1, sram_rdata_b2, sram_rdata_b3, sram_rdata_b4, 
        sram_rdata_b5, sram_rdata_b6, sram_rdata_b7, sram_rdata_b8, 
        sram_rdata_weight, sram_raddr_weight, sram_raddr_a0, sram_raddr_a1, 
        sram_raddr_a2, sram_raddr_a3, sram_raddr_a4, sram_raddr_a5, 
        sram_raddr_a6, sram_raddr_a7, sram_raddr_a8, sram_write_enable_b0, 
        sram_write_enable_b1, sram_write_enable_b2, sram_write_enable_b3, 
        sram_write_enable_b4, sram_write_enable_b5, sram_write_enable_b6, 
        sram_write_enable_b7, sram_write_enable_b8, sram_bytemask_b, 
        sram_waddr_b, sram_wdata_b, sram_raddr_b0, sram_raddr_b1, 
        sram_raddr_b2, sram_raddr_b3, sram_raddr_b4, sram_raddr_b5, 
        sram_raddr_b6, sram_raddr_b7, sram_raddr_b8, sram_write_enable_c0, 
        sram_write_enable_c1, sram_write_enable_c2, sram_write_enable_c3, 
        sram_write_enable_c4, sram_bytemask_c, sram_waddr_c, sram_wdata_c, 
        sram_write_enable_d0, sram_write_enable_d1, sram_write_enable_d2, 
        sram_write_enable_d3, sram_write_enable_d4, sram_bytemask_d, 
        sram_waddr_d, sram_wdata_d, conv1_done, conv_done, mem_sel );
  input [31:0] sram_rdata_a0;
  input [31:0] sram_rdata_a1;
  input [31:0] sram_rdata_a2;
  input [31:0] sram_rdata_a3;
  input [31:0] sram_rdata_a4;
  input [31:0] sram_rdata_a5;
  input [31:0] sram_rdata_a6;
  input [31:0] sram_rdata_a7;
  input [31:0] sram_rdata_a8;
  input [31:0] sram_rdata_b0;
  input [31:0] sram_rdata_b1;
  input [31:0] sram_rdata_b2;
  input [31:0] sram_rdata_b3;
  input [31:0] sram_rdata_b4;
  input [31:0] sram_rdata_b5;
  input [31:0] sram_rdata_b6;
  input [31:0] sram_rdata_b7;
  input [31:0] sram_rdata_b8;
  input [99:0] sram_rdata_weight;
  output [16:0] sram_raddr_weight;
  output [9:0] sram_raddr_a0;
  output [9:0] sram_raddr_a1;
  output [9:0] sram_raddr_a2;
  output [9:0] sram_raddr_a3;
  output [9:0] sram_raddr_a4;
  output [9:0] sram_raddr_a5;
  output [9:0] sram_raddr_a6;
  output [9:0] sram_raddr_a7;
  output [9:0] sram_raddr_a8;
  output [3:0] sram_bytemask_b;
  output [9:0] sram_waddr_b;
  output [7:0] sram_wdata_b;
  output [9:0] sram_raddr_b0;
  output [9:0] sram_raddr_b1;
  output [9:0] sram_raddr_b2;
  output [9:0] sram_raddr_b3;
  output [9:0] sram_raddr_b4;
  output [9:0] sram_raddr_b5;
  output [9:0] sram_raddr_b6;
  output [9:0] sram_raddr_b7;
  output [9:0] sram_raddr_b8;
  output [3:0] sram_bytemask_c;
  output [9:0] sram_waddr_c;
  output [7:0] sram_wdata_c;
  output [3:0] sram_bytemask_d;
  output [9:0] sram_waddr_d;
  output [7:0] sram_wdata_d;
  input clk, srstn, conv_start;
  output sram_write_enable_b0, sram_write_enable_b1, sram_write_enable_b2,
         sram_write_enable_b3, sram_write_enable_b4, sram_write_enable_b5,
         sram_write_enable_b6, sram_write_enable_b7, sram_write_enable_b8,
         sram_write_enable_c0, sram_write_enable_c1, sram_write_enable_c2,
         sram_write_enable_c3, sram_write_enable_c4, sram_write_enable_d0,
         sram_write_enable_d1, sram_write_enable_d2, sram_write_enable_d3,
         sram_write_enable_d4, conv1_done, conv_done, mem_sel;
  wire   load_conv1_bias_enable, conv1_bias_set_16_, conv1_bias_set_15_,
         conv1_bias_set_14_, conv1_bias_set_13_, conv1_bias_set_12_,
         conv1_bias_set_11_, conv1_bias_set_10_, conv1_bias_set_9_,
         conv1_bias_set_8_, conv1_bias_set_7_, conv1_bias_set_6_,
         conv1_bias_set_5_, conv1_bias_set_4_, conv1_bias_set_3_,
         conv1_bias_set_2_, conv1_bias_set_1_, conv1_bias_set_0_, set_7_,
         set_6_, set_5_, set_4_, set_3_, set_2_, set_1_, set_0_,
         load_conv2_bias0_enable, load_conv2_bias1_enable, data_out_31_,
         data_out_30_, data_out_29_, data_out_28_, data_out_27_, data_out_26_,
         data_out_25_, data_out_24_, data_out_23_, data_out_22_, data_out_21_,
         data_out_20_, data_out_19_, data_out_18_, data_out_17_, data_out_16_,
         data_out_15_, data_out_14_, data_out_13_, data_out_12_, data_out_11_,
         data_out_10_, data_out_9_, data_out_8_, data_out_7_, data_out_6_,
         data_out_5_, data_out_4_, data_out_3_, data_out_2_, data_out_1_,
         data_out_0_, n1;
  wire   [1:0] mode;
  wire   [3:0] box_sel;
  wire   [4:0] channel;
  wire   [99:0] conv1_weight;
  wire   [99:0] weight;
  wire   [287:0] src_window;
  wire   [3:0] bias_data;

  fsm fsm ( .clk(clk), .srstn(n1), .conv_start(conv_start), .conv1_done(
        conv1_done), .conv_done(conv_done), .mode(mode), .mem_sel(mem_sel) );
  conv_control conv_control ( .clk(clk), .srstn(srstn), .mode(mode), .mem_sel(
        mem_sel), .conv1_done(conv1_done), .sram_raddr_weight(
        sram_raddr_weight), .box_sel(box_sel), .load_conv1_bias_enable(
        load_conv1_bias_enable), .conv1_bias_set({conv1_bias_set_16_, 
        conv1_bias_set_15_, conv1_bias_set_14_, conv1_bias_set_13_, 
        conv1_bias_set_12_, conv1_bias_set_11_, conv1_bias_set_10_, 
        conv1_bias_set_9_, conv1_bias_set_8_, conv1_bias_set_7_, 
        conv1_bias_set_6_, conv1_bias_set_5_, conv1_bias_set_4_, 
        conv1_bias_set_3_, conv1_bias_set_2_, conv1_bias_set_1_, 
        conv1_bias_set_0_}), .sram_raddr_a0(sram_raddr_a0), .sram_raddr_a1(
        sram_raddr_a1), .sram_raddr_a2(sram_raddr_a2), .sram_raddr_a3(
        sram_raddr_a3), .sram_raddr_a4(sram_raddr_a4), .sram_raddr_a5(
        sram_raddr_a5), .sram_raddr_a6(sram_raddr_a6), .sram_raddr_a7(
        sram_raddr_a7), .sram_raddr_a8(sram_raddr_a8), .sram_write_enable_b0(
        sram_write_enable_b0), .sram_write_enable_b1(sram_write_enable_b1), 
        .sram_write_enable_b2(sram_write_enable_b2), .sram_write_enable_b3(
        sram_write_enable_b3), .sram_write_enable_b4(sram_write_enable_b4), 
        .sram_write_enable_b5(sram_write_enable_b5), .sram_write_enable_b6(
        sram_write_enable_b6), .sram_write_enable_b7(sram_write_enable_b7), 
        .sram_write_enable_b8(sram_write_enable_b8), .sram_bytemask_b(
        sram_bytemask_b), .sram_waddr_b(sram_waddr_b), .conv_done(conv_done), 
        .channel(channel), .set({set_7_, set_6_, set_5_, set_4_, set_3_, 
        set_2_, set_1_, set_0_}), .load_conv2_bias0_enable(
        load_conv2_bias0_enable), .load_conv2_bias1_enable(
        load_conv2_bias1_enable), .sram_raddr_b0(sram_raddr_b0), 
        .sram_raddr_b1(sram_raddr_b1), .sram_raddr_b2(sram_raddr_b2), 
        .sram_raddr_b3(sram_raddr_b3), .sram_raddr_b4(sram_raddr_b4), 
        .sram_raddr_b5(sram_raddr_b5), .sram_raddr_b6(sram_raddr_b6), 
        .sram_raddr_b7(sram_raddr_b7), .sram_raddr_b8(sram_raddr_b8), 
        .sram_write_enable_c0(sram_write_enable_c0), .sram_write_enable_c1(
        sram_write_enable_c1), .sram_write_enable_c2(sram_write_enable_c2), 
        .sram_write_enable_c3(sram_write_enable_c3), .sram_write_enable_c4(
        sram_write_enable_c4), .sram_bytemask_c(sram_bytemask_c), 
        .sram_waddr_c(sram_waddr_c), .sram_write_enable_d0(
        sram_write_enable_d0), .sram_write_enable_d1(sram_write_enable_d1), 
        .sram_write_enable_d2(sram_write_enable_d2), .sram_write_enable_d3(
        sram_write_enable_d3), .sram_write_enable_d4(sram_write_enable_d4), 
        .sram_bytemask_d(sram_bytemask_d), .sram_waddr_d(sram_waddr_d) );
  data_reg data_reg ( .clk(clk), .srstn(n1), .mode(mode), .box_sel(box_sel), 
        .sram_rdata_a0(sram_rdata_a0), .sram_rdata_a1(sram_rdata_a1), 
        .sram_rdata_a2(sram_rdata_a2), .sram_rdata_a3(sram_rdata_a3), 
        .sram_rdata_a4(sram_rdata_a4), .sram_rdata_a5(sram_rdata_a5), 
        .sram_rdata_a6(sram_rdata_a6), .sram_rdata_a7(sram_rdata_a7), 
        .sram_rdata_a8(sram_rdata_a8), .sram_rdata_b0(sram_rdata_b0), 
        .sram_rdata_b1(sram_rdata_b1), .sram_rdata_b2(sram_rdata_b2), 
        .sram_rdata_b3(sram_rdata_b3), .sram_rdata_b4(sram_rdata_b4), 
        .sram_rdata_b5(sram_rdata_b5), .sram_rdata_b6(sram_rdata_b6), 
        .sram_rdata_b7(sram_rdata_b7), .sram_rdata_b8(sram_rdata_b8), 
        .sram_rdata_weight(sram_rdata_weight), .conv1_weight(conv1_weight), 
        .weight(weight), .src_window(src_window) );
  bias_sel bias_sel ( .clk(clk), .srstn(srstn), .mode(mode), 
        .load_conv1_bias_enable(load_conv1_bias_enable), 
        .load_conv2_bias0_enable(load_conv2_bias0_enable), 
        .load_conv2_bias1_enable(load_conv2_bias1_enable), .sram_rdata_weight(
        sram_rdata_weight), .bias_data(bias_data), .conv1_bias_set_5_(
        conv1_bias_set_5_), .conv1_bias_set_4_(conv1_bias_set_4_), 
        .conv1_bias_set_3_(conv1_bias_set_3_), .conv1_bias_set_2_(
        conv1_bias_set_2_), .conv1_bias_set_1_(conv1_bias_set_1_), 
        .conv1_bias_set_0_(conv1_bias_set_0_), .set_5_(set_5_), .set_4_(set_4_), .set_3_(set_3_), .set_2_(set_2_), .set_1_(set_1_), .set_0_(set_0_) );
  multiply_compare multiply_compare ( .clk(clk), .srstn(n1), .mode(mode), 
        .channel(channel), .conv1_sram_rdata_weight(conv1_weight), 
        .conv2_sram_rdata_weight(weight), .src_window(src_window), .data_out({
        data_out_31_, data_out_30_, data_out_29_, data_out_28_, data_out_27_, 
        data_out_26_, data_out_25_, data_out_24_, data_out_23_, data_out_22_, 
        data_out_21_, data_out_20_, data_out_19_, data_out_18_, data_out_17_, 
        data_out_16_, data_out_15_, data_out_14_, data_out_13_, data_out_12_, 
        data_out_11_, data_out_10_, data_out_9_, data_out_8_, data_out_7_, 
        data_out_6_, data_out_5_, data_out_4_, data_out_3_, data_out_2_, 
        data_out_1_, data_out_0_}) );
  quantize quantize ( .clk(clk), .srstn(n1), .bias_data(bias_data), .mode(mode), .quantized_data(sram_wdata_c), .ori_data_31_(data_out_31_), .ori_data_30_(
        data_out_30_), .ori_data_29_(data_out_29_), .ori_data_28_(data_out_28_), .ori_data_27_(data_out_27_), .ori_data_26_(data_out_26_), .ori_data_25_(
        data_out_25_), .ori_data_24_(data_out_24_), .ori_data_23_(data_out_23_), .ori_data_22_(data_out_22_), .ori_data_21_(data_out_21_), .ori_data_20_(
        data_out_20_), .ori_data_19_(data_out_19_), .ori_data_18_(data_out_18_), .ori_data_17_(data_out_17_), .ori_data_16_(data_out_16_), .ori_data_15_(
        data_out_15_), .ori_data_14_(data_out_14_), .ori_data_13_(data_out_13_), .ori_data_12_(data_out_12_), .ori_data_11_(data_out_11_), .ori_data_10_(
        data_out_10_), .ori_data_9_(data_out_9_), .ori_data_8_(data_out_8_), 
        .ori_data_7_(data_out_7_), .ori_data_6_(data_out_6_), .ori_data_5_(
        data_out_5_) );
  NBUFFX2_HVT U1 ( .A(srstn), .Y(n1) );
  DELLN1X2_HVT U2 ( .A(sram_wdata_c[0]), .Y(sram_wdata_d[0]) );
  DELLN1X2_HVT U3 ( .A(sram_wdata_c[1]), .Y(sram_wdata_d[1]) );
  DELLN1X2_HVT U4 ( .A(sram_wdata_c[2]), .Y(sram_wdata_d[2]) );
  DELLN1X2_HVT U5 ( .A(sram_wdata_c[3]), .Y(sram_wdata_d[3]) );
  DELLN1X2_HVT U6 ( .A(sram_wdata_c[4]), .Y(sram_wdata_d[4]) );
  DELLN1X2_HVT U7 ( .A(sram_wdata_c[5]), .Y(sram_wdata_d[5]) );
  DELLN1X2_HVT U8 ( .A(sram_wdata_c[6]), .Y(sram_wdata_d[6]) );
  DELLN1X2_HVT U9 ( .A(sram_wdata_c[7]), .Y(sram_wdata_d[7]) );
  NBUFFX2_HVT U10 ( .A(sram_wdata_c[7]), .Y(sram_wdata_b[7]) );
  NBUFFX2_HVT U11 ( .A(sram_wdata_c[6]), .Y(sram_wdata_b[6]) );
  NBUFFX2_HVT U12 ( .A(sram_wdata_c[5]), .Y(sram_wdata_b[5]) );
  NBUFFX2_HVT U13 ( .A(sram_wdata_c[4]), .Y(sram_wdata_b[4]) );
  NBUFFX2_HVT U14 ( .A(sram_wdata_c[3]), .Y(sram_wdata_b[3]) );
  NBUFFX2_HVT U15 ( .A(sram_wdata_c[2]), .Y(sram_wdata_b[2]) );
  NBUFFX2_HVT U16 ( .A(sram_wdata_c[1]), .Y(sram_wdata_b[1]) );
  NBUFFX2_HVT U17 ( .A(sram_wdata_c[0]), .Y(sram_wdata_b[0]) );
endmodule

