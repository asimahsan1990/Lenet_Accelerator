/**
 * Editor : 
 * File : conv_top.v
 */
module conv_top(

);


endmodule