
module fsm ( clk, srstn, conv_start, conv1_done, conv_done, fc_done, mode, 
        mem_sel );
  output [1:0] mode;
  input clk, srstn, conv_start, conv1_done, conv_done, fc_done;
  output mem_sel;
  wire   n_mem_sel, done_control, n2, n6, n8, n3, n5, n7, n9, n10, n11;
  wire   [1:0] n_mode;

  DFFSSRX1_HVT mode_reg_0_ ( .D(1'b0), .SETB(n8), .RSTB(n_mode[0]), .CLK(clk), 
        .Q(mode[0]), .QN(n6) );
  DFFSSRX1_HVT mode_reg_1_ ( .D(1'b0), .SETB(n8), .RSTB(n_mode[1]), .CLK(clk), 
        .Q(mode[1]), .QN(n3) );
  DFFSSRX1_HVT done_control_reg ( .D(done_control), .SETB(n2), .RSTB(srstn), 
        .CLK(clk), .Q(done_control), .QN(n5) );
  DFFSSRX1_HVT mem_sel_reg ( .D(n_mem_sel), .SETB(srstn), .RSTB(1'b1), .CLK(
        clk), .Q(mem_sel) );
  OA222X1_HVT U4 ( .A1(n10), .A2(n3), .A3(n10), .A4(mode[0]), .A5(n10), .A6(
        conv1_done), .Y(n_mode[1]) );
  INVX0_HVT U5 ( .A(conv_done), .Y(n2) );
  INVX1_HVT U6 ( .A(srstn), .Y(n8) );
  INVX1_HVT U7 ( .A(conv1_done), .Y(n7) );
  AND2X1_HVT U8 ( .A1(mode[1]), .A2(n6), .Y(n10) );
  MUX21X1_HVT U9 ( .A1(n7), .A2(conv_start), .S0(n6), .Y(n9) );
  AO22X1_HVT U10 ( .A1(n10), .A2(conv_done), .A3(n9), .A4(n3), .Y(n_mode[0])
         );
  AO22X1_HVT U11 ( .A1(done_control), .A2(fc_done), .A3(n5), .A4(conv_done), 
        .Y(n11) );
  HADDX1_HVT U12 ( .A0(mem_sel), .B0(n11), .SO(n_mem_sel) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_0 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n1;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n1), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n1) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_26 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_25 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_24 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_23 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_22 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_21 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_20 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_19 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_18 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_17 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_16 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_15 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_14 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_13 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_12 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_11 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_10 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_9 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_8 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_7 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_6 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_5 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_4 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_3 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_2 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_1 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22628, n2;

  AND2X1_HVT main_gate ( .A1(net22628), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22628) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module conv_control ( clk, srstn, mode, mem_sel, conv1_done, sram_raddr_weight, 
        box_sel, load_conv1_bias_enable, conv1_bias_set, sram_raddr_a0, 
        sram_raddr_a1, sram_raddr_a2, sram_raddr_a3, sram_raddr_a4, 
        sram_raddr_a5, sram_raddr_a6, sram_raddr_a7, sram_raddr_a8, 
        sram_write_enable_b0, sram_write_enable_b1, sram_write_enable_b2, 
        sram_write_enable_b3, sram_write_enable_b4, sram_write_enable_b5, 
        sram_write_enable_b6, sram_write_enable_b7, sram_write_enable_b8, 
        sram_bytemask_b, sram_waddr_b, conv_done, channel, set, 
        load_conv2_bias0_enable, load_conv2_bias1_enable, sram_raddr_b0, 
        sram_raddr_b1, sram_raddr_b2, sram_raddr_b3, sram_raddr_b4, 
        sram_raddr_b5, sram_raddr_b6, sram_raddr_b7, sram_raddr_b8, 
        sram_write_enable_c0, sram_write_enable_c1, sram_write_enable_c2, 
        sram_write_enable_c3, sram_write_enable_c4, sram_bytemask_c, 
        sram_waddr_c, sram_write_enable_d0, sram_write_enable_d1, 
        sram_write_enable_d2, sram_write_enable_d3, sram_write_enable_d4, 
        sram_bytemask_d, sram_waddr_d );
  input [1:0] mode;
  output [16:0] sram_raddr_weight;
  output [3:0] box_sel;
  output [16:0] conv1_bias_set;
  output [9:0] sram_raddr_a0;
  output [9:0] sram_raddr_a1;
  output [9:0] sram_raddr_a2;
  output [9:0] sram_raddr_a3;
  output [9:0] sram_raddr_a4;
  output [9:0] sram_raddr_a5;
  output [9:0] sram_raddr_a6;
  output [9:0] sram_raddr_a7;
  output [9:0] sram_raddr_a8;
  output [3:0] sram_bytemask_b;
  output [9:0] sram_waddr_b;
  output [4:0] channel;
  output [7:0] set;
  output [9:0] sram_raddr_b0;
  output [9:0] sram_raddr_b1;
  output [9:0] sram_raddr_b2;
  output [9:0] sram_raddr_b3;
  output [9:0] sram_raddr_b4;
  output [9:0] sram_raddr_b5;
  output [9:0] sram_raddr_b6;
  output [9:0] sram_raddr_b7;
  output [9:0] sram_raddr_b8;
  output [3:0] sram_bytemask_c;
  output [9:0] sram_waddr_c;
  output [3:0] sram_bytemask_d;
  output [9:0] sram_waddr_d;
  input clk, srstn, mem_sel;
  output conv1_done, load_conv1_bias_enable, sram_write_enable_b0,
         sram_write_enable_b1, sram_write_enable_b2, sram_write_enable_b3,
         sram_write_enable_b4, sram_write_enable_b5, sram_write_enable_b6,
         sram_write_enable_b7, sram_write_enable_b8, conv_done,
         load_conv2_bias0_enable, load_conv2_bias1_enable,
         sram_write_enable_c0, sram_write_enable_c1, sram_write_enable_c2,
         sram_write_enable_c3, sram_write_enable_c4, sram_write_enable_d0,
         sram_write_enable_d1, sram_write_enable_d2, sram_write_enable_d3,
         sram_write_enable_d4;
  wire   n_conv1_done, n_conv_done, conv1_weight_done, conv2_weight_done,
         delay3_write_enable, load_data_enable, n_conv1_weight_done,
         n_write_enable, write_enable, delay_write_enable, delay2_write_enable,
         n_load_data_enable, n_box_sel_1_, n_addr_row_sel_cnt_0_,
         n_sram_write_enable_b0, n_sram_write_enable_b1,
         n_sram_write_enable_b2, n_sram_write_enable_b3,
         n_sram_write_enable_b4, n_sram_write_enable_b5,
         n_sram_write_enable_b6, n_sram_write_enable_b7,
         n_sram_write_enable_b8, n_sram_write_enable_c0,
         n_sram_write_enable_c1, n_sram_write_enable_c2,
         n_sram_write_enable_c3, n_sram_write_enable_c4,
         n_sram_write_enable_d0, n_sram_write_enable_d1,
         n_sram_write_enable_d2, n_sram_write_enable_d3,
         n_sram_write_enable_d4, N2914, net22462, net22639, net22644, net22649,
         net22654, net22655, net22658, net22663, net22692, net22699, net22706,
         net22713, net22720, net22727, net22734, net22748, net22755, net22758,
         net22776, net22783, net22790, net22797, net22811, net22818, net22825,
         net22839, net22853, net22856, net22861, net22864, net22867, net22870,
         net22873, net22876, net22879, net22882, net22885, net22888, net22891,
         net22894, net22899, net22901, net22902, net22903, net22904, net22905,
         net22906, net22907, net22908, net22909, net22910, net22913, net22917,
         net22918, net22919, net22920, net22921, net22922, net22923, net22924,
         net22925, net22926, net22929, net22933, net22934, net22935, net22936,
         net22937, net22938, net22941, net22944, net22946, net22947, net22948,
         net22949, net22950, net22953, net23434, net23879, net23893, net24316,
         net24761, net25206, net25220, net25643, net26089, net26535, net26550,
         net26973, net27507, net28022, net28537, net29052, net29567, net30082,
         net30597, net31112, net31204, net31627, n368, n369, n371, n392, n1020,
         n1021, n1022, n1023, n1024, n1027, n1051, n1052, n1053, n1061, n1062,
         n1063, n1655, n1662, n1667, n1, n2, n3, n5, n6, n7, n8, n10, n11, n12,
         n13, n14, n15, n17, n18, n20, n21, n23, n24, n25, n26, n28, n29, n31,
         n32, n33, n34, n35, n37, n38, n39, n40, n41, n42, n43, n47, n48, n49,
         n50, n51, n53, n54, n55, n57, n58, n59, n60, n62, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n77, n78, n79, n80, n81, n82, n83,
         n86, n89, n90, n91, n92, n93, n94, n95, n96, n98, n101, n103, n104,
         n105, n106, n107, n109, n111, n112, n113, n115, n117, n119, n120,
         n122, n124, n126, n128, n129, n130, n131, n132, n134, n135, n136,
         n138, n141, n142, n143, n144, n145, n146, n149, n151, n152, n155,
         n157, n158, n159, n160, n162, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n370, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1025, n1026,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1656, n1657, n1658, n1659, n1660, n1661, n1663, n1664, n1665,
         n1666, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003;
  wire   [7:0] conv1_weight_cnt;
  wire   [7:0] conv2_weight_cnt;
  wire   [3:0] state;
  wire   [3:0] n_state;
  wire   [4:0] channel_cnt;
  wire   [1:0] data_sel_col;
  wire   [1:0] data_sel_row;
  wire   [9:0] delay1_sram_waddr_b;
  wire   [3:0] write_row_conv1;
  wire   [1:0] write_col_conv1;
  wire   [4:0] delay3_addr_change;
  wire   [2:0] delay3_state;
  wire   [3:0] n_row;
  wire   [7:0] n_weight_cnt;
  wire   [7:0] weight_cnt;
  wire   [7:0] delay_set;
  wire   [1:0] n_addr_col_sel_cnt;
  wire   [1:0] addr_col_sel_cnt;
  wire   [1:0] addr_row_sel_cnt;
  wire   [3:0] n_sram_bytemask_b;
  wire   [3:0] row;
  wire   [3:0] col;
  wire   [3:0] row_delay;
  wire   [3:0] col_delay;
  wire   [3:0] write_row;
  wire   [3:0] write_col;
  wire   [3:0] row_enable;
  wire   [3:0] col_enable;
  wire   [9:0] delay1_sram_waddr_c;
  wire   [9:0] delay1_sram_waddr_d;
  wire   [3:0] n_sram_bytemask_c;
  wire   [3:0] n_sram_bytemask_d;
  wire   [4:0] addr_change;
  wire   [4:0] delay_addr_change;
  wire   [4:0] delay2_addr_change;
  wire   [4:0] delay_channel;
  wire   [4:0] delay2_channel;
  wire   [3:0] delay1_state;
  wire   [3:0] delay2_state;
  wire   [9:0] n_sram_raddr_a0;
  wire   [9:0] n_sram_raddr_a1;
  wire   [9:0] n_sram_raddr_a2;
  wire   [9:0] n_sram_raddr_a3;
  wire   [9:0] n_sram_raddr_a4;
  wire   [9:0] n_sram_raddr_a5;
  wire   [9:0] n_sram_raddr_a6;
  wire   [9:0] n_sram_raddr_a7;
  wire   [9:0] n_sram_raddr_a8;
  wire   [9:0] n_sram_raddr_b0;
  wire   [9:0] n_sram_raddr_b1;
  wire   [9:0] n_sram_raddr_b2;
  wire   [9:0] n_sram_raddr_b3;
  wire   [9:0] n_sram_raddr_b4;
  wire   [9:0] n_sram_raddr_b5;
  wire   [9:0] n_sram_raddr_b6;
  wire   [9:0] n_sram_raddr_b7;
  wire   [9:0] n_sram_raddr_b8;

  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_0 clk_gate_col_reg ( .CLK(clk), 
        .EN(net22462), .ENCLK(net22658) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_26 clk_gate_weight_cnt_reg ( 
        .CLK(clk), .EN(net22462), .ENCLK(net22663) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_25 clk_gate_sram_raddr_weight_reg ( 
        .CLK(clk), .EN(net22776), .ENCLK(net22758) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_24 clk_gate_sram_raddr_weight_reg_0 ( 
        .CLK(clk), .EN(net22776), .ENCLK(net22856) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_23 clk_gate_delay1_sram_waddr_b_reg ( 
        .CLK(clk), .EN(net22861), .ENCLK(net22894) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_22 clk_gate_delay1_sram_waddr_c_reg ( 
        .CLK(clk), .EN(net22899), .ENCLK(net22913) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_21 clk_gate_delay1_sram_waddr_d_reg ( 
        .CLK(clk), .EN(net22899), .ENCLK(net22929) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_20 clk_gate_channel_cnt_reg ( 
        .CLK(clk), .EN(net22933), .ENCLK(net22941) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_19 clk_gate_addr_change_reg ( 
        .CLK(clk), .EN(net22944), .ENCLK(net22953) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_18 clk_gate_sram_raddr_a7_reg ( 
        .CLK(clk), .EN(net23893), .ENCLK(net23434) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_17 clk_gate_sram_raddr_a1_reg ( 
        .CLK(clk), .EN(net23893), .ENCLK(net23879) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_16 clk_gate_sram_raddr_a4_reg ( 
        .CLK(clk), .EN(net23893), .ENCLK(net24316) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_15 clk_gate_sram_raddr_a8_reg ( 
        .CLK(clk), .EN(net25220), .ENCLK(net24761) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_14 clk_gate_sram_raddr_a2_reg ( 
        .CLK(clk), .EN(net25220), .ENCLK(net25206) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_13 clk_gate_sram_raddr_a5_reg ( 
        .CLK(clk), .EN(net25220), .ENCLK(net25643) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_12 clk_gate_sram_raddr_a0_reg ( 
        .CLK(clk), .EN(net26550), .ENCLK(net26089) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_11 clk_gate_sram_raddr_a3_reg ( 
        .CLK(clk), .EN(net26550), .ENCLK(net26535) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_10 clk_gate_sram_raddr_a6_reg ( 
        .CLK(clk), .EN(net26550), .ENCLK(net26973) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_9 clk_gate_sram_raddr_b7_reg ( 
        .CLK(clk), .EN(net31204), .ENCLK(net27507) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_8 clk_gate_sram_raddr_b8_reg ( 
        .CLK(clk), .EN(net31204), .ENCLK(net28022) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_7 clk_gate_sram_raddr_b0_reg ( 
        .CLK(clk), .EN(net31204), .ENCLK(net28537) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_6 clk_gate_sram_raddr_b1_reg ( 
        .CLK(clk), .EN(net31204), .ENCLK(net29052) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_5 clk_gate_sram_raddr_b2_reg ( 
        .CLK(clk), .EN(net31204), .ENCLK(net29567) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_4 clk_gate_sram_raddr_b3_reg ( 
        .CLK(clk), .EN(net31204), .ENCLK(net30082) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_3 clk_gate_sram_raddr_b4_reg ( 
        .CLK(clk), .EN(net31204), .ENCLK(net30597) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_2 clk_gate_sram_raddr_b5_reg ( 
        .CLK(clk), .EN(net31204), .ENCLK(net31112) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_1 clk_gate_sram_raddr_b6_reg ( 
        .CLK(clk), .EN(net31204), .ENCLK(net31627) );
  DFFSSRX1_HVT channel_cnt_reg_0_ ( .D(1'b0), .SETB(n198), .RSTB(net22938), 
        .CLK(net22941), .Q(channel_cnt[0]) );
  DFFSSRX1_HVT state_reg_0_ ( .D(1'b0), .SETB(n193), .RSTB(n_state[0]), .CLK(
        clk), .Q(state[0]), .QN(n253) );
  DFFSSRX1_HVT weight_cnt_reg_0_ ( .D(1'b0), .SETB(n201), .RSTB(
        n_weight_cnt[0]), .CLK(net22663), .Q(weight_cnt[0]), .QN(n308) );
  DFFSSRX1_HVT delay_set_reg_0_ ( .D(1'b0), .SETB(n195), .RSTB(weight_cnt[0]), 
        .CLK(clk), .Q(delay_set[0]) );
  DFFSSRX1_HVT set_reg_0_ ( .D(1'b0), .SETB(n212), .RSTB(delay_set[0]), .CLK(
        clk), .Q(set[0]) );
  DFFSSRX1_HVT conv2_weight_cnt_reg_0_ ( .D(1'b0), .SETB(n210), .RSTB(set[0]), 
        .CLK(clk), .Q(conv2_weight_cnt[0]) );
  DFFSSRX1_HVT conv1_weight_cnt_reg_0_ ( .D(1'b0), .SETB(n169), .RSTB(
        conv2_weight_cnt[0]), .CLK(clk), .Q(conv1_weight_cnt[0]) );
  DFFSSRX1_HVT conv_done_reg ( .D(1'b0), .SETB(n185), .RSTB(n_conv_done), 
        .CLK(clk), .Q(conv_done) );
  DFFSSRX1_HVT state_reg_1_ ( .D(1'b0), .SETB(n199), .RSTB(n_state[1]), .CLK(
        clk), .Q(state[1]), .QN(n240) );
  DFFSSRX1_HVT weight_cnt_reg_7_ ( .D(1'b0), .SETB(n194), .RSTB(
        n_weight_cnt[7]), .CLK(net22663), .Q(weight_cnt[7]), .QN(n461) );
  DFFSSRX1_HVT delay_set_reg_7_ ( .D(1'b0), .SETB(n202), .RSTB(weight_cnt[7]), 
        .CLK(clk), .Q(delay_set[7]) );
  DFFSSRX1_HVT set_reg_7_ ( .D(1'b0), .SETB(n196), .RSTB(delay_set[7]), .CLK(
        clk), .Q(set[7]) );
  DFFSSRX1_HVT conv2_weight_cnt_reg_7_ ( .D(1'b0), .SETB(n211), .RSTB(set[7]), 
        .CLK(clk), .Q(conv2_weight_cnt[7]) );
  DFFSSRX1_HVT conv1_weight_cnt_reg_7_ ( .D(1'b0), .SETB(n209), .RSTB(
        conv2_weight_cnt[7]), .CLK(clk), .Q(conv1_weight_cnt[7]) );
  DFFSSRX1_HVT weight_cnt_reg_6_ ( .D(1'b0), .SETB(n187), .RSTB(
        n_weight_cnt[6]), .CLK(net22663), .Q(weight_cnt[6]) );
  DFFSSRX1_HVT delay_set_reg_6_ ( .D(1'b0), .SETB(n184), .RSTB(weight_cnt[6]), 
        .CLK(clk), .Q(delay_set[6]) );
  DFFSSRX1_HVT set_reg_6_ ( .D(1'b0), .SETB(n177), .RSTB(delay_set[6]), .CLK(
        clk), .Q(set[6]) );
  DFFSSRX1_HVT conv2_weight_cnt_reg_6_ ( .D(1'b0), .SETB(n176), .RSTB(set[6]), 
        .CLK(clk), .Q(conv2_weight_cnt[6]) );
  DFFSSRX1_HVT conv1_weight_cnt_reg_6_ ( .D(1'b0), .SETB(n175), .RSTB(
        conv2_weight_cnt[6]), .CLK(clk), .Q(conv1_weight_cnt[6]) );
  DFFSSRX1_HVT weight_cnt_reg_5_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_weight_cnt[5]), .CLK(net22663), .Q(weight_cnt[5]), .QN(n453) );
  DFFSSRX1_HVT delay_set_reg_5_ ( .D(1'b0), .SETB(n212), .RSTB(weight_cnt[5]), 
        .CLK(clk), .Q(delay_set[5]) );
  DFFSSRX1_HVT set_reg_5_ ( .D(1'b0), .SETB(n210), .RSTB(delay_set[5]), .CLK(
        clk), .Q(set[5]) );
  DFFSSRX1_HVT conv2_weight_cnt_reg_5_ ( .D(1'b0), .SETB(n169), .RSTB(set[5]), 
        .CLK(clk), .Q(conv2_weight_cnt[5]) );
  DFFSSRX1_HVT conv1_weight_cnt_reg_5_ ( .D(1'b0), .SETB(n186), .RSTB(
        conv2_weight_cnt[5]), .CLK(clk), .Q(conv1_weight_cnt[5]) );
  DFFSSRX1_HVT weight_cnt_reg_4_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_weight_cnt[4]), .CLK(net22663), .Q(weight_cnt[4]) );
  DFFSSRX1_HVT delay_set_reg_4_ ( .D(1'b0), .SETB(n176), .RSTB(weight_cnt[4]), 
        .CLK(clk), .Q(delay_set[4]) );
  DFFSSRX1_HVT set_reg_4_ ( .D(1'b0), .SETB(n175), .RSTB(delay_set[4]), .CLK(
        clk), .Q(set[4]) );
  DFFSSRX1_HVT conv2_weight_cnt_reg_4_ ( .D(1'b0), .SETB(n174), .RSTB(set[4]), 
        .CLK(clk), .Q(conv2_weight_cnt[4]) );
  DFFSSRX1_HVT conv1_weight_cnt_reg_4_ ( .D(1'b0), .SETB(n211), .RSTB(
        conv2_weight_cnt[4]), .CLK(clk), .Q(conv1_weight_cnt[4]) );
  DFFSSRX1_HVT weight_cnt_reg_3_ ( .D(1'b0), .SETB(n209), .RSTB(
        n_weight_cnt[3]), .CLK(net22663), .Q(weight_cnt[3]), .QN(n439) );
  DFFSSRX1_HVT delay_set_reg_3_ ( .D(1'b0), .SETB(n169), .RSTB(weight_cnt[3]), 
        .CLK(clk), .Q(delay_set[3]) );
  DFFSSRX1_HVT set_reg_3_ ( .D(1'b0), .SETB(n185), .RSTB(delay_set[3]), .CLK(
        clk), .Q(set[3]) );
  DFFSSRX1_HVT conv2_weight_cnt_reg_3_ ( .D(1'b0), .SETB(n198), .RSTB(set[3]), 
        .CLK(clk), .Q(conv2_weight_cnt[3]) );
  DFFSSRX1_HVT conv1_weight_cnt_reg_3_ ( .D(1'b0), .SETB(n193), .RSTB(
        conv2_weight_cnt[3]), .CLK(clk), .Q(conv1_weight_cnt[3]) );
  DFFSSRX1_HVT weight_cnt_reg_2_ ( .D(1'b0), .SETB(n201), .RSTB(
        n_weight_cnt[2]), .CLK(net22663), .Q(weight_cnt[2]) );
  DFFSSRX1_HVT delay_set_reg_2_ ( .D(1'b0), .SETB(n195), .RSTB(weight_cnt[2]), 
        .CLK(clk), .Q(delay_set[2]) );
  DFFSSRX1_HVT set_reg_2_ ( .D(1'b0), .SETB(n212), .RSTB(delay_set[2]), .CLK(
        clk), .Q(set[2]) );
  DFFSSRX1_HVT conv2_weight_cnt_reg_2_ ( .D(1'b0), .SETB(n210), .RSTB(set[2]), 
        .CLK(clk), .Q(conv2_weight_cnt[2]) );
  DFFSSRX1_HVT conv1_weight_cnt_reg_2_ ( .D(1'b0), .SETB(n187), .RSTB(
        conv2_weight_cnt[2]), .CLK(clk), .Q(conv1_weight_cnt[2]) );
  DFFSSRX1_HVT weight_cnt_reg_1_ ( .D(1'b0), .SETB(n184), .RSTB(
        n_weight_cnt[1]), .CLK(net22663), .Q(weight_cnt[1]), .QN(n444) );
  DFFSSRX1_HVT delay_set_reg_1_ ( .D(1'b0), .SETB(n199), .RSTB(weight_cnt[1]), 
        .CLK(clk), .Q(delay_set[1]) );
  DFFSSRX1_HVT set_reg_1_ ( .D(1'b0), .SETB(n194), .RSTB(delay_set[1]), .CLK(
        clk), .Q(set[1]) );
  DFFSSRX1_HVT conv2_weight_cnt_reg_1_ ( .D(1'b0), .SETB(n202), .RSTB(set[1]), 
        .CLK(clk), .Q(conv2_weight_cnt[1]) );
  DFFSSRX1_HVT conv1_weight_cnt_reg_1_ ( .D(1'b0), .SETB(n196), .RSTB(
        conv2_weight_cnt[1]), .CLK(clk), .Q(conv1_weight_cnt[1]) );
  DFFSSRX1_HVT conv1_done_reg ( .D(1'b0), .SETB(n211), .RSTB(n_conv1_done), 
        .CLK(clk), .Q(conv1_done), .QN(n462) );
  DFFSSRX1_HVT col_reg_0_ ( .D(1'b0), .SETB(n209), .RSTB(net22654), .CLK(
        net22658), .Q(col[0]), .QN(n262) );
  DFFSSRX1_HVT col_delay_reg_0_ ( .D(1'b0), .SETB(n169), .RSTB(col[0]), .CLK(
        clk), .Q(col_delay[0]) );
  DFFSSRX1_HVT write_col_reg_0_ ( .D(1'b0), .SETB(n186), .RSTB(col_delay[0]), 
        .CLK(clk), .Q(write_col[0]) );
  DFFSSRX1_HVT col_enable_reg_0_ ( .D(1'b0), .SETB(n177), .RSTB(write_col[0]), 
        .CLK(clk), .Q(col_enable[0]) );
  DFFSSRX1_HVT write_col_conv1_reg_0_ ( .D(1'b0), .SETB(n176), .RSTB(
        col_enable[0]), .CLK(clk), .Q(write_col_conv1[0]) );
  DFFSSRX1_HVT col_reg_1_ ( .D(1'b0), .SETB(n175), .RSTB(net22649), .CLK(
        net22658), .Q(col[1]), .QN(n319) );
  DFFSSRX1_HVT col_delay_reg_1_ ( .D(1'b0), .SETB(n174), .RSTB(col[1]), .CLK(
        clk), .Q(col_delay[1]) );
  DFFSSRX1_HVT write_col_reg_1_ ( .D(1'b0), .SETB(n212), .RSTB(col_delay[1]), 
        .CLK(clk), .Q(write_col[1]) );
  DFFSSRX1_HVT col_enable_reg_1_ ( .D(1'b0), .SETB(n210), .RSTB(write_col[1]), 
        .CLK(clk), .Q(col_enable[1]) );
  DFFSSRX1_HVT write_col_conv1_reg_1_ ( .D(1'b0), .SETB(n169), .RSTB(
        col_enable[1]), .CLK(clk), .Q(write_col_conv1[1]), .QN(n312) );
  DFFSSRX1_HVT col_reg_2_ ( .D(1'b0), .SETB(n185), .RSTB(net22644), .CLK(
        net22658), .Q(col[2]), .QN(n235) );
  DFFSSRX1_HVT col_delay_reg_2_ ( .D(1'b0), .SETB(n177), .RSTB(col[2]), .CLK(
        clk), .Q(col_delay[2]) );
  DFFSSRX1_HVT write_col_reg_2_ ( .D(1'b0), .SETB(n176), .RSTB(col_delay[2]), 
        .CLK(clk), .Q(write_col[2]) );
  DFFSSRX1_HVT col_enable_reg_2_ ( .D(1'b0), .SETB(n175), .RSTB(write_col[2]), 
        .CLK(clk), .Q(col_enable[2]) );
  DFFSSRX1_HVT write_col_conv1_reg_2_ ( .D(1'b0), .SETB(n174), .RSTB(
        col_enable[2]), .CLK(clk), .Q(n257), .QN(n1063) );
  DFFSSRX1_HVT col_reg_3_ ( .D(1'b0), .SETB(n211), .RSTB(net22639), .CLK(
        net22658), .Q(col[3]), .QN(n241) );
  DFFSSRX1_HVT col_delay_reg_3_ ( .D(1'b0), .SETB(n209), .RSTB(col[3]), .CLK(
        clk), .Q(col_delay[3]) );
  DFFSSRX1_HVT write_col_reg_3_ ( .D(1'b0), .SETB(n187), .RSTB(col_delay[3]), 
        .CLK(clk), .Q(write_col[3]) );
  DFFSSRX1_HVT col_enable_reg_3_ ( .D(1'b0), .SETB(n184), .RSTB(write_col[3]), 
        .CLK(clk), .Q(col_enable[3]) );
  DFFSSRX1_HVT write_col_conv1_reg_3_ ( .D(1'b0), .SETB(n198), .RSTB(
        col_enable[3]), .CLK(clk), .Q(n258), .QN(n1062) );
  DFFSSRX1_HVT addr_col_sel_cnt_reg_0_ ( .D(1'b0), .SETB(n193), .RSTB(
        n_addr_col_sel_cnt[0]), .CLK(clk), .Q(addr_col_sel_cnt[0]), .QN(n1052)
         );
  DFFSSRX1_HVT data_sel_col_reg_0_ ( .D(1'b0), .SETB(n201), .RSTB(
        addr_col_sel_cnt[0]), .CLK(clk), .Q(data_sel_col[0]) );
  DFFSSRX1_HVT addr_col_sel_cnt_reg_1_ ( .D(1'b0), .SETB(n195), .RSTB(
        n_addr_col_sel_cnt[1]), .CLK(clk), .Q(addr_col_sel_cnt[1]), .QN(n1051)
         );
  DFFSSRX1_HVT data_sel_col_reg_1_ ( .D(1'b0), .SETB(n212), .RSTB(
        addr_col_sel_cnt[1]), .CLK(clk), .Q(data_sel_col[1]) );
  DFFSSRX1_HVT addr_row_sel_cnt_reg_0_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_addr_row_sel_cnt_0_), .CLK(clk), .Q(addr_row_sel_cnt[0]), .QN(n338)
         );
  DFFSSRX1_HVT data_sel_row_reg_0_ ( .D(1'b0), .SETB(n169), .RSTB(
        addr_row_sel_cnt[0]), .CLK(clk), .Q(data_sel_row[0]) );
  DFFSSRX1_HVT addr_row_sel_cnt_reg_1_ ( .D(n392), .SETB(n1667), .RSTB(n183), 
        .CLK(clk), .Q(addr_row_sel_cnt[1]), .QN(n1053) );
  DFFSSRX1_HVT data_sel_row_reg_1_ ( .D(1'b0), .SETB(n186), .RSTB(
        addr_row_sel_cnt[1]), .CLK(clk), .Q(data_sel_row[1]) );
  DFFSSRX1_HVT conv2_weight_done_reg ( .D(1'b0), .SETB(n199), .RSTB(net22655), 
        .CLK(net22658), .Q(conv2_weight_done) );
  DFFSSRX1_HVT row_reg_0_ ( .D(1'b0), .SETB(n194), .RSTB(n_row[0]), .CLK(
        net22658), .Q(row[0]), .QN(n259) );
  DFFSSRX1_HVT row_delay_reg_0_ ( .D(1'b0), .SETB(n202), .RSTB(row[0]), .CLK(
        clk), .Q(row_delay[0]) );
  DFFSSRX1_HVT write_row_reg_0_ ( .D(1'b0), .SETB(n196), .RSTB(row_delay[0]), 
        .CLK(clk), .Q(write_row[0]) );
  DFFSSRX1_HVT row_enable_reg_0_ ( .D(1'b0), .SETB(n211), .RSTB(write_row[0]), 
        .CLK(clk), .Q(row_enable[0]) );
  DFFSSRX1_HVT write_row_conv1_reg_0_ ( .D(1'b0), .SETB(n209), .RSTB(
        row_enable[0]), .CLK(clk), .Q(write_row_conv1[0]) );
  DFFSSRX1_HVT sram_bytemask_d_reg_1_ ( .D(1'b0), .SETB(n169), .RSTB(
        n_sram_bytemask_d[1]), .CLK(clk), .Q(sram_bytemask_d[1]) );
  DFFSSRX1_HVT sram_bytemask_c_reg_1_ ( .D(1'b0), .SETB(n185), .RSTB(
        n_sram_bytemask_c[1]), .CLK(clk), .Q(sram_bytemask_c[1]) );
  DFFSSRX1_HVT sram_bytemask_d_reg_0_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_bytemask_d[0]), .CLK(clk), .Q(sram_bytemask_d[0]) );
  DFFSSRX1_HVT sram_bytemask_c_reg_0_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_bytemask_c[0]), .CLK(clk), .Q(sram_bytemask_c[0]) );
  DFFSSRX1_HVT sram_bytemask_c_reg_2_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_bytemask_c[2]), .CLK(clk), .Q(sram_bytemask_c[2]) );
  DFFSSRX1_HVT sram_bytemask_c_reg_3_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_bytemask_c[3]), .CLK(clk), .Q(sram_bytemask_c[3]) );
  DFFSSRX1_HVT sram_bytemask_d_reg_2_ ( .D(1'b0), .SETB(n212), .RSTB(
        n_sram_bytemask_d[2]), .CLK(clk), .Q(sram_bytemask_d[2]) );
  DFFSSRX1_HVT sram_bytemask_d_reg_3_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_bytemask_d[3]), .CLK(clk), .Q(sram_bytemask_d[3]) );
  DFFSSRX1_HVT row_reg_1_ ( .D(1'b0), .SETB(n187), .RSTB(n_row[1]), .CLK(
        net22658), .Q(row[1]), .QN(n349) );
  DFFSSRX1_HVT row_delay_reg_1_ ( .D(1'b0), .SETB(n184), .RSTB(row[1]), .CLK(
        clk), .Q(row_delay[1]) );
  DFFSSRX1_HVT write_row_reg_1_ ( .D(1'b0), .SETB(n177), .RSTB(row_delay[1]), 
        .CLK(clk), .Q(write_row[1]) );
  DFFSSRX1_HVT row_enable_reg_1_ ( .D(1'b0), .SETB(n176), .RSTB(write_row[1]), 
        .CLK(clk), .Q(row_enable[1]) );
  DFFSSRX1_HVT write_row_conv1_reg_1_ ( .D(1'b0), .SETB(n175), .RSTB(
        row_enable[1]), .CLK(clk), .Q(n249), .QN(n1061) );
  DFFSSRX1_HVT box_sel_reg_2_ ( .D(n371), .SETB(n1655), .RSTB(n182), .CLK(clk), 
        .Q(box_sel[2]) );
  DFFSSRX1_HVT box_sel_reg_1_ ( .D(1'b0), .SETB(n174), .RSTB(n_box_sel_1_), 
        .CLK(clk), .Q(box_sel[1]) );
  DFFSSRX1_HVT box_sel_reg_0_ ( .D(n369), .SETB(n1662), .RSTB(n231), .CLK(clk), 
        .Q(box_sel[0]) );
  DFFSSRX1_HVT box_sel_reg_3_ ( .D(n368), .SETB(n1655), .RSTB(n183), .CLK(clk), 
        .Q(box_sel[3]) );
  DFFSSRX1_HVT row_reg_2_ ( .D(1'b0), .SETB(n211), .RSTB(n_row[2]), .CLK(
        net22658), .Q(row[2]), .QN(n256) );
  DFFSSRX1_HVT row_delay_reg_2_ ( .D(1'b0), .SETB(n209), .RSTB(row[2]), .CLK(
        clk), .Q(row_delay[2]) );
  DFFSSRX1_HVT write_row_reg_2_ ( .D(1'b0), .SETB(n169), .RSTB(row_delay[2]), 
        .CLK(clk), .Q(write_row[2]) );
  DFFSSRX1_HVT row_enable_reg_2_ ( .D(1'b0), .SETB(n186), .RSTB(write_row[2]), 
        .CLK(clk), .Q(row_enable[2]) );
  DFFSSRX1_HVT write_row_conv1_reg_2_ ( .D(1'b0), .SETB(n198), .RSTB(
        row_enable[2]), .CLK(clk), .Q(write_row_conv1[2]), .QN(n289) );
  DFFSSRX1_HVT row_reg_3_ ( .D(1'b0), .SETB(n193), .RSTB(n_row[3]), .CLK(
        net22658), .Q(row[3]), .QN(n313) );
  DFFSSRX1_HVT row_delay_reg_3_ ( .D(1'b0), .SETB(n201), .RSTB(row[3]), .CLK(
        clk), .Q(row_delay[3]) );
  DFFSSRX1_HVT write_row_reg_3_ ( .D(1'b0), .SETB(n195), .RSTB(row_delay[3]), 
        .CLK(clk), .Q(write_row[3]) );
  DFFSSRX1_HVT row_enable_reg_3_ ( .D(1'b0), .SETB(n212), .RSTB(write_row[3]), 
        .CLK(clk), .Q(row_enable[3]) );
  DFFSSRX1_HVT write_row_conv1_reg_3_ ( .D(1'b0), .SETB(n210), .RSTB(
        row_enable[3]), .CLK(clk), .Q(write_row_conv1[3]), .QN(n357) );
  DFFSSRX1_HVT channel_cnt_reg_4_ ( .D(1'b0), .SETB(n169), .RSTB(net22934), 
        .CLK(net22941), .Q(channel_cnt[4]), .QN(n314) );
  DFFSSRX1_HVT channel_cnt_reg_3_ ( .D(1'b0), .SETB(n185), .RSTB(net22935), 
        .CLK(net22941), .Q(channel_cnt[3]) );
  DFFSSRX1_HVT channel_cnt_reg_2_ ( .D(1'b0), .SETB(n199), .RSTB(net22936), 
        .CLK(net22941), .Q(channel_cnt[2]), .QN(n435) );
  DFFSSRX1_HVT channel_cnt_reg_1_ ( .D(1'b0), .SETB(n194), .RSTB(net22937), 
        .CLK(net22941), .Q(channel_cnt[1]) );
  DFFSSRX1_HVT load_conv1_bias_enable_reg ( .D(1'b0), .SETB(n202), .RSTB(n1020), .CLK(clk), .Q(load_conv1_bias_enable) );
  DFFSSRX1_HVT sram_raddr_weight_reg_7_ ( .D(1'b0), .SETB(n196), .RSTB(
        net22783), .CLK(net22856), .Q(sram_raddr_weight[7]), .QN(n359) );
  DFFSSRX1_HVT conv1_bias_set_reg_7_ ( .D(1'b0), .SETB(n211), .RSTB(
        sram_raddr_weight[7]), .CLK(clk), .Q(conv1_bias_set[7]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_6_ ( .D(1'b0), .SETB(n209), .RSTB(
        net22790), .CLK(net22856), .Q(sram_raddr_weight[6]), .QN(n358) );
  DFFSSRX1_HVT conv1_bias_set_reg_6_ ( .D(1'b0), .SETB(n187), .RSTB(
        sram_raddr_weight[6]), .CLK(clk), .Q(conv1_bias_set[6]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_5_ ( .D(1'b0), .SETB(n184), .RSTB(
        net22797), .CLK(net22856), .Q(sram_raddr_weight[5]), .QN(n437) );
  DFFSSRX1_HVT conv1_bias_set_reg_5_ ( .D(1'b0), .SETB(n177), .RSTB(
        sram_raddr_weight[5]), .CLK(clk), .Q(conv1_bias_set[5]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_3_ ( .D(1'b0), .SETB(n176), .RSTB(
        net22818), .CLK(net22856), .Q(sram_raddr_weight[3]), .QN(n432) );
  DFFSSRX1_HVT conv1_bias_set_reg_3_ ( .D(1'b0), .SETB(n175), .RSTB(
        sram_raddr_weight[3]), .CLK(clk), .Q(conv1_bias_set[3]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_16_ ( .D(1'b0), .SETB(n174), .RSTB(
        net22692), .CLK(net22758), .Q(sram_raddr_weight[16]), .QN(n463) );
  DFFSSRX1_HVT conv1_bias_set_reg_16_ ( .D(1'b0), .SETB(n212), .RSTB(
        sram_raddr_weight[16]), .CLK(clk), .Q(conv1_bias_set[16]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_15_ ( .D(1'b0), .SETB(n210), .RSTB(
        net22699), .CLK(net22758), .Q(sram_raddr_weight[15]), .QN(n304) );
  DFFSSRX1_HVT conv1_bias_set_reg_15_ ( .D(1'b0), .SETB(n169), .RSTB(
        sram_raddr_weight[15]), .CLK(clk), .Q(conv1_bias_set[15]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_14_ ( .D(1'b0), .SETB(n186), .RSTB(
        net22706), .CLK(net22758), .Q(sram_raddr_weight[14]), .QN(n403) );
  DFFSSRX1_HVT conv1_bias_set_reg_14_ ( .D(1'b0), .SETB(n177), .RSTB(
        sram_raddr_weight[14]), .CLK(clk), .Q(conv1_bias_set[14]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_13_ ( .D(1'b0), .SETB(n176), .RSTB(
        net22713), .CLK(net22758), .Q(sram_raddr_weight[13]) );
  DFFSSRX1_HVT conv1_bias_set_reg_13_ ( .D(1'b0), .SETB(n175), .RSTB(
        sram_raddr_weight[13]), .CLK(clk), .Q(conv1_bias_set[13]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_12_ ( .D(1'b0), .SETB(n174), .RSTB(
        net22720), .CLK(net22758), .Q(sram_raddr_weight[12]), .QN(n429) );
  DFFSSRX1_HVT conv1_bias_set_reg_12_ ( .D(1'b0), .SETB(n211), .RSTB(
        sram_raddr_weight[12]), .CLK(clk), .Q(conv1_bias_set[12]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_11_ ( .D(1'b0), .SETB(n209), .RSTB(
        net22727), .CLK(net22758), .Q(sram_raddr_weight[11]) );
  DFFSSRX1_HVT conv1_bias_set_reg_11_ ( .D(1'b0), .SETB(n169), .RSTB(
        sram_raddr_weight[11]), .CLK(clk), .Q(conv1_bias_set[11]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_10_ ( .D(1'b0), .SETB(n185), .RSTB(
        net22734), .CLK(net22758), .Q(sram_raddr_weight[10]), .QN(n430) );
  DFFSSRX1_HVT conv1_bias_set_reg_10_ ( .D(1'b0), .SETB(n198), .RSTB(
        sram_raddr_weight[10]), .CLK(clk), .Q(conv1_bias_set[10]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_9_ ( .D(1'b0), .SETB(n193), .RSTB(
        net22748), .CLK(net22758), .Q(sram_raddr_weight[9]), .QN(n288) );
  DFFSSRX1_HVT conv1_bias_set_reg_9_ ( .D(1'b0), .SETB(n201), .RSTB(
        sram_raddr_weight[9]), .CLK(clk), .Q(conv1_bias_set[9]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_8_ ( .D(1'b0), .SETB(n195), .RSTB(
        net22755), .CLK(net22758), .Q(sram_raddr_weight[8]), .QN(n355) );
  DFFSSRX1_HVT conv1_bias_set_reg_8_ ( .D(1'b0), .SETB(n212), .RSTB(
        sram_raddr_weight[8]), .CLK(clk), .Q(conv1_bias_set[8]) );
  DFFSSRX1_HVT load_conv2_bias0_enable_reg ( .D(1'b0), .SETB(n210), .RSTB(
        n1021), .CLK(clk), .Q(load_conv2_bias0_enable) );
  DFFSSRX1_HVT conv1_weight_done_reg ( .D(1'b0), .SETB(n187), .RSTB(
        n_conv1_weight_done), .CLK(clk), .Q(conv1_weight_done), .QN(n254) );
  DFFSSRX1_HVT load_data_enable_reg ( .D(1'b0), .SETB(n184), .RSTB(
        n_load_data_enable), .CLK(clk), .Q(load_data_enable) );
  DFFSSRX1_HVT write_enable_reg ( .D(1'b0), .SETB(n199), .RSTB(n_write_enable), 
        .CLK(clk), .Q(write_enable) );
  DFFSSRX1_HVT delay_write_enable_reg ( .D(1'b0), .SETB(n194), .RSTB(
        write_enable), .CLK(clk), .Q(delay_write_enable) );
  DFFSSRX1_HVT delay2_write_enable_reg ( .D(1'b0), .SETB(n202), .RSTB(
        delay_write_enable), .CLK(clk), .Q(delay2_write_enable) );
  DFFSSRX1_HVT delay3_write_enable_reg ( .D(1'b0), .SETB(n196), .RSTB(
        delay2_write_enable), .CLK(clk), .Q(delay3_write_enable) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_9_ ( .D(1'b0), .SETB(N2914), .RSTB(
        net22864), .CLK(net22894), .Q(delay1_sram_waddr_b[9]) );
  DFFSSRX1_HVT sram_waddr_b_reg_9_ ( .D(1'b0), .SETB(n211), .RSTB(
        delay1_sram_waddr_b[9]), .CLK(clk), .Q(sram_waddr_b[9]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_8_ ( .D(1'b0), .SETB(N2914), .RSTB(
        net22867), .CLK(net22894), .Q(delay1_sram_waddr_b[8]), .QN(n445) );
  DFFSSRX1_HVT sram_waddr_b_reg_8_ ( .D(1'b0), .SETB(n209), .RSTB(
        delay1_sram_waddr_b[8]), .CLK(clk), .Q(sram_waddr_b[8]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_7_ ( .D(1'b0), .SETB(N2914), .RSTB(
        net22870), .CLK(net22894), .Q(delay1_sram_waddr_b[7]) );
  DFFSSRX1_HVT sram_waddr_b_reg_7_ ( .D(1'b0), .SETB(n169), .RSTB(
        delay1_sram_waddr_b[7]), .CLK(clk), .Q(sram_waddr_b[7]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_6_ ( .D(1'b0), .SETB(N2914), .RSTB(
        net22873), .CLK(net22894), .Q(delay1_sram_waddr_b[6]), .QN(n408) );
  DFFSSRX1_HVT sram_waddr_b_reg_6_ ( .D(1'b0), .SETB(n186), .RSTB(
        delay1_sram_waddr_b[6]), .CLK(clk), .Q(sram_waddr_b[6]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_5_ ( .D(1'b0), .SETB(N2914), .RSTB(
        net22876), .CLK(net22894), .Q(delay1_sram_waddr_b[5]) );
  DFFSSRX1_HVT sram_waddr_b_reg_5_ ( .D(1'b0), .SETB(n177), .RSTB(
        delay1_sram_waddr_b[5]), .CLK(clk), .Q(sram_waddr_b[5]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_4_ ( .D(1'b0), .SETB(N2914), .RSTB(
        net22879), .CLK(net22894), .Q(delay1_sram_waddr_b[4]), .QN(n344) );
  DFFSSRX1_HVT sram_waddr_b_reg_4_ ( .D(1'b0), .SETB(n176), .RSTB(
        delay1_sram_waddr_b[4]), .CLK(clk), .Q(sram_waddr_b[4]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_3_ ( .D(1'b0), .SETB(N2914), .RSTB(
        net22882), .CLK(net22894), .Q(delay1_sram_waddr_b[3]) );
  DFFSSRX1_HVT sram_waddr_b_reg_3_ ( .D(1'b0), .SETB(n175), .RSTB(
        delay1_sram_waddr_b[3]), .CLK(clk), .Q(sram_waddr_b[3]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_2_ ( .D(1'b0), .SETB(N2914), .RSTB(
        net22885), .CLK(net22894), .Q(delay1_sram_waddr_b[2]), .QN(n428) );
  DFFSSRX1_HVT sram_waddr_b_reg_2_ ( .D(1'b0), .SETB(n174), .RSTB(
        delay1_sram_waddr_b[2]), .CLK(clk), .Q(sram_waddr_b[2]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_1_ ( .D(1'b0), .SETB(N2914), .RSTB(
        net22888), .CLK(net22894), .Q(delay1_sram_waddr_b[1]) );
  DFFSSRX1_HVT sram_waddr_b_reg_1_ ( .D(1'b0), .SETB(n212), .RSTB(
        delay1_sram_waddr_b[1]), .CLK(clk), .Q(sram_waddr_b[1]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_0_ ( .D(1'b0), .SETB(N2914), .RSTB(
        net22891), .CLK(net22894), .Q(delay1_sram_waddr_b[0]) );
  DFFSSRX1_HVT sram_waddr_b_reg_0_ ( .D(1'b0), .SETB(n210), .RSTB(
        delay1_sram_waddr_b[0]), .CLK(clk), .Q(sram_waddr_b[0]) );
  DFFSSRX1_HVT sram_bytemask_b_reg_3_ ( .D(1'b0), .SETB(n169), .RSTB(
        n_sram_bytemask_b[3]), .CLK(clk), .Q(sram_bytemask_b[3]) );
  DFFSSRX1_HVT sram_bytemask_b_reg_2_ ( .D(1'b0), .SETB(n185), .RSTB(
        n_sram_bytemask_b[2]), .CLK(clk), .Q(sram_bytemask_b[2]) );
  DFFSSRX1_HVT sram_bytemask_b_reg_1_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_bytemask_b[1]), .CLK(clk), .Q(sram_bytemask_b[1]) );
  DFFSSRX1_HVT sram_bytemask_b_reg_0_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_bytemask_b[0]), .CLK(clk), .Q(sram_bytemask_b[0]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_1_ ( .D(1'b0), .SETB(n175), .RSTB(
        net22839), .CLK(net22856), .Q(sram_raddr_weight[1]), .QN(n436) );
  DFFSSRX1_HVT conv1_bias_set_reg_1_ ( .D(1'b0), .SETB(n174), .RSTB(
        sram_raddr_weight[1]), .CLK(clk), .Q(conv1_bias_set[1]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_0_ ( .D(1'b0), .SETB(n211), .RSTB(
        net22853), .CLK(net22856), .Q(sram_raddr_weight[0]), .QN(n309) );
  DFFSSRX1_HVT conv1_bias_set_reg_0_ ( .D(1'b0), .SETB(n209), .RSTB(
        sram_raddr_weight[0]), .CLK(clk), .Q(conv1_bias_set[0]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_2_ ( .D(1'b0), .SETB(n187), .RSTB(
        net22825), .CLK(net22856), .Q(sram_raddr_weight[2]), .QN(n305) );
  DFFSSRX1_HVT conv1_bias_set_reg_2_ ( .D(1'b0), .SETB(n184), .RSTB(
        sram_raddr_weight[2]), .CLK(clk), .Q(conv1_bias_set[2]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_4_ ( .D(1'b0), .SETB(n198), .RSTB(
        net22811), .CLK(net22856), .Q(sram_raddr_weight[4]), .QN(n447) );
  DFFSSRX1_HVT conv1_bias_set_reg_4_ ( .D(1'b0), .SETB(n193), .RSTB(
        sram_raddr_weight[4]), .CLK(clk), .Q(conv1_bias_set[4]) );
  DFFSSRX1_HVT load_conv2_bias1_enable_reg ( .D(1'b0), .SETB(n201), .RSTB(
        n1022), .CLK(clk), .Q(load_conv2_bias1_enable) );
  DFFSSRX1_HVT addr_change_reg_0_ ( .D(1'b0), .SETB(n195), .RSTB(net22950), 
        .CLK(net22953), .Q(addr_change[0]) );
  DFFSSRX1_HVT addr_change_reg_1_ ( .D(1'b0), .SETB(n212), .RSTB(net22949), 
        .CLK(net22953), .Q(addr_change[1]) );
  DFFSSRX1_HVT addr_change_reg_2_ ( .D(1'b0), .SETB(n210), .RSTB(net22948), 
        .CLK(net22953), .Q(addr_change[2]) );
  DFFSSRX1_HVT addr_change_reg_3_ ( .D(1'b0), .SETB(n169), .RSTB(net22947), 
        .CLK(net22953), .Q(addr_change[3]), .QN(n454) );
  DFFSSRX1_HVT addr_change_reg_4_ ( .D(1'b0), .SETB(n186), .RSTB(net22946), 
        .CLK(net22953), .Q(addr_change[4]), .QN(n460) );
  DFFSSRX1_HVT delay_addr_change_reg_4_ ( .D(1'b0), .SETB(n199), .RSTB(
        addr_change[4]), .CLK(clk), .Q(delay_addr_change[4]) );
  DFFSSRX1_HVT delay_addr_change_reg_3_ ( .D(1'b0), .SETB(n194), .RSTB(
        addr_change[3]), .CLK(clk), .Q(delay_addr_change[3]) );
  DFFSSRX1_HVT delay_addr_change_reg_2_ ( .D(1'b0), .SETB(n202), .RSTB(
        addr_change[2]), .CLK(clk), .Q(delay_addr_change[2]) );
  DFFSSRX1_HVT delay_addr_change_reg_1_ ( .D(1'b0), .SETB(n196), .RSTB(
        addr_change[1]), .CLK(clk), .Q(delay_addr_change[1]) );
  DFFSSRX1_HVT delay_addr_change_reg_0_ ( .D(1'b0), .SETB(n211), .RSTB(
        addr_change[0]), .CLK(clk), .Q(delay_addr_change[0]) );
  DFFSSRX1_HVT delay2_addr_change_reg_4_ ( .D(1'b0), .SETB(n209), .RSTB(
        delay_addr_change[4]), .CLK(clk), .Q(delay2_addr_change[4]) );
  DFFSSRX1_HVT delay2_addr_change_reg_3_ ( .D(1'b0), .SETB(n169), .RSTB(
        delay_addr_change[3]), .CLK(clk), .Q(delay2_addr_change[3]) );
  DFFSSRX1_HVT delay2_addr_change_reg_2_ ( .D(1'b0), .SETB(n185), .RSTB(
        delay_addr_change[2]), .CLK(clk), .Q(delay2_addr_change[2]) );
  DFFSSRX1_HVT delay2_addr_change_reg_1_ ( .D(1'b0), .SETB(n177), .RSTB(
        delay_addr_change[1]), .CLK(clk), .Q(delay2_addr_change[1]) );
  DFFSSRX1_HVT delay2_addr_change_reg_0_ ( .D(1'b0), .SETB(n176), .RSTB(
        delay_addr_change[0]), .CLK(clk), .Q(delay2_addr_change[0]) );
  DFFSSRX1_HVT delay3_addr_change_reg_4_ ( .D(1'b0), .SETB(n175), .RSTB(
        delay2_addr_change[4]), .CLK(clk), .Q(delay3_addr_change[4]), .QN(n469) );
  DFFSSRX1_HVT delay3_addr_change_reg_3_ ( .D(1'b0), .SETB(n174), .RSTB(
        delay2_addr_change[3]), .CLK(clk), .Q(delay3_addr_change[3]), .QN(n311) );
  DFFSSRX1_HVT delay3_addr_change_reg_2_ ( .D(1'b0), .SETB(n212), .RSTB(
        delay2_addr_change[2]), .CLK(clk), .Q(delay3_addr_change[2]), .QN(n255) );
  DFFSSRX1_HVT delay3_addr_change_reg_1_ ( .D(1'b0), .SETB(n210), .RSTB(
        delay2_addr_change[1]), .CLK(clk), .Q(delay3_addr_change[1]) );
  DFFSSRX1_HVT delay3_addr_change_reg_0_ ( .D(1'b0), .SETB(n187), .RSTB(
        delay2_addr_change[0]), .CLK(clk), .Q(delay3_addr_change[0]) );
  DFFSSRX1_HVT delay_channel_reg_4_ ( .D(1'b0), .SETB(n208), .RSTB(
        channel_cnt[4]), .CLK(clk), .Q(delay_channel[4]) );
  DFFSSRX1_HVT delay_channel_reg_3_ ( .D(1'b0), .SETB(n201), .RSTB(
        channel_cnt[3]), .CLK(clk), .Q(delay_channel[3]) );
  DFFSSRX1_HVT delay_channel_reg_2_ ( .D(1'b0), .SETB(n186), .RSTB(
        channel_cnt[2]), .CLK(clk), .Q(delay_channel[2]) );
  DFFSSRX1_HVT delay_channel_reg_1_ ( .D(1'b0), .SETB(n199), .RSTB(
        channel_cnt[1]), .CLK(clk), .Q(delay_channel[1]) );
  DFFSSRX1_HVT delay_channel_reg_0_ ( .D(1'b0), .SETB(n196), .RSTB(
        channel_cnt[0]), .CLK(clk), .Q(delay_channel[0]) );
  DFFSSRX1_HVT delay2_channel_reg_4_ ( .D(1'b0), .SETB(n198), .RSTB(
        delay_channel[4]), .CLK(clk), .Q(delay2_channel[4]) );
  DFFSSRX1_HVT delay2_channel_reg_3_ ( .D(1'b0), .SETB(n195), .RSTB(
        delay_channel[3]), .CLK(clk), .Q(delay2_channel[3]) );
  DFFSSRX1_HVT delay2_channel_reg_2_ ( .D(1'b0), .SETB(n177), .RSTB(
        delay_channel[2]), .CLK(clk), .Q(delay2_channel[2]) );
  DFFSSRX1_HVT delay2_channel_reg_1_ ( .D(1'b0), .SETB(n194), .RSTB(
        delay_channel[1]), .CLK(clk), .Q(delay2_channel[1]) );
  DFFSSRX1_HVT delay2_channel_reg_0_ ( .D(1'b0), .SETB(n187), .RSTB(
        delay_channel[0]), .CLK(clk), .Q(delay2_channel[0]) );
  DFFSSRX1_HVT channel_reg_4_ ( .D(1'b0), .SETB(n193), .RSTB(delay2_channel[4]), .CLK(clk), .Q(channel[4]) );
  DFFSSRX1_HVT channel_reg_3_ ( .D(1'b0), .SETB(n169), .RSTB(delay2_channel[3]), .CLK(clk), .Q(channel[3]) );
  DFFSSRX1_HVT channel_reg_2_ ( .D(1'b0), .SETB(n208), .RSTB(delay2_channel[2]), .CLK(clk), .Q(channel[2]) );
  DFFSSRX1_HVT channel_reg_1_ ( .D(1'b0), .SETB(n202), .RSTB(delay2_channel[1]), .CLK(clk), .Q(channel[1]) );
  DFFSSRX1_HVT channel_reg_0_ ( .D(1'b0), .SETB(n184), .RSTB(delay2_channel[0]), .CLK(clk), .Q(channel[0]) );
  DFFSSRX1_HVT delay1_state_reg_3_ ( .D(1'b0), .SETB(n184), .RSTB(state[3]), 
        .CLK(clk), .Q(delay1_state[3]) );
  DFFSSRX1_HVT delay2_state_reg_3_ ( .D(1'b0), .SETB(n177), .RSTB(
        delay1_state[3]), .CLK(clk), .Q(delay2_state[3]) );
  DFFSSRX1_HVT delay3_state_reg_3_ ( .D(1'b0), .SETB(n176), .RSTB(
        delay2_state[3]), .CLK(clk), .QN(n1027) );
  DFFSSRX1_HVT delay1_state_reg_2_ ( .D(1'b0), .SETB(n175), .RSTB(state[2]), 
        .CLK(clk), .Q(delay1_state[2]) );
  DFFSSRX1_HVT delay2_state_reg_2_ ( .D(1'b0), .SETB(n174), .RSTB(
        delay1_state[2]), .CLK(clk), .Q(delay2_state[2]) );
  DFFSSRX1_HVT delay3_state_reg_2_ ( .D(1'b0), .SETB(n211), .RSTB(
        delay2_state[2]), .CLK(clk), .Q(delay3_state[2]) );
  DFFSSRX1_HVT delay1_state_reg_1_ ( .D(1'b0), .SETB(n209), .RSTB(state[1]), 
        .CLK(clk), .Q(delay1_state[1]) );
  DFFSSRX1_HVT delay2_state_reg_1_ ( .D(1'b0), .SETB(n169), .RSTB(
        delay1_state[1]), .CLK(clk), .Q(delay2_state[1]) );
  DFFSSRX1_HVT delay3_state_reg_1_ ( .D(1'b0), .SETB(n186), .RSTB(
        delay2_state[1]), .CLK(clk), .Q(delay3_state[1]) );
  DFFSSRX1_HVT delay1_state_reg_0_ ( .D(1'b0), .SETB(n198), .RSTB(state[0]), 
        .CLK(clk), .Q(delay1_state[0]) );
  DFFSSRX1_HVT delay2_state_reg_0_ ( .D(1'b0), .SETB(n193), .RSTB(
        delay1_state[0]), .CLK(clk), .Q(delay2_state[0]) );
  DFFSSRX1_HVT delay3_state_reg_0_ ( .D(1'b0), .SETB(n201), .RSTB(
        delay2_state[0]), .CLK(clk), .Q(delay3_state[0]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_9_ ( .D(1'b0), .SETB(n195), .RSTB(
        net22917), .CLK(net22929), .Q(delay1_sram_waddr_d[9]), .QN(n468) );
  DFFSSRX1_HVT sram_waddr_d_reg_9_ ( .D(1'b0), .SETB(n212), .RSTB(
        delay1_sram_waddr_d[9]), .CLK(clk), .Q(sram_waddr_d[9]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_8_ ( .D(1'b0), .SETB(n210), .RSTB(
        net22918), .CLK(net22929), .Q(delay1_sram_waddr_d[8]) );
  DFFSSRX1_HVT sram_waddr_d_reg_8_ ( .D(1'b0), .SETB(n169), .RSTB(
        delay1_sram_waddr_d[8]), .CLK(clk), .Q(sram_waddr_d[8]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_7_ ( .D(1'b0), .SETB(n185), .RSTB(
        net22919), .CLK(net22929), .Q(delay1_sram_waddr_d[7]) );
  DFFSSRX1_HVT sram_waddr_d_reg_7_ ( .D(1'b0), .SETB(n199), .RSTB(
        delay1_sram_waddr_d[7]), .CLK(clk), .Q(sram_waddr_d[7]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_6_ ( .D(1'b0), .SETB(n194), .RSTB(
        net22920), .CLK(net22929), .Q(delay1_sram_waddr_d[6]) );
  DFFSSRX1_HVT sram_waddr_d_reg_6_ ( .D(1'b0), .SETB(n202), .RSTB(
        delay1_sram_waddr_d[6]), .CLK(clk), .Q(sram_waddr_d[6]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_5_ ( .D(1'b0), .SETB(n196), .RSTB(
        net22921), .CLK(net22929), .Q(delay1_sram_waddr_d[5]) );
  DFFSSRX1_HVT sram_waddr_d_reg_5_ ( .D(1'b0), .SETB(n211), .RSTB(
        delay1_sram_waddr_d[5]), .CLK(clk), .Q(sram_waddr_d[5]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_4_ ( .D(1'b0), .SETB(n209), .RSTB(
        net22922), .CLK(net22929), .Q(delay1_sram_waddr_d[4]) );
  DFFSSRX1_HVT sram_waddr_d_reg_4_ ( .D(1'b0), .SETB(n187), .RSTB(
        delay1_sram_waddr_d[4]), .CLK(clk), .Q(sram_waddr_d[4]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_3_ ( .D(1'b0), .SETB(n184), .RSTB(
        net22923), .CLK(net22929), .Q(delay1_sram_waddr_d[3]) );
  DFFSSRX1_HVT sram_waddr_d_reg_3_ ( .D(1'b0), .SETB(n177), .RSTB(
        delay1_sram_waddr_d[3]), .CLK(clk), .Q(sram_waddr_d[3]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_2_ ( .D(1'b0), .SETB(n176), .RSTB(
        net22924), .CLK(net22929), .Q(delay1_sram_waddr_d[2]) );
  DFFSSRX1_HVT sram_waddr_d_reg_2_ ( .D(1'b0), .SETB(n175), .RSTB(
        delay1_sram_waddr_d[2]), .CLK(clk), .Q(sram_waddr_d[2]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_1_ ( .D(1'b0), .SETB(n174), .RSTB(
        net22925), .CLK(net22929), .Q(delay1_sram_waddr_d[1]) );
  DFFSSRX1_HVT sram_waddr_d_reg_1_ ( .D(1'b0), .SETB(n212), .RSTB(
        delay1_sram_waddr_d[1]), .CLK(clk), .Q(sram_waddr_d[1]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_0_ ( .D(1'b0), .SETB(n210), .RSTB(
        net22926), .CLK(net22929), .Q(delay1_sram_waddr_d[0]), .QN(n441) );
  DFFSSRX1_HVT sram_waddr_d_reg_0_ ( .D(1'b0), .SETB(n186), .RSTB(
        delay1_sram_waddr_d[0]), .CLK(clk), .Q(sram_waddr_d[0]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_9_ ( .D(1'b0), .SETB(n208), .RSTB(
        net22901), .CLK(net22913), .Q(delay1_sram_waddr_c[9]), .QN(n467) );
  DFFSSRX1_HVT sram_waddr_c_reg_9_ ( .D(1'b0), .SETB(n177), .RSTB(
        delay1_sram_waddr_c[9]), .CLK(clk), .Q(sram_waddr_c[9]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_8_ ( .D(1'b0), .SETB(n176), .RSTB(
        net22902), .CLK(net22913), .Q(delay1_sram_waddr_c[8]) );
  DFFSSRX1_HVT sram_waddr_c_reg_8_ ( .D(1'b0), .SETB(n175), .RSTB(
        delay1_sram_waddr_c[8]), .CLK(clk), .Q(sram_waddr_c[8]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_7_ ( .D(1'b0), .SETB(n174), .RSTB(
        net22903), .CLK(net22913), .Q(delay1_sram_waddr_c[7]) );
  DFFSSRX1_HVT sram_waddr_c_reg_7_ ( .D(1'b0), .SETB(n211), .RSTB(
        delay1_sram_waddr_c[7]), .CLK(clk), .Q(sram_waddr_c[7]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_6_ ( .D(1'b0), .SETB(n209), .RSTB(
        net22904), .CLK(net22913), .Q(delay1_sram_waddr_c[6]) );
  DFFSSRX1_HVT sram_waddr_c_reg_6_ ( .D(1'b0), .SETB(n185), .RSTB(
        delay1_sram_waddr_c[6]), .CLK(clk), .Q(sram_waddr_c[6]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_5_ ( .D(1'b0), .SETB(n208), .RSTB(
        net22905), .CLK(net22913), .Q(delay1_sram_waddr_c[5]) );
  DFFSSRX1_HVT sram_waddr_c_reg_5_ ( .D(1'b0), .SETB(n198), .RSTB(
        delay1_sram_waddr_c[5]), .CLK(clk), .Q(sram_waddr_c[5]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_4_ ( .D(1'b0), .SETB(n193), .RSTB(
        net22906), .CLK(net22913), .Q(delay1_sram_waddr_c[4]) );
  DFFSSRX1_HVT sram_waddr_c_reg_4_ ( .D(1'b0), .SETB(n201), .RSTB(
        delay1_sram_waddr_c[4]), .CLK(clk), .Q(sram_waddr_c[4]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_3_ ( .D(1'b0), .SETB(n195), .RSTB(
        net22907), .CLK(net22913), .Q(delay1_sram_waddr_c[3]) );
  DFFSSRX1_HVT sram_waddr_c_reg_3_ ( .D(1'b0), .SETB(n212), .RSTB(
        delay1_sram_waddr_c[3]), .CLK(clk), .Q(sram_waddr_c[3]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_2_ ( .D(1'b0), .SETB(n210), .RSTB(
        net22908), .CLK(net22913), .Q(delay1_sram_waddr_c[2]) );
  DFFSSRX1_HVT sram_waddr_c_reg_2_ ( .D(1'b0), .SETB(n186), .RSTB(
        delay1_sram_waddr_c[2]), .CLK(clk), .Q(sram_waddr_c[2]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_1_ ( .D(1'b0), .SETB(n208), .RSTB(
        net22909), .CLK(net22913), .Q(delay1_sram_waddr_c[1]) );
  DFFSSRX1_HVT sram_waddr_c_reg_1_ ( .D(1'b0), .SETB(n199), .RSTB(
        delay1_sram_waddr_c[1]), .CLK(clk), .Q(sram_waddr_c[1]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_0_ ( .D(1'b0), .SETB(n194), .RSTB(
        net22910), .CLK(net22913), .Q(delay1_sram_waddr_c[0]), .QN(n440) );
  DFFSSRX1_HVT sram_waddr_c_reg_0_ ( .D(1'b0), .SETB(n202), .RSTB(
        delay1_sram_waddr_c[0]), .CLK(clk), .Q(sram_waddr_c[0]) );
  DFFSSRX1_HVT sram_raddr_a7_reg_9_ ( .D(1'b0), .SETB(n196), .RSTB(
        n_sram_raddr_a7[9]), .CLK(net23434), .Q(sram_raddr_a7[9]) );
  DFFSSRX1_HVT sram_raddr_a7_reg_8_ ( .D(1'b0), .SETB(n211), .RSTB(
        n_sram_raddr_a7[8]), .CLK(net23434), .Q(sram_raddr_a7[8]) );
  DFFSSRX1_HVT sram_raddr_a7_reg_7_ ( .D(1'b0), .SETB(n209), .RSTB(
        n_sram_raddr_a7[7]), .CLK(net23434), .Q(sram_raddr_a7[7]) );
  DFFSSRX1_HVT sram_raddr_a7_reg_6_ ( .D(1'b0), .SETB(n185), .RSTB(
        n_sram_raddr_a7[6]), .CLK(net23434), .Q(sram_raddr_a7[6]) );
  DFFSSRX1_HVT sram_raddr_a7_reg_5_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_a7[5]), .CLK(net23434), .Q(sram_raddr_a7[5]) );
  DFFSSRX1_HVT sram_raddr_a7_reg_4_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_a7[4]), .CLK(net23434), .Q(sram_raddr_a7[4]) );
  DFFSSRX1_HVT sram_raddr_a7_reg_3_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_a7[3]), .CLK(net23434), .Q(sram_raddr_a7[3]), .QN(n466)
         );
  DFFSSRX1_HVT sram_raddr_a7_reg_2_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_a7[2]), .CLK(net23434), .Q(sram_raddr_a7[2]) );
  DFFSSRX1_HVT sram_raddr_a7_reg_1_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_raddr_a7[1]), .CLK(net23434), .Q(sram_raddr_a7[1]), .QN(n443)
         );
  DFFSSRX1_HVT sram_raddr_a7_reg_0_ ( .D(1'b0), .SETB(n212), .RSTB(
        n_sram_raddr_a7[0]), .CLK(net23434), .Q(sram_raddr_a7[0]), .QN(n303)
         );
  DFFSSRX1_HVT sram_raddr_a8_reg_9_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_a8[9]), .CLK(net24761), .Q(sram_raddr_a8[9]) );
  DFFSSRX1_HVT sram_raddr_a8_reg_8_ ( .D(1'b0), .SETB(n186), .RSTB(
        n_sram_raddr_a8[8]), .CLK(net24761), .Q(sram_raddr_a8[8]) );
  DFFSSRX1_HVT sram_raddr_a8_reg_7_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_a8[7]), .CLK(net24761), .Q(sram_raddr_a8[7]) );
  DFFSSRX1_HVT sram_raddr_a8_reg_6_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_a8[6]), .CLK(net24761), .Q(sram_raddr_a8[6]) );
  DFFSSRX1_HVT sram_raddr_a8_reg_5_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_a8[5]), .CLK(net24761), .Q(sram_raddr_a8[5]) );
  DFFSSRX1_HVT sram_raddr_a8_reg_4_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_a8[4]), .CLK(net24761), .Q(sram_raddr_a8[4]) );
  DFFSSRX1_HVT sram_raddr_a8_reg_3_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_raddr_a8[3]), .CLK(net24761), .Q(sram_raddr_a8[3]) );
  DFFSSRX1_HVT sram_raddr_a8_reg_2_ ( .D(1'b0), .SETB(n211), .RSTB(
        n_sram_raddr_a8[2]), .CLK(net24761), .Q(sram_raddr_a8[2]), .QN(n452)
         );
  DFFSSRX1_HVT sram_raddr_a8_reg_1_ ( .D(1'b0), .SETB(n209), .RSTB(
        n_sram_raddr_a8[1]), .CLK(net24761), .Q(sram_raddr_a8[1]), .QN(n451)
         );
  DFFSSRX1_HVT sram_raddr_a8_reg_0_ ( .D(1'b0), .SETB(n185), .RSTB(
        n_sram_raddr_a8[0]), .CLK(net24761), .Q(sram_raddr_a8[0]), .QN(n302)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_9_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_a0[9]), .CLK(net26089), .Q(sram_raddr_a0[9]), .QN(n457)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_8_ ( .D(1'b0), .SETB(n198), .RSTB(
        n_sram_raddr_a0[8]), .CLK(net26089), .Q(sram_raddr_a0[8]), .QN(n424)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_7_ ( .D(1'b0), .SETB(n193), .RSTB(
        n_sram_raddr_a0[7]), .CLK(net26089), .Q(sram_raddr_a0[7]), .QN(n397)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_6_ ( .D(1'b0), .SETB(n201), .RSTB(
        n_sram_raddr_a0[6]), .CLK(net26089), .Q(sram_raddr_a0[6]), .QN(n446)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_5_ ( .D(1'b0), .SETB(n195), .RSTB(
        n_sram_raddr_a0[5]), .CLK(net26089), .Q(sram_raddr_a0[5]), .QN(n284)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_4_ ( .D(1'b0), .SETB(n212), .RSTB(
        n_sram_raddr_a0[4]), .CLK(net26089), .Q(sram_raddr_a0[4]), .QN(n342)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_3_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_a0[3]), .CLK(net26089), .Q(sram_raddr_a0[3]), .QN(n239)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_2_ ( .D(1'b0), .SETB(n186), .RSTB(
        n_sram_raddr_a0[2]), .CLK(net26089), .Q(sram_raddr_a0[2]), .QN(n248)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_1_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_a0[1]), .CLK(net26089), .Q(sram_raddr_a0[1]), .QN(n422)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_0_ ( .D(1'b0), .SETB(n199), .RSTB(
        n_sram_raddr_a0[0]), .CLK(net26089), .Q(sram_raddr_a0[0]), .QN(n431)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_9_ ( .D(1'b0), .SETB(n194), .RSTB(
        n_sram_raddr_a1[9]), .CLK(net23879), .Q(sram_raddr_a1[9]), .QN(n458)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_8_ ( .D(1'b0), .SETB(n202), .RSTB(
        n_sram_raddr_a1[8]), .CLK(net23879), .Q(sram_raddr_a1[8]), .QN(n425)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_7_ ( .D(1'b0), .SETB(n196), .RSTB(
        n_sram_raddr_a1[7]), .CLK(net23879), .Q(sram_raddr_a1[7]), .QN(n438)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_6_ ( .D(1'b0), .SETB(n211), .RSTB(
        n_sram_raddr_a1[6]), .CLK(net23879), .Q(sram_raddr_a1[6]), .QN(n448)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_5_ ( .D(1'b0), .SETB(n209), .RSTB(
        n_sram_raddr_a1[5]), .CLK(net23879), .Q(sram_raddr_a1[5]), .QN(n345)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_4_ ( .D(1'b0), .SETB(n185), .RSTB(
        n_sram_raddr_a1[4]), .CLK(net23879), .Q(sram_raddr_a1[4]), .QN(n278)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_3_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_a1[3]), .CLK(net23879), .Q(sram_raddr_a1[3]), .QN(n238)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_2_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_a1[2]), .CLK(net23879), .Q(sram_raddr_a1[2]), .QN(n247)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_1_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_a1[1]), .CLK(net23879), .Q(sram_raddr_a1[1]), .QN(n450)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_0_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_a1[0]), .CLK(net23879), .Q(sram_raddr_a1[0]), .QN(n310)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_9_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_raddr_a2[9]), .CLK(net25206), .Q(sram_raddr_a2[9]), .QN(n459)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_8_ ( .D(1'b0), .SETB(n212), .RSTB(
        n_sram_raddr_a2[8]), .CLK(net25206), .Q(sram_raddr_a2[8]), .QN(n449)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_7_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_a2[7]), .CLK(net25206), .Q(sram_raddr_a2[7]), .QN(n398)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_6_ ( .D(1'b0), .SETB(n184), .RSTB(
        n_sram_raddr_a2[6]), .CLK(net25206), .Q(sram_raddr_a2[6]), .QN(n410)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_5_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_a2[5]), .CLK(net25206), .Q(sram_raddr_a2[5]), .QN(n348)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_4_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_a2[4]), .CLK(net25206), .Q(sram_raddr_a2[4]), .QN(n341)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_3_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_a2[3]), .CLK(net25206), .Q(sram_raddr_a2[3]), .QN(n343)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_2_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_a2[2]), .CLK(net25206), .Q(sram_raddr_a2[2]), .QN(n366)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_1_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_raddr_a2[1]), .CLK(net25206), .Q(sram_raddr_a2[1]) );
  DFFSSRX1_HVT sram_raddr_a2_reg_0_ ( .D(1'b0), .SETB(n211), .RSTB(
        n_sram_raddr_a2[0]), .CLK(net25206), .Q(sram_raddr_a2[0]), .QN(n442)
         );
  DFFSSRX1_HVT sram_raddr_a3_reg_9_ ( .D(1'b0), .SETB(n209), .RSTB(
        n_sram_raddr_a3[9]), .CLK(net26535), .Q(sram_raddr_a3[9]) );
  DFFSSRX1_HVT sram_raddr_a3_reg_8_ ( .D(1'b0), .SETB(n186), .RSTB(
        n_sram_raddr_a3[8]), .CLK(net26535), .Q(sram_raddr_a3[8]) );
  DFFSSRX1_HVT sram_raddr_a3_reg_7_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_a3[7]), .CLK(net26535), .Q(sram_raddr_a3[7]), .QN(n412)
         );
  DFFSSRX1_HVT sram_raddr_a3_reg_6_ ( .D(1'b0), .SETB(n198), .RSTB(
        n_sram_raddr_a3[6]), .CLK(net26535), .Q(sram_raddr_a3[6]), .QN(n331)
         );
  DFFSSRX1_HVT sram_raddr_a3_reg_5_ ( .D(1'b0), .SETB(n193), .RSTB(
        n_sram_raddr_a3[5]), .CLK(net26535), .Q(sram_raddr_a3[5]), .QN(n363)
         );
  DFFSSRX1_HVT sram_raddr_a3_reg_4_ ( .D(1'b0), .SETB(n201), .RSTB(
        n_sram_raddr_a3[4]), .CLK(net26535), .Q(sram_raddr_a3[4]), .QN(n275)
         );
  DFFSSRX1_HVT sram_raddr_a3_reg_3_ ( .D(1'b0), .SETB(n195), .RSTB(
        n_sram_raddr_a3[3]), .CLK(net26535), .Q(sram_raddr_a3[3]), .QN(n244)
         );
  DFFSSRX1_HVT sram_raddr_a3_reg_2_ ( .D(1'b0), .SETB(n212), .RSTB(
        n_sram_raddr_a3[2]), .CLK(net26535), .Q(sram_raddr_a3[2]), .QN(n236)
         );
  DFFSSRX1_HVT sram_raddr_a3_reg_1_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_a3[1]), .CLK(net26535), .Q(sram_raddr_a3[1]) );
  DFFSSRX1_HVT sram_raddr_a3_reg_0_ ( .D(1'b0), .SETB(n185), .RSTB(
        n_sram_raddr_a3[0]), .CLK(net26535), .Q(sram_raddr_a3[0]), .QN(n433)
         );
  DFFSSRX1_HVT sram_raddr_a4_reg_9_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_a4[9]), .CLK(net24316), .Q(sram_raddr_a4[9]) );
  DFFSSRX1_HVT sram_raddr_a4_reg_8_ ( .D(1'b0), .SETB(n199), .RSTB(
        n_sram_raddr_a4[8]), .CLK(net24316), .Q(sram_raddr_a4[8]) );
  DFFSSRX1_HVT sram_raddr_a4_reg_7_ ( .D(1'b0), .SETB(n194), .RSTB(
        n_sram_raddr_a4[7]), .CLK(net24316), .Q(sram_raddr_a4[7]) );
  DFFSSRX1_HVT sram_raddr_a4_reg_6_ ( .D(1'b0), .SETB(n202), .RSTB(
        n_sram_raddr_a4[6]), .CLK(net24316), .Q(sram_raddr_a4[6]), .QN(n333)
         );
  DFFSSRX1_HVT sram_raddr_a4_reg_5_ ( .D(1'b0), .SETB(n196), .RSTB(
        n_sram_raddr_a4[5]), .CLK(net24316), .Q(sram_raddr_a4[5]), .QN(n356)
         );
  DFFSSRX1_HVT sram_raddr_a4_reg_4_ ( .D(1'b0), .SETB(n211), .RSTB(
        n_sram_raddr_a4[4]), .CLK(net24316), .Q(sram_raddr_a4[4]), .QN(n246)
         );
  DFFSSRX1_HVT sram_raddr_a4_reg_3_ ( .D(1'b0), .SETB(n209), .RSTB(
        n_sram_raddr_a4[3]), .CLK(net24316), .Q(sram_raddr_a4[3]), .QN(n283)
         );
  DFFSSRX1_HVT sram_raddr_a4_reg_2_ ( .D(1'b0), .SETB(n184), .RSTB(
        n_sram_raddr_a4[2]), .CLK(net24316), .Q(sram_raddr_a4[2]), .QN(n237)
         );
  DFFSSRX1_HVT sram_raddr_a4_reg_1_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_a4[1]), .CLK(net24316), .Q(sram_raddr_a4[1]), .QN(n307)
         );
  DFFSSRX1_HVT sram_raddr_a4_reg_0_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_a4[0]), .CLK(net24316), .Q(sram_raddr_a4[0]), .QN(n417)
         );
  DFFSSRX1_HVT sram_raddr_a5_reg_9_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_a5[9]), .CLK(net25643), .Q(sram_raddr_a5[9]), .QN(n455)
         );
  DFFSSRX1_HVT sram_raddr_a5_reg_8_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_a5[8]), .CLK(net25643), .Q(sram_raddr_a5[8]) );
  DFFSSRX1_HVT sram_raddr_a5_reg_7_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_raddr_a5[7]), .CLK(net25643), .Q(sram_raddr_a5[7]), .QN(n396)
         );
  DFFSSRX1_HVT sram_raddr_a5_reg_6_ ( .D(1'b0), .SETB(n212), .RSTB(
        n_sram_raddr_a5[6]), .CLK(net25643), .Q(sram_raddr_a5[6]), .QN(n362)
         );
  DFFSSRX1_HVT sram_raddr_a5_reg_5_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_a5[5]), .CLK(net25643), .Q(sram_raddr_a5[5]), .QN(n332)
         );
  DFFSSRX1_HVT sram_raddr_a5_reg_4_ ( .D(1'b0), .SETB(n184), .RSTB(
        n_sram_raddr_a5[4]), .CLK(net25643), .Q(sram_raddr_a5[4]), .QN(n361)
         );
  DFFSSRX1_HVT sram_raddr_a5_reg_3_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_a5[3]), .CLK(net25643), .Q(sram_raddr_a5[3]), .QN(n274)
         );
  DFFSSRX1_HVT sram_raddr_a5_reg_2_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_a5[2]), .CLK(net25643), .Q(sram_raddr_a5[2]), .QN(n360)
         );
  DFFSSRX1_HVT sram_raddr_a5_reg_1_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_a5[1]), .CLK(net25643), .Q(sram_raddr_a5[1]) );
  DFFSSRX1_HVT sram_raddr_a5_reg_0_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_a5[0]), .CLK(net25643), .Q(sram_raddr_a5[0]), .QN(n416)
         );
  DFFSSRX1_HVT sram_raddr_a6_reg_9_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_raddr_a6[9]), .CLK(net26973), .Q(sram_raddr_a6[9]) );
  DFFSSRX1_HVT sram_raddr_a6_reg_8_ ( .D(1'b0), .SETB(n211), .RSTB(
        n_sram_raddr_a6[8]), .CLK(net26973), .Q(sram_raddr_a6[8]) );
  DFFSSRX1_HVT sram_raddr_a6_reg_7_ ( .D(1'b0), .SETB(n209), .RSTB(
        n_sram_raddr_a6[7]), .CLK(net26973), .Q(sram_raddr_a6[7]) );
  DFFSSRX1_HVT sram_raddr_a6_reg_6_ ( .D(1'b0), .SETB(n184), .RSTB(
        n_sram_raddr_a6[6]), .CLK(net26973), .Q(sram_raddr_a6[6]), .QN(n464)
         );
  DFFSSRX1_HVT sram_raddr_a6_reg_5_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_a6[5]), .CLK(net26973), .Q(sram_raddr_a6[5]) );
  DFFSSRX1_HVT sram_raddr_a6_reg_4_ ( .D(1'b0), .SETB(n198), .RSTB(
        n_sram_raddr_a6[4]), .CLK(net26973), .Q(sram_raddr_a6[4]) );
  DFFSSRX1_HVT sram_raddr_a6_reg_3_ ( .D(1'b0), .SETB(n193), .RSTB(
        n_sram_raddr_a6[3]), .CLK(net26973), .Q(sram_raddr_a6[3]) );
  DFFSSRX1_HVT sram_raddr_a6_reg_2_ ( .D(1'b0), .SETB(n201), .RSTB(
        n_sram_raddr_a6[2]), .CLK(net26973), .Q(sram_raddr_a6[2]), .QN(n456)
         );
  DFFSSRX1_HVT sram_raddr_a6_reg_1_ ( .D(1'b0), .SETB(n195), .RSTB(
        n_sram_raddr_a6[1]), .CLK(net26973), .Q(sram_raddr_a6[1]) );
  DFFSSRX1_HVT sram_raddr_a6_reg_0_ ( .D(1'b0), .SETB(n212), .RSTB(
        n_sram_raddr_a6[0]), .CLK(net26973), .Q(sram_raddr_a6[0]), .QN(n306)
         );
  DFFSSRX1_HVT sram_raddr_b7_reg_9_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_b7[9]), .CLK(net27507), .Q(sram_raddr_b7[9]), .QN(n405)
         );
  DFFSSRX1_HVT sram_raddr_b7_reg_8_ ( .D(1'b0), .SETB(n169), .RSTB(
        n_sram_raddr_b7[8]), .CLK(net27507), .Q(sram_raddr_b7[8]), .QN(n353)
         );
  DFFSSRX1_HVT sram_raddr_b7_reg_7_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_b7[7]), .CLK(net27507), .Q(sram_raddr_b7[7]), .QN(n330)
         );
  DFFSSRX1_HVT sram_raddr_b7_reg_6_ ( .D(1'b0), .SETB(n199), .RSTB(
        n_sram_raddr_b7[6]), .CLK(net27507), .Q(sram_raddr_b7[6]) );
  DFFSSRX1_HVT sram_raddr_b7_reg_5_ ( .D(1'b0), .SETB(n194), .RSTB(
        n_sram_raddr_b7[5]), .CLK(net27507), .Q(sram_raddr_b7[5]), .QN(n340)
         );
  DFFSSRX1_HVT sram_raddr_b7_reg_4_ ( .D(1'b0), .SETB(n202), .RSTB(
        n_sram_raddr_b7[4]), .CLK(net27507), .Q(sram_raddr_b7[4]), .QN(n277)
         );
  DFFSSRX1_HVT sram_raddr_b7_reg_3_ ( .D(1'b0), .SETB(n196), .RSTB(
        n_sram_raddr_b7[3]), .CLK(net27507), .Q(sram_raddr_b7[3]), .QN(n347)
         );
  DFFSSRX1_HVT sram_raddr_b7_reg_2_ ( .D(1'b0), .SETB(n211), .RSTB(
        n_sram_raddr_b7[2]), .CLK(net27507), .Q(sram_raddr_b7[2]), .QN(n243)
         );
  DFFSSRX1_HVT sram_raddr_b7_reg_1_ ( .D(1'b0), .SETB(n209), .RSTB(
        n_sram_raddr_b7[1]), .CLK(net27507), .Q(sram_raddr_b7[1]) );
  DFFSSRX1_HVT sram_raddr_b7_reg_0_ ( .D(1'b0), .SETB(n169), .RSTB(
        n_sram_raddr_b7[0]), .CLK(net27507), .Q(sram_raddr_b7[0]), .QN(n419)
         );
  DFFSSRX1_HVT sram_raddr_b8_reg_9_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_b8[9]), .CLK(net28022), .Q(sram_raddr_b8[9]), .QN(n407)
         );
  DFFSSRX1_HVT sram_raddr_b8_reg_8_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_b8[8]), .CLK(net28022), .Q(sram_raddr_b8[8]), .QN(n337)
         );
  DFFSSRX1_HVT sram_raddr_b8_reg_7_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_b8[7]), .CLK(net28022), .Q(sram_raddr_b8[7]), .QN(n269)
         );
  DFFSSRX1_HVT sram_raddr_b8_reg_6_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_b8[6]), .CLK(net28022), .Q(sram_raddr_b8[6]) );
  DFFSSRX1_HVT sram_raddr_b8_reg_5_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_raddr_b8[5]), .CLK(net28022), .Q(sram_raddr_b8[5]), .QN(n325)
         );
  DFFSSRX1_HVT sram_raddr_b8_reg_4_ ( .D(1'b0), .SETB(n212), .RSTB(
        n_sram_raddr_b8[4]), .CLK(net28022), .Q(sram_raddr_b8[4]), .QN(n346)
         );
  DFFSSRX1_HVT sram_raddr_b8_reg_3_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_b8[3]), .CLK(net28022), .Q(sram_raddr_b8[3]), .QN(n282)
         );
  DFFSSRX1_HVT sram_raddr_b8_reg_2_ ( .D(1'b0), .SETB(n169), .RSTB(
        n_sram_raddr_b8[2]), .CLK(net28022), .Q(sram_raddr_b8[2]), .QN(n245)
         );
  DFFSSRX1_HVT sram_raddr_b8_reg_1_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_b8[1]), .CLK(net28022), .Q(sram_raddr_b8[1]) );
  DFFSSRX1_HVT sram_raddr_b8_reg_0_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_b8[0]), .CLK(net28022), .Q(sram_raddr_b8[0]), .QN(n420)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_9_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_b0[9]), .CLK(net28537), .Q(sram_raddr_b0[9]), .QN(n423)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_8_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_b0[8]), .CLK(net28537), .Q(sram_raddr_b0[8]), .QN(n329)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_7_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_raddr_b0[7]), .CLK(net28537), .Q(sram_raddr_b0[7]), .QN(n263)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_6_ ( .D(1'b0), .SETB(n211), .RSTB(
        n_sram_raddr_b0[6]), .CLK(net28537), .Q(sram_raddr_b0[6]), .QN(n391)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_5_ ( .D(1'b0), .SETB(n209), .RSTB(
        n_sram_raddr_b0[5]), .CLK(net28537), .Q(sram_raddr_b0[5]), .QN(n272)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_4_ ( .D(1'b0), .SETB(n169), .RSTB(
        n_sram_raddr_b0[4]), .CLK(net28537), .Q(sram_raddr_b0[4]), .QN(n323)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_3_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_b0[3]), .CLK(net28537), .Q(sram_raddr_b0[3]), .QN(n411)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_2_ ( .D(1'b0), .SETB(n198), .RSTB(
        n_sram_raddr_b0[2]), .CLK(net28537), .Q(sram_raddr_b0[2]), .QN(n279)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_1_ ( .D(1'b0), .SETB(n193), .RSTB(
        n_sram_raddr_b0[1]), .CLK(net28537), .Q(sram_raddr_b0[1]), .QN(n364)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_0_ ( .D(1'b0), .SETB(n201), .RSTB(
        n_sram_raddr_b0[0]), .CLK(net28537), .Q(sram_raddr_b0[0]), .QN(n250)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_9_ ( .D(1'b0), .SETB(n195), .RSTB(
        n_sram_raddr_b1[9]), .CLK(net29052), .Q(sram_raddr_b1[9]), .QN(n409)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_8_ ( .D(1'b0), .SETB(n212), .RSTB(
        n_sram_raddr_b1[8]), .CLK(net29052), .Q(sram_raddr_b1[8]), .QN(n267)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_7_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_b1[7]), .CLK(net29052), .Q(sram_raddr_b1[7]), .QN(n317)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_6_ ( .D(1'b0), .SETB(n169), .RSTB(
        n_sram_raddr_b1[6]), .CLK(net29052), .Q(sram_raddr_b1[6]), .QN(n327)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_5_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_b1[5]), .CLK(net29052), .Q(sram_raddr_b1[5]), .QN(n265)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_4_ ( .D(1'b0), .SETB(n199), .RSTB(
        n_sram_raddr_b1[4]), .CLK(net29052), .Q(sram_raddr_b1[4]), .QN(n335)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_3_ ( .D(1'b0), .SETB(n194), .RSTB(
        n_sram_raddr_b1[3]), .CLK(net29052), .Q(sram_raddr_b1[3]), .QN(n414)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_2_ ( .D(1'b0), .SETB(n202), .RSTB(
        n_sram_raddr_b1[2]), .CLK(net29052), .Q(sram_raddr_b1[2]), .QN(n273)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_1_ ( .D(1'b0), .SETB(n196), .RSTB(
        n_sram_raddr_b1[1]), .CLK(net29052), .Q(sram_raddr_b1[1]), .QN(n365)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_0_ ( .D(1'b0), .SETB(n211), .RSTB(
        n_sram_raddr_b1[0]), .CLK(net29052), .Q(sram_raddr_b1[0]), .QN(n251)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_9_ ( .D(1'b0), .SETB(n209), .RSTB(
        n_sram_raddr_b2[9]), .CLK(net29567), .Q(sram_raddr_b2[9]), .QN(n434)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_8_ ( .D(1'b0), .SETB(n169), .RSTB(
        n_sram_raddr_b2[8]), .CLK(net29567), .Q(sram_raddr_b2[8]), .QN(n401)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_7_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_b2[7]), .CLK(net29567), .Q(sram_raddr_b2[7]), .QN(n260)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_6_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_b2[6]), .CLK(net29567), .Q(sram_raddr_b2[6]), .QN(n390)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_5_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_b2[5]), .CLK(net29567), .Q(sram_raddr_b2[5]), .QN(n318)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_4_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_b2[4]), .CLK(net29567), .Q(sram_raddr_b2[4]), .QN(n264)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_3_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_raddr_b2[3]), .CLK(net29567), .Q(sram_raddr_b2[3]), .QN(n426)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_2_ ( .D(1'b0), .SETB(n212), .RSTB(
        n_sram_raddr_b2[2]), .CLK(net29567), .Q(sram_raddr_b2[2]), .QN(n334)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_1_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_b2[1]), .CLK(net29567), .Q(sram_raddr_b2[1]), .QN(n370)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_0_ ( .D(1'b0), .SETB(n169), .RSTB(
        n_sram_raddr_b2[0]), .CLK(net29567), .Q(sram_raddr_b2[0]), .QN(n287)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_9_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_b3[9]), .CLK(net30082), .Q(sram_raddr_b3[9]), .QN(n402)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_8_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_b3[8]), .CLK(net30082), .Q(sram_raddr_b3[8]), .QN(n268)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_7_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_b3[7]), .CLK(net30082), .Q(sram_raddr_b3[7]), .QN(n350)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_6_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_b3[6]), .CLK(net30082), .Q(sram_raddr_b3[6]), .QN(n400)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_5_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_raddr_b3[5]), .CLK(net30082), .Q(sram_raddr_b3[5]), .QN(n261)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_4_ ( .D(1'b0), .SETB(n211), .RSTB(
        n_sram_raddr_b3[4]), .CLK(net30082), .Q(sram_raddr_b3[4]), .QN(n320)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_3_ ( .D(1'b0), .SETB(n209), .RSTB(
        n_sram_raddr_b3[3]), .CLK(net30082), .Q(sram_raddr_b3[3]), .QN(n393)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_2_ ( .D(1'b0), .SETB(n187), .RSTB(
        n_sram_raddr_b3[2]), .CLK(net30082), .Q(sram_raddr_b3[2]), .QN(n326)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_1_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_b3[1]), .CLK(net30082), .Q(sram_raddr_b3[1]), .QN(n367)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_0_ ( .D(1'b0), .SETB(n198), .RSTB(
        n_sram_raddr_b3[0]), .CLK(net30082), .Q(sram_raddr_b3[0]), .QN(n285)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_9_ ( .D(1'b0), .SETB(n193), .RSTB(
        n_sram_raddr_b4[9]), .CLK(net30597), .Q(sram_raddr_b4[9]), .QN(n395)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_8_ ( .D(1'b0), .SETB(n201), .RSTB(
        n_sram_raddr_b4[8]), .CLK(net30597), .Q(sram_raddr_b4[8]), .QN(n328)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_7_ ( .D(1'b0), .SETB(n195), .RSTB(
        n_sram_raddr_b4[7]), .CLK(net30597), .Q(sram_raddr_b4[7]), .QN(n316)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_6_ ( .D(1'b0), .SETB(n212), .RSTB(
        n_sram_raddr_b4[6]), .CLK(net30597), .Q(sram_raddr_b4[6]), .QN(n415)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_5_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_b4[5]), .CLK(net30597), .Q(sram_raddr_b4[5]), .QN(n271)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_4_ ( .D(1'b0), .SETB(n187), .RSTB(
        n_sram_raddr_b4[4]), .CLK(net30597), .Q(sram_raddr_b4[4]), .QN(n336)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_3_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_b4[3]), .CLK(net30597), .Q(sram_raddr_b4[3]), .QN(n389)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_2_ ( .D(1'b0), .SETB(n199), .RSTB(
        n_sram_raddr_b4[2]), .CLK(net30597), .Q(sram_raddr_b4[2]), .QN(n322)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_1_ ( .D(1'b0), .SETB(n194), .RSTB(
        n_sram_raddr_b4[1]), .CLK(net30597), .Q(sram_raddr_b4[1]), .QN(n372)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_0_ ( .D(1'b0), .SETB(n202), .RSTB(
        n_sram_raddr_b4[0]), .CLK(net30597), .Q(sram_raddr_b4[0]), .QN(n286)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_9_ ( .D(1'b0), .SETB(n196), .RSTB(
        n_sram_raddr_b5[9]), .CLK(net31112), .Q(sram_raddr_b5[9]), .QN(n394)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_8_ ( .D(1'b0), .SETB(n211), .RSTB(
        n_sram_raddr_b5[8]), .CLK(net31112), .Q(sram_raddr_b5[8]), .QN(n281)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_7_ ( .D(1'b0), .SETB(n209), .RSTB(
        n_sram_raddr_b5[7]), .CLK(net31112), .Q(sram_raddr_b5[7]), .QN(n354)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_6_ ( .D(1'b0), .SETB(n187), .RSTB(
        n_sram_raddr_b5[6]), .CLK(net31112), .Q(sram_raddr_b5[6]), .QN(n404)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_5_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_b5[5]), .CLK(net31112), .Q(sram_raddr_b5[5]), .QN(n266)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_4_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_b5[4]), .CLK(net31112), .Q(sram_raddr_b5[4]), .QN(n324)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_3_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_b5[3]), .CLK(net31112), .Q(sram_raddr_b5[3]), .QN(n413)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_2_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_b5[2]), .CLK(net31112), .Q(sram_raddr_b5[2]), .QN(n321)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_1_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_raddr_b5[1]), .CLK(net31112), .Q(sram_raddr_b5[1]), .QN(n373)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_0_ ( .D(1'b0), .SETB(n187), .RSTB(
        n_sram_raddr_b5[0]), .CLK(net31112), .Q(sram_raddr_b5[0]), .QN(n252)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_9_ ( .D(1'b0), .SETB(n184), .RSTB(
        n_sram_raddr_b6[9]), .CLK(net31627), .Q(sram_raddr_b6[9]), .QN(n406)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_8_ ( .D(1'b0), .SETB(n187), .RSTB(
        n_sram_raddr_b6[8]), .CLK(net31627), .Q(sram_raddr_b6[8]), .QN(n388)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_7_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_b6[7]), .CLK(net31627), .Q(sram_raddr_b6[7]), .QN(n270)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_6_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_b6[6]), .CLK(net31627), .Q(sram_raddr_b6[6]), .QN(n427)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_5_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_b6[5]), .CLK(net31627), .Q(sram_raddr_b6[5]), .QN(n339)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_4_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_b6[4]), .CLK(net31627), .Q(sram_raddr_b6[4]), .QN(n276)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_3_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_raddr_b6[3]), .CLK(net31627), .Q(sram_raddr_b6[3]), .QN(n351)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_2_ ( .D(1'b0), .SETB(n169), .RSTB(
        n_sram_raddr_b6[2]), .CLK(net31627), .Q(sram_raddr_b6[2]), .QN(n242)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_1_ ( .D(1'b0), .SETB(n185), .RSTB(
        n_sram_raddr_b6[1]), .CLK(net31627), .Q(sram_raddr_b6[1]) );
  DFFSSRX1_HVT sram_raddr_b6_reg_0_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_b6[0]), .CLK(net31627), .Q(sram_raddr_b6[0]), .QN(n418)
         );
  DFFSSRX1_HVT sram_write_enable_b7_reg ( .D(n_sram_write_enable_b7), .SETB(
        n197), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b7) );
  DFFSSRX1_HVT sram_write_enable_b8_reg ( .D(n_sram_write_enable_b8), .SETB(
        n182), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b8) );
  DFFSSRX1_HVT sram_write_enable_b0_reg ( .D(n_sram_write_enable_b0), .SETB(
        n183), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b0) );
  DFFSSRX1_HVT sram_write_enable_b1_reg ( .D(n_sram_write_enable_b1), .SETB(
        n182), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b1) );
  DFFSSRX1_HVT sram_write_enable_b2_reg ( .D(n_sram_write_enable_b2), .SETB(
        n231), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b2) );
  DFFSSRX1_HVT sram_write_enable_b3_reg ( .D(n_sram_write_enable_b3), .SETB(
        n183), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b3) );
  DFFSSRX1_HVT sram_write_enable_b4_reg ( .D(n_sram_write_enable_b4), .SETB(
        n182), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b4) );
  DFFSSRX1_HVT sram_write_enable_b5_reg ( .D(n_sram_write_enable_b5), .SETB(
        n231), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b5) );
  DFFSSRX1_HVT sram_write_enable_b6_reg ( .D(n_sram_write_enable_b6), .SETB(
        n183), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b6) );
  DFFSSRX1_HVT sram_write_enable_d3_reg ( .D(n_sram_write_enable_d3), .SETB(
        n182), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_d3) );
  DFFSSRX1_HVT sram_write_enable_d4_reg ( .D(n_sram_write_enable_d4), .SETB(
        n231), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_d4) );
  DFFSSRX1_HVT sram_write_enable_c0_reg ( .D(n_sram_write_enable_c0), .SETB(
        n183), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_c0) );
  DFFSSRX1_HVT sram_write_enable_c1_reg ( .D(n_sram_write_enable_c1), .SETB(
        n182), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_c1) );
  DFFSSRX1_HVT sram_write_enable_c2_reg ( .D(n_sram_write_enable_c2), .SETB(
        n231), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_c2) );
  DFFSSRX1_HVT sram_write_enable_c3_reg ( .D(n_sram_write_enable_c3), .SETB(
        n183), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_c3) );
  DFFSSRX1_HVT sram_write_enable_c4_reg ( .D(n_sram_write_enable_c4), .SETB(
        n182), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_c4) );
  DFFSSRX1_HVT sram_write_enable_d0_reg ( .D(n_sram_write_enable_d0), .SETB(
        n231), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_d0) );
  DFFSSRX1_HVT sram_write_enable_d1_reg ( .D(n_sram_write_enable_d1), .SETB(
        n182), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_d1) );
  DFFSSRX1_HVT sram_write_enable_d2_reg ( .D(n_sram_write_enable_d2), .SETB(
        n231), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_d2) );
  DFFSSRX1_HVT state_reg_2_ ( .D(1'b0), .SETB(n186), .RSTB(n_state[2]), .CLK(
        clk), .Q(state[2]), .QN(n1024) );
  DFFSSRX1_HVT state_reg_3_ ( .D(1'b0), .SETB(n169), .RSTB(n_state[3]), .CLK(
        clk), .Q(state[3]), .QN(n1023) );
  AO221X1_HVT U3 ( .A1(1'b1), .A2(n1487), .A3(n1489), .A4(n408), .A5(n155), 
        .Y(n157) );
  AO221X1_HVT U4 ( .A1(1'b1), .A2(n1928), .A3(n1925), .A4(n167), .A5(n149), 
        .Y(n_sram_raddr_a4[8]) );
  AO221X1_HVT U5 ( .A1(1'b1), .A2(n1493), .A3(n1495), .A4(n344), .A5(n141), 
        .Y(n142) );
  AO221X1_HVT U6 ( .A1(1'b1), .A2(n905), .A3(n918), .A4(n273), .A5(n132), .Y(
        n1183) );
  AO221X1_HVT U7 ( .A1(1'b1), .A2(n1501), .A3(n428), .A4(n1502), .A5(n126), 
        .Y(n128) );
  AO221X1_HVT U8 ( .A1(1'b1), .A2(n1637), .A3(n450), .A4(n310), .A5(n120), .Y(
        n122) );
  AO222X1_HVT U9 ( .A1(sram_raddr_b8[7]), .A2(n234), .A3(n68), .A4(n1316), 
        .A5(1'b1), .A6(n74), .Y(n_sram_raddr_b8[7]) );
  AO221X1_HVT U10 ( .A1(1'b1), .A2(n1434), .A3(n358), .A4(n112), .A5(n113), 
        .Y(n115) );
  AO221X1_HVT U11 ( .A1(1'b1), .A2(n1883), .A3(n1880), .A4(n1838), .A5(n109), 
        .Y(n_sram_raddr_a3[8]) );
  AO221X1_HVT U12 ( .A1(1'b1), .A2(n1923), .A3(n1922), .A4(n167), .A5(n101), 
        .Y(n_sram_raddr_a4[7]) );
  AO222X1_HVT U13 ( .A1(sram_raddr_b7[7]), .A2(n233), .A3(n91), .A4(n1231), 
        .A5(1'b1), .A6(n96), .Y(n_sram_raddr_b7[7]) );
  AO222X1_HVT U14 ( .A1(sram_raddr_b7[5]), .A2(n232), .A3(n77), .A4(n1219), 
        .A5(1'b1), .A6(n83), .Y(n_sram_raddr_b7[5]) );
  AO221X1_HVT U15 ( .A1(1'b1), .A2(n402), .A3(n268), .A4(n880), .A5(n1158), 
        .Y(n62) );
  AO221X1_HVT U16 ( .A1(1'b1), .A2(n48), .A3(n1336), .A4(n1308), .A5(n51), .Y(
        n53) );
  AO22X1_HVT U17 ( .A1(n325), .A2(n1304), .A3(n1309), .A4(1'b1), .Y(n38) );
  OA221X1_HVT U18 ( .A1(1'b0), .A2(n1566), .A3(n1565), .A4(col[2]), .A5(n1564), 
        .Y(net22644) );
  OA221X1_HVT U19 ( .A1(1'b0), .A2(n539), .A3(row[2]), .A4(n538), .A5(n537), 
        .Y(n_row[2]) );
  OA221X1_HVT U20 ( .A1(1'b0), .A2(n1549), .A3(channel_cnt[1]), .A4(
        channel_cnt[0]), .A5(n1548), .Y(net22937) );
  OA221X1_HVT U21 ( .A1(1'b0), .A2(sram_raddr_weight[13]), .A3(
        sram_raddr_weight[12]), .A4(n1405), .A5(n203), .Y(n162) );
  OA221X1_HVT U22 ( .A1(1'b0), .A2(n1556), .A3(addr_change[0]), .A4(
        addr_change[1]), .A5(n1555), .Y(net22949) );
  OA221X1_HVT U23 ( .A1(1'b0), .A2(n1543), .A3(n1531), .A4(
        delay1_sram_waddr_d[8]), .A5(n1530), .Y(net22918) );
  OA221X1_HVT U24 ( .A1(1'b0), .A2(n1260), .A3(sram_raddr_b1[6]), .A4(n933), 
        .A5(n942), .Y(n1224) );
  OA221X1_HVT U25 ( .A1(1'b0), .A2(n192), .A3(sram_raddr_b8[3]), .A4(n1275), 
        .A5(n1274), .Y(n997) );
  OA221X1_HVT U26 ( .A1(1'b0), .A2(n1556), .A3(addr_change[2]), .A4(n138), 
        .A5(n1554), .Y(net22948) );
  OA221X1_HVT U27 ( .A1(1'b0), .A2(n1543), .A3(n1533), .A4(
        delay1_sram_waddr_d[7]), .A5(n1532), .Y(net22919) );
  OA221X1_HVT U28 ( .A1(1'b0), .A2(n1556), .A3(addr_change[3]), .A4(n124), 
        .A5(n1553), .Y(net22947) );
  OA221X1_HVT U29 ( .A1(1'b0), .A2(n1543), .A3(n1535), .A4(
        delay1_sram_waddr_d[6]), .A5(n1534), .Y(net22920) );
  OA21X1_HVT U30 ( .A1(n1317), .A2(sram_raddr_b8[7]), .A3(n224), .Y(n68) );
  OA221X1_HVT U31 ( .A1(1'b0), .A2(n1469), .A3(n249), .A4(n289), .A5(n357), 
        .Y(n117) );
  OA221X1_HVT U32 ( .A1(1'b0), .A2(n1543), .A3(n1537), .A4(
        delay1_sram_waddr_d[5]), .A5(n1536), .Y(net22921) );
  OA221X1_HVT U33 ( .A1(1'b0), .A2(n1543), .A3(n1539), .A4(
        delay1_sram_waddr_d[4]), .A5(n1538), .Y(net22922) );
  OA21X1_HVT U34 ( .A1(n1232), .A2(sram_raddr_b7[7]), .A3(n179), .Y(n91) );
  OA221X1_HVT U35 ( .A1(1'b0), .A2(n1543), .A3(delay1_sram_waddr_d[3]), .A4(
        n98), .A5(n1540), .Y(net22923) );
  OA221X1_HVT U36 ( .A1(1'b0), .A2(n1543), .A3(delay1_sram_waddr_d[2]), .A4(
        n89), .A5(n1541), .Y(net22924) );
  OA21X1_HVT U37 ( .A1(n1213), .A2(sram_raddr_b7[5]), .A3(n225), .Y(n77) );
  OA221X1_HVT U38 ( .A1(1'b0), .A2(n696), .A3(sram_raddr_b1[8]), .A4(n1366), 
        .A5(n1303), .Y(n701) );
  OA221X1_HVT U39 ( .A1(1'b0), .A2(n1543), .A3(delay1_sram_waddr_d[0]), .A4(
        delay1_sram_waddr_d[1]), .A5(n1542), .Y(net22925) );
  OA221X1_HVT U40 ( .A1(1'b0), .A2(n1303), .A3(sram_raddr_b4[8]), .A4(n1366), 
        .A5(n953), .Y(n977) );
  OA221X1_HVT U41 ( .A1(1'b0), .A2(n1527), .A3(n1515), .A4(
        delay1_sram_waddr_c[8]), .A5(n1514), .Y(net22902) );
  OA221X1_HVT U42 ( .A1(1'b0), .A2(n1168), .A3(sram_raddr_b3[9]), .A4(n883), 
        .A5(n62), .Y(n64) );
  OA221X1_HVT U43 ( .A1(1'b0), .A2(n64), .A3(n886), .A4(n885), .A5(n884), .Y(
        n65) );
  OA221X1_HVT U44 ( .A1(1'b0), .A2(n1527), .A3(n1517), .A4(
        delay1_sram_waddr_c[7]), .A5(n1516), .Y(net22903) );
  OA221X1_HVT U45 ( .A1(1'b0), .A2(n1527), .A3(n1519), .A4(
        delay1_sram_waddr_c[6]), .A5(n1518), .Y(net22904) );
  OA221X1_HVT U46 ( .A1(1'b0), .A2(n1527), .A3(n1521), .A4(
        delay1_sram_waddr_c[5]), .A5(n1520), .Y(net22905) );
  OA221X1_HVT U47 ( .A1(1'b0), .A2(n1527), .A3(n1523), .A4(
        delay1_sram_waddr_c[4]), .A5(n1522), .Y(net22906) );
  OA221X1_HVT U48 ( .A1(1'b0), .A2(n587), .A3(n323), .A4(n626), .A5(n29), .Y(
        n31) );
  OA221X1_HVT U49 ( .A1(1'b0), .A2(n1527), .A3(delay1_sram_waddr_c[3]), .A4(
        n28), .A5(n1524), .Y(net22907) );
  OA221X1_HVT U50 ( .A1(1'b0), .A2(n21), .A3(n173), .A4(n934), .A5(n938), .Y(
        n23) );
  OA221X1_HVT U51 ( .A1(1'b0), .A2(n1527), .A3(delay1_sram_waddr_c[2]), .A4(
        n17), .A5(n1525), .Y(net22908) );
  OA221X1_HVT U52 ( .A1(1'b0), .A2(n1527), .A3(delay1_sram_waddr_c[0]), .A4(
        delay1_sram_waddr_c[1]), .A5(n1526), .Y(net22909) );
  OA221X1_HVT U53 ( .A1(1'b0), .A2(n1302), .A3(n1025), .A4(n1299), .A5(n3), 
        .Y(n5) );
  OA221X1_HVT U54 ( .A1(1'b0), .A2(n5), .A3(n1071), .A4(n1015), .A5(n1014), 
        .Y(n6) );
  INVX1_HVT U55 ( .A(n1832), .Y(n172) );
  INVX1_HVT U56 ( .A(n1266), .Y(n168) );
  INVX1_HVT U57 ( .A(n1320), .Y(n173) );
  AO22X1_HVT U58 ( .A1(n266), .A2(n1016), .A3(sram_raddr_b5[5]), .A4(n1290), 
        .Y(n1) );
  AO21X1_HVT U59 ( .A1(n1013), .A2(n319), .A3(n1306), .Y(n2) );
  NAND2X0_HVT U60 ( .A1(n2), .A2(sram_raddr_b5[5]), .Y(n3) );
  OAI222X1_HVT U62 ( .A1(n1), .A2(n1366), .A3(n6), .A4(n221), .A5(n1303), .A6(
        n266), .Y(n_sram_raddr_b5[5]) );
  OA22X1_HVT U63 ( .A1(n644), .A2(n273), .A3(n899), .A4(n226), .Y(n7) );
  NAND3X0_HVT U64 ( .A1(n898), .A2(n646), .A3(n7), .Y(n8) );
  AO222X1_HVT U65 ( .A1(n8), .A2(n206), .A3(sram_raddr_b1[2]), .A4(n232), .A5(
        n273), .A6(n223), .Y(n_sram_raddr_b1[2]) );
  INVX0_HVT U67 ( .A(n664), .Y(n10) );
  OA221X1_HVT U68 ( .A1(n10), .A2(col[0]), .A3(n10), .A4(n707), .A5(n665), .Y(
        n11) );
  OA22X1_HVT U69 ( .A1(n265), .A2(n11), .A3(n929), .A4(n226), .Y(n12) );
  NAND3X0_HVT U70 ( .A1(n928), .A2(n670), .A3(n12), .Y(n13) );
  NAND2X0_HVT U71 ( .A1(n917), .A2(n265), .Y(n14) );
  AND2X1_HVT U72 ( .A1(n14), .A2(n673), .Y(n15) );
  AO222X1_HVT U73 ( .A1(n13), .A2(n1557), .A3(sram_raddr_b1[5]), .A4(n234), 
        .A5(n188), .A6(n15), .Y(n_sram_raddr_b1[5]) );
  INVX0_HVT U75 ( .A(n1526), .Y(n17) );
  AND2X1_HVT U76 ( .A1(n670), .A2(n215), .Y(n18) );
  AO222X1_HVT U77 ( .A1(n707), .A2(n676), .A3(n707), .A4(n1198), .A5(n676), 
        .A6(n675), .Y(n20) );
  OA22X1_HVT U78 ( .A1(n327), .A2(n18), .A3(sram_raddr_b1[6]), .A4(n20), .Y(
        n21) );
  OA22X1_HVT U80 ( .A1(n327), .A2(n1303), .A3(n23), .A4(n221), .Y(n24) );
  NAND2X0_HVT U81 ( .A1(n673), .A2(n327), .Y(n25) );
  NAND3X0_HVT U82 ( .A1(n25), .A2(n684), .A3(n179), .Y(n26) );
  NAND2X0_HVT U83 ( .A1(n24), .A2(n26), .Y(n_sram_raddr_b1[6]) );
  INVX0_HVT U85 ( .A(n1525), .Y(n28) );
  NAND2X0_HVT U86 ( .A1(n586), .A2(n1148), .Y(n29) );
  OA22X1_HVT U88 ( .A1(n272), .A2(n31), .A3(n838), .A4(n227), .Y(n32) );
  NAND3X0_HVT U89 ( .A1(n841), .A2(n594), .A3(n32), .Y(n33) );
  NAND2X0_HVT U90 ( .A1(n598), .A2(n272), .Y(n34) );
  AND2X1_HVT U91 ( .A1(n34), .A2(n597), .Y(n35) );
  AO222X1_HVT U92 ( .A1(n33), .A2(n1557), .A3(sram_raddr_b0[5]), .A4(n232), 
        .A5(n224), .A6(n35), .Y(n_sram_raddr_b0[5]) );
  INVX0_HVT U94 ( .A(n179), .Y(n37) );
  OA21X1_HVT U95 ( .A1(n1298), .A2(col[1]), .A3(n216), .Y(n39) );
  OA22X1_HVT U96 ( .A1(n325), .A2(n39), .A3(n1299), .A4(n1305), .Y(n40) );
  NAND2X0_HVT U97 ( .A1(n1336), .A2(n1300), .Y(n41) );
  AO221X1_HVT U98 ( .A1(n1310), .A2(n1301), .A3(n1310), .A4(n266), .A5(n227), 
        .Y(n42) );
  AND4X1_HVT U99 ( .A1(n40), .A2(n1302), .A3(n41), .A4(n42), .Y(n43) );
  OAI222X1_HVT U100 ( .A1(n37), .A2(n38), .A3(n43), .A4(n221), .A5(n325), .A6(
        n1303), .Y(n_sram_raddr_b8[5]) );
  AND2X1_HVT U104 ( .A1(n1322), .A2(n1318), .Y(n47) );
  AO222X1_HVT U105 ( .A1(n47), .A2(sram_raddr_b8[6]), .A3(n47), .A4(n1305), 
        .A5(sram_raddr_b8[6]), .A6(n1306), .Y(n48) );
  INVX0_HVT U106 ( .A(n1310), .Y(n49) );
  AO221X1_HVT U107 ( .A1(n1310), .A2(sram_raddr_b5[6]), .A3(n49), .A4(n404), 
        .A5(n227), .Y(n50) );
  NAND2X0_HVT U108 ( .A1(n1307), .A2(n50), .Y(n51) );
  OR2X1_HVT U110 ( .A1(sram_raddr_b8[6]), .A2(n1309), .Y(n54) );
  AND2X1_HVT U111 ( .A1(n224), .A2(n1314), .Y(n55) );
  AO222X1_HVT U112 ( .A1(n53), .A2(n206), .A3(n54), .A4(n55), .A5(n233), .A6(
        sram_raddr_b8[6]), .Y(n_sram_raddr_b8[6]) );
  NAND4X0_HVT U114 ( .A1(row[0]), .A2(col[2]), .A3(row[1]), .A4(col[3]), .Y(
        n57) );
  NAND3X0_HVT U115 ( .A1(row[0]), .A2(n235), .A3(n532), .Y(n58) );
  NAND3X0_HVT U116 ( .A1(n531), .A2(n57), .A3(n58), .Y(n59) );
  AO221X1_HVT U117 ( .A1(n59), .A2(n259), .A3(n59), .A4(n550), .A5(n1570), .Y(
        n60) );
  NAND3X0_HVT U118 ( .A1(row[3]), .A2(n537), .A3(n60), .Y(n533) );
  OA22X1_HVT U121 ( .A1(n402), .A2(n887), .A3(n65), .A4(n221), .Y(n66) );
  NAND4X0_HVT U122 ( .A1(n402), .A2(n888), .A3(sram_raddr_b3[8]), .A4(
        sram_raddr_b3[7]), .Y(n67) );
  NAND2X0_HVT U123 ( .A1(n66), .A2(n67), .Y(n_sram_raddr_b3[9]) );
  OA21X1_HVT U124 ( .A1(n354), .A2(n1311), .A3(n1319), .Y(n69) );
  AO22X1_HVT U125 ( .A1(n1322), .A2(n215), .A3(n213), .A4(col[1]), .Y(n70) );
  OA22X1_HVT U126 ( .A1(n173), .A2(n69), .A3(n269), .A4(n70), .Y(n71) );
  NAND3X0_HVT U127 ( .A1(n269), .A2(n1318), .A3(n1322), .Y(n72) );
  NAND3X0_HVT U128 ( .A1(n71), .A2(n1312), .A3(n72), .Y(n73) );
  OA221X1_HVT U129 ( .A1(n73), .A2(n1313), .A3(n73), .A4(n1336), .A5(n207), 
        .Y(n74) );
  OA21X1_HVT U132 ( .A1(n1210), .A2(n271), .A3(n1214), .Y(n78) );
  AO22X1_HVT U133 ( .A1(n1215), .A2(n214), .A3(n215), .A4(col[0]), .Y(n79) );
  OA22X1_HVT U134 ( .A1(n226), .A2(n78), .A3(n340), .A4(n79), .Y(n80) );
  NAND3X0_HVT U135 ( .A1(n340), .A2(n1226), .A3(n1215), .Y(n81) );
  NAND3X0_HVT U136 ( .A1(n80), .A2(n1211), .A3(n81), .Y(n82) );
  OA221X1_HVT U137 ( .A1(n82), .A2(n1212), .A3(n82), .A4(n1248), .A5(n205), 
        .Y(n83) );
  NAND4X0_HVT U140 ( .A1(state[0]), .A2(n1024), .A3(state[3]), .A4(n240), .Y(
        n86) );
  AO21X1_HVT U141 ( .A1(n1389), .A2(n86), .A3(n230), .Y(net22776) );
  INVX0_HVT U144 ( .A(n1542), .Y(n89) );
  OA21X1_HVT U145 ( .A1(n916), .A2(n918), .A3(n1260), .Y(n90) );
  OA21X1_HVT U146 ( .A1(sram_raddr_b1[3]), .A2(n905), .A3(n90), .Y(n1193) );
  OA21X1_HVT U147 ( .A1(n316), .A2(n1227), .A3(n1233), .Y(n92) );
  AO22X1_HVT U148 ( .A1(n1244), .A2(n213), .A3(n214), .A4(col[0]), .Y(n93) );
  OA22X1_HVT U149 ( .A1(n227), .A2(n92), .A3(n330), .A4(n93), .Y(n94) );
  NAND3X0_HVT U150 ( .A1(n1228), .A2(n94), .A3(n1235), .Y(n95) );
  OA221X1_HVT U151 ( .A1(n95), .A2(n1229), .A3(n95), .A4(n1248), .A5(n1557), 
        .Y(n96) );
  INVX0_HVT U153 ( .A(n1541), .Y(n98) );
  AO22X1_HVT U156 ( .A1(n1934), .A2(sram_raddr_a4[7]), .A3(n1803), .A4(n1797), 
        .Y(n101) );
  OA222X1_HVT U158 ( .A1(sram_raddr_weight[11]), .A2(sram_raddr_weight[9]), 
        .A3(sram_raddr_weight[11]), .A4(sram_raddr_weight[10]), .A5(
        sram_raddr_weight[11]), .A6(n1417), .Y(n103) );
  AND2X1_HVT U159 ( .A1(n1409), .A2(n1455), .Y(n104) );
  OA21X1_HVT U160 ( .A1(sram_raddr_weight[10]), .A2(n1412), .A3(
        sram_raddr_weight[11]), .Y(n105) );
  AO222X1_HVT U161 ( .A1(n103), .A2(n104), .A3(n105), .A4(n207), .A5(n1410), 
        .A6(n206), .Y(net22727) );
  NAND2X0_HVT U162 ( .A1(n669), .A2(n277), .Y(n106) );
  NAND2X0_HVT U163 ( .A1(n106), .A2(sram_raddr_b7[5]), .Y(n107) );
  NAND2X0_HVT U164 ( .A1(n107), .A2(n672), .Y(n1212) );
  AO22X1_HVT U166 ( .A1(n1887), .A2(sram_raddr_a3[8]), .A3(n1769), .A4(n1765), 
        .Y(n109) );
  AO221X1_HVT U168 ( .A1(n1433), .A2(n1439), .A3(n1433), .A4(n358), .A5(n228), 
        .Y(n111) );
  NAND2X0_HVT U169 ( .A1(sram_raddr_weight[5]), .A2(n1438), .Y(n112) );
  INVX0_HVT U170 ( .A(n1455), .Y(n113) );
  NAND3X0_HVT U172 ( .A1(n399), .A2(n111), .A3(n115), .Y(net22790) );
  OA21X1_HVT U174 ( .A1(write_row_conv1[2]), .A2(n1061), .A3(n117), .Y(n1347)
         );
  OA22X1_HVT U176 ( .A1(n450), .A2(n1892), .A3(n189), .A4(n1774), .Y(n119) );
  INVX0_HVT U177 ( .A(n1664), .Y(n120) );
  NAND3X0_HVT U179 ( .A1(n119), .A2(n1775), .A3(n122), .Y(n_sram_raddr_a1[1])
         );
  INVX0_HVT U181 ( .A(n1554), .Y(n124) );
  INVX0_HVT U183 ( .A(n1506), .Y(n126) );
  INVX0_HVT U185 ( .A(n1503), .Y(n129) );
  AO221X1_HVT U186 ( .A1(n1499), .A2(n428), .A3(n1499), .A4(n129), .A5(n1498), 
        .Y(n130) );
  NAND2X0_HVT U187 ( .A1(n128), .A2(n130), .Y(net22885) );
  AO21X1_HVT U188 ( .A1(channel_cnt[2]), .A2(n1547), .A3(channel_cnt[3]), .Y(
        n131) );
  AND3X1_HVT U189 ( .A1(n1549), .A2(n1546), .A3(n131), .Y(net22935) );
  INVX0_HVT U190 ( .A(n1260), .Y(n132) );
  NAND2X0_HVT U192 ( .A1(n1921), .A2(sram_raddr_a4[7]), .Y(n134) );
  NAND2X0_HVT U193 ( .A1(n1924), .A2(n134), .Y(n135) );
  AO222X1_HVT U194 ( .A1(n135), .A2(n1974), .A3(n1931), .A4(n1922), .A5(
        sram_raddr_a7[7]), .A6(n1934), .Y(n136) );
  OR2X1_HVT U195 ( .A1(n1923), .A2(n136), .Y(n_sram_raddr_a7[7]) );
  INVX0_HVT U197 ( .A(n1555), .Y(n138) );
  INVX0_HVT U200 ( .A(n1506), .Y(n141) );
  AO221X1_HVT U201 ( .A1(n1492), .A2(n344), .A3(n1492), .A4(n1494), .A5(n1498), 
        .Y(n143) );
  NAND2X0_HVT U202 ( .A1(n142), .A2(n143), .Y(net22879) );
  AOI22X1_HVT U203 ( .A1(n1995), .A2(n1997), .A3(n2001), .A4(n1996), .Y(n144)
         );
  OAI221X1_HVT U204 ( .A1(n144), .A2(n1995), .A3(n144), .A4(n1996), .A5(n1662), 
        .Y(n_box_sel_1_) );
  NAND2X0_HVT U205 ( .A1(n591), .A2(n276), .Y(n145) );
  NAND2X0_HVT U206 ( .A1(n145), .A2(sram_raddr_b6[5]), .Y(n146) );
  NAND2X0_HVT U207 ( .A1(n146), .A2(n593), .Y(n1121) );
  AO22X1_HVT U210 ( .A1(n1934), .A2(sram_raddr_a4[8]), .A3(n1803), .A4(n1799), 
        .Y(n149) );
  INVX0_HVT U212 ( .A(n1585), .Y(n151) );
  OR2X1_HVT U213 ( .A1(n1581), .A2(sram_raddr_a0[2]), .Y(n152) );
  AO222X1_HVT U214 ( .A1(n151), .A2(n152), .A3(n1974), .A4(n1738), .A5(n519), 
        .A6(n1851), .Y(n_sram_raddr_a0[2]) );
  INVX0_HVT U217 ( .A(n1506), .Y(n155) );
  AO221X1_HVT U219 ( .A1(n1486), .A2(n408), .A3(n1486), .A4(n1488), .A5(n1498), 
        .Y(n158) );
  NAND2X0_HVT U220 ( .A1(n157), .A2(n158), .Y(net22873) );
  INVX0_HVT U221 ( .A(n1403), .Y(n159) );
  OA221X1_HVT U222 ( .A1(sram_raddr_weight[13]), .A2(sram_raddr_weight[12]), 
        .A3(sram_raddr_weight[13]), .A4(n1406), .A5(n159), .Y(n160) );
  OR3X1_HVT U224 ( .A1(n1404), .A2(n160), .A3(n162), .Y(net22713) );
  AND3X1_HVT U228 ( .A1(n1382), .A2(weight_cnt[0]), .A3(weight_cnt[1]), .Y(
        n166) );
  OA21X1_HVT U229 ( .A1(n166), .A2(weight_cnt[2]), .A3(n1372), .Y(
        n_weight_cnt[2]) );
  INVX1_HVT U230 ( .A(n180), .Y(n181) );
  INVX2_HVT U231 ( .A(srstn), .Y(n180) );
  INVX1_HVT U232 ( .A(n189), .Y(n170) );
  INVX1_HVT U233 ( .A(n1942), .Y(n167) );
  INVX1_HVT U234 ( .A(n1846), .Y(n479) );
  NOR2X0_HVT U235 ( .A1(n1388), .A2(n1387), .Y(net22649) );
  INVX0_HVT U236 ( .A(n1935), .Y(n470) );
  INVX0_HVT U237 ( .A(n200), .Y(n184) );
  INVX1_HVT U238 ( .A(n212), .Y(n200) );
  INVX1_HVT U239 ( .A(n211), .Y(n197) );
  INVX0_HVT U240 ( .A(n1658), .Y(n1659) );
  INVX1_HVT U241 ( .A(n226), .Y(n178) );
  INVX2_HVT U242 ( .A(n231), .Y(n169) );
  NOR2X0_HVT U243 ( .A1(n1482), .A2(n1500), .Y(n1485) );
  INVX1_HVT U244 ( .A(n1669), .Y(n1670) );
  INVX0_HVT U245 ( .A(n1651), .Y(n1652) );
  INVX2_HVT U246 ( .A(n1974), .Y(n171) );
  NOR2X1_HVT U247 ( .A1(n396), .A2(n1713), .Y(n1725) );
  NOR2X1_HVT U248 ( .A1(n1879), .A2(sram_raddr_a3[8]), .Y(n1884) );
  INVX1_HVT U249 ( .A(n181), .Y(n229) );
  INVX1_HVT U250 ( .A(n181), .Y(n230) );
  NBUFFX2_HVT U251 ( .A(n181), .Y(n231) );
  INVX0_HVT U252 ( .A(n899), .Y(n900) );
  INVX1_HVT U253 ( .A(n674), .Y(n676) );
  INVX1_HVT U254 ( .A(n1109), .Y(n1107) );
  INVX1_HVT U255 ( .A(n1557), .Y(n228) );
  INVX1_HVT U256 ( .A(n1219), .Y(n1220) );
  INVX0_HVT U257 ( .A(n1916), .Y(n1920) );
  INVX1_HVT U258 ( .A(n1440), .Y(n1444) );
  INVX0_HVT U259 ( .A(n1806), .Y(n481) );
  INVX0_HVT U260 ( .A(n1772), .Y(n484) );
  AOI22X1_HVT U261 ( .A1(n1932), .A2(n1931), .A3(n170), .A4(n1930), .Y(n1933)
         );
  INVX0_HVT U262 ( .A(n1073), .Y(n1058) );
  INVX0_HVT U263 ( .A(n1405), .Y(n1410) );
  INVX0_HVT U264 ( .A(n887), .Y(n878) );
  INVX0_HVT U265 ( .A(n1727), .Y(n1728) );
  INVX0_HVT U266 ( .A(n1530), .Y(n1529) );
  INVX0_HVT U267 ( .A(n1514), .Y(n1513) );
  INVX0_HVT U268 ( .A(n1672), .Y(n1673) );
  INVX0_HVT U269 ( .A(n1620), .Y(n1621) );
  INVX0_HVT U270 ( .A(n997), .Y(n495) );
  INVX0_HVT U271 ( .A(n1889), .Y(n473) );
  INVX0_HVT U272 ( .A(n1723), .Y(n1724) );
  INVX0_HVT U273 ( .A(n701), .Y(n699) );
  INVX0_HVT U274 ( .A(n862), .Y(n863) );
  INVX1_HVT U275 ( .A(n228), .Y(n203) );
  INVX0_HVT U276 ( .A(n1457), .Y(n1443) );
  INVX0_HVT U277 ( .A(n1456), .Y(net22655) );
  INVX0_HVT U278 ( .A(n881), .Y(n882) );
  INVX0_HVT U279 ( .A(n1614), .Y(n1577) );
  INVX0_HVT U280 ( .A(n1622), .Y(n1623) );
  INVX0_HVT U281 ( .A(n1616), .Y(n1617) );
  INVX0_HVT U282 ( .A(n564), .Y(n565) );
  INVX0_HVT U283 ( .A(n1193), .Y(n908) );
  INVX0_HVT U284 ( .A(n968), .Y(n969) );
  INVX0_HVT U285 ( .A(n1164), .Y(n1165) );
  INVX0_HVT U286 ( .A(n1987), .Y(n1944) );
  INVX0_HVT U287 ( .A(n1666), .Y(n1668) );
  INVX0_HVT U288 ( .A(n1721), .Y(n1692) );
  INVX1_HVT U289 ( .A(n231), .Y(n196) );
  INVX1_HVT U290 ( .A(n200), .Y(n202) );
  INVX1_HVT U291 ( .A(n231), .Y(n187) );
  INVX1_HVT U292 ( .A(n197), .Y(n198) );
  INVX1_HVT U293 ( .A(n231), .Y(n193) );
  INVX1_HVT U294 ( .A(n200), .Y(n201) );
  INVX1_HVT U295 ( .A(n197), .Y(n194) );
  INVX1_HVT U296 ( .A(n231), .Y(n195) );
  INVX1_HVT U297 ( .A(n197), .Y(n185) );
  INVX1_HVT U298 ( .A(n197), .Y(n199) );
  INVX1_HVT U299 ( .A(n197), .Y(n186) );
  INVX0_HVT U300 ( .A(n1714), .Y(n1715) );
  INVX0_HVT U301 ( .A(n1368), .Y(n534) );
  INVX1_HVT U302 ( .A(n1259), .Y(n190) );
  INVX0_HVT U303 ( .A(n953), .Y(n950) );
  INVX1_HVT U304 ( .A(n1259), .Y(n192) );
  INVX0_HVT U305 ( .A(n929), .Y(n930) );
  INVX0_HVT U306 ( .A(n1065), .Y(n1066) );
  INVX1_HVT U307 ( .A(n1259), .Y(n191) );
  INVX0_HVT U308 ( .A(n1674), .Y(n1675) );
  INVX0_HVT U309 ( .A(n590), .Y(n582) );
  INVX0_HVT U310 ( .A(n750), .Y(n739) );
  INVX0_HVT U311 ( .A(n668), .Y(n660) );
  AND2X1_HVT U312 ( .A1(n1366), .A2(n1303), .Y(n1266) );
  INVX0_HVT U313 ( .A(n696), .Y(n686) );
  INVX1_HVT U314 ( .A(n222), .Y(n188) );
  INVX2_HVT U315 ( .A(n231), .Y(n174) );
  INVX2_HVT U316 ( .A(n200), .Y(n175) );
  INVX2_HVT U317 ( .A(n197), .Y(n176) );
  INVX2_HVT U318 ( .A(n197), .Y(n177) );
  INVX1_HVT U319 ( .A(n1974), .Y(n189) );
  INVX0_HVT U320 ( .A(n1332), .Y(n982) );
  INVX0_HVT U321 ( .A(n690), .Y(n708) );
  INVX0_HVT U322 ( .A(n1236), .Y(n891) );
  INVX1_HVT U323 ( .A(n228), .Y(n204) );
  INVX1_HVT U324 ( .A(n228), .Y(n207) );
  INVX0_HVT U325 ( .A(n1729), .Y(n1730) );
  INVX0_HVT U326 ( .A(n1941), .Y(n1981) );
  INVX0_HVT U327 ( .A(n1767), .Y(n1768) );
  INVX1_HVT U328 ( .A(n228), .Y(n205) );
  INVX0_HVT U329 ( .A(n1849), .Y(n1868) );
  INVX1_HVT U330 ( .A(n228), .Y(n206) );
  INVX1_HVT U331 ( .A(n1315), .Y(n233) );
  INVX0_HVT U332 ( .A(n1601), .Y(n1607) );
  INVX0_HVT U333 ( .A(n1913), .Y(n1915) );
  INVX0_HVT U334 ( .A(n1334), .Y(n1340) );
  INVX0_HVT U335 ( .A(n1801), .Y(n1802) );
  INVX1_HVT U336 ( .A(n1315), .Y(n232) );
  NOR2X0_HVT U337 ( .A1(conv1_weight_done), .A2(n1667), .Y(n1974) );
  INVX0_HVT U338 ( .A(n847), .Y(n849) );
  INVX0_HVT U339 ( .A(n1034), .Y(n1017) );
  INVX0_HVT U340 ( .A(n1764), .Y(n1766) );
  AND2X1_HVT U341 ( .A1(n1567), .A2(n254), .Y(n1832) );
  INVX0_HVT U342 ( .A(n1380), .Y(n1383) );
  INVX0_HVT U343 ( .A(n1568), .Y(n1679) );
  NOR2X1_HVT U344 ( .A1(n1924), .A2(sram_raddr_a4[8]), .Y(n1929) );
  INVX0_HVT U345 ( .A(n1137), .Y(n1126) );
  INVX0_HVT U346 ( .A(n1326), .Y(n1328) );
  NOR2X1_HVT U347 ( .A1(n333), .A2(n1649), .Y(n1660) );
  INVX0_HVT U348 ( .A(n583), .Y(n584) );
  INVX0_HVT U349 ( .A(n591), .Y(n580) );
  INVX0_HVT U350 ( .A(n1078), .Y(n1132) );
  INVX0_HVT U351 ( .A(n661), .Y(n662) );
  INVX0_HVT U352 ( .A(n1546), .Y(n1545) );
  INVX0_HVT U353 ( .A(n556), .Y(n549) );
  AOI22X1_HVT U354 ( .A1(sram_raddr_b7[6]), .A2(n1306), .A3(n1216), .A4(n1226), 
        .Y(n1217) );
  INVX0_HVT U355 ( .A(n740), .Y(n741) );
  INVX0_HVT U356 ( .A(n1999), .Y(n2002) );
  INVX0_HVT U357 ( .A(n1995), .Y(n1998) );
  INVX0_HVT U358 ( .A(n1089), .Y(n1090) );
  INVX0_HVT U359 ( .A(n1996), .Y(n524) );
  INVX0_HVT U360 ( .A(n1374), .Y(n1375) );
  INVX0_HVT U361 ( .A(n669), .Y(n658) );
  INVX0_HVT U362 ( .A(n924), .Y(n919) );
  INVX0_HVT U363 ( .A(n1507), .Y(n1470) );
  AND4X1_HVT U364 ( .A1(n552), .A2(row[0]), .A3(n551), .A4(n550), .Y(n1320) );
  INVX0_HVT U365 ( .A(n1951), .Y(n1956) );
  AND4X1_HVT U366 ( .A1(n552), .A2(n551), .A3(n349), .A4(n259), .Y(n1064) );
  INVX1_HVT U367 ( .A(n1366), .Y(n179) );
  INVX0_HVT U368 ( .A(n1025), .Y(n1026) );
  INVX0_HVT U369 ( .A(n1564), .Y(n1386) );
  INVX0_HVT U370 ( .A(n1782), .Y(n1783) );
  INVX0_HVT U371 ( .A(n797), .Y(n800) );
  INVX0_HVT U372 ( .A(n1631), .Y(n1632) );
  INVX0_HVT U373 ( .A(n647), .Y(n645) );
  INVX0_HVT U374 ( .A(n576), .Y(n722) );
  INVX0_HVT U375 ( .A(n1548), .Y(n1547) );
  INVX0_HVT U376 ( .A(n1748), .Y(n1749) );
  INVX0_HVT U377 ( .A(n1291), .Y(n1289) );
  INVX0_HVT U378 ( .A(n546), .Y(n552) );
  INVX0_HVT U379 ( .A(n1203), .Y(n1201) );
  INVX0_HVT U380 ( .A(n1580), .Y(n1579) );
  INVX0_HVT U381 ( .A(n1298), .Y(n1286) );
  INVX0_HVT U382 ( .A(n729), .Y(n723) );
  INVX0_HVT U383 ( .A(n1553), .Y(n1552) );
  INVX0_HVT U384 ( .A(n1578), .Y(n1582) );
  INVX0_HVT U385 ( .A(n1903), .Y(n1904) );
  INVX0_HVT U386 ( .A(n1857), .Y(n1858) );
  INVX0_HVT U387 ( .A(n732), .Y(n725) );
  INVX0_HVT U388 ( .A(n1471), .Y(n1473) );
  INVX0_HVT U389 ( .A(n1562), .Y(n1021) );
  INVX0_HVT U390 ( .A(mode[1]), .Y(n522) );
  AND4X1_HVT U391 ( .A1(state[1]), .A2(state[0]), .A3(n1023), .A4(state[2]), 
        .Y(n1557) );
  INVX1_HVT U392 ( .A(n180), .Y(n182) );
  INVX1_HVT U393 ( .A(n180), .Y(n183) );
  INVX2_HVT U394 ( .A(n197), .Y(n208) );
  INVX2_HVT U395 ( .A(n200), .Y(n210) );
  INVX2_HVT U396 ( .A(n200), .Y(n209) );
  INVX2_HVT U397 ( .A(n231), .Y(n212) );
  INVX2_HVT U398 ( .A(n231), .Y(n211) );
  NAND2X2_HVT U399 ( .A1(n554), .A2(n1355), .Y(n1455) );
  INVX1_HVT U400 ( .A(n1306), .Y(n213) );
  INVX1_HVT U401 ( .A(n1306), .Y(n214) );
  INVX2_HVT U402 ( .A(n1306), .Y(n215) );
  INVX2_HVT U403 ( .A(n1306), .Y(n216) );
  INVX1_HVT U404 ( .A(n1266), .Y(n217) );
  INVX1_HVT U405 ( .A(n1832), .Y(n218) );
  INVX1_HVT U406 ( .A(n1064), .Y(n219) );
  INVX1_HVT U407 ( .A(n1064), .Y(n220) );
  INVX1_HVT U408 ( .A(n1557), .Y(n221) );
  INVX1_HVT U409 ( .A(n179), .Y(n222) );
  INVX1_HVT U410 ( .A(n222), .Y(n223) );
  INVX1_HVT U411 ( .A(n222), .Y(n224) );
  INVX1_HVT U412 ( .A(n222), .Y(n225) );
  INVX1_HVT U413 ( .A(n1320), .Y(n226) );
  INVX1_HVT U414 ( .A(n1320), .Y(n227) );
  AND2X2_HVT U415 ( .A1(mode[1]), .A2(n521), .Y(n1354) );
  OAI21X1_HVT U416 ( .A1(n557), .A2(n556), .A3(n1544), .Y(n1315) );
  INVX0_HVT U417 ( .A(n1315), .Y(n234) );
  INVX1_HVT U418 ( .A(n1389), .Y(n2003) );
  INVX1_HVT U419 ( .A(n233), .Y(n1303) );
  OR2X1_HVT U420 ( .A1(n554), .A2(n555), .Y(n1366) );
  INVX1_HVT U421 ( .A(n1198), .Y(n1226) );
  INVX1_HVT U422 ( .A(n1945), .Y(n1989) );
  INVX1_HVT U423 ( .A(n218), .Y(n1896) );
  INVX1_HVT U424 ( .A(n219), .Y(n1260) );
  INVX1_HVT U425 ( .A(n1357), .Y(n1363) );
  NAND4X0_HVT U426 ( .A1(state[0]), .A2(state[1]), .A3(n1023), .A4(n1024), .Y(
        n1389) );
  INVX1_HVT U427 ( .A(n1299), .Y(n1318) );
  OA221X1_HVT U428 ( .A1(n1568), .A2(n1052), .A3(n1568), .A4(
        addr_col_sel_cnt[1]), .A5(n1559), .Y(n1945) );
  OAI21X1_HVT U429 ( .A1(n254), .A2(n1355), .A3(n1369), .Y(n_conv1_weight_done) );
  INVX1_HVT U430 ( .A(n1500), .Y(n1506) );
  INVX1_HVT U431 ( .A(n1455), .Y(n1465) );
  OAI21X1_HVT U432 ( .A1(n770), .A2(n269), .A3(n793), .Y(n1313) );
  OA221X1_HVT U433 ( .A1(n1568), .A2(n1052), .A3(n1568), .A4(n1051), .A5(n1559), .Y(n1759) );
  INVX1_HVT U434 ( .A(n554), .Y(n1549) );
  NAND3X0_HVT U435 ( .A1(n1024), .A2(n1445), .A3(state[3]), .Y(n554) );
  INVX1_HVT U436 ( .A(n542), .Y(n544) );
  INVX1_HVT U437 ( .A(n543), .Y(n545) );
  INVX1_HVT U438 ( .A(mem_sel), .Y(n1512) );
  INVX1_HVT U439 ( .A(n1798), .Y(n1800) );
  INVX1_HVT U440 ( .A(n1243), .Y(n1258) );
  INVX1_HVT U441 ( .A(n1331), .Y(n1346) );
  OAI21X1_HVT U442 ( .A1(n1274), .A2(n346), .A3(n751), .Y(n1287) );
  AO221X1_HVT U443 ( .A1(sram_raddr_b1[9]), .A2(n969), .A3(n409), .A4(n968), 
        .A5(n220), .Y(n1243) );
  OAI21X1_HVT U444 ( .A1(sram_raddr_a4[5]), .A2(n1642), .A3(n1649), .Y(n1786)
         );
  OAI21X1_HVT U445 ( .A1(n681), .A2(n330), .A3(n690), .Y(n1229) );
  OAI21X1_HVT U446 ( .A1(sram_raddr_a5[4]), .A2(n1693), .A3(n1699), .Y(n1816)
         );
  AO221X1_HVT U447 ( .A1(sram_raddr_b2[9]), .A2(n1066), .A3(n434), .A4(n1065), 
        .A5(n219), .Y(n1331) );
  OAI21X1_HVT U448 ( .A1(sram_raddr_b4[6]), .A2(n671), .A3(n680), .Y(n934) );
  OAI21X1_HVT U449 ( .A1(sram_raddr_a5[6]), .A2(n1706), .A3(n1713), .Y(n1825)
         );
  OAI21X1_HVT U450 ( .A1(n604), .A2(n270), .A3(n627), .Y(n1143) );
  AO22X1_HVT U451 ( .A1(write_row_conv1[0]), .A2(n1363), .A3(n1354), .A4(
        col_enable[1]), .Y(n542) );
  AO22X1_HVT U452 ( .A1(write_col_conv1[0]), .A2(n1363), .A3(n1354), .A4(
        col_enable[0]), .Y(n543) );
  AND2X1_HVT U453 ( .A1(n1528), .A2(mem_sel), .Y(n1543) );
  AND2X1_HVT U454 ( .A1(n1528), .A2(n1512), .Y(n1527) );
  INVX1_HVT U455 ( .A(n1498), .Y(n1505) );
  AO21X1_HVT U456 ( .A1(n1476), .A2(n1475), .A3(n1507), .Y(n1500) );
  AND4X1_HVT U457 ( .A1(n1569), .A2(n1053), .A3(n2003), .A4(n338), .Y(n1567)
         );
  INVX1_HVT U458 ( .A(n1361), .Y(n1544) );
  NAND2X0_HVT U459 ( .A1(channel_cnt[1]), .A2(channel_cnt[0]), .Y(n1548) );
  NAND3X0_HVT U460 ( .A1(n551), .A2(n256), .A3(n313), .Y(n556) );
  AND3X1_HVT U461 ( .A1(n1565), .A2(n241), .A3(n235), .Y(n551) );
  NAND2X0_HVT U462 ( .A1(row[1]), .A2(row[0]), .Y(n557) );
  INVX2_HVT U463 ( .A(n1759), .Y(n1887) );
  INVX2_HVT U464 ( .A(n1892), .Y(n1934) );
  INVX1_HVT U465 ( .A(n520), .Y(n1569) );
  NAND2X0_HVT U466 ( .A1(n1993), .A2(n254), .Y(n1568) );
  AND2X1_HVT U467 ( .A1(n2003), .A2(n520), .Y(n1993) );
  INVX1_HVT U468 ( .A(mode[0]), .Y(n521) );
  AND2X1_HVT U469 ( .A1(n1363), .A2(delay2_write_enable), .Y(n1469) );
  NAND2X0_HVT U470 ( .A1(mode[0]), .A2(n522), .Y(n1357) );
  NAND4X0_HVT U471 ( .A1(n1053), .A2(n1569), .A3(n2003), .A4(
        addr_row_sel_cnt[0]), .Y(n1667) );
  INVX1_HVT U472 ( .A(n1563), .Y(n1020) );
  NOR4X1_HVT U473 ( .A1(conv2_weight_cnt[7]), .A2(conv2_weight_cnt[6]), .A3(
        n528), .A4(n527), .Y(n_conv_done) );
  NOR4X1_HVT U474 ( .A1(conv1_weight_cnt[7]), .A2(conv1_weight_cnt[6]), .A3(
        conv1_weight_cnt[5]), .A4(n1357), .Y(n525) );
  NOR4X1_HVT U475 ( .A1(conv1_done), .A2(conv1_weight_cnt[1]), .A3(
        conv1_weight_cnt[0]), .A4(conv1_weight_cnt[3]), .Y(n526) );
  NOR4X1_HVT U476 ( .A1(channel_cnt[1]), .A2(channel_cnt[4]), .A3(
        conv2_weight_done), .A4(n529), .Y(n530) );
  INVX1_HVT U477 ( .A(n2000), .Y(n1994) );
  INVX1_HVT U478 ( .A(n1532), .Y(n1531) );
  INVX1_HVT U479 ( .A(n1534), .Y(n1533) );
  INVX1_HVT U480 ( .A(n1536), .Y(n1535) );
  INVX1_HVT U481 ( .A(n1538), .Y(n1537) );
  INVX1_HVT U482 ( .A(n1540), .Y(n1539) );
  INVX1_HVT U483 ( .A(n1516), .Y(n1515) );
  INVX1_HVT U484 ( .A(n1518), .Y(n1517) );
  INVX1_HVT U485 ( .A(n1520), .Y(n1519) );
  INVX1_HVT U486 ( .A(n1522), .Y(n1521) );
  INVX1_HVT U487 ( .A(n1524), .Y(n1523) );
  NOR4X1_HVT U488 ( .A1(delay1_sram_waddr_b[0]), .A2(delay1_sram_waddr_b[1]), 
        .A3(delay1_sram_waddr_b[2]), .A4(delay1_sram_waddr_b[3]), .Y(n1494) );
  INVX1_HVT U489 ( .A(n1388), .Y(n1566) );
  INVX1_HVT U490 ( .A(n1371), .Y(n1377) );
  INVX1_HVT U491 ( .A(n1803), .Y(n1794) );
  INVX1_HVT U492 ( .A(n1869), .Y(n1874) );
  INVX1_HVT U493 ( .A(n1628), .Y(n1629) );
  INVX1_HVT U494 ( .A(n977), .Y(n964) );
  INVX1_HVT U495 ( .A(n1843), .Y(n1830) );
  INVX1_HVT U496 ( .A(n1390), .Y(n1441) );
  INVX1_HVT U497 ( .A(n1838), .Y(n1942) );
  INVX1_HVT U498 ( .A(n1985), .Y(n1986) );
  INVX1_HVT U499 ( .A(n1973), .Y(n1975) );
  INVX1_HVT U500 ( .A(n1962), .Y(n1967) );
  INVX1_HVT U501 ( .A(n1841), .Y(n1842) );
  INVX1_HVT U502 ( .A(n1826), .Y(n1831) );
  INVX1_HVT U503 ( .A(n1817), .Y(n1821) );
  INVX1_HVT U504 ( .A(n1760), .Y(n1761) );
  INVX1_HVT U505 ( .A(n1769), .Y(n1758) );
  INVX1_HVT U506 ( .A(n1149), .Y(n1150) );
  INVX1_HVT U507 ( .A(n1145), .Y(n1147) );
  INVX1_HVT U508 ( .A(n1134), .Y(n1135) );
  INVX1_HVT U509 ( .A(n1230), .Y(n1232) );
  INVX1_HVT U510 ( .A(n1233), .Y(n1234) );
  INVX1_HVT U511 ( .A(n1246), .Y(n1252) );
  NAND2X0_HVT U512 ( .A1(n1259), .A2(n1174), .Y(n1248) );
  NAND2X0_HVT U513 ( .A1(n1259), .A2(n1078), .Y(n1162) );
  NAND2X0_HVT U514 ( .A1(n1259), .A2(n1326), .Y(n1336) );
  INVX1_HVT U515 ( .A(n955), .Y(n956) );
  INVX1_HVT U516 ( .A(n684), .Y(n697) );
  INVX1_HVT U517 ( .A(n693), .Y(n712) );
  INVX1_HVT U518 ( .A(n948), .Y(n954) );
  INVX1_HVT U519 ( .A(n932), .Y(n1202) );
  INVX1_HVT U520 ( .A(n897), .Y(n918) );
  INVX1_HVT U521 ( .A(n961), .Y(n974) );
  NAND2X0_HVT U522 ( .A1(col[1]), .A2(n213), .Y(n1332) );
  INVX1_HVT U523 ( .A(n1319), .Y(n1321) );
  INVX1_HVT U524 ( .A(n1314), .Y(n1317) );
  INVX1_HVT U525 ( .A(n1041), .Y(n1056) );
  INVX1_HVT U526 ( .A(n1016), .Y(n1290) );
  INVX1_HVT U527 ( .A(n1018), .Y(n1071) );
  INVX1_HVT U528 ( .A(n1005), .Y(n1003) );
  INVX1_HVT U529 ( .A(n844), .Y(n1108) );
  INVX1_HVT U530 ( .A(n864), .Y(n886) );
  INVX1_HVT U531 ( .A(n868), .Y(n869) );
  INVX1_HVT U532 ( .A(n830), .Y(n828) );
  INVX1_HVT U533 ( .A(n1084), .Y(n1158) );
  INVX1_HVT U534 ( .A(n764), .Y(n1004) );
  INVX1_HVT U535 ( .A(n751), .Y(n759) );
  NAND2X0_HVT U536 ( .A1(n722), .A2(n319), .Y(n1299) );
  INVX1_HVT U537 ( .A(n747), .Y(n748) );
  INVX1_HVT U538 ( .A(n788), .Y(n745) );
  NAND2X0_HVT U539 ( .A1(n219), .A2(n1326), .Y(n788) );
  INVX1_HVT U540 ( .A(n666), .Y(n667) );
  INVX1_HVT U541 ( .A(n1148), .Y(n1125) );
  INVX1_HVT U542 ( .A(n609), .Y(n607) );
  INVX1_HVT U543 ( .A(n598), .Y(n829) );
  INVX1_HVT U544 ( .A(n778), .Y(n691) );
  INVX1_HVT U545 ( .A(n678), .Y(n707) );
  INVX1_HVT U546 ( .A(n1644), .Y(n1645) );
  INVX1_HVT U547 ( .A(n588), .Y(n589) );
  INVX1_HVT U548 ( .A(n610), .Y(n626) );
  NAND3X0_HVT U549 ( .A1(n241), .A2(n262), .A3(n235), .Y(n1198) );
  NAND2X0_HVT U550 ( .A1(n1174), .A2(n1326), .Y(n1148) );
  INVX1_HVT U551 ( .A(n1429), .Y(n1424) );
  INVX1_HVT U552 ( .A(n1433), .Y(n1428) );
  INVX1_HVT U553 ( .A(n1409), .Y(n1406) );
  INVX1_HVT U554 ( .A(n1411), .Y(n1417) );
  INVX1_HVT U555 ( .A(n1435), .Y(n1438) );
  INVX1_HVT U556 ( .A(n1708), .Y(n1709) );
  INVX1_HVT U557 ( .A(n1701), .Y(n1702) );
  INVX1_HVT U558 ( .A(n1694), .Y(n1695) );
  NAND2X0_HVT U559 ( .A1(n172), .A2(n1941), .Y(n1721) );
  INVX1_HVT U560 ( .A(n1606), .Y(n1605) );
  INVX1_HVT U561 ( .A(n1587), .Y(n1586) );
  INVX1_HVT U562 ( .A(n1592), .Y(n1593) );
  INVX1_HVT U563 ( .A(n1588), .Y(n1589) );
  NAND2X0_HVT U564 ( .A1(n172), .A2(n1849), .Y(n1614) );
  NAND2X0_HVT U565 ( .A1(n183), .A2(n1560), .Y(net31204) );
  NOR4X1_HVT U566 ( .A1(n1548), .A2(n314), .A3(channel_cnt[3]), .A4(
        channel_cnt[2]), .Y(n555) );
  AND4X1_HVT U567 ( .A1(n1356), .A2(n1446), .A3(n1361), .A4(n1365), .Y(n280)
         );
  OAI222X1_HVT U568 ( .A1(sram_raddr_weight[5]), .A2(n1438), .A3(
        sram_raddr_weight[5]), .A4(n1455), .A5(n437), .A6(n1437), .Y(n290) );
  OAI221X1_HVT U569 ( .A1(sram_raddr_b4[5]), .A2(n1202), .A3(n271), .A4(n932), 
        .A5(n225), .Y(n291) );
  OAI221X1_HVT U570 ( .A1(n1133), .A2(n1132), .A3(n1133), .A4(n1131), .A5(n205), .Y(n292) );
  OAI221X1_HVT U571 ( .A1(n1144), .A2(n1162), .A3(n1144), .A4(n1143), .A5(n206), .Y(n293) );
  OAI221X1_HVT U572 ( .A1(n1122), .A2(n1162), .A3(n1122), .A4(n1121), .A5(n203), .Y(n294) );
  OAI221X1_HVT U573 ( .A1(n734), .A2(n1320), .A3(n734), .A4(n996), .A5(n204), 
        .Y(n295) );
  AOI22X1_HVT U574 ( .A1(n178), .A2(n1083), .A3(n1082), .A4(n1162), .Y(n296)
         );
  AOI22X1_HVT U575 ( .A1(n1777), .A2(n1803), .A3(sram_raddr_a4[2]), .A4(n1934), 
        .Y(n297) );
  AOI22X1_HVT U576 ( .A1(sram_raddr_b7[1]), .A2(n1236), .A3(n1178), .A4(n1248), 
        .Y(n298) );
  AOI22X1_HVT U577 ( .A1(n1974), .A2(n237), .A3(n1897), .A4(n1931), .Y(n299)
         );
  AOI22X1_HVT U578 ( .A1(sram_raddr_a6[2]), .A2(n1887), .A3(n1851), .A4(n1885), 
        .Y(n300) );
  AOI22X1_HVT U579 ( .A1(sram_raddr_b8[1]), .A2(n1332), .A3(n1264), .A4(n1336), 
        .Y(n301) );
  AOI22X1_HVT U580 ( .A1(sram_raddr_a0[9]), .A2(n1626), .A3(n1625), .A4(n1624), 
        .Y(n315) );
  AND3X1_HVT U581 ( .A1(n1280), .A2(n995), .A3(n994), .Y(n352) );
  OAI221X1_HVT U582 ( .A1(sram_raddr_a1[2]), .A2(n1637), .A3(sram_raddr_a1[2]), 
        .A4(n1664), .A5(n1630), .Y(n374) );
  OAI221X1_HVT U583 ( .A1(n931), .A2(n961), .A3(n931), .A4(n930), .A5(n1557), 
        .Y(n375) );
  AOI22X1_HVT U584 ( .A1(n1738), .A2(n1769), .A3(sram_raddr_a3[2]), .A4(n1887), 
        .Y(n376) );
  AOI22X1_HVT U585 ( .A1(sram_raddr_a2[9]), .A2(n1733), .A3(n1732), .A4(n1731), 
        .Y(n377) );
  AOI22X1_HVT U586 ( .A1(sram_raddr_a1[9]), .A2(n1678), .A3(n1677), .A4(n1676), 
        .Y(n378) );
  AOI22X1_HVT U587 ( .A1(sram_raddr_a6[1]), .A2(n1887), .A3(n1868), .A4(n1850), 
        .Y(n379) );
  AOI22X1_HVT U588 ( .A1(sram_raddr_a6[9]), .A2(n1887), .A3(n1886), .A4(n1885), 
        .Y(n380) );
  NAND2X0_HVT U589 ( .A1(n167), .A2(n1897), .Y(n381) );
  NAND2X0_HVT U590 ( .A1(n1896), .A2(n248), .Y(n382) );
  NAND2X0_HVT U591 ( .A1(n172), .A2(n1913), .Y(n1664) );
  NAND2X0_HVT U592 ( .A1(n515), .A2(n516), .Y(n383) );
  NAND2X0_HVT U593 ( .A1(n507), .A2(n508), .Y(n384) );
  NAND2X0_HVT U594 ( .A1(n503), .A2(n504), .Y(n385) );
  NAND2X0_HVT U595 ( .A1(n505), .A2(n506), .Y(n386) );
  NAND2X0_HVT U596 ( .A1(n501), .A2(n502), .Y(n387) );
  AND3X1_HVT U597 ( .A1(n1416), .A2(n1466), .A3(n1562), .Y(n399) );
  AND2X1_HVT U598 ( .A1(n1355), .A2(n1563), .Y(n421) );
  NAND2X0_HVT U599 ( .A1(sram_raddr_a7[9]), .A2(n1934), .Y(n471) );
  NAND3X0_HVT U600 ( .A1(n1933), .A2(n470), .A3(n471), .Y(n_sram_raddr_a7[9])
         );
  NAND2X0_HVT U601 ( .A1(sram_raddr_a7[2]), .A2(n1934), .Y(n472) );
  NAND3X0_HVT U602 ( .A1(n299), .A2(n477), .A3(n472), .Y(n_sram_raddr_a7[2])
         );
  NAND2X0_HVT U603 ( .A1(n1974), .A2(n1888), .Y(n474) );
  NAND3X0_HVT U604 ( .A1(n380), .A2(n473), .A3(n474), .Y(n_sram_raddr_a6[9])
         );
  NAND2X0_HVT U605 ( .A1(n1974), .A2(n236), .Y(n475) );
  NAND3X0_HVT U606 ( .A1(n300), .A2(n382), .A3(n475), .Y(n_sram_raddr_a6[2])
         );
  NAND2X0_HVT U607 ( .A1(n170), .A2(sram_raddr_a3[1]), .Y(n476) );
  NAND3X0_HVT U608 ( .A1(n379), .A2(n1848), .A3(n476), .Y(n_sram_raddr_a6[1])
         );
  NAND2X0_HVT U609 ( .A1(n1896), .A2(n247), .Y(n477) );
  NAND3X0_HVT U610 ( .A1(n297), .A2(n381), .A3(n477), .Y(n_sram_raddr_a4[2])
         );
  NAND2X0_HVT U611 ( .A1(n1851), .A2(n167), .Y(n478) );
  NAND3X0_HVT U612 ( .A1(n376), .A2(n382), .A3(n478), .Y(n_sram_raddr_a3[2])
         );
  NAND2X0_HVT U613 ( .A1(n170), .A2(n1844), .Y(n480) );
  NAND3X0_HVT U614 ( .A1(n377), .A2(n479), .A3(n480), .Y(n_sram_raddr_a2[9])
         );
  NAND2X0_HVT U615 ( .A1(n170), .A2(n1804), .Y(n482) );
  NAND3X0_HVT U616 ( .A1(n378), .A2(n481), .A3(n482), .Y(n_sram_raddr_a1[9])
         );
  NAND2X0_HVT U617 ( .A1(n1974), .A2(n1777), .Y(n483) );
  NAND3X0_HVT U618 ( .A1(n381), .A2(n374), .A3(n483), .Y(n_sram_raddr_a1[2])
         );
  NAND2X0_HVT U619 ( .A1(n170), .A2(n1770), .Y(n485) );
  NAND3X0_HVT U620 ( .A1(n315), .A2(n484), .A3(n485), .Y(n_sram_raddr_a0[9])
         );
  NAND2X0_HVT U621 ( .A1(n206), .A2(n1439), .Y(n486) );
  NAND3X0_HVT U622 ( .A1(n290), .A2(n399), .A3(n486), .Y(net22797) );
  NAND2X0_HVT U623 ( .A1(n1558), .A2(n462), .Y(n487) );
  NAND3X0_HVT U624 ( .A1(n280), .A2(n421), .A3(n487), .Y(n_state[0]) );
  NAND2X0_HVT U625 ( .A1(n178), .A2(n1265), .Y(n488) );
  NAND3X0_HVT U626 ( .A1(n301), .A2(n1263), .A3(n488), .Y(n1267) );
  NAND2X0_HVT U627 ( .A1(n1218), .A2(n1248), .Y(n489) );
  NAND3X0_HVT U628 ( .A1(n1217), .A2(n387), .A3(n489), .Y(n1223) );
  NAND2X0_HVT U629 ( .A1(n178), .A2(n1179), .Y(n490) );
  NAND3X0_HVT U630 ( .A1(n298), .A2(n1177), .A3(n490), .Y(n1180) );
  NAND2X0_HVT U631 ( .A1(sram_raddr_b6[7]), .A2(n232), .Y(n491) );
  NAND3X0_HVT U632 ( .A1(n385), .A2(n293), .A3(n491), .Y(n_sram_raddr_b6[7])
         );
  NAND2X0_HVT U633 ( .A1(sram_raddr_b6[6]), .A2(n233), .Y(n492) );
  NAND3X0_HVT U634 ( .A1(n386), .A2(n292), .A3(n492), .Y(n_sram_raddr_b6[6])
         );
  NAND2X0_HVT U635 ( .A1(sram_raddr_b6[5]), .A2(n233), .Y(n493) );
  NAND3X0_HVT U636 ( .A1(n384), .A2(n294), .A3(n493), .Y(n_sram_raddr_b6[5])
         );
  NAND2X0_HVT U637 ( .A1(sram_raddr_b6[1]), .A2(n1084), .Y(n494) );
  NAND3X0_HVT U638 ( .A1(n296), .A2(n1081), .A3(n494), .Y(n1085) );
  NAND2X0_HVT U639 ( .A1(n996), .A2(n1018), .Y(n496) );
  NAND3X0_HVT U640 ( .A1(n352), .A2(n495), .A3(n496), .Y(n1001) );
  NAND2X0_HVT U641 ( .A1(sram_raddr_b4[5]), .A2(n234), .Y(n497) );
  NAND3X0_HVT U642 ( .A1(n291), .A2(n375), .A3(n497), .Y(n_sram_raddr_b4[5])
         );
  NAND2X0_HVT U643 ( .A1(sram_raddr_b2[3]), .A2(n233), .Y(n498) );
  NAND3X0_HVT U644 ( .A1(n383), .A2(n295), .A3(n498), .Y(n_sram_raddr_b2[3])
         );
  AND2X1_HVT U645 ( .A1(n517), .A2(n518), .Y(n1838) );
  AND2X1_HVT U646 ( .A1(n1391), .A2(n1400), .Y(n499) );
  OR2X1_HVT U647 ( .A1(n403), .A2(n228), .Y(n500) );
  AND2X1_HVT U648 ( .A1(n499), .A2(n500), .Y(n1396) );
  AND2X1_HVT U649 ( .A1(n1227), .A2(n178), .Y(n501) );
  OR2X1_HVT U650 ( .A1(n1214), .A2(sram_raddr_b4[6]), .Y(n502) );
  AND2X1_HVT U651 ( .A1(n1146), .A2(n225), .Y(n503) );
  OR2X1_HVT U652 ( .A1(n1147), .A2(sram_raddr_b6[7]), .Y(n504) );
  AND2X1_HVT U653 ( .A1(n1145), .A2(n223), .Y(n505) );
  OR2X1_HVT U654 ( .A1(n1135), .A2(sram_raddr_b6[6]), .Y(n506) );
  AND2X1_HVT U655 ( .A1(n1134), .A2(n225), .Y(n507) );
  OR2X1_HVT U656 ( .A1(n1123), .A2(sram_raddr_b6[5]), .Y(n508) );
  AND2X1_HVT U657 ( .A1(n1069), .A2(n1072), .Y(n509) );
  OR2X1_HVT U658 ( .A1(n1070), .A2(n1071), .Y(n510) );
  AND2X1_HVT U659 ( .A1(n509), .A2(n510), .Y(n1074) );
  AND2X1_HVT U660 ( .A1(n972), .A2(n975), .Y(n511) );
  OR2X1_HVT U661 ( .A1(n973), .A2(n974), .Y(n512) );
  AND2X1_HVT U662 ( .A1(n511), .A2(n512), .Y(n976) );
  AND2X1_HVT U663 ( .A1(n744), .A2(n746), .Y(n513) );
  OR2X1_HVT U664 ( .A1(n264), .A2(n745), .Y(n514) );
  AND2X1_HVT U665 ( .A1(n513), .A2(n514), .Y(n749) );
  AND2X1_HVT U666 ( .A1(n1002), .A2(n188), .Y(n515) );
  OR2X1_HVT U667 ( .A1(sram_raddr_b2[2]), .A2(sram_raddr_b2[3]), .Y(n516) );
  AND2X1_HVT U668 ( .A1(n338), .A2(n1571), .Y(n517) );
  OR2X1_HVT U669 ( .A1(n1570), .A2(n259), .Y(n518) );
  AND2X1_HVT U670 ( .A1(n517), .A2(n518), .Y(n519) );
  AO21X1_HVT U671 ( .A1(n521), .A2(n522), .A3(n229), .Y(N2914) );
  AND2X1_HVT U672 ( .A1(col[1]), .A2(col[0]), .Y(n1565) );
  NAND3X0_HVT U673 ( .A1(n1565), .A2(col[3]), .A3(n235), .Y(n520) );
  AND3X1_HVT U674 ( .A1(n1993), .A2(n1051), .A3(n1052), .Y(
        n_addr_col_sel_cnt[0]) );
  AND3X1_HVT U675 ( .A1(n1051), .A2(n1993), .A3(addr_col_sel_cnt[0]), .Y(
        n_addr_col_sel_cnt[1]) );
  AO21X1_HVT U676 ( .A1(addr_row_sel_cnt[0]), .A2(n1993), .A3(n1567), .Y(
        n_addr_row_sel_cnt_0_) );
  AO22X1_HVT U677 ( .A1(col[1]), .A2(n1354), .A3(n1363), .A4(data_sel_col[1]), 
        .Y(n1996) );
  AO22X1_HVT U678 ( .A1(row[1]), .A2(n1354), .A3(n1363), .A4(data_sel_row[1]), 
        .Y(n2000) );
  AO22X1_HVT U679 ( .A1(row[0]), .A2(n1354), .A3(n1363), .A4(data_sel_row[0]), 
        .Y(n1999) );
  NAND2X0_HVT U680 ( .A1(n2003), .A2(n1999), .Y(n523) );
  OA22X1_HVT U681 ( .A1(n524), .A2(n1389), .A3(n1994), .A4(n523), .Y(n1662) );
  AO22X1_HVT U682 ( .A1(col[0]), .A2(n1354), .A3(n1363), .A4(data_sel_col[0]), 
        .Y(n1995) );
  AND2X1_HVT U683 ( .A1(n253), .A2(n240), .Y(n1445) );
  NAND3X0_HVT U684 ( .A1(n228), .A2(n554), .A3(n1389), .Y(n1997) );
  NAND2X0_HVT U685 ( .A1(n221), .A2(n554), .Y(n2001) );
  NAND3X0_HVT U686 ( .A1(n2003), .A2(n1996), .A3(n1995), .Y(n1655) );
  AND4X1_HVT U687 ( .A1(conv1_weight_cnt[2]), .A2(conv1_weight_cnt[4]), .A3(
        n526), .A4(n525), .Y(n_conv1_done) );
  NAND4X0_HVT U688 ( .A1(state[1]), .A2(n1023), .A3(n1024), .A4(n253), .Y(
        n1355) );
  AO22X1_HVT U689 ( .A1(row[1]), .A2(col[3]), .A3(row[0]), .A4(col[2]), .Y(
        n531) );
  OA21X1_HVT U690 ( .A1(row[0]), .A2(col[2]), .A3(n1565), .Y(n532) );
  NAND2X0_HVT U691 ( .A1(n349), .A2(n241), .Y(n548) );
  NAND2X0_HVT U692 ( .A1(row[1]), .A2(col[3]), .Y(n547) );
  NAND2X0_HVT U693 ( .A1(n548), .A2(n547), .Y(n550) );
  NAND3X0_HVT U694 ( .A1(row[1]), .A2(row[3]), .A3(n256), .Y(n1570) );
  NAND2X0_HVT U695 ( .A1(n256), .A2(n557), .Y(n537) );
  OR2X1_HVT U696 ( .A1(n1389), .A2(n533), .Y(n1369) );
  OR4X1_HVT U697 ( .A1(conv_done), .A2(conv2_weight_cnt[3]), .A3(
        conv2_weight_cnt[0]), .A4(conv2_weight_cnt[2]), .Y(n528) );
  NAND4X0_HVT U698 ( .A1(n1354), .A2(conv2_weight_cnt[5]), .A3(
        conv2_weight_cnt[1]), .A4(conv2_weight_cnt[4]), .Y(n527) );
  AND2X1_HVT U699 ( .A1(n2003), .A2(n254), .Y(n1558) );
  NAND2X0_HVT U700 ( .A1(n1226), .A2(n319), .Y(n1078) );
  NOR2X0_HVT U701 ( .A1(n554), .A2(channel_cnt[0]), .Y(net22938) );
  OR2X1_HVT U702 ( .A1(channel_cnt[2]), .A2(channel_cnt[3]), .Y(n529) );
  AO22X1_HVT U703 ( .A1(n1558), .A2(n1132), .A3(net22938), .A4(n530), .Y(
        n_load_data_enable) );
  NAND2X0_HVT U704 ( .A1(n256), .A2(n313), .Y(n546) );
  AO221X1_HVT U705 ( .A1(n548), .A2(n532), .A3(n548), .A4(n531), .A5(n546), 
        .Y(n1390) );
  NAND2X0_HVT U706 ( .A1(n207), .A2(n1441), .Y(n1457) );
  NAND2X0_HVT U707 ( .A1(n2003), .A2(n533), .Y(n1368) );
  OA22X1_HVT U708 ( .A1(n551), .A2(n1457), .A3(n1569), .A4(n1368), .Y(n1388)
         );
  NAND2X0_HVT U709 ( .A1(n1465), .A2(n1388), .Y(n536) );
  AO22X1_HVT U710 ( .A1(n1569), .A2(n534), .A3(n551), .A4(n1443), .Y(n538) );
  AO22X1_HVT U711 ( .A1(row[0]), .A2(n536), .A3(n259), .A4(n538), .Y(n_row[0])
         );
  AO21X1_HVT U712 ( .A1(row[0]), .A2(n538), .A3(row[1]), .Y(n535) );
  OA221X1_HVT U713 ( .A1(n536), .A2(n557), .A3(n536), .A4(n538), .A5(n535), 
        .Y(n_row[1]) );
  AO221X1_HVT U715 ( .A1(n538), .A2(n256), .A3(n538), .A4(n557), .A5(n536), 
        .Y(n539) );
  AND3X1_HVT U716 ( .A1(row[0]), .A2(row[1]), .A3(n538), .Y(n540) );
  AO22X1_HVT U717 ( .A1(row[2]), .A2(n540), .A3(row[3]), .A4(n539), .Y(
        n_row[3]) );
  AND2X1_HVT U718 ( .A1(n543), .A2(n542), .Y(n541) );
  AND2X1_HVT U719 ( .A1(n1469), .A2(n541), .Y(n_sram_bytemask_b[0]) );
  AND3X1_HVT U720 ( .A1(n545), .A2(n1469), .A3(n542), .Y(n_sram_bytemask_b[1])
         );
  AND3X1_HVT U721 ( .A1(n1469), .A2(n544), .A3(n543), .Y(n_sram_bytemask_b[2])
         );
  AND3X1_HVT U722 ( .A1(n1469), .A2(n545), .A3(n544), .Y(n_sram_bytemask_b[3])
         );
  AND3X1_HVT U723 ( .A1(n1354), .A2(n541), .A3(n1512), .Y(n_sram_bytemask_c[0]) );
  AND4X1_HVT U724 ( .A1(n1354), .A2(n545), .A3(n1512), .A4(n542), .Y(
        n_sram_bytemask_c[1]) );
  AND4X1_HVT U725 ( .A1(n1354), .A2(n544), .A3(n1512), .A4(n543), .Y(
        n_sram_bytemask_c[2]) );
  AND4X1_HVT U726 ( .A1(n1354), .A2(n545), .A3(n544), .A4(n1512), .Y(
        n_sram_bytemask_c[3]) );
  AND3X1_HVT U727 ( .A1(mem_sel), .A2(n1354), .A3(n541), .Y(
        n_sram_bytemask_d[0]) );
  AND4X1_HVT U728 ( .A1(n1354), .A2(mem_sel), .A3(n545), .A4(n542), .Y(
        n_sram_bytemask_d[1]) );
  AND4X1_HVT U729 ( .A1(n1354), .A2(mem_sel), .A3(n544), .A4(n543), .Y(
        n_sram_bytemask_d[2]) );
  AND4X1_HVT U730 ( .A1(mem_sel), .A2(n1354), .A3(n545), .A4(n544), .Y(
        n_sram_bytemask_d[3]) );
  NAND2X0_HVT U731 ( .A1(n241), .A2(n235), .Y(n576) );
  AO21X1_HVT U732 ( .A1(n1565), .A2(n546), .A3(n576), .Y(n1306) );
  AO22X1_HVT U733 ( .A1(col[1]), .A2(col[0]), .A3(n319), .A4(n262), .Y(n1387)
         );
  NAND2X0_HVT U734 ( .A1(n214), .A2(n1387), .Y(n1084) );
  NAND2X0_HVT U735 ( .A1(n219), .A2(n1078), .Y(n610) );
  NAND4X0_HVT U736 ( .A1(n549), .A2(n548), .A3(n259), .A4(n547), .Y(n1259) );
  AO22X1_HVT U737 ( .A1(n191), .A2(n418), .A3(n178), .A4(n285), .Y(n553) );
  AO221X1_HVT U738 ( .A1(sram_raddr_b0[0]), .A2(n1084), .A3(n250), .A4(n610), 
        .A5(n553), .Y(n558) );
  NAND2X0_HVT U739 ( .A1(n1549), .A2(n555), .Y(n1361) );
  AO22X1_HVT U740 ( .A1(n203), .A2(n558), .A3(sram_raddr_b0[0]), .A4(n168), 
        .Y(n_sram_raddr_b0[0]) );
  NAND2X0_HVT U741 ( .A1(sram_raddr_b3[0]), .A2(sram_raddr_b3[1]), .Y(n563) );
  NAND2X0_HVT U742 ( .A1(n285), .A2(n367), .Y(n1109) );
  NAND2X0_HVT U743 ( .A1(n563), .A2(n1109), .Y(n1083) );
  OA22X1_HVT U744 ( .A1(n1158), .A2(n364), .A3(n173), .A4(n1083), .Y(n560) );
  NAND2X0_HVT U745 ( .A1(sram_raddr_b6[1]), .A2(sram_raddr_b6[0]), .Y(n562) );
  OA21X1_HVT U746 ( .A1(sram_raddr_b6[1]), .A2(sram_raddr_b6[0]), .A3(n562), 
        .Y(n1082) );
  NAND2X0_HVT U747 ( .A1(n192), .A2(n1082), .Y(n807) );
  NAND2X0_HVT U748 ( .A1(sram_raddr_b0[0]), .A2(sram_raddr_b0[1]), .Y(n805) );
  NAND2X0_HVT U749 ( .A1(n250), .A2(n364), .Y(n830) );
  NAND3X0_HVT U750 ( .A1(n805), .A2(n610), .A3(n830), .Y(n559) );
  NAND3X0_HVT U751 ( .A1(n560), .A2(n807), .A3(n559), .Y(n561) );
  AO22X1_HVT U752 ( .A1(n204), .A2(n561), .A3(sram_raddr_b0[1]), .A4(n217), 
        .Y(n_sram_raddr_b0[1]) );
  NAND2X0_HVT U753 ( .A1(n242), .A2(n562), .Y(n569) );
  OA21X1_HVT U754 ( .A1(n562), .A2(n242), .A3(n569), .Y(n1089) );
  NAND2X0_HVT U755 ( .A1(n326), .A2(n563), .Y(n578) );
  OA21X1_HVT U756 ( .A1(n563), .A2(n326), .A3(n578), .Y(n810) );
  OA22X1_HVT U757 ( .A1(n1089), .A2(n1259), .A3(n810), .A4(n226), .Y(n813) );
  OA21X1_HVT U758 ( .A1(n626), .A2(n805), .A3(n215), .Y(n564) );
  NAND4X0_HVT U759 ( .A1(col[0]), .A2(n241), .A3(n319), .A4(n235), .Y(n1174)
         );
  NAND2X0_HVT U760 ( .A1(n219), .A2(n1174), .Y(n678) );
  NAND2X0_HVT U761 ( .A1(n707), .A2(n1198), .Y(n778) );
  NAND3X0_HVT U762 ( .A1(n564), .A2(n279), .A3(n778), .Y(n568) );
  NAND2X0_HVT U763 ( .A1(n813), .A2(n568), .Y(n566) );
  OA221X1_HVT U764 ( .A1(n566), .A2(sram_raddr_b0[2]), .A3(n566), .A4(n565), 
        .A5(n207), .Y(n567) );
  AO221X1_HVT U765 ( .A1(sram_raddr_b0[2]), .A2(n233), .A3(n279), .A4(n224), 
        .A5(n567), .Y(n_sram_raddr_b0[2]) );
  NAND2X0_HVT U766 ( .A1(sram_raddr_b0[3]), .A2(n234), .Y(n575) );
  AND2X1_HVT U767 ( .A1(n216), .A2(n568), .Y(n570) );
  NAND2X0_HVT U768 ( .A1(n411), .A2(n570), .Y(n571) );
  NAND2X0_HVT U769 ( .A1(sram_raddr_b6[3]), .A2(n569), .Y(n591) );
  OA21X1_HVT U770 ( .A1(sram_raddr_b6[3]), .A2(n569), .A3(n591), .Y(n1095) );
  NAND2X0_HVT U771 ( .A1(n192), .A2(n1095), .Y(n821) );
  OA221X1_HVT U772 ( .A1(n691), .A2(n571), .A3(n570), .A4(n411), .A5(n821), 
        .Y(n572) );
  HADDX1_HVT U773 ( .A0(n393), .B0(n578), .SO(n818) );
  AO221X1_HVT U774 ( .A1(n572), .A2(n227), .A3(n572), .A4(n818), .A5(n228), 
        .Y(n574) );
  AO221X1_HVT U775 ( .A1(sram_raddr_b0[3]), .A2(sram_raddr_b0[2]), .A3(n411), 
        .A4(n279), .A5(n1366), .Y(n573) );
  NAND3X0_HVT U776 ( .A1(n575), .A2(n574), .A3(n573), .Y(n_sram_raddr_b0[3])
         );
  NAND2X0_HVT U777 ( .A1(sram_raddr_b0[3]), .A2(sram_raddr_b0[2]), .Y(n827) );
  NAND3X0_HVT U778 ( .A1(sram_raddr_b0[3]), .A2(sram_raddr_b0[0]), .A3(
        sram_raddr_b0[1]), .Y(n606) );
  AND3X1_HVT U779 ( .A1(n827), .A2(n323), .A3(n606), .Y(n577) );
  NAND3X0_HVT U780 ( .A1(col[1]), .A2(n722), .A3(n262), .Y(n1326) );
  NAND2X0_HVT U781 ( .A1(n827), .A2(n323), .Y(n586) );
  NAND3X0_HVT U782 ( .A1(sram_raddr_b0[3]), .A2(sram_raddr_b0[2]), .A3(
        sram_raddr_b0[4]), .Y(n598) );
  NAND2X0_HVT U783 ( .A1(n586), .A2(n598), .Y(n583) );
  AO22X1_HVT U784 ( .A1(n577), .A2(n610), .A3(n1148), .A4(n583), .Y(n590) );
  OA221X1_HVT U785 ( .A1(n626), .A2(n827), .A3(n626), .A4(n606), .A5(n213), 
        .Y(n587) );
  NAND2X0_HVT U786 ( .A1(sram_raddr_b3[3]), .A2(n578), .Y(n579) );
  NAND2X0_HVT U787 ( .A1(n579), .A2(n320), .Y(n588) );
  OA21X1_HVT U788 ( .A1(n320), .A2(n579), .A3(n588), .Y(n831) );
  OA22X1_HVT U789 ( .A1(n587), .A2(n323), .A3(n831), .A4(n226), .Y(n581) );
  AO22X1_HVT U790 ( .A1(n580), .A2(sram_raddr_b6[4]), .A3(n591), .A4(n276), 
        .Y(n1105) );
  NAND2X0_HVT U791 ( .A1(n190), .A2(n1105), .Y(n833) );
  NAND3X0_HVT U792 ( .A1(n582), .A2(n581), .A3(n833), .Y(n585) );
  AO222X1_HVT U793 ( .A1(n585), .A2(n203), .A3(n233), .A4(sram_raddr_b0[4]), 
        .A5(n223), .A6(n584), .Y(n_sram_raddr_b0[4]) );
  NAND2X0_HVT U794 ( .A1(n589), .A2(n261), .Y(n592) );
  OA21X1_HVT U795 ( .A1(n589), .A2(n261), .A3(n592), .Y(n838) );
  NAND3X0_HVT U796 ( .A1(n272), .A2(n598), .A3(n590), .Y(n594) );
  NAND3X0_HVT U797 ( .A1(n591), .A2(n339), .A3(n276), .Y(n593) );
  NAND2X0_HVT U798 ( .A1(n191), .A2(n1121), .Y(n841) );
  NAND4X0_HVT U799 ( .A1(sram_raddr_b0[3]), .A2(sram_raddr_b0[2]), .A3(
        sram_raddr_b0[5]), .A4(sram_raddr_b0[4]), .Y(n597) );
  NAND2X0_HVT U800 ( .A1(sram_raddr_b3[6]), .A2(n592), .Y(n603) );
  OA21X1_HVT U801 ( .A1(sram_raddr_b3[6]), .A2(n592), .A3(n603), .Y(n851) );
  NAND2X0_HVT U802 ( .A1(n851), .A2(n178), .Y(n596) );
  NAND2X0_HVT U803 ( .A1(sram_raddr_b6[6]), .A2(n593), .Y(n604) );
  OA21X1_HVT U804 ( .A1(sram_raddr_b6[6]), .A2(n593), .A3(n604), .Y(n1131) );
  NAND2X0_HVT U805 ( .A1(n190), .A2(n1131), .Y(n848) );
  NAND3X0_HVT U806 ( .A1(n827), .A2(n272), .A3(n323), .Y(n609) );
  AO222X1_HVT U807 ( .A1(n626), .A2(n607), .A3(n626), .A4(n1125), .A5(n607), 
        .A6(n606), .Y(n602) );
  OA222X1_HVT U808 ( .A1(n391), .A2(n215), .A3(n391), .A4(n594), .A5(
        sram_raddr_b0[6]), .A6(n602), .Y(n595) );
  NAND3X0_HVT U809 ( .A1(n596), .A2(n848), .A3(n595), .Y(n601) );
  AO221X1_HVT U810 ( .A1(n188), .A2(n391), .A3(n188), .A4(n597), .A5(n233), 
        .Y(n617) );
  NAND3X0_HVT U811 ( .A1(n225), .A2(sram_raddr_b0[5]), .A3(n829), .Y(n599) );
  NAND2X0_HVT U812 ( .A1(n391), .A2(n599), .Y(n600) );
  AO22X1_HVT U813 ( .A1(n1557), .A2(n601), .A3(n617), .A4(n600), .Y(
        n_sram_raddr_b0[6]) );
  AND4X1_HVT U814 ( .A1(n188), .A2(sram_raddr_b0[6]), .A3(sram_raddr_b0[5]), 
        .A4(n829), .Y(n634) );
  OA21X1_HVT U815 ( .A1(n602), .A2(n391), .A3(n214), .Y(n613) );
  NAND2X0_HVT U816 ( .A1(n350), .A2(n603), .Y(n631) );
  OA21X1_HVT U817 ( .A1(n603), .A2(n350), .A3(n631), .Y(n862) );
  OA22X1_HVT U818 ( .A1(n613), .A2(n263), .A3(n862), .A4(n173), .Y(n605) );
  NAND2X0_HVT U819 ( .A1(n270), .A2(n604), .Y(n627) );
  NAND2X0_HVT U820 ( .A1(n192), .A2(n1143), .Y(n860) );
  NAND2X0_HVT U821 ( .A1(n605), .A2(n860), .Y(n611) );
  NAND2X0_HVT U822 ( .A1(n607), .A2(n606), .Y(n608) );
  NAND2X0_HVT U823 ( .A1(sram_raddr_b0[6]), .A2(n608), .Y(n624) );
  NAND2X0_HVT U824 ( .A1(sram_raddr_b0[6]), .A2(n609), .Y(n622) );
  AO22X1_HVT U825 ( .A1(n610), .A2(n624), .A3(n1148), .A4(n622), .Y(n614) );
  OA221X1_HVT U826 ( .A1(n611), .A2(n263), .A3(n611), .A4(n614), .A5(n204), 
        .Y(n612) );
  AO221X1_HVT U827 ( .A1(sram_raddr_b0[7]), .A2(n617), .A3(n263), .A4(n634), 
        .A5(n612), .Y(n_sram_raddr_b0[7]) );
  HADDX1_HVT U828 ( .A0(sram_raddr_b3[8]), .B0(n631), .SO(n870) );
  OA22X1_HVT U829 ( .A1(n613), .A2(n329), .A3(n870), .A4(n227), .Y(n616) );
  HADDX1_HVT U830 ( .A0(n388), .B0(n627), .SO(n1155) );
  NAND2X0_HVT U831 ( .A1(n190), .A2(n1155), .Y(n873) );
  NAND3X0_HVT U832 ( .A1(n329), .A2(n263), .A3(n614), .Y(n630) );
  NAND3X0_HVT U833 ( .A1(sram_raddr_b0[8]), .A2(sram_raddr_b0[7]), .A3(n778), 
        .Y(n615) );
  NAND4X0_HVT U834 ( .A1(n616), .A2(n873), .A3(n630), .A4(n615), .Y(n620) );
  AO21X1_HVT U835 ( .A1(sram_raddr_b0[7]), .A2(n634), .A3(sram_raddr_b0[8]), 
        .Y(n619) );
  NAND2X0_HVT U836 ( .A1(sram_raddr_b0[8]), .A2(sram_raddr_b0[7]), .Y(n618) );
  AO21X1_HVT U837 ( .A1(n618), .A2(n168), .A3(n617), .Y(n621) );
  AO22X1_HVT U838 ( .A1(n205), .A2(n620), .A3(n619), .A4(n621), .Y(
        n_sram_raddr_b0[8]) );
  NAND2X0_HVT U839 ( .A1(sram_raddr_b0[9]), .A2(n621), .Y(n637) );
  AND2X1_HVT U840 ( .A1(n329), .A2(n263), .Y(n625) );
  OA221X1_HVT U841 ( .A1(n1125), .A2(n625), .A3(n1125), .A4(n622), .A5(n216), 
        .Y(n623) );
  OA221X1_HVT U842 ( .A1(n626), .A2(n625), .A3(n626), .A4(n624), .A5(n623), 
        .Y(n629) );
  OR2X1_HVT U843 ( .A1(n627), .A2(sram_raddr_b6[8]), .Y(n628) );
  HADDX1_HVT U844 ( .A0(n628), .B0(n406), .SO(n1163) );
  NAND2X0_HVT U845 ( .A1(n190), .A2(n1163), .Y(n884) );
  OA221X1_HVT U846 ( .A1(sram_raddr_b0[9]), .A2(n630), .A3(n423), .A4(n629), 
        .A5(n884), .Y(n633) );
  OR2X1_HVT U847 ( .A1(n631), .A2(sram_raddr_b3[8]), .Y(n632) );
  HADDX1_HVT U848 ( .A0(sram_raddr_b3[9]), .B0(n632), .SO(n885) );
  AO221X1_HVT U849 ( .A1(n633), .A2(n226), .A3(n633), .A4(n885), .A5(n228), 
        .Y(n636) );
  NAND4X0_HVT U850 ( .A1(sram_raddr_b0[7]), .A2(sram_raddr_b0[8]), .A3(n634), 
        .A4(n423), .Y(n635) );
  NAND3X0_HVT U851 ( .A1(n637), .A2(n636), .A3(n635), .Y(n_sram_raddr_b0[9])
         );
  NAND2X0_HVT U852 ( .A1(col[0]), .A2(n214), .Y(n1236) );
  AO22X1_HVT U853 ( .A1(n192), .A2(n419), .A3(n178), .A4(n286), .Y(n638) );
  AO221X1_HVT U854 ( .A1(sram_raddr_b1[0]), .A2(n1236), .A3(n251), .A4(n678), 
        .A5(n638), .Y(n639) );
  AO22X1_HVT U855 ( .A1(n205), .A2(n639), .A3(sram_raddr_b1[0]), .A4(n168), 
        .Y(n_sram_raddr_b1[0]) );
  NAND2X0_HVT U856 ( .A1(sram_raddr_b4[0]), .A2(sram_raddr_b4[1]), .Y(n643) );
  NAND2X0_HVT U857 ( .A1(n286), .A2(n372), .Y(n1203) );
  NAND2X0_HVT U858 ( .A1(n643), .A2(n1203), .Y(n1179) );
  OA22X1_HVT U859 ( .A1(n891), .A2(n365), .A3(n226), .A4(n1179), .Y(n641) );
  NAND2X0_HVT U860 ( .A1(sram_raddr_b7[1]), .A2(sram_raddr_b7[0]), .Y(n647) );
  OA21X1_HVT U861 ( .A1(sram_raddr_b7[1]), .A2(sram_raddr_b7[0]), .A3(n647), 
        .Y(n1178) );
  NAND2X0_HVT U862 ( .A1(n192), .A2(n1178), .Y(n894) );
  NAND2X0_HVT U863 ( .A1(sram_raddr_b1[0]), .A2(sram_raddr_b1[1]), .Y(n892) );
  NAND2X0_HVT U864 ( .A1(n251), .A2(n365), .Y(n897) );
  NAND3X0_HVT U865 ( .A1(n678), .A2(n892), .A3(n897), .Y(n640) );
  NAND3X0_HVT U866 ( .A1(n641), .A2(n894), .A3(n640), .Y(n642) );
  AO22X1_HVT U867 ( .A1(n1557), .A2(n642), .A3(sram_raddr_b1[1]), .A4(n217), 
        .Y(n_sram_raddr_b1[1]) );
  OA21X1_HVT U868 ( .A1(n707), .A2(n892), .A3(n216), .Y(n644) );
  NAND2X0_HVT U869 ( .A1(n322), .A2(n643), .Y(n656) );
  OA21X1_HVT U870 ( .A1(n643), .A2(n322), .A3(n656), .Y(n899) );
  NAND3X0_HVT U871 ( .A1(n644), .A2(n778), .A3(n273), .Y(n646) );
  AO22X1_HVT U872 ( .A1(sram_raddr_b7[2]), .A2(n645), .A3(n243), .A4(n647), 
        .Y(n1184) );
  NAND2X0_HVT U873 ( .A1(n191), .A2(n1184), .Y(n898) );
  NAND2X0_HVT U874 ( .A1(sram_raddr_b1[3]), .A2(n233), .Y(n654) );
  AO221X1_HVT U875 ( .A1(sram_raddr_b1[3]), .A2(sram_raddr_b1[2]), .A3(n414), 
        .A4(n273), .A5(n1366), .Y(n653) );
  AND2X1_HVT U876 ( .A1(n215), .A2(n646), .Y(n649) );
  NAND2X0_HVT U877 ( .A1(n414), .A2(n649), .Y(n650) );
  NAND2X0_HVT U878 ( .A1(n243), .A2(n647), .Y(n648) );
  NAND2X0_HVT U879 ( .A1(sram_raddr_b7[3]), .A2(n648), .Y(n669) );
  OA21X1_HVT U880 ( .A1(sram_raddr_b7[3]), .A2(n648), .A3(n669), .Y(n1189) );
  NAND2X0_HVT U881 ( .A1(n190), .A2(n1189), .Y(n909) );
  OA221X1_HVT U882 ( .A1(n691), .A2(n650), .A3(n649), .A4(n414), .A5(n909), 
        .Y(n651) );
  HADDX1_HVT U883 ( .A0(n389), .B0(n656), .SO(n906) );
  AO221X1_HVT U884 ( .A1(n651), .A2(n173), .A3(n651), .A4(n906), .A5(n228), 
        .Y(n652) );
  NAND3X0_HVT U885 ( .A1(n654), .A2(n653), .A3(n652), .Y(n_sram_raddr_b1[3])
         );
  NAND3X0_HVT U886 ( .A1(sram_raddr_b1[3]), .A2(sram_raddr_b1[2]), .A3(
        sram_raddr_b1[4]), .Y(n917) );
  NAND2X0_HVT U887 ( .A1(sram_raddr_b1[3]), .A2(sram_raddr_b1[2]), .Y(n916) );
  NAND2X0_HVT U888 ( .A1(n916), .A2(n335), .Y(n664) );
  NAND2X0_HVT U889 ( .A1(n917), .A2(n664), .Y(n661) );
  NAND3X0_HVT U890 ( .A1(sram_raddr_b1[3]), .A2(sram_raddr_b1[0]), .A3(
        sram_raddr_b1[1]), .Y(n675) );
  AND3X1_HVT U891 ( .A1(n916), .A2(n335), .A3(n675), .Y(n655) );
  AO22X1_HVT U892 ( .A1(n1226), .A2(n661), .A3(n655), .A4(n678), .Y(n668) );
  OA221X1_HVT U893 ( .A1(n707), .A2(n916), .A3(n707), .A4(n675), .A5(n213), 
        .Y(n665) );
  NAND2X0_HVT U894 ( .A1(sram_raddr_b4[3]), .A2(n656), .Y(n657) );
  NAND2X0_HVT U895 ( .A1(n657), .A2(n336), .Y(n666) );
  OA21X1_HVT U896 ( .A1(n336), .A2(n657), .A3(n666), .Y(n915) );
  OA22X1_HVT U897 ( .A1(n665), .A2(n335), .A3(n915), .A4(n227), .Y(n659) );
  AO22X1_HVT U898 ( .A1(n658), .A2(sram_raddr_b7[4]), .A3(n669), .A4(n277), 
        .Y(n1199) );
  NAND2X0_HVT U899 ( .A1(n192), .A2(n1199), .Y(n920) );
  NAND3X0_HVT U900 ( .A1(n660), .A2(n659), .A3(n920), .Y(n663) );
  AO222X1_HVT U901 ( .A1(n663), .A2(n204), .A3(n234), .A4(sram_raddr_b1[4]), 
        .A5(n224), .A6(n662), .Y(n_sram_raddr_b1[4]) );
  NAND2X0_HVT U902 ( .A1(n667), .A2(n271), .Y(n671) );
  OA21X1_HVT U903 ( .A1(n667), .A2(n271), .A3(n671), .Y(n929) );
  NAND3X0_HVT U904 ( .A1(n265), .A2(n917), .A3(n668), .Y(n670) );
  NAND3X0_HVT U905 ( .A1(n669), .A2(n340), .A3(n277), .Y(n672) );
  NAND2X0_HVT U906 ( .A1(n190), .A2(n1212), .Y(n928) );
  NAND4X0_HVT U907 ( .A1(sram_raddr_b1[3]), .A2(sram_raddr_b1[2]), .A3(
        sram_raddr_b1[5]), .A4(sram_raddr_b1[4]), .Y(n673) );
  NAND3X0_HVT U908 ( .A1(n916), .A2(n265), .A3(n335), .Y(n674) );
  NAND2X0_HVT U909 ( .A1(sram_raddr_b4[6]), .A2(n671), .Y(n680) );
  NAND2X0_HVT U910 ( .A1(sram_raddr_b7[6]), .A2(n672), .Y(n681) );
  OA21X1_HVT U911 ( .A1(sram_raddr_b7[6]), .A2(n672), .A3(n681), .Y(n1218) );
  NAND2X0_HVT U912 ( .A1(n190), .A2(n1218), .Y(n938) );
  OR3X1_HVT U914 ( .A1(n327), .A2(n265), .A3(n917), .Y(n684) );
  NAND2X0_HVT U915 ( .A1(sram_raddr_b1[6]), .A2(n674), .Y(n703) );
  NAND2X0_HVT U916 ( .A1(n676), .A2(n675), .Y(n677) );
  NAND2X0_HVT U917 ( .A1(sram_raddr_b1[6]), .A2(n677), .Y(n705) );
  AO22X1_HVT U918 ( .A1(n1226), .A2(n703), .A3(n678), .A4(n705), .Y(n689) );
  NAND2X0_HVT U919 ( .A1(n689), .A2(n317), .Y(n683) );
  AND2X1_HVT U920 ( .A1(n1226), .A2(n703), .Y(n679) );
  OA22X1_HVT U921 ( .A1(n891), .A2(n679), .A3(n707), .A4(n705), .Y(n692) );
  NAND2X0_HVT U922 ( .A1(n316), .A2(n680), .Y(n693) );
  OA21X1_HVT U923 ( .A1(n680), .A2(n316), .A3(n693), .Y(n943) );
  OA22X1_HVT U924 ( .A1(n692), .A2(n317), .A3(n943), .A4(n173), .Y(n682) );
  NAND2X0_HVT U925 ( .A1(n330), .A2(n681), .Y(n690) );
  NAND2X0_HVT U926 ( .A1(n192), .A2(n1229), .Y(n946) );
  NAND3X0_HVT U927 ( .A1(n683), .A2(n682), .A3(n946), .Y(n688) );
  NAND2X0_HVT U928 ( .A1(n317), .A2(n684), .Y(n687) );
  NAND2X0_HVT U929 ( .A1(sram_raddr_b1[7]), .A2(n697), .Y(n685) );
  NAND2X0_HVT U930 ( .A1(n223), .A2(n685), .Y(n696) );
  AO222X1_HVT U931 ( .A1(n688), .A2(n203), .A3(n687), .A4(n686), .A5(
        sram_raddr_b1[7]), .A6(n233), .Y(n_sram_raddr_b1[7]) );
  NAND3X0_HVT U932 ( .A1(n317), .A2(n267), .A3(n689), .Y(n711) );
  AO22X1_HVT U933 ( .A1(sram_raddr_b7[8]), .A2(n690), .A3(n353), .A4(n708), 
        .Y(n1240) );
  NAND2X0_HVT U934 ( .A1(n190), .A2(n1240), .Y(n959) );
  AO221X1_HVT U935 ( .A1(n692), .A2(n691), .A3(n692), .A4(n317), .A5(n267), 
        .Y(n695) );
  AO22X1_HVT U936 ( .A1(sram_raddr_b4[8]), .A2(n693), .A3(n328), .A4(n712), 
        .Y(n960) );
  NAND2X0_HVT U937 ( .A1(n178), .A2(n960), .Y(n694) );
  NAND4X0_HVT U938 ( .A1(n711), .A2(n959), .A3(n695), .A4(n694), .Y(n700) );
  NAND3X0_HVT U939 ( .A1(n225), .A2(sram_raddr_b1[7]), .A3(n697), .Y(n702) );
  NAND2X0_HVT U940 ( .A1(n267), .A2(n702), .Y(n698) );
  AO22X1_HVT U941 ( .A1(n207), .A2(n700), .A3(n699), .A4(n698), .Y(
        n_sram_raddr_b1[8]) );
  AO222X1_HVT U942 ( .A1(n409), .A2(n267), .A3(n409), .A4(n702), .A5(
        sram_raddr_b1[9]), .A6(n701), .Y(n716) );
  AND2X1_HVT U943 ( .A1(n317), .A2(n267), .Y(n706) );
  OA221X1_HVT U944 ( .A1(col[0]), .A2(n706), .A3(col[0]), .A4(n703), .A5(n214), 
        .Y(n704) );
  OA221X1_HVT U945 ( .A1(n707), .A2(n706), .A3(n707), .A4(n705), .A5(n704), 
        .Y(n710) );
  NAND2X0_HVT U946 ( .A1(n708), .A2(n353), .Y(n709) );
  HADDX1_HVT U947 ( .A0(n405), .B0(n709), .SO(n1249) );
  NAND2X0_HVT U948 ( .A1(n192), .A2(n1249), .Y(n972) );
  OA221X1_HVT U949 ( .A1(sram_raddr_b1[9]), .A2(n711), .A3(n409), .A4(n710), 
        .A5(n972), .Y(n714) );
  NAND2X0_HVT U950 ( .A1(n712), .A2(n328), .Y(n713) );
  HADDX1_HVT U951 ( .A0(sram_raddr_b4[9]), .B0(n713), .SO(n973) );
  AO221X1_HVT U952 ( .A1(n714), .A2(n226), .A3(n714), .A4(n973), .A5(n221), 
        .Y(n715) );
  NAND2X0_HVT U953 ( .A1(n716), .A2(n715), .Y(n_sram_raddr_b1[9]) );
  AO22X1_HVT U954 ( .A1(n191), .A2(n420), .A3(n1320), .A4(n252), .Y(n717) );
  AO221X1_HVT U955 ( .A1(sram_raddr_b2[0]), .A2(n1332), .A3(n287), .A4(n788), 
        .A5(n717), .Y(n718) );
  AO22X1_HVT U956 ( .A1(n207), .A2(n718), .A3(sram_raddr_b2[0]), .A4(n168), 
        .Y(n_sram_raddr_b2[0]) );
  NAND2X0_HVT U957 ( .A1(sram_raddr_b5[0]), .A2(sram_raddr_b5[1]), .Y(n732) );
  NAND2X0_HVT U958 ( .A1(n252), .A2(n373), .Y(n1291) );
  NAND2X0_HVT U959 ( .A1(n732), .A2(n1291), .Y(n1265) );
  OA22X1_HVT U960 ( .A1(n982), .A2(n370), .A3(n227), .A4(n1265), .Y(n720) );
  NAND2X0_HVT U961 ( .A1(sram_raddr_b8[1]), .A2(sram_raddr_b8[0]), .Y(n729) );
  OA21X1_HVT U962 ( .A1(sram_raddr_b8[1]), .A2(sram_raddr_b8[0]), .A3(n729), 
        .Y(n1264) );
  NAND2X0_HVT U963 ( .A1(n191), .A2(n1264), .Y(n985) );
  NAND2X0_HVT U964 ( .A1(sram_raddr_b2[0]), .A2(sram_raddr_b2[1]), .Y(n983) );
  NAND2X0_HVT U965 ( .A1(n287), .A2(n370), .Y(n1005) );
  NAND3X0_HVT U966 ( .A1(n788), .A2(n983), .A3(n1005), .Y(n719) );
  NAND3X0_HVT U967 ( .A1(n720), .A2(n985), .A3(n719), .Y(n721) );
  AO22X1_HVT U968 ( .A1(n206), .A2(n721), .A3(sram_raddr_b2[1]), .A4(n217), 
        .Y(n_sram_raddr_b2[1]) );
  NAND2X0_HVT U969 ( .A1(n334), .A2(n983), .Y(n735) );
  OA22X1_HVT U970 ( .A1(sram_raddr_b2[2]), .A2(n1299), .A3(n745), .A4(n735), 
        .Y(n728) );
  AO22X1_HVT U971 ( .A1(sram_raddr_b8[2]), .A2(n723), .A3(n245), .A4(n729), 
        .Y(n1271) );
  NAND2X0_HVT U972 ( .A1(n190), .A2(n1271), .Y(n988) );
  AO221X1_HVT U973 ( .A1(n213), .A2(n745), .A3(n214), .A4(n983), .A5(n334), 
        .Y(n724) );
  NAND3X0_HVT U974 ( .A1(n728), .A2(n988), .A3(n724), .Y(n726) );
  AO22X1_HVT U975 ( .A1(sram_raddr_b5[2]), .A2(n725), .A3(n321), .A4(n732), 
        .Y(n990) );
  OA221X1_HVT U976 ( .A1(n726), .A2(n178), .A3(n726), .A4(n990), .A5(n207), 
        .Y(n727) );
  AO221X1_HVT U977 ( .A1(sram_raddr_b2[2]), .A2(n232), .A3(n334), .A4(n224), 
        .A5(n727), .Y(n_sram_raddr_b2[2]) );
  NAND2X0_HVT U978 ( .A1(n215), .A2(n728), .Y(n731) );
  OA221X1_HVT U979 ( .A1(n788), .A2(sram_raddr_b2[2]), .A3(n788), .A4(n1318), 
        .A5(n735), .Y(n730) );
  NAND2X0_HVT U980 ( .A1(n245), .A2(n729), .Y(n1275) );
  NAND2X0_HVT U981 ( .A1(sram_raddr_b8[3]), .A2(n1275), .Y(n1274) );
  AO221X1_HVT U982 ( .A1(sram_raddr_b2[3]), .A2(n731), .A3(n426), .A4(n730), 
        .A5(n997), .Y(n734) );
  NAND2X0_HVT U983 ( .A1(n321), .A2(n732), .Y(n733) );
  NAND2X0_HVT U984 ( .A1(sram_raddr_b5[3]), .A2(n733), .Y(n737) );
  OA21X1_HVT U985 ( .A1(sram_raddr_b5[3]), .A2(n733), .A3(n737), .Y(n996) );
  NAND2X0_HVT U986 ( .A1(sram_raddr_b2[3]), .A2(sram_raddr_b2[2]), .Y(n1002)
         );
  NAND2X0_HVT U987 ( .A1(n264), .A2(n1002), .Y(n743) );
  NAND3X0_HVT U988 ( .A1(sram_raddr_b2[4]), .A2(sram_raddr_b2[3]), .A3(
        sram_raddr_b2[2]), .Y(n764) );
  NAND2X0_HVT U989 ( .A1(n743), .A2(n764), .Y(n740) );
  NAND2X0_HVT U990 ( .A1(sram_raddr_b2[3]), .A2(n735), .Y(n757) );
  AND2X1_HVT U991 ( .A1(n264), .A2(n757), .Y(n736) );
  AO22X1_HVT U992 ( .A1(n1318), .A2(n740), .A3(n736), .A4(n788), .Y(n750) );
  OA21X1_HVT U993 ( .A1(n745), .A2(n757), .A3(n213), .Y(n746) );
  NAND2X0_HVT U994 ( .A1(n324), .A2(n737), .Y(n747) );
  OA21X1_HVT U995 ( .A1(n737), .A2(n324), .A3(n747), .Y(n1006) );
  OA22X1_HVT U996 ( .A1(n746), .A2(n264), .A3(n1006), .A4(n173), .Y(n738) );
  NAND2X0_HVT U997 ( .A1(n346), .A2(n1274), .Y(n751) );
  NAND2X0_HVT U998 ( .A1(n191), .A2(n1287), .Y(n1008) );
  NAND3X0_HVT U999 ( .A1(n739), .A2(n738), .A3(n1008), .Y(n742) );
  AO222X1_HVT U1000 ( .A1(n742), .A2(n205), .A3(n234), .A4(sram_raddr_b2[4]), 
        .A5(n179), .A6(n741), .Y(n_sram_raddr_b2[4]) );
  NAND2X0_HVT U1001 ( .A1(n319), .A2(n743), .Y(n744) );
  NAND2X0_HVT U1002 ( .A1(n748), .A2(n266), .Y(n756) );
  OA21X1_HVT U1003 ( .A1(n748), .A2(n266), .A3(n756), .Y(n1015) );
  OA22X1_HVT U1004 ( .A1(n749), .A2(n318), .A3(n1015), .A4(n173), .Y(n752) );
  NAND3X0_HVT U1005 ( .A1(n318), .A2(n764), .A3(n750), .Y(n758) );
  AO22X1_HVT U1006 ( .A1(sram_raddr_b8[5]), .A2(n751), .A3(n325), .A4(n759), 
        .Y(n1300) );
  NAND2X0_HVT U1007 ( .A1(n190), .A2(n1300), .Y(n1014) );
  NAND3X0_HVT U1008 ( .A1(n752), .A2(n758), .A3(n1014), .Y(n753) );
  AO22X1_HVT U1009 ( .A1(n204), .A2(n753), .A3(n233), .A4(sram_raddr_b2[5]), 
        .Y(n755) );
  NAND4X0_HVT U1010 ( .A1(sram_raddr_b2[5]), .A2(sram_raddr_b2[4]), .A3(
        sram_raddr_b2[3]), .A4(sram_raddr_b2[2]), .Y(n763) );
  NAND2X0_HVT U1011 ( .A1(n318), .A2(n764), .Y(n754) );
  OA222X1_HVT U1012 ( .A1(n755), .A2(n225), .A3(n755), .A4(n763), .A5(n755), 
        .A6(n754), .Y(n_sram_raddr_b2[5]) );
  NAND2X0_HVT U1013 ( .A1(sram_raddr_b5[6]), .A2(n756), .Y(n769) );
  OA21X1_HVT U1014 ( .A1(sram_raddr_b5[6]), .A2(n756), .A3(n769), .Y(n1019) );
  NAND2X0_HVT U1015 ( .A1(n1019), .A2(n1320), .Y(n762) );
  NAND3X0_HVT U1016 ( .A1(n318), .A2(n264), .A3(n1002), .Y(n772) );
  NAND3X0_HVT U1017 ( .A1(n318), .A2(n264), .A3(n757), .Y(n773) );
  AOI22X1_HVT U1018 ( .A1(n1318), .A2(n772), .A3(n788), .A4(n773), .Y(n768) );
  OA222X1_HVT U1019 ( .A1(n390), .A2(n213), .A3(n390), .A4(n758), .A5(
        sram_raddr_b2[6]), .A6(n768), .Y(n761) );
  NAND2X0_HVT U1020 ( .A1(n759), .A2(n325), .Y(n760) );
  NAND2X0_HVT U1021 ( .A1(sram_raddr_b8[6]), .A2(n760), .Y(n770) );
  OA21X1_HVT U1022 ( .A1(sram_raddr_b8[6]), .A2(n760), .A3(n770), .Y(n1308) );
  NAND2X0_HVT U1023 ( .A1(n190), .A2(n1308), .Y(n1031) );
  NAND3X0_HVT U1024 ( .A1(n762), .A2(n761), .A3(n1031), .Y(n767) );
  AO221X1_HVT U1025 ( .A1(n225), .A2(n390), .A3(n188), .A4(n763), .A5(n234), 
        .Y(n781) );
  NAND3X0_HVT U1026 ( .A1(n223), .A2(sram_raddr_b2[5]), .A3(n1004), .Y(n765)
         );
  NAND2X0_HVT U1027 ( .A1(n390), .A2(n765), .Y(n766) );
  AO22X1_HVT U1028 ( .A1(n206), .A2(n767), .A3(n781), .A4(n766), .Y(
        n_sram_raddr_b2[6]) );
  AND4X1_HVT U1029 ( .A1(n188), .A2(sram_raddr_b2[6]), .A3(sram_raddr_b2[5]), 
        .A4(n1004), .Y(n799) );
  OA21X1_HVT U1030 ( .A1(n768), .A2(n390), .A3(n216), .Y(n776) );
  NAND2X0_HVT U1031 ( .A1(n354), .A2(n769), .Y(n790) );
  OA21X1_HVT U1032 ( .A1(n769), .A2(n354), .A3(n790), .Y(n1036) );
  OA22X1_HVT U1033 ( .A1(n776), .A2(n260), .A3(n1036), .A4(n226), .Y(n771) );
  NAND2X0_HVT U1034 ( .A1(n269), .A2(n770), .Y(n793) );
  NAND2X0_HVT U1035 ( .A1(n191), .A2(n1313), .Y(n1038) );
  NAND2X0_HVT U1036 ( .A1(n771), .A2(n1038), .Y(n774) );
  NAND2X0_HVT U1037 ( .A1(sram_raddr_b2[6]), .A2(n772), .Y(n785) );
  NAND2X0_HVT U1038 ( .A1(sram_raddr_b2[6]), .A2(n773), .Y(n784) );
  AO22X1_HVT U1039 ( .A1(n1318), .A2(n785), .A3(n788), .A4(n784), .Y(n777) );
  OA221X1_HVT U1040 ( .A1(n774), .A2(n260), .A3(n774), .A4(n777), .A5(n207), 
        .Y(n775) );
  AO221X1_HVT U1041 ( .A1(sram_raddr_b2[7]), .A2(n781), .A3(n260), .A4(n799), 
        .A5(n775), .Y(n_sram_raddr_b2[7]) );
  HADDX1_HVT U1042 ( .A0(sram_raddr_b5[8]), .B0(n790), .SO(n1048) );
  OA22X1_HVT U1043 ( .A1(n1048), .A2(n226), .A3(n776), .A4(n401), .Y(n780) );
  HADDX1_HVT U1044 ( .A0(n337), .B0(n793), .SO(n1327) );
  NAND2X0_HVT U1045 ( .A1(n191), .A2(n1327), .Y(n1046) );
  NAND3X0_HVT U1046 ( .A1(n401), .A2(n260), .A3(n777), .Y(n792) );
  NAND3X0_HVT U1047 ( .A1(sram_raddr_b2[8]), .A2(sram_raddr_b2[7]), .A3(n778), 
        .Y(n779) );
  NAND4X0_HVT U1048 ( .A1(n780), .A2(n1046), .A3(n792), .A4(n779), .Y(n783) );
  AO21X1_HVT U1049 ( .A1(sram_raddr_b2[7]), .A2(n799), .A3(sram_raddr_b2[8]), 
        .Y(n782) );
  NAND2X0_HVT U1050 ( .A1(sram_raddr_b2[8]), .A2(sram_raddr_b2[7]), .Y(n797)
         );
  AO21X1_HVT U1051 ( .A1(n188), .A2(n797), .A3(n781), .Y(n798) );
  AO22X1_HVT U1052 ( .A1(n203), .A2(n783), .A3(n782), .A4(n798), .Y(
        n_sram_raddr_b2[8]) );
  NAND3X0_HVT U1053 ( .A1(n401), .A2(n260), .A3(n784), .Y(n787) );
  NAND4X0_HVT U1054 ( .A1(n214), .A2(n260), .A3(n401), .A4(n785), .Y(n786) );
  AO22X1_HVT U1055 ( .A1(n788), .A2(n787), .A3(n1332), .A4(n786), .Y(n789) );
  NAND2X0_HVT U1056 ( .A1(sram_raddr_b2[9]), .A2(n789), .Y(n796) );
  OR2X1_HVT U1057 ( .A1(n790), .A2(sram_raddr_b5[8]), .Y(n791) );
  HADDX1_HVT U1058 ( .A0(sram_raddr_b5[9]), .B0(n791), .SO(n1070) );
  OA22X1_HVT U1059 ( .A1(sram_raddr_b2[9]), .A2(n792), .A3(n227), .A4(n1070), 
        .Y(n795) );
  OR2X1_HVT U1060 ( .A1(n793), .A2(sram_raddr_b8[8]), .Y(n794) );
  HADDX1_HVT U1061 ( .A0(n794), .B0(n407), .SO(n1337) );
  NAND2X0_HVT U1062 ( .A1(n190), .A2(n1337), .Y(n1069) );
  NAND3X0_HVT U1063 ( .A1(n796), .A2(n795), .A3(n1069), .Y(n802) );
  OA222X1_HVT U1064 ( .A1(sram_raddr_b2[9]), .A2(n800), .A3(sram_raddr_b2[9]), 
        .A4(n799), .A5(n434), .A6(n798), .Y(n801) );
  AO21X1_HVT U1065 ( .A1(n204), .A2(n802), .A3(n801), .Y(n_sram_raddr_b2[9])
         );
  NAND2X0_HVT U1066 ( .A1(n1078), .A2(n173), .Y(n864) );
  AO22X1_HVT U1067 ( .A1(n192), .A2(n418), .A3(n1260), .A4(n250), .Y(n803) );
  AO221X1_HVT U1068 ( .A1(sram_raddr_b3[0]), .A2(n1084), .A3(n285), .A4(n864), 
        .A5(n803), .Y(n804) );
  AO22X1_HVT U1069 ( .A1(n204), .A2(n804), .A3(sram_raddr_b3[0]), .A4(n217), 
        .Y(n_sram_raddr_b3[0]) );
  OA22X1_HVT U1070 ( .A1(n886), .A2(n1083), .A3(n1158), .A4(n367), .Y(n808) );
  NAND2X0_HVT U1071 ( .A1(n805), .A2(n830), .Y(n806) );
  NAND2X0_HVT U1072 ( .A1(n1260), .A2(n806), .Y(n1081) );
  NAND3X0_HVT U1073 ( .A1(n808), .A2(n807), .A3(n1081), .Y(n809) );
  AO22X1_HVT U1074 ( .A1(n203), .A2(n809), .A3(sram_raddr_b3[1]), .A4(n168), 
        .Y(n_sram_raddr_b3[1]) );
  OA22X1_HVT U1075 ( .A1(sram_raddr_b3[2]), .A2(n1125), .A3(n810), .A4(n1078), 
        .Y(n812) );
  NAND2X0_HVT U1076 ( .A1(sram_raddr_b3[2]), .A2(n1306), .Y(n811) );
  AO221X1_HVT U1077 ( .A1(sram_raddr_b0[2]), .A2(n830), .A3(n279), .A4(n828), 
        .A5(n220), .Y(n1086) );
  NAND4X0_HVT U1078 ( .A1(n813), .A2(n812), .A3(n811), .A4(n1086), .Y(n816) );
  NAND2X0_HVT U1079 ( .A1(n188), .A2(n326), .Y(n814) );
  NAND2X0_HVT U1080 ( .A1(n1303), .A2(n814), .Y(n825) );
  NAND2X0_HVT U1081 ( .A1(n326), .A2(n1366), .Y(n815) );
  AO22X1_HVT U1082 ( .A1(n204), .A2(n816), .A3(n825), .A4(n815), .Y(
        n_sram_raddr_b3[2]) );
  OA21X1_HVT U1083 ( .A1(sram_raddr_b3[2]), .A2(n1125), .A3(n215), .Y(n817) );
  OA22X1_HVT U1084 ( .A1(n886), .A2(n818), .A3(n817), .A4(n393), .Y(n822) );
  OA222X1_HVT U1085 ( .A1(sram_raddr_b0[3]), .A2(sram_raddr_b0[2]), .A3(
        sram_raddr_b0[3]), .A4(n830), .A5(n828), .A6(n827), .Y(n819) );
  NAND2X0_HVT U1086 ( .A1(n1260), .A2(n819), .Y(n1100) );
  NAND3X0_HVT U1087 ( .A1(sram_raddr_b3[2]), .A2(n393), .A3(n1148), .Y(n820)
         );
  NAND4X0_HVT U1088 ( .A1(n822), .A2(n821), .A3(n1100), .A4(n820), .Y(n824) );
  AND2X1_HVT U1089 ( .A1(sram_raddr_b3[2]), .A2(n393), .Y(n823) );
  AO222X1_HVT U1090 ( .A1(n825), .A2(sram_raddr_b3[3]), .A3(n824), .A4(n205), 
        .A5(n823), .A6(n224), .Y(n_sram_raddr_b3[3]) );
  NAND3X0_HVT U1091 ( .A1(sram_raddr_b3[3]), .A2(sram_raddr_b3[2]), .A3(
        sram_raddr_b3[4]), .Y(n844) );
  NAND2X0_HVT U1092 ( .A1(sram_raddr_b3[3]), .A2(sram_raddr_b3[2]), .Y(n1106)
         );
  NAND2X0_HVT U1093 ( .A1(n320), .A2(n1106), .Y(n826) );
  AND2X1_HVT U1094 ( .A1(n844), .A2(n826), .Y(n835) );
  OA22X1_HVT U1095 ( .A1(n1125), .A2(n835), .A3(n215), .A4(n320), .Y(n834) );
  OA21X1_HVT U1096 ( .A1(n828), .A2(n827), .A3(n323), .Y(n839) );
  OAI221X1_HVT U1097 ( .A1(n839), .A2(n830), .A3(n839), .A4(n829), .A5(n1260), 
        .Y(n1112) );
  OR2X1_HVT U1098 ( .A1(n886), .A2(n831), .Y(n832) );
  NAND4X0_HVT U1099 ( .A1(n834), .A2(n833), .A3(n1112), .A4(n832), .Y(n836) );
  AO222X1_HVT U1100 ( .A1(n836), .A2(n206), .A3(n232), .A4(sram_raddr_b3[4]), 
        .A5(n225), .A6(n835), .Y(n_sram_raddr_b3[4]) );
  OA221X1_HVT U1101 ( .A1(n1387), .A2(n320), .A3(n1387), .A4(n1106), .A5(n215), 
        .Y(n837) );
  OA22X1_HVT U1102 ( .A1(n886), .A2(n838), .A3(n261), .A4(n837), .Y(n842) );
  NAND3X0_HVT U1103 ( .A1(n261), .A2(n320), .A3(n1106), .Y(n857) );
  OR2X1_HVT U1104 ( .A1(n857), .A2(n1125), .Y(n840) );
  NAND2X0_HVT U1105 ( .A1(n839), .A2(n272), .Y(n847) );
  AO221X1_HVT U1106 ( .A1(n847), .A2(n839), .A3(n847), .A4(n272), .A5(n220), 
        .Y(n1119) );
  AND4X1_HVT U1107 ( .A1(n842), .A2(n841), .A3(n840), .A4(n1119), .Y(n843) );
  OA22X1_HVT U1108 ( .A1(n843), .A2(n221), .A3(n1303), .A4(n261), .Y(n846) );
  AO221X1_HVT U1109 ( .A1(sram_raddr_b3[5]), .A2(n1108), .A3(n261), .A4(n844), 
        .A5(n1366), .Y(n845) );
  NAND2X0_HVT U1110 ( .A1(n846), .A2(n845), .Y(n_sram_raddr_b3[5]) );
  NAND2X0_HVT U1111 ( .A1(sram_raddr_b0[6]), .A2(n847), .Y(n858) );
  NAND2X0_HVT U1112 ( .A1(n1260), .A2(n858), .Y(n850) );
  OA221X1_HVT U1113 ( .A1(n850), .A2(n849), .A3(n850), .A4(n391), .A5(n848), 
        .Y(n1130) );
  AO221X1_HVT U1114 ( .A1(n213), .A2(n1125), .A3(n216), .A4(n857), .A5(n400), 
        .Y(n854) );
  NAND2X0_HVT U1115 ( .A1(n851), .A2(n864), .Y(n853) );
  NAND3X0_HVT U1116 ( .A1(n1148), .A2(n400), .A3(n857), .Y(n852) );
  NAND4X0_HVT U1117 ( .A1(n1130), .A2(n854), .A3(n853), .A4(n852), .Y(n856) );
  NAND4X0_HVT U1118 ( .A1(sram_raddr_b3[6]), .A2(sram_raddr_b3[5]), .A3(n1108), 
        .A4(n1303), .Y(n875) );
  AND2X1_HVT U1119 ( .A1(n168), .A2(n875), .Y(n867) );
  OA222X1_HVT U1120 ( .A1(sram_raddr_b3[6]), .A2(n225), .A3(sram_raddr_b3[6]), 
        .A4(sram_raddr_b3[5]), .A5(sram_raddr_b3[6]), .A6(n1108), .Y(n855) );
  AO22X1_HVT U1121 ( .A1(n205), .A2(n856), .A3(n867), .A4(n855), .Y(
        n_sram_raddr_b3[6]) );
  AND4X1_HVT U1122 ( .A1(n188), .A2(sram_raddr_b3[6]), .A3(sram_raddr_b3[5]), 
        .A4(n1108), .Y(n888) );
  NAND2X0_HVT U1123 ( .A1(sram_raddr_b3[6]), .A2(n857), .Y(n871) );
  NAND3X0_HVT U1124 ( .A1(n1148), .A2(n350), .A3(n871), .Y(n861) );
  NAND2X0_HVT U1125 ( .A1(n263), .A2(n858), .Y(n868) );
  AO221X1_HVT U1126 ( .A1(n868), .A2(n858), .A3(n868), .A4(n263), .A5(n220), 
        .Y(n1141) );
  AO221X1_HVT U1127 ( .A1(n214), .A2(n1387), .A3(n213), .A4(n871), .A5(n350), 
        .Y(n859) );
  NAND4X0_HVT U1128 ( .A1(n861), .A2(n860), .A3(n1141), .A4(n859), .Y(n865) );
  OA221X1_HVT U1129 ( .A1(n865), .A2(n864), .A3(n865), .A4(n863), .A5(n207), 
        .Y(n866) );
  AO221X1_HVT U1130 ( .A1(sram_raddr_b3[7]), .A2(n867), .A3(n350), .A4(n888), 
        .A5(n866), .Y(n_sram_raddr_b3[7]) );
  NAND2X0_HVT U1131 ( .A1(n869), .A2(n329), .Y(n881) );
  AO221X1_HVT U1132 ( .A1(n881), .A2(n869), .A3(n881), .A4(n329), .A5(n220), 
        .Y(n1154) );
  OA21X1_HVT U1133 ( .A1(n870), .A2(n886), .A3(n1154), .Y(n874) );
  NAND4X0_HVT U1134 ( .A1(n1148), .A2(n268), .A3(n350), .A4(n871), .Y(n883) );
  AND3X1_HVT U1135 ( .A1(n214), .A2(n350), .A3(n871), .Y(n880) );
  OR3X1_HVT U1136 ( .A1(n1158), .A2(n880), .A3(n268), .Y(n872) );
  NAND4X0_HVT U1137 ( .A1(n874), .A2(n873), .A3(n883), .A4(n872), .Y(n879) );
  OR3X1_HVT U1138 ( .A1(n350), .A2(n875), .A3(n268), .Y(n876) );
  NAND2X0_HVT U1139 ( .A1(n876), .A2(n168), .Y(n887) );
  AO21X1_HVT U1140 ( .A1(sram_raddr_b3[7]), .A2(n888), .A3(sram_raddr_b3[8]), 
        .Y(n877) );
  AO22X1_HVT U1141 ( .A1(n205), .A2(n879), .A3(n878), .A4(n877), .Y(
        n_sram_raddr_b3[8]) );
  AO221X1_HVT U1142 ( .A1(sram_raddr_b0[9]), .A2(n882), .A3(n423), .A4(n881), 
        .A5(n219), .Y(n1168) );
  NAND2X0_HVT U1143 ( .A1(n1174), .A2(n173), .Y(n961) );
  AO22X1_HVT U1144 ( .A1(n190), .A2(n419), .A3(n1260), .A4(n251), .Y(n889) );
  AO221X1_HVT U1145 ( .A1(sram_raddr_b4[0]), .A2(n1236), .A3(n286), .A4(n961), 
        .A5(n889), .Y(n890) );
  AO22X1_HVT U1146 ( .A1(n207), .A2(n890), .A3(sram_raddr_b4[0]), .A4(n168), 
        .Y(n_sram_raddr_b4[0]) );
  OA22X1_HVT U1147 ( .A1(n891), .A2(n372), .A3(n974), .A4(n1179), .Y(n895) );
  NAND2X0_HVT U1148 ( .A1(n892), .A2(n897), .Y(n893) );
  NAND2X0_HVT U1149 ( .A1(n1260), .A2(n893), .Y(n1177) );
  NAND3X0_HVT U1150 ( .A1(n895), .A2(n894), .A3(n1177), .Y(n896) );
  AO22X1_HVT U1151 ( .A1(n207), .A2(n896), .A3(sram_raddr_b4[1]), .A4(n168), 
        .Y(n_sram_raddr_b4[1]) );
  AO21X1_HVT U1152 ( .A1(n205), .A2(n1306), .A3(n232), .Y(n1560) );
  AND2X1_HVT U1153 ( .A1(sram_raddr_b1[2]), .A2(n897), .Y(n905) );
  NAND2X0_HVT U1154 ( .A1(n1226), .A2(n322), .Y(n904) );
  NAND3X0_HVT U1155 ( .A1(n898), .A2(n1183), .A3(n904), .Y(n901) );
  OA221X1_HVT U1156 ( .A1(n901), .A2(n961), .A3(n901), .A4(n900), .A5(n203), 
        .Y(n902) );
  AO221X1_HVT U1157 ( .A1(sram_raddr_b4[2]), .A2(n1560), .A3(n322), .A4(n223), 
        .A5(n902), .Y(n_sram_raddr_b4[2]) );
  NAND3X0_HVT U1158 ( .A1(n1226), .A2(sram_raddr_b4[2]), .A3(n389), .Y(n903)
         );
  OA221X1_HVT U1159 ( .A1(n389), .A2(n216), .A3(n389), .A4(n904), .A5(n903), 
        .Y(n910) );
  OR2X1_HVT U1160 ( .A1(n974), .A2(n906), .Y(n907) );
  NAND4X0_HVT U1161 ( .A1(n910), .A2(n909), .A3(n908), .A4(n907), .Y(n914) );
  NAND2X0_HVT U1162 ( .A1(n225), .A2(n322), .Y(n911) );
  NAND2X0_HVT U1163 ( .A1(n1303), .A2(n911), .Y(n913) );
  AND2X1_HVT U1164 ( .A1(sram_raddr_b4[2]), .A2(n389), .Y(n912) );
  AO222X1_HVT U1165 ( .A1(n914), .A2(n207), .A3(n913), .A4(sram_raddr_b4[3]), 
        .A5(n912), .A6(n188), .Y(n_sram_raddr_b4[3]) );
  NAND3X0_HVT U1166 ( .A1(sram_raddr_b4[3]), .A2(sram_raddr_b4[2]), .A3(
        sram_raddr_b4[4]), .Y(n932) );
  NAND2X0_HVT U1167 ( .A1(sram_raddr_b4[3]), .A2(sram_raddr_b4[2]), .Y(n1200)
         );
  NAND2X0_HVT U1168 ( .A1(n336), .A2(n1200), .Y(n925) );
  AND2X1_HVT U1169 ( .A1(n932), .A2(n925), .Y(n922) );
  OA22X1_HVT U1170 ( .A1(n974), .A2(n915), .A3(n922), .A4(n1198), .Y(n921) );
  OA21X1_HVT U1171 ( .A1(n918), .A2(n916), .A3(n335), .Y(n924) );
  AO221X1_HVT U1172 ( .A1(n919), .A2(n918), .A3(n919), .A4(n917), .A5(n220), 
        .Y(n1206) );
  NAND3X0_HVT U1173 ( .A1(n921), .A2(n920), .A3(n1206), .Y(n923) );
  AO222X1_HVT U1174 ( .A1(n923), .A2(n205), .A3(n1560), .A4(sram_raddr_b4[4]), 
        .A5(n922), .A6(n225), .Y(n_sram_raddr_b4[4]) );
  NAND3X0_HVT U1175 ( .A1(n271), .A2(n336), .A3(n1200), .Y(n944) );
  OR2X1_HVT U1176 ( .A1(n1198), .A2(n944), .Y(n927) );
  NAND2X0_HVT U1177 ( .A1(n924), .A2(n265), .Y(n933) );
  AO221X1_HVT U1178 ( .A1(n933), .A2(n924), .A3(n933), .A4(n265), .A5(n220), 
        .Y(n1211) );
  OAI221X1_HVT U1179 ( .A1(n1306), .A2(n262), .A3(n1306), .A4(n925), .A5(
        sram_raddr_b4[5]), .Y(n926) );
  NAND4X0_HVT U1180 ( .A1(n928), .A2(n927), .A3(n1211), .A4(n926), .Y(n931) );
  NAND2X0_HVT U1181 ( .A1(sram_raddr_b1[6]), .A2(n933), .Y(n942) );
  OR2X1_HVT U1182 ( .A1(n974), .A2(n934), .Y(n937) );
  AO221X1_HVT U1183 ( .A1(n215), .A2(n1198), .A3(n214), .A4(n944), .A5(n415), 
        .Y(n936) );
  NAND3X0_HVT U1184 ( .A1(n1226), .A2(n415), .A3(n944), .Y(n935) );
  NAND4X0_HVT U1185 ( .A1(n938), .A2(n937), .A3(n936), .A4(n935), .Y(n941) );
  NAND3X0_HVT U1186 ( .A1(sram_raddr_b4[6]), .A2(sram_raddr_b4[5]), .A3(n1202), 
        .Y(n948) );
  OA221X1_HVT U1187 ( .A1(sram_raddr_b4[6]), .A2(sram_raddr_b4[5]), .A3(
        sram_raddr_b4[6]), .A4(n1202), .A5(n948), .Y(n939) );
  AO22X1_HVT U1188 ( .A1(n224), .A2(n939), .A3(n234), .A4(sram_raddr_b4[6]), 
        .Y(n940) );
  AO221X1_HVT U1189 ( .A1(n207), .A2(n1224), .A3(n203), .A4(n941), .A5(n940), 
        .Y(n_sram_raddr_b4[6]) );
  NAND2X0_HVT U1190 ( .A1(n317), .A2(n942), .Y(n955) );
  AO221X1_HVT U1191 ( .A1(n955), .A2(n942), .A3(n955), .A4(n317), .A5(n220), 
        .Y(n1228) );
  OA21X1_HVT U1192 ( .A1(n974), .A2(n943), .A3(n1228), .Y(n947) );
  NAND2X0_HVT U1193 ( .A1(sram_raddr_b4[6]), .A2(n944), .Y(n966) );
  NAND3X0_HVT U1194 ( .A1(n1226), .A2(n316), .A3(n966), .Y(n957) );
  AO221X1_HVT U1195 ( .A1(n213), .A2(col[0]), .A3(n213), .A4(n966), .A5(n316), 
        .Y(n945) );
  NAND4X0_HVT U1196 ( .A1(n947), .A2(n957), .A3(n946), .A4(n945), .Y(n952) );
  NAND2X0_HVT U1197 ( .A1(n316), .A2(n948), .Y(n951) );
  NAND2X0_HVT U1198 ( .A1(sram_raddr_b4[7]), .A2(n954), .Y(n949) );
  NAND2X0_HVT U1199 ( .A1(n224), .A2(n949), .Y(n953) );
  AO222X1_HVT U1200 ( .A1(n952), .A2(n207), .A3(n951), .A4(n950), .A5(
        sram_raddr_b4[7]), .A6(n232), .Y(n_sram_raddr_b4[7]) );
  AND3X1_HVT U1201 ( .A1(n223), .A2(sram_raddr_b4[7]), .A3(n954), .Y(n965) );
  OR2X1_HVT U1202 ( .A1(n957), .A2(sram_raddr_b4[8]), .Y(n971) );
  NAND2X0_HVT U1203 ( .A1(n956), .A2(n267), .Y(n968) );
  AO221X1_HVT U1204 ( .A1(n968), .A2(n956), .A3(n968), .A4(n267), .A5(n220), 
        .Y(n1239) );
  NAND3X0_HVT U1205 ( .A1(n1236), .A2(n957), .A3(sram_raddr_b4[8]), .Y(n958)
         );
  NAND4X0_HVT U1206 ( .A1(n971), .A2(n959), .A3(n1239), .A4(n958), .Y(n962) );
  OA221X1_HVT U1207 ( .A1(n962), .A2(n961), .A3(n962), .A4(n960), .A5(n204), 
        .Y(n963) );
  AO221X1_HVT U1208 ( .A1(n964), .A2(sram_raddr_b4[8]), .A3(n964), .A4(n965), 
        .A5(n963), .Y(n_sram_raddr_b4[8]) );
  NAND3X0_HVT U1209 ( .A1(n395), .A2(n965), .A3(sram_raddr_b4[8]), .Y(n979) );
  AND2X1_HVT U1210 ( .A1(n316), .A2(n966), .Y(n967) );
  OA221X1_HVT U1211 ( .A1(n1198), .A2(n967), .A3(n1198), .A4(n328), .A5(n213), 
        .Y(n970) );
  OA221X1_HVT U1212 ( .A1(sram_raddr_b4[9]), .A2(n971), .A3(n395), .A4(n970), 
        .A5(n1243), .Y(n975) );
  OA22X1_HVT U1213 ( .A1(n977), .A2(n395), .A3(n976), .A4(n221), .Y(n978) );
  NAND2X0_HVT U1214 ( .A1(n979), .A2(n978), .Y(n_sram_raddr_b4[9]) );
  NAND2X0_HVT U1215 ( .A1(n227), .A2(n1326), .Y(n1018) );
  AO22X1_HVT U1216 ( .A1(n190), .A2(n420), .A3(n1260), .A4(n287), .Y(n980) );
  AO221X1_HVT U1217 ( .A1(sram_raddr_b5[0]), .A2(n1332), .A3(n252), .A4(n1018), 
        .A5(n980), .Y(n981) );
  AO22X1_HVT U1218 ( .A1(n205), .A2(n981), .A3(sram_raddr_b5[0]), .A4(n217), 
        .Y(n_sram_raddr_b5[0]) );
  OA22X1_HVT U1219 ( .A1(n982), .A2(n373), .A3(n1071), .A4(n1265), .Y(n986) );
  NAND2X0_HVT U1220 ( .A1(n983), .A2(n1005), .Y(n984) );
  NAND2X0_HVT U1221 ( .A1(n1260), .A2(n984), .Y(n1263) );
  NAND3X0_HVT U1222 ( .A1(n986), .A2(n985), .A3(n1263), .Y(n987) );
  AO22X1_HVT U1223 ( .A1(n206), .A2(n987), .A3(sram_raddr_b5[1]), .A4(n217), 
        .Y(n_sram_raddr_b5[1]) );
  AO22X1_HVT U1224 ( .A1(sram_raddr_b5[2]), .A2(n215), .A3(n321), .A4(n1299), 
        .Y(n989) );
  AO221X1_HVT U1225 ( .A1(sram_raddr_b2[2]), .A2(n1005), .A3(n334), .A4(n1003), 
        .A5(n220), .Y(n1269) );
  NAND3X0_HVT U1226 ( .A1(n989), .A2(n988), .A3(n1269), .Y(n991) );
  OA221X1_HVT U1227 ( .A1(n991), .A2(n1018), .A3(n991), .A4(n990), .A5(n1557), 
        .Y(n992) );
  AO221X1_HVT U1228 ( .A1(sram_raddr_b5[2]), .A2(n234), .A3(n321), .A4(n188), 
        .A5(n992), .Y(n_sram_raddr_b5[2]) );
  OA222X1_HVT U1229 ( .A1(sram_raddr_b2[3]), .A2(sram_raddr_b2[2]), .A3(
        sram_raddr_b2[3]), .A4(n1005), .A5(n1003), .A6(n1002), .Y(n993) );
  NAND2X0_HVT U1230 ( .A1(n1260), .A2(n993), .Y(n1280) );
  AO221X1_HVT U1231 ( .A1(n214), .A2(sram_raddr_b5[2]), .A3(n216), .A4(n1299), 
        .A5(n413), .Y(n995) );
  NAND3X0_HVT U1232 ( .A1(sram_raddr_b5[2]), .A2(n1318), .A3(n413), .Y(n994)
         );
  NAND2X0_HVT U1233 ( .A1(n224), .A2(n321), .Y(n998) );
  NAND2X0_HVT U1234 ( .A1(n1303), .A2(n998), .Y(n1000) );
  AND2X1_HVT U1235 ( .A1(sram_raddr_b5[2]), .A2(n413), .Y(n999) );
  AO222X1_HVT U1236 ( .A1(n1001), .A2(n207), .A3(n1000), .A4(sram_raddr_b5[3]), 
        .A5(n999), .A6(n224), .Y(n_sram_raddr_b5[3]) );
  NAND3X0_HVT U1237 ( .A1(sram_raddr_b5[4]), .A2(sram_raddr_b5[3]), .A3(
        sram_raddr_b5[2]), .Y(n1016) );
  NAND2X0_HVT U1238 ( .A1(sram_raddr_b5[3]), .A2(sram_raddr_b5[2]), .Y(n1288)
         );
  NAND2X0_HVT U1239 ( .A1(n324), .A2(n1288), .Y(n1013) );
  AND2X1_HVT U1240 ( .A1(n1016), .A2(n1013), .Y(n1010) );
  OA22X1_HVT U1241 ( .A1(n213), .A2(n324), .A3(n1010), .A4(n1299), .Y(n1009)
         );
  OA21X1_HVT U1242 ( .A1(n1003), .A2(n1002), .A3(n264), .Y(n1012) );
  OAI221X1_HVT U1243 ( .A1(n1012), .A2(n1005), .A3(n1012), .A4(n1004), .A5(
        n1260), .Y(n1294) );
  OR2X1_HVT U1244 ( .A1(n1071), .A2(n1006), .Y(n1007) );
  NAND4X0_HVT U1245 ( .A1(n1009), .A2(n1008), .A3(n1294), .A4(n1007), .Y(n1011) );
  AO222X1_HVT U1246 ( .A1(n1011), .A2(n1557), .A3(n233), .A4(sram_raddr_b5[4]), 
        .A5(n224), .A6(n1010), .Y(n_sram_raddr_b5[4]) );
  NAND2X0_HVT U1247 ( .A1(n1012), .A2(n318), .Y(n1034) );
  AO221X1_HVT U1248 ( .A1(n1034), .A2(n1012), .A3(n1034), .A4(n318), .A5(n219), 
        .Y(n1302) );
  NAND3X0_HVT U1249 ( .A1(n266), .A2(n324), .A3(n1288), .Y(n1025) );
  AO221X1_HVT U1250 ( .A1(sram_raddr_b2[6]), .A2(n1034), .A3(n390), .A4(n1017), 
        .A5(n220), .Y(n1307) );
  NAND2X0_HVT U1251 ( .A1(n1019), .A2(n1018), .Y(n1030) );
  NAND2X0_HVT U1252 ( .A1(sram_raddr_b5[6]), .A2(n1025), .Y(n1050) );
  NAND2X0_HVT U1253 ( .A1(n1318), .A2(n1050), .Y(n1028) );
  AO222X1_HVT U1254 ( .A1(n404), .A2(n1028), .A3(n404), .A4(n1026), .A5(n1028), 
        .A6(n215), .Y(n1029) );
  NAND4X0_HVT U1255 ( .A1(n1031), .A2(n1307), .A3(n1030), .A4(n1029), .Y(n1033) );
  NAND3X0_HVT U1256 ( .A1(sram_raddr_b5[6]), .A2(sram_raddr_b5[5]), .A3(n1290), 
        .Y(n1041) );
  AO21X1_HVT U1257 ( .A1(n223), .A2(n1041), .A3(n234), .Y(n1042) );
  OA222X1_HVT U1258 ( .A1(sram_raddr_b5[6]), .A2(n224), .A3(sram_raddr_b5[6]), 
        .A4(sram_raddr_b5[5]), .A5(sram_raddr_b5[6]), .A6(n1290), .Y(n1032) );
  AO22X1_HVT U1259 ( .A1(n206), .A2(n1033), .A3(n1042), .A4(n1032), .Y(
        n_sram_raddr_b5[6]) );
  NAND2X0_HVT U1260 ( .A1(sram_raddr_b2[6]), .A2(n1034), .Y(n1035) );
  NAND2X0_HVT U1261 ( .A1(n260), .A2(n1035), .Y(n1045) );
  AO221X1_HVT U1262 ( .A1(n1045), .A2(n1035), .A3(n1045), .A4(n260), .A5(n220), 
        .Y(n1312) );
  OA21X1_HVT U1263 ( .A1(n1071), .A2(n1036), .A3(n1312), .Y(n1040) );
  NAND3X0_HVT U1264 ( .A1(n1318), .A2(n354), .A3(n1050), .Y(n1039) );
  AO221X1_HVT U1265 ( .A1(n216), .A2(col[1]), .A3(n214), .A4(n1050), .A5(n354), 
        .Y(n1037) );
  NAND4X0_HVT U1266 ( .A1(n1040), .A2(n1039), .A3(n1038), .A4(n1037), .Y(n1044) );
  OA222X1_HVT U1267 ( .A1(sram_raddr_b5[7]), .A2(n223), .A3(sram_raddr_b5[7]), 
        .A4(n1056), .A5(n1042), .A6(n354), .Y(n1043) );
  AO21X1_HVT U1268 ( .A1(n203), .A2(n1044), .A3(n1043), .Y(n_sram_raddr_b5[7])
         );
  OR2X1_HVT U1269 ( .A1(n1045), .A2(sram_raddr_b2[8]), .Y(n1065) );
  NAND2X0_HVT U1270 ( .A1(sram_raddr_b2[8]), .A2(n1045), .Y(n1047) );
  OA221X1_HVT U1271 ( .A1(n220), .A2(n1065), .A3(n220), .A4(n1047), .A5(n1046), 
        .Y(n1325) );
  AND3X1_HVT U1272 ( .A1(n214), .A2(n354), .A3(n1050), .Y(n1060) );
  NAND2X0_HVT U1273 ( .A1(sram_raddr_b5[8]), .A2(n1332), .Y(n1049) );
  OA22X1_HVT U1274 ( .A1(n1060), .A2(n1049), .A3(n1048), .A4(n1071), .Y(n1054)
         );
  NAND4X0_HVT U1275 ( .A1(n1318), .A2(n281), .A3(n354), .A4(n1050), .Y(n1068)
         );
  NAND3X0_HVT U1276 ( .A1(n1325), .A2(n1054), .A3(n1068), .Y(n1059) );
  NAND4X0_HVT U1277 ( .A1(sram_raddr_b5[8]), .A2(sram_raddr_b5[7]), .A3(n1056), 
        .A4(n1303), .Y(n1055) );
  NAND2X0_HVT U1278 ( .A1(n168), .A2(n1055), .Y(n1073) );
  AND3X1_HVT U1279 ( .A1(n223), .A2(sram_raddr_b5[7]), .A3(n1056), .Y(n1075)
         );
  OR2X1_HVT U1280 ( .A1(sram_raddr_b5[8]), .A2(n1075), .Y(n1057) );
  AO22X1_HVT U1281 ( .A1(n204), .A2(n1059), .A3(n1058), .A4(n1057), .Y(
        n_sram_raddr_b5[8]) );
  AO22X1_HVT U1282 ( .A1(col[1]), .A2(n213), .A3(n1060), .A4(n281), .Y(n1067)
         );
  OA221X1_HVT U1283 ( .A1(sram_raddr_b5[9]), .A2(n1068), .A3(n394), .A4(n1067), 
        .A5(n1331), .Y(n1072) );
  OA22X1_HVT U1284 ( .A1(n1074), .A2(n221), .A3(n394), .A4(n1073), .Y(n1077)
         );
  NAND3X0_HVT U1285 ( .A1(sram_raddr_b5[8]), .A2(n1075), .A3(n394), .Y(n1076)
         );
  NAND2X0_HVT U1286 ( .A1(n1077), .A2(n1076), .Y(n_sram_raddr_b5[9]) );
  AO22X1_HVT U1287 ( .A1(n1260), .A2(n250), .A3(n1320), .A4(n285), .Y(n1079)
         );
  AO221X1_HVT U1288 ( .A1(sram_raddr_b6[0]), .A2(n1084), .A3(n418), .A4(n1162), 
        .A5(n1079), .Y(n1080) );
  AO22X1_HVT U1289 ( .A1(n203), .A2(n1080), .A3(sram_raddr_b6[0]), .A4(n168), 
        .Y(n_sram_raddr_b6[0]) );
  AO22X1_HVT U1290 ( .A1(n204), .A2(n1085), .A3(sram_raddr_b6[1]), .A4(n217), 
        .Y(n_sram_raddr_b6[1]) );
  AO22X1_HVT U1291 ( .A1(sram_raddr_b6[2]), .A2(n216), .A3(n242), .A4(n1125), 
        .Y(n1088) );
  AO221X1_HVT U1292 ( .A1(sram_raddr_b3[2]), .A2(n1109), .A3(n326), .A4(n1107), 
        .A5(n173), .Y(n1087) );
  NAND3X0_HVT U1293 ( .A1(n1088), .A2(n1087), .A3(n1086), .Y(n1091) );
  OA221X1_HVT U1294 ( .A1(n1091), .A2(n1162), .A3(n1091), .A4(n1090), .A5(n203), .Y(n1092) );
  AO221X1_HVT U1295 ( .A1(sram_raddr_b6[2]), .A2(n233), .A3(n242), .A4(n224), 
        .A5(n1092), .Y(n_sram_raddr_b6[2]) );
  NAND2X0_HVT U1296 ( .A1(n225), .A2(n242), .Y(n1093) );
  NAND2X0_HVT U1297 ( .A1(n1303), .A2(n1093), .Y(n1104) );
  NAND2X0_HVT U1298 ( .A1(n242), .A2(n1148), .Y(n1094) );
  NAND2X0_HVT U1299 ( .A1(n213), .A2(n1094), .Y(n1096) );
  AOI22X1_HVT U1300 ( .A1(sram_raddr_b6[3]), .A2(n1096), .A3(n1095), .A4(n1162), .Y(n1101) );
  NAND3X0_HVT U1301 ( .A1(sram_raddr_b6[2]), .A2(n351), .A3(n1148), .Y(n1099)
         );
  OA222X1_HVT U1302 ( .A1(sram_raddr_b3[3]), .A2(sram_raddr_b3[2]), .A3(
        sram_raddr_b3[3]), .A4(n1109), .A5(n1107), .A6(n1106), .Y(n1097) );
  NAND2X0_HVT U1303 ( .A1(n1320), .A2(n1097), .Y(n1098) );
  NAND4X0_HVT U1304 ( .A1(n1101), .A2(n1100), .A3(n1099), .A4(n1098), .Y(n1103) );
  AND2X1_HVT U1305 ( .A1(sram_raddr_b6[2]), .A2(n351), .Y(n1102) );
  AO222X1_HVT U1306 ( .A1(n1104), .A2(sram_raddr_b6[3]), .A3(n1103), .A4(n204), 
        .A5(n1102), .A6(n223), .Y(n_sram_raddr_b6[3]) );
  AND3X1_HVT U1307 ( .A1(sram_raddr_b6[3]), .A2(sram_raddr_b6[2]), .A3(
        sram_raddr_b6[4]), .Y(n1123) );
  OA21X1_HVT U1308 ( .A1(n242), .A2(n351), .A3(n276), .Y(n1124) );
  NOR2X0_HVT U1309 ( .A1(n1123), .A2(n1124), .Y(n1114) );
  OA22X1_HVT U1310 ( .A1(n1125), .A2(n1114), .A3(n216), .A4(n276), .Y(n1113)
         );
  NAND2X0_HVT U1311 ( .A1(n1162), .A2(n1105), .Y(n1111) );
  OA21X1_HVT U1312 ( .A1(n1107), .A2(n1106), .A3(n320), .Y(n1116) );
  OAI221X1_HVT U1313 ( .A1(n1116), .A2(n1109), .A3(n1116), .A4(n1108), .A5(
        n178), .Y(n1110) );
  NAND4X0_HVT U1314 ( .A1(n1113), .A2(n1112), .A3(n1111), .A4(n1110), .Y(n1115) );
  AO222X1_HVT U1315 ( .A1(n1115), .A2(n206), .A3(n234), .A4(sram_raddr_b6[4]), 
        .A5(n223), .A6(n1114), .Y(n_sram_raddr_b6[4]) );
  NAND3X0_HVT U1316 ( .A1(n1124), .A2(n339), .A3(n1148), .Y(n1120) );
  AO221X1_HVT U1317 ( .A1(n216), .A2(n1125), .A3(n216), .A4(n1124), .A5(n339), 
        .Y(n1118) );
  NAND2X0_HVT U1318 ( .A1(n1116), .A2(n261), .Y(n1137) );
  AO221X1_HVT U1319 ( .A1(n1137), .A2(n1116), .A3(n1137), .A4(n261), .A5(n226), 
        .Y(n1117) );
  NAND4X0_HVT U1320 ( .A1(n1120), .A2(n1119), .A3(n1118), .A4(n1117), .Y(n1122) );
  NAND4X0_HVT U1321 ( .A1(sram_raddr_b6[3]), .A2(sram_raddr_b6[2]), .A3(
        sram_raddr_b6[5]), .A4(sram_raddr_b6[4]), .Y(n1134) );
  NAND2X0_HVT U1322 ( .A1(n1124), .A2(n339), .Y(n1136) );
  AO221X1_HVT U1323 ( .A1(n215), .A2(n1125), .A3(n215), .A4(n1136), .A5(n427), 
        .Y(n1129) );
  AO221X1_HVT U1324 ( .A1(sram_raddr_b3[6]), .A2(n1137), .A3(n400), .A4(n1126), 
        .A5(n227), .Y(n1128) );
  NAND3X0_HVT U1325 ( .A1(n427), .A2(n1148), .A3(n1136), .Y(n1127) );
  NAND4X0_HVT U1326 ( .A1(n1130), .A2(n1129), .A3(n1128), .A4(n1127), .Y(n1133) );
  NAND2X0_HVT U1327 ( .A1(sram_raddr_b6[6]), .A2(n1135), .Y(n1145) );
  NAND2X0_HVT U1328 ( .A1(sram_raddr_b6[6]), .A2(n1136), .Y(n1151) );
  NAND3X0_HVT U1329 ( .A1(n270), .A2(n1148), .A3(n1151), .Y(n1142) );
  NAND2X0_HVT U1330 ( .A1(sram_raddr_b3[6]), .A2(n1137), .Y(n1138) );
  NAND2X0_HVT U1331 ( .A1(n350), .A2(n1138), .Y(n1149) );
  AO221X1_HVT U1332 ( .A1(n1149), .A2(n1138), .A3(n1149), .A4(n350), .A5(n173), 
        .Y(n1140) );
  AO221X1_HVT U1333 ( .A1(n216), .A2(n1387), .A3(n216), .A4(n1151), .A5(n270), 
        .Y(n1139) );
  NAND4X0_HVT U1334 ( .A1(n1142), .A2(n1141), .A3(n1140), .A4(n1139), .Y(n1144) );
  NAND2X0_HVT U1335 ( .A1(sram_raddr_b6[7]), .A2(n1147), .Y(n1146) );
  AO221X1_HVT U1336 ( .A1(n188), .A2(n388), .A3(n223), .A4(n1146), .A5(n234), 
        .Y(n1170) );
  AND3X1_HVT U1337 ( .A1(n223), .A2(sram_raddr_b6[7]), .A3(n1147), .Y(n1171)
         );
  NAND4X0_HVT U1338 ( .A1(n388), .A2(n270), .A3(n1148), .A4(n1151), .Y(n1160)
         );
  NAND2X0_HVT U1339 ( .A1(n1150), .A2(n268), .Y(n1164) );
  AO221X1_HVT U1340 ( .A1(n1164), .A2(n1150), .A3(n1164), .A4(n268), .A5(n173), 
        .Y(n1153) );
  AND3X1_HVT U1341 ( .A1(n215), .A2(n270), .A3(n1151), .Y(n1159) );
  OR3X1_HVT U1342 ( .A1(n1158), .A2(n1159), .A3(n388), .Y(n1152) );
  NAND4X0_HVT U1343 ( .A1(n1160), .A2(n1154), .A3(n1153), .A4(n1152), .Y(n1156) );
  OA221X1_HVT U1344 ( .A1(n1156), .A2(n1155), .A3(n1156), .A4(n1162), .A5(
        n1557), .Y(n1157) );
  AO221X1_HVT U1345 ( .A1(n1170), .A2(sram_raddr_b6[8]), .A3(n1170), .A4(n1171), .A5(n1157), .Y(n_sram_raddr_b6[8]) );
  AO21X1_HVT U1346 ( .A1(n1159), .A2(n388), .A3(n1158), .Y(n1161) );
  AO22X1_HVT U1347 ( .A1(sram_raddr_b6[9]), .A2(n1161), .A3(n406), .A4(n1160), 
        .Y(n1169) );
  NAND2X0_HVT U1348 ( .A1(n1163), .A2(n1162), .Y(n1167) );
  AO221X1_HVT U1349 ( .A1(sram_raddr_b3[9]), .A2(n1165), .A3(n402), .A4(n1164), 
        .A5(n227), .Y(n1166) );
  NAND4X0_HVT U1350 ( .A1(n1169), .A2(n1168), .A3(n1167), .A4(n1166), .Y(n1173) );
  OA222X1_HVT U1351 ( .A1(sram_raddr_b6[9]), .A2(sram_raddr_b6[8]), .A3(
        sram_raddr_b6[9]), .A4(n1171), .A5(n406), .A6(n1170), .Y(n1172) );
  AO21X1_HVT U1352 ( .A1(n206), .A2(n1173), .A3(n1172), .Y(n_sram_raddr_b6[9])
         );
  AO22X1_HVT U1353 ( .A1(n1260), .A2(n251), .A3(n178), .A4(n286), .Y(n1175) );
  AO221X1_HVT U1354 ( .A1(sram_raddr_b7[0]), .A2(n1236), .A3(n419), .A4(n1248), 
        .A5(n1175), .Y(n1176) );
  AO22X1_HVT U1355 ( .A1(n205), .A2(n1176), .A3(sram_raddr_b7[0]), .A4(n168), 
        .Y(n_sram_raddr_b7[0]) );
  AO22X1_HVT U1356 ( .A1(n205), .A2(n1180), .A3(sram_raddr_b7[1]), .A4(n217), 
        .Y(n_sram_raddr_b7[1]) );
  NAND2X0_HVT U1357 ( .A1(n1226), .A2(n243), .Y(n1187) );
  OA21X1_HVT U1358 ( .A1(n214), .A2(n243), .A3(n1187), .Y(n1182) );
  AO221X1_HVT U1359 ( .A1(sram_raddr_b4[2]), .A2(n1203), .A3(n322), .A4(n1201), 
        .A5(n173), .Y(n1181) );
  NAND3X0_HVT U1360 ( .A1(n1183), .A2(n1182), .A3(n1181), .Y(n1185) );
  OA221X1_HVT U1361 ( .A1(n1185), .A2(n1248), .A3(n1185), .A4(n1184), .A5(n204), .Y(n1186) );
  AO221X1_HVT U1362 ( .A1(sram_raddr_b7[2]), .A2(n234), .A3(n243), .A4(n225), 
        .A5(n1186), .Y(n_sram_raddr_b7[2]) );
  NAND2X0_HVT U1363 ( .A1(n216), .A2(n1187), .Y(n1188) );
  OA222X1_HVT U1364 ( .A1(sram_raddr_b7[3]), .A2(n1226), .A3(sram_raddr_b7[3]), 
        .A4(sram_raddr_b7[2]), .A5(n347), .A6(n1188), .Y(n1192) );
  OA222X1_HVT U1365 ( .A1(sram_raddr_b4[3]), .A2(sram_raddr_b4[2]), .A3(
        sram_raddr_b4[3]), .A4(n1203), .A5(n1201), .A6(n1200), .Y(n1190) );
  AO22X1_HVT U1366 ( .A1(n178), .A2(n1190), .A3(n1189), .A4(n1248), .Y(n1191)
         );
  OR3X1_HVT U1367 ( .A1(n1193), .A2(n1192), .A3(n1191), .Y(n1197) );
  NAND2X0_HVT U1368 ( .A1(n223), .A2(n243), .Y(n1194) );
  NAND2X0_HVT U1369 ( .A1(n1303), .A2(n1194), .Y(n1196) );
  AND2X1_HVT U1370 ( .A1(sram_raddr_b7[2]), .A2(n347), .Y(n1195) );
  AO222X1_HVT U1371 ( .A1(n1197), .A2(n206), .A3(n1196), .A4(sram_raddr_b7[3]), 
        .A5(n1195), .A6(n223), .Y(n_sram_raddr_b7[3]) );
  AND3X1_HVT U1372 ( .A1(sram_raddr_b7[3]), .A2(sram_raddr_b7[2]), .A3(
        sram_raddr_b7[4]), .Y(n1213) );
  OA21X1_HVT U1373 ( .A1(n243), .A2(n347), .A3(n277), .Y(n1215) );
  NOR2X0_HVT U1374 ( .A1(n1213), .A2(n1215), .Y(n1208) );
  OA22X1_HVT U1375 ( .A1(n215), .A2(n277), .A3(n1208), .A4(n1198), .Y(n1207)
         );
  NAND2X0_HVT U1376 ( .A1(n1248), .A2(n1199), .Y(n1205) );
  OA21X1_HVT U1377 ( .A1(n1201), .A2(n1200), .A3(n336), .Y(n1210) );
  OAI221X1_HVT U1378 ( .A1(n1210), .A2(n1203), .A3(n1210), .A4(n1202), .A5(
        n178), .Y(n1204) );
  NAND4X0_HVT U1379 ( .A1(n1207), .A2(n1206), .A3(n1205), .A4(n1204), .Y(n1209) );
  AO222X1_HVT U1380 ( .A1(n1209), .A2(n1557), .A3(n234), .A4(sram_raddr_b7[4]), 
        .A5(n225), .A6(n1208), .Y(n_sram_raddr_b7[4]) );
  NAND2X0_HVT U1381 ( .A1(n1210), .A2(n271), .Y(n1214) );
  NAND4X0_HVT U1382 ( .A1(sram_raddr_b7[3]), .A2(sram_raddr_b7[2]), .A3(
        sram_raddr_b7[5]), .A4(sram_raddr_b7[4]), .Y(n1219) );
  NAND2X0_HVT U1383 ( .A1(sram_raddr_b4[6]), .A2(n1214), .Y(n1227) );
  NAND2X0_HVT U1384 ( .A1(n1215), .A2(n340), .Y(n1225) );
  HADDX1_HVT U1385 ( .A0(sram_raddr_b7[6]), .B0(n1225), .SO(n1216) );
  NAND2X0_HVT U1386 ( .A1(sram_raddr_b7[6]), .A2(n1220), .Y(n1230) );
  OA21X1_HVT U1387 ( .A1(sram_raddr_b7[6]), .A2(n1220), .A3(n1230), .Y(n1221)
         );
  AO22X1_HVT U1388 ( .A1(n188), .A2(n1221), .A3(n232), .A4(sram_raddr_b7[6]), 
        .Y(n1222) );
  AO221X1_HVT U1389 ( .A1(n205), .A2(n1224), .A3(n206), .A4(n1223), .A5(n1222), 
        .Y(n_sram_raddr_b7[6]) );
  NAND2X0_HVT U1390 ( .A1(sram_raddr_b7[6]), .A2(n1225), .Y(n1244) );
  NAND3X0_HVT U1391 ( .A1(n1226), .A2(n330), .A3(n1244), .Y(n1235) );
  NAND2X0_HVT U1392 ( .A1(n316), .A2(n1227), .Y(n1233) );
  NAND2X0_HVT U1393 ( .A1(sram_raddr_b7[7]), .A2(n1232), .Y(n1231) );
  AO221X1_HVT U1394 ( .A1(n224), .A2(n353), .A3(n224), .A4(n1231), .A5(n234), 
        .Y(n1254) );
  AND3X1_HVT U1395 ( .A1(n224), .A2(sram_raddr_b7[7]), .A3(n1232), .Y(n1255)
         );
  OR2X1_HVT U1396 ( .A1(n1235), .A2(sram_raddr_b7[8]), .Y(n1246) );
  NAND2X0_HVT U1397 ( .A1(n1234), .A2(n328), .Y(n1247) );
  AO221X1_HVT U1398 ( .A1(n1247), .A2(n1234), .A3(n1247), .A4(n328), .A5(n173), 
        .Y(n1238) );
  NAND3X0_HVT U1399 ( .A1(n1236), .A2(n1235), .A3(sram_raddr_b7[8]), .Y(n1237)
         );
  NAND4X0_HVT U1400 ( .A1(n1246), .A2(n1239), .A3(n1238), .A4(n1237), .Y(n1241) );
  OA221X1_HVT U1401 ( .A1(n1241), .A2(n1248), .A3(n1241), .A4(n1240), .A5(n203), .Y(n1242) );
  AO221X1_HVT U1402 ( .A1(n1254), .A2(sram_raddr_b7[8]), .A3(n1254), .A4(n1255), .A5(n1242), .Y(n_sram_raddr_b7[8]) );
  NAND2X0_HVT U1403 ( .A1(n330), .A2(n1244), .Y(n1245) );
  AO221X1_HVT U1404 ( .A1(n262), .A2(sram_raddr_b7[8]), .A3(n262), .A4(n1245), 
        .A5(n1306), .Y(n1253) );
  HADDX1_HVT U1405 ( .A0(n395), .B0(n1247), .SO(n1250) );
  AO22X1_HVT U1406 ( .A1(n178), .A2(n1250), .A3(n1249), .A4(n1248), .Y(n1251)
         );
  AO221X1_HVT U1407 ( .A1(sram_raddr_b7[9]), .A2(n1253), .A3(n405), .A4(n1252), 
        .A5(n1251), .Y(n1257) );
  OA222X1_HVT U1408 ( .A1(sram_raddr_b7[9]), .A2(sram_raddr_b7[8]), .A3(
        sram_raddr_b7[9]), .A4(n1255), .A5(n405), .A6(n1254), .Y(n1256) );
  AO221X1_HVT U1409 ( .A1(n1557), .A2(n1258), .A3(n207), .A4(n1257), .A5(n1256), .Y(n_sram_raddr_b7[9]) );
  AO22X1_HVT U1410 ( .A1(n1260), .A2(n287), .A3(n178), .A4(n252), .Y(n1261) );
  AO221X1_HVT U1411 ( .A1(sram_raddr_b8[0]), .A2(n1332), .A3(n420), .A4(n1336), 
        .A5(n1261), .Y(n1262) );
  AO22X1_HVT U1412 ( .A1(n203), .A2(n1262), .A3(sram_raddr_b8[0]), .A4(n168), 
        .Y(n_sram_raddr_b8[0]) );
  AO22X1_HVT U1413 ( .A1(n207), .A2(n1267), .A3(sram_raddr_b8[1]), .A4(n217), 
        .Y(n_sram_raddr_b8[1]) );
  AO22X1_HVT U1414 ( .A1(sram_raddr_b8[2]), .A2(n216), .A3(n245), .A4(n1299), 
        .Y(n1270) );
  AO221X1_HVT U1415 ( .A1(sram_raddr_b5[2]), .A2(n1291), .A3(n321), .A4(n1289), 
        .A5(n227), .Y(n1268) );
  NAND3X0_HVT U1416 ( .A1(n1270), .A2(n1269), .A3(n1268), .Y(n1272) );
  OA221X1_HVT U1417 ( .A1(n1272), .A2(n1336), .A3(n1272), .A4(n1271), .A5(
        n1557), .Y(n1273) );
  AO221X1_HVT U1418 ( .A1(sram_raddr_b8[2]), .A2(n234), .A3(n245), .A4(n225), 
        .A5(n1273), .Y(n_sram_raddr_b8[2]) );
  OA222X1_HVT U1419 ( .A1(sram_raddr_b5[3]), .A2(sram_raddr_b5[2]), .A3(
        sram_raddr_b5[3]), .A4(n1291), .A5(n1289), .A6(n1288), .Y(n1277) );
  OA21X1_HVT U1420 ( .A1(sram_raddr_b8[3]), .A2(n1275), .A3(n1274), .Y(n1276)
         );
  AOI22X1_HVT U1421 ( .A1(n178), .A2(n1277), .A3(n1276), .A4(n1336), .Y(n1281)
         );
  AO221X1_HVT U1422 ( .A1(n216), .A2(sram_raddr_b8[2]), .A3(n216), .A4(n1299), 
        .A5(n282), .Y(n1279) );
  NAND3X0_HVT U1423 ( .A1(sram_raddr_b8[2]), .A2(n1318), .A3(n282), .Y(n1278)
         );
  NAND4X0_HVT U1424 ( .A1(n1281), .A2(n1280), .A3(n1279), .A4(n1278), .Y(n1285) );
  NAND2X0_HVT U1425 ( .A1(n223), .A2(n245), .Y(n1282) );
  NAND2X0_HVT U1426 ( .A1(n1303), .A2(n1282), .Y(n1284) );
  AND2X1_HVT U1427 ( .A1(sram_raddr_b8[2]), .A2(n282), .Y(n1283) );
  AO222X1_HVT U1428 ( .A1(n1285), .A2(n206), .A3(n1284), .A4(sram_raddr_b8[3]), 
        .A5(n1283), .A6(n179), .Y(n_sram_raddr_b8[3]) );
  NAND3X0_HVT U1429 ( .A1(sram_raddr_b8[4]), .A2(sram_raddr_b8[3]), .A3(
        sram_raddr_b8[2]), .Y(n1304) );
  OA21X1_HVT U1430 ( .A1(n282), .A2(n245), .A3(n346), .Y(n1298) );
  AND2X1_HVT U1431 ( .A1(n1304), .A2(n1286), .Y(n1296) );
  OA22X1_HVT U1432 ( .A1(n215), .A2(n346), .A3(n1296), .A4(n1299), .Y(n1295)
         );
  NAND2X0_HVT U1433 ( .A1(n1336), .A2(n1287), .Y(n1293) );
  OA21X1_HVT U1434 ( .A1(n1289), .A2(n1288), .A3(n324), .Y(n1301) );
  OAI221X1_HVT U1435 ( .A1(n1301), .A2(n1291), .A3(n1301), .A4(n1290), .A5(
        n178), .Y(n1292) );
  NAND4X0_HVT U1436 ( .A1(n1295), .A2(n1294), .A3(n1293), .A4(n1292), .Y(n1297) );
  AO222X1_HVT U1437 ( .A1(n1297), .A2(n204), .A3(n232), .A4(sram_raddr_b8[4]), 
        .A5(n179), .A6(n1296), .Y(n_sram_raddr_b8[4]) );
  NAND2X0_HVT U1438 ( .A1(n1298), .A2(n325), .Y(n1305) );
  NAND2X0_HVT U1439 ( .A1(n1301), .A2(n266), .Y(n1310) );
  AND4X1_HVT U1440 ( .A1(sram_raddr_b8[5]), .A2(sram_raddr_b8[4]), .A3(
        sram_raddr_b8[3]), .A4(sram_raddr_b8[2]), .Y(n1309) );
  NAND2X0_HVT U1441 ( .A1(sram_raddr_b8[6]), .A2(n1305), .Y(n1322) );
  NAND2X0_HVT U1442 ( .A1(sram_raddr_b8[6]), .A2(n1309), .Y(n1314) );
  NAND2X0_HVT U1443 ( .A1(sram_raddr_b5[6]), .A2(n1310), .Y(n1311) );
  NAND2X0_HVT U1444 ( .A1(n354), .A2(n1311), .Y(n1319) );
  NAND2X0_HVT U1445 ( .A1(sram_raddr_b8[7]), .A2(n1317), .Y(n1316) );
  AO221X1_HVT U1446 ( .A1(n188), .A2(n337), .A3(n188), .A4(n1316), .A5(n232), 
        .Y(n1342) );
  AND3X1_HVT U1447 ( .A1(n188), .A2(sram_raddr_b8[7]), .A3(n1317), .Y(n1343)
         );
  NAND4X0_HVT U1448 ( .A1(n1318), .A2(n337), .A3(n269), .A4(n1322), .Y(n1334)
         );
  NAND2X0_HVT U1449 ( .A1(n1321), .A2(n281), .Y(n1335) );
  AO221X1_HVT U1450 ( .A1(n1335), .A2(n1321), .A3(n1335), .A4(n281), .A5(n227), 
        .Y(n1324) );
  NAND3X0_HVT U1451 ( .A1(n215), .A2(n269), .A3(n1322), .Y(n1333) );
  NAND3X0_HVT U1452 ( .A1(sram_raddr_b8[8]), .A2(n1332), .A3(n1333), .Y(n1323)
         );
  NAND4X0_HVT U1453 ( .A1(n1325), .A2(n1334), .A3(n1324), .A4(n1323), .Y(n1329) );
  OA221X1_HVT U1454 ( .A1(n1329), .A2(n1328), .A3(n1329), .A4(n1327), .A5(
        n1557), .Y(n1330) );
  AO221X1_HVT U1455 ( .A1(n1342), .A2(sram_raddr_b8[8]), .A3(n1342), .A4(n1343), .A5(n1330), .Y(n_sram_raddr_b8[8]) );
  OA21X1_HVT U1456 ( .A1(sram_raddr_b8[8]), .A2(n1333), .A3(n1332), .Y(n1341)
         );
  HADDX1_HVT U1457 ( .A0(n394), .B0(n1335), .SO(n1338) );
  AO22X1_HVT U1458 ( .A1(n178), .A2(n1338), .A3(n1337), .A4(n1336), .Y(n1339)
         );
  AO221X1_HVT U1459 ( .A1(sram_raddr_b8[9]), .A2(n1341), .A3(n407), .A4(n1340), 
        .A5(n1339), .Y(n1345) );
  OA222X1_HVT U1460 ( .A1(sram_raddr_b8[9]), .A2(sram_raddr_b8[8]), .A3(
        sram_raddr_b8[9]), .A4(n1343), .A5(n407), .A6(n1342), .Y(n1344) );
  AO221X1_HVT U1461 ( .A1(n204), .A2(n1346), .A3(n206), .A4(n1345), .A5(n1344), 
        .Y(n_sram_raddr_b8[9]) );
  OA221X1_HVT U1462 ( .A1(n1063), .A2(write_col_conv1[1]), .A3(n257), .A4(n312), .A5(n1062), .Y(n1350) );
  NAND2X0_HVT U1463 ( .A1(n1350), .A2(n1347), .Y(n_sram_write_enable_b0) );
  OA221X1_HVT U1464 ( .A1(write_col_conv1[1]), .A2(n258), .A3(n312), .A4(n1062), .A5(n1063), .Y(n1351) );
  NAND2X0_HVT U1465 ( .A1(n1351), .A2(n1347), .Y(n_sram_write_enable_b1) );
  NAND3X0_HVT U1466 ( .A1(write_col_conv1[1]), .A2(n1063), .A3(n258), .Y(n1471) );
  NAND3X0_HVT U1467 ( .A1(n1062), .A2(n257), .A3(n312), .Y(n1475) );
  NAND2X0_HVT U1468 ( .A1(n1471), .A2(n1475), .Y(n1468) );
  NAND2X0_HVT U1469 ( .A1(n1347), .A2(n1468), .Y(n_sram_write_enable_b2) );
  AO222X1_HVT U1470 ( .A1(write_row_conv1[3]), .A2(n1061), .A3(
        write_row_conv1[3]), .A4(write_row_conv1[2]), .A5(n249), .A6(n357), 
        .Y(n1348) );
  AND3X1_HVT U1471 ( .A1(n1348), .A2(n1469), .A3(n289), .Y(n1349) );
  NAND2X0_HVT U1472 ( .A1(n1350), .A2(n1349), .Y(n_sram_write_enable_b3) );
  NAND2X0_HVT U1473 ( .A1(n1351), .A2(n1349), .Y(n_sram_write_enable_b4) );
  NAND2X0_HVT U1474 ( .A1(n1349), .A2(n1468), .Y(n_sram_write_enable_b5) );
  OA222X1_HVT U1475 ( .A1(n1061), .A2(write_row_conv1[3]), .A3(n249), .A4(
        write_row_conv1[2]), .A5(n357), .A6(n289), .Y(n1472) );
  NAND4X0_HVT U1476 ( .A1(n1472), .A2(n1363), .A3(delay2_write_enable), .A4(
        n1350), .Y(n_sram_write_enable_b6) );
  NAND4X0_HVT U1477 ( .A1(n1472), .A2(n1363), .A3(delay2_write_enable), .A4(
        n1351), .Y(n_sram_write_enable_b7) );
  NAND4X0_HVT U1478 ( .A1(n1472), .A2(n1363), .A3(delay2_write_enable), .A4(
        n1468), .Y(n_sram_write_enable_b8) );
  AND3X1_HVT U1479 ( .A1(n1354), .A2(delay3_write_enable), .A3(n469), .Y(n1353) );
  NAND4X0_HVT U1480 ( .A1(n1353), .A2(n1512), .A3(n311), .A4(n255), .Y(
        n_sram_write_enable_c0) );
  AND3X1_HVT U1481 ( .A1(delay3_addr_change[2]), .A2(n1353), .A3(n311), .Y(
        n1352) );
  NAND2X0_HVT U1482 ( .A1(n1352), .A2(n1512), .Y(n_sram_write_enable_c1) );
  NAND4X0_HVT U1483 ( .A1(delay3_addr_change[3]), .A2(n1353), .A3(n1512), .A4(
        n255), .Y(n_sram_write_enable_c2) );
  NAND4X0_HVT U1484 ( .A1(delay3_addr_change[3]), .A2(delay3_addr_change[2]), 
        .A3(n1353), .A4(n1512), .Y(n_sram_write_enable_c3) );
  AND3X1_HVT U1485 ( .A1(delay3_addr_change[4]), .A2(n311), .A3(n255), .Y(
        n1508) );
  NAND4X0_HVT U1486 ( .A1(n1354), .A2(delay3_write_enable), .A3(n1508), .A4(
        n1512), .Y(n_sram_write_enable_c4) );
  NAND4X0_HVT U1487 ( .A1(mem_sel), .A2(n1353), .A3(n255), .A4(n311), .Y(
        n_sram_write_enable_d0) );
  NAND2X0_HVT U1488 ( .A1(mem_sel), .A2(n1352), .Y(n_sram_write_enable_d1) );
  NAND4X0_HVT U1489 ( .A1(delay3_addr_change[3]), .A2(mem_sel), .A3(n1353), 
        .A4(n255), .Y(n_sram_write_enable_d2) );
  NAND4X0_HVT U1490 ( .A1(mem_sel), .A2(delay3_addr_change[3]), .A3(
        delay3_addr_change[2]), .A4(n1353), .Y(n_sram_write_enable_d3) );
  NAND4X0_HVT U1491 ( .A1(mem_sel), .A2(n1354), .A3(delay3_write_enable), .A4(
        n1508), .Y(n_sram_write_enable_d4) );
  NAND4X0_HVT U1492 ( .A1(state[0]), .A2(n1023), .A3(n1024), .A4(n240), .Y(
        n1563) );
  NAND3X0_HVT U1493 ( .A1(n1023), .A2(n1445), .A3(state[2]), .Y(n1356) );
  NAND3X0_HVT U1494 ( .A1(state[1]), .A2(n1024), .A3(state[3]), .Y(n1446) );
  NAND2X0_HVT U1495 ( .A1(n1549), .A2(conv_done), .Y(n1365) );
  NAND3X0_HVT U1496 ( .A1(n1023), .A2(n1024), .A3(n253), .Y(n1358) );
  OA22X1_HVT U1497 ( .A1(conv_done), .A2(n1361), .A3(n1358), .A4(n1357), .Y(
        n1360) );
  NAND2X0_HVT U1498 ( .A1(n1445), .A2(state[2]), .Y(n1416) );
  NAND2X0_HVT U1499 ( .A1(n2003), .A2(n462), .Y(n1359) );
  NAND4X0_HVT U1500 ( .A1(n421), .A2(n1360), .A3(n1416), .A4(n1359), .Y(
        n_state[1]) );
  NAND4X0_HVT U1501 ( .A1(state[0]), .A2(n1023), .A3(n240), .A4(state[2]), .Y(
        n1562) );
  OA21X1_HVT U1502 ( .A1(n1023), .A2(n1416), .A3(n1562), .Y(n1464) );
  OA22X1_HVT U1503 ( .A1(conv_done), .A2(n1361), .A3(n1389), .A4(n462), .Y(
        n1362) );
  NAND4X0_HVT U1504 ( .A1(state[1]), .A2(state[0]), .A3(n1024), .A4(state[3]), 
        .Y(n1466) );
  NAND3X0_HVT U1505 ( .A1(n1464), .A2(n1362), .A3(n1466), .Y(n_state[2]) );
  NAND2X0_HVT U1506 ( .A1(n1023), .A2(state[2]), .Y(n1367) );
  NAND3X0_HVT U1507 ( .A1(n1023), .A2(n1445), .A3(n1363), .Y(n1364) );
  NAND4X0_HVT U1508 ( .A1(n1367), .A2(n1366), .A3(n1365), .A4(n1364), .Y(
        n_state[3]) );
  NAND2X0_HVT U1509 ( .A1(n204), .A2(n1390), .Y(n1456) );
  NAND3X0_HVT U1510 ( .A1(n1465), .A2(n1457), .A3(n1368), .Y(n1378) );
  NAND2X0_HVT U1511 ( .A1(n1456), .A2(n1369), .Y(n1382) );
  AO22X1_HVT U1512 ( .A1(weight_cnt[0]), .A2(n1378), .A3(n308), .A4(n1382), 
        .Y(n_weight_cnt[0]) );
  AO22X1_HVT U1513 ( .A1(weight_cnt[1]), .A2(n308), .A3(n444), .A4(
        weight_cnt[0]), .Y(n1370) );
  AO22X1_HVT U1514 ( .A1(n1370), .A2(n1382), .A3(weight_cnt[1]), .A4(n1378), 
        .Y(n_weight_cnt[1]) );
  NAND3X0_HVT U1515 ( .A1(weight_cnt[1]), .A2(weight_cnt[0]), .A3(
        weight_cnt[2]), .Y(n1371) );
  AO21X1_HVT U1516 ( .A1(n1382), .A2(n1371), .A3(n1378), .Y(n1372) );
  OA222X1_HVT U1517 ( .A1(weight_cnt[3]), .A2(n1377), .A3(weight_cnt[3]), .A4(
        n1382), .A5(n439), .A6(n1372), .Y(n_weight_cnt[3]) );
  NAND3X0_HVT U1518 ( .A1(weight_cnt[3]), .A2(n1377), .A3(weight_cnt[4]), .Y(
        n1374) );
  OA221X1_HVT U1519 ( .A1(weight_cnt[4]), .A2(n1377), .A3(weight_cnt[4]), .A4(
        weight_cnt[3]), .A5(n1374), .Y(n1373) );
  AO22X1_HVT U1520 ( .A1(n1373), .A2(n1382), .A3(weight_cnt[4]), .A4(n1378), 
        .Y(n_weight_cnt[4]) );
  AO22X1_HVT U1521 ( .A1(n1375), .A2(n453), .A3(n1374), .A4(weight_cnt[5]), 
        .Y(n1376) );
  AO22X1_HVT U1522 ( .A1(n1376), .A2(n1382), .A3(weight_cnt[5]), .A4(n1378), 
        .Y(n_weight_cnt[5]) );
  AND4X1_HVT U1523 ( .A1(weight_cnt[3]), .A2(n1377), .A3(weight_cnt[4]), .A4(
        weight_cnt[5]), .Y(n1379) );
  NAND2X0_HVT U1524 ( .A1(n1379), .A2(weight_cnt[6]), .Y(n1380) );
  AO21X1_HVT U1525 ( .A1(n1382), .A2(n1380), .A3(n1378), .Y(n1381) );
  OA221X1_HVT U1526 ( .A1(weight_cnt[6]), .A2(n1379), .A3(weight_cnt[6]), .A4(
        n1382), .A5(n1381), .Y(n_weight_cnt[6]) );
  OA222X1_HVT U1527 ( .A1(weight_cnt[7]), .A2(n1383), .A3(weight_cnt[7]), .A4(
        n1382), .A5(n461), .A6(n1381), .Y(n_weight_cnt[7]) );
  OR3X1_HVT U1528 ( .A1(conv2_weight_done), .A2(write_enable), .A3(
        load_data_enable), .Y(n1385) );
  OR3X1_HVT U1529 ( .A1(conv1_weight_done), .A2(write_enable), .A3(
        load_data_enable), .Y(n1384) );
  AO22X1_HVT U1530 ( .A1(n1549), .A2(n1385), .A3(n2003), .A4(n1384), .Y(
        n_write_enable) );
  NAND2X0_HVT U1531 ( .A1(n1549), .A2(n181), .Y(net22462) );
  NAND2X0_HVT U1532 ( .A1(n1565), .A2(col[2]), .Y(n1564) );
  OA221X1_HVT U1533 ( .A1(n1386), .A2(col[3]), .A3(n1564), .A4(n241), .A5(
        n1566), .Y(net22639) );
  AND2X1_HVT U1534 ( .A1(n262), .A2(n1566), .Y(net22654) );
  AO221X1_HVT U1535 ( .A1(sram_raddr_weight[4]), .A2(sram_raddr_weight[3]), 
        .A3(sram_raddr_weight[4]), .A4(sram_raddr_weight[2]), .A5(n1390), .Y(
        n1436) );
  NOR2X0_HVT U1536 ( .A1(n1436), .A2(sram_raddr_weight[5]), .Y(n1439) );
  NAND2X0_HVT U1537 ( .A1(n1439), .A2(n358), .Y(n1433) );
  NAND2X0_HVT U1538 ( .A1(n1428), .A2(n359), .Y(n1429) );
  NAND3X0_HVT U1539 ( .A1(n288), .A2(n355), .A3(n1424), .Y(n1412) );
  OR3X1_HVT U1540 ( .A1(sram_raddr_weight[11]), .A2(sram_raddr_weight[10]), 
        .A3(n1412), .Y(n1405) );
  OR3X1_HVT U1541 ( .A1(sram_raddr_weight[13]), .A2(sram_raddr_weight[12]), 
        .A3(n1405), .Y(n1392) );
  NAND2X0_HVT U1542 ( .A1(n203), .A2(n1392), .Y(n1400) );
  NAND4X0_HVT U1543 ( .A1(sram_raddr_weight[3]), .A2(sram_raddr_weight[2]), 
        .A3(sram_raddr_weight[0]), .A4(sram_raddr_weight[1]), .Y(n1440) );
  NAND2X0_HVT U1544 ( .A1(sram_raddr_weight[4]), .A2(n1444), .Y(n1435) );
  AND3X1_HVT U1545 ( .A1(sram_raddr_weight[5]), .A2(sram_raddr_weight[6]), 
        .A3(n1438), .Y(n1434) );
  AND2X1_HVT U1546 ( .A1(sram_raddr_weight[7]), .A2(n1434), .Y(n1423) );
  NAND2X0_HVT U1547 ( .A1(sram_raddr_weight[8]), .A2(n1423), .Y(n1411) );
  NAND4X0_HVT U1548 ( .A1(sram_raddr_weight[11]), .A2(sram_raddr_weight[9]), 
        .A3(sram_raddr_weight[10]), .A4(n1417), .Y(n1409) );
  AND4X1_HVT U1549 ( .A1(sram_raddr_weight[12]), .A2(sram_raddr_weight[13]), 
        .A3(n1406), .A4(n1455), .Y(n1402) );
  NAND2X0_HVT U1550 ( .A1(sram_raddr_weight[14]), .A2(n1402), .Y(n1398) );
  OR2X1_HVT U1551 ( .A1(n304), .A2(n1398), .Y(n1393) );
  NAND2X0_HVT U1552 ( .A1(n1455), .A2(n1393), .Y(n1391) );
  AO221X1_HVT U1553 ( .A1(n1396), .A2(n304), .A3(n1396), .A4(n221), .A5(n463), 
        .Y(n1395) );
  NOR2X0_HVT U1554 ( .A1(n221), .A2(n1392), .Y(n1404) );
  NAND2X0_HVT U1555 ( .A1(n1404), .A2(n403), .Y(n1397) );
  AO221X1_HVT U1556 ( .A1(n1393), .A2(sram_raddr_weight[15]), .A3(n1393), .A4(
        n1397), .A5(sram_raddr_weight[16]), .Y(n1394) );
  NAND2X0_HVT U1557 ( .A1(n1395), .A2(n1394), .Y(net22692) );
  OAI222X1_HVT U1558 ( .A1(sram_raddr_weight[15]), .A2(n1398), .A3(
        sram_raddr_weight[15]), .A4(n1397), .A5(n304), .A6(n1396), .Y(net22699) );
  NAND3X0_HVT U1559 ( .A1(sram_raddr_weight[13]), .A2(sram_raddr_weight[12]), 
        .A3(n1406), .Y(n1399) );
  NAND2X0_HVT U1560 ( .A1(n1455), .A2(n1399), .Y(n1403) );
  NAND2X0_HVT U1561 ( .A1(n1400), .A2(n1403), .Y(n1401) );
  AO222X1_HVT U1562 ( .A1(n403), .A2(n1402), .A3(n403), .A4(n1404), .A5(
        sram_raddr_weight[14]), .A6(n1401), .Y(net22706) );
  AO22X1_HVT U1563 ( .A1(n204), .A2(n1405), .A3(n1455), .A4(n1409), .Y(n1408)
         );
  AO22X1_HVT U1564 ( .A1(n207), .A2(n1410), .A3(n1406), .A4(n1455), .Y(n1407)
         );
  AO22X1_HVT U1565 ( .A1(sram_raddr_weight[12]), .A2(n1408), .A3(n429), .A4(
        n1407), .Y(net22720) );
  AND2X1_HVT U1566 ( .A1(n1455), .A2(n1411), .Y(n1422) );
  AO22X1_HVT U1567 ( .A1(n203), .A2(n1412), .A3(n288), .A4(n1455), .Y(n1415)
         );
  OR2X1_HVT U1568 ( .A1(n221), .A2(n1412), .Y(n1421) );
  NAND3X0_HVT U1569 ( .A1(sram_raddr_weight[9]), .A2(n1417), .A3(n1455), .Y(
        n1413) );
  NAND2X0_HVT U1570 ( .A1(n1421), .A2(n1413), .Y(n1414) );
  AO222X1_HVT U1571 ( .A1(sram_raddr_weight[10]), .A2(n1422), .A3(
        sram_raddr_weight[10]), .A4(n1415), .A5(n430), .A6(n1414), .Y(net22734) );
  NAND3X0_HVT U1572 ( .A1(n1417), .A2(n288), .A3(n1455), .Y(n1420) );
  AO221X1_HVT U1573 ( .A1(n204), .A2(sram_raddr_weight[8]), .A3(n1557), .A4(
        n1429), .A5(n1422), .Y(n1418) );
  NAND2X0_HVT U1574 ( .A1(sram_raddr_weight[9]), .A2(n1418), .Y(n1419) );
  NAND4X0_HVT U1575 ( .A1(n399), .A2(n1421), .A3(n1420), .A4(n1419), .Y(
        net22748) );
  NAND2X0_HVT U1576 ( .A1(n1422), .A2(n1423), .Y(n1427) );
  OA22X1_HVT U1577 ( .A1(n1424), .A2(n228), .A3(n1465), .A4(n1423), .Y(n1425)
         );
  AO222X1_HVT U1578 ( .A1(n355), .A2(n221), .A3(n355), .A4(n1429), .A5(
        sram_raddr_weight[8]), .A6(n1425), .Y(n1426) );
  NAND3X0_HVT U1579 ( .A1(n1427), .A2(n1426), .A3(n399), .Y(net22755) );
  OA22X1_HVT U1580 ( .A1(n1428), .A2(n228), .A3(n1465), .A4(n1434), .Y(n1430)
         );
  OA22X1_HVT U1581 ( .A1(n1430), .A2(n359), .A3(n221), .A4(n1429), .Y(n1432)
         );
  NAND3X0_HVT U1582 ( .A1(n1434), .A2(n359), .A3(n1455), .Y(n1431) );
  NAND3X0_HVT U1583 ( .A1(n399), .A2(n1432), .A3(n1431), .Y(net22783) );
  AO22X1_HVT U1584 ( .A1(n203), .A2(n1436), .A3(n1455), .A4(n1435), .Y(n1437)
         );
  NAND2X0_HVT U1585 ( .A1(n1455), .A2(n1440), .Y(n1450) );
  NAND4X0_HVT U1586 ( .A1(n205), .A2(n1441), .A3(n432), .A4(n305), .Y(n1453)
         );
  NAND3X0_HVT U1587 ( .A1(n1456), .A2(n1450), .A3(n1453), .Y(n1448) );
  NAND2X0_HVT U1588 ( .A1(n1441), .A2(n305), .Y(n1449) );
  OR2X1_HVT U1589 ( .A1(sram_raddr_weight[3]), .A2(n1449), .Y(n1442) );
  AO22X1_HVT U1590 ( .A1(n1444), .A2(n1455), .A3(n1443), .A4(n1442), .Y(n1447)
         );
  NAND3X0_HVT U1591 ( .A1(n1023), .A2(n253), .A3(state[2]), .Y(n1561) );
  NAND3X0_HVT U1592 ( .A1(n1023), .A2(n1024), .A3(n1445), .Y(n1550) );
  NAND4X0_HVT U1593 ( .A1(n1464), .A2(n1446), .A3(n1561), .A4(n1550), .Y(n1459) );
  AO221X1_HVT U1594 ( .A1(sram_raddr_weight[4]), .A2(n1448), .A3(n447), .A4(
        n1447), .A5(n1459), .Y(net22811) );
  NAND3X0_HVT U1595 ( .A1(sram_raddr_weight[2]), .A2(sram_raddr_weight[0]), 
        .A3(sram_raddr_weight[1]), .Y(n1451) );
  AOI22X1_HVT U1596 ( .A1(n203), .A2(n1449), .A3(n1455), .A4(n1451), .Y(n1452)
         );
  OA22X1_HVT U1597 ( .A1(n1452), .A2(n432), .A3(n1451), .A4(n1450), .Y(n1454)
         );
  NAND3X0_HVT U1598 ( .A1(n399), .A2(n1454), .A3(n1453), .Y(net22818) );
  NAND2X0_HVT U1599 ( .A1(sram_raddr_weight[0]), .A2(sram_raddr_weight[1]), 
        .Y(n1458) );
  NAND2X0_HVT U1600 ( .A1(n1455), .A2(n1458), .Y(n1462) );
  NAND2X0_HVT U1601 ( .A1(n1456), .A2(n1462), .Y(n1461) );
  OAI21X1_HVT U1602 ( .A1(n1458), .A2(n1465), .A3(n1457), .Y(n1460) );
  AO221X1_HVT U1603 ( .A1(sram_raddr_weight[2]), .A2(n1461), .A3(n305), .A4(
        n1460), .A5(n1459), .Y(net22825) );
  AO222X1_HVT U1604 ( .A1(n436), .A2(n1462), .A3(n436), .A4(n309), .A5(n1462), 
        .A6(n221), .Y(n1463) );
  NAND2X0_HVT U1605 ( .A1(n1464), .A2(n1463), .Y(net22839) );
  AO22X1_HVT U1606 ( .A1(sram_raddr_weight[0]), .A2(n221), .A3(n309), .A4(
        n1465), .Y(n1467) );
  NAND3X0_HVT U1607 ( .A1(n1467), .A2(n1466), .A3(n1561), .Y(net22853) );
  NAND2X0_HVT U1608 ( .A1(write_col_conv1[0]), .A2(n1468), .Y(n1507) );
  AO21X1_HVT U1609 ( .A1(n1470), .A2(n1469), .A3(N2914), .Y(net22861) );
  NAND2X0_HVT U1610 ( .A1(n1472), .A2(write_row_conv1[0]), .Y(n1476) );
  NAND3X0_HVT U1611 ( .A1(write_col_conv1[0]), .A2(n1473), .A3(n1476), .Y(
        n1498) );
  NAND2X0_HVT U1612 ( .A1(n1494), .A2(n344), .Y(n1492) );
  NOR2X0_HVT U1613 ( .A1(n1492), .A2(delay1_sram_waddr_b[5]), .Y(n1488) );
  NAND2X0_HVT U1614 ( .A1(n1488), .A2(n408), .Y(n1486) );
  NOR2X0_HVT U1615 ( .A1(n1486), .A2(delay1_sram_waddr_b[7]), .Y(n1483) );
  NAND2X0_HVT U1616 ( .A1(n1483), .A2(n445), .Y(n1474) );
  HADDX1_HVT U1617 ( .A0(delay1_sram_waddr_b[9]), .B0(n1474), .SO(n1479) );
  NAND4X0_HVT U1618 ( .A1(delay1_sram_waddr_b[0]), .A2(delay1_sram_waddr_b[1]), 
        .A3(delay1_sram_waddr_b[2]), .A4(delay1_sram_waddr_b[3]), .Y(n1495) );
  NOR2X0_HVT U1619 ( .A1(n344), .A2(n1495), .Y(n1493) );
  NAND2X0_HVT U1620 ( .A1(delay1_sram_waddr_b[5]), .A2(n1493), .Y(n1489) );
  NOR2X0_HVT U1621 ( .A1(n408), .A2(n1489), .Y(n1487) );
  AND2X1_HVT U1622 ( .A1(delay1_sram_waddr_b[7]), .A2(n1487), .Y(n1482) );
  NAND2X0_HVT U1623 ( .A1(delay1_sram_waddr_b[8]), .A2(n1482), .Y(n1477) );
  HADDX1_HVT U1624 ( .A0(delay1_sram_waddr_b[9]), .B0(n1477), .SO(n1478) );
  OAI22X1_HVT U1625 ( .A1(n1498), .A2(n1479), .A3(n1500), .A4(n1478), .Y(
        net22864) );
  OAI22X1_HVT U1626 ( .A1(n1483), .A2(n1498), .A3(n1482), .A4(n1500), .Y(n1481) );
  AO22X1_HVT U1627 ( .A1(n1505), .A2(n1483), .A3(n1506), .A4(n1482), .Y(n1480)
         );
  AO22X1_HVT U1628 ( .A1(delay1_sram_waddr_b[8]), .A2(n1481), .A3(n445), .A4(
        n1480), .Y(net22867) );
  OA221X1_HVT U1629 ( .A1(n1483), .A2(delay1_sram_waddr_b[7]), .A3(n1483), 
        .A4(n1486), .A5(n1505), .Y(n1484) );
  AO221X1_HVT U1630 ( .A1(n1485), .A2(delay1_sram_waddr_b[7]), .A3(n1485), 
        .A4(n1487), .A5(n1484), .Y(net22870) );
  AO21X1_HVT U1631 ( .A1(delay1_sram_waddr_b[5]), .A2(n1492), .A3(n1488), .Y(
        n1491) );
  OA21X1_HVT U1632 ( .A1(delay1_sram_waddr_b[5]), .A2(n1493), .A3(n1489), .Y(
        n1490) );
  AO22X1_HVT U1633 ( .A1(n1505), .A2(n1491), .A3(n1506), .A4(n1490), .Y(
        net22876) );
  OR3X1_HVT U1634 ( .A1(delay1_sram_waddr_b[0]), .A2(delay1_sram_waddr_b[1]), 
        .A3(delay1_sram_waddr_b[2]), .Y(n1499) );
  AO21X1_HVT U1635 ( .A1(delay1_sram_waddr_b[3]), .A2(n1499), .A3(n1494), .Y(
        n1497) );
  AND3X1_HVT U1636 ( .A1(delay1_sram_waddr_b[0]), .A2(delay1_sram_waddr_b[1]), 
        .A3(delay1_sram_waddr_b[2]), .Y(n1501) );
  OA21X1_HVT U1637 ( .A1(delay1_sram_waddr_b[3]), .A2(n1501), .A3(n1495), .Y(
        n1496) );
  AO22X1_HVT U1638 ( .A1(n1505), .A2(n1497), .A3(n1506), .A4(n1496), .Y(
        net22882) );
  OR2X1_HVT U1639 ( .A1(delay1_sram_waddr_b[0]), .A2(delay1_sram_waddr_b[1]), 
        .Y(n1503) );
  NAND2X0_HVT U1640 ( .A1(delay1_sram_waddr_b[0]), .A2(delay1_sram_waddr_b[1]), 
        .Y(n1502) );
  NAND2X0_HVT U1641 ( .A1(n1503), .A2(n1502), .Y(n1504) );
  MUX21X1_HVT U1642 ( .A1(n1506), .A2(n1505), .S0(n1504), .Y(net22888) );
  NOR2X0_HVT U1643 ( .A1(n1507), .A2(delay1_sram_waddr_b[0]), .Y(net22891) );
  AND4X1_HVT U1644 ( .A1(delay3_state[2]), .A2(n1027), .A3(delay3_state[0]), 
        .A4(delay3_state[1]), .Y(n1528) );
  NAND4X0_HVT U1645 ( .A1(n1528), .A2(delay3_addr_change[0]), .A3(
        delay3_addr_change[1]), .A4(n1508), .Y(n1511) );
  NAND2X0_HVT U1646 ( .A1(delay3_state[2]), .A2(n1027), .Y(n1509) );
  OR3X1_HVT U1647 ( .A1(delay3_state[0]), .A2(delay3_state[1]), .A3(n1509), 
        .Y(n1510) );
  NAND3X0_HVT U1648 ( .A1(n182), .A2(n1511), .A3(n1510), .Y(net22899) );
  NAND4X0_HVT U1649 ( .A1(delay1_sram_waddr_c[0]), .A2(delay1_sram_waddr_c[1]), 
        .A3(delay1_sram_waddr_c[2]), .A4(delay1_sram_waddr_c[3]), .Y(n1524) );
  NAND2X0_HVT U1650 ( .A1(n1523), .A2(delay1_sram_waddr_c[4]), .Y(n1522) );
  NAND2X0_HVT U1651 ( .A1(n1521), .A2(delay1_sram_waddr_c[5]), .Y(n1520) );
  NAND2X0_HVT U1652 ( .A1(n1519), .A2(delay1_sram_waddr_c[6]), .Y(n1518) );
  NAND2X0_HVT U1653 ( .A1(n1517), .A2(delay1_sram_waddr_c[7]), .Y(n1516) );
  NAND2X0_HVT U1654 ( .A1(n1515), .A2(delay1_sram_waddr_c[8]), .Y(n1514) );
  OA221X1_HVT U1655 ( .A1(n1513), .A2(delay1_sram_waddr_c[9]), .A3(n1514), 
        .A4(n467), .A5(n1527), .Y(net22901) );
  NAND3X0_HVT U1656 ( .A1(delay1_sram_waddr_c[0]), .A2(delay1_sram_waddr_c[1]), 
        .A3(delay1_sram_waddr_c[2]), .Y(n1525) );
  NAND2X0_HVT U1657 ( .A1(delay1_sram_waddr_c[0]), .A2(delay1_sram_waddr_c[1]), 
        .Y(n1526) );
  AND2X1_HVT U1658 ( .A1(n1527), .A2(n440), .Y(net22910) );
  NAND4X0_HVT U1659 ( .A1(delay1_sram_waddr_d[0]), .A2(delay1_sram_waddr_d[1]), 
        .A3(delay1_sram_waddr_d[2]), .A4(delay1_sram_waddr_d[3]), .Y(n1540) );
  NAND2X0_HVT U1660 ( .A1(n1539), .A2(delay1_sram_waddr_d[4]), .Y(n1538) );
  NAND2X0_HVT U1661 ( .A1(n1537), .A2(delay1_sram_waddr_d[5]), .Y(n1536) );
  NAND2X0_HVT U1662 ( .A1(n1535), .A2(delay1_sram_waddr_d[6]), .Y(n1534) );
  NAND2X0_HVT U1663 ( .A1(n1533), .A2(delay1_sram_waddr_d[7]), .Y(n1532) );
  NAND2X0_HVT U1664 ( .A1(n1531), .A2(delay1_sram_waddr_d[8]), .Y(n1530) );
  OA221X1_HVT U1665 ( .A1(n1529), .A2(delay1_sram_waddr_d[9]), .A3(n1530), 
        .A4(n468), .A5(n1543), .Y(net22917) );
  NAND3X0_HVT U1666 ( .A1(delay1_sram_waddr_d[0]), .A2(delay1_sram_waddr_d[1]), 
        .A3(delay1_sram_waddr_d[2]), .Y(n1541) );
  NAND2X0_HVT U1667 ( .A1(delay1_sram_waddr_d[0]), .A2(delay1_sram_waddr_d[1]), 
        .Y(n1542) );
  AND2X1_HVT U1668 ( .A1(n1543), .A2(n441), .Y(net22926) );
  NAND2X0_HVT U1669 ( .A1(n1544), .A2(n182), .Y(net22933) );
  NAND3X0_HVT U1670 ( .A1(n1547), .A2(channel_cnt[2]), .A3(channel_cnt[3]), 
        .Y(n1546) );
  OA221X1_HVT U1671 ( .A1(channel_cnt[4]), .A2(n1545), .A3(n314), .A4(n1546), 
        .A5(n1549), .Y(net22934) );
  OA221X1_HVT U1672 ( .A1(n1547), .A2(channel_cnt[2]), .A3(n1548), .A4(n435), 
        .A5(n1549), .Y(net22936) );
  NAND3X0_HVT U1673 ( .A1(n183), .A2(n221), .A3(n1550), .Y(net22944) );
  NAND4X0_HVT U1674 ( .A1(addr_change[0]), .A2(addr_change[1]), .A3(
        addr_change[2]), .A4(addr_change[3]), .Y(n1553) );
  NAND4X0_HVT U1675 ( .A1(addr_change[1]), .A2(addr_change[0]), .A3(
        addr_change[4]), .A4(n454), .Y(n1551) );
  OA21X1_HVT U1676 ( .A1(addr_change[2]), .A2(n1551), .A3(n1557), .Y(n1556) );
  OA221X1_HVT U1677 ( .A1(addr_change[4]), .A2(n1552), .A3(n460), .A4(n1553), 
        .A5(n1556), .Y(net22946) );
  NAND3X0_HVT U1678 ( .A1(addr_change[0]), .A2(addr_change[1]), .A3(
        addr_change[2]), .Y(n1554) );
  NAND2X0_HVT U1679 ( .A1(addr_change[0]), .A2(addr_change[1]), .Y(n1555) );
  NOR2X0_HVT U1680 ( .A1(n228), .A2(addr_change[0]), .Y(net22950) );
  NAND4X0_HVT U1681 ( .A1(n1569), .A2(n1558), .A3(addr_row_sel_cnt[0]), .A4(
        addr_row_sel_cnt[1]), .Y(n1559) );
  OA221X1_HVT U1682 ( .A1(n1568), .A2(n1051), .A3(n1568), .A4(
        addr_col_sel_cnt[0]), .A5(n1559), .Y(n1892) );
  NAND2X0_HVT U1683 ( .A1(n181), .A2(n1934), .Y(net23893) );
  NAND2X0_HVT U1684 ( .A1(n182), .A2(n1989), .Y(net25220) );
  NAND2X0_HVT U1685 ( .A1(n183), .A2(n1887), .Y(net26550) );
  NOR2X0_HVT U1686 ( .A1(n240), .A2(n1561), .Y(n1022) );
  NAND3X0_HVT U1687 ( .A1(n1051), .A2(n1052), .A3(n1679), .Y(n1849) );
  AND4X1_HVT U1688 ( .A1(n1569), .A2(n2003), .A3(addr_row_sel_cnt[1]), .A4(
        n254), .Y(n1571) );
  AO22X1_HVT U1689 ( .A1(n1838), .A2(n306), .A3(n170), .A4(n433), .Y(n1572) );
  AO221X1_HVT U1690 ( .A1(sram_raddr_a0[0]), .A2(n1887), .A3(n431), .A4(n1614), 
        .A5(n1572), .Y(n_sram_raddr_a0[0]) );
  NAND2X0_HVT U1691 ( .A1(sram_raddr_a6[1]), .A2(sram_raddr_a6[0]), .Y(n1578)
         );
  OA21X1_HVT U1692 ( .A1(sram_raddr_a6[1]), .A2(sram_raddr_a6[0]), .A3(n1578), 
        .Y(n1850) );
  NAND2X0_HVT U1693 ( .A1(n519), .A2(n1850), .Y(n1735) );
  AO221X1_HVT U1694 ( .A1(n1759), .A2(n1577), .A3(n1759), .A4(sram_raddr_a0[0]), .A5(n422), .Y(n1575) );
  NAND3X0_HVT U1695 ( .A1(sram_raddr_a0[0]), .A2(n1614), .A3(n422), .Y(n1574)
         );
  NAND2X0_HVT U1696 ( .A1(sram_raddr_a3[1]), .A2(sram_raddr_a3[0]), .Y(n1580)
         );
  OA21X1_HVT U1697 ( .A1(sram_raddr_a3[1]), .A2(sram_raddr_a3[0]), .A3(n1580), 
        .Y(n1736) );
  NAND2X0_HVT U1698 ( .A1(n1974), .A2(n1736), .Y(n1573) );
  NAND4X0_HVT U1699 ( .A1(n1735), .A2(n1575), .A3(n1574), .A4(n1573), .Y(
        n_sram_raddr_a0[1]) );
  AND3X1_HVT U1700 ( .A1(sram_raddr_a0[2]), .A2(sram_raddr_a0[1]), .A3(
        sram_raddr_a0[0]), .Y(n1576) );
  OA21X1_HVT U1701 ( .A1(n1577), .A2(n1576), .A3(n1759), .Y(n1585) );
  AND3X1_HVT U1702 ( .A1(sram_raddr_a0[1]), .A2(sram_raddr_a0[0]), .A3(n1614), 
        .Y(n1581) );
  AO22X1_HVT U1703 ( .A1(n1582), .A2(n456), .A3(n1578), .A4(sram_raddr_a6[2]), 
        .Y(n1851) );
  AO22X1_HVT U1704 ( .A1(sram_raddr_a3[2]), .A2(n1580), .A3(n236), .A4(n1579), 
        .Y(n1738) );
  NAND4X0_HVT U1705 ( .A1(sram_raddr_a3[2]), .A2(sram_raddr_a3[3]), .A3(
        sram_raddr_a3[1]), .A4(sram_raddr_a3[0]), .Y(n1587) );
  AO221X1_HVT U1706 ( .A1(n244), .A2(n236), .A3(n244), .A4(n1580), .A5(n1586), 
        .Y(n1739) );
  OA22X1_HVT U1707 ( .A1(n1585), .A2(n239), .A3(n171), .A4(n1739), .Y(n1583)
         );
  NAND3X0_HVT U1708 ( .A1(sram_raddr_a0[2]), .A2(n1581), .A3(n239), .Y(n1584)
         );
  NAND4X0_HVT U1709 ( .A1(sram_raddr_a6[1]), .A2(sram_raddr_a6[0]), .A3(
        sram_raddr_a6[2]), .A4(sram_raddr_a6[3]), .Y(n1588) );
  OA221X1_HVT U1710 ( .A1(sram_raddr_a6[3]), .A2(sram_raddr_a6[2]), .A3(
        sram_raddr_a6[3]), .A4(n1582), .A5(n1588), .Y(n1852) );
  NAND2X0_HVT U1711 ( .A1(n167), .A2(n1852), .Y(n1740) );
  NAND3X0_HVT U1712 ( .A1(n1583), .A2(n1584), .A3(n1740), .Y(
        n_sram_raddr_a0[3]) );
  AND2X1_HVT U1713 ( .A1(n1585), .A2(n1584), .Y(n1595) );
  AND2X1_HVT U1714 ( .A1(sram_raddr_a3[4]), .A2(n1586), .Y(n1591) );
  AO21X1_HVT U1715 ( .A1(n275), .A2(n1587), .A3(n1591), .Y(n1745) );
  OA22X1_HVT U1716 ( .A1(n1595), .A2(n342), .A3(n189), .A4(n1745), .Y(n1590)
         );
  AND4X1_HVT U1717 ( .A1(sram_raddr_a0[3]), .A2(sram_raddr_a0[2]), .A3(
        sram_raddr_a0[1]), .A4(sram_raddr_a0[0]), .Y(n1600) );
  NAND3X0_HVT U1718 ( .A1(n1600), .A2(n1614), .A3(n342), .Y(n1594) );
  NAND2X0_HVT U1719 ( .A1(n1589), .A2(sram_raddr_a6[4]), .Y(n1592) );
  OA21X1_HVT U1720 ( .A1(n1589), .A2(sram_raddr_a6[4]), .A3(n1592), .Y(n1856)
         );
  NAND2X0_HVT U1721 ( .A1(n519), .A2(n1856), .Y(n1743) );
  NAND3X0_HVT U1722 ( .A1(n1590), .A2(n1594), .A3(n1743), .Y(
        n_sram_raddr_a0[4]) );
  NAND2X0_HVT U1723 ( .A1(sram_raddr_a3[5]), .A2(n1591), .Y(n1599) );
  OA21X1_HVT U1724 ( .A1(sram_raddr_a3[5]), .A2(n1591), .A3(n1599), .Y(n1747)
         );
  NAND2X0_HVT U1725 ( .A1(n170), .A2(n1747), .Y(n1598) );
  NAND2X0_HVT U1726 ( .A1(n1593), .A2(sram_raddr_a6[5]), .Y(n1601) );
  OA21X1_HVT U1727 ( .A1(n1593), .A2(sram_raddr_a6[5]), .A3(n1601), .Y(n1862)
         );
  NAND2X0_HVT U1728 ( .A1(n167), .A2(n1862), .Y(n1750) );
  NAND4X0_HVT U1729 ( .A1(sram_raddr_a0[4]), .A2(n1600), .A3(n1614), .A4(n284), 
        .Y(n1596) );
  AND3X1_HVT U1730 ( .A1(n1595), .A2(n1596), .A3(n1594), .Y(n1604) );
  AO21X1_HVT U1731 ( .A1(n284), .A2(n1596), .A3(n1604), .Y(n1597) );
  NAND3X0_HVT U1732 ( .A1(n1598), .A2(n1750), .A3(n1597), .Y(
        n_sram_raddr_a0[5]) );
  OR2X1_HVT U1733 ( .A1(n331), .A2(n1599), .Y(n1606) );
  AO21X1_HVT U1734 ( .A1(n331), .A2(n1599), .A3(n1605), .Y(n1755) );
  OA22X1_HVT U1735 ( .A1(n1604), .A2(n446), .A3(n189), .A4(n1755), .Y(n1602)
         );
  AND3X1_HVT U1736 ( .A1(sram_raddr_a0[5]), .A2(sram_raddr_a0[4]), .A3(n1600), 
        .Y(n1609) );
  NAND3X0_HVT U1737 ( .A1(n1609), .A2(n1614), .A3(n446), .Y(n1603) );
  AO22X1_HVT U1738 ( .A1(n1607), .A2(n464), .A3(n1601), .A4(sram_raddr_a6[6]), 
        .Y(n1867) );
  NAND2X0_HVT U1739 ( .A1(n1838), .A2(n1867), .Y(n1753) );
  NAND3X0_HVT U1740 ( .A1(n1602), .A2(n1603), .A3(n1753), .Y(
        n_sram_raddr_a0[6]) );
  AND2X1_HVT U1741 ( .A1(n1604), .A2(n1603), .Y(n1613) );
  AND2X1_HVT U1742 ( .A1(sram_raddr_a3[7]), .A2(n1605), .Y(n1618) );
  AO21X1_HVT U1743 ( .A1(n412), .A2(n1606), .A3(n1618), .Y(n1757) );
  OA22X1_HVT U1744 ( .A1(n1613), .A2(n397), .A3(n189), .A4(n1757), .Y(n1611)
         );
  AND2X1_HVT U1745 ( .A1(n1607), .A2(sram_raddr_a6[6]), .Y(n1608) );
  NAND2X0_HVT U1746 ( .A1(n1608), .A2(sram_raddr_a6[7]), .Y(n1616) );
  OA21X1_HVT U1747 ( .A1(n1608), .A2(sram_raddr_a6[7]), .A3(n1616), .Y(n1873)
         );
  NAND2X0_HVT U1748 ( .A1(n167), .A2(n1873), .Y(n1762) );
  AND2X1_HVT U1749 ( .A1(sram_raddr_a0[6]), .A2(n1609), .Y(n1615) );
  NAND3X0_HVT U1750 ( .A1(n1615), .A2(n397), .A3(n1614), .Y(n1610) );
  NAND3X0_HVT U1751 ( .A1(n1611), .A2(n1762), .A3(n1610), .Y(
        n_sram_raddr_a0[7]) );
  NAND2X0_HVT U1752 ( .A1(n397), .A2(n1614), .Y(n1612) );
  NAND2X0_HVT U1753 ( .A1(n1613), .A2(n1612), .Y(n1626) );
  AND3X1_HVT U1754 ( .A1(sram_raddr_a0[7]), .A2(n1615), .A3(n1614), .Y(n1624)
         );
  NAND2X0_HVT U1755 ( .A1(n1617), .A2(sram_raddr_a6[8]), .Y(n1620) );
  OA21X1_HVT U1756 ( .A1(n1617), .A2(sram_raddr_a6[8]), .A3(n1620), .Y(n1880)
         );
  NAND2X0_HVT U1757 ( .A1(sram_raddr_a3[8]), .A2(n1618), .Y(n1622) );
  OA21X1_HVT U1758 ( .A1(sram_raddr_a3[8]), .A2(n1618), .A3(n1622), .Y(n1765)
         );
  AO22X1_HVT U1759 ( .A1(n519), .A2(n1880), .A3(n170), .A4(n1765), .Y(n1619)
         );
  AO221X1_HVT U1760 ( .A1(sram_raddr_a0[8]), .A2(n1626), .A3(n424), .A4(n1624), 
        .A5(n1619), .Y(n_sram_raddr_a0[8]) );
  HADDX1_HVT U1761 ( .A0(sram_raddr_a6[9]), .B0(n1621), .SO(n1886) );
  AND2X1_HVT U1762 ( .A1(n519), .A2(n1886), .Y(n1772) );
  HADDX1_HVT U1763 ( .A0(sram_raddr_a3[9]), .B0(n1623), .SO(n1770) );
  HADDX1_HVT U1764 ( .A0(sram_raddr_a0[9]), .B0(sram_raddr_a0[8]), .SO(n1625)
         );
  NAND2X0_HVT U1765 ( .A1(n_addr_col_sel_cnt[1]), .A2(n254), .Y(n1913) );
  AO22X1_HVT U1766 ( .A1(n1838), .A2(n303), .A3(n170), .A4(n417), .Y(n1627) );
  AO221X1_HVT U1767 ( .A1(sram_raddr_a1[0]), .A2(n1934), .A3(n310), .A4(n1664), 
        .A5(n1627), .Y(n_sram_raddr_a1[0]) );
  NAND2X0_HVT U1768 ( .A1(sram_raddr_a4[1]), .A2(sram_raddr_a4[0]), .Y(n1628)
         );
  AO21X1_HVT U1769 ( .A1(n307), .A2(n417), .A3(n1629), .Y(n1774) );
  AO22X1_HVT U1770 ( .A1(sram_raddr_a7[1]), .A2(n303), .A3(n443), .A4(
        sram_raddr_a7[0]), .Y(n1891) );
  NAND2X0_HVT U1771 ( .A1(n167), .A2(n1891), .Y(n1775) );
  AND2X1_HVT U1772 ( .A1(sram_raddr_a1[1]), .A2(sram_raddr_a1[0]), .Y(n1637)
         );
  NAND3X0_HVT U1773 ( .A1(sram_raddr_a1[2]), .A2(sram_raddr_a1[1]), .A3(
        sram_raddr_a1[0]), .Y(n1635) );
  AO21X1_HVT U1774 ( .A1(n1664), .A2(n1635), .A3(n1934), .Y(n1630) );
  AO22X1_HVT U1775 ( .A1(sram_raddr_a4[2]), .A2(n1628), .A3(n237), .A4(n1629), 
        .Y(n1777) );
  NAND3X0_HVT U1776 ( .A1(sram_raddr_a7[1]), .A2(sram_raddr_a7[0]), .A3(
        sram_raddr_a7[2]), .Y(n1631) );
  OA221X1_HVT U1777 ( .A1(sram_raddr_a7[2]), .A2(sram_raddr_a7[0]), .A3(
        sram_raddr_a7[2]), .A4(sram_raddr_a7[1]), .A5(n1631), .Y(n1897) );
  NAND4X0_HVT U1778 ( .A1(sram_raddr_a4[2]), .A2(sram_raddr_a4[3]), .A3(
        sram_raddr_a4[1]), .A4(sram_raddr_a4[0]), .Y(n1636) );
  OA221X1_HVT U1779 ( .A1(sram_raddr_a4[3]), .A2(sram_raddr_a4[2]), .A3(
        sram_raddr_a4[3]), .A4(n1629), .A5(n1636), .Y(n1778) );
  AOI22X1_HVT U1780 ( .A1(sram_raddr_a1[3]), .A2(n1630), .A3(n170), .A4(n1778), 
        .Y(n1634) );
  NAND4X0_HVT U1781 ( .A1(sram_raddr_a1[2]), .A2(n1637), .A3(n1664), .A4(n238), 
        .Y(n1633) );
  AO22X1_HVT U1782 ( .A1(n1632), .A2(n466), .A3(n1631), .A4(sram_raddr_a7[3]), 
        .Y(n1898) );
  NAND2X0_HVT U1783 ( .A1(n1838), .A2(n1898), .Y(n1779) );
  NAND3X0_HVT U1784 ( .A1(n1634), .A2(n1633), .A3(n1779), .Y(
        n_sram_raddr_a1[3]) );
  AOI221X1_HVT U1785 ( .A1(n1664), .A2(n238), .A3(n1664), .A4(n1635), .A5(
        n1934), .Y(n1641) );
  NOR2X0_HVT U1786 ( .A1(n246), .A2(n1636), .Y(n1642) );
  AO21X1_HVT U1787 ( .A1(n246), .A2(n1636), .A3(n1642), .Y(n1781) );
  OA22X1_HVT U1788 ( .A1(n1641), .A2(n278), .A3(n171), .A4(n1781), .Y(n1639)
         );
  AND4X1_HVT U1789 ( .A1(sram_raddr_a1[3]), .A2(sram_raddr_a1[2]), .A3(n1637), 
        .A4(n1664), .Y(n1643) );
  NAND2X0_HVT U1790 ( .A1(n1643), .A2(n278), .Y(n1640) );
  AND4X1_HVT U1791 ( .A1(sram_raddr_a7[1]), .A2(sram_raddr_a7[0]), .A3(
        sram_raddr_a7[2]), .A4(sram_raddr_a7[3]), .Y(n1638) );
  NAND2X0_HVT U1792 ( .A1(n1638), .A2(sram_raddr_a7[4]), .Y(n1644) );
  OA21X1_HVT U1793 ( .A1(n1638), .A2(sram_raddr_a7[4]), .A3(n1644), .Y(n1902)
         );
  NAND2X0_HVT U1794 ( .A1(n167), .A2(n1902), .Y(n1784) );
  NAND3X0_HVT U1795 ( .A1(n1639), .A2(n1640), .A3(n1784), .Y(
        n_sram_raddr_a1[4]) );
  AND2X1_HVT U1796 ( .A1(n1641), .A2(n1640), .Y(n1648) );
  NAND2X0_HVT U1797 ( .A1(sram_raddr_a4[5]), .A2(n1642), .Y(n1649) );
  OA22X1_HVT U1798 ( .A1(n1648), .A2(n345), .A3(n189), .A4(n1786), .Y(n1646)
         );
  AND2X1_HVT U1799 ( .A1(sram_raddr_a1[4]), .A2(n1643), .Y(n1650) );
  NAND2X0_HVT U1800 ( .A1(n1650), .A2(n345), .Y(n1647) );
  NAND2X0_HVT U1801 ( .A1(n1645), .A2(sram_raddr_a7[5]), .Y(n1651) );
  OA21X1_HVT U1802 ( .A1(n1645), .A2(sram_raddr_a7[5]), .A3(n1651), .Y(n1908)
         );
  NAND2X0_HVT U1803 ( .A1(n167), .A2(n1908), .Y(n1788) );
  NAND3X0_HVT U1804 ( .A1(n1646), .A2(n1647), .A3(n1788), .Y(
        n_sram_raddr_a1[5]) );
  AND2X1_HVT U1805 ( .A1(n1648), .A2(n1647), .Y(n1656) );
  AO21X1_HVT U1806 ( .A1(n333), .A2(n1649), .A3(n1660), .Y(n1793) );
  OA22X1_HVT U1807 ( .A1(n1656), .A2(n448), .A3(n189), .A4(n1793), .Y(n1653)
         );
  AND2X1_HVT U1808 ( .A1(sram_raddr_a1[5]), .A2(n1650), .Y(n1657) );
  NAND2X0_HVT U1809 ( .A1(n1657), .A2(n448), .Y(n1654) );
  NAND2X0_HVT U1810 ( .A1(n1652), .A2(sram_raddr_a7[6]), .Y(n1658) );
  OA21X1_HVT U1811 ( .A1(n1652), .A2(sram_raddr_a7[6]), .A3(n1658), .Y(n1914)
         );
  NAND2X0_HVT U1812 ( .A1(n1838), .A2(n1914), .Y(n1791) );
  NAND3X0_HVT U1813 ( .A1(n1653), .A2(n1654), .A3(n1791), .Y(
        n_sram_raddr_a1[6]) );
  NAND2X0_HVT U1814 ( .A1(n1656), .A2(n1654), .Y(n1663) );
  AND2X1_HVT U1815 ( .A1(sram_raddr_a1[6]), .A2(n1657), .Y(n1665) );
  NAND2X0_HVT U1816 ( .A1(n1659), .A2(sram_raddr_a7[7]), .Y(n1666) );
  OA21X1_HVT U1817 ( .A1(n1659), .A2(sram_raddr_a7[7]), .A3(n1666), .Y(n1922)
         );
  NAND2X0_HVT U1818 ( .A1(sram_raddr_a4[7]), .A2(n1660), .Y(n1669) );
  OA21X1_HVT U1819 ( .A1(sram_raddr_a4[7]), .A2(n1660), .A3(n1669), .Y(n1797)
         );
  AO22X1_HVT U1820 ( .A1(n519), .A2(n1922), .A3(n1974), .A4(n1797), .Y(n1661)
         );
  AO221X1_HVT U1821 ( .A1(sram_raddr_a1[7]), .A2(n1663), .A3(n438), .A4(n1665), 
        .A5(n1661), .Y(n_sram_raddr_a1[7]) );
  AO21X1_HVT U1822 ( .A1(n438), .A2(n1664), .A3(n1663), .Y(n1678) );
  AND2X1_HVT U1823 ( .A1(sram_raddr_a1[7]), .A2(n1665), .Y(n1676) );
  NAND2X0_HVT U1824 ( .A1(n1668), .A2(sram_raddr_a7[8]), .Y(n1672) );
  OA21X1_HVT U1825 ( .A1(n1668), .A2(sram_raddr_a7[8]), .A3(n1672), .Y(n1925)
         );
  NAND2X0_HVT U1826 ( .A1(sram_raddr_a4[8]), .A2(n1670), .Y(n1674) );
  OA21X1_HVT U1827 ( .A1(sram_raddr_a4[8]), .A2(n1670), .A3(n1674), .Y(n1799)
         );
  AO22X1_HVT U1828 ( .A1(n519), .A2(n1925), .A3(n170), .A4(n1799), .Y(n1671)
         );
  AO221X1_HVT U1829 ( .A1(sram_raddr_a1[8]), .A2(n1678), .A3(n425), .A4(n1676), 
        .A5(n1671), .Y(n_sram_raddr_a1[8]) );
  HADDX1_HVT U1830 ( .A0(sram_raddr_a7[9]), .B0(n1673), .SO(n1932) );
  AND2X1_HVT U1831 ( .A1(n1838), .A2(n1932), .Y(n1806) );
  HADDX1_HVT U1832 ( .A0(sram_raddr_a4[9]), .B0(n1675), .SO(n1804) );
  HADDX1_HVT U1833 ( .A0(sram_raddr_a1[9]), .B0(sram_raddr_a1[8]), .SO(n1677)
         );
  NAND3X0_HVT U1834 ( .A1(n1052), .A2(n1679), .A3(addr_col_sel_cnt[1]), .Y(
        n1941) );
  AO22X1_HVT U1835 ( .A1(n1838), .A2(n302), .A3(n1974), .A4(n416), .Y(n1680)
         );
  AO221X1_HVT U1836 ( .A1(sram_raddr_a2[0]), .A2(n1989), .A3(n442), .A4(n1721), 
        .A5(n1680), .Y(n_sram_raddr_a2[0]) );
  AO22X1_HVT U1837 ( .A1(sram_raddr_a8[1]), .A2(n302), .A3(n451), .A4(
        sram_raddr_a8[0]), .Y(n1938) );
  NAND2X0_HVT U1838 ( .A1(sram_raddr_a5[1]), .A2(sram_raddr_a5[0]), .Y(n1687)
         );
  OA21X1_HVT U1839 ( .A1(sram_raddr_a5[1]), .A2(sram_raddr_a5[0]), .A3(n1687), 
        .Y(n1807) );
  NAND2X0_HVT U1840 ( .A1(sram_raddr_a2[1]), .A2(sram_raddr_a2[0]), .Y(n1685)
         );
  OA21X1_HVT U1841 ( .A1(sram_raddr_a2[1]), .A2(sram_raddr_a2[0]), .A3(n1685), 
        .Y(n1681) );
  AO222X1_HVT U1842 ( .A1(n1838), .A2(n1938), .A3(n170), .A4(n1807), .A5(n1681), .A6(n1896), .Y(n1940) );
  AO22X1_HVT U1843 ( .A1(n1981), .A2(n1681), .A3(sram_raddr_a2[1]), .A4(n1989), 
        .Y(n1682) );
  OR2X1_HVT U1844 ( .A1(n1940), .A2(n1682), .Y(n_sram_raddr_a2[1]) );
  NAND2X0_HVT U1845 ( .A1(sram_raddr_a8[1]), .A2(sram_raddr_a8[0]), .Y(n1683)
         );
  AND3X1_HVT U1846 ( .A1(sram_raddr_a8[1]), .A2(sram_raddr_a8[0]), .A3(
        sram_raddr_a8[2]), .Y(n1689) );
  AO21X1_HVT U1847 ( .A1(n1683), .A2(n452), .A3(n1689), .Y(n1943) );
  NAND3X0_HVT U1848 ( .A1(sram_raddr_a5[2]), .A2(sram_raddr_a5[1]), .A3(
        sram_raddr_a5[0]), .Y(n1684) );
  NAND2X0_HVT U1849 ( .A1(n360), .A2(n1687), .Y(n1951) );
  NAND2X0_HVT U1850 ( .A1(n1684), .A2(n1951), .Y(n1946) );
  OA22X1_HVT U1851 ( .A1(n1942), .A2(n1943), .A3(n171), .A4(n1946), .Y(n1811)
         );
  AND3X1_HVT U1852 ( .A1(sram_raddr_a2[2]), .A2(sram_raddr_a2[1]), .A3(
        sram_raddr_a2[0]), .Y(n1707) );
  AND2X1_HVT U1853 ( .A1(n366), .A2(n1685), .Y(n1813) );
  OR2X1_HVT U1854 ( .A1(n1707), .A2(n1813), .Y(n1809) );
  OA22X1_HVT U1855 ( .A1(n1692), .A2(n1809), .A3(n1945), .A4(n366), .Y(n1686)
         );
  NAND2X0_HVT U1856 ( .A1(n1811), .A2(n1686), .Y(n_sram_raddr_a2[2]) );
  OA21X1_HVT U1857 ( .A1(n1692), .A2(n1707), .A3(n1945), .Y(n1688) );
  AND4X1_HVT U1858 ( .A1(sram_raddr_a5[3]), .A2(sram_raddr_a5[2]), .A3(
        sram_raddr_a5[1]), .A4(sram_raddr_a5[0]), .Y(n1693) );
  AO221X1_HVT U1859 ( .A1(n274), .A2(n360), .A3(n274), .A4(n1687), .A5(n1693), 
        .Y(n1812) );
  OA22X1_HVT U1860 ( .A1(n1688), .A2(n343), .A3(n171), .A4(n1812), .Y(n1691)
         );
  NAND3X0_HVT U1861 ( .A1(n1707), .A2(n1721), .A3(n343), .Y(n1690) );
  NAND4X0_HVT U1862 ( .A1(sram_raddr_a8[1]), .A2(sram_raddr_a8[0]), .A3(
        sram_raddr_a8[2]), .A4(sram_raddr_a8[3]), .Y(n1694) );
  OA21X1_HVT U1863 ( .A1(n1689), .A2(sram_raddr_a8[3]), .A3(n1694), .Y(n1950)
         );
  NAND2X0_HVT U1864 ( .A1(n167), .A2(n1950), .Y(n1814) );
  NAND3X0_HVT U1865 ( .A1(n1691), .A2(n1690), .A3(n1814), .Y(
        n_sram_raddr_a2[3]) );
  OA221X1_HVT U1866 ( .A1(n1692), .A2(sram_raddr_a2[3]), .A3(n1692), .A4(n1707), .A5(n1945), .Y(n1698) );
  NAND2X0_HVT U1867 ( .A1(sram_raddr_a5[4]), .A2(n1693), .Y(n1699) );
  OA22X1_HVT U1868 ( .A1(n1698), .A2(n341), .A3(n171), .A4(n1816), .Y(n1696)
         );
  NAND4X0_HVT U1869 ( .A1(sram_raddr_a2[3]), .A2(n1707), .A3(n1721), .A4(n341), 
        .Y(n1697) );
  NAND2X0_HVT U1870 ( .A1(n1695), .A2(sram_raddr_a8[4]), .Y(n1701) );
  OA21X1_HVT U1871 ( .A1(n1695), .A2(sram_raddr_a8[4]), .A3(n1701), .Y(n1955)
         );
  NAND2X0_HVT U1872 ( .A1(n519), .A2(n1955), .Y(n1818) );
  NAND3X0_HVT U1873 ( .A1(n1696), .A2(n1697), .A3(n1818), .Y(
        n_sram_raddr_a2[4]) );
  AND2X1_HVT U1874 ( .A1(n1698), .A2(n1697), .Y(n1705) );
  NOR2X0_HVT U1875 ( .A1(n332), .A2(n1699), .Y(n1706) );
  AO21X1_HVT U1876 ( .A1(n332), .A2(n1699), .A3(n1706), .Y(n1820) );
  OA22X1_HVT U1877 ( .A1(n1705), .A2(n348), .A3(n171), .A4(n1820), .Y(n1703)
         );
  AND3X1_HVT U1878 ( .A1(sram_raddr_a2[4]), .A2(sram_raddr_a2[3]), .A3(n1707), 
        .Y(n1700) );
  NAND3X0_HVT U1879 ( .A1(n1700), .A2(n1721), .A3(n348), .Y(n1704) );
  NAND2X0_HVT U1880 ( .A1(n1702), .A2(sram_raddr_a8[5]), .Y(n1708) );
  OA21X1_HVT U1881 ( .A1(n1702), .A2(sram_raddr_a8[5]), .A3(n1708), .Y(n1961)
         );
  NAND2X0_HVT U1882 ( .A1(n1838), .A2(n1961), .Y(n1823) );
  NAND3X0_HVT U1883 ( .A1(n1703), .A2(n1704), .A3(n1823), .Y(
        n_sram_raddr_a2[5]) );
  AND2X1_HVT U1884 ( .A1(n1705), .A2(n1704), .Y(n1712) );
  NAND2X0_HVT U1885 ( .A1(sram_raddr_a5[6]), .A2(n1706), .Y(n1713) );
  OA22X1_HVT U1886 ( .A1(n1712), .A2(n410), .A3(n189), .A4(n1825), .Y(n1710)
         );
  AND4X1_HVT U1887 ( .A1(sram_raddr_a2[5]), .A2(sram_raddr_a2[4]), .A3(
        sram_raddr_a2[3]), .A4(n1707), .Y(n1716) );
  NAND3X0_HVT U1888 ( .A1(n1716), .A2(n1721), .A3(n410), .Y(n1711) );
  NAND2X0_HVT U1889 ( .A1(n1709), .A2(sram_raddr_a8[6]), .Y(n1714) );
  OA21X1_HVT U1890 ( .A1(n1709), .A2(sram_raddr_a8[6]), .A3(n1714), .Y(n1966)
         );
  NAND2X0_HVT U1891 ( .A1(n519), .A2(n1966), .Y(n1827) );
  NAND3X0_HVT U1892 ( .A1(n1710), .A2(n1711), .A3(n1827), .Y(
        n_sram_raddr_a2[6]) );
  AND2X1_HVT U1893 ( .A1(n1712), .A2(n1711), .Y(n1720) );
  AO21X1_HVT U1894 ( .A1(n396), .A2(n1713), .A3(n1725), .Y(n1829) );
  OA22X1_HVT U1895 ( .A1(n1720), .A2(n398), .A3(n171), .A4(n1829), .Y(n1718)
         );
  NAND2X0_HVT U1896 ( .A1(n1715), .A2(sram_raddr_a8[7]), .Y(n1723) );
  OA21X1_HVT U1897 ( .A1(n1715), .A2(sram_raddr_a8[7]), .A3(n1723), .Y(n1972)
         );
  NAND2X0_HVT U1898 ( .A1(n167), .A2(n1972), .Y(n1834) );
  AND2X1_HVT U1899 ( .A1(sram_raddr_a2[6]), .A2(n1716), .Y(n1722) );
  NAND3X0_HVT U1900 ( .A1(n1722), .A2(n398), .A3(n1721), .Y(n1717) );
  NAND3X0_HVT U1901 ( .A1(n1718), .A2(n1834), .A3(n1717), .Y(
        n_sram_raddr_a2[7]) );
  NAND2X0_HVT U1902 ( .A1(n398), .A2(n1721), .Y(n1719) );
  NAND2X0_HVT U1903 ( .A1(n1720), .A2(n1719), .Y(n1733) );
  AND3X1_HVT U1904 ( .A1(sram_raddr_a2[7]), .A2(n1722), .A3(n1721), .Y(n1731)
         );
  NAND2X0_HVT U1905 ( .A1(n1724), .A2(sram_raddr_a8[8]), .Y(n1727) );
  OA21X1_HVT U1906 ( .A1(n1724), .A2(sram_raddr_a8[8]), .A3(n1727), .Y(n1980)
         );
  NAND2X0_HVT U1907 ( .A1(sram_raddr_a5[8]), .A2(n1725), .Y(n1729) );
  OA21X1_HVT U1908 ( .A1(sram_raddr_a5[8]), .A2(n1725), .A3(n1729), .Y(n1839)
         );
  AO22X1_HVT U1909 ( .A1(n519), .A2(n1980), .A3(n1974), .A4(n1839), .Y(n1726)
         );
  AO221X1_HVT U1910 ( .A1(sram_raddr_a2[8]), .A2(n1733), .A3(n449), .A4(n1731), 
        .A5(n1726), .Y(n_sram_raddr_a2[8]) );
  HADDX1_HVT U1911 ( .A0(sram_raddr_a8[9]), .B0(n1728), .SO(n1988) );
  AND2X1_HVT U1912 ( .A1(n519), .A2(n1988), .Y(n1846) );
  HADDX1_HVT U1913 ( .A0(sram_raddr_a5[9]), .B0(n1730), .SO(n1844) );
  HADDX1_HVT U1914 ( .A0(sram_raddr_a2[9]), .B0(sram_raddr_a2[8]), .SO(n1732)
         );
  NAND2X0_HVT U1915 ( .A1(n189), .A2(n1849), .Y(n1769) );
  AO22X1_HVT U1916 ( .A1(n519), .A2(n306), .A3(n1896), .A4(sram_raddr_a0[0]), 
        .Y(n1734) );
  AO221X1_HVT U1917 ( .A1(sram_raddr_a3[0]), .A2(n1887), .A3(n433), .A4(n1769), 
        .A5(n1734), .Y(n_sram_raddr_a3[0]) );
  OA21X1_HVT U1918 ( .A1(n422), .A2(n218), .A3(n1735), .Y(n1848) );
  AOI22X1_HVT U1919 ( .A1(n1736), .A2(n1769), .A3(sram_raddr_a3[1]), .A4(n1887), .Y(n1737) );
  NAND2X0_HVT U1920 ( .A1(n1848), .A2(n1737), .Y(n_sram_raddr_a3[1]) );
  OA22X1_HVT U1921 ( .A1(n1759), .A2(n244), .A3(n1758), .A4(n1739), .Y(n1741)
         );
  AO221X1_HVT U1922 ( .A1(sram_raddr_a0[3]), .A2(n248), .A3(n239), .A4(
        sram_raddr_a0[2]), .A5(n218), .Y(n1854) );
  NAND3X0_HVT U1923 ( .A1(n1741), .A2(n1740), .A3(n1854), .Y(
        n_sram_raddr_a3[3]) );
  NAND3X0_HVT U1924 ( .A1(n342), .A2(n239), .A3(n248), .Y(n1748) );
  NAND2X0_HVT U1925 ( .A1(n239), .A2(n248), .Y(n1742) );
  NAND2X0_HVT U1926 ( .A1(sram_raddr_a0[4]), .A2(n1742), .Y(n1744) );
  OA221X1_HVT U1927 ( .A1(n172), .A2(n1748), .A3(n218), .A4(n1744), .A5(n1743), 
        .Y(n1861) );
  OA22X1_HVT U1928 ( .A1(n1759), .A2(n275), .A3(n1758), .A4(n1745), .Y(n1746)
         );
  NAND2X0_HVT U1929 ( .A1(n1861), .A2(n1746), .Y(n_sram_raddr_a3[4]) );
  AOI22X1_HVT U1930 ( .A1(n1747), .A2(n1769), .A3(sram_raddr_a3[5]), .A4(n1887), .Y(n1751) );
  AO221X1_HVT U1931 ( .A1(sram_raddr_a0[5]), .A2(n1749), .A3(n284), .A4(n1748), 
        .A5(n172), .Y(n1865) );
  NAND3X0_HVT U1932 ( .A1(n1751), .A2(n1750), .A3(n1865), .Y(
        n_sram_raddr_a3[5]) );
  NAND4X0_HVT U1933 ( .A1(n284), .A2(n342), .A3(n239), .A4(n248), .Y(n1752) );
  OR2X1_HVT U1934 ( .A1(n1752), .A2(sram_raddr_a0[6]), .Y(n1760) );
  NAND2X0_HVT U1935 ( .A1(sram_raddr_a0[6]), .A2(n1752), .Y(n1754) );
  OA221X1_HVT U1936 ( .A1(n172), .A2(n1760), .A3(n218), .A4(n1754), .A5(n1753), 
        .Y(n1872) );
  OA22X1_HVT U1937 ( .A1(n1759), .A2(n331), .A3(n1758), .A4(n1755), .Y(n1756)
         );
  NAND2X0_HVT U1938 ( .A1(n1872), .A2(n1756), .Y(n_sram_raddr_a3[6]) );
  OA22X1_HVT U1939 ( .A1(n1759), .A2(n412), .A3(n1758), .A4(n1757), .Y(n1763)
         );
  NAND2X0_HVT U1940 ( .A1(n1761), .A2(n397), .Y(n1764) );
  AO221X1_HVT U1941 ( .A1(n1764), .A2(n1761), .A3(n1764), .A4(n397), .A5(n172), 
        .Y(n1877) );
  NAND3X0_HVT U1942 ( .A1(n1763), .A2(n1762), .A3(n1877), .Y(
        n_sram_raddr_a3[7]) );
  OA221X1_HVT U1943 ( .A1(sram_raddr_a0[8]), .A2(n1766), .A3(n424), .A4(n1764), 
        .A5(n1896), .Y(n1883) );
  NAND2X0_HVT U1944 ( .A1(n1766), .A2(n424), .Y(n1767) );
  OA221X1_HVT U1945 ( .A1(sram_raddr_a0[9]), .A2(n1768), .A3(n457), .A4(n1767), 
        .A5(n1896), .Y(n1889) );
  AO22X1_HVT U1946 ( .A1(n1770), .A2(n1769), .A3(sram_raddr_a3[9]), .A4(n1887), 
        .Y(n1771) );
  OR3X1_HVT U1947 ( .A1(n1772), .A2(n1889), .A3(n1771), .Y(n_sram_raddr_a3[9])
         );
  NAND2X0_HVT U1948 ( .A1(n1913), .A2(n171), .Y(n1803) );
  AO22X1_HVT U1949 ( .A1(n1838), .A2(n303), .A3(n1896), .A4(sram_raddr_a1[0]), 
        .Y(n1773) );
  AO221X1_HVT U1950 ( .A1(sram_raddr_a4[0]), .A2(n1934), .A3(n417), .A4(n1803), 
        .A5(n1773), .Y(n_sram_raddr_a4[0]) );
  OA22X1_HVT U1951 ( .A1(n1794), .A2(n1774), .A3(n1892), .A4(n307), .Y(n1776)
         );
  NAND2X0_HVT U1952 ( .A1(n1896), .A2(sram_raddr_a1[1]), .Y(n1893) );
  NAND3X0_HVT U1953 ( .A1(n1776), .A2(n1775), .A3(n1893), .Y(
        n_sram_raddr_a4[1]) );
  AOI22X1_HVT U1954 ( .A1(n1778), .A2(n1803), .A3(sram_raddr_a4[3]), .A4(n1934), .Y(n1780) );
  AO221X1_HVT U1955 ( .A1(sram_raddr_a1[2]), .A2(n238), .A3(n247), .A4(
        sram_raddr_a1[3]), .A5(n172), .Y(n1900) );
  NAND3X0_HVT U1956 ( .A1(n1780), .A2(n1779), .A3(n1900), .Y(
        n_sram_raddr_a4[3]) );
  OA22X1_HVT U1957 ( .A1(n1892), .A2(n246), .A3(n1794), .A4(n1781), .Y(n1785)
         );
  NAND2X0_HVT U1958 ( .A1(n247), .A2(n238), .Y(n1782) );
  AO221X1_HVT U1959 ( .A1(sram_raddr_a1[4]), .A2(n1783), .A3(n278), .A4(n1782), 
        .A5(n218), .Y(n1906) );
  NAND3X0_HVT U1960 ( .A1(n1785), .A2(n1784), .A3(n1906), .Y(
        n_sram_raddr_a4[4]) );
  OA22X1_HVT U1961 ( .A1(n1892), .A2(n356), .A3(n1794), .A4(n1786), .Y(n1789)
         );
  NAND4X0_HVT U1962 ( .A1(n345), .A2(n278), .A3(n247), .A4(n238), .Y(n1790) );
  AND3X1_HVT U1963 ( .A1(n278), .A2(n247), .A3(n238), .Y(n1787) );
  AO221X1_HVT U1964 ( .A1(n1790), .A2(n1787), .A3(n1790), .A4(n345), .A5(n172), 
        .Y(n1911) );
  NAND3X0_HVT U1965 ( .A1(n1789), .A2(n1788), .A3(n1911), .Y(
        n_sram_raddr_a4[5]) );
  OR2X1_HVT U1966 ( .A1(n1790), .A2(sram_raddr_a1[6]), .Y(n1796) );
  NAND2X0_HVT U1967 ( .A1(sram_raddr_a1[6]), .A2(n1790), .Y(n1792) );
  OA221X1_HVT U1968 ( .A1(n218), .A2(n1796), .A3(n218), .A4(n1792), .A5(n1791), 
        .Y(n1919) );
  OA22X1_HVT U1969 ( .A1(n1892), .A2(n333), .A3(n1794), .A4(n1793), .Y(n1795)
         );
  NAND2X0_HVT U1970 ( .A1(n1919), .A2(n1795), .Y(n_sram_raddr_a4[6]) );
  OR2X1_HVT U1971 ( .A1(n1796), .A2(sram_raddr_a1[7]), .Y(n1798) );
  OA221X1_HVT U1972 ( .A1(n1800), .A2(sram_raddr_a1[7]), .A3(n1800), .A4(n1796), .A5(n1896), .Y(n1923) );
  OA221X1_HVT U1973 ( .A1(sram_raddr_a1[8]), .A2(n1800), .A3(n425), .A4(n1798), 
        .A5(n1896), .Y(n1928) );
  NAND2X0_HVT U1974 ( .A1(n1800), .A2(n425), .Y(n1801) );
  OA221X1_HVT U1975 ( .A1(sram_raddr_a1[9]), .A2(n1802), .A3(n458), .A4(n1801), 
        .A5(n1896), .Y(n1935) );
  AO22X1_HVT U1976 ( .A1(n1804), .A2(n1803), .A3(sram_raddr_a4[9]), .A4(n1934), 
        .Y(n1805) );
  OR3X1_HVT U1977 ( .A1(n1806), .A2(n1935), .A3(n1805), .Y(n_sram_raddr_a4[9])
         );
  NAND2X0_HVT U1978 ( .A1(n171), .A2(n1941), .Y(n1843) );
  AO22X1_HVT U1979 ( .A1(n519), .A2(n302), .A3(n1896), .A4(n442), .Y(n1936) );
  AO221X1_HVT U1980 ( .A1(sram_raddr_a5[0]), .A2(n1989), .A3(n416), .A4(n1843), 
        .A5(n1936), .Y(n_sram_raddr_a5[0]) );
  AO22X1_HVT U1981 ( .A1(n1981), .A2(n1807), .A3(sram_raddr_a5[1]), .A4(n1989), 
        .Y(n1808) );
  OR2X1_HVT U1982 ( .A1(n1940), .A2(n1808), .Y(n_sram_raddr_a5[1]) );
  OA22X1_HVT U1983 ( .A1(n1945), .A2(n360), .A3(n1941), .A4(n1946), .Y(n1810)
         );
  NAND2X0_HVT U1984 ( .A1(n1896), .A2(n1809), .Y(n1948) );
  NAND3X0_HVT U1985 ( .A1(n1811), .A2(n1810), .A3(n1948), .Y(
        n_sram_raddr_a5[2]) );
  OA22X1_HVT U1986 ( .A1(n1830), .A2(n1812), .A3(n1945), .A4(n274), .Y(n1815)
         );
  NAND2X0_HVT U1987 ( .A1(n1813), .A2(n343), .Y(n1817) );
  AO221X1_HVT U1988 ( .A1(n1817), .A2(n1813), .A3(n1817), .A4(n343), .A5(n172), 
        .Y(n1953) );
  NAND3X0_HVT U1989 ( .A1(n1815), .A2(n1814), .A3(n1953), .Y(
        n_sram_raddr_a5[3]) );
  OA22X1_HVT U1990 ( .A1(n1945), .A2(n361), .A3(n1830), .A4(n1816), .Y(n1819)
         );
  AO221X1_HVT U1991 ( .A1(sram_raddr_a2[4]), .A2(n1821), .A3(n341), .A4(n1817), 
        .A5(n218), .Y(n1959) );
  NAND3X0_HVT U1992 ( .A1(n1819), .A2(n1818), .A3(n1959), .Y(
        n_sram_raddr_a5[4]) );
  OA22X1_HVT U1993 ( .A1(n1945), .A2(n332), .A3(n1830), .A4(n1820), .Y(n1824)
         );
  AND2X1_HVT U1994 ( .A1(n1821), .A2(n341), .Y(n1822) );
  NAND2X0_HVT U1995 ( .A1(n1822), .A2(n348), .Y(n1826) );
  AO221X1_HVT U1996 ( .A1(n1826), .A2(n1822), .A3(n1826), .A4(n348), .A5(n218), 
        .Y(n1964) );
  NAND3X0_HVT U1997 ( .A1(n1824), .A2(n1823), .A3(n1964), .Y(
        n_sram_raddr_a5[5]) );
  OA22X1_HVT U1998 ( .A1(n1945), .A2(n362), .A3(n1830), .A4(n1825), .Y(n1828)
         );
  AO221X1_HVT U1999 ( .A1(sram_raddr_a2[6]), .A2(n1831), .A3(n410), .A4(n1826), 
        .A5(n172), .Y(n1970) );
  NAND3X0_HVT U2000 ( .A1(n1828), .A2(n1827), .A3(n1970), .Y(
        n_sram_raddr_a5[6]) );
  OA22X1_HVT U2001 ( .A1(n1945), .A2(n396), .A3(n1830), .A4(n1829), .Y(n1835)
         );
  AND2X1_HVT U2002 ( .A1(n1831), .A2(n410), .Y(n1833) );
  NAND2X0_HVT U2003 ( .A1(n1833), .A2(n398), .Y(n1836) );
  AO221X1_HVT U2004 ( .A1(n1836), .A2(n1833), .A3(n1836), .A4(n398), .A5(n172), 
        .Y(n1977) );
  NAND3X0_HVT U2005 ( .A1(n1835), .A2(n1834), .A3(n1977), .Y(
        n_sram_raddr_a5[7]) );
  OR2X1_HVT U2006 ( .A1(n1836), .A2(sram_raddr_a2[8]), .Y(n1841) );
  AO21X1_HVT U2007 ( .A1(sram_raddr_a2[8]), .A2(n1836), .A3(n1842), .Y(n1837)
         );
  AO22X1_HVT U2008 ( .A1(n519), .A2(n1980), .A3(n1896), .A4(n1837), .Y(n1983)
         );
  AO22X1_HVT U2009 ( .A1(n1839), .A2(n1843), .A3(sram_raddr_a5[8]), .A4(n1989), 
        .Y(n1840) );
  OR2X1_HVT U2010 ( .A1(n1983), .A2(n1840), .Y(n_sram_raddr_a5[8]) );
  OA221X1_HVT U2011 ( .A1(sram_raddr_a2[9]), .A2(n1842), .A3(n459), .A4(n1841), 
        .A5(n1896), .Y(n1992) );
  AO22X1_HVT U2012 ( .A1(n1844), .A2(n1843), .A3(sram_raddr_a5[9]), .A4(n1989), 
        .Y(n1845) );
  OR3X1_HVT U2013 ( .A1(n1846), .A2(n1992), .A3(n1845), .Y(n_sram_raddr_a5[9])
         );
  NAND2X0_HVT U2014 ( .A1(n1942), .A2(n1849), .Y(n1885) );
  AO22X1_HVT U2015 ( .A1(n1896), .A2(sram_raddr_a0[0]), .A3(n1974), .A4(
        sram_raddr_a3[0]), .Y(n1847) );
  AO221X1_HVT U2016 ( .A1(sram_raddr_a6[0]), .A2(n1887), .A3(n306), .A4(n1885), 
        .A5(n1847), .Y(n_sram_raddr_a6[0]) );
  AOI22X1_HVT U2017 ( .A1(sram_raddr_a6[3]), .A2(n1887), .A3(n1852), .A4(n1885), .Y(n1855) );
  AO221X1_HVT U2018 ( .A1(sram_raddr_a3[2]), .A2(n244), .A3(n236), .A4(
        sram_raddr_a3[3]), .A5(n189), .Y(n1853) );
  NAND3X0_HVT U2019 ( .A1(n1855), .A2(n1854), .A3(n1853), .Y(
        n_sram_raddr_a6[3]) );
  AOI22X1_HVT U2020 ( .A1(sram_raddr_a6[4]), .A2(n1887), .A3(n1868), .A4(n1856), .Y(n1860) );
  NAND2X0_HVT U2021 ( .A1(n236), .A2(n244), .Y(n1857) );
  AO221X1_HVT U2022 ( .A1(sram_raddr_a3[4]), .A2(n1858), .A3(n275), .A4(n1857), 
        .A5(n189), .Y(n1859) );
  NAND3X0_HVT U2023 ( .A1(n1861), .A2(n1860), .A3(n1859), .Y(
        n_sram_raddr_a6[4]) );
  AOI22X1_HVT U2024 ( .A1(sram_raddr_a6[5]), .A2(n1887), .A3(n1862), .A4(n1885), .Y(n1866) );
  NAND4X0_HVT U2025 ( .A1(n363), .A2(n275), .A3(n236), .A4(n244), .Y(n1869) );
  AND3X1_HVT U2026 ( .A1(n275), .A2(n236), .A3(n244), .Y(n1863) );
  AO221X1_HVT U2027 ( .A1(n1869), .A2(n1863), .A3(n1869), .A4(n363), .A5(n171), 
        .Y(n1864) );
  NAND3X0_HVT U2028 ( .A1(n1866), .A2(n1865), .A3(n1864), .Y(
        n_sram_raddr_a6[5]) );
  AOI22X1_HVT U2029 ( .A1(sram_raddr_a6[6]), .A2(n1887), .A3(n1868), .A4(n1867), .Y(n1871) );
  AO221X1_HVT U2030 ( .A1(sram_raddr_a3[6]), .A2(n1874), .A3(n331), .A4(n1869), 
        .A5(n189), .Y(n1870) );
  NAND3X0_HVT U2031 ( .A1(n1872), .A2(n1871), .A3(n1870), .Y(
        n_sram_raddr_a6[6]) );
  AOI22X1_HVT U2032 ( .A1(sram_raddr_a6[7]), .A2(n1887), .A3(n1873), .A4(n1885), .Y(n1878) );
  AND2X1_HVT U2033 ( .A1(n1874), .A2(n331), .Y(n1875) );
  NAND2X0_HVT U2034 ( .A1(n1875), .A2(n412), .Y(n1879) );
  AO221X1_HVT U2035 ( .A1(n1879), .A2(n1875), .A3(n1879), .A4(n412), .A5(n189), 
        .Y(n1876) );
  NAND3X0_HVT U2036 ( .A1(n1878), .A2(n1877), .A3(n1876), .Y(
        n_sram_raddr_a6[7]) );
  OA221X1_HVT U2037 ( .A1(n1884), .A2(sram_raddr_a3[8]), .A3(n1884), .A4(n1879), .A5(n170), .Y(n1882) );
  AO22X1_HVT U2038 ( .A1(sram_raddr_a6[8]), .A2(n1887), .A3(n1880), .A4(n1885), 
        .Y(n1881) );
  OR3X1_HVT U2039 ( .A1(n1883), .A2(n1882), .A3(n1881), .Y(n_sram_raddr_a6[8])
         );
  HADDX1_HVT U2040 ( .A0(sram_raddr_a3[9]), .B0(n1884), .SO(n1888) );
  NAND2X0_HVT U2041 ( .A1(n1942), .A2(n1913), .Y(n1931) );
  AO22X1_HVT U2042 ( .A1(n1896), .A2(sram_raddr_a1[0]), .A3(n1974), .A4(
        sram_raddr_a4[0]), .Y(n1890) );
  AO221X1_HVT U2043 ( .A1(sram_raddr_a7[0]), .A2(n1934), .A3(n303), .A4(n1931), 
        .A5(n1890), .Y(n_sram_raddr_a7[0]) );
  NAND2X0_HVT U2044 ( .A1(n1891), .A2(n1931), .Y(n1895) );
  OA22X1_HVT U2045 ( .A1(n1892), .A2(n443), .A3(n171), .A4(n307), .Y(n1894) );
  NAND3X0_HVT U2046 ( .A1(n1895), .A2(n1894), .A3(n1893), .Y(
        n_sram_raddr_a7[1]) );
  AOI22X1_HVT U2047 ( .A1(sram_raddr_a7[3]), .A2(n1934), .A3(n1898), .A4(n1931), .Y(n1901) );
  AO221X1_HVT U2048 ( .A1(sram_raddr_a4[2]), .A2(n283), .A3(n237), .A4(
        sram_raddr_a4[3]), .A5(n171), .Y(n1899) );
  NAND3X0_HVT U2049 ( .A1(n1901), .A2(n1900), .A3(n1899), .Y(
        n_sram_raddr_a7[3]) );
  AOI22X1_HVT U2050 ( .A1(sram_raddr_a7[4]), .A2(n1934), .A3(n1902), .A4(n1931), .Y(n1907) );
  NAND2X0_HVT U2051 ( .A1(n237), .A2(n283), .Y(n1903) );
  AO221X1_HVT U2052 ( .A1(sram_raddr_a4[4]), .A2(n1904), .A3(n246), .A4(n1903), 
        .A5(n189), .Y(n1905) );
  NAND3X0_HVT U2053 ( .A1(n1907), .A2(n1906), .A3(n1905), .Y(
        n_sram_raddr_a7[4]) );
  AOI22X1_HVT U2054 ( .A1(sram_raddr_a7[5]), .A2(n1934), .A3(n1908), .A4(n1931), .Y(n1912) );
  NAND4X0_HVT U2055 ( .A1(n356), .A2(n246), .A3(n237), .A4(n283), .Y(n1916) );
  AND3X1_HVT U2056 ( .A1(n246), .A2(n237), .A3(n283), .Y(n1909) );
  AO221X1_HVT U2057 ( .A1(n1916), .A2(n1909), .A3(n1916), .A4(n356), .A5(n189), 
        .Y(n1910) );
  NAND3X0_HVT U2058 ( .A1(n1912), .A2(n1911), .A3(n1910), .Y(
        n_sram_raddr_a7[5]) );
  AOI22X1_HVT U2059 ( .A1(sram_raddr_a7[6]), .A2(n1934), .A3(n1915), .A4(n1914), .Y(n1918) );
  AO221X1_HVT U2060 ( .A1(sram_raddr_a4[6]), .A2(n1920), .A3(n333), .A4(n1916), 
        .A5(n171), .Y(n1917) );
  NAND3X0_HVT U2061 ( .A1(n1919), .A2(n1918), .A3(n1917), .Y(
        n_sram_raddr_a7[6]) );
  NAND2X0_HVT U2062 ( .A1(n1920), .A2(n333), .Y(n1921) );
  OR2X1_HVT U2063 ( .A1(n1921), .A2(sram_raddr_a4[7]), .Y(n1924) );
  OA221X1_HVT U2064 ( .A1(n1929), .A2(sram_raddr_a4[8]), .A3(n1929), .A4(n1924), .A5(n170), .Y(n1927) );
  AO22X1_HVT U2065 ( .A1(sram_raddr_a7[8]), .A2(n1934), .A3(n1925), .A4(n1931), 
        .Y(n1926) );
  OR3X1_HVT U2066 ( .A1(n1928), .A2(n1927), .A3(n1926), .Y(n_sram_raddr_a7[8])
         );
  HADDX1_HVT U2067 ( .A0(sram_raddr_a4[9]), .B0(n1929), .SO(n1930) );
  AO221X1_HVT U2068 ( .A1(sram_raddr_a8[0]), .A2(n1989), .A3(n302), .A4(n1981), 
        .A5(n1936), .Y(n1937) );
  AO21X1_HVT U2069 ( .A1(n170), .A2(n416), .A3(n1937), .Y(n_sram_raddr_a8[0])
         );
  AO22X1_HVT U2070 ( .A1(sram_raddr_a8[1]), .A2(n1989), .A3(n1981), .A4(n1938), 
        .Y(n1939) );
  OR2X1_HVT U2071 ( .A1(n1940), .A2(n1939), .Y(n_sram_raddr_a8[1]) );
  NAND2X0_HVT U2072 ( .A1(n1942), .A2(n1941), .Y(n1987) );
  OA22X1_HVT U2073 ( .A1(n1945), .A2(n452), .A3(n1944), .A4(n1943), .Y(n1949)
         );
  NAND2X0_HVT U2074 ( .A1(n170), .A2(n1946), .Y(n1947) );
  NAND3X0_HVT U2075 ( .A1(n1949), .A2(n1948), .A3(n1947), .Y(
        n_sram_raddr_a8[2]) );
  AOI22X1_HVT U2076 ( .A1(sram_raddr_a8[3]), .A2(n1989), .A3(n1950), .A4(n1987), .Y(n1954) );
  AO221X1_HVT U2077 ( .A1(sram_raddr_a5[3]), .A2(n1956), .A3(n274), .A4(n1951), 
        .A5(n171), .Y(n1952) );
  NAND3X0_HVT U2078 ( .A1(n1954), .A2(n1953), .A3(n1952), .Y(
        n_sram_raddr_a8[3]) );
  AOI22X1_HVT U2079 ( .A1(sram_raddr_a8[4]), .A2(n1989), .A3(n1955), .A4(n1987), .Y(n1960) );
  AND2X1_HVT U2080 ( .A1(n1956), .A2(n274), .Y(n1957) );
  NAND2X0_HVT U2081 ( .A1(n1957), .A2(n361), .Y(n1962) );
  AO221X1_HVT U2082 ( .A1(n1962), .A2(n1957), .A3(n1962), .A4(n361), .A5(n171), 
        .Y(n1958) );
  NAND3X0_HVT U2083 ( .A1(n1960), .A2(n1959), .A3(n1958), .Y(
        n_sram_raddr_a8[4]) );
  AOI22X1_HVT U2084 ( .A1(sram_raddr_a8[5]), .A2(n1989), .A3(n1961), .A4(n1987), .Y(n1965) );
  AO221X1_HVT U2085 ( .A1(sram_raddr_a5[5]), .A2(n1967), .A3(n332), .A4(n1962), 
        .A5(n171), .Y(n1963) );
  NAND3X0_HVT U2086 ( .A1(n1965), .A2(n1964), .A3(n1963), .Y(
        n_sram_raddr_a8[5]) );
  AOI22X1_HVT U2087 ( .A1(sram_raddr_a8[6]), .A2(n1989), .A3(n1966), .A4(n1987), .Y(n1971) );
  AND2X1_HVT U2088 ( .A1(n1967), .A2(n332), .Y(n1968) );
  NAND2X0_HVT U2089 ( .A1(n1968), .A2(n362), .Y(n1973) );
  AO221X1_HVT U2090 ( .A1(n1973), .A2(n1968), .A3(n1973), .A4(n362), .A5(n189), 
        .Y(n1969) );
  NAND3X0_HVT U2091 ( .A1(n1971), .A2(n1970), .A3(n1969), .Y(
        n_sram_raddr_a8[6]) );
  AOI22X1_HVT U2092 ( .A1(sram_raddr_a8[7]), .A2(n1989), .A3(n1972), .A4(n1987), .Y(n1978) );
  NAND2X0_HVT U2093 ( .A1(n1975), .A2(n396), .Y(n1979) );
  AO221X1_HVT U2094 ( .A1(n1979), .A2(n1975), .A3(n1979), .A4(n396), .A5(n171), 
        .Y(n1976) );
  NAND3X0_HVT U2095 ( .A1(n1978), .A2(n1977), .A3(n1976), .Y(
        n_sram_raddr_a8[7]) );
  OR2X1_HVT U2096 ( .A1(n1979), .A2(sram_raddr_a5[8]), .Y(n1985) );
  OA221X1_HVT U2097 ( .A1(n1986), .A2(sram_raddr_a5[8]), .A3(n1986), .A4(n1979), .A5(n170), .Y(n1984) );
  AO22X1_HVT U2098 ( .A1(sram_raddr_a8[8]), .A2(n1989), .A3(n1981), .A4(n1980), 
        .Y(n1982) );
  OR3X1_HVT U2099 ( .A1(n1984), .A2(n1983), .A3(n1982), .Y(n_sram_raddr_a8[8])
         );
  OA221X1_HVT U2100 ( .A1(sram_raddr_a5[9]), .A2(n1986), .A3(n455), .A4(n1985), 
        .A5(n170), .Y(n1991) );
  AO22X1_HVT U2101 ( .A1(sram_raddr_a8[9]), .A2(n1989), .A3(n1988), .A4(n1987), 
        .Y(n1990) );
  OR3X1_HVT U2102 ( .A1(n1992), .A2(n1991), .A3(n1990), .Y(n_sram_raddr_a8[9])
         );
  AND2X1_HVT U2103 ( .A1(n1993), .A2(addr_row_sel_cnt[1]), .Y(n392) );
  OA221X1_HVT U2104 ( .A1(n2003), .A2(n1994), .A3(n2003), .A4(n2001), .A5(
        n1999), .Y(n371) );
  AO22X1_HVT U2105 ( .A1(n1998), .A2(n1997), .A3(n1996), .A4(n2001), .Y(n369)
         );
  OA221X1_HVT U2106 ( .A1(n2003), .A2(n2002), .A3(n2003), .A4(n2001), .A5(
        n2000), .Y(n368) );
endmodule


module data_reg ( clk, srstn, mode, box_sel, sram_rdata_a0, sram_rdata_a1, 
        sram_rdata_a2, sram_rdata_a3, sram_rdata_a4, sram_rdata_a5, 
        sram_rdata_a6, sram_rdata_a7, sram_rdata_a8, sram_rdata_b0, 
        sram_rdata_b1, sram_rdata_b2, sram_rdata_b3, sram_rdata_b4, 
        sram_rdata_b5, sram_rdata_b6, sram_rdata_b7, sram_rdata_b8, 
        sram_rdata_weight, conv1_weight, weight, src_window );
  input [1:0] mode;
  input [3:0] box_sel;
  input [31:0] sram_rdata_a0;
  input [31:0] sram_rdata_a1;
  input [31:0] sram_rdata_a2;
  input [31:0] sram_rdata_a3;
  input [31:0] sram_rdata_a4;
  input [31:0] sram_rdata_a5;
  input [31:0] sram_rdata_a6;
  input [31:0] sram_rdata_a7;
  input [31:0] sram_rdata_a8;
  input [31:0] sram_rdata_b0;
  input [31:0] sram_rdata_b1;
  input [31:0] sram_rdata_b2;
  input [31:0] sram_rdata_b3;
  input [31:0] sram_rdata_b4;
  input [31:0] sram_rdata_b5;
  input [31:0] sram_rdata_b6;
  input [31:0] sram_rdata_b7;
  input [31:0] sram_rdata_b8;
  input [99:0] sram_rdata_weight;
  output [99:0] conv1_weight;
  output [99:0] weight;
  output [287:0] src_window;
  input clk, srstn;
  wire   N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52,
         N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66,
         N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80,
         N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94,
         N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139,
         N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161,
         N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172,
         N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183,
         N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194,
         N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205,
         N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216,
         N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227,
         N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238,
         N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249,
         N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260,
         N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271,
         N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282,
         N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293,
         N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304,
         N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315,
         N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326,
         N346, n2, n3, n5, n6, n8, n9, n11, n12, n14, n15, n17, n18, n20, n21,
         n23, n24, n26, n27, n29, n30, n32, n33, n35, n36, n38, n3900, n4100,
         n4200, n4400, n4500, n4700, n4800, n5000, n5100, n5300, n5400, n5600,
         n5700, n5900, n6000, n6200, n6300, n6500, n6600, n6800, n6900, n7100,
         n7200, n7400, n7500, n7700, n7800, n8000, n8100, n8300, n8400, n8600,
         n8700, n8900, n9000, n9200, n9300, n9400, n9500, n9700, n9800, n9900,
         n10000, n10100, n10200, n10300, n10400, n10500, n10600, n10700,
         n10800, n10900, n11000, n11100, n11200, n11300, n11400, n11500,
         n11600, n11700, n11800, n11900, n12000, n12100, n12200, n12300,
         n12400, n12500, n12600, n12700, n12800, n12900, n13000, n13100,
         n13200, n13300, n13400, n13500, n13600, n13700, n13800, n13900,
         n14000, n14100, n14200, n14300, n14400, n14500, n14600, n14700,
         n14800, n14900, n15000, n15100, n15200, n15300, n15400, n15500,
         n15600, n15700, n15800, n15900, n16000, n16100, n16200, n16300,
         n16400, n16500, n16600, n1670, n1680, n1690, n1700, n1710, n1720,
         n1730, n1740, n1750, n1760, n1770, n1780, n1790, n1800, n1810, n1820,
         n1830, n1840, n1850, n1860, n1870, n1880, n1890, n1900, n1910, n1920,
         n1930, n1940, n1950, n1960, n1970, n1980, n1990, n2000, n2010, n2020,
         n2030, n2040, n2050, n2060, n2070, n2080, n2090, n2100, n2110, n2120,
         n2130, n2140, n2150, n2160, n2170, n2180, n2190, n2200, n2210, n2220,
         n2230, n2240, n2250, n2260, n2270, n2280, n2290, n2300, n2310, n2320,
         n2330, n2340, n2350, n2360, n2370, n2380, n2390, n2400, n2410, n2420,
         n2430, n2440, n2450, n2460, n2470, n2480, n2490, n2500, n2510, n2520,
         n2530, n2540, n2550, n2560, n2570, n2580, n2590, n2600, n2610, n2620,
         n2630, n2640, n2650, n2660, n2670, n2680, n2690, n2700, n2710, n2720,
         n2730, n2740, n2750, n2760, n2770, n2780, n2790, n2800, n2810, n2820,
         n2830, n2840, n2850, n2860, n2870, n2880, n2890, n2900, n2910, n2920,
         n2930, n2940, n2950, n2960, n2970, n2980, n2990, n3000, n3010, n3020,
         n3030, n3040, n3050, n3060, n3070, n3080, n3090, n3100, n3110, n3120,
         n3130, n3140, n3150, n3160, n3170, n3180, n3190, n3200, n3210, n3220,
         n3230, n3240, n3250, n3260, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n3460, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n3901, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n4001, n401, n402, n403, n404, n405, n406, n407, n408, n409, n4101,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n4201, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n4301, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n4401, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n4501, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n4601, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n4701, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n4801, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n4901, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n5001, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n5101, n511, n512, n513, n514, n515, n516, n517, n518, n519, n5201,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n5301, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n5401, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n5501, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n5601, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n5701, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n5801, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n5901, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n6001, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n6101, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n6201, n621, n622, n623, n624, n625, n626, n627, n628, n629, n6301,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n6401, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n6501, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n6601, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n6701, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n6801, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n6901, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n7001, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n7101, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n7201, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n7301, n731, n732, n733, n734, n735, n736, n737, n738, n739, n7401,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n7501, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n7601, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n7701, n771, n772, n773,
         n774, n775, n777, n778, n779, n7801, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n7901, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n8001, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n8101, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n8201, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n8301, n831, n832, n833, n834, n835, n836, n837, n838, n839, n8401,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n8501, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n8601, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n8701, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n8801, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n8901, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n9001, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n9101, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n9201, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n9301, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n9401, n941, n942, n943, n944, n945, n946, n947, n948, n949, n9501,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n9601, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n9701, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n9801, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n9901, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n10001, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n10101, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n10201, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n10301, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n10401, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n10501, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n10601, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n10701, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n10801, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n10901, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n11001, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n11101, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n11201, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n11301, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n11401, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n11501, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n11601, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n11701, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n11801, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n11901, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n12001, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n12101, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n12201, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n12301, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n12401, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n12501, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n12601, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n12701, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n12801, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n12901, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n13001, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n13101, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n13201, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n13301, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n13401, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n13501, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n13601, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n13701, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n13801, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n13901, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n14001, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n14101, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n14201, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n14301, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n14401, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n14501, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n14601, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n14701, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n14801, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n14901, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n15001, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n15101, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n15201, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n15301, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n15401, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n15501, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n15601, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n15701, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n15801, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n15901, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n16001, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n16101, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n16201, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n16301, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n16401, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n16501, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n16601, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667;
  wire   [287:0] n_src_aox;
  wire   [31:0] sram_rdata_0;
  wire   [31:0] sram_rdata_1;
  wire   [31:0] sram_rdata_2;
  wire   [31:0] sram_rdata_3;
  wire   [31:0] sram_rdata_4;
  wire   [31:0] sram_rdata_5;
  wire   [31:0] sram_rdata_6;
  wire   [31:0] sram_rdata_7;
  wire   [31:0] sram_rdata_8;

  DFFSSRX1_HVT src_aox_reg_0__7_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[287]), .CLK(clk), .Q(src_window[287]) );
  DFFSSRX1_HVT src_aox_reg_0__6_ ( .D(1'b0), .SETB(n2560), .RSTB(
        n_src_aox[286]), .CLK(clk), .Q(src_window[286]) );
  DFFSSRX1_HVT src_aox_reg_0__5_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[285]), .CLK(clk), .Q(src_window[285]) );
  DFFSSRX1_HVT src_aox_reg_0__4_ ( .D(1'b0), .SETB(n579), .RSTB(n_src_aox[284]), .CLK(clk), .Q(src_window[284]) );
  DFFSSRX1_HVT src_aox_reg_0__3_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[283]), .CLK(clk), .Q(src_window[283]) );
  DFFSSRX1_HVT src_aox_reg_0__2_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[282]), .CLK(clk), .Q(src_window[282]) );
  DFFSSRX1_HVT src_aox_reg_0__1_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[281]), .CLK(clk), .Q(src_window[281]) );
  DFFSSRX1_HVT src_aox_reg_0__0_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[280]), .CLK(clk), .Q(src_window[280]) );
  DFFSSRX1_HVT src_aox_reg_1__7_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[279]), .CLK(clk), .Q(src_window[279]) );
  DFFSSRX1_HVT src_aox_reg_1__6_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[278]), .CLK(clk), .Q(src_window[278]) );
  DFFSSRX1_HVT src_aox_reg_1__5_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[277]), .CLK(clk), .Q(src_window[277]) );
  DFFSSRX1_HVT src_aox_reg_1__4_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[276]), .CLK(clk), .Q(src_window[276]) );
  DFFSSRX1_HVT src_aox_reg_1__3_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[275]), .CLK(clk), .Q(src_window[275]) );
  DFFSSRX1_HVT src_aox_reg_1__2_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[274]), .CLK(clk), .Q(src_window[274]) );
  DFFSSRX1_HVT src_aox_reg_1__1_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[273]), .CLK(clk), .Q(src_window[273]) );
  DFFSSRX1_HVT src_aox_reg_1__0_ ( .D(1'b0), .SETB(n579), .RSTB(n_src_aox[272]), .CLK(clk), .Q(src_window[272]) );
  DFFSSRX1_HVT src_aox_reg_2__7_ ( .D(1'b0), .SETB(N346), .RSTB(n_src_aox[271]), .CLK(clk), .Q(src_window[271]) );
  DFFSSRX1_HVT src_aox_reg_2__6_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[270]), .CLK(clk), .Q(src_window[270]) );
  DFFSSRX1_HVT src_aox_reg_2__5_ ( .D(1'b0), .SETB(n579), .RSTB(n_src_aox[269]), .CLK(clk), .Q(src_window[269]) );
  DFFSSRX1_HVT src_aox_reg_2__4_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[268]), .CLK(clk), .Q(src_window[268]) );
  DFFSSRX1_HVT src_aox_reg_2__3_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[267]), .CLK(clk), .Q(src_window[267]) );
  DFFSSRX1_HVT src_aox_reg_2__2_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[266]), .CLK(clk), .Q(src_window[266]) );
  DFFSSRX1_HVT src_aox_reg_2__1_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[265]), .CLK(clk), .Q(src_window[265]) );
  DFFSSRX1_HVT src_aox_reg_2__0_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[264]), .CLK(clk), .Q(src_window[264]) );
  DFFSSRX1_HVT src_aox_reg_3__7_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[263]), .CLK(clk), .Q(src_window[263]) );
  DFFSSRX1_HVT src_aox_reg_3__6_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[262]), .CLK(clk), .Q(src_window[262]) );
  DFFSSRX1_HVT src_aox_reg_3__5_ ( .D(1'b0), .SETB(N346), .RSTB(n_src_aox[261]), .CLK(clk), .Q(src_window[261]) );
  DFFSSRX1_HVT src_aox_reg_3__4_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[260]), .CLK(clk), .Q(src_window[260]) );
  DFFSSRX1_HVT src_aox_reg_3__3_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[259]), .CLK(clk), .Q(src_window[259]) );
  DFFSSRX1_HVT src_aox_reg_3__2_ ( .D(1'b0), .SETB(n13200), .RSTB(
        n_src_aox[258]), .CLK(clk), .Q(src_window[258]) );
  DFFSSRX1_HVT src_aox_reg_3__1_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[257]), .CLK(clk), .Q(src_window[257]) );
  DFFSSRX1_HVT src_aox_reg_3__0_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[256]), .CLK(clk), .Q(src_window[256]) );
  DFFSSRX1_HVT src_aox_reg_4__7_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[255]), .CLK(clk), .Q(src_window[255]) );
  DFFSSRX1_HVT src_aox_reg_4__6_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[254]), .CLK(clk), .Q(src_window[254]) );
  DFFSSRX1_HVT src_aox_reg_4__5_ ( .D(1'b0), .SETB(n13200), .RSTB(
        n_src_aox[253]), .CLK(clk), .Q(src_window[253]) );
  DFFSSRX1_HVT src_aox_reg_4__4_ ( .D(1'b0), .SETB(n579), .RSTB(n_src_aox[252]), .CLK(clk), .Q(src_window[252]) );
  DFFSSRX1_HVT src_aox_reg_4__3_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[251]), .CLK(clk), .Q(src_window[251]) );
  DFFSSRX1_HVT src_aox_reg_4__2_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[250]), .CLK(clk), .Q(src_window[250]) );
  DFFSSRX1_HVT src_aox_reg_4__1_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[249]), .CLK(clk), .Q(src_window[249]) );
  DFFSSRX1_HVT src_aox_reg_4__0_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[248]), .CLK(clk), .Q(src_window[248]) );
  DFFSSRX1_HVT src_aox_reg_5__7_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[247]), .CLK(clk), .Q(src_window[247]) );
  DFFSSRX1_HVT src_aox_reg_5__6_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[246]), .CLK(clk), .Q(src_window[246]) );
  DFFSSRX1_HVT src_aox_reg_5__5_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[245]), .CLK(clk), .Q(src_window[245]) );
  DFFSSRX1_HVT src_aox_reg_5__4_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[244]), .CLK(clk), .Q(src_window[244]) );
  DFFSSRX1_HVT src_aox_reg_5__3_ ( .D(1'b0), .SETB(n2560), .RSTB(
        n_src_aox[243]), .CLK(clk), .Q(src_window[243]) );
  DFFSSRX1_HVT src_aox_reg_5__2_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[242]), .CLK(clk), .Q(src_window[242]) );
  DFFSSRX1_HVT src_aox_reg_5__1_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[241]), .CLK(clk), .Q(src_window[241]) );
  DFFSSRX1_HVT src_aox_reg_5__0_ ( .D(1'b0), .SETB(n579), .RSTB(n_src_aox[240]), .CLK(clk), .Q(src_window[240]) );
  DFFSSRX1_HVT src_aox_reg_6__7_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[239]), .CLK(clk), .Q(src_window[239]) );
  DFFSSRX1_HVT src_aox_reg_6__6_ ( .D(1'b0), .SETB(n2560), .RSTB(
        n_src_aox[238]), .CLK(clk), .Q(src_window[238]) );
  DFFSSRX1_HVT src_aox_reg_6__5_ ( .D(1'b0), .SETB(n579), .RSTB(n_src_aox[237]), .CLK(clk), .Q(src_window[237]) );
  DFFSSRX1_HVT src_aox_reg_6__4_ ( .D(1'b0), .SETB(n13200), .RSTB(
        n_src_aox[236]), .CLK(clk), .Q(src_window[236]) );
  DFFSSRX1_HVT src_aox_reg_6__3_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[235]), .CLK(clk), .Q(src_window[235]) );
  DFFSSRX1_HVT src_aox_reg_6__2_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[234]), .CLK(clk), .Q(src_window[234]) );
  DFFSSRX1_HVT src_aox_reg_6__1_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[233]), .CLK(clk), .Q(src_window[233]) );
  DFFSSRX1_HVT src_aox_reg_6__0_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[232]), .CLK(clk), .Q(src_window[232]) );
  DFFSSRX1_HVT src_aox_reg_7__7_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[231]), .CLK(clk), .Q(src_window[231]) );
  DFFSSRX1_HVT src_aox_reg_7__6_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[230]), .CLK(clk), .Q(src_window[230]) );
  DFFSSRX1_HVT src_aox_reg_7__5_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[229]), .CLK(clk), .Q(src_window[229]) );
  DFFSSRX1_HVT src_aox_reg_7__4_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[228]), .CLK(clk), .Q(src_window[228]) );
  DFFSSRX1_HVT src_aox_reg_7__3_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[227]), .CLK(clk), .Q(src_window[227]) );
  DFFSSRX1_HVT src_aox_reg_7__2_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[226]), .CLK(clk), .Q(src_window[226]) );
  DFFSSRX1_HVT src_aox_reg_7__1_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[225]), .CLK(clk), .Q(src_window[225]) );
  DFFSSRX1_HVT src_aox_reg_7__0_ ( .D(1'b0), .SETB(n13200), .RSTB(
        n_src_aox[224]), .CLK(clk), .Q(src_window[224]) );
  DFFSSRX1_HVT src_aox_reg_8__7_ ( .D(1'b0), .SETB(n13200), .RSTB(
        n_src_aox[223]), .CLK(clk), .Q(src_window[223]) );
  DFFSSRX1_HVT src_aox_reg_8__6_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[222]), .CLK(clk), .Q(src_window[222]) );
  DFFSSRX1_HVT src_aox_reg_8__5_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[221]), .CLK(clk), .Q(src_window[221]) );
  DFFSSRX1_HVT src_aox_reg_8__4_ ( .D(1'b0), .SETB(n579), .RSTB(n_src_aox[220]), .CLK(clk), .Q(src_window[220]) );
  DFFSSRX1_HVT src_aox_reg_8__3_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[219]), .CLK(clk), .Q(src_window[219]) );
  DFFSSRX1_HVT src_aox_reg_8__2_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[218]), .CLK(clk), .Q(src_window[218]) );
  DFFSSRX1_HVT src_aox_reg_8__1_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[217]), .CLK(clk), .Q(src_window[217]) );
  DFFSSRX1_HVT src_aox_reg_8__0_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[216]), .CLK(clk), .Q(src_window[216]) );
  DFFSSRX1_HVT src_aox_reg_9__7_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[215]), .CLK(clk), .Q(src_window[215]) );
  DFFSSRX1_HVT src_aox_reg_9__6_ ( .D(1'b0), .SETB(n13200), .RSTB(
        n_src_aox[214]), .CLK(clk), .Q(src_window[214]) );
  DFFSSRX1_HVT src_aox_reg_9__5_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[213]), .CLK(clk), .Q(src_window[213]) );
  DFFSSRX1_HVT src_aox_reg_9__4_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[212]), .CLK(clk), .Q(src_window[212]) );
  DFFSSRX1_HVT src_aox_reg_9__3_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[211]), .CLK(clk), .Q(src_window[211]) );
  DFFSSRX1_HVT src_aox_reg_9__2_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[210]), .CLK(clk), .Q(src_window[210]) );
  DFFSSRX1_HVT src_aox_reg_9__1_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[209]), .CLK(clk), .Q(src_window[209]) );
  DFFSSRX1_HVT src_aox_reg_9__0_ ( .D(1'b0), .SETB(n579), .RSTB(n_src_aox[208]), .CLK(clk), .Q(src_window[208]) );
  DFFSSRX1_HVT src_aox_reg_10__7_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[207]), .CLK(clk), .Q(src_window[207]) );
  DFFSSRX1_HVT src_aox_reg_10__6_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[206]), .CLK(clk), .Q(src_window[206]) );
  DFFSSRX1_HVT src_aox_reg_10__5_ ( .D(1'b0), .SETB(n579), .RSTB(
        n_src_aox[205]), .CLK(clk), .Q(src_window[205]) );
  DFFSSRX1_HVT src_aox_reg_10__4_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[204]), .CLK(clk), .Q(src_window[204]) );
  DFFSSRX1_HVT src_aox_reg_10__3_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[203]), .CLK(clk), .Q(src_window[203]) );
  DFFSSRX1_HVT src_aox_reg_10__2_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[202]), .CLK(clk), .Q(src_window[202]) );
  DFFSSRX1_HVT src_aox_reg_10__1_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[201]), .CLK(clk), .Q(src_window[201]) );
  DFFSSRX1_HVT src_aox_reg_10__0_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[200]), .CLK(clk), .Q(src_window[200]) );
  DFFSSRX1_HVT src_aox_reg_11__7_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[199]), .CLK(clk), .Q(src_window[199]) );
  DFFSSRX1_HVT src_aox_reg_11__6_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[198]), .CLK(clk), .Q(src_window[198]) );
  DFFSSRX1_HVT src_aox_reg_11__5_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[197]), .CLK(clk), .Q(src_window[197]) );
  DFFSSRX1_HVT src_aox_reg_11__4_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[196]), .CLK(clk), .Q(src_window[196]) );
  DFFSSRX1_HVT src_aox_reg_11__3_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[195]), .CLK(clk), .Q(src_window[195]) );
  DFFSSRX1_HVT src_aox_reg_11__2_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[194]), .CLK(clk), .Q(src_window[194]) );
  DFFSSRX1_HVT src_aox_reg_11__1_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[193]), .CLK(clk), .Q(src_window[193]) );
  DFFSSRX1_HVT src_aox_reg_11__0_ ( .D(1'b0), .SETB(n2560), .RSTB(
        n_src_aox[192]), .CLK(clk), .Q(src_window[192]) );
  DFFSSRX1_HVT src_aox_reg_12__7_ ( .D(1'b0), .SETB(N346), .RSTB(
        n_src_aox[191]), .CLK(clk), .Q(src_window[191]) );
  DFFSSRX1_HVT src_aox_reg_12__6_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[190]), .CLK(clk), .Q(src_window[190]) );
  DFFSSRX1_HVT src_aox_reg_12__5_ ( .D(1'b0), .SETB(n2560), .RSTB(
        n_src_aox[189]), .CLK(clk), .Q(src_window[189]) );
  DFFSSRX1_HVT src_aox_reg_12__4_ ( .D(1'b0), .SETB(n579), .RSTB(
        n_src_aox[188]), .CLK(clk), .Q(src_window[188]) );
  DFFSSRX1_HVT src_aox_reg_12__3_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[187]), .CLK(clk), .Q(src_window[187]) );
  DFFSSRX1_HVT src_aox_reg_12__2_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[186]), .CLK(clk), .Q(src_window[186]) );
  DFFSSRX1_HVT src_aox_reg_12__1_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[185]), .CLK(clk), .Q(src_window[185]) );
  DFFSSRX1_HVT src_aox_reg_12__0_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[184]), .CLK(clk), .Q(src_window[184]) );
  DFFSSRX1_HVT src_aox_reg_13__7_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[183]), .CLK(clk), .Q(src_window[183]) );
  DFFSSRX1_HVT src_aox_reg_13__6_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[182]), .CLK(clk), .Q(src_window[182]) );
  DFFSSRX1_HVT src_aox_reg_13__5_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[181]), .CLK(clk), .Q(src_window[181]) );
  DFFSSRX1_HVT src_aox_reg_13__4_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[180]), .CLK(clk), .Q(src_window[180]) );
  DFFSSRX1_HVT src_aox_reg_13__3_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[179]), .CLK(clk), .Q(src_window[179]) );
  DFFSSRX1_HVT src_aox_reg_13__2_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[178]), .CLK(clk), .Q(src_window[178]) );
  DFFSSRX1_HVT src_aox_reg_13__1_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[177]), .CLK(clk), .Q(src_window[177]) );
  DFFSSRX1_HVT src_aox_reg_13__0_ ( .D(1'b0), .SETB(n579), .RSTB(
        n_src_aox[176]), .CLK(clk), .Q(src_window[176]) );
  DFFSSRX1_HVT src_aox_reg_14__7_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[175]), .CLK(clk), .Q(src_window[175]) );
  DFFSSRX1_HVT src_aox_reg_14__6_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[174]), .CLK(clk), .Q(src_window[174]) );
  DFFSSRX1_HVT src_aox_reg_14__5_ ( .D(1'b0), .SETB(n579), .RSTB(
        n_src_aox[173]), .CLK(clk), .Q(src_window[173]) );
  DFFSSRX1_HVT src_aox_reg_14__4_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[172]), .CLK(clk), .Q(src_window[172]) );
  DFFSSRX1_HVT src_aox_reg_14__3_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[171]), .CLK(clk), .Q(src_window[171]) );
  DFFSSRX1_HVT src_aox_reg_14__2_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[170]), .CLK(clk), .Q(src_window[170]) );
  DFFSSRX1_HVT src_aox_reg_14__1_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[169]), .CLK(clk), .Q(src_window[169]) );
  DFFSSRX1_HVT src_aox_reg_14__0_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[168]), .CLK(clk), .Q(src_window[168]) );
  DFFSSRX1_HVT src_aox_reg_15__7_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[167]), .CLK(clk), .Q(src_window[167]) );
  DFFSSRX1_HVT src_aox_reg_15__6_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[166]), .CLK(clk), .Q(src_window[166]) );
  DFFSSRX1_HVT src_aox_reg_15__5_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[165]), .CLK(clk), .Q(src_window[165]) );
  DFFSSRX1_HVT src_aox_reg_15__4_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[164]), .CLK(clk), .Q(src_window[164]) );
  DFFSSRX1_HVT src_aox_reg_15__3_ ( .D(1'b0), .SETB(n2560), .RSTB(
        n_src_aox[163]), .CLK(clk), .Q(src_window[163]) );
  DFFSSRX1_HVT src_aox_reg_15__2_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[162]), .CLK(clk), .Q(src_window[162]) );
  DFFSSRX1_HVT src_aox_reg_15__1_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[161]), .CLK(clk), .Q(src_window[161]) );
  DFFSSRX1_HVT src_aox_reg_15__0_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[160]), .CLK(clk), .Q(src_window[160]) );
  DFFSSRX1_HVT src_aox_reg_16__7_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[159]), .CLK(clk), .Q(src_window[159]) );
  DFFSSRX1_HVT src_aox_reg_16__6_ ( .D(1'b0), .SETB(n2560), .RSTB(
        n_src_aox[158]), .CLK(clk), .Q(src_window[158]) );
  DFFSSRX1_HVT src_aox_reg_16__5_ ( .D(1'b0), .SETB(n13200), .RSTB(
        n_src_aox[157]), .CLK(clk), .Q(src_window[157]) );
  DFFSSRX1_HVT src_aox_reg_16__4_ ( .D(1'b0), .SETB(n579), .RSTB(
        n_src_aox[156]), .CLK(clk), .Q(src_window[156]) );
  DFFSSRX1_HVT src_aox_reg_16__3_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[155]), .CLK(clk), .Q(src_window[155]) );
  DFFSSRX1_HVT src_aox_reg_16__2_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[154]), .CLK(clk), .Q(src_window[154]) );
  DFFSSRX1_HVT src_aox_reg_16__1_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[153]), .CLK(clk), .Q(src_window[153]) );
  DFFSSRX1_HVT src_aox_reg_16__0_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[152]), .CLK(clk), .Q(src_window[152]) );
  DFFSSRX1_HVT src_aox_reg_17__7_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[151]), .CLK(clk), .Q(src_window[151]) );
  DFFSSRX1_HVT src_aox_reg_17__6_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[150]), .CLK(clk), .Q(src_window[150]) );
  DFFSSRX1_HVT src_aox_reg_17__5_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[149]), .CLK(clk), .Q(src_window[149]) );
  DFFSSRX1_HVT src_aox_reg_17__4_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[148]), .CLK(clk), .Q(src_window[148]) );
  DFFSSRX1_HVT src_aox_reg_17__3_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[147]), .CLK(clk), .Q(src_window[147]) );
  DFFSSRX1_HVT src_aox_reg_17__2_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[146]), .CLK(clk), .Q(src_window[146]) );
  DFFSSRX1_HVT src_aox_reg_17__1_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[145]), .CLK(clk), .Q(src_window[145]) );
  DFFSSRX1_HVT src_aox_reg_17__0_ ( .D(1'b0), .SETB(n579), .RSTB(
        n_src_aox[144]), .CLK(clk), .Q(src_window[144]) );
  DFFSSRX1_HVT src_aox_reg_18__7_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[143]), .CLK(clk), .Q(src_window[143]) );
  DFFSSRX1_HVT src_aox_reg_18__6_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[142]), .CLK(clk), .Q(src_window[142]) );
  DFFSSRX1_HVT src_aox_reg_18__5_ ( .D(1'b0), .SETB(n579), .RSTB(
        n_src_aox[141]), .CLK(clk), .Q(src_window[141]) );
  DFFSSRX1_HVT src_aox_reg_18__4_ ( .D(1'b0), .SETB(n13200), .RSTB(
        n_src_aox[140]), .CLK(clk), .Q(src_window[140]) );
  DFFSSRX1_HVT src_aox_reg_18__3_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[139]), .CLK(clk), .Q(src_window[139]) );
  DFFSSRX1_HVT src_aox_reg_18__2_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[138]), .CLK(clk), .Q(src_window[138]) );
  DFFSSRX1_HVT src_aox_reg_18__1_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[137]), .CLK(clk), .Q(src_window[137]) );
  DFFSSRX1_HVT src_aox_reg_18__0_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[136]), .CLK(clk), .Q(src_window[136]) );
  DFFSSRX1_HVT src_aox_reg_19__7_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[135]), .CLK(clk), .Q(src_window[135]) );
  DFFSSRX1_HVT src_aox_reg_19__6_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[134]), .CLK(clk), .Q(src_window[134]) );
  DFFSSRX1_HVT src_aox_reg_19__5_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[133]), .CLK(clk), .Q(src_window[133]) );
  DFFSSRX1_HVT src_aox_reg_19__4_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[132]), .CLK(clk), .Q(src_window[132]) );
  DFFSSRX1_HVT src_aox_reg_19__3_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[131]), .CLK(clk), .Q(src_window[131]) );
  DFFSSRX1_HVT src_aox_reg_19__2_ ( .D(1'b0), .SETB(n2560), .RSTB(
        n_src_aox[130]), .CLK(clk), .Q(src_window[130]) );
  DFFSSRX1_HVT src_aox_reg_19__1_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[129]), .CLK(clk), .Q(src_window[129]) );
  DFFSSRX1_HVT src_aox_reg_19__0_ ( .D(1'b0), .SETB(n13200), .RSTB(
        n_src_aox[128]), .CLK(clk), .Q(src_window[128]) );
  DFFSSRX1_HVT src_aox_reg_20__7_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[127]), .CLK(clk), .Q(src_window[127]) );
  DFFSSRX1_HVT src_aox_reg_20__6_ ( .D(1'b0), .SETB(n13200), .RSTB(
        n_src_aox[126]), .CLK(clk), .Q(src_window[126]) );
  DFFSSRX1_HVT src_aox_reg_20__5_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[125]), .CLK(clk), .Q(src_window[125]) );
  DFFSSRX1_HVT src_aox_reg_20__4_ ( .D(1'b0), .SETB(n579), .RSTB(
        n_src_aox[124]), .CLK(clk), .Q(src_window[124]) );
  DFFSSRX1_HVT src_aox_reg_20__3_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[123]), .CLK(clk), .Q(src_window[123]) );
  DFFSSRX1_HVT src_aox_reg_20__2_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[122]), .CLK(clk), .Q(src_window[122]) );
  DFFSSRX1_HVT src_aox_reg_20__1_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[121]), .CLK(clk), .Q(src_window[121]) );
  DFFSSRX1_HVT src_aox_reg_20__0_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[120]), .CLK(clk), .Q(src_window[120]) );
  DFFSSRX1_HVT src_aox_reg_21__7_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[119]), .CLK(clk), .Q(src_window[119]) );
  DFFSSRX1_HVT src_aox_reg_21__6_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[118]), .CLK(clk), .Q(src_window[118]) );
  DFFSSRX1_HVT src_aox_reg_21__5_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[117]), .CLK(clk), .Q(src_window[117]) );
  DFFSSRX1_HVT src_aox_reg_21__4_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[116]), .CLK(clk), .Q(src_window[116]) );
  DFFSSRX1_HVT src_aox_reg_21__3_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[115]), .CLK(clk), .Q(src_window[115]) );
  DFFSSRX1_HVT src_aox_reg_21__2_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[114]), .CLK(clk), .Q(src_window[114]) );
  DFFSSRX1_HVT src_aox_reg_21__1_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[113]), .CLK(clk), .Q(src_window[113]) );
  DFFSSRX1_HVT src_aox_reg_21__0_ ( .D(1'b0), .SETB(n579), .RSTB(
        n_src_aox[112]), .CLK(clk), .Q(src_window[112]) );
  DFFSSRX1_HVT src_aox_reg_22__7_ ( .D(1'b0), .SETB(N346), .RSTB(
        n_src_aox[111]), .CLK(clk), .Q(src_window[111]) );
  DFFSSRX1_HVT src_aox_reg_22__6_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[110]), .CLK(clk), .Q(src_window[110]) );
  DFFSSRX1_HVT src_aox_reg_22__5_ ( .D(1'b0), .SETB(n579), .RSTB(
        n_src_aox[109]), .CLK(clk), .Q(src_window[109]) );
  DFFSSRX1_HVT src_aox_reg_22__4_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[108]), .CLK(clk), .Q(src_window[108]) );
  DFFSSRX1_HVT src_aox_reg_22__3_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[107]), .CLK(clk), .Q(src_window[107]) );
  DFFSSRX1_HVT src_aox_reg_22__2_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[106]), .CLK(clk), .Q(src_window[106]) );
  DFFSSRX1_HVT src_aox_reg_22__1_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[105]), .CLK(clk), .Q(src_window[105]) );
  DFFSSRX1_HVT src_aox_reg_22__0_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[104]), .CLK(clk), .Q(src_window[104]) );
  DFFSSRX1_HVT src_aox_reg_23__7_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[103]), .CLK(clk), .Q(src_window[103]) );
  DFFSSRX1_HVT src_aox_reg_23__6_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[102]), .CLK(clk), .Q(src_window[102]) );
  DFFSSRX1_HVT src_aox_reg_23__5_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[101]), .CLK(clk), .Q(src_window[101]) );
  DFFSSRX1_HVT src_aox_reg_23__4_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[100]), .CLK(clk), .Q(src_window[100]) );
  DFFSSRX1_HVT src_aox_reg_23__3_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[99]), .CLK(clk), .Q(src_window[99]) );
  DFFSSRX1_HVT src_aox_reg_23__2_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[98]), .CLK(clk), .Q(src_window[98]) );
  DFFSSRX1_HVT src_aox_reg_23__1_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[97]), .CLK(clk), .Q(src_window[97]) );
  DFFSSRX1_HVT src_aox_reg_23__0_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[96]), .CLK(clk), .Q(src_window[96]) );
  DFFSSRX1_HVT src_aox_reg_24__7_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[95]), .CLK(clk), .Q(src_window[95]) );
  DFFSSRX1_HVT src_aox_reg_24__6_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[94]), .CLK(clk), .Q(src_window[94]) );
  DFFSSRX1_HVT src_aox_reg_24__5_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[93]), .CLK(clk), .Q(src_window[93]) );
  DFFSSRX1_HVT src_aox_reg_24__4_ ( .D(1'b0), .SETB(n579), .RSTB(n_src_aox[92]), .CLK(clk), .Q(src_window[92]) );
  DFFSSRX1_HVT src_aox_reg_24__3_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[91]), .CLK(clk), .Q(src_window[91]) );
  DFFSSRX1_HVT src_aox_reg_24__2_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[90]), .CLK(clk), .Q(src_window[90]) );
  DFFSSRX1_HVT src_aox_reg_24__1_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[89]), .CLK(clk), .Q(src_window[89]) );
  DFFSSRX1_HVT src_aox_reg_24__0_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[88]), .CLK(clk), .Q(src_window[88]) );
  DFFSSRX1_HVT src_aox_reg_25__7_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[87]), .CLK(clk), .Q(src_window[87]) );
  DFFSSRX1_HVT src_aox_reg_25__6_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[86]), .CLK(clk), .Q(src_window[86]) );
  DFFSSRX1_HVT src_aox_reg_25__5_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[85]), .CLK(clk), .Q(src_window[85]) );
  DFFSSRX1_HVT src_aox_reg_25__4_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[84]), .CLK(clk), .Q(src_window[84]) );
  DFFSSRX1_HVT src_aox_reg_25__3_ ( .D(1'b0), .SETB(n2560), .RSTB(
        n_src_aox[83]), .CLK(clk), .Q(src_window[83]) );
  DFFSSRX1_HVT src_aox_reg_25__2_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[82]), .CLK(clk), .Q(src_window[82]) );
  DFFSSRX1_HVT src_aox_reg_25__1_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[81]), .CLK(clk), .Q(src_window[81]) );
  DFFSSRX1_HVT src_aox_reg_25__0_ ( .D(1'b0), .SETB(n579), .RSTB(n_src_aox[80]), .CLK(clk), .Q(src_window[80]) );
  DFFSSRX1_HVT src_aox_reg_26__7_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[79]), .CLK(clk), .Q(src_window[79]) );
  DFFSSRX1_HVT src_aox_reg_26__6_ ( .D(1'b0), .SETB(n2560), .RSTB(
        n_src_aox[78]), .CLK(clk), .Q(src_window[78]) );
  DFFSSRX1_HVT src_aox_reg_26__5_ ( .D(1'b0), .SETB(n579), .RSTB(n_src_aox[77]), .CLK(clk), .Q(src_window[77]) );
  DFFSSRX1_HVT src_aox_reg_26__4_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[76]), .CLK(clk), .Q(src_window[76]) );
  DFFSSRX1_HVT src_aox_reg_26__3_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[75]), .CLK(clk), .Q(src_window[75]) );
  DFFSSRX1_HVT src_aox_reg_26__2_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[74]), .CLK(clk), .Q(src_window[74]) );
  DFFSSRX1_HVT src_aox_reg_26__1_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[73]), .CLK(clk), .Q(src_window[73]) );
  DFFSSRX1_HVT src_aox_reg_26__0_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[72]), .CLK(clk), .Q(src_window[72]) );
  DFFSSRX1_HVT src_aox_reg_27__7_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[71]), .CLK(clk), .Q(src_window[71]) );
  DFFSSRX1_HVT src_aox_reg_27__6_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[70]), .CLK(clk), .Q(src_window[70]) );
  DFFSSRX1_HVT src_aox_reg_27__5_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[69]), .CLK(clk), .Q(src_window[69]) );
  DFFSSRX1_HVT src_aox_reg_27__4_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[68]), .CLK(clk), .Q(src_window[68]) );
  DFFSSRX1_HVT src_aox_reg_27__3_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[67]), .CLK(clk), .Q(src_window[67]) );
  DFFSSRX1_HVT src_aox_reg_27__2_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[66]), .CLK(clk), .Q(src_window[66]) );
  DFFSSRX1_HVT src_aox_reg_27__1_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[65]), .CLK(clk), .Q(src_window[65]) );
  DFFSSRX1_HVT src_aox_reg_27__0_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[64]), .CLK(clk), .Q(src_window[64]) );
  DFFSSRX1_HVT src_aox_reg_28__7_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[63]), .CLK(clk), .Q(src_window[63]) );
  DFFSSRX1_HVT src_aox_reg_28__6_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[62]), .CLK(clk), .Q(src_window[62]) );
  DFFSSRX1_HVT src_aox_reg_28__5_ ( .D(1'b0), .SETB(n13200), .RSTB(
        n_src_aox[61]), .CLK(clk), .Q(src_window[61]) );
  DFFSSRX1_HVT src_aox_reg_28__4_ ( .D(1'b0), .SETB(N346), .RSTB(n_src_aox[60]), .CLK(clk), .Q(src_window[60]) );
  DFFSSRX1_HVT src_aox_reg_28__3_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[59]), .CLK(clk), .Q(src_window[59]) );
  DFFSSRX1_HVT src_aox_reg_28__2_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[58]), .CLK(clk), .Q(src_window[58]) );
  DFFSSRX1_HVT src_aox_reg_28__1_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[57]), .CLK(clk), .Q(src_window[57]) );
  DFFSSRX1_HVT src_aox_reg_28__0_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[56]), .CLK(clk), .Q(src_window[56]) );
  DFFSSRX1_HVT src_aox_reg_29__7_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[55]), .CLK(clk), .Q(src_window[55]) );
  DFFSSRX1_HVT src_aox_reg_29__6_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[54]), .CLK(clk), .Q(src_window[54]) );
  DFFSSRX1_HVT src_aox_reg_29__5_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[53]), .CLK(clk), .Q(src_window[53]) );
  DFFSSRX1_HVT src_aox_reg_29__4_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[52]), .CLK(clk), .Q(src_window[52]) );
  DFFSSRX1_HVT src_aox_reg_29__3_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[51]), .CLK(clk), .Q(src_window[51]) );
  DFFSSRX1_HVT src_aox_reg_29__2_ ( .D(1'b0), .SETB(N346), .RSTB(n_src_aox[50]), .CLK(clk), .Q(src_window[50]) );
  DFFSSRX1_HVT src_aox_reg_29__1_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[49]), .CLK(clk), .Q(src_window[49]) );
  DFFSSRX1_HVT src_aox_reg_29__0_ ( .D(1'b0), .SETB(n579), .RSTB(n_src_aox[48]), .CLK(clk), .Q(src_window[48]) );
  DFFSSRX1_HVT src_aox_reg_30__7_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[47]), .CLK(clk), .Q(src_window[47]) );
  DFFSSRX1_HVT src_aox_reg_30__6_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[46]), .CLK(clk), .Q(src_window[46]) );
  DFFSSRX1_HVT src_aox_reg_30__5_ ( .D(1'b0), .SETB(n579), .RSTB(n_src_aox[45]), .CLK(clk), .Q(src_window[45]) );
  DFFSSRX1_HVT src_aox_reg_30__4_ ( .D(1'b0), .SETB(n13200), .RSTB(
        n_src_aox[44]), .CLK(clk), .Q(src_window[44]) );
  DFFSSRX1_HVT src_aox_reg_30__3_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[43]), .CLK(clk), .Q(src_window[43]) );
  DFFSSRX1_HVT src_aox_reg_30__2_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[42]), .CLK(clk), .Q(src_window[42]) );
  DFFSSRX1_HVT src_aox_reg_30__1_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[41]), .CLK(clk), .Q(src_window[41]) );
  DFFSSRX1_HVT src_aox_reg_30__0_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[40]), .CLK(clk), .Q(src_window[40]) );
  DFFSSRX1_HVT src_aox_reg_31__7_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[39]), .CLK(clk), .Q(src_window[39]) );
  DFFSSRX1_HVT src_aox_reg_31__6_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[38]), .CLK(clk), .Q(src_window[38]) );
  DFFSSRX1_HVT src_aox_reg_31__5_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[37]), .CLK(clk), .Q(src_window[37]) );
  DFFSSRX1_HVT src_aox_reg_31__4_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[36]), .CLK(clk), .Q(src_window[36]) );
  DFFSSRX1_HVT src_aox_reg_31__3_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[35]), .CLK(clk), .Q(src_window[35]) );
  DFFSSRX1_HVT src_aox_reg_31__2_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[34]), .CLK(clk), .Q(src_window[34]) );
  DFFSSRX1_HVT src_aox_reg_31__1_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[33]), .CLK(clk), .Q(src_window[33]) );
  DFFSSRX1_HVT src_aox_reg_31__0_ ( .D(1'b0), .SETB(n13200), .RSTB(
        n_src_aox[32]), .CLK(clk), .Q(src_window[32]) );
  DFFSSRX1_HVT src_aox_reg_32__7_ ( .D(1'b0), .SETB(N346), .RSTB(n_src_aox[31]), .CLK(clk), .Q(src_window[31]) );
  DFFSSRX1_HVT src_aox_reg_32__6_ ( .D(1'b0), .SETB(n2540), .RSTB(
        n_src_aox[30]), .CLK(clk), .Q(src_window[30]) );
  DFFSSRX1_HVT src_aox_reg_32__5_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[29]), .CLK(clk), .Q(src_window[29]) );
  DFFSSRX1_HVT src_aox_reg_32__4_ ( .D(1'b0), .SETB(N346), .RSTB(n_src_aox[28]), .CLK(clk), .Q(src_window[28]) );
  DFFSSRX1_HVT src_aox_reg_32__3_ ( .D(1'b0), .SETB(n13200), .RSTB(
        n_src_aox[27]), .CLK(clk), .Q(src_window[27]) );
  DFFSSRX1_HVT src_aox_reg_32__2_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[26]), .CLK(clk), .Q(src_window[26]) );
  DFFSSRX1_HVT src_aox_reg_32__1_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[25]), .CLK(clk), .Q(src_window[25]) );
  DFFSSRX1_HVT src_aox_reg_32__0_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[24]), .CLK(clk), .Q(src_window[24]) );
  DFFSSRX1_HVT src_aox_reg_33__7_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[23]), .CLK(clk), .Q(src_window[23]) );
  DFFSSRX1_HVT src_aox_reg_33__6_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[22]), .CLK(clk), .Q(src_window[22]) );
  DFFSSRX1_HVT src_aox_reg_33__5_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[21]), .CLK(clk), .Q(src_window[21]) );
  DFFSSRX1_HVT src_aox_reg_33__4_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[20]), .CLK(clk), .Q(src_window[20]) );
  DFFSSRX1_HVT src_aox_reg_33__3_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[19]), .CLK(clk), .Q(src_window[19]) );
  DFFSSRX1_HVT src_aox_reg_33__2_ ( .D(1'b0), .SETB(n13200), .RSTB(
        n_src_aox[18]), .CLK(clk), .Q(src_window[18]) );
  DFFSSRX1_HVT src_aox_reg_33__1_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[17]), .CLK(clk), .Q(src_window[17]) );
  DFFSSRX1_HVT src_aox_reg_33__0_ ( .D(1'b0), .SETB(n579), .RSTB(n_src_aox[16]), .CLK(clk), .Q(src_window[16]) );
  DFFSSRX1_HVT src_aox_reg_34__7_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[15]), .CLK(clk), .Q(src_window[15]) );
  DFFSSRX1_HVT src_aox_reg_34__6_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[14]), .CLK(clk), .Q(src_window[14]) );
  DFFSSRX1_HVT src_aox_reg_34__5_ ( .D(1'b0), .SETB(n579), .RSTB(n_src_aox[13]), .CLK(clk), .Q(src_window[13]) );
  DFFSSRX1_HVT src_aox_reg_34__4_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[12]), .CLK(clk), .Q(src_window[12]) );
  DFFSSRX1_HVT src_aox_reg_34__3_ ( .D(1'b0), .SETB(n2550), .RSTB(
        n_src_aox[11]), .CLK(clk), .Q(src_window[11]) );
  DFFSSRX1_HVT src_aox_reg_34__2_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[10]), .CLK(clk), .Q(src_window[10]) );
  DFFSSRX1_HVT src_aox_reg_34__1_ ( .D(1'b0), .SETB(n9900), .RSTB(n_src_aox[9]), .CLK(clk), .Q(src_window[9]) );
  DFFSSRX1_HVT src_aox_reg_34__0_ ( .D(1'b0), .SETB(n2590), .RSTB(n_src_aox[8]), .CLK(clk), .Q(src_window[8]) );
  DFFSSRX1_HVT src_aox_reg_35__7_ ( .D(1'b0), .SETB(n11500), .RSTB(
        n_src_aox[7]), .CLK(clk), .Q(src_window[7]) );
  DFFSSRX1_HVT src_aox_reg_35__6_ ( .D(1'b0), .SETB(n9800), .RSTB(n_src_aox[6]), .CLK(clk), .Q(src_window[6]) );
  DFFSSRX1_HVT src_aox_reg_35__5_ ( .D(1'b0), .SETB(n2590), .RSTB(n_src_aox[5]), .CLK(clk), .Q(src_window[5]) );
  DFFSSRX1_HVT src_aox_reg_35__4_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[4]), .CLK(clk), .Q(src_window[4]) );
  DFFSSRX1_HVT src_aox_reg_35__3_ ( .D(1'b0), .SETB(n2560), .RSTB(n_src_aox[3]), .CLK(clk), .Q(src_window[3]) );
  DFFSSRX1_HVT src_aox_reg_35__2_ ( .D(1'b0), .SETB(n2540), .RSTB(n_src_aox[2]), .CLK(clk), .Q(src_window[2]) );
  DFFSSRX1_HVT src_aox_reg_35__1_ ( .D(1'b0), .SETB(n2580), .RSTB(n_src_aox[1]), .CLK(clk), .Q(src_window[1]) );
  DFFSSRX1_HVT src_aox_reg_35__0_ ( .D(1'b0), .SETB(n9800), .RSTB(n_src_aox[0]), .CLK(clk), .Q(src_window[0]) );
  DFFSSRX1_HVT conv1_weight_reg_99_ ( .D(1'b0), .SETB(n12100), .RSTB(
        sram_rdata_weight[99]), .CLK(clk), .Q(conv1_weight[99]) );
  DFFSSRX1_HVT weight_reg_99_ ( .D(1'b0), .SETB(n13500), .RSTB(
        conv1_weight[99]), .CLK(clk), .Q(weight[99]) );
  DFFSSRX1_HVT conv1_weight_reg_98_ ( .D(1'b0), .SETB(n13300), .RSTB(
        sram_rdata_weight[98]), .CLK(clk), .Q(conv1_weight[98]) );
  DFFSSRX1_HVT weight_reg_98_ ( .D(1'b0), .SETB(n2430), .RSTB(conv1_weight[98]), .CLK(clk), .Q(weight[98]) );
  DFFSSRX1_HVT conv1_weight_reg_97_ ( .D(1'b0), .SETB(n12100), .RSTB(
        sram_rdata_weight[97]), .CLK(clk), .Q(conv1_weight[97]) );
  DFFSSRX1_HVT weight_reg_97_ ( .D(1'b0), .SETB(n2500), .RSTB(conv1_weight[97]), .CLK(clk), .Q(weight[97]) );
  DFFSSRX1_HVT conv1_weight_reg_96_ ( .D(1'b0), .SETB(n2390), .RSTB(
        sram_rdata_weight[96]), .CLK(clk), .Q(conv1_weight[96]) );
  DFFSSRX1_HVT weight_reg_96_ ( .D(1'b0), .SETB(n2420), .RSTB(conv1_weight[96]), .CLK(clk), .Q(weight[96]) );
  DFFSSRX1_HVT conv1_weight_reg_95_ ( .D(1'b0), .SETB(n2830), .RSTB(
        sram_rdata_weight[95]), .CLK(clk), .Q(conv1_weight[95]) );
  DFFSSRX1_HVT weight_reg_95_ ( .D(1'b0), .SETB(n2490), .RSTB(conv1_weight[95]), .CLK(clk), .Q(weight[95]) );
  DFFSSRX1_HVT conv1_weight_reg_94_ ( .D(1'b0), .SETB(n2380), .RSTB(
        sram_rdata_weight[94]), .CLK(clk), .Q(conv1_weight[94]) );
  DFFSSRX1_HVT weight_reg_94_ ( .D(1'b0), .SETB(n2440), .RSTB(conv1_weight[94]), .CLK(clk), .Q(weight[94]) );
  DFFSSRX1_HVT conv1_weight_reg_93_ ( .D(1'b0), .SETB(n2470), .RSTB(
        sram_rdata_weight[93]), .CLK(clk), .Q(conv1_weight[93]) );
  DFFSSRX1_HVT weight_reg_93_ ( .D(1'b0), .SETB(n2510), .RSTB(conv1_weight[93]), .CLK(clk), .Q(weight[93]) );
  DFFSSRX1_HVT conv1_weight_reg_92_ ( .D(1'b0), .SETB(n2400), .RSTB(
        sram_rdata_weight[92]), .CLK(clk), .Q(conv1_weight[92]) );
  DFFSSRX1_HVT weight_reg_92_ ( .D(1'b0), .SETB(n12100), .RSTB(
        conv1_weight[92]), .CLK(clk), .Q(weight[92]) );
  DFFSSRX1_HVT conv1_weight_reg_91_ ( .D(1'b0), .SETB(n12300), .RSTB(
        sram_rdata_weight[91]), .CLK(clk), .Q(conv1_weight[91]) );
  DFFSSRX1_HVT weight_reg_91_ ( .D(1'b0), .SETB(n12000), .RSTB(
        conv1_weight[91]), .CLK(clk), .Q(weight[91]) );
  DFFSSRX1_HVT conv1_weight_reg_90_ ( .D(1'b0), .SETB(n12200), .RSTB(
        sram_rdata_weight[90]), .CLK(clk), .Q(conv1_weight[90]) );
  DFFSSRX1_HVT weight_reg_90_ ( .D(1'b0), .SETB(n2430), .RSTB(conv1_weight[90]), .CLK(clk), .Q(weight[90]) );
  DFFSSRX1_HVT conv1_weight_reg_89_ ( .D(1'b0), .SETB(n12300), .RSTB(
        sram_rdata_weight[89]), .CLK(clk), .Q(conv1_weight[89]) );
  DFFSSRX1_HVT weight_reg_89_ ( .D(1'b0), .SETB(n2500), .RSTB(conv1_weight[89]), .CLK(clk), .Q(weight[89]) );
  DFFSSRX1_HVT conv1_weight_reg_88_ ( .D(1'b0), .SETB(n2390), .RSTB(
        sram_rdata_weight[88]), .CLK(clk), .Q(conv1_weight[88]) );
  DFFSSRX1_HVT weight_reg_88_ ( .D(1'b0), .SETB(n2450), .RSTB(conv1_weight[88]), .CLK(clk), .Q(weight[88]) );
  DFFSSRX1_HVT conv1_weight_reg_87_ ( .D(1'b0), .SETB(n2400), .RSTB(
        sram_rdata_weight[87]), .CLK(clk), .Q(conv1_weight[87]) );
  DFFSSRX1_HVT weight_reg_87_ ( .D(1'b0), .SETB(n2520), .RSTB(conv1_weight[87]), .CLK(clk), .Q(weight[87]) );
  DFFSSRX1_HVT conv1_weight_reg_86_ ( .D(1'b0), .SETB(n2410), .RSTB(
        sram_rdata_weight[86]), .CLK(clk), .Q(conv1_weight[86]) );
  DFFSSRX1_HVT weight_reg_86_ ( .D(1'b0), .SETB(n2440), .RSTB(conv1_weight[86]), .CLK(clk), .Q(weight[86]) );
  DFFSSRX1_HVT conv1_weight_reg_85_ ( .D(1'b0), .SETB(n2470), .RSTB(
        sram_rdata_weight[85]), .CLK(clk), .Q(conv1_weight[85]) );
  DFFSSRX1_HVT weight_reg_85_ ( .D(1'b0), .SETB(n2510), .RSTB(conv1_weight[85]), .CLK(clk), .Q(weight[85]) );
  DFFSSRX1_HVT conv1_weight_reg_84_ ( .D(1'b0), .SETB(n2400), .RSTB(
        sram_rdata_weight[84]), .CLK(clk), .Q(conv1_weight[84]) );
  DFFSSRX1_HVT weight_reg_84_ ( .D(1'b0), .SETB(n12100), .RSTB(
        conv1_weight[84]), .CLK(clk), .Q(weight[84]) );
  DFFSSRX1_HVT conv1_weight_reg_83_ ( .D(1'b0), .SETB(n12300), .RSTB(
        sram_rdata_weight[83]), .CLK(clk), .Q(conv1_weight[83]) );
  DFFSSRX1_HVT weight_reg_83_ ( .D(1'b0), .SETB(n12000), .RSTB(
        conv1_weight[83]), .CLK(clk), .Q(weight[83]) );
  DFFSSRX1_HVT conv1_weight_reg_82_ ( .D(1'b0), .SETB(n12200), .RSTB(
        sram_rdata_weight[82]), .CLK(clk), .Q(conv1_weight[82]) );
  DFFSSRX1_HVT weight_reg_82_ ( .D(1'b0), .SETB(n2420), .RSTB(conv1_weight[82]), .CLK(clk), .Q(weight[82]) );
  DFFSSRX1_HVT conv1_weight_reg_81_ ( .D(1'b0), .SETB(n2850), .RSTB(
        sram_rdata_weight[81]), .CLK(clk), .Q(conv1_weight[81]) );
  DFFSSRX1_HVT weight_reg_81_ ( .D(1'b0), .SETB(n2490), .RSTB(conv1_weight[81]), .CLK(clk), .Q(weight[81]) );
  DFFSSRX1_HVT conv1_weight_reg_80_ ( .D(1'b0), .SETB(n2380), .RSTB(
        sram_rdata_weight[80]), .CLK(clk), .Q(conv1_weight[80]) );
  DFFSSRX1_HVT weight_reg_80_ ( .D(1'b0), .SETB(n2420), .RSTB(conv1_weight[80]), .CLK(clk), .Q(weight[80]) );
  DFFSSRX1_HVT conv1_weight_reg_79_ ( .D(1'b0), .SETB(n2850), .RSTB(
        sram_rdata_weight[79]), .CLK(clk), .Q(conv1_weight[79]) );
  DFFSSRX1_HVT weight_reg_79_ ( .D(1'b0), .SETB(n2490), .RSTB(conv1_weight[79]), .CLK(clk), .Q(weight[79]) );
  DFFSSRX1_HVT conv1_weight_reg_78_ ( .D(1'b0), .SETB(n2380), .RSTB(
        sram_rdata_weight[78]), .CLK(clk), .Q(conv1_weight[78]) );
  DFFSSRX1_HVT weight_reg_78_ ( .D(1'b0), .SETB(n2440), .RSTB(conv1_weight[78]), .CLK(clk), .Q(weight[78]) );
  DFFSSRX1_HVT conv1_weight_reg_77_ ( .D(1'b0), .SETB(n2470), .RSTB(
        sram_rdata_weight[77]), .CLK(clk), .Q(conv1_weight[77]) );
  DFFSSRX1_HVT weight_reg_77_ ( .D(1'b0), .SETB(n2510), .RSTB(conv1_weight[77]), .CLK(clk), .Q(weight[77]) );
  DFFSSRX1_HVT conv1_weight_reg_76_ ( .D(1'b0), .SETB(n2400), .RSTB(
        sram_rdata_weight[76]), .CLK(clk), .Q(conv1_weight[76]) );
  DFFSSRX1_HVT weight_reg_76_ ( .D(1'b0), .SETB(n13400), .RSTB(
        conv1_weight[76]), .CLK(clk), .Q(weight[76]) );
  DFFSSRX1_HVT conv1_weight_reg_75_ ( .D(1'b0), .SETB(n12200), .RSTB(
        sram_rdata_weight[75]), .CLK(clk), .Q(conv1_weight[75]) );
  DFFSSRX1_HVT weight_reg_75_ ( .D(1'b0), .SETB(n13500), .RSTB(
        conv1_weight[75]), .CLK(clk), .Q(weight[75]) );
  DFFSSRX1_HVT conv1_weight_reg_74_ ( .D(1'b0), .SETB(n13300), .RSTB(
        sram_rdata_weight[74]), .CLK(clk), .Q(conv1_weight[74]) );
  DFFSSRX1_HVT weight_reg_74_ ( .D(1'b0), .SETB(n2450), .RSTB(conv1_weight[74]), .CLK(clk), .Q(weight[74]) );
  DFFSSRX1_HVT conv1_weight_reg_73_ ( .D(1'b0), .SETB(n12300), .RSTB(
        sram_rdata_weight[73]), .CLK(clk), .Q(conv1_weight[73]) );
  DFFSSRX1_HVT weight_reg_73_ ( .D(1'b0), .SETB(n2520), .RSTB(conv1_weight[73]), .CLK(clk), .Q(weight[73]) );
  DFFSSRX1_HVT conv1_weight_reg_72_ ( .D(1'b0), .SETB(n2410), .RSTB(
        sram_rdata_weight[72]), .CLK(clk), .Q(conv1_weight[72]) );
  DFFSSRX1_HVT weight_reg_72_ ( .D(1'b0), .SETB(n2450), .RSTB(conv1_weight[72]), .CLK(clk), .Q(weight[72]) );
  DFFSSRX1_HVT conv1_weight_reg_71_ ( .D(1'b0), .SETB(n2440), .RSTB(
        sram_rdata_weight[71]), .CLK(clk), .Q(conv1_weight[71]) );
  DFFSSRX1_HVT weight_reg_71_ ( .D(1'b0), .SETB(n2520), .RSTB(conv1_weight[71]), .CLK(clk), .Q(weight[71]) );
  DFFSSRX1_HVT conv1_weight_reg_70_ ( .D(1'b0), .SETB(n2410), .RSTB(
        sram_rdata_weight[70]), .CLK(clk), .Q(conv1_weight[70]) );
  DFFSSRX1_HVT weight_reg_70_ ( .D(1'b0), .SETB(n2440), .RSTB(conv1_weight[70]), .CLK(clk), .Q(weight[70]) );
  DFFSSRX1_HVT conv1_weight_reg_69_ ( .D(1'b0), .SETB(n2470), .RSTB(
        sram_rdata_weight[69]), .CLK(clk), .Q(conv1_weight[69]) );
  DFFSSRX1_HVT weight_reg_69_ ( .D(1'b0), .SETB(n2510), .RSTB(conv1_weight[69]), .CLK(clk), .Q(weight[69]) );
  DFFSSRX1_HVT conv1_weight_reg_68_ ( .D(1'b0), .SETB(n2400), .RSTB(
        sram_rdata_weight[68]), .CLK(clk), .Q(conv1_weight[68]) );
  DFFSSRX1_HVT weight_reg_68_ ( .D(1'b0), .SETB(n12100), .RSTB(
        conv1_weight[68]), .CLK(clk), .Q(weight[68]) );
  DFFSSRX1_HVT conv1_weight_reg_67_ ( .D(1'b0), .SETB(n12300), .RSTB(
        sram_rdata_weight[67]), .CLK(clk), .Q(conv1_weight[67]) );
  DFFSSRX1_HVT weight_reg_67_ ( .D(1'b0), .SETB(n12000), .RSTB(
        conv1_weight[67]), .CLK(clk), .Q(weight[67]) );
  DFFSSRX1_HVT conv1_weight_reg_66_ ( .D(1'b0), .SETB(n12200), .RSTB(
        sram_rdata_weight[66]), .CLK(clk), .Q(conv1_weight[66]) );
  DFFSSRX1_HVT weight_reg_66_ ( .D(1'b0), .SETB(n2430), .RSTB(conv1_weight[66]), .CLK(clk), .Q(weight[66]) );
  DFFSSRX1_HVT conv1_weight_reg_65_ ( .D(1'b0), .SETB(n12200), .RSTB(
        sram_rdata_weight[65]), .CLK(clk), .Q(conv1_weight[65]) );
  DFFSSRX1_HVT weight_reg_65_ ( .D(1'b0), .SETB(n2500), .RSTB(conv1_weight[65]), .CLK(clk), .Q(weight[65]) );
  DFFSSRX1_HVT conv1_weight_reg_64_ ( .D(1'b0), .SETB(n2390), .RSTB(
        sram_rdata_weight[64]), .CLK(clk), .Q(conv1_weight[64]) );
  DFFSSRX1_HVT weight_reg_64_ ( .D(1'b0), .SETB(n2420), .RSTB(conv1_weight[64]), .CLK(clk), .Q(weight[64]) );
  DFFSSRX1_HVT conv1_weight_reg_63_ ( .D(1'b0), .SETB(n2840), .RSTB(
        sram_rdata_weight[63]), .CLK(clk), .Q(conv1_weight[63]) );
  DFFSSRX1_HVT weight_reg_63_ ( .D(1'b0), .SETB(n2490), .RSTB(conv1_weight[63]), .CLK(clk), .Q(weight[63]) );
  DFFSSRX1_HVT conv1_weight_reg_62_ ( .D(1'b0), .SETB(n2380), .RSTB(
        sram_rdata_weight[62]), .CLK(clk), .Q(conv1_weight[62]) );
  DFFSSRX1_HVT weight_reg_62_ ( .D(1'b0), .SETB(n2440), .RSTB(conv1_weight[62]), .CLK(clk), .Q(weight[62]) );
  DFFSSRX1_HVT conv1_weight_reg_61_ ( .D(1'b0), .SETB(n2470), .RSTB(
        sram_rdata_weight[61]), .CLK(clk), .Q(conv1_weight[61]) );
  DFFSSRX1_HVT weight_reg_61_ ( .D(1'b0), .SETB(n2510), .RSTB(conv1_weight[61]), .CLK(clk), .Q(weight[61]) );
  DFFSSRX1_HVT conv1_weight_reg_60_ ( .D(1'b0), .SETB(n2400), .RSTB(
        sram_rdata_weight[60]), .CLK(clk), .Q(conv1_weight[60]) );
  DFFSSRX1_HVT weight_reg_60_ ( .D(1'b0), .SETB(n12100), .RSTB(
        conv1_weight[60]), .CLK(clk), .Q(weight[60]) );
  DFFSSRX1_HVT conv1_weight_reg_59_ ( .D(1'b0), .SETB(n12300), .RSTB(
        sram_rdata_weight[59]), .CLK(clk), .Q(conv1_weight[59]) );
  DFFSSRX1_HVT weight_reg_59_ ( .D(1'b0), .SETB(n12000), .RSTB(
        conv1_weight[59]), .CLK(clk), .Q(weight[59]) );
  DFFSSRX1_HVT conv1_weight_reg_58_ ( .D(1'b0), .SETB(n12200), .RSTB(
        sram_rdata_weight[58]), .CLK(clk), .Q(conv1_weight[58]) );
  DFFSSRX1_HVT weight_reg_58_ ( .D(1'b0), .SETB(n2430), .RSTB(conv1_weight[58]), .CLK(clk), .Q(weight[58]) );
  DFFSSRX1_HVT conv1_weight_reg_57_ ( .D(1'b0), .SETB(n12000), .RSTB(
        sram_rdata_weight[57]), .CLK(clk), .Q(conv1_weight[57]) );
  DFFSSRX1_HVT weight_reg_57_ ( .D(1'b0), .SETB(n2500), .RSTB(conv1_weight[57]), .CLK(clk), .Q(weight[57]) );
  DFFSSRX1_HVT conv1_weight_reg_56_ ( .D(1'b0), .SETB(n2390), .RSTB(
        sram_rdata_weight[56]), .CLK(clk), .Q(conv1_weight[56]) );
  DFFSSRX1_HVT weight_reg_56_ ( .D(1'b0), .SETB(n2450), .RSTB(conv1_weight[56]), .CLK(clk), .Q(weight[56]) );
  DFFSSRX1_HVT conv1_weight_reg_55_ ( .D(1'b0), .SETB(n2840), .RSTB(
        sram_rdata_weight[55]), .CLK(clk), .Q(conv1_weight[55]) );
  DFFSSRX1_HVT weight_reg_55_ ( .D(1'b0), .SETB(n2520), .RSTB(conv1_weight[55]), .CLK(clk), .Q(weight[55]) );
  DFFSSRX1_HVT conv1_weight_reg_54_ ( .D(1'b0), .SETB(n2410), .RSTB(
        sram_rdata_weight[54]), .CLK(clk), .Q(conv1_weight[54]) );
  DFFSSRX1_HVT weight_reg_54_ ( .D(1'b0), .SETB(n2440), .RSTB(conv1_weight[54]), .CLK(clk), .Q(weight[54]) );
  DFFSSRX1_HVT conv1_weight_reg_53_ ( .D(1'b0), .SETB(n2470), .RSTB(
        sram_rdata_weight[53]), .CLK(clk), .Q(conv1_weight[53]) );
  DFFSSRX1_HVT weight_reg_53_ ( .D(1'b0), .SETB(n2510), .RSTB(conv1_weight[53]), .CLK(clk), .Q(weight[53]) );
  DFFSSRX1_HVT conv1_weight_reg_52_ ( .D(1'b0), .SETB(n2400), .RSTB(
        sram_rdata_weight[52]), .CLK(clk), .Q(conv1_weight[52]) );
  DFFSSRX1_HVT weight_reg_52_ ( .D(1'b0), .SETB(n13400), .RSTB(
        conv1_weight[52]), .CLK(clk), .Q(weight[52]) );
  DFFSSRX1_HVT conv1_weight_reg_51_ ( .D(1'b0), .SETB(n12300), .RSTB(
        sram_rdata_weight[51]), .CLK(clk), .Q(conv1_weight[51]) );
  DFFSSRX1_HVT weight_reg_51_ ( .D(1'b0), .SETB(n13500), .RSTB(
        conv1_weight[51]), .CLK(clk), .Q(weight[51]) );
  DFFSSRX1_HVT conv1_weight_reg_50_ ( .D(1'b0), .SETB(n13300), .RSTB(
        sram_rdata_weight[50]), .CLK(clk), .Q(conv1_weight[50]) );
  DFFSSRX1_HVT weight_reg_50_ ( .D(1'b0), .SETB(n2420), .RSTB(conv1_weight[50]), .CLK(clk), .Q(weight[50]) );
  DFFSSRX1_HVT conv1_weight_reg_49_ ( .D(1'b0), .SETB(n2830), .RSTB(
        sram_rdata_weight[49]), .CLK(clk), .Q(conv1_weight[49]) );
  DFFSSRX1_HVT weight_reg_49_ ( .D(1'b0), .SETB(n2490), .RSTB(conv1_weight[49]), .CLK(clk), .Q(weight[49]) );
  DFFSSRX1_HVT conv1_weight_reg_48_ ( .D(1'b0), .SETB(n2380), .RSTB(
        sram_rdata_weight[48]), .CLK(clk), .Q(conv1_weight[48]) );
  DFFSSRX1_HVT weight_reg_48_ ( .D(1'b0), .SETB(n2420), .RSTB(conv1_weight[48]), .CLK(clk), .Q(weight[48]) );
  DFFSSRX1_HVT conv1_weight_reg_47_ ( .D(1'b0), .SETB(n2830), .RSTB(
        sram_rdata_weight[47]), .CLK(clk), .Q(conv1_weight[47]) );
  DFFSSRX1_HVT weight_reg_47_ ( .D(1'b0), .SETB(n2490), .RSTB(conv1_weight[47]), .CLK(clk), .Q(weight[47]) );
  DFFSSRX1_HVT conv1_weight_reg_46_ ( .D(1'b0), .SETB(n2380), .RSTB(
        sram_rdata_weight[46]), .CLK(clk), .Q(conv1_weight[46]) );
  DFFSSRX1_HVT weight_reg_46_ ( .D(1'b0), .SETB(n2440), .RSTB(conv1_weight[46]), .CLK(clk), .Q(weight[46]) );
  DFFSSRX1_HVT conv1_weight_reg_45_ ( .D(1'b0), .SETB(n2470), .RSTB(
        sram_rdata_weight[45]), .CLK(clk), .Q(conv1_weight[45]) );
  DFFSSRX1_HVT weight_reg_45_ ( .D(1'b0), .SETB(n2510), .RSTB(conv1_weight[45]), .CLK(clk), .Q(weight[45]) );
  DFFSSRX1_HVT conv1_weight_reg_44_ ( .D(1'b0), .SETB(n2400), .RSTB(
        sram_rdata_weight[44]), .CLK(clk), .Q(conv1_weight[44]) );
  DFFSSRX1_HVT weight_reg_44_ ( .D(1'b0), .SETB(n12100), .RSTB(
        conv1_weight[44]), .CLK(clk), .Q(weight[44]) );
  DFFSSRX1_HVT conv1_weight_reg_43_ ( .D(1'b0), .SETB(n12300), .RSTB(
        sram_rdata_weight[43]), .CLK(clk), .Q(conv1_weight[43]) );
  DFFSSRX1_HVT weight_reg_43_ ( .D(1'b0), .SETB(n12000), .RSTB(
        conv1_weight[43]), .CLK(clk), .Q(weight[43]) );
  DFFSSRX1_HVT conv1_weight_reg_42_ ( .D(1'b0), .SETB(n12200), .RSTB(
        sram_rdata_weight[42]), .CLK(clk), .Q(conv1_weight[42]) );
  DFFSSRX1_HVT weight_reg_42_ ( .D(1'b0), .SETB(n2450), .RSTB(conv1_weight[42]), .CLK(clk), .Q(weight[42]) );
  DFFSSRX1_HVT conv1_weight_reg_41_ ( .D(1'b0), .SETB(n2840), .RSTB(
        sram_rdata_weight[41]), .CLK(clk), .Q(conv1_weight[41]) );
  DFFSSRX1_HVT weight_reg_41_ ( .D(1'b0), .SETB(n2520), .RSTB(conv1_weight[41]), .CLK(clk), .Q(weight[41]) );
  DFFSSRX1_HVT conv1_weight_reg_40_ ( .D(1'b0), .SETB(n2410), .RSTB(
        sram_rdata_weight[40]), .CLK(clk), .Q(conv1_weight[40]) );
  DFFSSRX1_HVT weight_reg_40_ ( .D(1'b0), .SETB(n2450), .RSTB(conv1_weight[40]), .CLK(clk), .Q(weight[40]) );
  DFFSSRX1_HVT conv1_weight_reg_39_ ( .D(1'b0), .SETB(n2850), .RSTB(
        sram_rdata_weight[39]), .CLK(clk), .Q(conv1_weight[39]) );
  DFFSSRX1_HVT weight_reg_39_ ( .D(1'b0), .SETB(n2520), .RSTB(conv1_weight[39]), .CLK(clk), .Q(weight[39]) );
  DFFSSRX1_HVT conv1_weight_reg_38_ ( .D(1'b0), .SETB(n2410), .RSTB(
        sram_rdata_weight[38]), .CLK(clk), .Q(conv1_weight[38]) );
  DFFSSRX1_HVT weight_reg_38_ ( .D(1'b0), .SETB(n2440), .RSTB(conv1_weight[38]), .CLK(clk), .Q(weight[38]) );
  DFFSSRX1_HVT conv1_weight_reg_37_ ( .D(1'b0), .SETB(n2470), .RSTB(
        sram_rdata_weight[37]), .CLK(clk), .Q(conv1_weight[37]) );
  DFFSSRX1_HVT weight_reg_37_ ( .D(1'b0), .SETB(n2510), .RSTB(conv1_weight[37]), .CLK(clk), .Q(weight[37]) );
  DFFSSRX1_HVT conv1_weight_reg_36_ ( .D(1'b0), .SETB(n2400), .RSTB(
        sram_rdata_weight[36]), .CLK(clk), .Q(conv1_weight[36]) );
  DFFSSRX1_HVT weight_reg_36_ ( .D(1'b0), .SETB(n12100), .RSTB(
        conv1_weight[36]), .CLK(clk), .Q(weight[36]) );
  DFFSSRX1_HVT conv1_weight_reg_35_ ( .D(1'b0), .SETB(n12300), .RSTB(
        sram_rdata_weight[35]), .CLK(clk), .Q(conv1_weight[35]) );
  DFFSSRX1_HVT weight_reg_35_ ( .D(1'b0), .SETB(n12000), .RSTB(
        conv1_weight[35]), .CLK(clk), .Q(weight[35]) );
  DFFSSRX1_HVT conv1_weight_reg_34_ ( .D(1'b0), .SETB(n12200), .RSTB(
        sram_rdata_weight[34]), .CLK(clk), .Q(conv1_weight[34]) );
  DFFSSRX1_HVT weight_reg_34_ ( .D(1'b0), .SETB(n2430), .RSTB(conv1_weight[34]), .CLK(clk), .Q(weight[34]) );
  DFFSSRX1_HVT conv1_weight_reg_33_ ( .D(1'b0), .SETB(n12100), .RSTB(
        sram_rdata_weight[33]), .CLK(clk), .Q(conv1_weight[33]) );
  DFFSSRX1_HVT weight_reg_33_ ( .D(1'b0), .SETB(n2500), .RSTB(conv1_weight[33]), .CLK(clk), .Q(weight[33]) );
  DFFSSRX1_HVT conv1_weight_reg_32_ ( .D(1'b0), .SETB(n2390), .RSTB(
        sram_rdata_weight[32]), .CLK(clk), .Q(conv1_weight[32]) );
  DFFSSRX1_HVT weight_reg_32_ ( .D(1'b0), .SETB(n2420), .RSTB(conv1_weight[32]), .CLK(clk), .Q(weight[32]) );
  DFFSSRX1_HVT conv1_weight_reg_31_ ( .D(1'b0), .SETB(n2850), .RSTB(
        sram_rdata_weight[31]), .CLK(clk), .Q(conv1_weight[31]) );
  DFFSSRX1_HVT weight_reg_31_ ( .D(1'b0), .SETB(n2490), .RSTB(conv1_weight[31]), .CLK(clk), .Q(weight[31]) );
  DFFSSRX1_HVT conv1_weight_reg_30_ ( .D(1'b0), .SETB(n2380), .RSTB(
        sram_rdata_weight[30]), .CLK(clk), .Q(conv1_weight[30]) );
  DFFSSRX1_HVT weight_reg_30_ ( .D(1'b0), .SETB(n2440), .RSTB(conv1_weight[30]), .CLK(clk), .Q(weight[30]) );
  DFFSSRX1_HVT conv1_weight_reg_29_ ( .D(1'b0), .SETB(n2470), .RSTB(
        sram_rdata_weight[29]), .CLK(clk), .Q(conv1_weight[29]) );
  DFFSSRX1_HVT weight_reg_29_ ( .D(1'b0), .SETB(n2510), .RSTB(conv1_weight[29]), .CLK(clk), .Q(weight[29]) );
  DFFSSRX1_HVT conv1_weight_reg_28_ ( .D(1'b0), .SETB(n2400), .RSTB(
        sram_rdata_weight[28]), .CLK(clk), .Q(conv1_weight[28]) );
  DFFSSRX1_HVT weight_reg_28_ ( .D(1'b0), .SETB(n13400), .RSTB(
        conv1_weight[28]), .CLK(clk), .Q(weight[28]) );
  DFFSSRX1_HVT conv1_weight_reg_27_ ( .D(1'b0), .SETB(n12100), .RSTB(
        sram_rdata_weight[27]), .CLK(clk), .Q(conv1_weight[27]) );
  DFFSSRX1_HVT weight_reg_27_ ( .D(1'b0), .SETB(n13500), .RSTB(
        conv1_weight[27]), .CLK(clk), .Q(weight[27]) );
  DFFSSRX1_HVT conv1_weight_reg_26_ ( .D(1'b0), .SETB(n13300), .RSTB(
        sram_rdata_weight[26]), .CLK(clk), .Q(conv1_weight[26]) );
  DFFSSRX1_HVT weight_reg_26_ ( .D(1'b0), .SETB(n2430), .RSTB(conv1_weight[26]), .CLK(clk), .Q(weight[26]) );
  DFFSSRX1_HVT conv1_weight_reg_25_ ( .D(1'b0), .SETB(n2830), .RSTB(
        sram_rdata_weight[25]), .CLK(clk), .Q(conv1_weight[25]) );
  DFFSSRX1_HVT weight_reg_25_ ( .D(1'b0), .SETB(n2500), .RSTB(conv1_weight[25]), .CLK(clk), .Q(weight[25]) );
  DFFSSRX1_HVT conv1_weight_reg_24_ ( .D(1'b0), .SETB(n2390), .RSTB(
        sram_rdata_weight[24]), .CLK(clk), .Q(conv1_weight[24]) );
  DFFSSRX1_HVT weight_reg_24_ ( .D(1'b0), .SETB(n2450), .RSTB(conv1_weight[24]), .CLK(clk), .Q(weight[24]) );
  DFFSSRX1_HVT conv1_weight_reg_23_ ( .D(1'b0), .SETB(n2830), .RSTB(
        sram_rdata_weight[23]), .CLK(clk), .Q(conv1_weight[23]) );
  DFFSSRX1_HVT weight_reg_23_ ( .D(1'b0), .SETB(n2520), .RSTB(conv1_weight[23]), .CLK(clk), .Q(weight[23]) );
  DFFSSRX1_HVT conv1_weight_reg_22_ ( .D(1'b0), .SETB(n2410), .RSTB(
        sram_rdata_weight[22]), .CLK(clk), .Q(conv1_weight[22]) );
  DFFSSRX1_HVT weight_reg_22_ ( .D(1'b0), .SETB(n2440), .RSTB(conv1_weight[22]), .CLK(clk), .Q(weight[22]) );
  DFFSSRX1_HVT conv1_weight_reg_21_ ( .D(1'b0), .SETB(n2470), .RSTB(
        sram_rdata_weight[21]), .CLK(clk), .Q(conv1_weight[21]) );
  DFFSSRX1_HVT weight_reg_21_ ( .D(1'b0), .SETB(n2510), .RSTB(conv1_weight[21]), .CLK(clk), .Q(weight[21]) );
  DFFSSRX1_HVT conv1_weight_reg_20_ ( .D(1'b0), .SETB(n2400), .RSTB(
        sram_rdata_weight[20]), .CLK(clk), .Q(conv1_weight[20]) );
  DFFSSRX1_HVT weight_reg_20_ ( .D(1'b0), .SETB(n12100), .RSTB(
        conv1_weight[20]), .CLK(clk), .Q(weight[20]) );
  DFFSSRX1_HVT conv1_weight_reg_19_ ( .D(1'b0), .SETB(n12300), .RSTB(
        sram_rdata_weight[19]), .CLK(clk), .Q(conv1_weight[19]) );
  DFFSSRX1_HVT weight_reg_19_ ( .D(1'b0), .SETB(n12000), .RSTB(
        conv1_weight[19]), .CLK(clk), .Q(weight[19]) );
  DFFSSRX1_HVT conv1_weight_reg_18_ ( .D(1'b0), .SETB(n12200), .RSTB(
        sram_rdata_weight[18]), .CLK(clk), .Q(conv1_weight[18]) );
  DFFSSRX1_HVT weight_reg_18_ ( .D(1'b0), .SETB(n2420), .RSTB(conv1_weight[18]), .CLK(clk), .Q(weight[18]) );
  DFFSSRX1_HVT conv1_weight_reg_17_ ( .D(1'b0), .SETB(n2840), .RSTB(
        sram_rdata_weight[17]), .CLK(clk), .Q(conv1_weight[17]) );
  DFFSSRX1_HVT weight_reg_17_ ( .D(1'b0), .SETB(n2490), .RSTB(conv1_weight[17]), .CLK(clk), .Q(weight[17]) );
  DFFSSRX1_HVT conv1_weight_reg_16_ ( .D(1'b0), .SETB(n2380), .RSTB(
        sram_rdata_weight[16]), .CLK(clk), .Q(conv1_weight[16]) );
  DFFSSRX1_HVT weight_reg_16_ ( .D(1'b0), .SETB(n2430), .RSTB(conv1_weight[16]), .CLK(clk), .Q(weight[16]) );
  DFFSSRX1_HVT conv1_weight_reg_15_ ( .D(1'b0), .SETB(n13300), .RSTB(
        sram_rdata_weight[15]), .CLK(clk), .Q(conv1_weight[15]) );
  DFFSSRX1_HVT weight_reg_15_ ( .D(1'b0), .SETB(n2500), .RSTB(conv1_weight[15]), .CLK(clk), .Q(weight[15]) );
  DFFSSRX1_HVT conv1_weight_reg_14_ ( .D(1'b0), .SETB(n2390), .RSTB(
        sram_rdata_weight[14]), .CLK(clk), .Q(conv1_weight[14]) );
  DFFSSRX1_HVT weight_reg_14_ ( .D(1'b0), .SETB(n2420), .RSTB(conv1_weight[14]), .CLK(clk), .Q(weight[14]) );
  DFFSSRX1_HVT conv1_weight_reg_13_ ( .D(1'b0), .SETB(n2840), .RSTB(
        sram_rdata_weight[13]), .CLK(clk), .Q(conv1_weight[13]) );
  DFFSSRX1_HVT weight_reg_13_ ( .D(1'b0), .SETB(n2490), .RSTB(conv1_weight[13]), .CLK(clk), .Q(weight[13]) );
  DFFSSRX1_HVT conv1_weight_reg_12_ ( .D(1'b0), .SETB(n2380), .RSTB(
        sram_rdata_weight[12]), .CLK(clk), .Q(conv1_weight[12]) );
  DFFSSRX1_HVT weight_reg_12_ ( .D(1'b0), .SETB(n12100), .RSTB(
        conv1_weight[12]), .CLK(clk), .Q(weight[12]) );
  DFFSSRX1_HVT conv1_weight_reg_11_ ( .D(1'b0), .SETB(n12300), .RSTB(
        sram_rdata_weight[11]), .CLK(clk), .Q(conv1_weight[11]) );
  DFFSSRX1_HVT weight_reg_11_ ( .D(1'b0), .SETB(n12000), .RSTB(
        conv1_weight[11]), .CLK(clk), .Q(weight[11]) );
  DFFSSRX1_HVT conv1_weight_reg_10_ ( .D(1'b0), .SETB(n12200), .RSTB(
        sram_rdata_weight[10]), .CLK(clk), .Q(conv1_weight[10]) );
  DFFSSRX1_HVT weight_reg_10_ ( .D(1'b0), .SETB(n2450), .RSTB(conv1_weight[10]), .CLK(clk), .Q(weight[10]) );
  DFFSSRX1_HVT conv1_weight_reg_9_ ( .D(1'b0), .SETB(n2470), .RSTB(
        sram_rdata_weight[9]), .CLK(clk), .Q(conv1_weight[9]) );
  DFFSSRX1_HVT weight_reg_9_ ( .D(1'b0), .SETB(n2520), .RSTB(conv1_weight[9]), 
        .CLK(clk), .Q(weight[9]) );
  DFFSSRX1_HVT conv1_weight_reg_8_ ( .D(1'b0), .SETB(n2410), .RSTB(
        sram_rdata_weight[8]), .CLK(clk), .Q(conv1_weight[8]) );
  DFFSSRX1_HVT weight_reg_8_ ( .D(1'b0), .SETB(n2430), .RSTB(conv1_weight[8]), 
        .CLK(clk), .Q(weight[8]) );
  DFFSSRX1_HVT conv1_weight_reg_7_ ( .D(1'b0), .SETB(n13500), .RSTB(
        sram_rdata_weight[7]), .CLK(clk), .Q(conv1_weight[7]) );
  DFFSSRX1_HVT weight_reg_7_ ( .D(1'b0), .SETB(n2500), .RSTB(conv1_weight[7]), 
        .CLK(clk), .Q(weight[7]) );
  DFFSSRX1_HVT conv1_weight_reg_6_ ( .D(1'b0), .SETB(n2390), .RSTB(
        sram_rdata_weight[6]), .CLK(clk), .Q(conv1_weight[6]) );
  DFFSSRX1_HVT weight_reg_6_ ( .D(1'b0), .SETB(n2450), .RSTB(conv1_weight[6]), 
        .CLK(clk), .Q(weight[6]) );
  DFFSSRX1_HVT conv1_weight_reg_5_ ( .D(1'b0), .SETB(n2830), .RSTB(
        sram_rdata_weight[5]), .CLK(clk), .Q(conv1_weight[5]) );
  DFFSSRX1_HVT weight_reg_5_ ( .D(1'b0), .SETB(n2520), .RSTB(conv1_weight[5]), 
        .CLK(clk), .Q(weight[5]) );
  DFFSSRX1_HVT conv1_weight_reg_4_ ( .D(1'b0), .SETB(n2410), .RSTB(
        sram_rdata_weight[4]), .CLK(clk), .Q(conv1_weight[4]) );
  DFFSSRX1_HVT weight_reg_4_ ( .D(1'b0), .SETB(n13400), .RSTB(conv1_weight[4]), 
        .CLK(clk), .Q(weight[4]) );
  DFFSSRX1_HVT conv1_weight_reg_3_ ( .D(1'b0), .SETB(n12200), .RSTB(
        sram_rdata_weight[3]), .CLK(clk), .Q(conv1_weight[3]) );
  DFFSSRX1_HVT weight_reg_3_ ( .D(1'b0), .SETB(n13500), .RSTB(conv1_weight[3]), 
        .CLK(clk), .Q(weight[3]) );
  DFFSSRX1_HVT conv1_weight_reg_2_ ( .D(1'b0), .SETB(n13300), .RSTB(
        sram_rdata_weight[2]), .CLK(clk), .Q(conv1_weight[2]) );
  DFFSSRX1_HVT weight_reg_2_ ( .D(1'b0), .SETB(n2430), .RSTB(conv1_weight[2]), 
        .CLK(clk), .Q(weight[2]) );
  DFFSSRX1_HVT conv1_weight_reg_1_ ( .D(1'b0), .SETB(n2510), .RSTB(
        sram_rdata_weight[1]), .CLK(clk), .Q(conv1_weight[1]) );
  DFFSSRX1_HVT weight_reg_1_ ( .D(1'b0), .SETB(n2500), .RSTB(conv1_weight[1]), 
        .CLK(clk), .Q(weight[1]) );
  DFFSSRX1_HVT conv1_weight_reg_0_ ( .D(1'b0), .SETB(n2390), .RSTB(
        sram_rdata_weight[0]), .CLK(clk), .Q(conv1_weight[0]) );
  DFFSSRX1_HVT weight_reg_0_ ( .D(1'b0), .SETB(n2420), .RSTB(conv1_weight[0]), 
        .CLK(clk), .Q(weight[0]) );
  DFFSSRX1_HVT sram_rdata_8_reg_31_ ( .D(1'b0), .SETB(n2840), .RSTB(N326), 
        .CLK(clk), .Q(sram_rdata_8[31]), .QN(n3170) );
  DFFSSRX1_HVT sram_rdata_8_reg_30_ ( .D(1'b0), .SETB(n12000), .RSTB(N325), 
        .CLK(clk), .Q(sram_rdata_8[30]), .QN(n3160) );
  DFFSSRX1_HVT sram_rdata_8_reg_29_ ( .D(1'b0), .SETB(n2410), .RSTB(N324), 
        .CLK(clk), .Q(sram_rdata_8[29]), .QN(n3150) );
  DFFSSRX1_HVT sram_rdata_8_reg_28_ ( .D(1'b0), .SETB(n2420), .RSTB(N323), 
        .CLK(clk), .Q(sram_rdata_8[28]), .QN(n3140) );
  DFFSSRX1_HVT sram_rdata_8_reg_27_ ( .D(1'b0), .SETB(n2830), .RSTB(N322), 
        .CLK(clk), .Q(sram_rdata_8[27]), .QN(n3130) );
  DFFSSRX1_HVT sram_rdata_8_reg_26_ ( .D(1'b0), .SETB(n2520), .RSTB(N321), 
        .CLK(clk), .Q(sram_rdata_8[26]), .QN(n3120) );
  DFFSSRX1_HVT sram_rdata_8_reg_25_ ( .D(1'b0), .SETB(n2410), .RSTB(N320), 
        .CLK(clk), .Q(sram_rdata_8[25]), .QN(n3110) );
  DFFSSRX1_HVT sram_rdata_8_reg_24_ ( .D(1'b0), .SETB(n2420), .RSTB(N319), 
        .CLK(clk), .Q(sram_rdata_8[24]), .QN(n3100) );
  DFFSSRX1_HVT sram_rdata_8_reg_23_ ( .D(1'b0), .SETB(n12300), .RSTB(N318), 
        .CLK(clk), .Q(sram_rdata_8[23]), .QN(n3090) );
  DFFSSRX1_HVT sram_rdata_8_reg_22_ ( .D(1'b0), .SETB(n2520), .RSTB(N317), 
        .CLK(clk), .Q(sram_rdata_8[22]), .QN(n3080) );
  DFFSSRX1_HVT sram_rdata_8_reg_21_ ( .D(1'b0), .SETB(n13300), .RSTB(N316), 
        .CLK(clk), .Q(sram_rdata_8[21]), .QN(n3070) );
  DFFSSRX1_HVT sram_rdata_8_reg_20_ ( .D(1'b0), .SETB(n2420), .RSTB(N315), 
        .CLK(clk), .Q(sram_rdata_8[20]), .QN(n3060) );
  DFFSSRX1_HVT sram_rdata_8_reg_19_ ( .D(1'b0), .SETB(n2850), .RSTB(N314), 
        .CLK(clk), .Q(sram_rdata_8[19]), .QN(n3050) );
  DFFSSRX1_HVT sram_rdata_8_reg_18_ ( .D(1'b0), .SETB(n2520), .RSTB(N313), 
        .CLK(clk), .Q(sram_rdata_8[18]), .QN(n3040) );
  DFFSSRX1_HVT sram_rdata_8_reg_17_ ( .D(1'b0), .SETB(n2390), .RSTB(N312), 
        .CLK(clk), .Q(sram_rdata_8[17]), .QN(n3030) );
  DFFSSRX1_HVT sram_rdata_8_reg_16_ ( .D(1'b0), .SETB(n13400), .RSTB(N311), 
        .CLK(clk), .Q(sram_rdata_8[16]), .QN(n3020) );
  DFFSSRX1_HVT sram_rdata_8_reg_15_ ( .D(1'b0), .SETB(n2400), .RSTB(N310), 
        .CLK(clk), .Q(sram_rdata_8[15]), .QN(n3010) );
  DFFSSRX1_HVT sram_rdata_8_reg_14_ ( .D(1'b0), .SETB(n12000), .RSTB(N309), 
        .CLK(clk), .Q(sram_rdata_8[14]), .QN(n3000) );
  DFFSSRX1_HVT sram_rdata_8_reg_13_ ( .D(1'b0), .SETB(n2390), .RSTB(N308), 
        .CLK(clk), .Q(sram_rdata_8[13]), .QN(n2990) );
  DFFSSRX1_HVT sram_rdata_8_reg_12_ ( .D(1'b0), .SETB(n2450), .RSTB(N307), 
        .CLK(clk), .Q(sram_rdata_8[12]), .QN(n2980) );
  DFFSSRX1_HVT sram_rdata_8_reg_11_ ( .D(1'b0), .SETB(n13400), .RSTB(N306), 
        .CLK(clk), .Q(sram_rdata_8[11]), .QN(n2970) );
  DFFSSRX1_HVT sram_rdata_8_reg_10_ ( .D(1'b0), .SETB(n2500), .RSTB(N305), 
        .CLK(clk), .Q(sram_rdata_8[10]), .QN(n2960) );
  DFFSSRX1_HVT sram_rdata_8_reg_9_ ( .D(1'b0), .SETB(n2380), .RSTB(N304), 
        .CLK(clk), .Q(sram_rdata_8[9]), .QN(n2950) );
  DFFSSRX1_HVT sram_rdata_8_reg_8_ ( .D(1'b0), .SETB(n2450), .RSTB(N303), 
        .CLK(clk), .Q(sram_rdata_8[8]), .QN(n2940) );
  DFFSSRX1_HVT sram_rdata_8_reg_7_ ( .D(1'b0), .SETB(n12300), .RSTB(N302), 
        .CLK(clk), .Q(sram_rdata_8[7]), .QN(n2930) );
  DFFSSRX1_HVT sram_rdata_8_reg_6_ ( .D(1'b0), .SETB(n2500), .RSTB(N301), 
        .CLK(clk), .Q(sram_rdata_8[6]), .QN(n2920) );
  DFFSSRX1_HVT sram_rdata_8_reg_5_ ( .D(1'b0), .SETB(n13300), .RSTB(N300), 
        .CLK(clk), .Q(sram_rdata_8[5]), .QN(n2910) );
  DFFSSRX1_HVT sram_rdata_8_reg_4_ ( .D(1'b0), .SETB(n2450), .RSTB(N299), 
        .CLK(clk), .Q(sram_rdata_8[4]), .QN(n2900) );
  DFFSSRX1_HVT sram_rdata_8_reg_3_ ( .D(1'b0), .SETB(n13500), .RSTB(N298), 
        .CLK(clk), .Q(sram_rdata_8[3]), .QN(n2890) );
  DFFSSRX1_HVT sram_rdata_8_reg_2_ ( .D(1'b0), .SETB(n2490), .RSTB(N297), 
        .CLK(clk), .Q(sram_rdata_8[2]), .QN(n2880) );
  DFFSSRX1_HVT sram_rdata_8_reg_1_ ( .D(1'b0), .SETB(n2390), .RSTB(N296), 
        .CLK(clk), .Q(sram_rdata_8[1]), .QN(n2870) );
  DFFSSRX1_HVT sram_rdata_8_reg_0_ ( .D(1'b0), .SETB(n13400), .RSTB(N295), 
        .CLK(clk), .Q(sram_rdata_8[0]), .QN(n573) );
  DFFSSRX1_HVT sram_rdata_0_reg_31_ ( .D(1'b0), .SETB(n2420), .RSTB(N70), 
        .CLK(clk), .Q(sram_rdata_0[31]), .QN(n476) );
  DFFSSRX1_HVT sram_rdata_0_reg_30_ ( .D(1'b0), .SETB(n2850), .RSTB(N69), 
        .CLK(clk), .Q(sram_rdata_0[30]), .QN(n475) );
  DFFSSRX1_HVT sram_rdata_0_reg_29_ ( .D(1'b0), .SETB(n2520), .RSTB(N68), 
        .CLK(clk), .Q(sram_rdata_0[29]), .QN(n474) );
  DFFSSRX1_HVT sram_rdata_0_reg_28_ ( .D(1'b0), .SETB(n2380), .RSTB(N67), 
        .CLK(clk), .Q(sram_rdata_0[28]), .QN(n473) );
  DFFSSRX1_HVT sram_rdata_0_reg_27_ ( .D(1'b0), .SETB(n13400), .RSTB(N66), 
        .CLK(clk), .Q(sram_rdata_0[27]), .QN(n472) );
  DFFSSRX1_HVT sram_rdata_0_reg_26_ ( .D(1'b0), .SETB(n2440), .RSTB(N65), 
        .CLK(clk), .Q(sram_rdata_0[26]), .QN(n471) );
  DFFSSRX1_HVT sram_rdata_0_reg_25_ ( .D(1'b0), .SETB(n12000), .RSTB(N64), 
        .CLK(clk), .Q(sram_rdata_0[25]), .QN(n4701) );
  DFFSSRX1_HVT sram_rdata_0_reg_24_ ( .D(1'b0), .SETB(n2380), .RSTB(N63), 
        .CLK(clk), .Q(sram_rdata_0[24]), .QN(n469) );
  DFFSSRX1_HVT sram_rdata_0_reg_23_ ( .D(1'b0), .SETB(n2430), .RSTB(N62), 
        .CLK(clk), .Q(sram_rdata_0[23]), .QN(n468) );
  DFFSSRX1_HVT sram_rdata_0_reg_22_ ( .D(1'b0), .SETB(n2470), .RSTB(N61), 
        .CLK(clk), .Q(sram_rdata_0[22]), .QN(n467) );
  DFFSSRX1_HVT sram_rdata_0_reg_21_ ( .D(1'b0), .SETB(n2490), .RSTB(N60), 
        .CLK(clk), .Q(sram_rdata_0[21]), .QN(n466) );
  DFFSSRX1_HVT sram_rdata_0_reg_20_ ( .D(1'b0), .SETB(n2380), .RSTB(N59), 
        .CLK(clk), .Q(sram_rdata_0[20]), .QN(n465) );
  DFFSSRX1_HVT sram_rdata_0_reg_19_ ( .D(1'b0), .SETB(n2430), .RSTB(N58), 
        .CLK(clk), .Q(sram_rdata_0[19]), .QN(n464) );
  DFFSSRX1_HVT sram_rdata_0_reg_18_ ( .D(1'b0), .SETB(n12300), .RSTB(N57), 
        .CLK(clk), .Q(sram_rdata_0[18]), .QN(n463) );
  DFFSSRX1_HVT sram_rdata_0_reg_17_ ( .D(1'b0), .SETB(n2490), .RSTB(N56), 
        .CLK(clk), .Q(sram_rdata_0[17]), .QN(n462) );
  DFFSSRX1_HVT sram_rdata_0_reg_16_ ( .D(1'b0), .SETB(n13300), .RSTB(N55), 
        .CLK(clk), .Q(sram_rdata_0[16]), .QN(n461) );
  DFFSSRX1_HVT sram_rdata_0_reg_15_ ( .D(1'b0), .SETB(n2450), .RSTB(N54), 
        .CLK(clk), .Q(sram_rdata_0[15]), .QN(n4601) );
  DFFSSRX1_HVT sram_rdata_0_reg_14_ ( .D(1'b0), .SETB(n2840), .RSTB(N53), 
        .CLK(clk), .Q(sram_rdata_0[14]), .QN(n459) );
  DFFSSRX1_HVT sram_rdata_0_reg_13_ ( .D(1'b0), .SETB(n2490), .RSTB(N52), 
        .CLK(clk), .Q(sram_rdata_0[13]), .QN(n458) );
  DFFSSRX1_HVT sram_rdata_0_reg_12_ ( .D(1'b0), .SETB(n2410), .RSTB(N51), 
        .CLK(clk), .Q(sram_rdata_0[12]), .QN(n457) );
  DFFSSRX1_HVT sram_rdata_0_reg_11_ ( .D(1'b0), .SETB(n13400), .RSTB(N50), 
        .CLK(clk), .Q(sram_rdata_0[11]), .QN(n456) );
  DFFSSRX1_HVT sram_rdata_0_reg_10_ ( .D(1'b0), .SETB(n2840), .RSTB(N49), 
        .CLK(clk), .Q(sram_rdata_0[10]), .QN(n455) );
  DFFSSRX1_HVT sram_rdata_0_reg_9_ ( .D(1'b0), .SETB(n12000), .RSTB(N48), 
        .CLK(clk), .Q(sram_rdata_0[9]), .QN(n454) );
  DFFSSRX1_HVT sram_rdata_0_reg_8_ ( .D(1'b0), .SETB(n2410), .RSTB(N47), .CLK(
        clk), .Q(sram_rdata_0[8]), .QN(n453) );
  DFFSSRX1_HVT sram_rdata_0_reg_7_ ( .D(1'b0), .SETB(n2420), .RSTB(N46), .CLK(
        clk), .Q(sram_rdata_0[7]), .QN(n452) );
  DFFSSRX1_HVT sram_rdata_0_reg_6_ ( .D(1'b0), .SETB(n2830), .RSTB(N45), .CLK(
        clk), .Q(sram_rdata_0[6]), .QN(n451) );
  DFFSSRX1_HVT sram_rdata_0_reg_5_ ( .D(1'b0), .SETB(n2520), .RSTB(N44), .CLK(
        clk), .Q(sram_rdata_0[5]), .QN(n4501) );
  DFFSSRX1_HVT sram_rdata_0_reg_4_ ( .D(1'b0), .SETB(n2410), .RSTB(N43), .CLK(
        clk), .Q(sram_rdata_0[4]), .QN(n449) );
  DFFSSRX1_HVT sram_rdata_0_reg_3_ ( .D(1'b0), .SETB(n2420), .RSTB(N42), .CLK(
        clk), .Q(sram_rdata_0[3]), .QN(n448) );
  DFFSSRX1_HVT sram_rdata_0_reg_2_ ( .D(1'b0), .SETB(n12300), .RSTB(N41), 
        .CLK(clk), .Q(sram_rdata_0[2]), .QN(n447) );
  DFFSSRX1_HVT sram_rdata_0_reg_1_ ( .D(1'b0), .SETB(n2520), .RSTB(N40), .CLK(
        clk), .Q(sram_rdata_0[1]), .QN(n446) );
  DFFSSRX1_HVT sram_rdata_0_reg_0_ ( .D(1'b0), .SETB(n13500), .RSTB(N39), 
        .CLK(clk), .Q(sram_rdata_0[0]), .QN(n445) );
  DFFSSRX1_HVT sram_rdata_1_reg_31_ ( .D(1'b0), .SETB(n2490), .RSTB(N102), 
        .CLK(clk), .Q(sram_rdata_1[31]), .QN(n381) );
  DFFSSRX1_HVT sram_rdata_1_reg_30_ ( .D(1'b0), .SETB(n2390), .RSTB(N101), 
        .CLK(clk), .Q(sram_rdata_1[30]), .QN(n380) );
  DFFSSRX1_HVT sram_rdata_1_reg_29_ ( .D(1'b0), .SETB(n12100), .RSTB(N100), 
        .CLK(clk), .Q(sram_rdata_1[29]), .QN(n379) );
  DFFSSRX1_HVT sram_rdata_1_reg_28_ ( .D(1'b0), .SETB(n2400), .RSTB(N99), 
        .CLK(clk), .Q(sram_rdata_1[28]), .QN(n378) );
  DFFSSRX1_HVT sram_rdata_1_reg_27_ ( .D(1'b0), .SETB(n13500), .RSTB(N98), 
        .CLK(clk), .Q(sram_rdata_1[27]), .QN(n377) );
  DFFSSRX1_HVT sram_rdata_1_reg_26_ ( .D(1'b0), .SETB(n2390), .RSTB(N97), 
        .CLK(clk), .Q(sram_rdata_1[26]), .QN(n376) );
  DFFSSRX1_HVT sram_rdata_1_reg_25_ ( .D(1'b0), .SETB(n2430), .RSTB(N96), 
        .CLK(clk), .Q(sram_rdata_1[25]), .QN(n375) );
  DFFSSRX1_HVT sram_rdata_1_reg_24_ ( .D(1'b0), .SETB(n2840), .RSTB(N95), 
        .CLK(clk), .Q(sram_rdata_1[24]), .QN(n374) );
  DFFSSRX1_HVT sram_rdata_1_reg_23_ ( .D(1'b0), .SETB(n2500), .RSTB(N94), 
        .CLK(clk), .Q(sram_rdata_1[23]), .QN(n373) );
  DFFSSRX1_HVT sram_rdata_1_reg_22_ ( .D(1'b0), .SETB(n2410), .RSTB(N93), 
        .CLK(clk), .Q(sram_rdata_1[22]), .QN(n372) );
  DFFSSRX1_HVT sram_rdata_1_reg_21_ ( .D(1'b0), .SETB(n2430), .RSTB(N92), 
        .CLK(clk), .Q(sram_rdata_1[21]), .QN(n371) );
  DFFSSRX1_HVT sram_rdata_1_reg_20_ ( .D(1'b0), .SETB(n12300), .RSTB(N91), 
        .CLK(clk), .Q(sram_rdata_1[20]), .QN(n370) );
  DFFSSRX1_HVT sram_rdata_1_reg_19_ ( .D(1'b0), .SETB(n2500), .RSTB(N90), 
        .CLK(clk), .Q(sram_rdata_1[19]), .QN(n369) );
  DFFSSRX1_HVT sram_rdata_1_reg_18_ ( .D(1'b0), .SETB(n12200), .RSTB(N89), 
        .CLK(clk), .Q(sram_rdata_1[18]), .QN(n368) );
  DFFSSRX1_HVT sram_rdata_1_reg_17_ ( .D(1'b0), .SETB(n2420), .RSTB(N88), 
        .CLK(clk), .Q(sram_rdata_1[17]), .QN(n367) );
  DFFSSRX1_HVT sram_rdata_1_reg_16_ ( .D(1'b0), .SETB(n13400), .RSTB(N87), 
        .CLK(clk), .Q(sram_rdata_1[16]), .QN(n366) );
  DFFSSRX1_HVT sram_rdata_1_reg_15_ ( .D(1'b0), .SETB(n2520), .RSTB(N86), 
        .CLK(clk), .Q(sram_rdata_1[15]), .QN(n365) );
  DFFSSRX1_HVT sram_rdata_1_reg_14_ ( .D(1'b0), .SETB(n2380), .RSTB(N85), 
        .CLK(clk), .Q(sram_rdata_1[14]), .QN(n364) );
  DFFSSRX1_HVT sram_rdata_1_reg_13_ ( .D(1'b0), .SETB(n12100), .RSTB(N84), 
        .CLK(clk), .Q(sram_rdata_1[13]), .QN(n363) );
  DFFSSRX1_HVT sram_rdata_1_reg_12_ ( .D(1'b0), .SETB(n2470), .RSTB(N83), 
        .CLK(clk), .Q(sram_rdata_1[12]), .QN(n362) );
  DFFSSRX1_HVT sram_rdata_1_reg_11_ ( .D(1'b0), .SETB(n13500), .RSTB(N82), 
        .CLK(clk), .Q(sram_rdata_1[11]), .QN(n361) );
  DFFSSRX1_HVT sram_rdata_1_reg_10_ ( .D(1'b0), .SETB(n2380), .RSTB(N81), 
        .CLK(clk), .Q(sram_rdata_1[10]), .QN(n360) );
  DFFSSRX1_HVT sram_rdata_1_reg_9_ ( .D(1'b0), .SETB(n2430), .RSTB(N80), .CLK(
        clk), .Q(sram_rdata_1[9]), .QN(n359) );
  DFFSSRX1_HVT sram_rdata_1_reg_8_ ( .D(1'b0), .SETB(n2440), .RSTB(N79), .CLK(
        clk), .Q(sram_rdata_1[8]), .QN(n358) );
  DFFSSRX1_HVT sram_rdata_1_reg_7_ ( .D(1'b0), .SETB(n2490), .RSTB(N78), .CLK(
        clk), .Q(sram_rdata_1[7]), .QN(n357) );
  DFFSSRX1_HVT sram_rdata_1_reg_6_ ( .D(1'b0), .SETB(n2380), .RSTB(N77), .CLK(
        clk), .Q(sram_rdata_1[6]), .QN(n356) );
  DFFSSRX1_HVT sram_rdata_1_reg_5_ ( .D(1'b0), .SETB(n2430), .RSTB(N76), .CLK(
        clk), .Q(sram_rdata_1[5]), .QN(n355) );
  DFFSSRX1_HVT sram_rdata_1_reg_4_ ( .D(1'b0), .SETB(n12300), .RSTB(N75), 
        .CLK(clk), .Q(sram_rdata_1[4]), .QN(n354) );
  DFFSSRX1_HVT sram_rdata_1_reg_3_ ( .D(1'b0), .SETB(n2490), .RSTB(N74), .CLK(
        clk), .Q(sram_rdata_1[3]), .QN(n353) );
  DFFSSRX1_HVT sram_rdata_1_reg_2_ ( .D(1'b0), .SETB(n12200), .RSTB(N73), 
        .CLK(clk), .Q(sram_rdata_1[2]), .QN(n352) );
  DFFSSRX1_HVT sram_rdata_1_reg_1_ ( .D(1'b0), .SETB(n2450), .RSTB(N72), .CLK(
        clk), .Q(sram_rdata_1[1]), .QN(n351) );
  DFFSSRX1_HVT sram_rdata_1_reg_0_ ( .D(1'b0), .SETB(n2430), .RSTB(N71), .CLK(
        clk), .Q(sram_rdata_1[0]), .QN(n350) );
  DFFSSRX1_HVT sram_rdata_2_reg_31_ ( .D(1'b0), .SETB(n2850), .RSTB(N134), 
        .CLK(clk), .Q(sram_rdata_2[31]), .QN(n572) );
  DFFSSRX1_HVT sram_rdata_2_reg_30_ ( .D(1'b0), .SETB(n2500), .RSTB(N133), 
        .CLK(clk), .Q(sram_rdata_2[30]), .QN(n571) );
  DFFSSRX1_HVT sram_rdata_2_reg_29_ ( .D(1'b0), .SETB(n2410), .RSTB(N132), 
        .CLK(clk), .Q(sram_rdata_2[29]), .QN(n5701) );
  DFFSSRX1_HVT sram_rdata_2_reg_28_ ( .D(1'b0), .SETB(n2430), .RSTB(N131), 
        .CLK(clk), .Q(sram_rdata_2[28]), .QN(n569) );
  DFFSSRX1_HVT sram_rdata_2_reg_27_ ( .D(1'b0), .SETB(n12300), .RSTB(N130), 
        .CLK(clk), .Q(sram_rdata_2[27]), .QN(n568) );
  DFFSSRX1_HVT sram_rdata_2_reg_26_ ( .D(1'b0), .SETB(n2500), .RSTB(N129), 
        .CLK(clk), .Q(sram_rdata_2[26]), .QN(n567) );
  DFFSSRX1_HVT sram_rdata_2_reg_25_ ( .D(1'b0), .SETB(n12200), .RSTB(N128), 
        .CLK(clk), .Q(sram_rdata_2[25]), .QN(n566) );
  DFFSSRX1_HVT sram_rdata_2_reg_24_ ( .D(1'b0), .SETB(n2420), .RSTB(N127), 
        .CLK(clk), .Q(sram_rdata_2[24]), .QN(n565) );
  DFFSSRX1_HVT sram_rdata_2_reg_23_ ( .D(1'b0), .SETB(n2840), .RSTB(N126), 
        .CLK(clk), .Q(sram_rdata_2[23]), .QN(n564) );
  DFFSSRX1_HVT sram_rdata_2_reg_22_ ( .D(1'b0), .SETB(n2520), .RSTB(N125), 
        .CLK(clk), .Q(sram_rdata_2[22]), .QN(n563) );
  DFFSSRX1_HVT sram_rdata_2_reg_21_ ( .D(1'b0), .SETB(n2380), .RSTB(N124), 
        .CLK(clk), .Q(sram_rdata_2[21]), .QN(n562) );
  DFFSSRX1_HVT sram_rdata_2_reg_20_ ( .D(1'b0), .SETB(n12100), .RSTB(N123), 
        .CLK(clk), .Q(sram_rdata_2[20]), .QN(n561) );
  DFFSSRX1_HVT sram_rdata_2_reg_19_ ( .D(1'b0), .SETB(n12300), .RSTB(N122), 
        .CLK(clk), .Q(sram_rdata_2[19]), .QN(n5601) );
  DFFSSRX1_HVT sram_rdata_2_reg_18_ ( .D(1'b0), .SETB(n12000), .RSTB(N121), 
        .CLK(clk), .Q(sram_rdata_2[18]), .QN(n559) );
  DFFSSRX1_HVT sram_rdata_2_reg_17_ ( .D(1'b0), .SETB(n2380), .RSTB(N120), 
        .CLK(clk), .Q(sram_rdata_2[17]), .QN(n558) );
  DFFSSRX1_HVT sram_rdata_2_reg_16_ ( .D(1'b0), .SETB(n2430), .RSTB(N119), 
        .CLK(clk), .Q(sram_rdata_2[16]), .QN(n557) );
  DFFSSRX1_HVT sram_rdata_2_reg_15_ ( .D(1'b0), .SETB(n12200), .RSTB(N118), 
        .CLK(clk), .Q(sram_rdata_2[15]), .QN(n556) );
  DFFSSRX1_HVT sram_rdata_2_reg_14_ ( .D(1'b0), .SETB(n2490), .RSTB(N117), 
        .CLK(clk), .Q(sram_rdata_2[14]), .QN(n555) );
  DFFSSRX1_HVT sram_rdata_2_reg_13_ ( .D(1'b0), .SETB(n2380), .RSTB(N116), 
        .CLK(clk), .Q(sram_rdata_2[13]), .QN(n554) );
  DFFSSRX1_HVT sram_rdata_2_reg_12_ ( .D(1'b0), .SETB(n2430), .RSTB(N115), 
        .CLK(clk), .Q(sram_rdata_2[12]), .QN(n553) );
  DFFSSRX1_HVT sram_rdata_2_reg_11_ ( .D(1'b0), .SETB(n12200), .RSTB(N114), 
        .CLK(clk), .Q(sram_rdata_2[11]), .QN(n552) );
  DFFSSRX1_HVT sram_rdata_2_reg_10_ ( .D(1'b0), .SETB(n2490), .RSTB(N113), 
        .CLK(clk), .Q(sram_rdata_2[10]), .QN(n551) );
  DFFSSRX1_HVT sram_rdata_2_reg_9_ ( .D(1'b0), .SETB(n12200), .RSTB(N112), 
        .CLK(clk), .Q(sram_rdata_2[9]), .QN(n5501) );
  DFFSSRX1_HVT sram_rdata_2_reg_8_ ( .D(1'b0), .SETB(n2450), .RSTB(N111), 
        .CLK(clk), .Q(sram_rdata_2[8]), .QN(n549) );
  DFFSSRX1_HVT sram_rdata_2_reg_7_ ( .D(1'b0), .SETB(n2850), .RSTB(N110), 
        .CLK(clk), .Q(sram_rdata_2[7]), .QN(n548) );
  DFFSSRX1_HVT sram_rdata_2_reg_6_ ( .D(1'b0), .SETB(n2490), .RSTB(N109), 
        .CLK(clk), .Q(sram_rdata_2[6]), .QN(n547) );
  DFFSSRX1_HVT sram_rdata_2_reg_5_ ( .D(1'b0), .SETB(n2410), .RSTB(N108), 
        .CLK(clk), .Q(sram_rdata_2[5]), .QN(n546) );
  DFFSSRX1_HVT sram_rdata_2_reg_4_ ( .D(1'b0), .SETB(n12100), .RSTB(N107), 
        .CLK(clk), .Q(sram_rdata_2[4]), .QN(n545) );
  DFFSSRX1_HVT sram_rdata_2_reg_3_ ( .D(1'b0), .SETB(n2830), .RSTB(N106), 
        .CLK(clk), .Q(sram_rdata_2[3]), .QN(n544) );
  DFFSSRX1_HVT sram_rdata_2_reg_2_ ( .D(1'b0), .SETB(n12000), .RSTB(N105), 
        .CLK(clk), .Q(sram_rdata_2[2]), .QN(n543) );
  DFFSSRX1_HVT sram_rdata_2_reg_1_ ( .D(1'b0), .SETB(n2410), .RSTB(N104), 
        .CLK(clk), .Q(sram_rdata_2[1]), .QN(n542) );
  DFFSSRX1_HVT sram_rdata_2_reg_0_ ( .D(1'b0), .SETB(n13300), .RSTB(N103), 
        .CLK(clk), .Q(sram_rdata_2[0]), .QN(n541) );
  DFFSSRX1_HVT sram_rdata_3_reg_31_ ( .D(1'b0), .SETB(n2380), .RSTB(N166), 
        .CLK(clk), .Q(sram_rdata_3[31]), .QN(n444) );
  DFFSSRX1_HVT sram_rdata_3_reg_30_ ( .D(1'b0), .SETB(n2450), .RSTB(N165), 
        .CLK(clk), .Q(sram_rdata_3[30]), .QN(n443) );
  DFFSSRX1_HVT sram_rdata_3_reg_29_ ( .D(1'b0), .SETB(n12300), .RSTB(N164), 
        .CLK(clk), .Q(sram_rdata_3[29]), .QN(n442) );
  DFFSSRX1_HVT sram_rdata_3_reg_28_ ( .D(1'b0), .SETB(n2500), .RSTB(N163), 
        .CLK(clk), .Q(sram_rdata_3[28]), .QN(n441) );
  DFFSSRX1_HVT sram_rdata_3_reg_27_ ( .D(1'b0), .SETB(n13300), .RSTB(N162), 
        .CLK(clk), .Q(sram_rdata_3[27]), .QN(n4401) );
  DFFSSRX1_HVT sram_rdata_3_reg_26_ ( .D(1'b0), .SETB(n2450), .RSTB(N161), 
        .CLK(clk), .Q(sram_rdata_3[26]), .QN(n439) );
  DFFSSRX1_HVT sram_rdata_3_reg_25_ ( .D(1'b0), .SETB(n2470), .RSTB(N160), 
        .CLK(clk), .Q(sram_rdata_3[25]), .QN(n438) );
  DFFSSRX1_HVT sram_rdata_3_reg_24_ ( .D(1'b0), .SETB(n2490), .RSTB(N159), 
        .CLK(clk), .Q(sram_rdata_3[24]), .QN(n437) );
  DFFSSRX1_HVT sram_rdata_3_reg_23_ ( .D(1'b0), .SETB(n2390), .RSTB(N158), 
        .CLK(clk), .Q(sram_rdata_3[23]), .QN(n436) );
  DFFSSRX1_HVT sram_rdata_3_reg_22_ ( .D(1'b0), .SETB(n13400), .RSTB(N157), 
        .CLK(clk), .Q(sram_rdata_3[22]), .QN(n435) );
  DFFSSRX1_HVT sram_rdata_3_reg_21_ ( .D(1'b0), .SETB(n13400), .RSTB(N156), 
        .CLK(clk), .Q(sram_rdata_3[21]), .QN(n434) );
  DFFSSRX1_HVT sram_rdata_3_reg_20_ ( .D(1'b0), .SETB(n12000), .RSTB(N155), 
        .CLK(clk), .Q(sram_rdata_3[20]), .QN(n433) );
  DFFSSRX1_HVT sram_rdata_3_reg_19_ ( .D(1'b0), .SETB(n2390), .RSTB(N154), 
        .CLK(clk), .Q(sram_rdata_3[19]), .QN(n432) );
  DFFSSRX1_HVT sram_rdata_3_reg_18_ ( .D(1'b0), .SETB(n2430), .RSTB(N153), 
        .CLK(clk), .Q(sram_rdata_3[18]), .QN(n431) );
  DFFSSRX1_HVT sram_rdata_3_reg_17_ ( .D(1'b0), .SETB(n2830), .RSTB(N152), 
        .CLK(clk), .Q(sram_rdata_3[17]), .QN(n4301) );
  DFFSSRX1_HVT sram_rdata_3_reg_16_ ( .D(1'b0), .SETB(n2500), .RSTB(N151), 
        .CLK(clk), .Q(sram_rdata_3[16]), .QN(n429) );
  DFFSSRX1_HVT sram_rdata_3_reg_15_ ( .D(1'b0), .SETB(n2410), .RSTB(N150), 
        .CLK(clk), .Q(sram_rdata_3[15]), .QN(n428) );
  DFFSSRX1_HVT sram_rdata_3_reg_14_ ( .D(1'b0), .SETB(n2430), .RSTB(N149), 
        .CLK(clk), .Q(sram_rdata_3[14]), .QN(n427) );
  DFFSSRX1_HVT sram_rdata_3_reg_13_ ( .D(1'b0), .SETB(n12300), .RSTB(N148), 
        .CLK(clk), .Q(sram_rdata_3[13]), .QN(n426) );
  DFFSSRX1_HVT sram_rdata_3_reg_12_ ( .D(1'b0), .SETB(n2500), .RSTB(N147), 
        .CLK(clk), .Q(sram_rdata_3[12]), .QN(n425) );
  DFFSSRX1_HVT sram_rdata_3_reg_11_ ( .D(1'b0), .SETB(n13300), .RSTB(N146), 
        .CLK(clk), .Q(sram_rdata_3[11]), .QN(n424) );
  DFFSSRX1_HVT sram_rdata_3_reg_10_ ( .D(1'b0), .SETB(n2420), .RSTB(N145), 
        .CLK(clk), .Q(sram_rdata_3[10]), .QN(n423) );
  DFFSSRX1_HVT sram_rdata_3_reg_9_ ( .D(1'b0), .SETB(n2400), .RSTB(N144), 
        .CLK(clk), .Q(sram_rdata_3[9]), .QN(n422) );
  DFFSSRX1_HVT sram_rdata_3_reg_8_ ( .D(1'b0), .SETB(n2520), .RSTB(N143), 
        .CLK(clk), .Q(sram_rdata_3[8]), .QN(n421) );
  DFFSSRX1_HVT sram_rdata_3_reg_7_ ( .D(1'b0), .SETB(n2380), .RSTB(N142), 
        .CLK(clk), .Q(sram_rdata_3[7]), .QN(n4201) );
  DFFSSRX1_HVT sram_rdata_3_reg_6_ ( .D(1'b0), .SETB(n13400), .RSTB(N141), 
        .CLK(clk), .Q(sram_rdata_3[6]), .QN(n419) );
  DFFSSRX1_HVT sram_rdata_3_reg_5_ ( .D(1'b0), .SETB(n2510), .RSTB(N140), 
        .CLK(clk), .Q(sram_rdata_3[5]), .QN(n418) );
  DFFSSRX1_HVT sram_rdata_3_reg_4_ ( .D(1'b0), .SETB(n12000), .RSTB(N139), 
        .CLK(clk), .Q(sram_rdata_3[4]), .QN(n417) );
  DFFSSRX1_HVT sram_rdata_3_reg_3_ ( .D(1'b0), .SETB(n2380), .RSTB(N138), 
        .CLK(clk), .Q(sram_rdata_3[3]), .QN(n416) );
  DFFSSRX1_HVT sram_rdata_3_reg_2_ ( .D(1'b0), .SETB(n2430), .RSTB(N137), 
        .CLK(clk), .Q(sram_rdata_3[2]), .QN(n415) );
  DFFSSRX1_HVT sram_rdata_3_reg_1_ ( .D(1'b0), .SETB(n13500), .RSTB(N136), 
        .CLK(clk), .Q(sram_rdata_3[1]), .QN(n414) );
  DFFSSRX1_HVT sram_rdata_3_reg_0_ ( .D(1'b0), .SETB(n2830), .RSTB(N135), 
        .CLK(clk), .Q(sram_rdata_3[0]), .QN(n382) );
  DFFSSRX1_HVT sram_rdata_4_reg_31_ ( .D(1'b0), .SETB(n12300), .RSTB(N198), 
        .CLK(clk), .Q(sram_rdata_4[31]), .QN(n349) );
  DFFSSRX1_HVT sram_rdata_4_reg_30_ ( .D(1'b0), .SETB(n2520), .RSTB(N197), 
        .CLK(clk), .Q(sram_rdata_4[30]), .QN(n348) );
  DFFSSRX1_HVT sram_rdata_4_reg_29_ ( .D(1'b0), .SETB(n12200), .RSTB(N196), 
        .CLK(clk), .Q(sram_rdata_4[29]), .QN(n347) );
  DFFSSRX1_HVT sram_rdata_4_reg_28_ ( .D(1'b0), .SETB(n2420), .RSTB(N195), 
        .CLK(clk), .Q(sram_rdata_4[28]), .QN(n3460) );
  DFFSSRX1_HVT sram_rdata_4_reg_27_ ( .D(1'b0), .SETB(n2510), .RSTB(N194), 
        .CLK(clk), .Q(sram_rdata_4[27]), .QN(n345) );
  DFFSSRX1_HVT sram_rdata_4_reg_26_ ( .D(1'b0), .SETB(n2520), .RSTB(N193), 
        .CLK(clk), .Q(sram_rdata_4[26]), .QN(n344) );
  DFFSSRX1_HVT sram_rdata_4_reg_25_ ( .D(1'b0), .SETB(n2390), .RSTB(N192), 
        .CLK(clk), .Q(sram_rdata_4[25]), .QN(n343) );
  DFFSSRX1_HVT sram_rdata_4_reg_24_ ( .D(1'b0), .SETB(n12100), .RSTB(N191), 
        .CLK(clk), .Q(sram_rdata_4[24]), .QN(n342) );
  DFFSSRX1_HVT sram_rdata_4_reg_23_ ( .D(1'b0), .SETB(n13500), .RSTB(N190), 
        .CLK(clk), .Q(sram_rdata_4[23]), .QN(n341) );
  DFFSSRX1_HVT sram_rdata_4_reg_22_ ( .D(1'b0), .SETB(n13500), .RSTB(N189), 
        .CLK(clk), .Q(sram_rdata_4[22]), .QN(n340) );
  DFFSSRX1_HVT sram_rdata_4_reg_21_ ( .D(1'b0), .SETB(n2390), .RSTB(N188), 
        .CLK(clk), .Q(sram_rdata_4[21]), .QN(n339) );
  DFFSSRX1_HVT sram_rdata_4_reg_20_ ( .D(1'b0), .SETB(n2450), .RSTB(N187), 
        .CLK(clk), .Q(sram_rdata_4[20]), .QN(n338) );
  DFFSSRX1_HVT sram_rdata_4_reg_19_ ( .D(1'b0), .SETB(n2840), .RSTB(N186), 
        .CLK(clk), .Q(sram_rdata_4[19]), .QN(n337) );
  DFFSSRX1_HVT sram_rdata_4_reg_18_ ( .D(1'b0), .SETB(n2500), .RSTB(N185), 
        .CLK(clk), .Q(sram_rdata_4[18]), .QN(n336) );
  DFFSSRX1_HVT sram_rdata_4_reg_17_ ( .D(1'b0), .SETB(n2380), .RSTB(N184), 
        .CLK(clk), .Q(sram_rdata_4[17]), .QN(n335) );
  DFFSSRX1_HVT sram_rdata_4_reg_16_ ( .D(1'b0), .SETB(n2450), .RSTB(N183), 
        .CLK(clk), .Q(sram_rdata_4[16]), .QN(n334) );
  DFFSSRX1_HVT sram_rdata_4_reg_15_ ( .D(1'b0), .SETB(n12300), .RSTB(N182), 
        .CLK(clk), .Q(sram_rdata_4[15]), .QN(n333) );
  DFFSSRX1_HVT sram_rdata_4_reg_14_ ( .D(1'b0), .SETB(n2500), .RSTB(N181), 
        .CLK(clk), .Q(sram_rdata_4[14]), .QN(n332) );
  DFFSSRX1_HVT sram_rdata_4_reg_13_ ( .D(1'b0), .SETB(n12200), .RSTB(N180), 
        .CLK(clk), .Q(sram_rdata_4[13]), .QN(n331) );
  DFFSSRX1_HVT sram_rdata_4_reg_12_ ( .D(1'b0), .SETB(n2450), .RSTB(N179), 
        .CLK(clk), .Q(sram_rdata_4[12]), .QN(n330) );
  DFFSSRX1_HVT sram_rdata_4_reg_11_ ( .D(1'b0), .SETB(n2440), .RSTB(N178), 
        .CLK(clk), .Q(sram_rdata_4[11]), .QN(n329) );
  DFFSSRX1_HVT sram_rdata_4_reg_10_ ( .D(1'b0), .SETB(n2490), .RSTB(N177), 
        .CLK(clk), .Q(sram_rdata_4[10]), .QN(n328) );
  DFFSSRX1_HVT sram_rdata_4_reg_9_ ( .D(1'b0), .SETB(n2390), .RSTB(N176), 
        .CLK(clk), .Q(sram_rdata_4[9]), .QN(n327) );
  DFFSSRX1_HVT sram_rdata_4_reg_8_ ( .D(1'b0), .SETB(n12100), .RSTB(N175), 
        .CLK(clk), .Q(sram_rdata_4[8]), .QN(n3260) );
  DFFSSRX1_HVT sram_rdata_4_reg_7_ ( .D(1'b0), .SETB(n2850), .RSTB(N174), 
        .CLK(clk), .Q(sram_rdata_4[7]), .QN(n3250) );
  DFFSSRX1_HVT sram_rdata_4_reg_6_ ( .D(1'b0), .SETB(n13500), .RSTB(N173), 
        .CLK(clk), .Q(sram_rdata_4[6]), .QN(n3240) );
  DFFSSRX1_HVT sram_rdata_4_reg_5_ ( .D(1'b0), .SETB(n2390), .RSTB(N172), 
        .CLK(clk), .Q(sram_rdata_4[5]), .QN(n3230) );
  DFFSSRX1_HVT sram_rdata_4_reg_4_ ( .D(1'b0), .SETB(n2430), .RSTB(N171), 
        .CLK(clk), .Q(sram_rdata_4[4]), .QN(n3220) );
  DFFSSRX1_HVT sram_rdata_4_reg_3_ ( .D(1'b0), .SETB(n2840), .RSTB(N170), 
        .CLK(clk), .Q(sram_rdata_4[3]), .QN(n3210) );
  DFFSSRX1_HVT sram_rdata_4_reg_2_ ( .D(1'b0), .SETB(n2500), .RSTB(N169), 
        .CLK(clk), .Q(sram_rdata_4[2]), .QN(n3200) );
  DFFSSRX1_HVT sram_rdata_4_reg_1_ ( .D(1'b0), .SETB(n2410), .RSTB(N168), 
        .CLK(clk), .Q(sram_rdata_4[1]), .QN(n3190) );
  DFFSSRX1_HVT sram_rdata_4_reg_0_ ( .D(1'b0), .SETB(n2390), .RSTB(N167), 
        .CLK(clk), .Q(sram_rdata_4[0]), .QN(n3180) );
  DFFSSRX1_HVT sram_rdata_5_reg_31_ ( .D(1'b0), .SETB(n12100), .RSTB(N230), 
        .CLK(clk), .Q(sram_rdata_5[31]), .QN(n5401) );
  DFFSSRX1_HVT sram_rdata_5_reg_30_ ( .D(1'b0), .SETB(n13300), .RSTB(N229), 
        .CLK(clk), .Q(sram_rdata_5[30]), .QN(n539) );
  DFFSSRX1_HVT sram_rdata_5_reg_29_ ( .D(1'b0), .SETB(n12000), .RSTB(N228), 
        .CLK(clk), .Q(sram_rdata_5[29]), .QN(n538) );
  DFFSSRX1_HVT sram_rdata_5_reg_28_ ( .D(1'b0), .SETB(n2390), .RSTB(N227), 
        .CLK(clk), .Q(sram_rdata_5[28]), .QN(n537) );
  DFFSSRX1_HVT sram_rdata_5_reg_27_ ( .D(1'b0), .SETB(n2450), .RSTB(N226), 
        .CLK(clk), .Q(sram_rdata_5[27]), .QN(n536) );
  DFFSSRX1_HVT sram_rdata_5_reg_26_ ( .D(1'b0), .SETB(n2510), .RSTB(N225), 
        .CLK(clk), .Q(sram_rdata_5[26]), .QN(n535) );
  DFFSSRX1_HVT sram_rdata_5_reg_25_ ( .D(1'b0), .SETB(n2500), .RSTB(N224), 
        .CLK(clk), .Q(sram_rdata_5[25]), .QN(n534) );
  DFFSSRX1_HVT sram_rdata_5_reg_24_ ( .D(1'b0), .SETB(n2380), .RSTB(N223), 
        .CLK(clk), .Q(sram_rdata_5[24]), .QN(n533) );
  DFFSSRX1_HVT sram_rdata_5_reg_23_ ( .D(1'b0), .SETB(n2450), .RSTB(N222), 
        .CLK(clk), .Q(sram_rdata_5[23]), .QN(n532) );
  DFFSSRX1_HVT sram_rdata_5_reg_22_ ( .D(1'b0), .SETB(n2470), .RSTB(N221), 
        .CLK(clk), .Q(sram_rdata_5[22]), .QN(n531) );
  DFFSSRX1_HVT sram_rdata_5_reg_21_ ( .D(1'b0), .SETB(n2500), .RSTB(N220), 
        .CLK(clk), .Q(sram_rdata_5[21]), .QN(n5301) );
  DFFSSRX1_HVT sram_rdata_5_reg_20_ ( .D(1'b0), .SETB(n12200), .RSTB(N219), 
        .CLK(clk), .Q(sram_rdata_5[20]), .QN(n529) );
  DFFSSRX1_HVT sram_rdata_5_reg_19_ ( .D(1'b0), .SETB(n2450), .RSTB(N218), 
        .CLK(clk), .Q(sram_rdata_5[19]), .QN(n528) );
  DFFSSRX1_HVT sram_rdata_5_reg_18_ ( .D(1'b0), .SETB(n12200), .RSTB(N217), 
        .CLK(clk), .Q(sram_rdata_5[18]), .QN(n527) );
  DFFSSRX1_HVT sram_rdata_5_reg_17_ ( .D(1'b0), .SETB(n2490), .RSTB(N216), 
        .CLK(clk), .Q(sram_rdata_5[17]), .QN(n526) );
  DFFSSRX1_HVT sram_rdata_5_reg_16_ ( .D(1'b0), .SETB(n2390), .RSTB(N215), 
        .CLK(clk), .Q(sram_rdata_5[16]), .QN(n525) );
  DFFSSRX1_HVT sram_rdata_5_reg_15_ ( .D(1'b0), .SETB(n12100), .RSTB(N214), 
        .CLK(clk), .Q(sram_rdata_5[15]), .QN(n524) );
  DFFSSRX1_HVT sram_rdata_5_reg_14_ ( .D(1'b0), .SETB(n2840), .RSTB(N213), 
        .CLK(clk), .Q(sram_rdata_5[14]), .QN(n523) );
  DFFSSRX1_HVT sram_rdata_5_reg_13_ ( .D(1'b0), .SETB(n12000), .RSTB(N212), 
        .CLK(clk), .Q(sram_rdata_5[13]), .QN(n522) );
  DFFSSRX1_HVT sram_rdata_5_reg_12_ ( .D(1'b0), .SETB(n2390), .RSTB(N211), 
        .CLK(clk), .Q(sram_rdata_5[12]), .QN(n521) );
  DFFSSRX1_HVT sram_rdata_5_reg_11_ ( .D(1'b0), .SETB(n2430), .RSTB(N210), 
        .CLK(clk), .Q(sram_rdata_5[11]), .QN(n5201) );
  DFFSSRX1_HVT sram_rdata_5_reg_10_ ( .D(1'b0), .SETB(n2850), .RSTB(N209), 
        .CLK(clk), .Q(sram_rdata_5[10]), .QN(n519) );
  DFFSSRX1_HVT sram_rdata_5_reg_9_ ( .D(1'b0), .SETB(n2500), .RSTB(N208), 
        .CLK(clk), .Q(sram_rdata_5[9]), .QN(n518) );
  DFFSSRX1_HVT sram_rdata_5_reg_8_ ( .D(1'b0), .SETB(n2410), .RSTB(N207), 
        .CLK(clk), .Q(sram_rdata_5[8]), .QN(n517) );
  DFFSSRX1_HVT sram_rdata_5_reg_7_ ( .D(1'b0), .SETB(n2430), .RSTB(N206), 
        .CLK(clk), .Q(sram_rdata_5[7]), .QN(n516) );
  DFFSSRX1_HVT sram_rdata_5_reg_6_ ( .D(1'b0), .SETB(n12300), .RSTB(N205), 
        .CLK(clk), .Q(sram_rdata_5[6]), .QN(n515) );
  DFFSSRX1_HVT sram_rdata_5_reg_5_ ( .D(1'b0), .SETB(n2500), .RSTB(N204), 
        .CLK(clk), .Q(sram_rdata_5[5]), .QN(n514) );
  DFFSSRX1_HVT sram_rdata_5_reg_4_ ( .D(1'b0), .SETB(n12200), .RSTB(N203), 
        .CLK(clk), .Q(sram_rdata_5[4]), .QN(n513) );
  DFFSSRX1_HVT sram_rdata_5_reg_3_ ( .D(1'b0), .SETB(n2420), .RSTB(N202), 
        .CLK(clk), .Q(sram_rdata_5[3]), .QN(n512) );
  DFFSSRX1_HVT sram_rdata_5_reg_2_ ( .D(1'b0), .SETB(n13300), .RSTB(N201), 
        .CLK(clk), .Q(sram_rdata_5[2]), .QN(n511) );
  DFFSSRX1_HVT sram_rdata_5_reg_1_ ( .D(1'b0), .SETB(n2520), .RSTB(N200), 
        .CLK(clk), .Q(sram_rdata_5[1]), .QN(n5101) );
  DFFSSRX1_HVT sram_rdata_5_reg_0_ ( .D(1'b0), .SETB(n2500), .RSTB(N199), 
        .CLK(clk), .Q(sram_rdata_5[0]), .QN(n478) );
  DFFSSRX1_HVT sram_rdata_6_reg_31_ ( .D(1'b0), .SETB(n2380), .RSTB(N262), 
        .CLK(clk), .Q(sram_rdata_6[31]), .QN(n509) );
  DFFSSRX1_HVT sram_rdata_6_reg_30_ ( .D(1'b0), .SETB(n2430), .RSTB(N261), 
        .CLK(clk), .Q(sram_rdata_6[30]), .QN(n508) );
  DFFSSRX1_HVT sram_rdata_6_reg_29_ ( .D(1'b0), .SETB(n2850), .RSTB(N260), 
        .CLK(clk), .Q(sram_rdata_6[29]), .QN(n507) );
  DFFSSRX1_HVT sram_rdata_6_reg_28_ ( .D(1'b0), .SETB(n2490), .RSTB(N259), 
        .CLK(clk), .Q(sram_rdata_6[28]), .QN(n506) );
  DFFSSRX1_HVT sram_rdata_6_reg_27_ ( .D(1'b0), .SETB(n2380), .RSTB(N258), 
        .CLK(clk), .Q(sram_rdata_6[27]), .QN(n505) );
  DFFSSRX1_HVT sram_rdata_6_reg_26_ ( .D(1'b0), .SETB(n2430), .RSTB(N257), 
        .CLK(clk), .Q(sram_rdata_6[26]), .QN(n504) );
  DFFSSRX1_HVT sram_rdata_6_reg_25_ ( .D(1'b0), .SETB(n12300), .RSTB(N256), 
        .CLK(clk), .Q(sram_rdata_6[25]), .QN(n503) );
  DFFSSRX1_HVT sram_rdata_6_reg_24_ ( .D(1'b0), .SETB(n2490), .RSTB(N255), 
        .CLK(clk), .Q(sram_rdata_6[24]), .QN(n502) );
  DFFSSRX1_HVT sram_rdata_6_reg_23_ ( .D(1'b0), .SETB(n12200), .RSTB(N254), 
        .CLK(clk), .Q(sram_rdata_6[23]), .QN(n501) );
  DFFSSRX1_HVT sram_rdata_6_reg_22_ ( .D(1'b0), .SETB(n2450), .RSTB(N253), 
        .CLK(clk), .Q(sram_rdata_6[22]), .QN(n5001) );
  DFFSSRX1_HVT sram_rdata_6_reg_21_ ( .D(1'b0), .SETB(n2830), .RSTB(N252), 
        .CLK(clk), .Q(sram_rdata_6[21]), .QN(n499) );
  DFFSSRX1_HVT sram_rdata_6_reg_20_ ( .D(1'b0), .SETB(n2490), .RSTB(N251), 
        .CLK(clk), .Q(sram_rdata_6[20]), .QN(n498) );
  DFFSSRX1_HVT sram_rdata_6_reg_19_ ( .D(1'b0), .SETB(n2410), .RSTB(N250), 
        .CLK(clk), .Q(sram_rdata_6[19]), .QN(n497) );
  DFFSSRX1_HVT sram_rdata_6_reg_18_ ( .D(1'b0), .SETB(n12100), .RSTB(N249), 
        .CLK(clk), .Q(sram_rdata_6[18]), .QN(n496) );
  DFFSSRX1_HVT sram_rdata_6_reg_17_ ( .D(1'b0), .SETB(n2850), .RSTB(N248), 
        .CLK(clk), .Q(sram_rdata_6[17]), .QN(n495) );
  DFFSSRX1_HVT sram_rdata_6_reg_16_ ( .D(1'b0), .SETB(n13500), .RSTB(N247), 
        .CLK(clk), .Q(sram_rdata_6[16]), .QN(n494) );
  DFFSSRX1_HVT sram_rdata_6_reg_15_ ( .D(1'b0), .SETB(n2410), .RSTB(N246), 
        .CLK(clk), .Q(sram_rdata_6[15]), .QN(n493) );
  DFFSSRX1_HVT sram_rdata_6_reg_14_ ( .D(1'b0), .SETB(n2420), .RSTB(N245), 
        .CLK(clk), .Q(sram_rdata_6[14]), .QN(n492) );
  DFFSSRX1_HVT sram_rdata_6_reg_13_ ( .D(1'b0), .SETB(n2840), .RSTB(N244), 
        .CLK(clk), .Q(sram_rdata_6[13]), .QN(n491) );
  DFFSSRX1_HVT sram_rdata_6_reg_12_ ( .D(1'b0), .SETB(n2520), .RSTB(N243), 
        .CLK(clk), .Q(sram_rdata_6[12]), .QN(n4901) );
  DFFSSRX1_HVT sram_rdata_6_reg_11_ ( .D(1'b0), .SETB(n2410), .RSTB(N242), 
        .CLK(clk), .Q(sram_rdata_6[11]), .QN(n489) );
  DFFSSRX1_HVT sram_rdata_6_reg_10_ ( .D(1'b0), .SETB(n2420), .RSTB(N241), 
        .CLK(clk), .Q(sram_rdata_6[10]), .QN(n488) );
  DFFSSRX1_HVT sram_rdata_6_reg_9_ ( .D(1'b0), .SETB(n12300), .RSTB(N240), 
        .CLK(clk), .Q(sram_rdata_6[9]), .QN(n487) );
  DFFSSRX1_HVT sram_rdata_6_reg_8_ ( .D(1'b0), .SETB(n2520), .RSTB(N239), 
        .CLK(clk), .Q(sram_rdata_6[8]), .QN(n486) );
  DFFSSRX1_HVT sram_rdata_6_reg_7_ ( .D(1'b0), .SETB(n12200), .RSTB(N238), 
        .CLK(clk), .Q(sram_rdata_6[7]), .QN(n485) );
  DFFSSRX1_HVT sram_rdata_6_reg_6_ ( .D(1'b0), .SETB(n2420), .RSTB(N237), 
        .CLK(clk), .Q(sram_rdata_6[6]), .QN(n484) );
  DFFSSRX1_HVT sram_rdata_6_reg_5_ ( .D(1'b0), .SETB(n13300), .RSTB(N236), 
        .CLK(clk), .Q(sram_rdata_6[5]), .QN(n483) );
  DFFSSRX1_HVT sram_rdata_6_reg_4_ ( .D(1'b0), .SETB(n2520), .RSTB(N235), 
        .CLK(clk), .Q(sram_rdata_6[4]), .QN(n482) );
  DFFSSRX1_HVT sram_rdata_6_reg_3_ ( .D(1'b0), .SETB(n2390), .RSTB(N234), 
        .CLK(clk), .Q(sram_rdata_6[3]), .QN(n481) );
  DFFSSRX1_HVT sram_rdata_6_reg_2_ ( .D(1'b0), .SETB(n12100), .RSTB(N233), 
        .CLK(clk), .Q(sram_rdata_6[2]), .QN(n4801) );
  DFFSSRX1_HVT sram_rdata_6_reg_1_ ( .D(1'b0), .SETB(n13400), .RSTB(N232), 
        .CLK(clk), .Q(sram_rdata_6[1]), .QN(n479) );
  DFFSSRX1_HVT sram_rdata_6_reg_0_ ( .D(1'b0), .SETB(n13400), .RSTB(N231), 
        .CLK(clk), .Q(sram_rdata_6[0]), .QN(n477) );
  DFFSSRX1_HVT sram_rdata_7_reg_31_ ( .D(1'b0), .SETB(n2490), .RSTB(N294), 
        .CLK(clk), .Q(sram_rdata_7[31]), .QN(n413) );
  DFFSSRX1_HVT sram_rdata_7_reg_30_ ( .D(1'b0), .SETB(n12200), .RSTB(N293), 
        .CLK(clk), .Q(sram_rdata_7[30]), .QN(n412) );
  DFFSSRX1_HVT sram_rdata_7_reg_29_ ( .D(1'b0), .SETB(n2450), .RSTB(N292), 
        .CLK(clk), .Q(sram_rdata_7[29]), .QN(n411) );
  DFFSSRX1_HVT sram_rdata_7_reg_28_ ( .D(1'b0), .SETB(n2850), .RSTB(N291), 
        .CLK(clk), .Q(sram_rdata_7[28]), .QN(n4101) );
  DFFSSRX1_HVT sram_rdata_7_reg_27_ ( .D(1'b0), .SETB(n2490), .RSTB(N290), 
        .CLK(clk), .Q(sram_rdata_7[27]), .QN(n409) );
  DFFSSRX1_HVT sram_rdata_7_reg_26_ ( .D(1'b0), .SETB(n2410), .RSTB(N289), 
        .CLK(clk), .Q(sram_rdata_7[26]), .QN(n408) );
  DFFSSRX1_HVT sram_rdata_7_reg_25_ ( .D(1'b0), .SETB(n12100), .RSTB(N288), 
        .CLK(clk), .Q(sram_rdata_7[25]), .QN(n407) );
  DFFSSRX1_HVT sram_rdata_7_reg_24_ ( .D(1'b0), .SETB(n2830), .RSTB(N287), 
        .CLK(clk), .Q(sram_rdata_7[24]), .QN(n406) );
  DFFSSRX1_HVT sram_rdata_7_reg_23_ ( .D(1'b0), .SETB(n12000), .RSTB(N286), 
        .CLK(clk), .Q(sram_rdata_7[23]), .QN(n405) );
  DFFSSRX1_HVT sram_rdata_7_reg_22_ ( .D(1'b0), .SETB(n2410), .RSTB(N285), 
        .CLK(clk), .Q(sram_rdata_7[22]), .QN(n404) );
  DFFSSRX1_HVT sram_rdata_7_reg_21_ ( .D(1'b0), .SETB(n2420), .RSTB(N284), 
        .CLK(clk), .Q(sram_rdata_7[21]), .QN(n403) );
  DFFSSRX1_HVT sram_rdata_7_reg_20_ ( .D(1'b0), .SETB(n2850), .RSTB(N283), 
        .CLK(clk), .Q(sram_rdata_7[20]), .QN(n402) );
  DFFSSRX1_HVT sram_rdata_7_reg_19_ ( .D(1'b0), .SETB(n2520), .RSTB(N282), 
        .CLK(clk), .Q(sram_rdata_7[19]), .QN(n401) );
  DFFSSRX1_HVT sram_rdata_7_reg_18_ ( .D(1'b0), .SETB(n2410), .RSTB(N281), 
        .CLK(clk), .Q(sram_rdata_7[18]), .QN(n4001) );
  DFFSSRX1_HVT sram_rdata_7_reg_17_ ( .D(1'b0), .SETB(n2420), .RSTB(N280), 
        .CLK(clk), .Q(sram_rdata_7[17]), .QN(n399) );
  DFFSSRX1_HVT sram_rdata_7_reg_16_ ( .D(1'b0), .SETB(n12100), .RSTB(N279), 
        .CLK(clk), .Q(sram_rdata_7[16]), .QN(n398) );
  DFFSSRX1_HVT sram_rdata_7_reg_15_ ( .D(1'b0), .SETB(n2520), .RSTB(N278), 
        .CLK(clk), .Q(sram_rdata_7[15]), .QN(n397) );
  DFFSSRX1_HVT sram_rdata_7_reg_14_ ( .D(1'b0), .SETB(n12200), .RSTB(N277), 
        .CLK(clk), .Q(sram_rdata_7[14]), .QN(n396) );
  DFFSSRX1_HVT sram_rdata_7_reg_13_ ( .D(1'b0), .SETB(n2420), .RSTB(N276), 
        .CLK(clk), .Q(sram_rdata_7[13]), .QN(n395) );
  DFFSSRX1_HVT sram_rdata_7_reg_12_ ( .D(1'b0), .SETB(n2830), .RSTB(N275), 
        .CLK(clk), .Q(sram_rdata_7[12]), .QN(n394) );
  DFFSSRX1_HVT sram_rdata_7_reg_11_ ( .D(1'b0), .SETB(n2520), .RSTB(N274), 
        .CLK(clk), .Q(sram_rdata_7[11]), .QN(n393) );
  DFFSSRX1_HVT sram_rdata_7_reg_10_ ( .D(1'b0), .SETB(n2390), .RSTB(N273), 
        .CLK(clk), .Q(sram_rdata_7[10]), .QN(n392) );
  DFFSSRX1_HVT sram_rdata_7_reg_9_ ( .D(1'b0), .SETB(n12100), .RSTB(N272), 
        .CLK(clk), .Q(sram_rdata_7[9]), .QN(n391) );
  DFFSSRX1_HVT sram_rdata_7_reg_8_ ( .D(1'b0), .SETB(n2440), .RSTB(N271), 
        .CLK(clk), .Q(sram_rdata_7[8]), .QN(n3901) );
  DFFSSRX1_HVT sram_rdata_7_reg_7_ ( .D(1'b0), .SETB(n12000), .RSTB(N270), 
        .CLK(clk), .Q(sram_rdata_7[7]), .QN(n389) );
  DFFSSRX1_HVT sram_rdata_7_reg_6_ ( .D(1'b0), .SETB(n2390), .RSTB(N269), 
        .CLK(clk), .Q(sram_rdata_7[6]), .QN(n388) );
  DFFSSRX1_HVT sram_rdata_7_reg_5_ ( .D(1'b0), .SETB(n2450), .RSTB(N268), 
        .CLK(clk), .Q(sram_rdata_7[5]), .QN(n387) );
  DFFSSRX1_HVT sram_rdata_7_reg_4_ ( .D(1'b0), .SETB(n2400), .RSTB(N267), 
        .CLK(clk), .Q(sram_rdata_7[4]), .QN(n386) );
  DFFSSRX1_HVT sram_rdata_7_reg_3_ ( .D(1'b0), .SETB(n2500), .RSTB(N266), 
        .CLK(clk), .Q(sram_rdata_7[3]), .QN(n385) );
  DFFSSRX1_HVT sram_rdata_7_reg_2_ ( .D(1'b0), .SETB(n2380), .RSTB(N265), 
        .CLK(clk), .Q(sram_rdata_7[2]), .QN(n384) );
  DFFSSRX1_HVT sram_rdata_7_reg_1_ ( .D(1'b0), .SETB(n2450), .RSTB(N264), 
        .CLK(clk), .Q(sram_rdata_7[1]), .QN(n383) );
  DFFSSRX1_HVT sram_rdata_7_reg_0_ ( .D(1'b0), .SETB(n12100), .RSTB(N263), 
        .CLK(clk), .Q(sram_rdata_7[0]), .QN(n2860) );
  AO221X1_HVT U3 ( .A1(1'b1), .A2(n9400), .A3(sram_rdata_1[31]), .A4(n1760), 
        .A5(n9500), .Y(n_src_aox[287]) );
  AO221X1_HVT U4 ( .A1(1'b1), .A2(n9200), .A3(sram_rdata_2[21]), .A4(n1710), 
        .A5(n9300), .Y(n_src_aox[261]) );
  AO221X1_HVT U5 ( .A1(1'b1), .A2(n8900), .A3(sram_rdata_1[30]), .A4(n1730), 
        .A5(n9000), .Y(n_src_aox[286]) );
  AO221X1_HVT U6 ( .A1(1'b1), .A2(n8600), .A3(sram_rdata_1[20]), .A4(n575), 
        .A5(n8700), .Y(n_src_aox[276]) );
  AO221X1_HVT U7 ( .A1(1'b1), .A2(n8300), .A3(sram_rdata_1[28]), .A4(n1700), 
        .A5(n8400), .Y(n_src_aox[284]) );
  AO221X1_HVT U8 ( .A1(1'b1), .A2(n8000), .A3(sram_rdata_1[27]), .A4(n1770), 
        .A5(n8100), .Y(n_src_aox[283]) );
  AO221X1_HVT U9 ( .A1(1'b1), .A2(n7700), .A3(sram_rdata_1[24]), .A4(n575), 
        .A5(n7800), .Y(n_src_aox[280]) );
  AO221X1_HVT U10 ( .A1(1'b1), .A2(n7400), .A3(sram_rdata_5[30]), .A4(n2240), 
        .A5(n7500), .Y(n_src_aox[174]) );
  AO221X1_HVT U11 ( .A1(1'b1), .A2(n7100), .A3(sram_rdata_1[23]), .A4(n1800), 
        .A5(n7200), .Y(n_src_aox[279]) );
  AO221X1_HVT U12 ( .A1(1'b1), .A2(n6800), .A3(sram_rdata_0[2]), .A4(n578), 
        .A5(n6900), .Y(n_src_aox[194]) );
  AO221X1_HVT U13 ( .A1(1'b1), .A2(n6500), .A3(sram_rdata_1[18]), .A4(n2250), 
        .A5(n6600), .Y(n_src_aox[274]) );
  AO221X1_HVT U14 ( .A1(1'b1), .A2(n6200), .A3(sram_rdata_0[27]), .A4(n1740), 
        .A5(n6300), .Y(n_src_aox[251]) );
  AO221X1_HVT U15 ( .A1(1'b1), .A2(n5900), .A3(sram_rdata_2[28]), .A4(n1740), 
        .A5(n6000), .Y(n_src_aox[268]) );
  AO221X1_HVT U16 ( .A1(1'b1), .A2(n5600), .A3(sram_rdata_2[26]), .A4(n1710), 
        .A5(n5700), .Y(n_src_aox[266]) );
  AO221X1_HVT U17 ( .A1(1'b1), .A2(n5300), .A3(sram_rdata_2[27]), .A4(n2260), 
        .A5(n5400), .Y(n_src_aox[267]) );
  AO221X1_HVT U18 ( .A1(1'b1), .A2(n5000), .A3(sram_rdata_2[5]), .A4(n1730), 
        .A5(n5100), .Y(n_src_aox[213]) );
  AO221X1_HVT U19 ( .A1(1'b1), .A2(n4700), .A3(sram_rdata_2[24]), .A4(n2220), 
        .A5(n4800), .Y(n_src_aox[264]) );
  AO221X1_HVT U20 ( .A1(1'b1), .A2(n4400), .A3(sram_rdata_4[26]), .A4(n2250), 
        .A5(n4500), .Y(n_src_aox[186]) );
  AO221X1_HVT U21 ( .A1(1'b1), .A2(n4100), .A3(sram_rdata_2[22]), .A4(n1710), 
        .A5(n4200), .Y(n_src_aox[262]) );
  AO221X1_HVT U22 ( .A1(1'b1), .A2(n38), .A3(sram_rdata_4[28]), .A4(n2250), 
        .A5(n3900), .Y(n_src_aox[188]) );
  AO221X1_HVT U23 ( .A1(1'b1), .A2(n35), .A3(sram_rdata_2[17]), .A4(n1800), 
        .A5(n36), .Y(n_src_aox[257]) );
  AO221X1_HVT U24 ( .A1(1'b1), .A2(n32), .A3(sram_rdata_4[27]), .A4(n577), 
        .A5(n33), .Y(n_src_aox[187]) );
  AO221X1_HVT U25 ( .A1(1'b1), .A2(n29), .A3(sram_rdata_2[16]), .A4(n574), 
        .A5(n30), .Y(n_src_aox[256]) );
  AO221X1_HVT U26 ( .A1(1'b1), .A2(n26), .A3(sram_rdata_2[14]), .A4(n2260), 
        .A5(n27), .Y(n_src_aox[222]) );
  AO221X1_HVT U27 ( .A1(1'b1), .A2(n23), .A3(sram_rdata_0[29]), .A4(n2270), 
        .A5(n24), .Y(n_src_aox[253]) );
  AO221X1_HVT U28 ( .A1(1'b1), .A2(n20), .A3(sram_rdata_0[0]), .A4(n1740), 
        .A5(n21), .Y(n_src_aox[192]) );
  AO221X1_HVT U29 ( .A1(1'b1), .A2(n17), .A3(sram_rdata_0[20]), .A4(n576), 
        .A5(n18), .Y(n_src_aox[244]) );
  AO221X1_HVT U30 ( .A1(1'b1), .A2(n14), .A3(sram_rdata_1[14]), .A4(n2250), 
        .A5(n15), .Y(n_src_aox[238]) );
  AO221X1_HVT U31 ( .A1(1'b1), .A2(n11), .A3(sram_rdata_1[6]), .A4(n575), .A5(
        n12), .Y(n_src_aox[230]) );
  AO221X1_HVT U32 ( .A1(1'b1), .A2(n8), .A3(sram_rdata_1[0]), .A4(n2270), .A5(
        n9), .Y(n_src_aox[224]) );
  AO221X1_HVT U33 ( .A1(1'b1), .A2(n5), .A3(sram_rdata_1[3]), .A4(n2260), .A5(
        n6), .Y(n_src_aox[227]) );
  AO221X1_HVT U34 ( .A1(1'b1), .A2(n2), .A3(sram_rdata_5[29]), .A4(n2220), 
        .A5(n3), .Y(n_src_aox[173]) );
  INVX1_HVT U35 ( .A(n584), .Y(n10200) );
  INVX1_HVT U36 ( .A(n585), .Y(n10300) );
  NBUFFX2_HVT U37 ( .A(n1655), .Y(n2210) );
  AO22X1_HVT U39 ( .A1(n1583), .A2(n12400), .A3(n593), .A4(n1194), .Y(n2) );
  OAI22X1_HVT U40 ( .A1(n2690), .A2(n347), .A3(n10400), .A4(n442), .Y(n3) );
  AO22X1_HVT U42 ( .A1(n1415), .A2(n10900), .A3(n11100), .A4(n1416), .Y(n5) );
  OAI22X1_HVT U43 ( .A1(n14900), .A2(n448), .A3(n2780), .A4(n544), .Y(n6) );
  AO22X1_HVT U45 ( .A1(n1403), .A2(n11100), .A3(n5901), .A4(n1404), .Y(n8) );
  OAI22X1_HVT U46 ( .A1(n14800), .A2(n445), .A3(n10400), .A4(n541), .Y(n9) );
  AO22X1_HVT U48 ( .A1(n1427), .A2(n12700), .A3(n11000), .A4(n1428), .Y(n11)
         );
  OAI22X1_HVT U49 ( .A1(n2700), .A2(n451), .A3(n11800), .A4(n547), .Y(n12) );
  AO22X1_HVT U51 ( .A1(n1464), .A2(n10800), .A3(n13000), .A4(n1465), .Y(n14)
         );
  OAI22X1_HVT U52 ( .A1(n2710), .A2(n459), .A3(n2770), .A4(n555), .Y(n15) );
  AO22X1_HVT U54 ( .A1(n1491), .A2(n12800), .A3(n14400), .A4(n1492), .Y(n17)
         );
  OAI22X1_HVT U55 ( .A1(n2720), .A2(n561), .A3(n2800), .A4(n370), .Y(n18) );
  AO22X1_HVT U57 ( .A1(n1255), .A2(n12900), .A3(n10900), .A4(n1256), .Y(n20)
         );
  OAI22X1_HVT U58 ( .A1(n2750), .A2(n541), .A3(n11600), .A4(n350), .Y(n21) );
  AO22X1_HVT U60 ( .A1(n15301), .A2(n12700), .A3(n12900), .A4(n1531), .Y(n23)
         );
  OAI22X1_HVT U61 ( .A1(n14700), .A2(n5701), .A3(n10400), .A4(n379), .Y(n24)
         );
  AO22X1_HVT U63 ( .A1(n1396), .A2(n10900), .A3(n13000), .A4(n1397), .Y(n26)
         );
  OAI22X1_HVT U64 ( .A1(n14600), .A2(n364), .A3(n2780), .A4(n459), .Y(n27) );
  AO22X1_HVT U66 ( .A1(n1542), .A2(n10800), .A3(n10700), .A4(n1543), .Y(n29)
         );
  OAI22X1_HVT U67 ( .A1(n2720), .A2(n366), .A3(n10400), .A4(n461), .Y(n30) );
  AO22X1_HVT U69 ( .A1(n1641), .A2(n583), .A3(n10800), .A4(n1241), .Y(n32) );
  OAI22X1_HVT U70 ( .A1(n1662), .A2(n4401), .A3(n11800), .A4(n536), .Y(n33) );
  AO22X1_HVT U72 ( .A1(n1544), .A2(n10900), .A3(n14400), .A4(n1545), .Y(n35)
         );
  OAI22X1_HVT U73 ( .A1(n2700), .A2(n367), .A3(n10300), .A4(n462), .Y(n36) );
  AO22X1_HVT U75 ( .A1(n1643), .A2(n13000), .A3(n15100), .A4(n1242), .Y(n38)
         );
  OAI22X1_HVT U76 ( .A1(n14900), .A2(n441), .A3(n10300), .A4(n537), .Y(n3900)
         );
  AO22X1_HVT U78 ( .A1(n1563), .A2(n12800), .A3(n10700), .A4(n1564), .Y(n4100)
         );
  OAI22X1_HVT U79 ( .A1(n14700), .A2(n372), .A3(n10200), .A4(n467), .Y(n4200)
         );
  AO22X1_HVT U81 ( .A1(n1636), .A2(n12400), .A3(n592), .A4(n12401), .Y(n4400)
         );
  OAI22X1_HVT U82 ( .A1(n2700), .A2(n439), .A3(n2760), .A4(n535), .Y(n4500) );
  AO22X1_HVT U84 ( .A1(n15701), .A2(n12700), .A3(n10700), .A4(n1571), .Y(n4700) );
  OAI22X1_HVT U85 ( .A1(n2750), .A2(n374), .A3(n13900), .A4(n469), .Y(n4800)
         );
  AO22X1_HVT U87 ( .A1(n1354), .A2(n10800), .A3(n13000), .A4(n1355), .Y(n5000)
         );
  OAI22X1_HVT U88 ( .A1(n2710), .A2(n355), .A3(n2790), .A4(n4501), .Y(n5100)
         );
  AO22X1_HVT U90 ( .A1(n1579), .A2(n10900), .A3(n12400), .A4(n15801), .Y(n5300) );
  OAI22X1_HVT U91 ( .A1(n14900), .A2(n377), .A3(n10200), .A4(n472), .Y(n5400)
         );
  AO22X1_HVT U93 ( .A1(n1577), .A2(n10900), .A3(n10700), .A4(n1578), .Y(n5600)
         );
  OAI22X1_HVT U94 ( .A1(n10100), .A2(n376), .A3(n2760), .A4(n471), .Y(n5700)
         );
  AO22X1_HVT U96 ( .A1(n1581), .A2(n10800), .A3(n13000), .A4(n1582), .Y(n5900)
         );
  OAI22X1_HVT U97 ( .A1(n2730), .A2(n378), .A3(n11700), .A4(n473), .Y(n6000)
         );
  AO22X1_HVT U99 ( .A1(n1523), .A2(n10900), .A3(n12400), .A4(n1524), .Y(n6200)
         );
  OAI22X1_HVT U100 ( .A1(n1662), .A2(n568), .A3(n11800), .A4(n377), .Y(n6300)
         );
  AO22X1_HVT U102 ( .A1(n1608), .A2(n12800), .A3(n14400), .A4(n1609), .Y(n6500) );
  OAI22X1_HVT U103 ( .A1(n2690), .A2(n463), .A3(n13900), .A4(n559), .Y(n6600)
         );
  AO22X1_HVT U105 ( .A1(n1262), .A2(n12800), .A3(n13000), .A4(n1263), .Y(n6800) );
  OAI22X1_HVT U106 ( .A1(n2700), .A2(n543), .A3(n13900), .A4(n352), .Y(n6900)
         );
  AO22X1_HVT U108 ( .A1(n1627), .A2(n10900), .A3(n12900), .A4(n1628), .Y(n7100) );
  OAI22X1_HVT U109 ( .A1(n14900), .A2(n468), .A3(n2760), .A4(n564), .Y(n7200)
         );
  AO22X1_HVT U111 ( .A1(n1588), .A2(n12900), .A3(n1664), .A4(n1195), .Y(n7400)
         );
  OAI22X1_HVT U112 ( .A1(n2700), .A2(n348), .A3(n2780), .A4(n443), .Y(n7500)
         );
  AO22X1_HVT U114 ( .A1(n1629), .A2(n10800), .A3(n13000), .A4(n16301), .Y(
        n7700) );
  OAI22X1_HVT U115 ( .A1(n2740), .A2(n469), .A3(n2790), .A4(n565), .Y(n7800)
         );
  AO22X1_HVT U117 ( .A1(n1641), .A2(n12700), .A3(n13000), .A4(n1642), .Y(n8000) );
  OAI22X1_HVT U118 ( .A1(n2740), .A2(n472), .A3(n10200), .A4(n568), .Y(n8100)
         );
  AO22X1_HVT U120 ( .A1(n1643), .A2(n12700), .A3(n10700), .A4(n1644), .Y(n8300) );
  OAI22X1_HVT U121 ( .A1(n10000), .A2(n473), .A3(n10300), .A4(n569), .Y(n8400)
         );
  AO22X1_HVT U123 ( .A1(n1615), .A2(n594), .A3(n583), .A4(n1616), .Y(n8600) );
  OAI22X1_HVT U124 ( .A1(n2720), .A2(n465), .A3(n2800), .A4(n561), .Y(n8700)
         );
  AO22X1_HVT U126 ( .A1(n16501), .A2(n12800), .A3(n12400), .A4(n1651), .Y(
        n8900) );
  OAI22X1_HVT U127 ( .A1(n14600), .A2(n475), .A3(n2770), .A4(n571), .Y(n9000)
         );
  AO22X1_HVT U129 ( .A1(n1561), .A2(n5901), .A3(n11100), .A4(n1562), .Y(n9200)
         );
  OAI22X1_HVT U130 ( .A1(n11400), .A2(n371), .A3(n13800), .A4(n466), .Y(n9300)
         );
  AO22X1_HVT U131 ( .A1(n1652), .A2(n592), .A3(n581), .A4(n1654), .Y(n9400) );
  OAI22X1_HVT U132 ( .A1(n2740), .A2(n476), .A3(n13600), .A4(n572), .Y(n9500)
         );
  NAND2X0_HVT U134 ( .A1(box_sel[1]), .A2(n1659), .Y(n9700) );
  NAND2X0_HVT U135 ( .A1(mode[1]), .A2(n1665), .Y(n1666) );
  INVX1_HVT U136 ( .A(n1661), .Y(n11200) );
  INVX2_HVT U137 ( .A(n2530), .Y(n9800) );
  INVX2_HVT U138 ( .A(n2570), .Y(n9900) );
  INVX2_HVT U139 ( .A(n587), .Y(n10000) );
  INVX1_HVT U140 ( .A(n585), .Y(n11700) );
  INVX1_HVT U141 ( .A(n584), .Y(n11800) );
  INVX2_HVT U142 ( .A(n587), .Y(n10100) );
  INVX1_HVT U143 ( .A(n584), .Y(n11600) );
  INVX0_HVT U144 ( .A(n584), .Y(n13600) );
  INVX0_HVT U145 ( .A(n585), .Y(n13800) );
  INVX1_HVT U146 ( .A(n14100), .Y(n11900) );
  INVX0_HVT U147 ( .A(n585), .Y(n13900) );
  INVX1_HVT U148 ( .A(n586), .Y(n2750) );
  INVX0_HVT U149 ( .A(n584), .Y(n13700) );
  INVX2_HVT U150 ( .A(n585), .Y(n10400) );
  INVX2_HVT U151 ( .A(n14100), .Y(n10500) );
  INVX2_HVT U152 ( .A(n1662), .Y(n587) );
  INVX1_HVT U153 ( .A(n1662), .Y(n586) );
  INVX2_HVT U154 ( .A(n14100), .Y(n10600) );
  INVX2_HVT U155 ( .A(n14500), .Y(n10700) );
  INVX2_HVT U156 ( .A(n15200), .Y(n10800) );
  INVX2_HVT U157 ( .A(n15200), .Y(n10900) );
  INVX2_HVT U158 ( .A(n15300), .Y(n11000) );
  INVX2_HVT U159 ( .A(n15300), .Y(n11100) );
  INVX1_HVT U160 ( .A(srstn), .Y(n2850) );
  INVX1_HVT U161 ( .A(srstn), .Y(n2840) );
  INVX1_HVT U162 ( .A(srstn), .Y(n2830) );
  INVX1_HVT U163 ( .A(n2570), .Y(n13200) );
  INVX1_HVT U164 ( .A(n2570), .Y(n13100) );
  INVX2_HVT U165 ( .A(n2570), .Y(n11300) );
  INVX2_HVT U166 ( .A(n587), .Y(n11400) );
  INVX2_HVT U167 ( .A(n2530), .Y(n11500) );
  INVX1_HVT U168 ( .A(n2530), .Y(n2560) );
  INVX2_HVT U169 ( .A(n587), .Y(n2710) );
  INVX2_HVT U170 ( .A(n586), .Y(n2740) );
  INVX1_HVT U171 ( .A(N346), .Y(n2570) );
  INVX1_HVT U172 ( .A(n579), .Y(n2530) );
  INVX1_HVT U173 ( .A(n15800), .Y(n15700) );
  INVX1_HVT U174 ( .A(n15800), .Y(n15600) );
  INVX0_HVT U175 ( .A(n595), .Y(n2620) );
  INVX0_HVT U176 ( .A(n2640), .Y(n2670) );
  INVX1_HVT U177 ( .A(n15800), .Y(n15500) );
  INVX1_HVT U178 ( .A(n15800), .Y(n15400) );
  INVX1_HVT U179 ( .A(n2460), .Y(n13400) );
  INVX1_HVT U180 ( .A(n2480), .Y(n13300) );
  INVX1_HVT U181 ( .A(n2370), .Y(n13500) );
  INVX1_HVT U182 ( .A(n1663), .Y(n584) );
  INVX1_HVT U183 ( .A(n1663), .Y(n585) );
  INVX1_HVT U184 ( .A(n1850), .Y(n1870) );
  INVX1_HVT U185 ( .A(n1850), .Y(n1890) );
  INVX1_HVT U186 ( .A(n1850), .Y(n1860) );
  INVX1_HVT U187 ( .A(n1850), .Y(n1880) );
  INVX1_HVT U188 ( .A(n1667), .Y(n2640) );
  INVX2_HVT U189 ( .A(n2480), .Y(n12000) );
  INVX2_HVT U190 ( .A(n2460), .Y(n12100) );
  INVX2_HVT U191 ( .A(n2460), .Y(n12200) );
  INVX2_HVT U192 ( .A(n2460), .Y(n12300) );
  NAND3X0_HVT U193 ( .A1(n1657), .A2(n1656), .A3(n2070), .Y(n1662) );
  INVX1_HVT U194 ( .A(n15800), .Y(n16200) );
  INVX1_HVT U195 ( .A(n15800), .Y(n15900) );
  INVX1_HVT U196 ( .A(n1667), .Y(n595) );
  INVX1_HVT U197 ( .A(n15800), .Y(n16000) );
  INVX1_HVT U198 ( .A(n15800), .Y(n16100) );
  INVX1_HVT U199 ( .A(n14000), .Y(n1850) );
  INVX1_HVT U200 ( .A(n1720), .Y(n1790) );
  INVX1_HVT U201 ( .A(n2230), .Y(n1800) );
  INVX1_HVT U202 ( .A(n1940), .Y(n2010) );
  INVX1_HVT U203 ( .A(n9700), .Y(n1680) );
  INVX1_HVT U204 ( .A(n9700), .Y(n1910) );
  INVX1_HVT U205 ( .A(n9700), .Y(n1900) );
  INVX1_HVT U206 ( .A(n11200), .Y(n2070) );
  INVX1_HVT U207 ( .A(n2230), .Y(n2240) );
  INVX1_HVT U208 ( .A(n1720), .Y(n1730) );
  INVX1_HVT U209 ( .A(n1940), .Y(n2020) );
  INVX1_HVT U210 ( .A(n1720), .Y(n1740) );
  INVX1_HVT U211 ( .A(n9700), .Y(n1920) );
  INVX1_HVT U212 ( .A(n1940), .Y(n1980) );
  INVX1_HVT U213 ( .A(n9700), .Y(n1930) );
  INVX1_HVT U214 ( .A(n1940), .Y(n1970) );
  INVX1_HVT U215 ( .A(n2230), .Y(n2250) );
  INVX1_HVT U216 ( .A(n1720), .Y(n1780) );
  INVX1_HVT U217 ( .A(n1940), .Y(n2000) );
  INVX1_HVT U218 ( .A(n1940), .Y(n1960) );
  INVX1_HVT U219 ( .A(n11200), .Y(n14000) );
  INVX1_HVT U220 ( .A(n2230), .Y(n2260) );
  INVX1_HVT U221 ( .A(n1720), .Y(n1760) );
  INVX1_HVT U222 ( .A(n9700), .Y(n1990) );
  INVX1_HVT U223 ( .A(n1720), .Y(n1750) );
  INVX1_HVT U224 ( .A(n1940), .Y(n1950) );
  INVX1_HVT U225 ( .A(n9700), .Y(n16600) );
  INVX1_HVT U226 ( .A(n9700), .Y(n16400) );
  INVX1_HVT U227 ( .A(n9700), .Y(n16300) );
  INVX2_HVT U228 ( .A(n14500), .Y(n12400) );
  INVX1_HVT U229 ( .A(n9700), .Y(n1670) );
  INVX1_HVT U230 ( .A(n9700), .Y(n16500) );
  INVX1_HVT U231 ( .A(n2130), .Y(n15800) );
  INVX1_HVT U232 ( .A(n2230), .Y(n1770) );
  INVX1_HVT U233 ( .A(n2230), .Y(n2270) );
  NAND3X0_HVT U234 ( .A1(n1657), .A2(n1656), .A3(n2170), .Y(n1663) );
  INVX1_HVT U235 ( .A(n1940), .Y(n1690) );
  INVX1_HVT U236 ( .A(n2830), .Y(n2370) );
  INVX1_HVT U237 ( .A(n2850), .Y(n2480) );
  INVX1_HVT U238 ( .A(n2840), .Y(n2460) );
  INVX2_HVT U239 ( .A(n15300), .Y(n12500) );
  INVX1_HVT U240 ( .A(n2120), .Y(n2130) );
  INVX1_HVT U241 ( .A(n2120), .Y(n2160) );
  INVX1_HVT U242 ( .A(n1700), .Y(n1720) );
  INVX1_HVT U243 ( .A(n1900), .Y(n1940) );
  INVX1_HVT U244 ( .A(n2120), .Y(n2140) );
  INVX1_HVT U245 ( .A(n11200), .Y(n12600) );
  INVX2_HVT U246 ( .A(n15200), .Y(n12700) );
  INVX1_HVT U247 ( .A(n2120), .Y(n2170) );
  INVX2_HVT U248 ( .A(n15200), .Y(n12800) );
  INVX1_HVT U249 ( .A(n15300), .Y(n14400) );
  INVX1_HVT U250 ( .A(n2120), .Y(n2150) );
  INVX2_HVT U251 ( .A(n15300), .Y(n12900) );
  INVX1_HVT U252 ( .A(n575), .Y(n2230) );
  DELLN1X2_HVT U253 ( .A(n1655), .Y(n577) );
  DELLN1X2_HVT U254 ( .A(n1653), .Y(n5801) );
  INVX2_HVT U255 ( .A(n15300), .Y(n13000) );
  INVX1_HVT U256 ( .A(n589), .Y(n2120) );
  DELLN1X2_HVT U257 ( .A(n1653), .Y(n582) );
  NBUFFX2_HVT U258 ( .A(n1653), .Y(n581) );
  DELLN1X2_HVT U259 ( .A(n1664), .Y(n593) );
  NBUFFX2_HVT U260 ( .A(n1666), .Y(n2820) );
  DELLN1X2_HVT U261 ( .A(n1653), .Y(n583) );
  DELLN1X2_HVT U262 ( .A(n1655), .Y(n578) );
  NBUFFX2_HVT U263 ( .A(n16601), .Y(n589) );
  INVX2_HVT U264 ( .A(n2370), .Y(n2390) );
  INVX1_HVT U265 ( .A(n2370), .Y(n2400) );
  INVX2_HVT U266 ( .A(srstn), .Y(n2430) );
  INVX1_HVT U267 ( .A(srstn), .Y(n2440) );
  INVX1_HVT U268 ( .A(n2460), .Y(n2470) );
  INVX2_HVT U269 ( .A(n2480), .Y(n2500) );
  INVX1_HVT U270 ( .A(n2480), .Y(n2510) );
  DELLN1X2_HVT U271 ( .A(n16601), .Y(n588) );
  DELLN1X2_HVT U272 ( .A(n16601), .Y(n2110) );
  DELLN1X2_HVT U273 ( .A(n1664), .Y(n591) );
  DELLN1X2_HVT U274 ( .A(n1664), .Y(n592) );
  DELLN1X2_HVT U275 ( .A(n1664), .Y(n594) );
  DELLN1X2_HVT U276 ( .A(n1664), .Y(n5901) );
  DELLN1X2_HVT U277 ( .A(n1664), .Y(n15100) );
  DELLN1X2_HVT U278 ( .A(n1664), .Y(n15000) );
  INVX2_HVT U279 ( .A(n2530), .Y(n2550) );
  INVX2_HVT U280 ( .A(n2530), .Y(n2540) );
  INVX2_HVT U281 ( .A(n2570), .Y(n2590) );
  INVX2_HVT U282 ( .A(n2570), .Y(n2580) );
  NBUFFX2_HVT U283 ( .A(N346), .Y(n579) );
  INVX2_HVT U284 ( .A(n595), .Y(n2630) );
  INVX2_HVT U285 ( .A(n595), .Y(n2610) );
  INVX2_HVT U286 ( .A(n595), .Y(n2600) );
  INVX0_HVT U287 ( .A(n2620), .Y(n14100) );
  INVX2_HVT U288 ( .A(n2640), .Y(n14200) );
  INVX2_HVT U289 ( .A(n2640), .Y(n14300) );
  INVX2_HVT U290 ( .A(n2640), .Y(n2680) );
  INVX2_HVT U291 ( .A(n2640), .Y(n2660) );
  INVX2_HVT U292 ( .A(n2640), .Y(n2650) );
  DELLN1X2_HVT U293 ( .A(n1655), .Y(n575) );
  DELLN1X2_HVT U294 ( .A(n1655), .Y(n574) );
  DELLN1X2_HVT U295 ( .A(n1655), .Y(n576) );
  DELLN1X2_HVT U296 ( .A(n1655), .Y(n2220) );
  DELLN1X2_HVT U297 ( .A(n1655), .Y(n1710) );
  DELLN1X2_HVT U298 ( .A(n1655), .Y(n1700) );
  INVX0_HVT U299 ( .A(n14400), .Y(n14500) );
  INVX2_HVT U300 ( .A(n587), .Y(n14600) );
  INVX2_HVT U301 ( .A(n587), .Y(n14700) );
  INVX2_HVT U302 ( .A(n587), .Y(n2700) );
  INVX2_HVT U303 ( .A(n587), .Y(n2690) );
  INVX2_HVT U304 ( .A(n586), .Y(n14800) );
  INVX2_HVT U305 ( .A(n586), .Y(n14900) );
  INVX2_HVT U306 ( .A(n586), .Y(n2730) );
  INVX2_HVT U307 ( .A(n586), .Y(n2720) );
  INVX0_HVT U308 ( .A(n15100), .Y(n15200) );
  INVX0_HVT U309 ( .A(n581), .Y(n15300) );
  INVX1_HVT U310 ( .A(n584), .Y(n2770) );
  INVX1_HVT U311 ( .A(n584), .Y(n2780) );
  INVX1_HVT U312 ( .A(n584), .Y(n2760) );
  INVX1_HVT U313 ( .A(n585), .Y(n2800) );
  INVX1_HVT U314 ( .A(n585), .Y(n2810) );
  INVX1_HVT U315 ( .A(n585), .Y(n2790) );
  INVX0_HVT U316 ( .A(n11200), .Y(n1810) );
  INVX0_HVT U317 ( .A(n11200), .Y(n1820) );
  INVX0_HVT U318 ( .A(n11200), .Y(n1830) );
  INVX0_HVT U319 ( .A(n11200), .Y(n1840) );
  INVX0_HVT U320 ( .A(n11200), .Y(n2030) );
  INVX0_HVT U321 ( .A(n11200), .Y(n2040) );
  INVX0_HVT U322 ( .A(n11200), .Y(n2050) );
  INVX0_HVT U323 ( .A(n11200), .Y(n2060) );
  INVX0_HVT U324 ( .A(n1850), .Y(n2080) );
  INVX0_HVT U325 ( .A(n1850), .Y(n2090) );
  INVX0_HVT U326 ( .A(n1850), .Y(n2100) );
  INVX0_HVT U327 ( .A(n15800), .Y(n2180) );
  INVX0_HVT U328 ( .A(n15800), .Y(n2190) );
  INVX0_HVT U329 ( .A(n15800), .Y(n2200) );
  INVX2_HVT U330 ( .A(n2600), .Y(n2280) );
  INVX2_HVT U331 ( .A(n2610), .Y(n2290) );
  INVX2_HVT U332 ( .A(n2630), .Y(n2300) );
  INVX2_HVT U333 ( .A(n2680), .Y(n2310) );
  INVX2_HVT U334 ( .A(n10600), .Y(n2320) );
  INVX2_HVT U335 ( .A(n10600), .Y(n2330) );
  INVX2_HVT U336 ( .A(n2660), .Y(n2340) );
  INVX2_HVT U337 ( .A(n10500), .Y(n2350) );
  INVX2_HVT U338 ( .A(n10600), .Y(n2360) );
  INVX2_HVT U339 ( .A(n2370), .Y(n2380) );
  INVX2_HVT U340 ( .A(n2370), .Y(n2410) );
  INVX2_HVT U341 ( .A(srstn), .Y(n2420) );
  INVX2_HVT U342 ( .A(srstn), .Y(n2450) );
  INVX2_HVT U343 ( .A(n2480), .Y(n2490) );
  INVX2_HVT U344 ( .A(n2480), .Y(n2520) );
  INVX1_HVT U345 ( .A(n2820), .Y(n1667) );
  INVX1_HVT U346 ( .A(mode[0]), .Y(n1665) );
  INVX1_HVT U347 ( .A(box_sel[1]), .Y(n1658) );
  INVX1_HVT U348 ( .A(box_sel[2]), .Y(n1657) );
  INVX1_HVT U349 ( .A(box_sel[3]), .Y(n1656) );
  INVX1_HVT U350 ( .A(box_sel[0]), .Y(n1659) );
  NAND2X0_HVT U351 ( .A1(n1655), .A2(n1658), .Y(n596) );
  AND3X1_HVT U352 ( .A1(n1659), .A2(n1656), .A3(n1657), .Y(n1655) );
  NAND2X0_HVT U353 ( .A1(srstn), .A2(n596), .Y(N346) );
  AO222X1_HVT U354 ( .A1(n1810), .A2(sram_rdata_5[0]), .A3(n2000), .A4(
        sram_rdata_3[0]), .A5(n2110), .A6(sram_rdata_4[0]), .Y(n1255) );
  AND2X1_HVT U355 ( .A1(n1656), .A2(box_sel[2]), .Y(n1653) );
  AO222X1_HVT U356 ( .A1(n2050), .A2(sram_rdata_2[0]), .A3(n15500), .A4(
        sram_rdata_1[0]), .A5(sram_rdata_0[0]), .A6(n1920), .Y(n886) );
  AOI22X1_HVT U357 ( .A1(n1255), .A2(n12700), .A3(n12500), .A4(n886), .Y(n599)
         );
  OA22X1_HVT U358 ( .A1(n2800), .A2(n2860), .A3(n2690), .A4(n573), .Y(n598) );
  NAND2X0_HVT U359 ( .A1(n1760), .A2(sram_rdata_6[0]), .Y(n597) );
  NAND3X0_HVT U360 ( .A1(n599), .A2(n598), .A3(n597), .Y(n_src_aox[0]) );
  AO222X1_HVT U361 ( .A1(n12600), .A2(sram_rdata_5[1]), .A3(n2200), .A4(
        sram_rdata_4[1]), .A5(sram_rdata_3[1]), .A6(n16500), .Y(n1258) );
  AO222X1_HVT U362 ( .A1(n1820), .A2(sram_rdata_2[1]), .A3(n2130), .A4(
        sram_rdata_1[1]), .A5(sram_rdata_0[1]), .A6(n16300), .Y(n8901) );
  AOI22X1_HVT U363 ( .A1(n1258), .A2(n591), .A3(n11100), .A4(n8901), .Y(n602)
         );
  OA22X1_HVT U364 ( .A1(n11700), .A2(n383), .A3(n14800), .A4(n2870), .Y(n601)
         );
  NAND2X0_HVT U365 ( .A1(n2270), .A2(sram_rdata_6[1]), .Y(n6001) );
  NAND3X0_HVT U366 ( .A1(n602), .A2(n601), .A3(n6001), .Y(n_src_aox[1]) );
  AO222X1_HVT U367 ( .A1(n1820), .A2(sram_rdata_5[2]), .A3(n588), .A4(
        sram_rdata_4[2]), .A5(sram_rdata_3[2]), .A6(n1910), .Y(n1263) );
  AO222X1_HVT U368 ( .A1(n1820), .A2(sram_rdata_2[2]), .A3(n589), .A4(
        sram_rdata_1[2]), .A5(sram_rdata_0[2]), .A6(n1690), .Y(n894) );
  AOI22X1_HVT U369 ( .A1(n1263), .A2(n10900), .A3(n13000), .A4(n894), .Y(n605)
         );
  OA22X1_HVT U370 ( .A1(n11800), .A2(n384), .A3(n10000), .A4(n2880), .Y(n604)
         );
  NAND2X0_HVT U371 ( .A1(n1750), .A2(sram_rdata_6[2]), .Y(n603) );
  NAND3X0_HVT U372 ( .A1(n605), .A2(n604), .A3(n603), .Y(n_src_aox[2]) );
  AO222X1_HVT U373 ( .A1(n1810), .A2(sram_rdata_5[3]), .A3(n16100), .A4(
        sram_rdata_4[3]), .A5(sram_rdata_3[3]), .A6(n16500), .Y(n1265) );
  AO222X1_HVT U374 ( .A1(n1880), .A2(sram_rdata_2[3]), .A3(n2140), .A4(
        sram_rdata_1[3]), .A5(sram_rdata_0[3]), .A6(n1680), .Y(n898) );
  AOI22X1_HVT U375 ( .A1(n1265), .A2(n15100), .A3(n582), .A4(n898), .Y(n608)
         );
  OA22X1_HVT U376 ( .A1(n2770), .A2(n385), .A3(n10100), .A4(n2890), .Y(n607)
         );
  NAND2X0_HVT U377 ( .A1(n1770), .A2(sram_rdata_6[3]), .Y(n606) );
  NAND3X0_HVT U378 ( .A1(n608), .A2(n607), .A3(n606), .Y(n_src_aox[3]) );
  AO222X1_HVT U379 ( .A1(n2100), .A2(sram_rdata_5[4]), .A3(n588), .A4(
        sram_rdata_4[4]), .A5(sram_rdata_3[4]), .A6(n16500), .Y(n12701) );
  AO222X1_HVT U380 ( .A1(n2060), .A2(sram_rdata_2[4]), .A3(n15400), .A4(
        sram_rdata_1[4]), .A5(sram_rdata_0[4]), .A6(n2000), .Y(n902) );
  AOI22X1_HVT U381 ( .A1(n12701), .A2(n12800), .A3(n5801), .A4(n902), .Y(n611)
         );
  OA22X1_HVT U382 ( .A1(n13900), .A2(n386), .A3(n14600), .A4(n2900), .Y(n6101)
         );
  NAND2X0_HVT U383 ( .A1(n1760), .A2(sram_rdata_6[4]), .Y(n609) );
  NAND3X0_HVT U384 ( .A1(n611), .A2(n6101), .A3(n609), .Y(n_src_aox[4]) );
  AO222X1_HVT U385 ( .A1(n2060), .A2(sram_rdata_5[5]), .A3(n2180), .A4(
        sram_rdata_4[5]), .A5(sram_rdata_3[5]), .A6(n1950), .Y(n1275) );
  AO222X1_HVT U386 ( .A1(n2040), .A2(sram_rdata_2[5]), .A3(n2160), .A4(
        sram_rdata_1[5]), .A5(sram_rdata_0[5]), .A6(n1900), .Y(n906) );
  AOI22X1_HVT U387 ( .A1(n1275), .A2(n15000), .A3(n5801), .A4(n906), .Y(n614)
         );
  OA22X1_HVT U388 ( .A1(n2790), .A2(n387), .A3(n2720), .A4(n2910), .Y(n613) );
  NAND2X0_HVT U389 ( .A1(n1730), .A2(sram_rdata_6[5]), .Y(n612) );
  NAND3X0_HVT U390 ( .A1(n614), .A2(n613), .A3(n612), .Y(n_src_aox[5]) );
  AO222X1_HVT U391 ( .A1(n1870), .A2(sram_rdata_5[6]), .A3(n2160), .A4(
        sram_rdata_4[6]), .A5(sram_rdata_3[6]), .A6(n1990), .Y(n12801) );
  AO222X1_HVT U392 ( .A1(n2030), .A2(sram_rdata_2[6]), .A3(n16000), .A4(
        sram_rdata_1[6]), .A5(sram_rdata_0[6]), .A6(n2020), .Y(n9101) );
  AOI22X1_HVT U393 ( .A1(n12801), .A2(n15000), .A3(n10700), .A4(n9101), .Y(
        n617) );
  OA22X1_HVT U394 ( .A1(n13700), .A2(n388), .A3(n2740), .A4(n2920), .Y(n616)
         );
  NAND2X0_HVT U395 ( .A1(n1740), .A2(sram_rdata_6[6]), .Y(n615) );
  NAND3X0_HVT U396 ( .A1(n617), .A2(n616), .A3(n615), .Y(n_src_aox[6]) );
  AO222X1_HVT U397 ( .A1(n1890), .A2(sram_rdata_5[7]), .A3(n15500), .A4(
        sram_rdata_4[7]), .A5(sram_rdata_3[7]), .A6(n1980), .Y(n1285) );
  AO222X1_HVT U398 ( .A1(n1820), .A2(sram_rdata_2[7]), .A3(n2150), .A4(
        sram_rdata_1[7]), .A5(sram_rdata_0[7]), .A6(n1680), .Y(n914) );
  AOI22X1_HVT U399 ( .A1(n1285), .A2(n15100), .A3(n10700), .A4(n914), .Y(n6201) );
  OA22X1_HVT U400 ( .A1(n13700), .A2(n389), .A3(n10100), .A4(n2930), .Y(n619)
         );
  NAND2X0_HVT U401 ( .A1(n1700), .A2(sram_rdata_6[7]), .Y(n618) );
  NAND3X0_HVT U402 ( .A1(n6201), .A2(n619), .A3(n618), .Y(n_src_aox[7]) );
  AO222X1_HVT U403 ( .A1(n1840), .A2(sram_rdata_5[8]), .A3(n15900), .A4(
        sram_rdata_4[8]), .A5(sram_rdata_3[8]), .A6(n1680), .Y(n12901) );
  AO222X1_HVT U404 ( .A1(n14000), .A2(sram_rdata_2[8]), .A3(n2110), .A4(
        sram_rdata_1[8]), .A5(sram_rdata_0[8]), .A6(n16300), .Y(n918) );
  AOI22X1_HVT U405 ( .A1(n12901), .A2(n593), .A3(n583), .A4(n918), .Y(n623) );
  OA22X1_HVT U406 ( .A1(n10300), .A2(n3901), .A3(n14700), .A4(n2940), .Y(n622)
         );
  NAND2X0_HVT U407 ( .A1(n2270), .A2(sram_rdata_6[8]), .Y(n621) );
  NAND3X0_HVT U408 ( .A1(n623), .A2(n622), .A3(n621), .Y(n_src_aox[8]) );
  AO222X1_HVT U409 ( .A1(n2050), .A2(sram_rdata_5[9]), .A3(n16200), .A4(
        sram_rdata_4[9]), .A5(sram_rdata_3[9]), .A6(n1970), .Y(n1295) );
  AO222X1_HVT U410 ( .A1(n1820), .A2(sram_rdata_2[9]), .A3(n16100), .A4(
        sram_rdata_1[9]), .A5(sram_rdata_0[9]), .A6(n1930), .Y(n922) );
  AOI22X1_HVT U411 ( .A1(n1295), .A2(n12700), .A3(n11100), .A4(n922), .Y(n626)
         );
  OA22X1_HVT U412 ( .A1(n13800), .A2(n391), .A3(n2750), .A4(n2950), .Y(n625)
         );
  NAND2X0_HVT U413 ( .A1(n2220), .A2(sram_rdata_6[9]), .Y(n624) );
  NAND3X0_HVT U414 ( .A1(n626), .A2(n625), .A3(n624), .Y(n_src_aox[9]) );
  AO222X1_HVT U415 ( .A1(n2090), .A2(sram_rdata_5[10]), .A3(n16200), .A4(
        sram_rdata_4[10]), .A5(sram_rdata_3[10]), .A6(n1990), .Y(n13001) );
  AO222X1_HVT U416 ( .A1(n1870), .A2(sram_rdata_2[10]), .A3(n16200), .A4(
        sram_rdata_1[10]), .A5(sram_rdata_0[10]), .A6(n2010), .Y(n926) );
  AOI22X1_HVT U417 ( .A1(n13001), .A2(n10800), .A3(n12500), .A4(n926), .Y(n629) );
  OA22X1_HVT U418 ( .A1(n2780), .A2(n392), .A3(n1662), .A4(n2960), .Y(n628) );
  NAND2X0_HVT U419 ( .A1(n1710), .A2(sram_rdata_6[10]), .Y(n627) );
  NAND3X0_HVT U420 ( .A1(n629), .A2(n628), .A3(n627), .Y(n_src_aox[10]) );
  AO222X1_HVT U421 ( .A1(n14000), .A2(sram_rdata_5[11]), .A3(n2190), .A4(
        sram_rdata_4[11]), .A5(sram_rdata_3[11]), .A6(n1960), .Y(n1305) );
  AO222X1_HVT U422 ( .A1(n1810), .A2(sram_rdata_2[11]), .A3(n16100), .A4(
        sram_rdata_1[11]), .A5(sram_rdata_0[11]), .A6(n1910), .Y(n9301) );
  AOI22X1_HVT U423 ( .A1(n1305), .A2(n593), .A3(n12900), .A4(n9301), .Y(n632)
         );
  OA22X1_HVT U424 ( .A1(n11800), .A2(n393), .A3(n2700), .A4(n2970), .Y(n631)
         );
  NAND2X0_HVT U425 ( .A1(n2260), .A2(sram_rdata_6[11]), .Y(n6301) );
  NAND3X0_HVT U426 ( .A1(n632), .A2(n631), .A3(n6301), .Y(n_src_aox[11]) );
  AO222X1_HVT U427 ( .A1(n1810), .A2(sram_rdata_5[12]), .A3(n15900), .A4(
        sram_rdata_4[12]), .A5(sram_rdata_3[12]), .A6(n1930), .Y(n13101) );
  AO222X1_HVT U428 ( .A1(n2060), .A2(sram_rdata_2[12]), .A3(n15500), .A4(
        sram_rdata_1[12]), .A5(sram_rdata_0[12]), .A6(n1680), .Y(n934) );
  AOI22X1_HVT U429 ( .A1(n13101), .A2(n10900), .A3(n583), .A4(n934), .Y(n635)
         );
  OA22X1_HVT U430 ( .A1(n11600), .A2(n394), .A3(n10100), .A4(n2980), .Y(n634)
         );
  NAND2X0_HVT U431 ( .A1(n1700), .A2(sram_rdata_6[12]), .Y(n633) );
  NAND3X0_HVT U432 ( .A1(n635), .A2(n634), .A3(n633), .Y(n_src_aox[12]) );
  AO222X1_HVT U433 ( .A1(n1880), .A2(sram_rdata_5[13]), .A3(n16200), .A4(
        sram_rdata_4[13]), .A5(sram_rdata_3[13]), .A6(n16300), .Y(n1315) );
  AO222X1_HVT U434 ( .A1(n1890), .A2(sram_rdata_2[13]), .A3(n2140), .A4(
        sram_rdata_1[13]), .A5(sram_rdata_0[13]), .A6(n16400), .Y(n938) );
  AOI22X1_HVT U435 ( .A1(n1315), .A2(n593), .A3(n10700), .A4(n938), .Y(n638)
         );
  OA22X1_HVT U436 ( .A1(n10400), .A2(n395), .A3(n10000), .A4(n2990), .Y(n637)
         );
  NAND2X0_HVT U437 ( .A1(n1730), .A2(sram_rdata_6[13]), .Y(n636) );
  NAND3X0_HVT U438 ( .A1(n638), .A2(n637), .A3(n636), .Y(n_src_aox[13]) );
  AO222X1_HVT U439 ( .A1(n1810), .A2(sram_rdata_5[14]), .A3(n15700), .A4(
        sram_rdata_4[14]), .A5(sram_rdata_3[14]), .A6(n2020), .Y(n13201) );
  AO222X1_HVT U440 ( .A1(n1890), .A2(sram_rdata_2[14]), .A3(n16000), .A4(
        sram_rdata_1[14]), .A5(sram_rdata_0[14]), .A6(n16300), .Y(n942) );
  AOI22X1_HVT U441 ( .A1(n13201), .A2(n15000), .A3(n581), .A4(n942), .Y(n641)
         );
  OA22X1_HVT U442 ( .A1(n13800), .A2(n396), .A3(n2740), .A4(n3000), .Y(n6401)
         );
  NAND2X0_HVT U443 ( .A1(n1710), .A2(sram_rdata_6[14]), .Y(n639) );
  NAND3X0_HVT U444 ( .A1(n641), .A2(n6401), .A3(n639), .Y(n_src_aox[14]) );
  AO222X1_HVT U445 ( .A1(n1661), .A2(sram_rdata_5[15]), .A3(n2200), .A4(
        sram_rdata_4[15]), .A5(sram_rdata_3[15]), .A6(n16600), .Y(n1325) );
  AO222X1_HVT U446 ( .A1(n1880), .A2(sram_rdata_2[15]), .A3(n2200), .A4(
        sram_rdata_1[15]), .A5(sram_rdata_0[15]), .A6(n2010), .Y(n946) );
  AOI22X1_HVT U447 ( .A1(n1325), .A2(n593), .A3(n11000), .A4(n946), .Y(n644)
         );
  OA22X1_HVT U448 ( .A1(n1663), .A2(n397), .A3(n14600), .A4(n3010), .Y(n643)
         );
  NAND2X0_HVT U449 ( .A1(n2260), .A2(sram_rdata_6[15]), .Y(n642) );
  NAND3X0_HVT U450 ( .A1(n644), .A2(n643), .A3(n642), .Y(n_src_aox[15]) );
  AO222X1_HVT U451 ( .A1(n2070), .A2(sram_rdata_4[0]), .A3(n1950), .A4(
        sram_rdata_5[0]), .A5(n588), .A6(sram_rdata_3[0]), .Y(n1329) );
  AO222X1_HVT U452 ( .A1(n2100), .A2(sram_rdata_1[0]), .A3(n16000), .A4(
        sram_rdata_0[0]), .A5(sram_rdata_2[0]), .A6(n1950), .Y(n9501) );
  AOI22X1_HVT U453 ( .A1(n1329), .A2(n12800), .A3(n12500), .A4(n9501), .Y(n647) );
  OA22X1_HVT U454 ( .A1(n11600), .A2(n477), .A3(n2860), .A4(n11400), .Y(n646)
         );
  NAND2X0_HVT U455 ( .A1(n1790), .A2(sram_rdata_8[0]), .Y(n645) );
  NAND3X0_HVT U456 ( .A1(n647), .A2(n646), .A3(n645), .Y(n_src_aox[16]) );
  AO222X1_HVT U457 ( .A1(n2070), .A2(sram_rdata_4[1]), .A3(n2110), .A4(
        sram_rdata_3[1]), .A5(sram_rdata_5[1]), .A6(n2000), .Y(n1335) );
  AO222X1_HVT U458 ( .A1(n2100), .A2(sram_rdata_1[1]), .A3(n2170), .A4(
        sram_rdata_0[1]), .A5(sram_rdata_2[1]), .A6(n1960), .Y(n954) );
  AOI22X1_HVT U459 ( .A1(n1335), .A2(n593), .A3(n14400), .A4(n954), .Y(n6501)
         );
  OA22X1_HVT U460 ( .A1(n11700), .A2(n479), .A3(n2690), .A4(n383), .Y(n649) );
  NAND2X0_HVT U461 ( .A1(n2220), .A2(sram_rdata_8[1]), .Y(n648) );
  NAND3X0_HVT U462 ( .A1(n6501), .A2(n649), .A3(n648), .Y(n_src_aox[17]) );
  AO222X1_HVT U463 ( .A1(n1810), .A2(sram_rdata_4[2]), .A3(n2170), .A4(
        sram_rdata_3[2]), .A5(sram_rdata_5[2]), .A6(n1920), .Y(n13401) );
  AO222X1_HVT U464 ( .A1(n2050), .A2(sram_rdata_1[2]), .A3(n2180), .A4(
        sram_rdata_0[2]), .A5(sram_rdata_2[2]), .A6(n16300), .Y(n958) );
  AOI22X1_HVT U465 ( .A1(n13401), .A2(n591), .A3(n5801), .A4(n958), .Y(n653)
         );
  OA22X1_HVT U466 ( .A1(n2800), .A2(n4801), .A3(n2720), .A4(n384), .Y(n652) );
  NAND2X0_HVT U467 ( .A1(n1730), .A2(sram_rdata_8[2]), .Y(n651) );
  NAND3X0_HVT U468 ( .A1(n653), .A2(n652), .A3(n651), .Y(n_src_aox[18]) );
  AO222X1_HVT U469 ( .A1(n1880), .A2(sram_rdata_4[3]), .A3(n589), .A4(
        sram_rdata_3[3]), .A5(sram_rdata_5[3]), .A6(n1930), .Y(n1345) );
  AO222X1_HVT U470 ( .A1(n1810), .A2(sram_rdata_1[3]), .A3(n16000), .A4(
        sram_rdata_0[3]), .A5(sram_rdata_2[3]), .A6(n1670), .Y(n962) );
  AOI22X1_HVT U471 ( .A1(n1345), .A2(n10900), .A3(n11100), .A4(n962), .Y(n656)
         );
  OA22X1_HVT U472 ( .A1(n2780), .A2(n481), .A3(n14900), .A4(n385), .Y(n655) );
  NAND2X0_HVT U473 ( .A1(n1800), .A2(sram_rdata_8[3]), .Y(n654) );
  NAND3X0_HVT U474 ( .A1(n656), .A2(n655), .A3(n654), .Y(n_src_aox[19]) );
  AO222X1_HVT U475 ( .A1(n1661), .A2(sram_rdata_4[4]), .A3(n2130), .A4(
        sram_rdata_3[4]), .A5(sram_rdata_5[4]), .A6(n1990), .Y(n13501) );
  AO222X1_HVT U476 ( .A1(n1661), .A2(sram_rdata_1[4]), .A3(n15900), .A4(
        sram_rdata_0[4]), .A5(sram_rdata_2[4]), .A6(n16600), .Y(n966) );
  AOI22X1_HVT U477 ( .A1(n13501), .A2(n593), .A3(n582), .A4(n966), .Y(n659) );
  OA22X1_HVT U478 ( .A1(n10200), .A2(n482), .A3(n2700), .A4(n386), .Y(n658) );
  NAND2X0_HVT U479 ( .A1(n2270), .A2(sram_rdata_8[4]), .Y(n657) );
  NAND3X0_HVT U480 ( .A1(n659), .A2(n658), .A3(n657), .Y(n_src_aox[20]) );
  AO222X1_HVT U481 ( .A1(n1880), .A2(sram_rdata_4[5]), .A3(n15700), .A4(
        sram_rdata_3[5]), .A5(sram_rdata_5[5]), .A6(n1930), .Y(n1355) );
  AO222X1_HVT U482 ( .A1(n1860), .A2(sram_rdata_1[5]), .A3(n15600), .A4(
        sram_rdata_0[5]), .A5(sram_rdata_2[5]), .A6(n16400), .Y(n9701) );
  AOI22X1_HVT U483 ( .A1(n1355), .A2(n15000), .A3(n581), .A4(n9701), .Y(n662)
         );
  OA22X1_HVT U484 ( .A1(n2790), .A2(n483), .A3(n14700), .A4(n387), .Y(n661) );
  NAND2X0_HVT U485 ( .A1(n1800), .A2(sram_rdata_8[5]), .Y(n6601) );
  NAND3X0_HVT U486 ( .A1(n662), .A2(n661), .A3(n6601), .Y(n_src_aox[21]) );
  AO222X1_HVT U487 ( .A1(n2080), .A2(sram_rdata_4[6]), .A3(n2150), .A4(
        sram_rdata_3[6]), .A5(sram_rdata_5[6]), .A6(n16600), .Y(n1357) );
  AO222X1_HVT U488 ( .A1(n2060), .A2(sram_rdata_1[6]), .A3(n2110), .A4(
        sram_rdata_0[6]), .A5(sram_rdata_2[6]), .A6(n1690), .Y(n974) );
  AOI22X1_HVT U489 ( .A1(n1357), .A2(n10800), .A3(n11000), .A4(n974), .Y(n665)
         );
  OA22X1_HVT U490 ( .A1(n2790), .A2(n484), .A3(n2740), .A4(n388), .Y(n664) );
  NAND2X0_HVT U491 ( .A1(n2250), .A2(sram_rdata_8[6]), .Y(n663) );
  NAND3X0_HVT U492 ( .A1(n665), .A2(n664), .A3(n663), .Y(n_src_aox[22]) );
  AO222X1_HVT U493 ( .A1(n2060), .A2(sram_rdata_4[7]), .A3(n2160), .A4(
        sram_rdata_3[7]), .A5(sram_rdata_5[7]), .A6(n2000), .Y(n1362) );
  AO222X1_HVT U494 ( .A1(n2030), .A2(sram_rdata_1[7]), .A3(n2170), .A4(
        sram_rdata_0[7]), .A5(sram_rdata_2[7]), .A6(n1950), .Y(n978) );
  AOI22X1_HVT U495 ( .A1(n1362), .A2(n593), .A3(n11000), .A4(n978), .Y(n668)
         );
  OA22X1_HVT U496 ( .A1(n2760), .A2(n485), .A3(n2730), .A4(n389), .Y(n667) );
  NAND2X0_HVT U497 ( .A1(n575), .A2(sram_rdata_8[7]), .Y(n666) );
  NAND3X0_HVT U498 ( .A1(n668), .A2(n667), .A3(n666), .Y(n_src_aox[23]) );
  AO222X1_HVT U499 ( .A1(n1870), .A2(sram_rdata_4[8]), .A3(n2130), .A4(
        sram_rdata_3[8]), .A5(sram_rdata_5[8]), .A6(n1920), .Y(n1367) );
  AO222X1_HVT U500 ( .A1(n2050), .A2(sram_rdata_1[8]), .A3(n2160), .A4(
        sram_rdata_0[8]), .A5(sram_rdata_2[8]), .A6(n1990), .Y(n982) );
  AOI22X1_HVT U501 ( .A1(n1367), .A2(n15000), .A3(n582), .A4(n982), .Y(n671)
         );
  OA22X1_HVT U502 ( .A1(n2760), .A2(n486), .A3(n11400), .A4(n3901), .Y(n6701)
         );
  NAND2X0_HVT U503 ( .A1(n574), .A2(sram_rdata_8[8]), .Y(n669) );
  NAND3X0_HVT U504 ( .A1(n671), .A2(n6701), .A3(n669), .Y(n_src_aox[24]) );
  AO222X1_HVT U505 ( .A1(n1860), .A2(sram_rdata_4[9]), .A3(n589), .A4(
        sram_rdata_3[9]), .A5(sram_rdata_5[9]), .A6(n2020), .Y(n1372) );
  AO222X1_HVT U506 ( .A1(n1860), .A2(sram_rdata_1[9]), .A3(n15700), .A4(
        sram_rdata_0[9]), .A5(sram_rdata_2[9]), .A6(n1980), .Y(n986) );
  AOI22X1_HVT U507 ( .A1(n1372), .A2(n12700), .A3(n12400), .A4(n986), .Y(n674)
         );
  OA22X1_HVT U508 ( .A1(n2810), .A2(n487), .A3(n2710), .A4(n391), .Y(n673) );
  NAND2X0_HVT U509 ( .A1(n577), .A2(sram_rdata_8[9]), .Y(n672) );
  NAND3X0_HVT U510 ( .A1(n674), .A2(n673), .A3(n672), .Y(n_src_aox[25]) );
  AO222X1_HVT U511 ( .A1(n1810), .A2(sram_rdata_4[10]), .A3(n2150), .A4(
        sram_rdata_3[10]), .A5(sram_rdata_5[10]), .A6(n2020), .Y(n1377) );
  AO222X1_HVT U512 ( .A1(n1830), .A2(sram_rdata_1[10]), .A3(n15600), .A4(
        sram_rdata_0[10]), .A5(sram_rdata_2[10]), .A6(n16400), .Y(n9901) );
  AOI22X1_HVT U513 ( .A1(n1377), .A2(n15000), .A3(n13000), .A4(n9901), .Y(n677) );
  OA22X1_HVT U514 ( .A1(n10300), .A2(n488), .A3(n2730), .A4(n392), .Y(n676) );
  NAND2X0_HVT U515 ( .A1(n1760), .A2(sram_rdata_8[10]), .Y(n675) );
  NAND3X0_HVT U516 ( .A1(n677), .A2(n676), .A3(n675), .Y(n_src_aox[26]) );
  AO222X1_HVT U517 ( .A1(n12600), .A2(sram_rdata_4[11]), .A3(n15700), .A4(
        sram_rdata_3[11]), .A5(sram_rdata_5[11]), .A6(n1670), .Y(n1382) );
  AO222X1_HVT U518 ( .A1(n1810), .A2(sram_rdata_1[11]), .A3(n2190), .A4(
        sram_rdata_0[11]), .A5(sram_rdata_2[11]), .A6(n1960), .Y(n994) );
  AOI22X1_HVT U519 ( .A1(n1382), .A2(n593), .A3(n12900), .A4(n994), .Y(n6801)
         );
  OA22X1_HVT U520 ( .A1(n10200), .A2(n489), .A3(n10000), .A4(n393), .Y(n679)
         );
  NAND2X0_HVT U521 ( .A1(n2210), .A2(sram_rdata_8[11]), .Y(n678) );
  NAND3X0_HVT U522 ( .A1(n6801), .A2(n679), .A3(n678), .Y(n_src_aox[27]) );
  AO222X1_HVT U523 ( .A1(n2100), .A2(sram_rdata_4[12]), .A3(n15700), .A4(
        sram_rdata_3[12]), .A5(sram_rdata_5[12]), .A6(n1910), .Y(n1387) );
  AO222X1_HVT U524 ( .A1(n2030), .A2(sram_rdata_1[12]), .A3(n588), .A4(
        sram_rdata_0[12]), .A5(sram_rdata_2[12]), .A6(n1670), .Y(n998) );
  AOI22X1_HVT U525 ( .A1(n1387), .A2(n12800), .A3(n10700), .A4(n998), .Y(n683)
         );
  OA22X1_HVT U526 ( .A1(n2770), .A2(n4901), .A3(n14700), .A4(n394), .Y(n682)
         );
  NAND2X0_HVT U527 ( .A1(n578), .A2(sram_rdata_8[12]), .Y(n681) );
  NAND3X0_HVT U528 ( .A1(n683), .A2(n682), .A3(n681), .Y(n_src_aox[28]) );
  AO222X1_HVT U529 ( .A1(n1810), .A2(sram_rdata_4[13]), .A3(n15700), .A4(
        sram_rdata_3[13]), .A5(sram_rdata_5[13]), .A6(n1990), .Y(n1392) );
  AO222X1_HVT U530 ( .A1(n1880), .A2(sram_rdata_1[13]), .A3(n2200), .A4(
        sram_rdata_0[13]), .A5(sram_rdata_2[13]), .A6(n1960), .Y(n1002) );
  AOI22X1_HVT U531 ( .A1(n1392), .A2(n10900), .A3(n11100), .A4(n1002), .Y(n686) );
  OA22X1_HVT U532 ( .A1(n10400), .A2(n491), .A3(n2710), .A4(n395), .Y(n685) );
  NAND2X0_HVT U533 ( .A1(n577), .A2(sram_rdata_8[13]), .Y(n684) );
  NAND3X0_HVT U534 ( .A1(n686), .A2(n685), .A3(n684), .Y(n_src_aox[29]) );
  AO222X1_HVT U535 ( .A1(n1880), .A2(sram_rdata_4[14]), .A3(n15900), .A4(
        sram_rdata_3[14]), .A5(sram_rdata_5[14]), .A6(n1920), .Y(n1397) );
  AO222X1_HVT U536 ( .A1(n2040), .A2(sram_rdata_1[14]), .A3(n589), .A4(
        sram_rdata_0[14]), .A5(sram_rdata_2[14]), .A6(n1910), .Y(n1006) );
  AOI22X1_HVT U537 ( .A1(n1397), .A2(n591), .A3(n11000), .A4(n1006), .Y(n689)
         );
  OA22X1_HVT U538 ( .A1(n10400), .A2(n492), .A3(n2720), .A4(n396), .Y(n688) );
  NAND2X0_HVT U539 ( .A1(n2240), .A2(sram_rdata_8[14]), .Y(n687) );
  NAND3X0_HVT U540 ( .A1(n689), .A2(n688), .A3(n687), .Y(n_src_aox[30]) );
  AO222X1_HVT U541 ( .A1(n1830), .A2(sram_rdata_4[15]), .A3(n588), .A4(
        sram_rdata_3[15]), .A5(sram_rdata_5[15]), .A6(n2010), .Y(n1399) );
  AO222X1_HVT U542 ( .A1(n1810), .A2(sram_rdata_1[15]), .A3(n16000), .A4(
        sram_rdata_0[15]), .A5(sram_rdata_2[15]), .A6(n16600), .Y(n10101) );
  AOI22X1_HVT U543 ( .A1(n1399), .A2(n15000), .A3(n583), .A4(n10101), .Y(n692)
         );
  OA22X1_HVT U544 ( .A1(n13700), .A2(n493), .A3(n14800), .A4(n397), .Y(n691)
         );
  NAND2X0_HVT U545 ( .A1(n574), .A2(sram_rdata_8[15]), .Y(n6901) );
  NAND3X0_HVT U546 ( .A1(n692), .A2(n691), .A3(n6901), .Y(n_src_aox[31]) );
  AO222X1_HVT U547 ( .A1(n2040), .A2(sram_rdata_3[0]), .A3(n1900), .A4(
        sram_rdata_4[0]), .A5(n2170), .A6(sram_rdata_5[0]), .Y(n1403) );
  AO222X1_HVT U548 ( .A1(n2070), .A2(sram_rdata_0[0]), .A3(n2150), .A4(
        sram_rdata_2[0]), .A5(n1990), .A6(sram_rdata_1[0]), .Y(n1014) );
  AOI22X1_HVT U549 ( .A1(n1403), .A2(n1664), .A3(n582), .A4(n1014), .Y(n695)
         );
  OA22X1_HVT U550 ( .A1(n1663), .A2(n573), .A3(n477), .A4(n2750), .Y(n694) );
  NAND2X0_HVT U551 ( .A1(n575), .A2(sram_rdata_7[0]), .Y(n693) );
  NAND3X0_HVT U552 ( .A1(n695), .A2(n694), .A3(n693), .Y(n_src_aox[32]) );
  AO222X1_HVT U553 ( .A1(n2030), .A2(sram_rdata_3[1]), .A3(n16200), .A4(
        sram_rdata_5[1]), .A5(n1980), .A6(sram_rdata_4[1]), .Y(n1406) );
  AO222X1_HVT U554 ( .A1(n1840), .A2(sram_rdata_0[1]), .A3(n2140), .A4(
        sram_rdata_2[1]), .A5(n1920), .A6(sram_rdata_1[1]), .Y(n1018) );
  AOI22X1_HVT U555 ( .A1(n1406), .A2(n10900), .A3(n12400), .A4(n1018), .Y(n698) );
  OA22X1_HVT U556 ( .A1(n10300), .A2(n2870), .A3(n14600), .A4(n479), .Y(n697)
         );
  NAND2X0_HVT U557 ( .A1(n1710), .A2(sram_rdata_7[1]), .Y(n696) );
  NAND3X0_HVT U558 ( .A1(n698), .A2(n697), .A3(n696), .Y(n_src_aox[33]) );
  AO222X1_HVT U559 ( .A1(n2080), .A2(sram_rdata_3[2]), .A3(n16100), .A4(
        sram_rdata_5[2]), .A5(n1680), .A6(sram_rdata_4[2]), .Y(n1411) );
  AO222X1_HVT U560 ( .A1(n2090), .A2(sram_rdata_0[2]), .A3(n2190), .A4(
        sram_rdata_2[2]), .A5(n16300), .A6(sram_rdata_1[2]), .Y(n1022) );
  AOI22X1_HVT U561 ( .A1(n1411), .A2(n10800), .A3(n10700), .A4(n1022), .Y(n701) );
  OA22X1_HVT U562 ( .A1(n1663), .A2(n2880), .A3(n11400), .A4(n4801), .Y(n7001)
         );
  NAND2X0_HVT U563 ( .A1(n1780), .A2(sram_rdata_7[2]), .Y(n699) );
  NAND3X0_HVT U564 ( .A1(n701), .A2(n7001), .A3(n699), .Y(n_src_aox[34]) );
  AO222X1_HVT U565 ( .A1(n2070), .A2(sram_rdata_3[3]), .A3(n2140), .A4(
        sram_rdata_5[3]), .A5(n1950), .A6(sram_rdata_4[3]), .Y(n1416) );
  AO222X1_HVT U566 ( .A1(n2080), .A2(sram_rdata_0[3]), .A3(n589), .A4(
        sram_rdata_2[3]), .A5(n1920), .A6(sram_rdata_1[3]), .Y(n1026) );
  AOI22X1_HVT U567 ( .A1(n1416), .A2(n594), .A3(n11000), .A4(n1026), .Y(n704)
         );
  OA22X1_HVT U568 ( .A1(n2770), .A2(n2890), .A3(n2730), .A4(n481), .Y(n703) );
  NAND2X0_HVT U569 ( .A1(n1780), .A2(sram_rdata_7[3]), .Y(n702) );
  NAND3X0_HVT U570 ( .A1(n704), .A2(n703), .A3(n702), .Y(n_src_aox[35]) );
  AO222X1_HVT U571 ( .A1(n1860), .A2(sram_rdata_3[4]), .A3(n2170), .A4(
        sram_rdata_5[4]), .A5(n1670), .A6(sram_rdata_4[4]), .Y(n1418) );
  AO222X1_HVT U572 ( .A1(n2030), .A2(sram_rdata_0[4]), .A3(n2190), .A4(
        sram_rdata_2[4]), .A5(n2020), .A6(sram_rdata_1[4]), .Y(n10301) );
  AOI22X1_HVT U573 ( .A1(n1418), .A2(n593), .A3(n581), .A4(n10301), .Y(n707)
         );
  OA22X1_HVT U574 ( .A1(n2810), .A2(n2900), .A3(n14900), .A4(n482), .Y(n706)
         );
  NAND2X0_HVT U575 ( .A1(n1760), .A2(sram_rdata_7[4]), .Y(n705) );
  NAND3X0_HVT U576 ( .A1(n707), .A2(n706), .A3(n705), .Y(n_src_aox[36]) );
  AO222X1_HVT U577 ( .A1(n1830), .A2(sram_rdata_3[5]), .A3(n2200), .A4(
        sram_rdata_5[5]), .A5(n1980), .A6(sram_rdata_4[5]), .Y(n1423) );
  AO222X1_HVT U578 ( .A1(n1840), .A2(sram_rdata_0[5]), .A3(n588), .A4(
        sram_rdata_2[5]), .A5(n1910), .A6(sram_rdata_1[5]), .Y(n1034) );
  AOI22X1_HVT U579 ( .A1(n1423), .A2(n593), .A3(n12900), .A4(n1034), .Y(n7101)
         );
  OA22X1_HVT U580 ( .A1(n13800), .A2(n2910), .A3(n2700), .A4(n483), .Y(n709)
         );
  NAND2X0_HVT U581 ( .A1(n2270), .A2(sram_rdata_7[5]), .Y(n708) );
  NAND3X0_HVT U582 ( .A1(n7101), .A2(n709), .A3(n708), .Y(n_src_aox[37]) );
  AO222X1_HVT U583 ( .A1(n1860), .A2(sram_rdata_3[6]), .A3(n15700), .A4(
        sram_rdata_5[6]), .A5(n1930), .A6(sram_rdata_4[6]), .Y(n1428) );
  AO222X1_HVT U584 ( .A1(n2090), .A2(sram_rdata_0[6]), .A3(n2160), .A4(
        sram_rdata_2[6]), .A5(n1920), .A6(sram_rdata_1[6]), .Y(n1038) );
  AOI22X1_HVT U585 ( .A1(n1428), .A2(n591), .A3(n582), .A4(n1038), .Y(n713) );
  OA22X1_HVT U586 ( .A1(n10200), .A2(n2920), .A3(n2700), .A4(n484), .Y(n712)
         );
  NAND2X0_HVT U587 ( .A1(n1780), .A2(sram_rdata_7[6]), .Y(n711) );
  NAND3X0_HVT U588 ( .A1(n713), .A2(n712), .A3(n711), .Y(n_src_aox[38]) );
  AO222X1_HVT U589 ( .A1(n12600), .A2(sram_rdata_3[7]), .A3(n16000), .A4(
        sram_rdata_5[7]), .A5(n1670), .A6(sram_rdata_4[7]), .Y(n14301) );
  AO222X1_HVT U590 ( .A1(n1830), .A2(sram_rdata_0[7]), .A3(n2140), .A4(
        sram_rdata_2[7]), .A5(n1910), .A6(sram_rdata_1[7]), .Y(n1042) );
  AOI22X1_HVT U591 ( .A1(n14301), .A2(n15000), .A3(n5801), .A4(n1042), .Y(n716) );
  OA22X1_HVT U592 ( .A1(n13600), .A2(n2930), .A3(n2750), .A4(n485), .Y(n715)
         );
  NAND2X0_HVT U593 ( .A1(n1780), .A2(sram_rdata_7[7]), .Y(n714) );
  NAND3X0_HVT U594 ( .A1(n716), .A2(n715), .A3(n714), .Y(n_src_aox[39]) );
  AO222X1_HVT U595 ( .A1(n2090), .A2(sram_rdata_3[8]), .A3(n15400), .A4(
        sram_rdata_5[8]), .A5(n16600), .A6(sram_rdata_4[8]), .Y(n1435) );
  AO222X1_HVT U596 ( .A1(n2050), .A2(sram_rdata_0[8]), .A3(n2140), .A4(
        sram_rdata_2[8]), .A5(n1980), .A6(sram_rdata_1[8]), .Y(n1046) );
  AOI22X1_HVT U597 ( .A1(n1435), .A2(n12800), .A3(n11000), .A4(n1046), .Y(n719) );
  OA22X1_HVT U598 ( .A1(n13800), .A2(n2940), .A3(n14800), .A4(n486), .Y(n718)
         );
  NAND2X0_HVT U599 ( .A1(n1730), .A2(sram_rdata_7[8]), .Y(n717) );
  NAND3X0_HVT U600 ( .A1(n719), .A2(n718), .A3(n717), .Y(n_src_aox[40]) );
  AO222X1_HVT U601 ( .A1(n2050), .A2(sram_rdata_3[9]), .A3(n15600), .A4(
        sram_rdata_5[9]), .A5(n16500), .A6(sram_rdata_4[9]), .Y(n14401) );
  AO222X1_HVT U602 ( .A1(n2030), .A2(sram_rdata_0[9]), .A3(n15600), .A4(
        sram_rdata_2[9]), .A5(n2000), .A6(sram_rdata_1[9]), .Y(n10501) );
  AOI22X1_HVT U603 ( .A1(n14401), .A2(n591), .A3(n12500), .A4(n10501), .Y(n722) );
  OA22X1_HVT U604 ( .A1(n2800), .A2(n2950), .A3(n14700), .A4(n487), .Y(n721)
         );
  NAND2X0_HVT U605 ( .A1(n1780), .A2(sram_rdata_7[9]), .Y(n7201) );
  NAND3X0_HVT U606 ( .A1(n722), .A2(n721), .A3(n7201), .Y(n_src_aox[41]) );
  AO222X1_HVT U607 ( .A1(n1820), .A2(sram_rdata_3[10]), .A3(n2180), .A4(
        sram_rdata_5[10]), .A5(n1970), .A6(sram_rdata_4[10]), .Y(n1445) );
  AO222X1_HVT U608 ( .A1(n2060), .A2(sram_rdata_0[10]), .A3(n2150), .A4(
        sram_rdata_2[10]), .A5(n1990), .A6(sram_rdata_1[10]), .Y(n1054) );
  AOI22X1_HVT U609 ( .A1(n1445), .A2(n15100), .A3(n583), .A4(n1054), .Y(n725)
         );
  OA22X1_HVT U610 ( .A1(n13700), .A2(n2960), .A3(n14600), .A4(n488), .Y(n724)
         );
  NAND2X0_HVT U611 ( .A1(n2240), .A2(sram_rdata_7[10]), .Y(n723) );
  NAND3X0_HVT U612 ( .A1(n725), .A2(n724), .A3(n723), .Y(n_src_aox[42]) );
  AO222X1_HVT U613 ( .A1(n1840), .A2(sram_rdata_3[11]), .A3(n2160), .A4(
        sram_rdata_5[11]), .A5(n1970), .A6(sram_rdata_4[11]), .Y(n14501) );
  AO222X1_HVT U614 ( .A1(n2030), .A2(sram_rdata_0[11]), .A3(n15700), .A4(
        sram_rdata_2[11]), .A5(n1910), .A6(sram_rdata_1[11]), .Y(n1058) );
  AOI22X1_HVT U615 ( .A1(n14501), .A2(n1664), .A3(n5801), .A4(n1058), .Y(n728)
         );
  OA22X1_HVT U616 ( .A1(n11800), .A2(n2970), .A3(n2720), .A4(n489), .Y(n727)
         );
  NAND2X0_HVT U617 ( .A1(n1750), .A2(sram_rdata_7[11]), .Y(n726) );
  NAND3X0_HVT U618 ( .A1(n728), .A2(n727), .A3(n726), .Y(n_src_aox[43]) );
  AO222X1_HVT U619 ( .A1(n12600), .A2(sram_rdata_3[12]), .A3(n16000), .A4(
        sram_rdata_5[12]), .A5(n16400), .A6(sram_rdata_4[12]), .Y(n1455) );
  AO222X1_HVT U620 ( .A1(n1870), .A2(sram_rdata_0[12]), .A3(n2150), .A4(
        sram_rdata_2[12]), .A5(n1900), .A6(sram_rdata_1[12]), .Y(n1062) );
  AOI22X1_HVT U621 ( .A1(n1455), .A2(n12700), .A3(n5801), .A4(n1062), .Y(n731)
         );
  OA22X1_HVT U622 ( .A1(n11700), .A2(n2980), .A3(n2750), .A4(n4901), .Y(n7301)
         );
  NAND2X0_HVT U623 ( .A1(n2250), .A2(sram_rdata_7[12]), .Y(n729) );
  NAND3X0_HVT U624 ( .A1(n731), .A2(n7301), .A3(n729), .Y(n_src_aox[44]) );
  AO222X1_HVT U625 ( .A1(n1880), .A2(sram_rdata_3[13]), .A3(n15500), .A4(
        sram_rdata_5[13]), .A5(n16600), .A6(sram_rdata_4[13]), .Y(n14601) );
  AO222X1_HVT U626 ( .A1(n1870), .A2(sram_rdata_0[13]), .A3(n588), .A4(
        sram_rdata_2[13]), .A5(n1910), .A6(sram_rdata_1[13]), .Y(n1066) );
  AOI22X1_HVT U627 ( .A1(n14601), .A2(n593), .A3(n11100), .A4(n1066), .Y(n734)
         );
  OA22X1_HVT U628 ( .A1(n11600), .A2(n2990), .A3(n2690), .A4(n491), .Y(n733)
         );
  NAND2X0_HVT U629 ( .A1(n2210), .A2(sram_rdata_7[13]), .Y(n732) );
  NAND3X0_HVT U630 ( .A1(n734), .A2(n733), .A3(n732), .Y(n_src_aox[45]) );
  AO222X1_HVT U631 ( .A1(n2070), .A2(sram_rdata_3[14]), .A3(n15600), .A4(
        sram_rdata_5[14]), .A5(n2000), .A6(sram_rdata_4[14]), .Y(n1465) );
  AO222X1_HVT U632 ( .A1(n1820), .A2(sram_rdata_0[14]), .A3(n16100), .A4(
        sram_rdata_2[14]), .A5(n1960), .A6(sram_rdata_1[14]), .Y(n10701) );
  AOI22X1_HVT U633 ( .A1(n1465), .A2(n10800), .A3(n11000), .A4(n10701), .Y(
        n737) );
  OA22X1_HVT U634 ( .A1(n2780), .A2(n3000), .A3(n2690), .A4(n492), .Y(n736) );
  NAND2X0_HVT U635 ( .A1(n578), .A2(sram_rdata_7[14]), .Y(n735) );
  NAND3X0_HVT U636 ( .A1(n737), .A2(n736), .A3(n735), .Y(n_src_aox[46]) );
  AO222X1_HVT U637 ( .A1(n1661), .A2(sram_rdata_3[15]), .A3(n15900), .A4(
        sram_rdata_5[15]), .A5(n1680), .A6(sram_rdata_4[15]), .Y(n1467) );
  AO222X1_HVT U638 ( .A1(n1661), .A2(sram_rdata_0[15]), .A3(n16100), .A4(
        sram_rdata_2[15]), .A5(n2020), .A6(sram_rdata_1[15]), .Y(n1074) );
  AOI22X1_HVT U639 ( .A1(n1467), .A2(n591), .A3(n11100), .A4(n1074), .Y(n7401)
         );
  OA22X1_HVT U640 ( .A1(n13700), .A2(n3010), .A3(n14900), .A4(n493), .Y(n739)
         );
  NAND2X0_HVT U641 ( .A1(n2240), .A2(sram_rdata_7[15]), .Y(n738) );
  NAND3X0_HVT U642 ( .A1(n7401), .A2(n739), .A3(n738), .Y(n_src_aox[47]) );
  AO222X1_HVT U643 ( .A1(n1880), .A2(sram_rdata_5[16]), .A3(n2200), .A4(
        sram_rdata_4[16]), .A5(sram_rdata_3[16]), .A6(n2020), .Y(n1472) );
  AO222X1_HVT U644 ( .A1(n2050), .A2(sram_rdata_2[16]), .A3(n2200), .A4(
        sram_rdata_1[16]), .A5(sram_rdata_0[16]), .A6(n16400), .Y(n1078) );
  AOI22X1_HVT U645 ( .A1(n1472), .A2(n12700), .A3(n582), .A4(n1078), .Y(n743)
         );
  OA22X1_HVT U646 ( .A1(n10400), .A2(n398), .A3(n1662), .A4(n3020), .Y(n742)
         );
  NAND2X0_HVT U647 ( .A1(n577), .A2(sram_rdata_6[16]), .Y(n741) );
  NAND3X0_HVT U648 ( .A1(n743), .A2(n742), .A3(n741), .Y(n_src_aox[48]) );
  AO222X1_HVT U649 ( .A1(n12600), .A2(sram_rdata_5[17]), .A3(n16200), .A4(
        sram_rdata_4[17]), .A5(sram_rdata_3[17]), .A6(n16400), .Y(n1477) );
  AO222X1_HVT U650 ( .A1(n1840), .A2(sram_rdata_2[17]), .A3(n15900), .A4(
        sram_rdata_1[17]), .A5(sram_rdata_0[17]), .A6(n1670), .Y(n1082) );
  AOI22X1_HVT U651 ( .A1(n1477), .A2(n15100), .A3(n14400), .A4(n1082), .Y(n746) );
  OA22X1_HVT U652 ( .A1(n10300), .A2(n399), .A3(n11400), .A4(n3030), .Y(n745)
         );
  NAND2X0_HVT U653 ( .A1(n1770), .A2(sram_rdata_6[17]), .Y(n744) );
  NAND3X0_HVT U654 ( .A1(n746), .A2(n745), .A3(n744), .Y(n_src_aox[49]) );
  AO222X1_HVT U655 ( .A1(n1890), .A2(sram_rdata_5[18]), .A3(n589), .A4(
        sram_rdata_4[18]), .A5(sram_rdata_3[18]), .A6(n2010), .Y(n1482) );
  AO222X1_HVT U656 ( .A1(n1830), .A2(sram_rdata_2[18]), .A3(n2140), .A4(
        sram_rdata_1[18]), .A5(sram_rdata_0[18]), .A6(n1980), .Y(n1086) );
  AOI22X1_HVT U657 ( .A1(n1482), .A2(n10900), .A3(n12500), .A4(n1086), .Y(n749) );
  OA22X1_HVT U658 ( .A1(n13600), .A2(n4001), .A3(n2700), .A4(n3040), .Y(n748)
         );
  NAND2X0_HVT U659 ( .A1(n1710), .A2(sram_rdata_6[18]), .Y(n747) );
  NAND3X0_HVT U660 ( .A1(n749), .A2(n748), .A3(n747), .Y(n_src_aox[50]) );
  AO222X1_HVT U661 ( .A1(n1870), .A2(sram_rdata_5[19]), .A3(n15500), .A4(
        sram_rdata_4[19]), .A5(sram_rdata_3[19]), .A6(n2010), .Y(n1487) );
  AO222X1_HVT U662 ( .A1(n12600), .A2(sram_rdata_2[19]), .A3(n16200), .A4(
        sram_rdata_1[19]), .A5(sram_rdata_0[19]), .A6(n1970), .Y(n10901) );
  AOI22X1_HVT U663 ( .A1(n1487), .A2(n15100), .A3(n5801), .A4(n10901), .Y(n752) );
  OA22X1_HVT U664 ( .A1(n2780), .A2(n401), .A3(n1662), .A4(n3050), .Y(n751) );
  NAND2X0_HVT U665 ( .A1(n2260), .A2(sram_rdata_6[19]), .Y(n7501) );
  NAND3X0_HVT U666 ( .A1(n752), .A2(n751), .A3(n7501), .Y(n_src_aox[51]) );
  AO222X1_HVT U667 ( .A1(n2080), .A2(sram_rdata_5[20]), .A3(n16100), .A4(
        sram_rdata_4[20]), .A5(sram_rdata_3[20]), .A6(n1920), .Y(n1492) );
  AO222X1_HVT U668 ( .A1(n2090), .A2(sram_rdata_2[20]), .A3(n2190), .A4(
        sram_rdata_1[20]), .A5(sram_rdata_0[20]), .A6(n16500), .Y(n1094) );
  AOI22X1_HVT U669 ( .A1(n1492), .A2(n10800), .A3(n12400), .A4(n1094), .Y(n755) );
  OA22X1_HVT U670 ( .A1(n2810), .A2(n402), .A3(n2730), .A4(n3060), .Y(n754) );
  NAND2X0_HVT U671 ( .A1(n2210), .A2(sram_rdata_6[20]), .Y(n753) );
  NAND3X0_HVT U672 ( .A1(n755), .A2(n754), .A3(n753), .Y(n_src_aox[52]) );
  AO222X1_HVT U673 ( .A1(n2100), .A2(sram_rdata_5[21]), .A3(n2110), .A4(
        sram_rdata_4[21]), .A5(sram_rdata_3[21]), .A6(n1910), .Y(n1494) );
  AO222X1_HVT U674 ( .A1(n2070), .A2(sram_rdata_2[21]), .A3(n589), .A4(
        sram_rdata_1[21]), .A5(sram_rdata_0[21]), .A6(n16600), .Y(n1098) );
  AOI22X1_HVT U675 ( .A1(n1494), .A2(n15100), .A3(n583), .A4(n1098), .Y(n758)
         );
  OA22X1_HVT U676 ( .A1(n2790), .A2(n403), .A3(n2710), .A4(n3070), .Y(n757) );
  NAND2X0_HVT U677 ( .A1(n576), .A2(sram_rdata_6[21]), .Y(n756) );
  NAND3X0_HVT U678 ( .A1(n758), .A2(n757), .A3(n756), .Y(n_src_aox[53]) );
  AO222X1_HVT U679 ( .A1(n1890), .A2(sram_rdata_5[22]), .A3(n2180), .A4(
        sram_rdata_4[22]), .A5(sram_rdata_3[22]), .A6(n1670), .Y(n1499) );
  AO222X1_HVT U680 ( .A1(n2040), .A2(sram_rdata_2[22]), .A3(n2170), .A4(
        sram_rdata_1[22]), .A5(sram_rdata_0[22]), .A6(n16300), .Y(n1102) );
  AOI22X1_HVT U681 ( .A1(n1499), .A2(n15000), .A3(n582), .A4(n1102), .Y(n761)
         );
  OA22X1_HVT U682 ( .A1(n10200), .A2(n404), .A3(n10100), .A4(n3080), .Y(n7601)
         );
  NAND2X0_HVT U683 ( .A1(n1760), .A2(sram_rdata_6[22]), .Y(n759) );
  NAND3X0_HVT U684 ( .A1(n761), .A2(n7601), .A3(n759), .Y(n_src_aox[54]) );
  AO222X1_HVT U685 ( .A1(n2060), .A2(sram_rdata_5[23]), .A3(n2200), .A4(
        sram_rdata_4[23]), .A5(sram_rdata_3[23]), .A6(n1680), .Y(n1504) );
  AO222X1_HVT U686 ( .A1(n2040), .A2(sram_rdata_2[23]), .A3(n16000), .A4(
        sram_rdata_1[23]), .A5(sram_rdata_0[23]), .A6(n1670), .Y(n1106) );
  AOI22X1_HVT U687 ( .A1(n1504), .A2(n593), .A3(n12900), .A4(n1106), .Y(n764)
         );
  OA22X1_HVT U688 ( .A1(n13700), .A2(n405), .A3(n14800), .A4(n3090), .Y(n763)
         );
  NAND2X0_HVT U689 ( .A1(n1770), .A2(sram_rdata_6[23]), .Y(n762) );
  NAND3X0_HVT U690 ( .A1(n764), .A2(n763), .A3(n762), .Y(n_src_aox[55]) );
  AO222X1_HVT U691 ( .A1(n1661), .A2(sram_rdata_5[24]), .A3(n15700), .A4(
        sram_rdata_4[24]), .A5(sram_rdata_3[24]), .A6(n16300), .Y(n1509) );
  AO222X1_HVT U692 ( .A1(n12600), .A2(sram_rdata_2[24]), .A3(n2130), .A4(
        sram_rdata_1[24]), .A5(sram_rdata_0[24]), .A6(n16500), .Y(n11101) );
  AOI22X1_HVT U693 ( .A1(n1509), .A2(n15100), .A3(n582), .A4(n11101), .Y(n767)
         );
  OA22X1_HVT U694 ( .A1(n13800), .A2(n406), .A3(n14900), .A4(n3100), .Y(n766)
         );
  NAND2X0_HVT U695 ( .A1(n2220), .A2(sram_rdata_6[24]), .Y(n765) );
  NAND3X0_HVT U696 ( .A1(n767), .A2(n766), .A3(n765), .Y(n_src_aox[56]) );
  AO222X1_HVT U697 ( .A1(n1830), .A2(sram_rdata_5[25]), .A3(n15500), .A4(
        sram_rdata_4[25]), .A5(sram_rdata_3[25]), .A6(n2000), .Y(n1514) );
  AO222X1_HVT U698 ( .A1(n1840), .A2(sram_rdata_2[25]), .A3(n2110), .A4(
        sram_rdata_1[25]), .A5(sram_rdata_0[25]), .A6(n1970), .Y(n1114) );
  AOI22X1_HVT U699 ( .A1(n1514), .A2(n591), .A3(n13000), .A4(n1114), .Y(n7701)
         );
  OA22X1_HVT U700 ( .A1(n13800), .A2(n407), .A3(n2750), .A4(n3110), .Y(n769)
         );
  NAND2X0_HVT U701 ( .A1(n1780), .A2(sram_rdata_6[25]), .Y(n768) );
  NAND3X0_HVT U702 ( .A1(n7701), .A2(n769), .A3(n768), .Y(n_src_aox[57]) );
  AO222X1_HVT U703 ( .A1(n2100), .A2(sram_rdata_5[26]), .A3(n15400), .A4(
        sram_rdata_4[26]), .A5(sram_rdata_3[26]), .A6(n1930), .Y(n1519) );
  AO222X1_HVT U704 ( .A1(n2040), .A2(sram_rdata_2[26]), .A3(n2130), .A4(
        sram_rdata_1[26]), .A5(sram_rdata_0[26]), .A6(n1990), .Y(n1118) );
  AOI22X1_HVT U705 ( .A1(n1519), .A2(n12800), .A3(n583), .A4(n1118), .Y(n773)
         );
  OA22X1_HVT U706 ( .A1(n2760), .A2(n408), .A3(n2710), .A4(n3120), .Y(n772) );
  NAND2X0_HVT U707 ( .A1(n2250), .A2(sram_rdata_6[26]), .Y(n771) );
  NAND3X0_HVT U708 ( .A1(n773), .A2(n772), .A3(n771), .Y(n_src_aox[58]) );
  AO222X1_HVT U709 ( .A1(n2050), .A2(sram_rdata_5[27]), .A3(n15500), .A4(
        sram_rdata_4[27]), .A5(sram_rdata_3[27]), .A6(n2020), .Y(n1524) );
  AO222X1_HVT U710 ( .A1(n2050), .A2(sram_rdata_2[27]), .A3(n15600), .A4(
        sram_rdata_1[27]), .A5(sram_rdata_0[27]), .A6(n1950), .Y(n1122) );
  AOI22X1_HVT U711 ( .A1(n1524), .A2(n15100), .A3(n10700), .A4(n1122), .Y(n777) );
  OA22X1_HVT U712 ( .A1(n11800), .A2(n409), .A3(n10000), .A4(n3130), .Y(n775)
         );
  NAND2X0_HVT U713 ( .A1(n1760), .A2(sram_rdata_6[27]), .Y(n774) );
  NAND3X0_HVT U714 ( .A1(n777), .A2(n775), .A3(n774), .Y(n_src_aox[59]) );
  AO222X1_HVT U715 ( .A1(n1870), .A2(sram_rdata_5[28]), .A3(n2190), .A4(
        sram_rdata_4[28]), .A5(sram_rdata_3[28]), .A6(n1920), .Y(n1526) );
  AO222X1_HVT U716 ( .A1(n2040), .A2(sram_rdata_2[28]), .A3(n2150), .A4(
        sram_rdata_1[28]), .A5(sram_rdata_0[28]), .A6(n1690), .Y(n1126) );
  AOI22X1_HVT U717 ( .A1(n1526), .A2(n15000), .A3(n582), .A4(n1126), .Y(n7801)
         );
  OA22X1_HVT U718 ( .A1(n11700), .A2(n4101), .A3(n2740), .A4(n3140), .Y(n779)
         );
  NAND2X0_HVT U719 ( .A1(n2220), .A2(sram_rdata_6[28]), .Y(n778) );
  NAND3X0_HVT U720 ( .A1(n7801), .A2(n779), .A3(n778), .Y(n_src_aox[60]) );
  AO222X1_HVT U721 ( .A1(n1661), .A2(sram_rdata_5[29]), .A3(n2140), .A4(
        sram_rdata_4[29]), .A5(sram_rdata_3[29]), .A6(n1690), .Y(n1531) );
  AO222X1_HVT U722 ( .A1(n1661), .A2(sram_rdata_2[29]), .A3(n15500), .A4(
        sram_rdata_1[29]), .A5(sram_rdata_0[29]), .A6(n1970), .Y(n11301) );
  AOI22X1_HVT U723 ( .A1(n1531), .A2(n15100), .A3(n14400), .A4(n11301), .Y(
        n783) );
  OA22X1_HVT U724 ( .A1(n11600), .A2(n411), .A3(n14600), .A4(n3150), .Y(n782)
         );
  NAND2X0_HVT U725 ( .A1(n1700), .A2(sram_rdata_6[29]), .Y(n781) );
  NAND3X0_HVT U726 ( .A1(n783), .A2(n782), .A3(n781), .Y(n_src_aox[61]) );
  AO222X1_HVT U727 ( .A1(n1860), .A2(sram_rdata_5[30]), .A3(n15600), .A4(
        sram_rdata_4[30]), .A5(sram_rdata_3[30]), .A6(n1900), .Y(n1533) );
  AO222X1_HVT U728 ( .A1(n1830), .A2(sram_rdata_2[30]), .A3(n2140), .A4(
        sram_rdata_1[30]), .A5(sram_rdata_0[30]), .A6(n1990), .Y(n1134) );
  AOI22X1_HVT U729 ( .A1(n1533), .A2(n12700), .A3(n5801), .A4(n1134), .Y(n786)
         );
  OA22X1_HVT U730 ( .A1(n2770), .A2(n412), .A3(n11400), .A4(n3160), .Y(n785)
         );
  NAND2X0_HVT U731 ( .A1(n1770), .A2(sram_rdata_6[30]), .Y(n784) );
  NAND3X0_HVT U732 ( .A1(n786), .A2(n785), .A3(n784), .Y(n_src_aox[62]) );
  AO222X1_HVT U733 ( .A1(n1820), .A2(sram_rdata_5[31]), .A3(n16100), .A4(
        sram_rdata_4[31]), .A5(sram_rdata_3[31]), .A6(n2000), .Y(n1538) );
  AO222X1_HVT U734 ( .A1(n1661), .A2(sram_rdata_2[31]), .A3(n2150), .A4(
        sram_rdata_1[31]), .A5(sram_rdata_0[31]), .A6(n1980), .Y(n1138) );
  AOI22X1_HVT U735 ( .A1(n1538), .A2(n591), .A3(n12900), .A4(n1138), .Y(n789)
         );
  OA22X1_HVT U736 ( .A1(n13900), .A2(n413), .A3(n2730), .A4(n3170), .Y(n788)
         );
  NAND2X0_HVT U737 ( .A1(n576), .A2(sram_rdata_6[31]), .Y(n787) );
  NAND3X0_HVT U738 ( .A1(n789), .A2(n788), .A3(n787), .Y(n_src_aox[63]) );
  AO222X1_HVT U739 ( .A1(n2090), .A2(sram_rdata_4[16]), .A3(n589), .A4(
        sram_rdata_3[16]), .A5(sram_rdata_5[16]), .A6(n1900), .Y(n1543) );
  AO222X1_HVT U740 ( .A1(n1890), .A2(sram_rdata_1[16]), .A3(n588), .A4(
        sram_rdata_0[16]), .A5(sram_rdata_2[16]), .A6(n1920), .Y(n1142) );
  AOI22X1_HVT U741 ( .A1(n1543), .A2(n10800), .A3(n12500), .A4(n1142), .Y(n792) );
  OA22X1_HVT U742 ( .A1(n10400), .A2(n494), .A3(n2750), .A4(n398), .Y(n791) );
  NAND2X0_HVT U743 ( .A1(n575), .A2(sram_rdata_8[16]), .Y(n7901) );
  NAND3X0_HVT U744 ( .A1(n792), .A2(n791), .A3(n7901), .Y(n_src_aox[64]) );
  AO222X1_HVT U745 ( .A1(n2060), .A2(sram_rdata_4[17]), .A3(n2110), .A4(
        sram_rdata_3[17]), .A5(sram_rdata_5[17]), .A6(n1920), .Y(n1545) );
  AO222X1_HVT U746 ( .A1(n1870), .A2(sram_rdata_1[17]), .A3(n15700), .A4(
        sram_rdata_0[17]), .A5(sram_rdata_2[17]), .A6(n16500), .Y(n1146) );
  AOI22X1_HVT U747 ( .A1(n1545), .A2(n591), .A3(n11100), .A4(n1146), .Y(n795)
         );
  OA22X1_HVT U748 ( .A1(n10300), .A2(n495), .A3(n2700), .A4(n399), .Y(n794) );
  NAND2X0_HVT U749 ( .A1(n575), .A2(sram_rdata_8[17]), .Y(n793) );
  NAND3X0_HVT U750 ( .A1(n795), .A2(n794), .A3(n793), .Y(n_src_aox[65]) );
  AO222X1_HVT U751 ( .A1(n1830), .A2(sram_rdata_4[18]), .A3(n2200), .A4(
        sram_rdata_3[18]), .A5(sram_rdata_5[18]), .A6(n16400), .Y(n1547) );
  AO222X1_HVT U752 ( .A1(n2030), .A2(sram_rdata_1[18]), .A3(n589), .A4(
        sram_rdata_0[18]), .A5(sram_rdata_2[18]), .A6(n16500), .Y(n11501) );
  AOI22X1_HVT U753 ( .A1(n1547), .A2(n15100), .A3(n583), .A4(n11501), .Y(n798)
         );
  OA22X1_HVT U754 ( .A1(n13800), .A2(n496), .A3(n14700), .A4(n4001), .Y(n797)
         );
  NAND2X0_HVT U755 ( .A1(n2240), .A2(sram_rdata_8[18]), .Y(n796) );
  NAND3X0_HVT U756 ( .A1(n798), .A2(n797), .A3(n796), .Y(n_src_aox[66]) );
  AO222X1_HVT U757 ( .A1(n1890), .A2(sram_rdata_4[19]), .A3(n2110), .A4(
        sram_rdata_3[19]), .A5(sram_rdata_5[19]), .A6(n2010), .Y(n1552) );
  AO222X1_HVT U758 ( .A1(n1830), .A2(sram_rdata_1[19]), .A3(n15600), .A4(
        sram_rdata_0[19]), .A5(sram_rdata_2[19]), .A6(n16600), .Y(n1154) );
  AOI22X1_HVT U759 ( .A1(n1552), .A2(n5901), .A3(n5801), .A4(n1154), .Y(n801)
         );
  OA22X1_HVT U760 ( .A1(n2770), .A2(n497), .A3(n2720), .A4(n401), .Y(n8001) );
  NAND2X0_HVT U761 ( .A1(n2210), .A2(sram_rdata_8[19]), .Y(n799) );
  NAND3X0_HVT U762 ( .A1(n801), .A2(n8001), .A3(n799), .Y(n_src_aox[67]) );
  AO222X1_HVT U763 ( .A1(n1840), .A2(sram_rdata_4[20]), .A3(n16000), .A4(
        sram_rdata_3[20]), .A5(sram_rdata_5[20]), .A6(n2010), .Y(n1557) );
  AO222X1_HVT U764 ( .A1(n1661), .A2(sram_rdata_1[20]), .A3(n2130), .A4(
        sram_rdata_0[20]), .A5(sram_rdata_2[20]), .A6(n1960), .Y(n1158) );
  AOI22X1_HVT U765 ( .A1(n1557), .A2(n15000), .A3(n12400), .A4(n1158), .Y(n804) );
  OA22X1_HVT U766 ( .A1(n2800), .A2(n498), .A3(n10000), .A4(n402), .Y(n803) );
  NAND2X0_HVT U767 ( .A1(n577), .A2(sram_rdata_8[20]), .Y(n802) );
  NAND3X0_HVT U768 ( .A1(n804), .A2(n803), .A3(n802), .Y(n_src_aox[68]) );
  AO222X1_HVT U769 ( .A1(n1830), .A2(sram_rdata_4[21]), .A3(n589), .A4(
        sram_rdata_3[21]), .A5(sram_rdata_5[21]), .A6(n2020), .Y(n1562) );
  AO222X1_HVT U770 ( .A1(n2070), .A2(sram_rdata_1[21]), .A3(n589), .A4(
        sram_rdata_0[21]), .A5(sram_rdata_2[21]), .A6(n1950), .Y(n1162) );
  AOI22X1_HVT U771 ( .A1(n1562), .A2(n12700), .A3(n582), .A4(n1162), .Y(n807)
         );
  OA22X1_HVT U772 ( .A1(n2790), .A2(n499), .A3(n11400), .A4(n403), .Y(n806) );
  NAND2X0_HVT U773 ( .A1(n578), .A2(sram_rdata_8[21]), .Y(n805) );
  NAND3X0_HVT U774 ( .A1(n807), .A2(n806), .A3(n805), .Y(n_src_aox[69]) );
  AO222X1_HVT U775 ( .A1(n2070), .A2(sram_rdata_4[22]), .A3(n15900), .A4(
        sram_rdata_3[22]), .A5(sram_rdata_5[22]), .A6(n1910), .Y(n1564) );
  AO222X1_HVT U776 ( .A1(n2100), .A2(sram_rdata_1[22]), .A3(n2200), .A4(
        sram_rdata_0[22]), .A5(sram_rdata_2[22]), .A6(n16300), .Y(n1166) );
  AOI22X1_HVT U777 ( .A1(n1564), .A2(n12800), .A3(n11000), .A4(n1166), .Y(
        n8101) );
  OA22X1_HVT U778 ( .A1(n10200), .A2(n5001), .A3(n2710), .A4(n404), .Y(n809)
         );
  NAND2X0_HVT U779 ( .A1(n1790), .A2(sram_rdata_8[22]), .Y(n808) );
  NAND3X0_HVT U780 ( .A1(n8101), .A2(n809), .A3(n808), .Y(n_src_aox[70]) );
  AO222X1_HVT U781 ( .A1(n2100), .A2(sram_rdata_4[23]), .A3(n15600), .A4(
        sram_rdata_3[23]), .A5(sram_rdata_5[23]), .A6(n1900), .Y(n1566) );
  AO222X1_HVT U782 ( .A1(n2090), .A2(sram_rdata_1[23]), .A3(n589), .A4(
        sram_rdata_0[23]), .A5(sram_rdata_2[23]), .A6(n16600), .Y(n11701) );
  AOI22X1_HVT U783 ( .A1(n1566), .A2(n591), .A3(n583), .A4(n11701), .Y(n813)
         );
  OA22X1_HVT U784 ( .A1(n13700), .A2(n501), .A3(n2740), .A4(n405), .Y(n812) );
  NAND2X0_HVT U785 ( .A1(n1790), .A2(sram_rdata_8[23]), .Y(n811) );
  NAND3X0_HVT U786 ( .A1(n813), .A2(n812), .A3(n811), .Y(n_src_aox[71]) );
  AO222X1_HVT U787 ( .A1(n1820), .A2(sram_rdata_4[24]), .A3(n2170), .A4(
        sram_rdata_3[24]), .A5(sram_rdata_5[24]), .A6(n1930), .Y(n1571) );
  AO222X1_HVT U788 ( .A1(n2040), .A2(sram_rdata_1[24]), .A3(n2170), .A4(
        sram_rdata_0[24]), .A5(sram_rdata_2[24]), .A6(n1950), .Y(n1174) );
  AOI22X1_HVT U789 ( .A1(n1571), .A2(n1664), .A3(n12400), .A4(n1174), .Y(n816)
         );
  OA22X1_HVT U790 ( .A1(n13800), .A2(n502), .A3(n10000), .A4(n406), .Y(n815)
         );
  NAND2X0_HVT U791 ( .A1(n1730), .A2(sram_rdata_8[24]), .Y(n814) );
  NAND3X0_HVT U792 ( .A1(n816), .A2(n815), .A3(n814), .Y(n_src_aox[72]) );
  AO222X1_HVT U793 ( .A1(n1820), .A2(sram_rdata_4[25]), .A3(n2180), .A4(
        sram_rdata_3[25]), .A5(sram_rdata_5[25]), .A6(n16300), .Y(n1573) );
  AO222X1_HVT U794 ( .A1(n1830), .A2(sram_rdata_1[25]), .A3(n15500), .A4(
        sram_rdata_0[25]), .A5(sram_rdata_2[25]), .A6(n16400), .Y(n1178) );
  AOI22X1_HVT U795 ( .A1(n1573), .A2(n1664), .A3(n11100), .A4(n1178), .Y(n819)
         );
  OA22X1_HVT U796 ( .A1(n2810), .A2(n503), .A3(n10100), .A4(n407), .Y(n818) );
  NAND2X0_HVT U797 ( .A1(n2270), .A2(sram_rdata_8[25]), .Y(n817) );
  NAND3X0_HVT U798 ( .A1(n819), .A2(n818), .A3(n817), .Y(n_src_aox[73]) );
  AO222X1_HVT U799 ( .A1(n2100), .A2(sram_rdata_4[26]), .A3(n589), .A4(
        sram_rdata_3[26]), .A5(sram_rdata_5[26]), .A6(n2010), .Y(n1578) );
  AO222X1_HVT U800 ( .A1(n1820), .A2(sram_rdata_1[26]), .A3(n2150), .A4(
        sram_rdata_0[26]), .A5(sram_rdata_2[26]), .A6(n1680), .Y(n1182) );
  AOI22X1_HVT U801 ( .A1(n1578), .A2(n15100), .A3(n11000), .A4(n1182), .Y(n822) );
  OA22X1_HVT U802 ( .A1(n2760), .A2(n504), .A3(n11400), .A4(n408), .Y(n821) );
  NAND2X0_HVT U803 ( .A1(n576), .A2(sram_rdata_8[26]), .Y(n8201) );
  NAND3X0_HVT U804 ( .A1(n822), .A2(n821), .A3(n8201), .Y(n_src_aox[74]) );
  AO222X1_HVT U805 ( .A1(n1830), .A2(sram_rdata_4[27]), .A3(n15900), .A4(
        sram_rdata_3[27]), .A5(sram_rdata_5[27]), .A6(n1990), .Y(n15801) );
  AO222X1_HVT U806 ( .A1(n14000), .A2(sram_rdata_1[27]), .A3(n15900), .A4(
        sram_rdata_0[27]), .A5(sram_rdata_2[27]), .A6(n1970), .Y(n1186) );
  AOI22X1_HVT U807 ( .A1(n15801), .A2(n592), .A3(n12500), .A4(n1186), .Y(n825)
         );
  OA22X1_HVT U808 ( .A1(n10200), .A2(n505), .A3(n14900), .A4(n409), .Y(n824)
         );
  NAND2X0_HVT U809 ( .A1(n1790), .A2(sram_rdata_8[27]), .Y(n823) );
  NAND3X0_HVT U810 ( .A1(n825), .A2(n824), .A3(n823), .Y(n_src_aox[75]) );
  AO222X1_HVT U811 ( .A1(n2080), .A2(sram_rdata_4[28]), .A3(n15900), .A4(
        sram_rdata_3[28]), .A5(sram_rdata_5[28]), .A6(n1930), .Y(n1582) );
  AO222X1_HVT U812 ( .A1(n2050), .A2(sram_rdata_1[28]), .A3(n2140), .A4(
        sram_rdata_0[28]), .A5(sram_rdata_2[28]), .A6(n2020), .Y(n11901) );
  AOI22X1_HVT U813 ( .A1(n1582), .A2(n10800), .A3(n582), .A4(n11901), .Y(n828)
         );
  OA22X1_HVT U814 ( .A1(n10300), .A2(n506), .A3(n2740), .A4(n4101), .Y(n827)
         );
  NAND2X0_HVT U815 ( .A1(n1740), .A2(sram_rdata_8[28]), .Y(n826) );
  NAND3X0_HVT U816 ( .A1(n828), .A2(n827), .A3(n826), .Y(n_src_aox[76]) );
  AO222X1_HVT U817 ( .A1(n2030), .A2(sram_rdata_4[29]), .A3(n16000), .A4(
        sram_rdata_3[29]), .A5(sram_rdata_5[29]), .A6(n2010), .Y(n1584) );
  AO222X1_HVT U818 ( .A1(n2060), .A2(sram_rdata_1[29]), .A3(n15500), .A4(
        sram_rdata_0[29]), .A5(sram_rdata_2[29]), .A6(n1980), .Y(n1194) );
  AOI22X1_HVT U819 ( .A1(n1584), .A2(n593), .A3(n10700), .A4(n1194), .Y(n831)
         );
  OA22X1_HVT U820 ( .A1(n10400), .A2(n507), .A3(n14700), .A4(n411), .Y(n8301)
         );
  NAND2X0_HVT U821 ( .A1(n1740), .A2(sram_rdata_8[29]), .Y(n829) );
  NAND3X0_HVT U822 ( .A1(n831), .A2(n8301), .A3(n829), .Y(n_src_aox[77]) );
  AO222X1_HVT U823 ( .A1(n14000), .A2(sram_rdata_4[30]), .A3(n2190), .A4(
        sram_rdata_3[30]), .A5(sram_rdata_5[30]), .A6(n1670), .Y(n1589) );
  AO222X1_HVT U824 ( .A1(n2060), .A2(sram_rdata_1[30]), .A3(n2150), .A4(
        sram_rdata_0[30]), .A5(sram_rdata_2[30]), .A6(n1690), .Y(n1195) );
  AOI22X1_HVT U825 ( .A1(n1589), .A2(n592), .A3(n582), .A4(n1195), .Y(n834) );
  OA22X1_HVT U826 ( .A1(n13700), .A2(n508), .A3(n10000), .A4(n412), .Y(n833)
         );
  NAND2X0_HVT U827 ( .A1(n2270), .A2(sram_rdata_8[30]), .Y(n832) );
  NAND3X0_HVT U828 ( .A1(n834), .A2(n833), .A3(n832), .Y(n_src_aox[78]) );
  AO222X1_HVT U829 ( .A1(n1840), .A2(sram_rdata_4[31]), .A3(n2140), .A4(
        sram_rdata_3[31]), .A5(sram_rdata_5[31]), .A6(n16600), .Y(n1594) );
  AO222X1_HVT U830 ( .A1(n1840), .A2(sram_rdata_1[31]), .A3(n16000), .A4(
        sram_rdata_0[31]), .A5(sram_rdata_2[31]), .A6(n1950), .Y(n1196) );
  AOI22X1_HVT U831 ( .A1(n1594), .A2(n10900), .A3(n5801), .A4(n1196), .Y(n837)
         );
  OA22X1_HVT U832 ( .A1(n13700), .A2(n509), .A3(n10000), .A4(n413), .Y(n836)
         );
  NAND2X0_HVT U833 ( .A1(n577), .A2(sram_rdata_8[31]), .Y(n835) );
  NAND3X0_HVT U834 ( .A1(n837), .A2(n836), .A3(n835), .Y(n_src_aox[79]) );
  AO222X1_HVT U835 ( .A1(n1661), .A2(sram_rdata_3[16]), .A3(n2130), .A4(
        sram_rdata_5[16]), .A5(n1980), .A6(sram_rdata_4[16]), .Y(n1599) );
  AO222X1_HVT U836 ( .A1(n1870), .A2(sram_rdata_0[16]), .A3(n2130), .A4(
        sram_rdata_2[16]), .A5(n2020), .A6(sram_rdata_1[16]), .Y(n12001) );
  AOI22X1_HVT U837 ( .A1(n1599), .A2(n591), .A3(n583), .A4(n12001), .Y(n8401)
         );
  OA22X1_HVT U838 ( .A1(n11600), .A2(n3020), .A3(n2740), .A4(n494), .Y(n839)
         );
  NAND2X0_HVT U839 ( .A1(n2270), .A2(sram_rdata_7[16]), .Y(n838) );
  NAND3X0_HVT U840 ( .A1(n8401), .A2(n839), .A3(n838), .Y(n_src_aox[80]) );
  AO222X1_HVT U841 ( .A1(n1860), .A2(sram_rdata_3[17]), .A3(n15400), .A4(
        sram_rdata_5[17]), .A5(n1960), .A6(sram_rdata_4[17]), .Y(n1604) );
  AO222X1_HVT U842 ( .A1(n1880), .A2(sram_rdata_0[17]), .A3(n2110), .A4(
        sram_rdata_2[17]), .A5(n1930), .A6(sram_rdata_1[17]), .Y(n1204) );
  AOI22X1_HVT U843 ( .A1(n1604), .A2(n10800), .A3(n12900), .A4(n1204), .Y(n843) );
  OA22X1_HVT U844 ( .A1(n11700), .A2(n3030), .A3(n2710), .A4(n495), .Y(n842)
         );
  NAND2X0_HVT U845 ( .A1(n2220), .A2(sram_rdata_7[17]), .Y(n841) );
  NAND3X0_HVT U846 ( .A1(n843), .A2(n842), .A3(n841), .Y(n_src_aox[81]) );
  AO222X1_HVT U847 ( .A1(n2090), .A2(sram_rdata_3[18]), .A3(n589), .A4(
        sram_rdata_5[18]), .A5(n2010), .A6(sram_rdata_4[18]), .Y(n1609) );
  AO222X1_HVT U848 ( .A1(n12600), .A2(sram_rdata_0[18]), .A3(n16200), .A4(
        sram_rdata_2[18]), .A5(n2000), .A6(sram_rdata_1[18]), .Y(n1208) );
  AOI22X1_HVT U849 ( .A1(n1609), .A2(n12800), .A3(n5801), .A4(n1208), .Y(n846)
         );
  OA22X1_HVT U850 ( .A1(n13800), .A2(n3040), .A3(n2690), .A4(n496), .Y(n845)
         );
  NAND2X0_HVT U851 ( .A1(n575), .A2(sram_rdata_7[18]), .Y(n844) );
  NAND3X0_HVT U852 ( .A1(n846), .A2(n845), .A3(n844), .Y(n_src_aox[82]) );
  AO222X1_HVT U853 ( .A1(n1860), .A2(sram_rdata_3[19]), .A3(n2190), .A4(
        sram_rdata_5[19]), .A5(n1970), .A6(sram_rdata_4[19]), .Y(n1611) );
  AO222X1_HVT U854 ( .A1(n12600), .A2(sram_rdata_0[19]), .A3(n16200), .A4(
        sram_rdata_2[19]), .A5(n1970), .A6(sram_rdata_1[19]), .Y(n1212) );
  AOI22X1_HVT U855 ( .A1(n1611), .A2(n5901), .A3(n11100), .A4(n1212), .Y(n849)
         );
  OA22X1_HVT U856 ( .A1(n2770), .A2(n3050), .A3(n14800), .A4(n497), .Y(n848)
         );
  NAND2X0_HVT U857 ( .A1(n2260), .A2(sram_rdata_7[19]), .Y(n847) );
  NAND3X0_HVT U858 ( .A1(n849), .A2(n848), .A3(n847), .Y(n_src_aox[83]) );
  AO222X1_HVT U859 ( .A1(n1820), .A2(sram_rdata_3[20]), .A3(n2180), .A4(
        sram_rdata_5[20]), .A5(n16400), .A6(sram_rdata_4[20]), .Y(n1616) );
  AO222X1_HVT U860 ( .A1(n2030), .A2(sram_rdata_0[20]), .A3(n16100), .A4(
        sram_rdata_2[20]), .A5(n1930), .A6(sram_rdata_1[20]), .Y(n1216) );
  AOI22X1_HVT U861 ( .A1(n1616), .A2(n10900), .A3(n10700), .A4(n1216), .Y(n852) );
  OA22X1_HVT U862 ( .A1(n2810), .A2(n3060), .A3(n14900), .A4(n498), .Y(n851)
         );
  NAND2X0_HVT U863 ( .A1(n1700), .A2(sram_rdata_7[20]), .Y(n8501) );
  NAND3X0_HVT U864 ( .A1(n852), .A2(n851), .A3(n8501), .Y(n_src_aox[84]) );
  AO222X1_HVT U865 ( .A1(n1890), .A2(sram_rdata_3[21]), .A3(n15400), .A4(
        sram_rdata_5[21]), .A5(n1980), .A6(sram_rdata_4[21]), .Y(n1618) );
  AO222X1_HVT U866 ( .A1(n12600), .A2(sram_rdata_0[21]), .A3(n15400), .A4(
        sram_rdata_2[21]), .A5(n1900), .A6(sram_rdata_1[21]), .Y(n12201) );
  AOI22X1_HVT U867 ( .A1(n1618), .A2(n1664), .A3(n11000), .A4(n12201), .Y(n855) );
  OA22X1_HVT U868 ( .A1(n2790), .A2(n3070), .A3(n2700), .A4(n499), .Y(n854) );
  NAND2X0_HVT U869 ( .A1(n1750), .A2(sram_rdata_7[21]), .Y(n853) );
  NAND3X0_HVT U870 ( .A1(n855), .A2(n854), .A3(n853), .Y(n_src_aox[85]) );
  AO222X1_HVT U871 ( .A1(n1890), .A2(sram_rdata_3[22]), .A3(n15500), .A4(
        sram_rdata_5[22]), .A5(n16500), .A6(sram_rdata_4[22]), .Y(n1623) );
  AO222X1_HVT U872 ( .A1(n1870), .A2(sram_rdata_0[22]), .A3(n2130), .A4(
        sram_rdata_2[22]), .A5(n2010), .A6(sram_rdata_1[22]), .Y(n1224) );
  AOI22X1_HVT U873 ( .A1(n1623), .A2(n12700), .A3(n581), .A4(n1224), .Y(n858)
         );
  OA22X1_HVT U874 ( .A1(n11800), .A2(n3080), .A3(n14600), .A4(n5001), .Y(n857)
         );
  NAND2X0_HVT U875 ( .A1(n578), .A2(sram_rdata_7[22]), .Y(n856) );
  NAND3X0_HVT U876 ( .A1(n858), .A2(n857), .A3(n856), .Y(n_src_aox[86]) );
  AO222X1_HVT U877 ( .A1(n14000), .A2(sram_rdata_3[23]), .A3(n15900), .A4(
        sram_rdata_5[23]), .A5(n1960), .A6(sram_rdata_4[23]), .Y(n1628) );
  AO222X1_HVT U878 ( .A1(n1890), .A2(sram_rdata_0[23]), .A3(n16100), .A4(
        sram_rdata_2[23]), .A5(n1930), .A6(sram_rdata_1[23]), .Y(n1228) );
  AOI22X1_HVT U879 ( .A1(n1628), .A2(n592), .A3(n10700), .A4(n1228), .Y(n861)
         );
  OA22X1_HVT U880 ( .A1(n2760), .A2(n3090), .A3(n2720), .A4(n501), .Y(n8601)
         );
  NAND2X0_HVT U881 ( .A1(n2260), .A2(sram_rdata_7[23]), .Y(n859) );
  NAND3X0_HVT U882 ( .A1(n861), .A2(n8601), .A3(n859), .Y(n_src_aox[87]) );
  AO222X1_HVT U883 ( .A1(n2070), .A2(sram_rdata_3[24]), .A3(n2180), .A4(
        sram_rdata_5[24]), .A5(n1920), .A6(sram_rdata_4[24]), .Y(n16301) );
  AO222X1_HVT U884 ( .A1(n2080), .A2(sram_rdata_0[24]), .A3(n2180), .A4(
        sram_rdata_2[24]), .A5(n1930), .A6(sram_rdata_1[24]), .Y(n1232) );
  AOI22X1_HVT U885 ( .A1(n16301), .A2(n10800), .A3(n581), .A4(n1232), .Y(n864)
         );
  OA22X1_HVT U886 ( .A1(n2790), .A2(n3100), .A3(n2720), .A4(n502), .Y(n863) );
  NAND2X0_HVT U887 ( .A1(n574), .A2(sram_rdata_7[24]), .Y(n862) );
  NAND3X0_HVT U888 ( .A1(n864), .A2(n863), .A3(n862), .Y(n_src_aox[88]) );
  AO222X1_HVT U889 ( .A1(n2090), .A2(sram_rdata_3[25]), .A3(n588), .A4(
        sram_rdata_5[25]), .A5(n1680), .A6(sram_rdata_4[25]), .Y(n1632) );
  AO222X1_HVT U890 ( .A1(n2100), .A2(sram_rdata_0[25]), .A3(n15600), .A4(
        sram_rdata_2[25]), .A5(n1970), .A6(sram_rdata_1[25]), .Y(n1236) );
  AOI22X1_HVT U891 ( .A1(n1632), .A2(n10900), .A3(n12400), .A4(n1236), .Y(n867) );
  OA22X1_HVT U892 ( .A1(n2800), .A2(n3110), .A3(n14600), .A4(n503), .Y(n866)
         );
  NAND2X0_HVT U893 ( .A1(n2220), .A2(sram_rdata_7[25]), .Y(n865) );
  NAND3X0_HVT U894 ( .A1(n867), .A2(n866), .A3(n865), .Y(n_src_aox[89]) );
  AO222X1_HVT U895 ( .A1(n1840), .A2(sram_rdata_3[26]), .A3(n2170), .A4(
        sram_rdata_5[26]), .A5(n16400), .A6(sram_rdata_4[26]), .Y(n1637) );
  AO222X1_HVT U896 ( .A1(n2030), .A2(sram_rdata_0[26]), .A3(n2200), .A4(
        sram_rdata_2[26]), .A5(n1670), .A6(sram_rdata_1[26]), .Y(n12401) );
  AOI22X1_HVT U897 ( .A1(n1637), .A2(n1664), .A3(n11000), .A4(n12401), .Y(
        n8701) );
  OA22X1_HVT U898 ( .A1(n2760), .A2(n3120), .A3(n14600), .A4(n504), .Y(n869)
         );
  NAND2X0_HVT U899 ( .A1(n1750), .A2(sram_rdata_7[26]), .Y(n868) );
  NAND3X0_HVT U900 ( .A1(n8701), .A2(n869), .A3(n868), .Y(n_src_aox[90]) );
  AO222X1_HVT U901 ( .A1(n2050), .A2(sram_rdata_3[27]), .A3(n2190), .A4(
        sram_rdata_5[27]), .A5(n1910), .A6(sram_rdata_4[27]), .Y(n1642) );
  AO222X1_HVT U902 ( .A1(n1840), .A2(sram_rdata_0[27]), .A3(n588), .A4(
        sram_rdata_2[27]), .A5(n1990), .A6(sram_rdata_1[27]), .Y(n1241) );
  AOI22X1_HVT U903 ( .A1(n1642), .A2(n591), .A3(n12900), .A4(n1241), .Y(n873)
         );
  OA22X1_HVT U904 ( .A1(n11800), .A2(n3130), .A3(n14900), .A4(n505), .Y(n872)
         );
  NAND2X0_HVT U905 ( .A1(n1780), .A2(sram_rdata_7[27]), .Y(n871) );
  NAND3X0_HVT U906 ( .A1(n873), .A2(n872), .A3(n871), .Y(n_src_aox[91]) );
  AO222X1_HVT U907 ( .A1(n1661), .A2(sram_rdata_3[28]), .A3(n15400), .A4(
        sram_rdata_5[28]), .A5(n1960), .A6(sram_rdata_4[28]), .Y(n1644) );
  AO222X1_HVT U908 ( .A1(n1860), .A2(sram_rdata_0[28]), .A3(n2160), .A4(
        sram_rdata_2[28]), .A5(n2020), .A6(sram_rdata_1[28]), .Y(n1242) );
  AOI22X1_HVT U909 ( .A1(n1644), .A2(n15100), .A3(n12400), .A4(n1242), .Y(n876) );
  OA22X1_HVT U910 ( .A1(n11700), .A2(n3140), .A3(n10000), .A4(n506), .Y(n875)
         );
  NAND2X0_HVT U911 ( .A1(n2240), .A2(sram_rdata_7[28]), .Y(n874) );
  NAND3X0_HVT U912 ( .A1(n876), .A2(n875), .A3(n874), .Y(n_src_aox[92]) );
  AO222X1_HVT U913 ( .A1(n1870), .A2(sram_rdata_3[29]), .A3(n15400), .A4(
        sram_rdata_5[29]), .A5(n1950), .A6(sram_rdata_4[29]), .Y(n1646) );
  AO222X1_HVT U914 ( .A1(n1880), .A2(sram_rdata_0[29]), .A3(n2110), .A4(
        sram_rdata_2[29]), .A5(n1900), .A6(sram_rdata_1[29]), .Y(n1243) );
  AOI22X1_HVT U915 ( .A1(n1646), .A2(n15100), .A3(n12400), .A4(n1243), .Y(n879) );
  OA22X1_HVT U916 ( .A1(n11600), .A2(n3150), .A3(n10100), .A4(n507), .Y(n878)
         );
  NAND2X0_HVT U917 ( .A1(n1790), .A2(sram_rdata_7[29]), .Y(n877) );
  NAND3X0_HVT U918 ( .A1(n879), .A2(n878), .A3(n877), .Y(n_src_aox[93]) );
  AO222X1_HVT U919 ( .A1(n2080), .A2(sram_rdata_3[30]), .A3(n16200), .A4(
        sram_rdata_5[30]), .A5(n1960), .A6(sram_rdata_4[30]), .Y(n1651) );
  AO222X1_HVT U920 ( .A1(n2030), .A2(sram_rdata_0[30]), .A3(n2160), .A4(
        sram_rdata_2[30]), .A5(n1920), .A6(sram_rdata_1[30]), .Y(n1247) );
  AOI22X1_HVT U921 ( .A1(n1651), .A2(n12800), .A3(n11000), .A4(n1247), .Y(n882) );
  OA22X1_HVT U922 ( .A1(n2780), .A2(n3160), .A3(n14700), .A4(n508), .Y(n881)
         );
  NAND2X0_HVT U923 ( .A1(n2250), .A2(sram_rdata_7[30]), .Y(n8801) );
  NAND3X0_HVT U924 ( .A1(n882), .A2(n881), .A3(n8801), .Y(n_src_aox[94]) );
  AO222X1_HVT U925 ( .A1(n2040), .A2(sram_rdata_3[31]), .A3(n2190), .A4(
        sram_rdata_5[31]), .A5(n1670), .A6(sram_rdata_4[31]), .Y(n1654) );
  AO222X1_HVT U926 ( .A1(n2040), .A2(sram_rdata_0[31]), .A3(n2130), .A4(
        sram_rdata_2[31]), .A5(n16400), .A6(sram_rdata_1[31]), .Y(n1251) );
  AOI22X1_HVT U927 ( .A1(n1654), .A2(n15000), .A3(n13000), .A4(n1251), .Y(n885) );
  OA22X1_HVT U928 ( .A1(n13900), .A2(n3170), .A3(n2740), .A4(n509), .Y(n884)
         );
  NAND2X0_HVT U929 ( .A1(n1780), .A2(sram_rdata_7[31]), .Y(n883) );
  NAND3X0_HVT U930 ( .A1(n885), .A2(n884), .A3(n883), .Y(n_src_aox[95]) );
  AO222X1_HVT U931 ( .A1(sram_rdata_6[0]), .A2(n1990), .A3(sram_rdata_8[0]), 
        .A4(n2100), .A5(sram_rdata_7[0]), .A6(n2200), .Y(n1256) );
  AOI22X1_HVT U932 ( .A1(n1256), .A2(n11000), .A3(n594), .A4(n886), .Y(n889)
         );
  OA22X1_HVT U933 ( .A1(n11600), .A2(n3180), .A3(n14800), .A4(n478), .Y(n888)
         );
  NAND2X0_HVT U934 ( .A1(n2220), .A2(sram_rdata_3[0]), .Y(n887) );
  NAND3X0_HVT U935 ( .A1(n889), .A2(n888), .A3(n887), .Y(n_src_aox[96]) );
  AO222X1_HVT U936 ( .A1(n1880), .A2(sram_rdata_8[1]), .A3(n2170), .A4(
        sram_rdata_7[1]), .A5(sram_rdata_6[1]), .A6(n1920), .Y(n1257) );
  AOI22X1_HVT U937 ( .A1(n8901), .A2(n15100), .A3(n5801), .A4(n1257), .Y(n893)
         );
  OA22X1_HVT U938 ( .A1(n10300), .A2(n3190), .A3(n2700), .A4(n5101), .Y(n892)
         );
  NAND2X0_HVT U939 ( .A1(n577), .A2(sram_rdata_3[1]), .Y(n891) );
  NAND3X0_HVT U940 ( .A1(n893), .A2(n892), .A3(n891), .Y(n_src_aox[97]) );
  AO222X1_HVT U941 ( .A1(n2040), .A2(sram_rdata_8[2]), .A3(n2140), .A4(
        sram_rdata_7[2]), .A5(sram_rdata_6[2]), .A6(n1690), .Y(n1262) );
  AOI22X1_HVT U942 ( .A1(n894), .A2(n10900), .A3(n12400), .A4(n1262), .Y(n897)
         );
  OA22X1_HVT U943 ( .A1(n13900), .A2(n3200), .A3(n10100), .A4(n511), .Y(n896)
         );
  NAND2X0_HVT U944 ( .A1(n1730), .A2(sram_rdata_3[2]), .Y(n895) );
  NAND3X0_HVT U945 ( .A1(n897), .A2(n896), .A3(n895), .Y(n_src_aox[98]) );
  AO222X1_HVT U946 ( .A1(n1870), .A2(sram_rdata_8[3]), .A3(n2140), .A4(
        sram_rdata_7[3]), .A5(sram_rdata_6[3]), .A6(n1990), .Y(n1264) );
  AOI22X1_HVT U947 ( .A1(n898), .A2(n15000), .A3(n13000), .A4(n1264), .Y(n901)
         );
  OA22X1_HVT U948 ( .A1(n2780), .A2(n3210), .A3(n2720), .A4(n512), .Y(n9001)
         );
  NAND2X0_HVT U949 ( .A1(n1760), .A2(sram_rdata_3[3]), .Y(n899) );
  NAND3X0_HVT U950 ( .A1(n901), .A2(n9001), .A3(n899), .Y(n_src_aox[99]) );
  AO222X1_HVT U951 ( .A1(n14000), .A2(sram_rdata_8[4]), .A3(n16100), .A4(
        sram_rdata_7[4]), .A5(sram_rdata_6[4]), .A6(n1980), .Y(n1269) );
  AOI22X1_HVT U952 ( .A1(n902), .A2(n10900), .A3(n11100), .A4(n1269), .Y(n905)
         );
  OA22X1_HVT U953 ( .A1(n2800), .A2(n3220), .A3(n14900), .A4(n513), .Y(n904)
         );
  NAND2X0_HVT U954 ( .A1(n1710), .A2(sram_rdata_3[4]), .Y(n903) );
  NAND3X0_HVT U955 ( .A1(n905), .A2(n904), .A3(n903), .Y(n_src_aox[100]) );
  AO222X1_HVT U956 ( .A1(n12600), .A2(sram_rdata_8[5]), .A3(n15600), .A4(
        sram_rdata_7[5]), .A5(sram_rdata_6[5]), .A6(n1910), .Y(n1274) );
  AOI22X1_HVT U957 ( .A1(n906), .A2(n10800), .A3(n581), .A4(n1274), .Y(n909)
         );
  OA22X1_HVT U958 ( .A1(n2790), .A2(n3230), .A3(n14700), .A4(n514), .Y(n908)
         );
  NAND2X0_HVT U959 ( .A1(n1700), .A2(sram_rdata_3[5]), .Y(n907) );
  NAND3X0_HVT U960 ( .A1(n909), .A2(n908), .A3(n907), .Y(n_src_aox[101]) );
  AO222X1_HVT U961 ( .A1(n1820), .A2(sram_rdata_8[6]), .A3(n2130), .A4(
        sram_rdata_7[6]), .A5(sram_rdata_6[6]), .A6(n1920), .Y(n1279) );
  AOI22X1_HVT U962 ( .A1(n9101), .A2(n593), .A3(n12900), .A4(n1279), .Y(n913)
         );
  OA22X1_HVT U963 ( .A1(n11800), .A2(n3240), .A3(n2700), .A4(n515), .Y(n912)
         );
  NAND2X0_HVT U964 ( .A1(n2240), .A2(sram_rdata_3[6]), .Y(n911) );
  NAND3X0_HVT U965 ( .A1(n913), .A2(n912), .A3(n911), .Y(n_src_aox[102]) );
  AO222X1_HVT U966 ( .A1(n1890), .A2(sram_rdata_8[7]), .A3(n15700), .A4(
        sram_rdata_7[7]), .A5(sram_rdata_6[7]), .A6(n16300), .Y(n1284) );
  AOI22X1_HVT U967 ( .A1(n914), .A2(n15100), .A3(n583), .A4(n1284), .Y(n917)
         );
  OA22X1_HVT U968 ( .A1(n13600), .A2(n3250), .A3(n2750), .A4(n516), .Y(n916)
         );
  NAND2X0_HVT U969 ( .A1(n2210), .A2(sram_rdata_3[7]), .Y(n915) );
  NAND3X0_HVT U970 ( .A1(n917), .A2(n916), .A3(n915), .Y(n_src_aox[103]) );
  AO222X1_HVT U971 ( .A1(n1840), .A2(sram_rdata_8[8]), .A3(n15700), .A4(
        sram_rdata_7[8]), .A5(sram_rdata_6[8]), .A6(n16500), .Y(n1289) );
  AOI22X1_HVT U972 ( .A1(n918), .A2(n15000), .A3(n581), .A4(n1289), .Y(n921)
         );
  OA22X1_HVT U973 ( .A1(n13900), .A2(n3260), .A3(n14800), .A4(n517), .Y(n9201)
         );
  NAND2X0_HVT U974 ( .A1(n578), .A2(sram_rdata_3[8]), .Y(n919) );
  NAND3X0_HVT U975 ( .A1(n921), .A2(n9201), .A3(n919), .Y(n_src_aox[104]) );
  AO222X1_HVT U976 ( .A1(n2090), .A2(sram_rdata_8[9]), .A3(n15700), .A4(
        sram_rdata_7[9]), .A5(sram_rdata_6[9]), .A6(n16400), .Y(n1294) );
  AOI22X1_HVT U977 ( .A1(n922), .A2(n15100), .A3(n12400), .A4(n1294), .Y(n925)
         );
  OA22X1_HVT U978 ( .A1(n2810), .A2(n327), .A3(n14600), .A4(n518), .Y(n924) );
  NAND2X0_HVT U979 ( .A1(n1710), .A2(sram_rdata_3[9]), .Y(n923) );
  NAND3X0_HVT U980 ( .A1(n925), .A2(n924), .A3(n923), .Y(n_src_aox[105]) );
  AO222X1_HVT U981 ( .A1(n1870), .A2(sram_rdata_8[10]), .A3(n16200), .A4(
        sram_rdata_7[10]), .A5(sram_rdata_6[10]), .A6(n16500), .Y(n1299) );
  AOI22X1_HVT U982 ( .A1(n926), .A2(n5901), .A3(n582), .A4(n1299), .Y(n929) );
  OA22X1_HVT U983 ( .A1(n13600), .A2(n328), .A3(n2710), .A4(n519), .Y(n928) );
  NAND2X0_HVT U984 ( .A1(n1760), .A2(sram_rdata_3[10]), .Y(n927) );
  NAND3X0_HVT U985 ( .A1(n929), .A2(n928), .A3(n927), .Y(n_src_aox[106]) );
  AO222X1_HVT U986 ( .A1(n1661), .A2(sram_rdata_8[11]), .A3(n16601), .A4(
        sram_rdata_7[11]), .A5(sram_rdata_6[11]), .A6(n1960), .Y(n1304) );
  AOI22X1_HVT U987 ( .A1(n9301), .A2(n12800), .A3(n581), .A4(n1304), .Y(n933)
         );
  OA22X1_HVT U988 ( .A1(n10200), .A2(n329), .A3(n2720), .A4(n5201), .Y(n932)
         );
  NAND2X0_HVT U989 ( .A1(n1790), .A2(sram_rdata_3[11]), .Y(n931) );
  NAND3X0_HVT U990 ( .A1(n933), .A2(n932), .A3(n931), .Y(n_src_aox[107]) );
  AO222X1_HVT U991 ( .A1(n2060), .A2(sram_rdata_8[12]), .A3(n2110), .A4(
        sram_rdata_7[12]), .A5(sram_rdata_6[12]), .A6(n2000), .Y(n1309) );
  AOI22X1_HVT U992 ( .A1(n934), .A2(n591), .A3(n12500), .A4(n1309), .Y(n937)
         );
  OA22X1_HVT U993 ( .A1(n10300), .A2(n330), .A3(n2750), .A4(n521), .Y(n936) );
  NAND2X0_HVT U994 ( .A1(n1740), .A2(sram_rdata_3[12]), .Y(n935) );
  NAND3X0_HVT U995 ( .A1(n937), .A2(n936), .A3(n935), .Y(n_src_aox[108]) );
  AO222X1_HVT U996 ( .A1(n1830), .A2(sram_rdata_8[13]), .A3(n2200), .A4(
        sram_rdata_7[13]), .A5(sram_rdata_6[13]), .A6(n2010), .Y(n1314) );
  AOI22X1_HVT U997 ( .A1(n938), .A2(n12800), .A3(n5801), .A4(n1314), .Y(n941)
         );
  OA22X1_HVT U998 ( .A1(n10400), .A2(n331), .A3(n2690), .A4(n522), .Y(n9401)
         );
  NAND2X0_HVT U999 ( .A1(n2270), .A2(sram_rdata_3[13]), .Y(n939) );
  NAND3X0_HVT U1000 ( .A1(n941), .A2(n9401), .A3(n939), .Y(n_src_aox[109]) );
  AO222X1_HVT U1001 ( .A1(n2030), .A2(sram_rdata_8[14]), .A3(n15700), .A4(
        sram_rdata_7[14]), .A5(sram_rdata_6[14]), .A6(n1970), .Y(n1319) );
  AOI22X1_HVT U1002 ( .A1(n942), .A2(n593), .A3(n12900), .A4(n1319), .Y(n945)
         );
  OA22X1_HVT U1003 ( .A1(n2770), .A2(n332), .A3(n14700), .A4(n523), .Y(n944)
         );
  NAND2X0_HVT U1004 ( .A1(n574), .A2(sram_rdata_3[14]), .Y(n943) );
  NAND3X0_HVT U1005 ( .A1(n945), .A2(n944), .A3(n943), .Y(n_src_aox[110]) );
  AO222X1_HVT U1006 ( .A1(n2040), .A2(sram_rdata_8[15]), .A3(n15600), .A4(
        sram_rdata_7[15]), .A5(sram_rdata_6[15]), .A6(n2020), .Y(n1324) );
  AOI22X1_HVT U1007 ( .A1(n946), .A2(n593), .A3(n12500), .A4(n1324), .Y(n949)
         );
  OA22X1_HVT U1008 ( .A1(n13800), .A2(n333), .A3(n2740), .A4(n524), .Y(n948)
         );
  NAND2X0_HVT U1009 ( .A1(n1800), .A2(sram_rdata_3[15]), .Y(n947) );
  NAND3X0_HVT U1010 ( .A1(n949), .A2(n948), .A3(n947), .Y(n_src_aox[111]) );
  AO222X1_HVT U1011 ( .A1(sram_rdata_6[0]), .A2(n2180), .A3(sram_rdata_8[0]), 
        .A4(n1690), .A5(n2070), .A6(sram_rdata_7[0]), .Y(n13301) );
  AOI22X1_HVT U1012 ( .A1(n13301), .A2(n13000), .A3(n594), .A4(n9501), .Y(n953) );
  OA22X1_HVT U1013 ( .A1(n10400), .A2(n382), .A3(n1662), .A4(n3180), .Y(n952)
         );
  NAND2X0_HVT U1014 ( .A1(n1750), .A2(sram_rdata_5[0]), .Y(n951) );
  NAND3X0_HVT U1015 ( .A1(n953), .A2(n952), .A3(n951), .Y(n_src_aox[112]) );
  AO222X1_HVT U1016 ( .A1(n2050), .A2(sram_rdata_7[1]), .A3(n15600), .A4(
        sram_rdata_6[1]), .A5(n1690), .A6(sram_rdata_8[1]), .Y(n1334) );
  AOI22X1_HVT U1017 ( .A1(n954), .A2(n15000), .A3(n583), .A4(n1334), .Y(n957)
         );
  OA22X1_HVT U1018 ( .A1(n11700), .A2(n414), .A3(n11400), .A4(n3190), .Y(n956)
         );
  NAND2X0_HVT U1019 ( .A1(n1770), .A2(sram_rdata_5[1]), .Y(n955) );
  NAND3X0_HVT U1020 ( .A1(n957), .A2(n956), .A3(n955), .Y(n_src_aox[113]) );
  AO222X1_HVT U1021 ( .A1(n1870), .A2(sram_rdata_7[2]), .A3(n15400), .A4(
        sram_rdata_6[2]), .A5(n1900), .A6(sram_rdata_8[2]), .Y(n1339) );
  AOI22X1_HVT U1022 ( .A1(n958), .A2(n12800), .A3(n5801), .A4(n1339), .Y(n961)
         );
  OA22X1_HVT U1023 ( .A1(n13800), .A2(n415), .A3(n14600), .A4(n3200), .Y(n9601) );
  NAND2X0_HVT U1024 ( .A1(n2260), .A2(sram_rdata_5[2]), .Y(n959) );
  NAND3X0_HVT U1025 ( .A1(n961), .A2(n9601), .A3(n959), .Y(n_src_aox[114]) );
  AO222X1_HVT U1026 ( .A1(n1880), .A2(sram_rdata_7[3]), .A3(n2140), .A4(
        sram_rdata_6[3]), .A5(n16300), .A6(sram_rdata_8[3]), .Y(n1344) );
  AOI22X1_HVT U1027 ( .A1(n962), .A2(n12700), .A3(n5801), .A4(n1344), .Y(n965)
         );
  OA22X1_HVT U1028 ( .A1(n2770), .A2(n416), .A3(n1662), .A4(n3210), .Y(n964)
         );
  NAND2X0_HVT U1029 ( .A1(n1700), .A2(sram_rdata_5[3]), .Y(n963) );
  NAND3X0_HVT U1030 ( .A1(n965), .A2(n964), .A3(n963), .Y(n_src_aox[115]) );
  AO222X1_HVT U1031 ( .A1(n2100), .A2(sram_rdata_7[4]), .A3(n16100), .A4(
        sram_rdata_6[4]), .A5(n16300), .A6(sram_rdata_8[4]), .Y(n1349) );
  AOI22X1_HVT U1032 ( .A1(n966), .A2(n594), .A3(n10700), .A4(n1349), .Y(n969)
         );
  OA22X1_HVT U1033 ( .A1(n2800), .A2(n417), .A3(n2720), .A4(n3220), .Y(n968)
         );
  NAND2X0_HVT U1034 ( .A1(n2250), .A2(sram_rdata_5[4]), .Y(n967) );
  NAND3X0_HVT U1035 ( .A1(n969), .A2(n968), .A3(n967), .Y(n_src_aox[116]) );
  AO222X1_HVT U1036 ( .A1(n14000), .A2(sram_rdata_7[5]), .A3(n2160), .A4(
        sram_rdata_6[5]), .A5(n1680), .A6(sram_rdata_8[5]), .Y(n1354) );
  AOI22X1_HVT U1037 ( .A1(n9701), .A2(n15000), .A3(n5801), .A4(n1354), .Y(n973) );
  OA22X1_HVT U1038 ( .A1(n2790), .A2(n418), .A3(n2690), .A4(n3230), .Y(n972)
         );
  NAND2X0_HVT U1039 ( .A1(n576), .A2(sram_rdata_5[5]), .Y(n971) );
  NAND3X0_HVT U1040 ( .A1(n973), .A2(n972), .A3(n971), .Y(n_src_aox[117]) );
  AO222X1_HVT U1041 ( .A1(n2080), .A2(sram_rdata_7[6]), .A3(n16601), .A4(
        sram_rdata_6[6]), .A5(n2010), .A6(sram_rdata_8[6]), .Y(n1356) );
  AOI22X1_HVT U1042 ( .A1(n974), .A2(n15000), .A3(n5801), .A4(n1356), .Y(n977)
         );
  OA22X1_HVT U1043 ( .A1(n10200), .A2(n419), .A3(n10100), .A4(n3240), .Y(n976)
         );
  NAND2X0_HVT U1044 ( .A1(n1710), .A2(sram_rdata_5[6]), .Y(n975) );
  NAND3X0_HVT U1045 ( .A1(n977), .A2(n976), .A3(n975), .Y(n_src_aox[118]) );
  AO222X1_HVT U1046 ( .A1(n2070), .A2(sram_rdata_7[7]), .A3(n2190), .A4(
        sram_rdata_6[7]), .A5(n1960), .A6(sram_rdata_8[7]), .Y(n1361) );
  AOI22X1_HVT U1047 ( .A1(n978), .A2(n594), .A3(n11100), .A4(n1361), .Y(n981)
         );
  OA22X1_HVT U1048 ( .A1(n13700), .A2(n4201), .A3(n2730), .A4(n3250), .Y(n9801) );
  NAND2X0_HVT U1049 ( .A1(n2240), .A2(sram_rdata_5[7]), .Y(n979) );
  NAND3X0_HVT U1050 ( .A1(n981), .A2(n9801), .A3(n979), .Y(n_src_aox[119]) );
  AO222X1_HVT U1051 ( .A1(n2070), .A2(sram_rdata_7[8]), .A3(n588), .A4(
        sram_rdata_6[8]), .A5(n1920), .A6(sram_rdata_8[8]), .Y(n1366) );
  AOI22X1_HVT U1052 ( .A1(n982), .A2(n10800), .A3(n583), .A4(n1366), .Y(n985)
         );
  OA22X1_HVT U1053 ( .A1(n13800), .A2(n421), .A3(n2730), .A4(n3260), .Y(n984)
         );
  NAND2X0_HVT U1054 ( .A1(n577), .A2(sram_rdata_5[8]), .Y(n983) );
  NAND3X0_HVT U1055 ( .A1(n985), .A2(n984), .A3(n983), .Y(n_src_aox[120]) );
  AO222X1_HVT U1056 ( .A1(n2070), .A2(sram_rdata_7[9]), .A3(n15900), .A4(
        sram_rdata_6[9]), .A5(n2000), .A6(sram_rdata_8[9]), .Y(n1371) );
  AOI22X1_HVT U1057 ( .A1(n986), .A2(n1664), .A3(n12900), .A4(n1371), .Y(n989)
         );
  OA22X1_HVT U1058 ( .A1(n13900), .A2(n422), .A3(n10100), .A4(n327), .Y(n988)
         );
  NAND2X0_HVT U1059 ( .A1(n1780), .A2(sram_rdata_5[9]), .Y(n987) );
  NAND3X0_HVT U1060 ( .A1(n989), .A2(n988), .A3(n987), .Y(n_src_aox[121]) );
  AO222X1_HVT U1061 ( .A1(n1820), .A2(sram_rdata_7[10]), .A3(n2200), .A4(
        sram_rdata_6[10]), .A5(n2020), .A6(sram_rdata_8[10]), .Y(n1376) );
  AOI22X1_HVT U1062 ( .A1(n9901), .A2(n593), .A3(n12500), .A4(n1376), .Y(n993)
         );
  OA22X1_HVT U1063 ( .A1(n2760), .A2(n423), .A3(n2690), .A4(n328), .Y(n992) );
  NAND2X0_HVT U1064 ( .A1(n575), .A2(sram_rdata_5[10]), .Y(n991) );
  NAND3X0_HVT U1065 ( .A1(n993), .A2(n992), .A3(n991), .Y(n_src_aox[122]) );
  AO222X1_HVT U1066 ( .A1(n2060), .A2(sram_rdata_7[11]), .A3(n2180), .A4(
        sram_rdata_6[11]), .A5(n1950), .A6(sram_rdata_8[11]), .Y(n1381) );
  AOI22X1_HVT U1067 ( .A1(n994), .A2(n593), .A3(n11000), .A4(n1381), .Y(n997)
         );
  OA22X1_HVT U1068 ( .A1(n11800), .A2(n424), .A3(n1662), .A4(n329), .Y(n996)
         );
  NAND2X0_HVT U1069 ( .A1(n2260), .A2(sram_rdata_5[11]), .Y(n995) );
  NAND3X0_HVT U1070 ( .A1(n997), .A2(n996), .A3(n995), .Y(n_src_aox[123]) );
  AO222X1_HVT U1071 ( .A1(n12600), .A2(sram_rdata_7[12]), .A3(n2190), .A4(
        sram_rdata_6[12]), .A5(n1670), .A6(sram_rdata_8[12]), .Y(n1386) );
  AOI22X1_HVT U1072 ( .A1(n998), .A2(n10900), .A3(n583), .A4(n1386), .Y(n1001)
         );
  OA22X1_HVT U1073 ( .A1(n11700), .A2(n425), .A3(n2740), .A4(n330), .Y(n10001)
         );
  NAND2X0_HVT U1074 ( .A1(n574), .A2(sram_rdata_5[12]), .Y(n999) );
  NAND3X0_HVT U1075 ( .A1(n1001), .A2(n10001), .A3(n999), .Y(n_src_aox[124])
         );
  AO222X1_HVT U1076 ( .A1(n14000), .A2(sram_rdata_7[13]), .A3(n16601), .A4(
        sram_rdata_6[13]), .A5(n16500), .A6(sram_rdata_8[13]), .Y(n1391) );
  AOI22X1_HVT U1077 ( .A1(n1002), .A2(n1664), .A3(n582), .A4(n1391), .Y(n1005)
         );
  OA22X1_HVT U1078 ( .A1(n10400), .A2(n426), .A3(n2710), .A4(n331), .Y(n1004)
         );
  NAND2X0_HVT U1079 ( .A1(n2220), .A2(sram_rdata_5[13]), .Y(n1003) );
  NAND3X0_HVT U1080 ( .A1(n1005), .A2(n1004), .A3(n1003), .Y(n_src_aox[125])
         );
  AO222X1_HVT U1081 ( .A1(n1810), .A2(sram_rdata_7[14]), .A3(n2110), .A4(
        sram_rdata_6[14]), .A5(n1690), .A6(sram_rdata_8[14]), .Y(n1396) );
  AOI22X1_HVT U1082 ( .A1(n1006), .A2(n12800), .A3(n582), .A4(n1396), .Y(n1009) );
  OA22X1_HVT U1083 ( .A1(n2780), .A2(n427), .A3(n11400), .A4(n332), .Y(n1008)
         );
  NAND2X0_HVT U1084 ( .A1(n1740), .A2(sram_rdata_5[14]), .Y(n1007) );
  NAND3X0_HVT U1085 ( .A1(n1009), .A2(n1008), .A3(n1007), .Y(n_src_aox[126])
         );
  AO222X1_HVT U1086 ( .A1(n12600), .A2(sram_rdata_7[15]), .A3(n2130), .A4(
        sram_rdata_6[15]), .A5(n1970), .A6(sram_rdata_8[15]), .Y(n1398) );
  AOI22X1_HVT U1087 ( .A1(n10101), .A2(n594), .A3(n13000), .A4(n1398), .Y(
        n1013) );
  OA22X1_HVT U1088 ( .A1(n13700), .A2(n428), .A3(n2730), .A4(n333), .Y(n1012)
         );
  NAND2X0_HVT U1089 ( .A1(n1800), .A2(sram_rdata_5[15]), .Y(n1011) );
  NAND3X0_HVT U1090 ( .A1(n1013), .A2(n1012), .A3(n1011), .Y(n_src_aox[127])
         );
  AO222X1_HVT U1091 ( .A1(sram_rdata_6[0]), .A2(n2080), .A3(sram_rdata_8[0]), 
        .A4(n2190), .A5(n1910), .A6(sram_rdata_7[0]), .Y(n1404) );
  AOI22X1_HVT U1092 ( .A1(n1404), .A2(n10700), .A3(n594), .A4(n1014), .Y(n1017) );
  OA22X1_HVT U1093 ( .A1(n11600), .A2(n478), .A3(n2750), .A4(n382), .Y(n1016)
         );
  NAND2X0_HVT U1094 ( .A1(n2210), .A2(sram_rdata_4[0]), .Y(n1015) );
  NAND3X0_HVT U1095 ( .A1(n1017), .A2(n1016), .A3(n1015), .Y(n_src_aox[128])
         );
  AO222X1_HVT U1096 ( .A1(n1661), .A2(sram_rdata_6[1]), .A3(n15400), .A4(
        sram_rdata_8[1]), .A5(sram_rdata_7[1]), .A6(n1960), .Y(n1405) );
  AOI22X1_HVT U1097 ( .A1(n1018), .A2(n591), .A3(n13000), .A4(n1405), .Y(n1021) );
  OA22X1_HVT U1098 ( .A1(n11700), .A2(n5101), .A3(n2700), .A4(n414), .Y(n10201) );
  NAND2X0_HVT U1099 ( .A1(n1790), .A2(sram_rdata_4[1]), .Y(n1019) );
  NAND3X0_HVT U1100 ( .A1(n1021), .A2(n10201), .A3(n1019), .Y(n_src_aox[129])
         );
  AO222X1_HVT U1101 ( .A1(n2090), .A2(sram_rdata_6[2]), .A3(n15400), .A4(
        sram_rdata_8[2]), .A5(sram_rdata_7[2]), .A6(n1910), .Y(n14101) );
  AOI22X1_HVT U1102 ( .A1(n1022), .A2(n591), .A3(n12900), .A4(n14101), .Y(
        n1025) );
  OA22X1_HVT U1103 ( .A1(n13600), .A2(n511), .A3(n14600), .A4(n415), .Y(n1024)
         );
  NAND2X0_HVT U1104 ( .A1(n2250), .A2(sram_rdata_4[2]), .Y(n1023) );
  NAND3X0_HVT U1105 ( .A1(n1025), .A2(n1024), .A3(n1023), .Y(n_src_aox[130])
         );
  AO222X1_HVT U1106 ( .A1(n2100), .A2(sram_rdata_6[3]), .A3(n588), .A4(
        sram_rdata_8[3]), .A5(sram_rdata_7[3]), .A6(n16400), .Y(n1415) );
  AOI22X1_HVT U1107 ( .A1(n1026), .A2(n12700), .A3(n13000), .A4(n1415), .Y(
        n1029) );
  OA22X1_HVT U1108 ( .A1(n2780), .A2(n512), .A3(n2730), .A4(n416), .Y(n1028)
         );
  NAND2X0_HVT U1109 ( .A1(n1750), .A2(sram_rdata_4[3]), .Y(n1027) );
  NAND3X0_HVT U1110 ( .A1(n1029), .A2(n1028), .A3(n1027), .Y(n_src_aox[131])
         );
  AO222X1_HVT U1111 ( .A1(n2050), .A2(sram_rdata_6[4]), .A3(n2160), .A4(
        sram_rdata_8[4]), .A5(sram_rdata_7[4]), .A6(n1930), .Y(n1417) );
  AOI22X1_HVT U1112 ( .A1(n10301), .A2(n10900), .A3(n582), .A4(n1417), .Y(
        n1033) );
  OA22X1_HVT U1113 ( .A1(n2810), .A2(n513), .A3(n1662), .A4(n417), .Y(n1032)
         );
  NAND2X0_HVT U1114 ( .A1(n2210), .A2(sram_rdata_4[4]), .Y(n1031) );
  NAND3X0_HVT U1115 ( .A1(n1033), .A2(n1032), .A3(n1031), .Y(n_src_aox[132])
         );
  AO222X1_HVT U1116 ( .A1(n2050), .A2(sram_rdata_6[5]), .A3(n588), .A4(
        sram_rdata_8[5]), .A5(sram_rdata_7[5]), .A6(n1680), .Y(n1422) );
  AOI22X1_HVT U1117 ( .A1(n1034), .A2(n10800), .A3(n12500), .A4(n1422), .Y(
        n1037) );
  OA22X1_HVT U1118 ( .A1(n2790), .A2(n514), .A3(n11400), .A4(n418), .Y(n1036)
         );
  NAND2X0_HVT U1119 ( .A1(n1700), .A2(sram_rdata_4[5]), .Y(n1035) );
  NAND3X0_HVT U1120 ( .A1(n1037), .A2(n1036), .A3(n1035), .Y(n_src_aox[133])
         );
  AO222X1_HVT U1121 ( .A1(n2030), .A2(sram_rdata_6[6]), .A3(n16200), .A4(
        sram_rdata_8[6]), .A5(sram_rdata_7[6]), .A6(n16500), .Y(n1427) );
  AOI22X1_HVT U1122 ( .A1(n1038), .A2(n593), .A3(n12500), .A4(n1427), .Y(n1041) );
  OA22X1_HVT U1123 ( .A1(n11800), .A2(n515), .A3(n2710), .A4(n419), .Y(n10401)
         );
  NAND2X0_HVT U1124 ( .A1(n1780), .A2(sram_rdata_4[6]), .Y(n1039) );
  NAND3X0_HVT U1125 ( .A1(n1041), .A2(n10401), .A3(n1039), .Y(n_src_aox[134])
         );
  AO222X1_HVT U1126 ( .A1(n2030), .A2(sram_rdata_6[7]), .A3(n2180), .A4(
        sram_rdata_8[7]), .A5(sram_rdata_7[7]), .A6(n1690), .Y(n1429) );
  AOI22X1_HVT U1127 ( .A1(n1042), .A2(n591), .A3(n582), .A4(n1429), .Y(n1045)
         );
  OA22X1_HVT U1128 ( .A1(n13600), .A2(n516), .A3(n14800), .A4(n4201), .Y(n1044) );
  NAND2X0_HVT U1129 ( .A1(n1740), .A2(sram_rdata_4[7]), .Y(n1043) );
  NAND3X0_HVT U1130 ( .A1(n1045), .A2(n1044), .A3(n1043), .Y(n_src_aox[135])
         );
  AO222X1_HVT U1131 ( .A1(n2060), .A2(sram_rdata_6[8]), .A3(n2130), .A4(
        sram_rdata_8[8]), .A5(sram_rdata_7[8]), .A6(n16300), .Y(n1434) );
  AOI22X1_HVT U1132 ( .A1(n1046), .A2(n591), .A3(n5801), .A4(n1434), .Y(n1049)
         );
  OA22X1_HVT U1133 ( .A1(n13800), .A2(n517), .A3(n10000), .A4(n421), .Y(n1048)
         );
  NAND2X0_HVT U1134 ( .A1(n578), .A2(sram_rdata_4[8]), .Y(n1047) );
  NAND3X0_HVT U1135 ( .A1(n1049), .A2(n1048), .A3(n1047), .Y(n_src_aox[136])
         );
  AO222X1_HVT U1136 ( .A1(n1810), .A2(sram_rdata_6[9]), .A3(n2160), .A4(
        sram_rdata_8[9]), .A5(sram_rdata_7[9]), .A6(n16500), .Y(n1439) );
  AOI22X1_HVT U1137 ( .A1(n10501), .A2(n593), .A3(n12500), .A4(n1439), .Y(
        n1053) );
  OA22X1_HVT U1138 ( .A1(n2800), .A2(n518), .A3(n10100), .A4(n422), .Y(n1052)
         );
  NAND2X0_HVT U1139 ( .A1(n578), .A2(sram_rdata_4[9]), .Y(n1051) );
  NAND3X0_HVT U1140 ( .A1(n1053), .A2(n1052), .A3(n1051), .Y(n_src_aox[137])
         );
  AO222X1_HVT U1141 ( .A1(n1880), .A2(sram_rdata_6[10]), .A3(n15600), .A4(
        sram_rdata_8[10]), .A5(sram_rdata_7[10]), .A6(n16600), .Y(n1444) );
  AOI22X1_HVT U1142 ( .A1(n1054), .A2(n593), .A3(n11100), .A4(n1444), .Y(n1057) );
  OA22X1_HVT U1143 ( .A1(n13600), .A2(n519), .A3(n11400), .A4(n423), .Y(n1056)
         );
  NAND2X0_HVT U1144 ( .A1(n2240), .A2(sram_rdata_4[10]), .Y(n1055) );
  NAND3X0_HVT U1145 ( .A1(n1057), .A2(n1056), .A3(n1055), .Y(n_src_aox[138])
         );
  AO222X1_HVT U1146 ( .A1(n1860), .A2(sram_rdata_6[11]), .A3(n16200), .A4(
        sram_rdata_8[11]), .A5(sram_rdata_7[11]), .A6(n1680), .Y(n1449) );
  AOI22X1_HVT U1147 ( .A1(n1058), .A2(n12800), .A3(n5801), .A4(n1449), .Y(
        n1061) );
  OA22X1_HVT U1148 ( .A1(n10200), .A2(n5201), .A3(n2730), .A4(n424), .Y(n10601) );
  NAND2X0_HVT U1149 ( .A1(n576), .A2(sram_rdata_4[11]), .Y(n1059) );
  NAND3X0_HVT U1150 ( .A1(n1061), .A2(n10601), .A3(n1059), .Y(n_src_aox[139])
         );
  AO222X1_HVT U1151 ( .A1(n2050), .A2(sram_rdata_6[12]), .A3(n2130), .A4(
        sram_rdata_8[12]), .A5(sram_rdata_7[12]), .A6(n1990), .Y(n1454) );
  AOI22X1_HVT U1152 ( .A1(n1062), .A2(n12700), .A3(n12900), .A4(n1454), .Y(
        n1065) );
  OA22X1_HVT U1153 ( .A1(n10300), .A2(n521), .A3(n2720), .A4(n425), .Y(n1064)
         );
  NAND2X0_HVT U1154 ( .A1(n1700), .A2(sram_rdata_4[12]), .Y(n1063) );
  NAND3X0_HVT U1155 ( .A1(n1065), .A2(n1064), .A3(n1063), .Y(n_src_aox[140])
         );
  AO222X1_HVT U1156 ( .A1(n12600), .A2(sram_rdata_6[13]), .A3(n2110), .A4(
        sram_rdata_8[13]), .A5(sram_rdata_7[13]), .A6(n1950), .Y(n1459) );
  AOI22X1_HVT U1157 ( .A1(n1066), .A2(n12700), .A3(n582), .A4(n1459), .Y(n1069) );
  OA22X1_HVT U1158 ( .A1(n11600), .A2(n522), .A3(n2710), .A4(n426), .Y(n1068)
         );
  NAND2X0_HVT U1159 ( .A1(n578), .A2(sram_rdata_4[13]), .Y(n1067) );
  NAND3X0_HVT U1160 ( .A1(n1069), .A2(n1068), .A3(n1067), .Y(n_src_aox[141])
         );
  AO222X1_HVT U1161 ( .A1(n1840), .A2(sram_rdata_6[14]), .A3(n2180), .A4(
        sram_rdata_8[14]), .A5(sram_rdata_7[14]), .A6(n1900), .Y(n1464) );
  AOI22X1_HVT U1162 ( .A1(n10701), .A2(n1664), .A3(n11000), .A4(n1464), .Y(
        n1073) );
  OA22X1_HVT U1163 ( .A1(n13600), .A2(n523), .A3(n10100), .A4(n427), .Y(n1072)
         );
  NAND2X0_HVT U1164 ( .A1(n1740), .A2(sram_rdata_4[14]), .Y(n1071) );
  NAND3X0_HVT U1165 ( .A1(n1073), .A2(n1072), .A3(n1071), .Y(n_src_aox[142])
         );
  AO222X1_HVT U1166 ( .A1(n2090), .A2(sram_rdata_6[15]), .A3(n15400), .A4(
        sram_rdata_8[15]), .A5(sram_rdata_7[15]), .A6(n2010), .Y(n1466) );
  AOI22X1_HVT U1167 ( .A1(n1074), .A2(n15100), .A3(n5801), .A4(n1466), .Y(
        n1077) );
  OA22X1_HVT U1168 ( .A1(n13700), .A2(n524), .A3(n2750), .A4(n428), .Y(n1076)
         );
  NAND2X0_HVT U1169 ( .A1(n1800), .A2(sram_rdata_4[15]), .Y(n1075) );
  NAND3X0_HVT U1170 ( .A1(n1077), .A2(n1076), .A3(n1075), .Y(n_src_aox[143])
         );
  AO222X1_HVT U1171 ( .A1(n1890), .A2(sram_rdata_8[16]), .A3(n15500), .A4(
        sram_rdata_7[16]), .A5(sram_rdata_6[16]), .A6(n1990), .Y(n1471) );
  AOI22X1_HVT U1172 ( .A1(n1078), .A2(n15000), .A3(n582), .A4(n1471), .Y(n1081) );
  OA22X1_HVT U1173 ( .A1(n11600), .A2(n334), .A3(n14900), .A4(n525), .Y(n10801) );
  NAND2X0_HVT U1174 ( .A1(n1740), .A2(sram_rdata_3[16]), .Y(n1079) );
  NAND3X0_HVT U1175 ( .A1(n1081), .A2(n10801), .A3(n1079), .Y(n_src_aox[144])
         );
  AO222X1_HVT U1176 ( .A1(n1860), .A2(sram_rdata_8[17]), .A3(n16100), .A4(
        sram_rdata_7[17]), .A5(sram_rdata_6[17]), .A6(n1970), .Y(n1476) );
  AOI22X1_HVT U1177 ( .A1(n1082), .A2(n10800), .A3(n5801), .A4(n1476), .Y(
        n1085) );
  OA22X1_HVT U1178 ( .A1(n11700), .A2(n335), .A3(n2690), .A4(n526), .Y(n1084)
         );
  NAND2X0_HVT U1179 ( .A1(n2270), .A2(sram_rdata_3[17]), .Y(n1083) );
  NAND3X0_HVT U1180 ( .A1(n1085), .A2(n1084), .A3(n1083), .Y(n_src_aox[145])
         );
  AO222X1_HVT U1181 ( .A1(n1880), .A2(sram_rdata_8[18]), .A3(n15400), .A4(
        sram_rdata_7[18]), .A5(sram_rdata_6[18]), .A6(n1670), .Y(n1481) );
  AOI22X1_HVT U1182 ( .A1(n1086), .A2(n593), .A3(n582), .A4(n1481), .Y(n1089)
         );
  OA22X1_HVT U1183 ( .A1(n13700), .A2(n336), .A3(n2690), .A4(n527), .Y(n1088)
         );
  NAND2X0_HVT U1184 ( .A1(n576), .A2(sram_rdata_3[18]), .Y(n1087) );
  NAND3X0_HVT U1185 ( .A1(n1089), .A2(n1088), .A3(n1087), .Y(n_src_aox[146])
         );
  AO222X1_HVT U1186 ( .A1(n1661), .A2(sram_rdata_8[19]), .A3(n2170), .A4(
        sram_rdata_7[19]), .A5(sram_rdata_6[19]), .A6(n1690), .Y(n1486) );
  AOI22X1_HVT U1187 ( .A1(n10901), .A2(n15000), .A3(n12400), .A4(n1486), .Y(
        n1093) );
  OA22X1_HVT U1188 ( .A1(n2780), .A2(n337), .A3(n14800), .A4(n528), .Y(n1092)
         );
  NAND2X0_HVT U1189 ( .A1(n1770), .A2(sram_rdata_3[19]), .Y(n1091) );
  NAND3X0_HVT U1190 ( .A1(n1093), .A2(n1092), .A3(n1091), .Y(n_src_aox[147])
         );
  AO222X1_HVT U1191 ( .A1(n2050), .A2(sram_rdata_8[20]), .A3(n2150), .A4(
        sram_rdata_7[20]), .A5(sram_rdata_6[20]), .A6(n1950), .Y(n1491) );
  AOI22X1_HVT U1192 ( .A1(n1094), .A2(n592), .A3(n11100), .A4(n1491), .Y(n1097) );
  OA22X1_HVT U1193 ( .A1(n2800), .A2(n338), .A3(n2740), .A4(n529), .Y(n1096)
         );
  NAND2X0_HVT U1194 ( .A1(n1760), .A2(sram_rdata_3[20]), .Y(n1095) );
  NAND3X0_HVT U1195 ( .A1(n1097), .A2(n1096), .A3(n1095), .Y(n_src_aox[148])
         );
  AO222X1_HVT U1196 ( .A1(n1860), .A2(sram_rdata_8[21]), .A3(n16601), .A4(
        sram_rdata_7[21]), .A5(sram_rdata_6[21]), .A6(n1980), .Y(n1493) );
  AOI22X1_HVT U1197 ( .A1(n1098), .A2(n591), .A3(n11000), .A4(n1493), .Y(n1101) );
  OA22X1_HVT U1198 ( .A1(n2790), .A2(n339), .A3(n2690), .A4(n5301), .Y(n11001)
         );
  NAND2X0_HVT U1199 ( .A1(n1730), .A2(sram_rdata_3[21]), .Y(n1099) );
  NAND3X0_HVT U1200 ( .A1(n1101), .A2(n11001), .A3(n1099), .Y(n_src_aox[149])
         );
  AO222X1_HVT U1201 ( .A1(n1820), .A2(sram_rdata_8[22]), .A3(n16000), .A4(
        sram_rdata_7[22]), .A5(sram_rdata_6[22]), .A6(n1900), .Y(n1498) );
  AOI22X1_HVT U1202 ( .A1(n1102), .A2(n594), .A3(n12400), .A4(n1498), .Y(n1105) );
  OA22X1_HVT U1203 ( .A1(n11800), .A2(n340), .A3(n14700), .A4(n531), .Y(n1104)
         );
  NAND2X0_HVT U1204 ( .A1(n574), .A2(sram_rdata_3[22]), .Y(n1103) );
  NAND3X0_HVT U1205 ( .A1(n1105), .A2(n1104), .A3(n1103), .Y(n_src_aox[150])
         );
  AO222X1_HVT U1206 ( .A1(n1880), .A2(sram_rdata_8[23]), .A3(n16200), .A4(
        sram_rdata_7[23]), .A5(sram_rdata_6[23]), .A6(n16600), .Y(n1503) );
  AOI22X1_HVT U1207 ( .A1(n1106), .A2(n10800), .A3(n583), .A4(n1503), .Y(n1109) );
  OA22X1_HVT U1208 ( .A1(n2760), .A2(n341), .A3(n2730), .A4(n532), .Y(n1108)
         );
  NAND2X0_HVT U1209 ( .A1(n1770), .A2(sram_rdata_3[23]), .Y(n1107) );
  NAND3X0_HVT U1210 ( .A1(n1109), .A2(n1108), .A3(n1107), .Y(n_src_aox[151])
         );
  AO222X1_HVT U1211 ( .A1(n1860), .A2(sram_rdata_8[24]), .A3(n2160), .A4(
        sram_rdata_7[24]), .A5(sram_rdata_6[24]), .A6(n2000), .Y(n1508) );
  AOI22X1_HVT U1212 ( .A1(n11101), .A2(n591), .A3(n12400), .A4(n1508), .Y(
        n1113) );
  OA22X1_HVT U1213 ( .A1(n2790), .A2(n342), .A3(n2730), .A4(n533), .Y(n1112)
         );
  NAND2X0_HVT U1214 ( .A1(n2270), .A2(sram_rdata_3[24]), .Y(n1111) );
  NAND3X0_HVT U1215 ( .A1(n1113), .A2(n1112), .A3(n1111), .Y(n_src_aox[152])
         );
  AO222X1_HVT U1216 ( .A1(n1840), .A2(sram_rdata_8[25]), .A3(n2180), .A4(
        sram_rdata_7[25]), .A5(sram_rdata_6[25]), .A6(n1960), .Y(n1513) );
  AOI22X1_HVT U1217 ( .A1(n1114), .A2(n15000), .A3(n12500), .A4(n1513), .Y(
        n1117) );
  OA22X1_HVT U1218 ( .A1(n2810), .A2(n343), .A3(n14700), .A4(n534), .Y(n1116)
         );
  NAND2X0_HVT U1219 ( .A1(n2220), .A2(sram_rdata_3[25]), .Y(n1115) );
  NAND3X0_HVT U1220 ( .A1(n1117), .A2(n1116), .A3(n1115), .Y(n_src_aox[153])
         );
  AO222X1_HVT U1221 ( .A1(n1860), .A2(sram_rdata_8[26]), .A3(n15500), .A4(
        sram_rdata_7[26]), .A5(sram_rdata_6[26]), .A6(n1930), .Y(n1518) );
  AOI22X1_HVT U1222 ( .A1(n1118), .A2(n12700), .A3(n11000), .A4(n1518), .Y(
        n1121) );
  OA22X1_HVT U1223 ( .A1(n2760), .A2(n344), .A3(n2690), .A4(n535), .Y(n11201)
         );
  NAND2X0_HVT U1224 ( .A1(n578), .A2(sram_rdata_3[26]), .Y(n1119) );
  NAND3X0_HVT U1225 ( .A1(n1121), .A2(n11201), .A3(n1119), .Y(n_src_aox[154])
         );
  AO222X1_HVT U1226 ( .A1(n2080), .A2(sram_rdata_8[27]), .A3(n15500), .A4(
        sram_rdata_7[27]), .A5(sram_rdata_6[27]), .A6(n1910), .Y(n1523) );
  AOI22X1_HVT U1227 ( .A1(n1122), .A2(n593), .A3(n582), .A4(n1523), .Y(n1125)
         );
  OA22X1_HVT U1228 ( .A1(n10200), .A2(n345), .A3(n14900), .A4(n536), .Y(n1124)
         );
  NAND2X0_HVT U1229 ( .A1(n2260), .A2(sram_rdata_3[27]), .Y(n1123) );
  NAND3X0_HVT U1230 ( .A1(n1125), .A2(n1124), .A3(n1123), .Y(n_src_aox[155])
         );
  AO222X1_HVT U1231 ( .A1(n2090), .A2(sram_rdata_8[28]), .A3(n2190), .A4(
        sram_rdata_7[28]), .A5(sram_rdata_6[28]), .A6(n16600), .Y(n1525) );
  AOI22X1_HVT U1232 ( .A1(n1126), .A2(n591), .A3(n12900), .A4(n1525), .Y(n1129) );
  OA22X1_HVT U1233 ( .A1(n11700), .A2(n3460), .A3(n10000), .A4(n537), .Y(n1128) );
  NAND2X0_HVT U1234 ( .A1(n1700), .A2(sram_rdata_3[28]), .Y(n1127) );
  NAND3X0_HVT U1235 ( .A1(n1129), .A2(n1128), .A3(n1127), .Y(n_src_aox[156])
         );
  AO222X1_HVT U1236 ( .A1(n2080), .A2(sram_rdata_8[29]), .A3(n15700), .A4(
        sram_rdata_7[29]), .A5(sram_rdata_6[29]), .A6(n1960), .Y(n15301) );
  AOI22X1_HVT U1237 ( .A1(n11301), .A2(n12800), .A3(n583), .A4(n15301), .Y(
        n1133) );
  OA22X1_HVT U1238 ( .A1(n11600), .A2(n347), .A3(n11400), .A4(n538), .Y(n1132)
         );
  NAND2X0_HVT U1239 ( .A1(n1730), .A2(sram_rdata_3[29]), .Y(n1131) );
  NAND3X0_HVT U1240 ( .A1(n1133), .A2(n1132), .A3(n1131), .Y(n_src_aox[157])
         );
  AO222X1_HVT U1241 ( .A1(n2080), .A2(sram_rdata_8[30]), .A3(n2200), .A4(
        sram_rdata_7[30]), .A5(sram_rdata_6[30]), .A6(n16600), .Y(n1532) );
  AOI22X1_HVT U1242 ( .A1(n1134), .A2(n12700), .A3(n11100), .A4(n1532), .Y(
        n1137) );
  OA22X1_HVT U1243 ( .A1(n2770), .A2(n348), .A3(n2710), .A4(n539), .Y(n1136)
         );
  NAND2X0_HVT U1244 ( .A1(n577), .A2(sram_rdata_3[30]), .Y(n1135) );
  NAND3X0_HVT U1245 ( .A1(n1137), .A2(n1136), .A3(n1135), .Y(n_src_aox[158])
         );
  AO222X1_HVT U1246 ( .A1(n1890), .A2(sram_rdata_8[31]), .A3(n2200), .A4(
        sram_rdata_7[31]), .A5(sram_rdata_6[31]), .A6(n16300), .Y(n1537) );
  AOI22X1_HVT U1247 ( .A1(n1138), .A2(n15100), .A3(n583), .A4(n1537), .Y(n1141) );
  OA22X1_HVT U1248 ( .A1(n13600), .A2(n349), .A3(n14800), .A4(n5401), .Y(
        n11401) );
  NAND2X0_HVT U1249 ( .A1(n2260), .A2(sram_rdata_3[31]), .Y(n1139) );
  NAND3X0_HVT U1250 ( .A1(n1141), .A2(n11401), .A3(n1139), .Y(n_src_aox[159])
         );
  AO222X1_HVT U1251 ( .A1(n2060), .A2(sram_rdata_7[16]), .A3(n2180), .A4(
        sram_rdata_6[16]), .A5(n16400), .A6(sram_rdata_8[16]), .Y(n1542) );
  AOI22X1_HVT U1252 ( .A1(n1142), .A2(n15000), .A3(n583), .A4(n1542), .Y(n1145) );
  OA22X1_HVT U1253 ( .A1(n10400), .A2(n429), .A3(n14900), .A4(n334), .Y(n1144)
         );
  NAND2X0_HVT U1254 ( .A1(n2210), .A2(sram_rdata_5[16]), .Y(n1143) );
  NAND3X0_HVT U1255 ( .A1(n1145), .A2(n1144), .A3(n1143), .Y(n_src_aox[160])
         );
  AO222X1_HVT U1256 ( .A1(n2040), .A2(sram_rdata_7[17]), .A3(n2170), .A4(
        sram_rdata_6[17]), .A5(n2010), .A6(sram_rdata_8[17]), .Y(n1544) );
  AOI22X1_HVT U1257 ( .A1(n1146), .A2(n12700), .A3(n581), .A4(n1544), .Y(n1149) );
  OA22X1_HVT U1258 ( .A1(n10300), .A2(n4301), .A3(n14600), .A4(n335), .Y(n1148) );
  NAND2X0_HVT U1259 ( .A1(n2210), .A2(sram_rdata_5[17]), .Y(n1147) );
  NAND3X0_HVT U1260 ( .A1(n1149), .A2(n1148), .A3(n1147), .Y(n_src_aox[161])
         );
  AO222X1_HVT U1261 ( .A1(n2090), .A2(sram_rdata_7[18]), .A3(n588), .A4(
        sram_rdata_6[18]), .A5(n1970), .A6(sram_rdata_8[18]), .Y(n1546) );
  AOI22X1_HVT U1262 ( .A1(n11501), .A2(n15100), .A3(n5801), .A4(n1546), .Y(
        n1153) );
  OA22X1_HVT U1263 ( .A1(n1663), .A2(n431), .A3(n11400), .A4(n336), .Y(n1152)
         );
  NAND2X0_HVT U1264 ( .A1(n1730), .A2(sram_rdata_5[18]), .Y(n1151) );
  NAND3X0_HVT U1265 ( .A1(n1153), .A2(n1152), .A3(n1151), .Y(n_src_aox[162])
         );
  AO222X1_HVT U1266 ( .A1(n1870), .A2(sram_rdata_7[19]), .A3(n2160), .A4(
        sram_rdata_6[19]), .A5(n1910), .A6(sram_rdata_8[19]), .Y(n1551) );
  AOI22X1_HVT U1267 ( .A1(n1154), .A2(n10800), .A3(n12500), .A4(n1551), .Y(
        n1157) );
  OA22X1_HVT U1268 ( .A1(n2770), .A2(n432), .A3(n14800), .A4(n337), .Y(n1156)
         );
  NAND2X0_HVT U1269 ( .A1(n2210), .A2(sram_rdata_5[19]), .Y(n1155) );
  NAND3X0_HVT U1270 ( .A1(n1157), .A2(n1156), .A3(n1155), .Y(n_src_aox[163])
         );
  AO222X1_HVT U1271 ( .A1(n1860), .A2(sram_rdata_7[20]), .A3(n2160), .A4(
        sram_rdata_6[20]), .A5(n1900), .A6(sram_rdata_8[20]), .Y(n1556) );
  AOI22X1_HVT U1272 ( .A1(n1158), .A2(n15000), .A3(n583), .A4(n1556), .Y(n1161) );
  OA22X1_HVT U1273 ( .A1(n2810), .A2(n433), .A3(n14800), .A4(n338), .Y(n11601)
         );
  NAND2X0_HVT U1274 ( .A1(n576), .A2(sram_rdata_5[20]), .Y(n1159) );
  NAND3X0_HVT U1275 ( .A1(n1161), .A2(n11601), .A3(n1159), .Y(n_src_aox[164])
         );
  AO222X1_HVT U1276 ( .A1(n1840), .A2(sram_rdata_7[21]), .A3(n2170), .A4(
        sram_rdata_6[21]), .A5(n1680), .A6(sram_rdata_8[21]), .Y(n1561) );
  AOI22X1_HVT U1277 ( .A1(n1162), .A2(n591), .A3(n11000), .A4(n1561), .Y(n1165) );
  OA22X1_HVT U1278 ( .A1(n2790), .A2(n434), .A3(n14700), .A4(n339), .Y(n1164)
         );
  NAND2X0_HVT U1279 ( .A1(n1780), .A2(sram_rdata_5[21]), .Y(n1163) );
  NAND3X0_HVT U1280 ( .A1(n1165), .A2(n1164), .A3(n1163), .Y(n_src_aox[165])
         );
  AO222X1_HVT U1281 ( .A1(n1810), .A2(sram_rdata_7[22]), .A3(n15400), .A4(
        sram_rdata_6[22]), .A5(n1680), .A6(sram_rdata_8[22]), .Y(n1563) );
  AOI22X1_HVT U1282 ( .A1(n1166), .A2(n12700), .A3(n11100), .A4(n1563), .Y(
        n1169) );
  OA22X1_HVT U1283 ( .A1(n10200), .A2(n435), .A3(n2700), .A4(n340), .Y(n1168)
         );
  NAND2X0_HVT U1284 ( .A1(n2250), .A2(sram_rdata_5[22]), .Y(n1167) );
  NAND3X0_HVT U1285 ( .A1(n1169), .A2(n1168), .A3(n1167), .Y(n_src_aox[166])
         );
  AO222X1_HVT U1286 ( .A1(n2070), .A2(sram_rdata_7[23]), .A3(n16000), .A4(
        sram_rdata_6[23]), .A5(n1670), .A6(sram_rdata_8[23]), .Y(n1565) );
  AOI22X1_HVT U1287 ( .A1(n11701), .A2(n15100), .A3(n582), .A4(n1565), .Y(
        n1173) );
  OA22X1_HVT U1288 ( .A1(n13700), .A2(n436), .A3(n10000), .A4(n341), .Y(n1172)
         );
  NAND2X0_HVT U1289 ( .A1(n1790), .A2(sram_rdata_5[23]), .Y(n1171) );
  NAND3X0_HVT U1290 ( .A1(n1173), .A2(n1172), .A3(n1171), .Y(n_src_aox[167])
         );
  AO222X1_HVT U1291 ( .A1(n2040), .A2(sram_rdata_7[24]), .A3(n2150), .A4(
        sram_rdata_6[24]), .A5(n16500), .A6(sram_rdata_8[24]), .Y(n15701) );
  AOI22X1_HVT U1292 ( .A1(n1174), .A2(n591), .A3(n12500), .A4(n15701), .Y(
        n1177) );
  OA22X1_HVT U1293 ( .A1(n13900), .A2(n437), .A3(n2730), .A4(n342), .Y(n1176)
         );
  NAND2X0_HVT U1294 ( .A1(n576), .A2(sram_rdata_5[24]), .Y(n1175) );
  NAND3X0_HVT U1295 ( .A1(n1177), .A2(n1176), .A3(n1175), .Y(n_src_aox[168])
         );
  AO222X1_HVT U1296 ( .A1(n2040), .A2(sram_rdata_7[25]), .A3(n588), .A4(
        sram_rdata_6[25]), .A5(n16400), .A6(sram_rdata_8[25]), .Y(n1572) );
  AOI22X1_HVT U1297 ( .A1(n1178), .A2(n12800), .A3(n11000), .A4(n1572), .Y(
        n1181) );
  OA22X1_HVT U1298 ( .A1(n2800), .A2(n438), .A3(n14600), .A4(n343), .Y(n11801)
         );
  NAND2X0_HVT U1299 ( .A1(n577), .A2(sram_rdata_5[25]), .Y(n1179) );
  NAND3X0_HVT U1300 ( .A1(n1181), .A2(n11801), .A3(n1179), .Y(n_src_aox[169])
         );
  AO222X1_HVT U1301 ( .A1(n2060), .A2(sram_rdata_7[26]), .A3(n16000), .A4(
        sram_rdata_6[26]), .A5(n16600), .A6(sram_rdata_8[26]), .Y(n1577) );
  AOI22X1_HVT U1302 ( .A1(n1182), .A2(n10900), .A3(n582), .A4(n1577), .Y(n1185) );
  OA22X1_HVT U1303 ( .A1(n2760), .A2(n439), .A3(n2690), .A4(n344), .Y(n1184)
         );
  NAND2X0_HVT U1304 ( .A1(n1740), .A2(sram_rdata_5[26]), .Y(n1183) );
  NAND3X0_HVT U1305 ( .A1(n1185), .A2(n1184), .A3(n1183), .Y(n_src_aox[170])
         );
  AO222X1_HVT U1306 ( .A1(n1840), .A2(sram_rdata_7[27]), .A3(n2190), .A4(
        sram_rdata_6[27]), .A5(n2020), .A6(sram_rdata_8[27]), .Y(n1579) );
  AOI22X1_HVT U1307 ( .A1(n1186), .A2(n593), .A3(n14400), .A4(n1579), .Y(n1189) );
  OA22X1_HVT U1308 ( .A1(n11800), .A2(n4401), .A3(n2720), .A4(n345), .Y(n1188)
         );
  NAND2X0_HVT U1309 ( .A1(n1800), .A2(sram_rdata_5[27]), .Y(n1187) );
  NAND3X0_HVT U1310 ( .A1(n1189), .A2(n1188), .A3(n1187), .Y(n_src_aox[171])
         );
  AO222X1_HVT U1311 ( .A1(n2040), .A2(sram_rdata_7[28]), .A3(n2160), .A4(
        sram_rdata_6[28]), .A5(n1980), .A6(sram_rdata_8[28]), .Y(n1581) );
  AOI22X1_HVT U1312 ( .A1(n11901), .A2(n591), .A3(n13000), .A4(n1581), .Y(
        n1193) );
  OA22X1_HVT U1313 ( .A1(n11700), .A2(n441), .A3(n2750), .A4(n3460), .Y(n1192)
         );
  NAND2X0_HVT U1314 ( .A1(n575), .A2(sram_rdata_5[28]), .Y(n1191) );
  NAND3X0_HVT U1315 ( .A1(n1193), .A2(n1192), .A3(n1191), .Y(n_src_aox[172])
         );
  AO222X1_HVT U1316 ( .A1(n1870), .A2(sram_rdata_7[29]), .A3(n2150), .A4(
        sram_rdata_6[29]), .A5(n2000), .A6(sram_rdata_8[29]), .Y(n1583) );
  AO222X1_HVT U1317 ( .A1(n1830), .A2(sram_rdata_7[30]), .A3(n2110), .A4(
        sram_rdata_6[30]), .A5(n1980), .A6(sram_rdata_8[30]), .Y(n1588) );
  AO222X1_HVT U1318 ( .A1(n1810), .A2(sram_rdata_7[31]), .A3(n15400), .A4(
        sram_rdata_6[31]), .A5(n1930), .A6(sram_rdata_8[31]), .Y(n1593) );
  AOI22X1_HVT U1319 ( .A1(n1196), .A2(n10800), .A3(n14400), .A4(n1593), .Y(
        n1199) );
  OA22X1_HVT U1320 ( .A1(n13600), .A2(n444), .A3(n14900), .A4(n349), .Y(n1198)
         );
  NAND2X0_HVT U1321 ( .A1(n574), .A2(sram_rdata_5[31]), .Y(n1197) );
  NAND3X0_HVT U1322 ( .A1(n1199), .A2(n1198), .A3(n1197), .Y(n_src_aox[175])
         );
  AO222X1_HVT U1323 ( .A1(n2070), .A2(sram_rdata_6[16]), .A3(n2150), .A4(
        sram_rdata_8[16]), .A5(sram_rdata_7[16]), .A6(n1980), .Y(n1598) );
  AOI22X1_HVT U1324 ( .A1(n12001), .A2(n591), .A3(n11100), .A4(n1598), .Y(
        n1203) );
  OA22X1_HVT U1325 ( .A1(n11600), .A2(n525), .A3(n2750), .A4(n429), .Y(n1202)
         );
  NAND2X0_HVT U1326 ( .A1(n1710), .A2(sram_rdata_4[16]), .Y(n1201) );
  NAND3X0_HVT U1327 ( .A1(n1203), .A2(n1202), .A3(n1201), .Y(n_src_aox[176])
         );
  AO222X1_HVT U1328 ( .A1(n12600), .A2(sram_rdata_6[17]), .A3(n16000), .A4(
        sram_rdata_8[17]), .A5(sram_rdata_7[17]), .A6(n1670), .Y(n1603) );
  AOI22X1_HVT U1329 ( .A1(n1204), .A2(n10900), .A3(n5801), .A4(n1603), .Y(
        n1207) );
  OA22X1_HVT U1330 ( .A1(n11700), .A2(n526), .A3(n10100), .A4(n4301), .Y(n1206) );
  NAND2X0_HVT U1331 ( .A1(n1780), .A2(sram_rdata_4[17]), .Y(n1205) );
  NAND3X0_HVT U1332 ( .A1(n1207), .A2(n1206), .A3(n1205), .Y(n_src_aox[177])
         );
  AO222X1_HVT U1333 ( .A1(n12600), .A2(sram_rdata_6[18]), .A3(n15600), .A4(
        sram_rdata_8[18]), .A5(sram_rdata_7[18]), .A6(n2000), .Y(n1608) );
  AOI22X1_HVT U1334 ( .A1(n1208), .A2(n15100), .A3(n5801), .A4(n1608), .Y(
        n1211) );
  OA22X1_HVT U1335 ( .A1(n1663), .A2(n527), .A3(n14700), .A4(n431), .Y(n12101)
         );
  NAND2X0_HVT U1336 ( .A1(n1800), .A2(sram_rdata_4[18]), .Y(n1209) );
  NAND3X0_HVT U1337 ( .A1(n1211), .A2(n12101), .A3(n1209), .Y(n_src_aox[178])
         );
  AO222X1_HVT U1338 ( .A1(n2100), .A2(sram_rdata_6[19]), .A3(n16200), .A4(
        sram_rdata_8[19]), .A5(sram_rdata_7[19]), .A6(n1960), .Y(n16101) );
  AOI22X1_HVT U1339 ( .A1(n1212), .A2(n15000), .A3(n14400), .A4(n16101), .Y(
        n1215) );
  OA22X1_HVT U1340 ( .A1(n2780), .A2(n528), .A3(n10000), .A4(n432), .Y(n1214)
         );
  NAND2X0_HVT U1341 ( .A1(n1760), .A2(sram_rdata_4[19]), .Y(n1213) );
  NAND3X0_HVT U1342 ( .A1(n1215), .A2(n1214), .A3(n1213), .Y(n_src_aox[179])
         );
  AO222X1_HVT U1343 ( .A1(n1860), .A2(sram_rdata_6[20]), .A3(n588), .A4(
        sram_rdata_8[20]), .A5(sram_rdata_7[20]), .A6(n2020), .Y(n1615) );
  AOI22X1_HVT U1344 ( .A1(n1216), .A2(n593), .A3(n10700), .A4(n1615), .Y(n1219) );
  OA22X1_HVT U1345 ( .A1(n2810), .A2(n529), .A3(n2730), .A4(n433), .Y(n1218)
         );
  NAND2X0_HVT U1346 ( .A1(n1730), .A2(sram_rdata_4[20]), .Y(n1217) );
  NAND3X0_HVT U1347 ( .A1(n1219), .A2(n1218), .A3(n1217), .Y(n_src_aox[180])
         );
  AO222X1_HVT U1348 ( .A1(n1810), .A2(sram_rdata_6[21]), .A3(n2110), .A4(
        sram_rdata_8[21]), .A5(sram_rdata_7[21]), .A6(n1950), .Y(n1617) );
  AOI22X1_HVT U1349 ( .A1(n12201), .A2(n12800), .A3(n582), .A4(n1617), .Y(
        n1223) );
  OA22X1_HVT U1350 ( .A1(n13900), .A2(n5301), .A3(n2690), .A4(n434), .Y(n1222)
         );
  NAND2X0_HVT U1351 ( .A1(n2270), .A2(sram_rdata_4[21]), .Y(n1221) );
  NAND3X0_HVT U1352 ( .A1(n1223), .A2(n1222), .A3(n1221), .Y(n_src_aox[181])
         );
  AO222X1_HVT U1353 ( .A1(n1830), .A2(sram_rdata_6[22]), .A3(n15900), .A4(
        sram_rdata_8[22]), .A5(sram_rdata_7[22]), .A6(n1900), .Y(n1622) );
  AOI22X1_HVT U1354 ( .A1(n1224), .A2(n15100), .A3(n5801), .A4(n1622), .Y(
        n1227) );
  OA22X1_HVT U1355 ( .A1(n10200), .A2(n531), .A3(n10100), .A4(n435), .Y(n1226)
         );
  NAND2X0_HVT U1356 ( .A1(n1730), .A2(sram_rdata_4[22]), .Y(n1225) );
  NAND3X0_HVT U1357 ( .A1(n1227), .A2(n1226), .A3(n1225), .Y(n_src_aox[182])
         );
  AO222X1_HVT U1358 ( .A1(n2060), .A2(sram_rdata_6[23]), .A3(n2180), .A4(
        sram_rdata_8[23]), .A5(sram_rdata_7[23]), .A6(n1680), .Y(n1627) );
  AOI22X1_HVT U1359 ( .A1(n1228), .A2(n591), .A3(n12500), .A4(n1627), .Y(n1231) );
  OA22X1_HVT U1360 ( .A1(n13600), .A2(n532), .A3(n14900), .A4(n436), .Y(n12301) );
  NAND2X0_HVT U1361 ( .A1(n1780), .A2(sram_rdata_4[23]), .Y(n1229) );
  NAND3X0_HVT U1362 ( .A1(n1231), .A2(n12301), .A3(n1229), .Y(n_src_aox[183])
         );
  AO222X1_HVT U1363 ( .A1(n2030), .A2(sram_rdata_6[24]), .A3(n15900), .A4(
        sram_rdata_8[24]), .A5(sram_rdata_7[24]), .A6(n1930), .Y(n1629) );
  AOI22X1_HVT U1364 ( .A1(n1232), .A2(n12700), .A3(n12900), .A4(n1629), .Y(
        n1235) );
  OA22X1_HVT U1365 ( .A1(n13800), .A2(n533), .A3(n14800), .A4(n437), .Y(n1234)
         );
  NAND2X0_HVT U1366 ( .A1(n576), .A2(sram_rdata_4[24]), .Y(n1233) );
  NAND3X0_HVT U1367 ( .A1(n1235), .A2(n1234), .A3(n1233), .Y(n_src_aox[184])
         );
  AO222X1_HVT U1368 ( .A1(n1820), .A2(sram_rdata_6[25]), .A3(n16100), .A4(
        sram_rdata_8[25]), .A5(sram_rdata_7[25]), .A6(n1680), .Y(n1631) );
  AOI22X1_HVT U1369 ( .A1(n1236), .A2(n1664), .A3(n10700), .A4(n1631), .Y(
        n1239) );
  OA22X1_HVT U1370 ( .A1(n13900), .A2(n534), .A3(n10000), .A4(n438), .Y(n1238)
         );
  NAND2X0_HVT U1371 ( .A1(n1790), .A2(sram_rdata_4[25]), .Y(n1237) );
  NAND3X0_HVT U1372 ( .A1(n1239), .A2(n1238), .A3(n1237), .Y(n_src_aox[185])
         );
  AO222X1_HVT U1373 ( .A1(n1890), .A2(sram_rdata_6[26]), .A3(n15500), .A4(
        sram_rdata_8[26]), .A5(sram_rdata_7[26]), .A6(n1980), .Y(n1636) );
  AO222X1_HVT U1374 ( .A1(n1830), .A2(sram_rdata_6[27]), .A3(n16100), .A4(
        sram_rdata_8[27]), .A5(sram_rdata_7[27]), .A6(n1690), .Y(n1641) );
  AO222X1_HVT U1375 ( .A1(n1890), .A2(sram_rdata_6[28]), .A3(n2140), .A4(
        sram_rdata_8[28]), .A5(sram_rdata_7[28]), .A6(n1970), .Y(n1643) );
  AO222X1_HVT U1376 ( .A1(n2070), .A2(sram_rdata_6[29]), .A3(n2150), .A4(
        sram_rdata_8[29]), .A5(sram_rdata_7[29]), .A6(n16400), .Y(n1645) );
  AOI22X1_HVT U1377 ( .A1(n1243), .A2(n15100), .A3(n582), .A4(n1645), .Y(n1246) );
  OA22X1_HVT U1378 ( .A1(n10400), .A2(n538), .A3(n2700), .A4(n442), .Y(n1245)
         );
  NAND2X0_HVT U1379 ( .A1(n574), .A2(sram_rdata_4[29]), .Y(n1244) );
  NAND3X0_HVT U1380 ( .A1(n1246), .A2(n1245), .A3(n1244), .Y(n_src_aox[189])
         );
  AO222X1_HVT U1381 ( .A1(n1890), .A2(sram_rdata_6[30]), .A3(n15900), .A4(
        sram_rdata_8[30]), .A5(sram_rdata_7[30]), .A6(n1670), .Y(n16501) );
  AOI22X1_HVT U1382 ( .A1(n1247), .A2(n15000), .A3(n5801), .A4(n16501), .Y(
        n12501) );
  OA22X1_HVT U1383 ( .A1(n2770), .A2(n539), .A3(n10100), .A4(n443), .Y(n1249)
         );
  NAND2X0_HVT U1384 ( .A1(n1710), .A2(sram_rdata_4[30]), .Y(n1248) );
  NAND3X0_HVT U1385 ( .A1(n12501), .A2(n1249), .A3(n1248), .Y(n_src_aox[190])
         );
  AO222X1_HVT U1386 ( .A1(n2090), .A2(sram_rdata_6[31]), .A3(n2110), .A4(
        sram_rdata_8[31]), .A5(sram_rdata_7[31]), .A6(n1970), .Y(n1652) );
  AOI22X1_HVT U1387 ( .A1(n1251), .A2(n591), .A3(n12500), .A4(n1652), .Y(n1254) );
  OA22X1_HVT U1388 ( .A1(n2770), .A2(n5401), .A3(n2730), .A4(n444), .Y(n1253)
         );
  NAND2X0_HVT U1389 ( .A1(n2240), .A2(sram_rdata_4[31]), .Y(n1252) );
  NAND3X0_HVT U1390 ( .A1(n1254), .A2(n1253), .A3(n1252), .Y(n_src_aox[191])
         );
  AOI22X1_HVT U1391 ( .A1(n1258), .A2(n583), .A3(n5901), .A4(n1257), .Y(n1261)
         );
  OA22X1_HVT U1392 ( .A1(n11700), .A2(n351), .A3(n2700), .A4(n542), .Y(n12601)
         );
  NAND2X0_HVT U1393 ( .A1(n1770), .A2(sram_rdata_0[1]), .Y(n1259) );
  NAND3X0_HVT U1394 ( .A1(n1261), .A2(n12601), .A3(n1259), .Y(n_src_aox[193])
         );
  AOI22X1_HVT U1395 ( .A1(n1265), .A2(n10700), .A3(n5901), .A4(n1264), .Y(
        n1268) );
  OA22X1_HVT U1396 ( .A1(n2770), .A2(n353), .A3(n2720), .A4(n544), .Y(n1267)
         );
  NAND2X0_HVT U1397 ( .A1(n2260), .A2(sram_rdata_0[3]), .Y(n1266) );
  NAND3X0_HVT U1398 ( .A1(n1268), .A2(n1267), .A3(n1266), .Y(n_src_aox[195])
         );
  AOI22X1_HVT U1399 ( .A1(n12701), .A2(n13000), .A3(n12700), .A4(n1269), .Y(
        n1273) );
  OA22X1_HVT U1400 ( .A1(n2800), .A2(n354), .A3(n1662), .A4(n545), .Y(n1272)
         );
  NAND2X0_HVT U1401 ( .A1(n2220), .A2(sram_rdata_0[4]), .Y(n1271) );
  NAND3X0_HVT U1402 ( .A1(n1273), .A2(n1272), .A3(n1271), .Y(n_src_aox[196])
         );
  AOI22X1_HVT U1403 ( .A1(n1275), .A2(n11100), .A3(n594), .A4(n1274), .Y(n1278) );
  OA22X1_HVT U1404 ( .A1(n2790), .A2(n355), .A3(n11400), .A4(n546), .Y(n1277)
         );
  NAND2X0_HVT U1405 ( .A1(n2210), .A2(sram_rdata_0[5]), .Y(n1276) );
  NAND3X0_HVT U1406 ( .A1(n1278), .A2(n1277), .A3(n1276), .Y(n_src_aox[197])
         );
  AOI22X1_HVT U1407 ( .A1(n12801), .A2(n14400), .A3(n5901), .A4(n1279), .Y(
        n1283) );
  OA22X1_HVT U1408 ( .A1(n11800), .A2(n356), .A3(n14600), .A4(n547), .Y(n1282)
         );
  NAND2X0_HVT U1409 ( .A1(n1760), .A2(sram_rdata_0[6]), .Y(n1281) );
  NAND3X0_HVT U1410 ( .A1(n1283), .A2(n1282), .A3(n1281), .Y(n_src_aox[198])
         );
  AOI22X1_HVT U1411 ( .A1(n1285), .A2(n11000), .A3(n594), .A4(n1284), .Y(n1288) );
  OA22X1_HVT U1412 ( .A1(n13600), .A2(n357), .A3(n2740), .A4(n548), .Y(n1287)
         );
  NAND2X0_HVT U1413 ( .A1(n574), .A2(sram_rdata_0[7]), .Y(n1286) );
  NAND3X0_HVT U1414 ( .A1(n1288), .A2(n1287), .A3(n1286), .Y(n_src_aox[199])
         );
  AOI22X1_HVT U1415 ( .A1(n12901), .A2(n13000), .A3(n10800), .A4(n1289), .Y(
        n1293) );
  OA22X1_HVT U1416 ( .A1(n13900), .A2(n358), .A3(n2750), .A4(n549), .Y(n1292)
         );
  NAND2X0_HVT U1417 ( .A1(n2220), .A2(sram_rdata_0[8]), .Y(n1291) );
  NAND3X0_HVT U1418 ( .A1(n1293), .A2(n1292), .A3(n1291), .Y(n_src_aox[200])
         );
  AOI22X1_HVT U1419 ( .A1(n1295), .A2(n12500), .A3(n12700), .A4(n1294), .Y(
        n1298) );
  OA22X1_HVT U1420 ( .A1(n2810), .A2(n359), .A3(n11400), .A4(n5501), .Y(n1297)
         );
  NAND2X0_HVT U1421 ( .A1(n1770), .A2(sram_rdata_0[9]), .Y(n1296) );
  NAND3X0_HVT U1422 ( .A1(n1298), .A2(n1297), .A3(n1296), .Y(n_src_aox[201])
         );
  AOI22X1_HVT U1423 ( .A1(n13001), .A2(n581), .A3(n592), .A4(n1299), .Y(n1303)
         );
  OA22X1_HVT U1424 ( .A1(n13700), .A2(n360), .A3(n10100), .A4(n551), .Y(n1302)
         );
  NAND2X0_HVT U1425 ( .A1(n2250), .A2(sram_rdata_0[10]), .Y(n1301) );
  NAND3X0_HVT U1426 ( .A1(n1303), .A2(n1302), .A3(n1301), .Y(n_src_aox[202])
         );
  AOI22X1_HVT U1427 ( .A1(n1305), .A2(n581), .A3(n594), .A4(n1304), .Y(n1308)
         );
  OA22X1_HVT U1428 ( .A1(n10200), .A2(n361), .A3(n2740), .A4(n552), .Y(n1307)
         );
  NAND2X0_HVT U1429 ( .A1(n1750), .A2(sram_rdata_0[11]), .Y(n1306) );
  NAND3X0_HVT U1430 ( .A1(n1308), .A2(n1307), .A3(n1306), .Y(n_src_aox[203])
         );
  AOI22X1_HVT U1431 ( .A1(n13101), .A2(n12500), .A3(n592), .A4(n1309), .Y(
        n1313) );
  OA22X1_HVT U1432 ( .A1(n10300), .A2(n362), .A3(n2740), .A4(n553), .Y(n1312)
         );
  NAND2X0_HVT U1433 ( .A1(n2210), .A2(sram_rdata_0[12]), .Y(n1311) );
  NAND3X0_HVT U1434 ( .A1(n1313), .A2(n1312), .A3(n1311), .Y(n_src_aox[204])
         );
  AOI22X1_HVT U1435 ( .A1(n1315), .A2(n12900), .A3(n5901), .A4(n1314), .Y(
        n1318) );
  OA22X1_HVT U1436 ( .A1(n11600), .A2(n363), .A3(n2710), .A4(n554), .Y(n1317)
         );
  NAND2X0_HVT U1437 ( .A1(n1700), .A2(sram_rdata_0[13]), .Y(n1316) );
  NAND3X0_HVT U1438 ( .A1(n1318), .A2(n1317), .A3(n1316), .Y(n_src_aox[205])
         );
  AOI22X1_HVT U1439 ( .A1(n13201), .A2(n12500), .A3(n10800), .A4(n1319), .Y(
        n1323) );
  OA22X1_HVT U1440 ( .A1(n13600), .A2(n364), .A3(n2750), .A4(n555), .Y(n1322)
         );
  NAND2X0_HVT U1441 ( .A1(n1770), .A2(sram_rdata_0[14]), .Y(n1321) );
  NAND3X0_HVT U1442 ( .A1(n1323), .A2(n1322), .A3(n1321), .Y(n_src_aox[206])
         );
  AOI22X1_HVT U1443 ( .A1(n1325), .A2(n11100), .A3(n594), .A4(n1324), .Y(n1328) );
  OA22X1_HVT U1444 ( .A1(n1663), .A2(n365), .A3(n10000), .A4(n556), .Y(n1327)
         );
  NAND2X0_HVT U1445 ( .A1(n576), .A2(sram_rdata_0[15]), .Y(n1326) );
  NAND3X0_HVT U1446 ( .A1(n1328), .A2(n1327), .A3(n1326), .Y(n_src_aox[207])
         );
  AOI22X1_HVT U1447 ( .A1(n13301), .A2(n12800), .A3(n582), .A4(n1329), .Y(
        n1333) );
  OA22X1_HVT U1448 ( .A1(n10400), .A2(n445), .A3(n2720), .A4(n350), .Y(n1332)
         );
  NAND2X0_HVT U1449 ( .A1(n1710), .A2(sram_rdata_2[0]), .Y(n1331) );
  NAND3X0_HVT U1450 ( .A1(n1333), .A2(n1332), .A3(n1331), .Y(n_src_aox[208])
         );
  AOI22X1_HVT U1451 ( .A1(n1335), .A2(n12500), .A3(n592), .A4(n1334), .Y(n1338) );
  OA22X1_HVT U1452 ( .A1(n10300), .A2(n446), .A3(n2690), .A4(n351), .Y(n1337)
         );
  NAND2X0_HVT U1453 ( .A1(n1710), .A2(sram_rdata_2[1]), .Y(n1336) );
  NAND3X0_HVT U1454 ( .A1(n1338), .A2(n1337), .A3(n1336), .Y(n_src_aox[209])
         );
  AOI22X1_HVT U1455 ( .A1(n13401), .A2(n581), .A3(n592), .A4(n1339), .Y(n1343)
         );
  OA22X1_HVT U1456 ( .A1(n13900), .A2(n447), .A3(n2690), .A4(n352), .Y(n1342)
         );
  NAND2X0_HVT U1457 ( .A1(n2240), .A2(sram_rdata_2[2]), .Y(n1341) );
  NAND3X0_HVT U1458 ( .A1(n1343), .A2(n1342), .A3(n1341), .Y(n_src_aox[210])
         );
  AOI22X1_HVT U1459 ( .A1(n1345), .A2(n581), .A3(n592), .A4(n1344), .Y(n1348)
         );
  OA22X1_HVT U1460 ( .A1(n2770), .A2(n448), .A3(n2720), .A4(n353), .Y(n1347)
         );
  NAND2X0_HVT U1461 ( .A1(n1790), .A2(sram_rdata_2[3]), .Y(n1346) );
  NAND3X0_HVT U1462 ( .A1(n1348), .A2(n1347), .A3(n1346), .Y(n_src_aox[211])
         );
  AOI22X1_HVT U1463 ( .A1(n13501), .A2(n12400), .A3(n5901), .A4(n1349), .Y(
        n1353) );
  OA22X1_HVT U1464 ( .A1(n2810), .A2(n449), .A3(n14900), .A4(n354), .Y(n1352)
         );
  NAND2X0_HVT U1465 ( .A1(n577), .A2(sram_rdata_2[4]), .Y(n1351) );
  NAND3X0_HVT U1466 ( .A1(n1353), .A2(n1352), .A3(n1351), .Y(n_src_aox[212])
         );
  AOI22X1_HVT U1467 ( .A1(n1357), .A2(n13000), .A3(n5901), .A4(n1356), .Y(
        n13601) );
  OA22X1_HVT U1468 ( .A1(n10200), .A2(n451), .A3(n2710), .A4(n356), .Y(n1359)
         );
  NAND2X0_HVT U1469 ( .A1(n1750), .A2(sram_rdata_2[6]), .Y(n1358) );
  NAND3X0_HVT U1470 ( .A1(n13601), .A2(n1359), .A3(n1358), .Y(n_src_aox[214])
         );
  AOI22X1_HVT U1471 ( .A1(n1362), .A2(n12400), .A3(n594), .A4(n1361), .Y(n1365) );
  OA22X1_HVT U1472 ( .A1(n2760), .A2(n452), .A3(n14800), .A4(n357), .Y(n1364)
         );
  NAND2X0_HVT U1473 ( .A1(n1750), .A2(sram_rdata_2[7]), .Y(n1363) );
  NAND3X0_HVT U1474 ( .A1(n1365), .A2(n1364), .A3(n1363), .Y(n_src_aox[215])
         );
  AOI22X1_HVT U1475 ( .A1(n1367), .A2(n12900), .A3(n592), .A4(n1366), .Y(
        n13701) );
  OA22X1_HVT U1476 ( .A1(n2790), .A2(n453), .A3(n2720), .A4(n358), .Y(n1369)
         );
  NAND2X0_HVT U1477 ( .A1(n1750), .A2(sram_rdata_2[8]), .Y(n1368) );
  NAND3X0_HVT U1478 ( .A1(n13701), .A2(n1369), .A3(n1368), .Y(n_src_aox[216])
         );
  AOI22X1_HVT U1479 ( .A1(n1372), .A2(n14400), .A3(n5901), .A4(n1371), .Y(
        n1375) );
  OA22X1_HVT U1480 ( .A1(n2800), .A2(n454), .A3(n14700), .A4(n359), .Y(n1374)
         );
  NAND2X0_HVT U1481 ( .A1(n2270), .A2(sram_rdata_2[9]), .Y(n1373) );
  NAND3X0_HVT U1482 ( .A1(n1375), .A2(n1374), .A3(n1373), .Y(n_src_aox[217])
         );
  AOI22X1_HVT U1483 ( .A1(n1377), .A2(n13000), .A3(n5901), .A4(n1376), .Y(
        n13801) );
  OA22X1_HVT U1484 ( .A1(n2760), .A2(n455), .A3(n14700), .A4(n360), .Y(n1379)
         );
  NAND2X0_HVT U1485 ( .A1(n576), .A2(sram_rdata_2[10]), .Y(n1378) );
  NAND3X0_HVT U1486 ( .A1(n13801), .A2(n1379), .A3(n1378), .Y(n_src_aox[218])
         );
  AOI22X1_HVT U1487 ( .A1(n1382), .A2(n11000), .A3(n12800), .A4(n1381), .Y(
        n1385) );
  OA22X1_HVT U1488 ( .A1(n11800), .A2(n456), .A3(n2730), .A4(n361), .Y(n1384)
         );
  NAND2X0_HVT U1489 ( .A1(n1790), .A2(sram_rdata_2[11]), .Y(n1383) );
  NAND3X0_HVT U1490 ( .A1(n1385), .A2(n1384), .A3(n1383), .Y(n_src_aox[219])
         );
  AOI22X1_HVT U1491 ( .A1(n1387), .A2(n11000), .A3(n592), .A4(n1386), .Y(
        n13901) );
  OA22X1_HVT U1492 ( .A1(n11700), .A2(n457), .A3(n10000), .A4(n362), .Y(n1389)
         );
  NAND2X0_HVT U1493 ( .A1(n1760), .A2(sram_rdata_2[12]), .Y(n1388) );
  NAND3X0_HVT U1494 ( .A1(n13901), .A2(n1389), .A3(n1388), .Y(n_src_aox[220])
         );
  AOI22X1_HVT U1495 ( .A1(n1392), .A2(n581), .A3(n5901), .A4(n1391), .Y(n1395)
         );
  OA22X1_HVT U1496 ( .A1(n10400), .A2(n458), .A3(n10100), .A4(n363), .Y(n1394)
         );
  NAND2X0_HVT U1497 ( .A1(n1750), .A2(sram_rdata_2[13]), .Y(n1393) );
  NAND3X0_HVT U1498 ( .A1(n1395), .A2(n1394), .A3(n1393), .Y(n_src_aox[221])
         );
  AOI22X1_HVT U1499 ( .A1(n1399), .A2(n14400), .A3(n12700), .A4(n1398), .Y(
        n1402) );
  OA22X1_HVT U1500 ( .A1(n13900), .A2(n4601), .A3(n14800), .A4(n365), .Y(n1401) );
  NAND2X0_HVT U1501 ( .A1(n1700), .A2(sram_rdata_2[15]), .Y(n14001) );
  NAND3X0_HVT U1502 ( .A1(n1402), .A2(n1401), .A3(n14001), .Y(n_src_aox[223])
         );
  AOI22X1_HVT U1503 ( .A1(n1406), .A2(n12900), .A3(n5901), .A4(n1405), .Y(
        n1409) );
  OA22X1_HVT U1504 ( .A1(n11700), .A2(n542), .A3(n14600), .A4(n446), .Y(n1408)
         );
  NAND2X0_HVT U1505 ( .A1(n578), .A2(sram_rdata_1[1]), .Y(n1407) );
  NAND3X0_HVT U1506 ( .A1(n1409), .A2(n1408), .A3(n1407), .Y(n_src_aox[225])
         );
  AOI22X1_HVT U1507 ( .A1(n1411), .A2(n14400), .A3(n10800), .A4(n14101), .Y(
        n1414) );
  OA22X1_HVT U1508 ( .A1(n13600), .A2(n543), .A3(n11400), .A4(n447), .Y(n1413)
         );
  NAND2X0_HVT U1509 ( .A1(n578), .A2(sram_rdata_1[2]), .Y(n1412) );
  NAND3X0_HVT U1510 ( .A1(n1414), .A2(n1413), .A3(n1412), .Y(n_src_aox[226])
         );
  AOI22X1_HVT U1511 ( .A1(n1418), .A2(n13000), .A3(n592), .A4(n1417), .Y(n1421) );
  OA22X1_HVT U1512 ( .A1(n2800), .A2(n545), .A3(n2740), .A4(n449), .Y(n14201)
         );
  NAND2X0_HVT U1513 ( .A1(n577), .A2(sram_rdata_1[4]), .Y(n1419) );
  NAND3X0_HVT U1514 ( .A1(n1421), .A2(n14201), .A3(n1419), .Y(n_src_aox[228])
         );
  AOI22X1_HVT U1515 ( .A1(n1423), .A2(n13000), .A3(n592), .A4(n1422), .Y(n1426) );
  OA22X1_HVT U1516 ( .A1(n13900), .A2(n546), .A3(n2710), .A4(n4501), .Y(n1425)
         );
  NAND2X0_HVT U1517 ( .A1(n1790), .A2(sram_rdata_1[5]), .Y(n1424) );
  NAND3X0_HVT U1518 ( .A1(n1426), .A2(n1425), .A3(n1424), .Y(n_src_aox[229])
         );
  AOI22X1_HVT U1519 ( .A1(n14301), .A2(n581), .A3(n592), .A4(n1429), .Y(n1433)
         );
  OA22X1_HVT U1520 ( .A1(n13600), .A2(n548), .A3(n10000), .A4(n452), .Y(n1432)
         );
  NAND2X0_HVT U1521 ( .A1(n2260), .A2(sram_rdata_1[7]), .Y(n1431) );
  NAND3X0_HVT U1522 ( .A1(n1433), .A2(n1432), .A3(n1431), .Y(n_src_aox[231])
         );
  AOI22X1_HVT U1523 ( .A1(n1435), .A2(n10700), .A3(n12800), .A4(n1434), .Y(
        n1438) );
  OA22X1_HVT U1524 ( .A1(n13900), .A2(n549), .A3(n14900), .A4(n453), .Y(n1437)
         );
  NAND2X0_HVT U1525 ( .A1(n1730), .A2(sram_rdata_1[8]), .Y(n1436) );
  NAND3X0_HVT U1526 ( .A1(n1438), .A2(n1437), .A3(n1436), .Y(n_src_aox[232])
         );
  AOI22X1_HVT U1527 ( .A1(n14401), .A2(n10700), .A3(n594), .A4(n1439), .Y(
        n1443) );
  OA22X1_HVT U1528 ( .A1(n2810), .A2(n5501), .A3(n2710), .A4(n454), .Y(n1442)
         );
  NAND2X0_HVT U1529 ( .A1(n576), .A2(sram_rdata_1[9]), .Y(n1441) );
  NAND3X0_HVT U1530 ( .A1(n1443), .A2(n1442), .A3(n1441), .Y(n_src_aox[233])
         );
  AOI22X1_HVT U1531 ( .A1(n1445), .A2(n13000), .A3(n10900), .A4(n1444), .Y(
        n1448) );
  OA22X1_HVT U1532 ( .A1(n2760), .A2(n551), .A3(n14700), .A4(n455), .Y(n1447)
         );
  NAND2X0_HVT U1533 ( .A1(n1750), .A2(sram_rdata_1[10]), .Y(n1446) );
  NAND3X0_HVT U1534 ( .A1(n1448), .A2(n1447), .A3(n1446), .Y(n_src_aox[234])
         );
  AOI22X1_HVT U1535 ( .A1(n14501), .A2(n11100), .A3(n594), .A4(n1449), .Y(
        n1453) );
  OA22X1_HVT U1536 ( .A1(n10200), .A2(n552), .A3(n2720), .A4(n456), .Y(n1452)
         );
  NAND2X0_HVT U1537 ( .A1(n576), .A2(sram_rdata_1[11]), .Y(n1451) );
  NAND3X0_HVT U1538 ( .A1(n1453), .A2(n1452), .A3(n1451), .Y(n_src_aox[235])
         );
  AOI22X1_HVT U1539 ( .A1(n1455), .A2(n581), .A3(n592), .A4(n1454), .Y(n1458)
         );
  OA22X1_HVT U1540 ( .A1(n10300), .A2(n553), .A3(n2730), .A4(n457), .Y(n1457)
         );
  NAND2X0_HVT U1541 ( .A1(n577), .A2(sram_rdata_1[12]), .Y(n1456) );
  NAND3X0_HVT U1542 ( .A1(n1458), .A2(n1457), .A3(n1456), .Y(n_src_aox[236])
         );
  AOI22X1_HVT U1543 ( .A1(n14601), .A2(n12500), .A3(n5901), .A4(n1459), .Y(
        n1463) );
  OA22X1_HVT U1544 ( .A1(n11600), .A2(n554), .A3(n2690), .A4(n458), .Y(n1462)
         );
  NAND2X0_HVT U1545 ( .A1(n1780), .A2(sram_rdata_1[13]), .Y(n1461) );
  NAND3X0_HVT U1546 ( .A1(n1463), .A2(n1462), .A3(n1461), .Y(n_src_aox[237])
         );
  AOI22X1_HVT U1547 ( .A1(n1467), .A2(n14400), .A3(n5901), .A4(n1466), .Y(
        n14701) );
  OA22X1_HVT U1548 ( .A1(n13800), .A2(n556), .A3(n14800), .A4(n4601), .Y(n1469) );
  NAND2X0_HVT U1549 ( .A1(n1800), .A2(sram_rdata_1[15]), .Y(n1468) );
  NAND3X0_HVT U1550 ( .A1(n14701), .A2(n1469), .A3(n1468), .Y(n_src_aox[239])
         );
  AOI22X1_HVT U1551 ( .A1(n1472), .A2(n12400), .A3(n5901), .A4(n1471), .Y(
        n1475) );
  OA22X1_HVT U1552 ( .A1(n11600), .A2(n366), .A3(n10000), .A4(n557), .Y(n1474)
         );
  NAND2X0_HVT U1553 ( .A1(n575), .A2(sram_rdata_0[16]), .Y(n1473) );
  NAND3X0_HVT U1554 ( .A1(n1475), .A2(n1474), .A3(n1473), .Y(n_src_aox[240])
         );
  AOI22X1_HVT U1555 ( .A1(n1477), .A2(n581), .A3(n594), .A4(n1476), .Y(n14801)
         );
  OA22X1_HVT U1556 ( .A1(n10300), .A2(n367), .A3(n10100), .A4(n558), .Y(n1479)
         );
  NAND2X0_HVT U1557 ( .A1(n575), .A2(sram_rdata_0[17]), .Y(n1478) );
  NAND3X0_HVT U1558 ( .A1(n14801), .A2(n1479), .A3(n1478), .Y(n_src_aox[241])
         );
  AOI22X1_HVT U1559 ( .A1(n1482), .A2(n11000), .A3(n594), .A4(n1481), .Y(n1485) );
  OA22X1_HVT U1560 ( .A1(n13700), .A2(n368), .A3(n14600), .A4(n559), .Y(n1484)
         );
  NAND2X0_HVT U1561 ( .A1(n1750), .A2(sram_rdata_0[18]), .Y(n1483) );
  NAND3X0_HVT U1562 ( .A1(n1485), .A2(n1484), .A3(n1483), .Y(n_src_aox[242])
         );
  AOI22X1_HVT U1563 ( .A1(n1487), .A2(n12900), .A3(n594), .A4(n1486), .Y(
        n14901) );
  OA22X1_HVT U1564 ( .A1(n2770), .A2(n369), .A3(n1662), .A4(n5601), .Y(n1489)
         );
  NAND2X0_HVT U1565 ( .A1(n574), .A2(sram_rdata_0[19]), .Y(n1488) );
  NAND3X0_HVT U1566 ( .A1(n14901), .A2(n1489), .A3(n1488), .Y(n_src_aox[243])
         );
  AOI22X1_HVT U1567 ( .A1(n1494), .A2(n11100), .A3(n592), .A4(n1493), .Y(n1497) );
  OA22X1_HVT U1568 ( .A1(n13800), .A2(n371), .A3(n2700), .A4(n562), .Y(n1496)
         );
  NAND2X0_HVT U1569 ( .A1(n577), .A2(sram_rdata_0[21]), .Y(n1495) );
  NAND3X0_HVT U1570 ( .A1(n1497), .A2(n1496), .A3(n1495), .Y(n_src_aox[245])
         );
  AOI22X1_HVT U1571 ( .A1(n1499), .A2(n581), .A3(n594), .A4(n1498), .Y(n1502)
         );
  OA22X1_HVT U1572 ( .A1(n11800), .A2(n372), .A3(n10100), .A4(n563), .Y(n1501)
         );
  NAND2X0_HVT U1573 ( .A1(n2240), .A2(sram_rdata_0[22]), .Y(n15001) );
  NAND3X0_HVT U1574 ( .A1(n1502), .A2(n1501), .A3(n15001), .Y(n_src_aox[246])
         );
  AOI22X1_HVT U1575 ( .A1(n1504), .A2(n12500), .A3(n5901), .A4(n1503), .Y(
        n1507) );
  OA22X1_HVT U1576 ( .A1(n2760), .A2(n373), .A3(n2740), .A4(n564), .Y(n1506)
         );
  NAND2X0_HVT U1577 ( .A1(n1800), .A2(sram_rdata_0[23]), .Y(n1505) );
  NAND3X0_HVT U1578 ( .A1(n1507), .A2(n1506), .A3(n1505), .Y(n_src_aox[247])
         );
  AOI22X1_HVT U1579 ( .A1(n1509), .A2(n11000), .A3(n5901), .A4(n1508), .Y(
        n1512) );
  OA22X1_HVT U1580 ( .A1(n13900), .A2(n374), .A3(n14800), .A4(n565), .Y(n1511)
         );
  NAND2X0_HVT U1581 ( .A1(n578), .A2(sram_rdata_0[24]), .Y(n15101) );
  NAND3X0_HVT U1582 ( .A1(n1512), .A2(n1511), .A3(n15101), .Y(n_src_aox[248])
         );
  AOI22X1_HVT U1583 ( .A1(n1514), .A2(n581), .A3(n5901), .A4(n1513), .Y(n1517)
         );
  OA22X1_HVT U1584 ( .A1(n2810), .A2(n375), .A3(n2700), .A4(n566), .Y(n1516)
         );
  NAND2X0_HVT U1585 ( .A1(n2220), .A2(sram_rdata_0[25]), .Y(n1515) );
  NAND3X0_HVT U1586 ( .A1(n1517), .A2(n1516), .A3(n1515), .Y(n_src_aox[249])
         );
  AOI22X1_HVT U1587 ( .A1(n1519), .A2(n12400), .A3(n12800), .A4(n1518), .Y(
        n1522) );
  OA22X1_HVT U1588 ( .A1(n2760), .A2(n376), .A3(n14600), .A4(n567), .Y(n1521)
         );
  NAND2X0_HVT U1589 ( .A1(n1770), .A2(sram_rdata_0[26]), .Y(n15201) );
  NAND3X0_HVT U1590 ( .A1(n1522), .A2(n1521), .A3(n15201), .Y(n_src_aox[250])
         );
  AOI22X1_HVT U1591 ( .A1(n1526), .A2(n581), .A3(n594), .A4(n1525), .Y(n1529)
         );
  OA22X1_HVT U1592 ( .A1(n10300), .A2(n378), .A3(n14800), .A4(n569), .Y(n1528)
         );
  NAND2X0_HVT U1593 ( .A1(n1750), .A2(sram_rdata_0[28]), .Y(n1527) );
  NAND3X0_HVT U1594 ( .A1(n1529), .A2(n1528), .A3(n1527), .Y(n_src_aox[252])
         );
  AOI22X1_HVT U1595 ( .A1(n1533), .A2(n11000), .A3(n5901), .A4(n1532), .Y(
        n1536) );
  OA22X1_HVT U1596 ( .A1(n2780), .A2(n380), .A3(n11400), .A4(n571), .Y(n1535)
         );
  NAND2X0_HVT U1597 ( .A1(n1770), .A2(sram_rdata_0[30]), .Y(n1534) );
  NAND3X0_HVT U1598 ( .A1(n1536), .A2(n1535), .A3(n1534), .Y(n_src_aox[254])
         );
  AOI22X1_HVT U1599 ( .A1(n1538), .A2(n583), .A3(n592), .A4(n1537), .Y(n1541)
         );
  OA22X1_HVT U1600 ( .A1(n2770), .A2(n381), .A3(n2730), .A4(n572), .Y(n15401)
         );
  NAND2X0_HVT U1601 ( .A1(n1770), .A2(sram_rdata_0[31]), .Y(n1539) );
  NAND3X0_HVT U1602 ( .A1(n1541), .A2(n15401), .A3(n1539), .Y(n_src_aox[255])
         );
  AOI22X1_HVT U1603 ( .A1(n1547), .A2(n13000), .A3(n5901), .A4(n1546), .Y(
        n15501) );
  OA22X1_HVT U1604 ( .A1(n13600), .A2(n463), .A3(n14600), .A4(n368), .Y(n1549)
         );
  NAND2X0_HVT U1605 ( .A1(n2250), .A2(sram_rdata_2[18]), .Y(n1548) );
  NAND3X0_HVT U1606 ( .A1(n15501), .A2(n1549), .A3(n1548), .Y(n_src_aox[258])
         );
  AOI22X1_HVT U1607 ( .A1(n1552), .A2(n12500), .A3(n594), .A4(n1551), .Y(n1555) );
  OA22X1_HVT U1608 ( .A1(n2780), .A2(n464), .A3(n2730), .A4(n369), .Y(n1554)
         );
  NAND2X0_HVT U1609 ( .A1(n574), .A2(sram_rdata_2[19]), .Y(n1553) );
  NAND3X0_HVT U1610 ( .A1(n1555), .A2(n1554), .A3(n1553), .Y(n_src_aox[259])
         );
  AOI22X1_HVT U1611 ( .A1(n1557), .A2(n581), .A3(n594), .A4(n1556), .Y(n15601)
         );
  OA22X1_HVT U1612 ( .A1(n2810), .A2(n465), .A3(n1662), .A4(n370), .Y(n1559)
         );
  NAND2X0_HVT U1613 ( .A1(n2250), .A2(sram_rdata_2[20]), .Y(n1558) );
  NAND3X0_HVT U1614 ( .A1(n15601), .A2(n1559), .A3(n1558), .Y(n_src_aox[260])
         );
  AOI22X1_HVT U1615 ( .A1(n1566), .A2(n12900), .A3(n592), .A4(n1565), .Y(n1569) );
  OA22X1_HVT U1616 ( .A1(n13600), .A2(n468), .A3(n2740), .A4(n373), .Y(n1568)
         );
  NAND2X0_HVT U1617 ( .A1(n2240), .A2(sram_rdata_2[23]), .Y(n1567) );
  NAND3X0_HVT U1618 ( .A1(n1569), .A2(n1568), .A3(n1567), .Y(n_src_aox[263])
         );
  AOI22X1_HVT U1619 ( .A1(n1573), .A2(n12400), .A3(n592), .A4(n1572), .Y(n1576) );
  OA22X1_HVT U1620 ( .A1(n2800), .A2(n4701), .A3(n11400), .A4(n375), .Y(n1575)
         );
  NAND2X0_HVT U1621 ( .A1(n1800), .A2(sram_rdata_2[25]), .Y(n1574) );
  NAND3X0_HVT U1622 ( .A1(n1576), .A2(n1575), .A3(n1574), .Y(n_src_aox[265])
         );
  AOI22X1_HVT U1623 ( .A1(n1584), .A2(n10700), .A3(n594), .A4(n1583), .Y(n1587) );
  OA22X1_HVT U1624 ( .A1(n11600), .A2(n474), .A3(n2690), .A4(n379), .Y(n1586)
         );
  NAND2X0_HVT U1625 ( .A1(n574), .A2(sram_rdata_2[29]), .Y(n1585) );
  NAND3X0_HVT U1626 ( .A1(n1587), .A2(n1586), .A3(n1585), .Y(n_src_aox[269])
         );
  AOI22X1_HVT U1627 ( .A1(n1589), .A2(n583), .A3(n592), .A4(n1588), .Y(n1592)
         );
  OA22X1_HVT U1628 ( .A1(n13700), .A2(n475), .A3(n11400), .A4(n380), .Y(n1591)
         );
  NAND2X0_HVT U1629 ( .A1(n1740), .A2(sram_rdata_2[30]), .Y(n15901) );
  NAND3X0_HVT U1630 ( .A1(n1592), .A2(n1591), .A3(n15901), .Y(n_src_aox[270])
         );
  AOI22X1_HVT U1631 ( .A1(n1594), .A2(n11100), .A3(n592), .A4(n1593), .Y(n1597) );
  OA22X1_HVT U1632 ( .A1(n13800), .A2(n476), .A3(n10000), .A4(n381), .Y(n1596)
         );
  NAND2X0_HVT U1633 ( .A1(n1760), .A2(sram_rdata_2[31]), .Y(n1595) );
  NAND3X0_HVT U1634 ( .A1(n1597), .A2(n1596), .A3(n1595), .Y(n_src_aox[271])
         );
  AOI22X1_HVT U1635 ( .A1(n1599), .A2(n10700), .A3(n592), .A4(n1598), .Y(n1602) );
  OA22X1_HVT U1636 ( .A1(n11600), .A2(n557), .A3(n14800), .A4(n461), .Y(n1601)
         );
  NAND2X0_HVT U1637 ( .A1(n574), .A2(sram_rdata_1[16]), .Y(n16001) );
  NAND3X0_HVT U1638 ( .A1(n1602), .A2(n1601), .A3(n16001), .Y(n_src_aox[272])
         );
  AOI22X1_HVT U1639 ( .A1(n1604), .A2(n581), .A3(n592), .A4(n1603), .Y(n1607)
         );
  OA22X1_HVT U1640 ( .A1(n11700), .A2(n558), .A3(n14700), .A4(n462), .Y(n1606)
         );
  NAND2X0_HVT U1641 ( .A1(n1800), .A2(sram_rdata_1[17]), .Y(n1605) );
  NAND3X0_HVT U1642 ( .A1(n1607), .A2(n1606), .A3(n1605), .Y(n_src_aox[273])
         );
  AOI22X1_HVT U1643 ( .A1(n1611), .A2(n12500), .A3(n5901), .A4(n16101), .Y(
        n1614) );
  OA22X1_HVT U1644 ( .A1(n2780), .A2(n5601), .A3(n14900), .A4(n464), .Y(n1613)
         );
  NAND2X0_HVT U1645 ( .A1(n1740), .A2(sram_rdata_1[19]), .Y(n1612) );
  NAND3X0_HVT U1646 ( .A1(n1614), .A2(n1613), .A3(n1612), .Y(n_src_aox[275])
         );
  AOI22X1_HVT U1647 ( .A1(n1618), .A2(n581), .A3(n594), .A4(n1617), .Y(n1621)
         );
  OA22X1_HVT U1648 ( .A1(n2790), .A2(n562), .A3(n14700), .A4(n466), .Y(n16201)
         );
  NAND2X0_HVT U1649 ( .A1(n2210), .A2(sram_rdata_1[21]), .Y(n1619) );
  NAND3X0_HVT U1650 ( .A1(n1621), .A2(n16201), .A3(n1619), .Y(n_src_aox[277])
         );
  AOI22X1_HVT U1651 ( .A1(n1623), .A2(n12400), .A3(n594), .A4(n1622), .Y(n1626) );
  OA22X1_HVT U1652 ( .A1(n11800), .A2(n563), .A3(n2710), .A4(n467), .Y(n1625)
         );
  NAND2X0_HVT U1653 ( .A1(n1790), .A2(sram_rdata_1[22]), .Y(n1624) );
  NAND3X0_HVT U1654 ( .A1(n1626), .A2(n1625), .A3(n1624), .Y(n_src_aox[278])
         );
  AOI22X1_HVT U1655 ( .A1(n1632), .A2(n12900), .A3(n5901), .A4(n1631), .Y(
        n1635) );
  OA22X1_HVT U1656 ( .A1(n2810), .A2(n566), .A3(n2710), .A4(n4701), .Y(n1634)
         );
  NAND2X0_HVT U1657 ( .A1(n578), .A2(sram_rdata_1[25]), .Y(n1633) );
  NAND3X0_HVT U1658 ( .A1(n1635), .A2(n1634), .A3(n1633), .Y(n_src_aox[281])
         );
  AOI22X1_HVT U1659 ( .A1(n1637), .A2(n10700), .A3(n5901), .A4(n1636), .Y(
        n16401) );
  OA22X1_HVT U1660 ( .A1(n13700), .A2(n567), .A3(n2710), .A4(n471), .Y(n1639)
         );
  NAND2X0_HVT U1661 ( .A1(n2240), .A2(sram_rdata_1[26]), .Y(n1638) );
  NAND3X0_HVT U1662 ( .A1(n16401), .A2(n1639), .A3(n1638), .Y(n_src_aox[282])
         );
  AOI22X1_HVT U1663 ( .A1(n1646), .A2(n12400), .A3(n592), .A4(n1645), .Y(n1649) );
  OA22X1_HVT U1664 ( .A1(n10400), .A2(n5701), .A3(n10100), .A4(n474), .Y(n1648) );
  NAND2X0_HVT U1665 ( .A1(n2210), .A2(sram_rdata_1[29]), .Y(n1647) );
  NAND3X0_HVT U1666 ( .A1(n1649), .A2(n1648), .A3(n1647), .Y(n_src_aox[285])
         );
  AND2X1_HVT U1667 ( .A1(box_sel[1]), .A2(box_sel[0]), .Y(n16601) );
  AND2X1_HVT U1668 ( .A1(box_sel[0]), .A2(n1658), .Y(n1661) );
  AND2X1_HVT U1669 ( .A1(box_sel[3]), .A2(n1657), .Y(n1664) );
  AO22X1_HVT U1670 ( .A1(n2670), .A2(sram_rdata_b1[29]), .A3(n2330), .A4(
        sram_rdata_a1[29]), .Y(N100) );
  AO22X1_HVT U1671 ( .A1(n14200), .A2(sram_rdata_b1[30]), .A3(n2640), .A4(
        sram_rdata_a1[30]), .Y(N101) );
  AO22X1_HVT U1672 ( .A1(n2620), .A2(sram_rdata_b1[31]), .A3(n2290), .A4(
        sram_rdata_a1[31]), .Y(N102) );
  AO22X1_HVT U1673 ( .A1(n11900), .A2(sram_rdata_b2[0]), .A3(n2290), .A4(
        sram_rdata_a2[0]), .Y(N103) );
  AO22X1_HVT U1674 ( .A1(n2660), .A2(sram_rdata_b2[1]), .A3(n2360), .A4(
        sram_rdata_a2[1]), .Y(N104) );
  AO22X1_HVT U1675 ( .A1(n14300), .A2(sram_rdata_b2[2]), .A3(n2290), .A4(
        sram_rdata_a2[2]), .Y(N105) );
  AO22X1_HVT U1676 ( .A1(n1667), .A2(sram_rdata_b2[3]), .A3(n2330), .A4(
        sram_rdata_a2[3]), .Y(N106) );
  AO22X1_HVT U1677 ( .A1(n2610), .A2(sram_rdata_b2[4]), .A3(n2330), .A4(
        sram_rdata_a2[4]), .Y(N107) );
  AO22X1_HVT U1678 ( .A1(n14200), .A2(sram_rdata_b2[5]), .A3(n2300), .A4(
        sram_rdata_a2[5]), .Y(N108) );
  AO22X1_HVT U1679 ( .A1(n10500), .A2(sram_rdata_b2[6]), .A3(n2340), .A4(
        sram_rdata_a2[6]), .Y(N109) );
  AO22X1_HVT U1680 ( .A1(n10600), .A2(sram_rdata_b2[7]), .A3(n2360), .A4(
        sram_rdata_a2[7]), .Y(N110) );
  AO22X1_HVT U1681 ( .A1(n2670), .A2(sram_rdata_b2[8]), .A3(n2350), .A4(
        sram_rdata_a2[8]), .Y(N111) );
  AO22X1_HVT U1682 ( .A1(n2650), .A2(sram_rdata_b2[9]), .A3(n2330), .A4(
        sram_rdata_a2[9]), .Y(N112) );
  AO22X1_HVT U1683 ( .A1(n2650), .A2(sram_rdata_b2[10]), .A3(n2350), .A4(
        sram_rdata_a2[10]), .Y(N113) );
  AO22X1_HVT U1684 ( .A1(n2600), .A2(sram_rdata_b2[11]), .A3(n2310), .A4(
        sram_rdata_a2[11]), .Y(N114) );
  AO22X1_HVT U1685 ( .A1(n2600), .A2(sram_rdata_b2[12]), .A3(n2310), .A4(
        sram_rdata_a2[12]), .Y(N115) );
  AO22X1_HVT U1686 ( .A1(n10500), .A2(sram_rdata_b2[13]), .A3(n2820), .A4(
        sram_rdata_a2[13]), .Y(N116) );
  AO22X1_HVT U1687 ( .A1(n14300), .A2(sram_rdata_b2[14]), .A3(n2300), .A4(
        sram_rdata_a2[14]), .Y(N117) );
  AO22X1_HVT U1688 ( .A1(n1667), .A2(sram_rdata_b2[15]), .A3(n2820), .A4(
        sram_rdata_a2[15]), .Y(N118) );
  AO22X1_HVT U1689 ( .A1(n10600), .A2(sram_rdata_b2[16]), .A3(n14100), .A4(
        sram_rdata_a2[16]), .Y(N119) );
  AO22X1_HVT U1690 ( .A1(n2680), .A2(sram_rdata_b2[17]), .A3(n2290), .A4(
        sram_rdata_a2[17]), .Y(N120) );
  AO22X1_HVT U1691 ( .A1(n2680), .A2(sram_rdata_b2[18]), .A3(n2310), .A4(
        sram_rdata_a2[18]), .Y(N121) );
  AO22X1_HVT U1692 ( .A1(n2630), .A2(sram_rdata_b2[19]), .A3(n2360), .A4(
        sram_rdata_a2[19]), .Y(N122) );
  AO22X1_HVT U1693 ( .A1(n2630), .A2(sram_rdata_b2[20]), .A3(n2340), .A4(
        sram_rdata_a2[20]), .Y(N123) );
  AO22X1_HVT U1694 ( .A1(n2650), .A2(sram_rdata_b2[21]), .A3(n2820), .A4(
        sram_rdata_a2[21]), .Y(N124) );
  AO22X1_HVT U1695 ( .A1(n14300), .A2(sram_rdata_b2[22]), .A3(n2320), .A4(
        sram_rdata_a2[22]), .Y(N125) );
  AO22X1_HVT U1696 ( .A1(n11900), .A2(sram_rdata_b2[23]), .A3(n2350), .A4(
        sram_rdata_a2[23]), .Y(N126) );
  AO22X1_HVT U1697 ( .A1(n2600), .A2(sram_rdata_b2[24]), .A3(n595), .A4(
        sram_rdata_a2[24]), .Y(N127) );
  AO22X1_HVT U1698 ( .A1(n2660), .A2(sram_rdata_b2[25]), .A3(n2360), .A4(
        sram_rdata_a2[25]), .Y(N128) );
  AO22X1_HVT U1699 ( .A1(n14200), .A2(sram_rdata_b2[26]), .A3(n2280), .A4(
        sram_rdata_a2[26]), .Y(N129) );
  AO22X1_HVT U1700 ( .A1(n2670), .A2(sram_rdata_b2[27]), .A3(n2280), .A4(
        sram_rdata_a2[27]), .Y(N130) );
  AO22X1_HVT U1701 ( .A1(n2610), .A2(sram_rdata_b2[28]), .A3(n2280), .A4(
        sram_rdata_a2[28]), .Y(N131) );
  AO22X1_HVT U1702 ( .A1(n14200), .A2(sram_rdata_b2[29]), .A3(n2320), .A4(
        sram_rdata_a2[29]), .Y(N132) );
  AO22X1_HVT U1703 ( .A1(n2680), .A2(sram_rdata_b2[30]), .A3(n2290), .A4(
        sram_rdata_a2[30]), .Y(N133) );
  AO22X1_HVT U1704 ( .A1(n2630), .A2(sram_rdata_b2[31]), .A3(n2340), .A4(
        sram_rdata_a2[31]), .Y(N134) );
  AO22X1_HVT U1705 ( .A1(n11900), .A2(sram_rdata_b3[0]), .A3(n2360), .A4(
        sram_rdata_a3[0]), .Y(N135) );
  AO22X1_HVT U1706 ( .A1(n14300), .A2(sram_rdata_b3[1]), .A3(n2280), .A4(
        sram_rdata_a3[1]), .Y(N136) );
  AO22X1_HVT U1707 ( .A1(n2660), .A2(sram_rdata_b3[2]), .A3(n2310), .A4(
        sram_rdata_a3[2]), .Y(N137) );
  AO22X1_HVT U1708 ( .A1(n2610), .A2(sram_rdata_b3[3]), .A3(n2300), .A4(
        sram_rdata_a3[3]), .Y(N138) );
  AO22X1_HVT U1709 ( .A1(n10500), .A2(sram_rdata_b3[4]), .A3(n2340), .A4(
        sram_rdata_a3[4]), .Y(N139) );
  AO22X1_HVT U1710 ( .A1(n2660), .A2(sram_rdata_b3[5]), .A3(n2330), .A4(
        sram_rdata_a3[5]), .Y(N140) );
  AO22X1_HVT U1711 ( .A1(n10500), .A2(sram_rdata_b3[6]), .A3(n2330), .A4(
        sram_rdata_a3[6]), .Y(N141) );
  AO22X1_HVT U1712 ( .A1(n10600), .A2(sram_rdata_b3[7]), .A3(n2360), .A4(
        sram_rdata_a3[7]), .Y(N142) );
  AO22X1_HVT U1713 ( .A1(n2610), .A2(sram_rdata_b3[8]), .A3(n2820), .A4(
        sram_rdata_a3[8]), .Y(N143) );
  AO22X1_HVT U1714 ( .A1(n2680), .A2(sram_rdata_b3[9]), .A3(n2350), .A4(
        sram_rdata_a3[9]), .Y(N144) );
  AO22X1_HVT U1715 ( .A1(n14300), .A2(sram_rdata_b3[10]), .A3(n2820), .A4(
        sram_rdata_a3[10]), .Y(N145) );
  AO22X1_HVT U1716 ( .A1(n2620), .A2(sram_rdata_b3[11]), .A3(n2290), .A4(
        sram_rdata_a3[11]), .Y(N146) );
  AO22X1_HVT U1717 ( .A1(n2630), .A2(sram_rdata_b3[12]), .A3(n2290), .A4(
        sram_rdata_a3[12]), .Y(N147) );
  AO22X1_HVT U1718 ( .A1(n10500), .A2(sram_rdata_b3[13]), .A3(n2350), .A4(
        sram_rdata_a3[13]), .Y(N148) );
  AO22X1_HVT U1719 ( .A1(n2660), .A2(sram_rdata_b3[14]), .A3(n2350), .A4(
        sram_rdata_a3[14]), .Y(N149) );
  AO22X1_HVT U1720 ( .A1(n2610), .A2(sram_rdata_b3[15]), .A3(n2820), .A4(
        sram_rdata_a3[15]), .Y(N150) );
  AO22X1_HVT U1721 ( .A1(n10600), .A2(sram_rdata_b3[16]), .A3(n2300), .A4(
        sram_rdata_a3[16]), .Y(N151) );
  AO22X1_HVT U1722 ( .A1(n14200), .A2(sram_rdata_b3[17]), .A3(n2280), .A4(
        sram_rdata_a3[17]), .Y(N152) );
  AO22X1_HVT U1723 ( .A1(n2650), .A2(sram_rdata_b3[18]), .A3(n1666), .A4(
        sram_rdata_a3[18]), .Y(N153) );
  AO22X1_HVT U1724 ( .A1(n2600), .A2(sram_rdata_b3[19]), .A3(n2320), .A4(
        sram_rdata_a3[19]), .Y(N154) );
  AO22X1_HVT U1725 ( .A1(n2620), .A2(sram_rdata_b3[20]), .A3(n2320), .A4(
        sram_rdata_a3[20]), .Y(N155) );
  AO22X1_HVT U1726 ( .A1(n2680), .A2(sram_rdata_b3[21]), .A3(n2310), .A4(
        sram_rdata_a3[21]), .Y(N156) );
  AO22X1_HVT U1727 ( .A1(n2670), .A2(sram_rdata_b3[22]), .A3(n2290), .A4(
        sram_rdata_a3[22]), .Y(N157) );
  AO22X1_HVT U1728 ( .A1(n11900), .A2(sram_rdata_b3[23]), .A3(n2290), .A4(
        sram_rdata_a3[23]), .Y(N158) );
  AO22X1_HVT U1729 ( .A1(n2630), .A2(sram_rdata_b3[24]), .A3(n2340), .A4(
        sram_rdata_a3[24]), .Y(N159) );
  AO22X1_HVT U1730 ( .A1(n14300), .A2(sram_rdata_b3[25]), .A3(n2340), .A4(
        sram_rdata_a3[25]), .Y(N160) );
  AO22X1_HVT U1731 ( .A1(n2680), .A2(sram_rdata_b3[26]), .A3(n2330), .A4(
        sram_rdata_a3[26]), .Y(N161) );
  AO22X1_HVT U1732 ( .A1(n2630), .A2(sram_rdata_b3[27]), .A3(n2360), .A4(
        sram_rdata_a3[27]), .Y(N162) );
  AO22X1_HVT U1733 ( .A1(n2620), .A2(sram_rdata_b3[28]), .A3(n2360), .A4(
        sram_rdata_a3[28]), .Y(N163) );
  AO22X1_HVT U1734 ( .A1(n2670), .A2(sram_rdata_b3[29]), .A3(n2360), .A4(
        sram_rdata_a3[29]), .Y(N164) );
  AO22X1_HVT U1735 ( .A1(n2650), .A2(sram_rdata_b3[30]), .A3(n2280), .A4(
        sram_rdata_a3[30]), .Y(N165) );
  AO22X1_HVT U1736 ( .A1(n2600), .A2(sram_rdata_b3[31]), .A3(n2310), .A4(
        sram_rdata_a3[31]), .Y(N166) );
  AO22X1_HVT U1737 ( .A1(n11900), .A2(sram_rdata_b4[0]), .A3(n2300), .A4(
        sram_rdata_a4[0]), .Y(N167) );
  AO22X1_HVT U1738 ( .A1(n2650), .A2(sram_rdata_b4[1]), .A3(n2320), .A4(
        sram_rdata_a4[1]), .Y(N168) );
  AO22X1_HVT U1739 ( .A1(n2680), .A2(sram_rdata_b4[2]), .A3(n2360), .A4(
        sram_rdata_a4[2]), .Y(N169) );
  AO22X1_HVT U1740 ( .A1(n2630), .A2(sram_rdata_b4[3]), .A3(n2330), .A4(
        sram_rdata_a4[3]), .Y(N170) );
  AO22X1_HVT U1741 ( .A1(n2600), .A2(sram_rdata_b4[4]), .A3(n2310), .A4(
        sram_rdata_a4[4]), .Y(N171) );
  AO22X1_HVT U1742 ( .A1(n14300), .A2(sram_rdata_b4[5]), .A3(n2300), .A4(
        sram_rdata_a4[5]), .Y(N172) );
  AO22X1_HVT U1743 ( .A1(n10500), .A2(sram_rdata_b4[6]), .A3(n2290), .A4(
        sram_rdata_a4[6]), .Y(N173) );
  AO22X1_HVT U1744 ( .A1(n10600), .A2(sram_rdata_b4[7]), .A3(n2290), .A4(
        sram_rdata_a4[7]), .Y(N174) );
  AO22X1_HVT U1745 ( .A1(n1667), .A2(sram_rdata_b4[8]), .A3(n2330), .A4(
        sram_rdata_a4[8]), .Y(N175) );
  AO22X1_HVT U1746 ( .A1(n14200), .A2(sram_rdata_b4[9]), .A3(n595), .A4(
        sram_rdata_a4[9]), .Y(N176) );
  AO22X1_HVT U1747 ( .A1(n2660), .A2(sram_rdata_b4[10]), .A3(n2330), .A4(
        sram_rdata_a4[10]), .Y(N177) );
  AO22X1_HVT U1748 ( .A1(n2610), .A2(sram_rdata_b4[11]), .A3(n595), .A4(
        sram_rdata_a4[11]), .Y(N178) );
  AO22X1_HVT U1749 ( .A1(n1667), .A2(sram_rdata_b4[12]), .A3(n2640), .A4(
        sram_rdata_a4[12]), .Y(N179) );
  AO22X1_HVT U1750 ( .A1(n10500), .A2(sram_rdata_b4[13]), .A3(n2350), .A4(
        sram_rdata_a4[13]), .Y(N180) );
  AO22X1_HVT U1751 ( .A1(n14200), .A2(sram_rdata_b4[14]), .A3(n2340), .A4(
        sram_rdata_a4[14]), .Y(N181) );
  AO22X1_HVT U1752 ( .A1(n2670), .A2(sram_rdata_b4[15]), .A3(n2310), .A4(
        sram_rdata_a4[15]), .Y(N182) );
  AO22X1_HVT U1753 ( .A1(n10600), .A2(sram_rdata_b4[16]), .A3(n2300), .A4(
        sram_rdata_a4[16]), .Y(N183) );
  AO22X1_HVT U1754 ( .A1(n2660), .A2(sram_rdata_b4[17]), .A3(n2350), .A4(
        sram_rdata_a4[17]), .Y(N184) );
  AO22X1_HVT U1755 ( .A1(n2660), .A2(sram_rdata_b4[18]), .A3(n2820), .A4(
        sram_rdata_a4[18]), .Y(N185) );
  AO22X1_HVT U1756 ( .A1(n2610), .A2(sram_rdata_b4[19]), .A3(n2330), .A4(
        sram_rdata_a4[19]), .Y(N186) );
  AO22X1_HVT U1757 ( .A1(n2610), .A2(sram_rdata_b4[20]), .A3(n2280), .A4(
        sram_rdata_a4[20]), .Y(N187) );
  AO22X1_HVT U1758 ( .A1(n14200), .A2(sram_rdata_b4[21]), .A3(n2300), .A4(
        sram_rdata_a4[21]), .Y(N188) );
  AO22X1_HVT U1759 ( .A1(n2650), .A2(sram_rdata_b4[22]), .A3(n2360), .A4(
        sram_rdata_a4[22]), .Y(N189) );
  AO22X1_HVT U1760 ( .A1(n11900), .A2(sram_rdata_b4[23]), .A3(n14100), .A4(
        sram_rdata_a4[23]), .Y(N190) );
  AO22X1_HVT U1761 ( .A1(n2620), .A2(sram_rdata_b4[24]), .A3(n2820), .A4(
        sram_rdata_a4[24]), .Y(N191) );
  AO22X1_HVT U1762 ( .A1(n2650), .A2(sram_rdata_b4[25]), .A3(n2300), .A4(
        sram_rdata_a4[25]), .Y(N192) );
  AO22X1_HVT U1763 ( .A1(n2650), .A2(sram_rdata_b4[26]), .A3(n2300), .A4(
        sram_rdata_a4[26]), .Y(N193) );
  AO22X1_HVT U1764 ( .A1(n2600), .A2(sram_rdata_b4[27]), .A3(n2350), .A4(
        sram_rdata_a4[27]), .Y(N194) );
  AO22X1_HVT U1765 ( .A1(n2600), .A2(sram_rdata_b4[28]), .A3(n2820), .A4(
        sram_rdata_a4[28]), .Y(N195) );
  AO22X1_HVT U1766 ( .A1(n2650), .A2(sram_rdata_b4[29]), .A3(n2320), .A4(
        sram_rdata_a4[29]), .Y(N196) );
  AO22X1_HVT U1767 ( .A1(n14300), .A2(sram_rdata_b4[30]), .A3(n14100), .A4(
        sram_rdata_a4[30]), .Y(N197) );
  AO22X1_HVT U1768 ( .A1(n1667), .A2(sram_rdata_b4[31]), .A3(n1666), .A4(
        sram_rdata_a4[31]), .Y(N198) );
  AO22X1_HVT U1769 ( .A1(n11900), .A2(sram_rdata_b5[0]), .A3(n2350), .A4(
        sram_rdata_a5[0]), .Y(N199) );
  AO22X1_HVT U1770 ( .A1(n2680), .A2(sram_rdata_b5[1]), .A3(n14100), .A4(
        sram_rdata_a5[1]), .Y(N200) );
  AO22X1_HVT U1771 ( .A1(n2650), .A2(sram_rdata_b5[2]), .A3(n2310), .A4(
        sram_rdata_a5[2]), .Y(N201) );
  AO22X1_HVT U1772 ( .A1(n2600), .A2(sram_rdata_b5[3]), .A3(n2290), .A4(
        sram_rdata_a5[3]), .Y(N202) );
  AO22X1_HVT U1773 ( .A1(n2630), .A2(sram_rdata_b5[4]), .A3(n2280), .A4(
        sram_rdata_a5[4]), .Y(N203) );
  AO22X1_HVT U1774 ( .A1(n2650), .A2(sram_rdata_b5[5]), .A3(n2820), .A4(
        sram_rdata_a5[5]), .Y(N204) );
  AO22X1_HVT U1775 ( .A1(n10500), .A2(sram_rdata_b5[6]), .A3(n1666), .A4(
        sram_rdata_a5[6]), .Y(N205) );
  AO22X1_HVT U1776 ( .A1(n10600), .A2(sram_rdata_b5[7]), .A3(n2340), .A4(
        sram_rdata_a5[7]), .Y(N206) );
  AO22X1_HVT U1777 ( .A1(n2600), .A2(sram_rdata_b5[8]), .A3(n595), .A4(
        sram_rdata_a5[8]), .Y(N207) );
  AO22X1_HVT U1778 ( .A1(n2660), .A2(sram_rdata_b5[9]), .A3(n2310), .A4(
        sram_rdata_a5[9]), .Y(N208) );
  AO22X1_HVT U1779 ( .A1(n14200), .A2(sram_rdata_b5[10]), .A3(n2280), .A4(
        sram_rdata_a5[10]), .Y(N209) );
  AO22X1_HVT U1780 ( .A1(n2620), .A2(sram_rdata_b5[11]), .A3(n2310), .A4(
        sram_rdata_a5[11]), .Y(N210) );
  AO22X1_HVT U1781 ( .A1(n2610), .A2(sram_rdata_b5[12]), .A3(n2330), .A4(
        sram_rdata_a5[12]), .Y(N211) );
  AO22X1_HVT U1782 ( .A1(n10500), .A2(sram_rdata_b5[13]), .A3(n2340), .A4(
        sram_rdata_a5[13]), .Y(N212) );
  AO22X1_HVT U1783 ( .A1(n2680), .A2(sram_rdata_b5[14]), .A3(n2340), .A4(
        sram_rdata_a5[14]), .Y(N213) );
  AO22X1_HVT U1784 ( .A1(n2630), .A2(sram_rdata_b5[15]), .A3(n2360), .A4(
        sram_rdata_a5[15]), .Y(N214) );
  AO22X1_HVT U1785 ( .A1(n10600), .A2(sram_rdata_b5[16]), .A3(n2350), .A4(
        sram_rdata_a5[16]), .Y(N215) );
  AO22X1_HVT U1786 ( .A1(n14300), .A2(sram_rdata_b5[17]), .A3(n2350), .A4(
        sram_rdata_a5[17]), .Y(N216) );
  AO22X1_HVT U1787 ( .A1(n14200), .A2(sram_rdata_b5[18]), .A3(n2330), .A4(
        sram_rdata_a5[18]), .Y(N217) );
  AO22X1_HVT U1788 ( .A1(n2620), .A2(sram_rdata_b5[19]), .A3(n2290), .A4(
        sram_rdata_a5[19]), .Y(N218) );
  AO22X1_HVT U1789 ( .A1(n10500), .A2(sram_rdata_b5[20]), .A3(n2280), .A4(
        sram_rdata_a5[20]), .Y(N219) );
  AO22X1_HVT U1790 ( .A1(n2660), .A2(sram_rdata_b5[21]), .A3(n2350), .A4(
        sram_rdata_a5[21]), .Y(N220) );
  AO22X1_HVT U1791 ( .A1(n2670), .A2(sram_rdata_b5[22]), .A3(n2350), .A4(
        sram_rdata_a5[22]), .Y(N221) );
  AO22X1_HVT U1792 ( .A1(n11900), .A2(sram_rdata_b5[23]), .A3(n2320), .A4(
        sram_rdata_a5[23]), .Y(N222) );
  AO22X1_HVT U1793 ( .A1(n2610), .A2(sram_rdata_b5[24]), .A3(n2300), .A4(
        sram_rdata_a5[24]), .Y(N223) );
  AO22X1_HVT U1794 ( .A1(n2680), .A2(sram_rdata_b5[25]), .A3(n2290), .A4(
        sram_rdata_a5[25]), .Y(N224) );
  AO22X1_HVT U1795 ( .A1(n14300), .A2(sram_rdata_b5[26]), .A3(n595), .A4(
        sram_rdata_a5[26]), .Y(N225) );
  AO22X1_HVT U1796 ( .A1(n10500), .A2(sram_rdata_b5[27]), .A3(n2820), .A4(
        sram_rdata_a5[27]), .Y(N226) );
  AO22X1_HVT U1797 ( .A1(n2630), .A2(sram_rdata_b5[28]), .A3(n2820), .A4(
        sram_rdata_a5[28]), .Y(N227) );
  AO22X1_HVT U1798 ( .A1(n2670), .A2(sram_rdata_b5[29]), .A3(n2290), .A4(
        sram_rdata_a5[29]), .Y(N228) );
  AO22X1_HVT U1799 ( .A1(n2680), .A2(sram_rdata_b5[30]), .A3(n2280), .A4(
        sram_rdata_a5[30]), .Y(N229) );
  AO22X1_HVT U1800 ( .A1(n2630), .A2(sram_rdata_b5[31]), .A3(n2360), .A4(
        sram_rdata_a5[31]), .Y(N230) );
  AO22X1_HVT U1801 ( .A1(n11900), .A2(sram_rdata_b6[0]), .A3(n2330), .A4(
        sram_rdata_a6[0]), .Y(N231) );
  AO22X1_HVT U1802 ( .A1(n14200), .A2(sram_rdata_b6[1]), .A3(n2820), .A4(
        sram_rdata_a6[1]), .Y(N232) );
  AO22X1_HVT U1803 ( .A1(n2660), .A2(sram_rdata_b6[2]), .A3(n2320), .A4(
        sram_rdata_a6[2]), .Y(N233) );
  AO22X1_HVT U1804 ( .A1(n2610), .A2(sram_rdata_b6[3]), .A3(n2360), .A4(
        sram_rdata_a6[3]), .Y(N234) );
  AO22X1_HVT U1805 ( .A1(n2620), .A2(sram_rdata_b6[4]), .A3(n1666), .A4(
        sram_rdata_a6[4]), .Y(N235) );
  AO22X1_HVT U1806 ( .A1(n2680), .A2(sram_rdata_b6[5]), .A3(n2360), .A4(
        sram_rdata_a6[5]), .Y(N236) );
  AO22X1_HVT U1807 ( .A1(n14300), .A2(sram_rdata_b6[6]), .A3(n2300), .A4(
        sram_rdata_a6[6]), .Y(N237) );
  AO22X1_HVT U1808 ( .A1(n1667), .A2(sram_rdata_b6[7]), .A3(n2310), .A4(
        sram_rdata_a6[7]), .Y(N238) );
  AO22X1_HVT U1809 ( .A1(n2630), .A2(sram_rdata_b6[8]), .A3(n2300), .A4(
        sram_rdata_a6[8]), .Y(N239) );
  AO22X1_HVT U1810 ( .A1(n14300), .A2(sram_rdata_b6[9]), .A3(n2340), .A4(
        sram_rdata_a6[9]), .Y(N240) );
  AO22X1_HVT U1811 ( .A1(n10500), .A2(sram_rdata_b6[10]), .A3(n2360), .A4(
        sram_rdata_a6[10]), .Y(N241) );
  AO22X1_HVT U1812 ( .A1(n10600), .A2(sram_rdata_b6[11]), .A3(n2320), .A4(
        sram_rdata_a6[11]), .Y(N242) );
  AO22X1_HVT U1813 ( .A1(n14300), .A2(sram_rdata_b6[12]), .A3(n14100), .A4(
        sram_rdata_a6[12]), .Y(N243) );
  AO22X1_HVT U1814 ( .A1(n10500), .A2(sram_rdata_b6[13]), .A3(n2310), .A4(
        sram_rdata_a6[13]), .Y(N244) );
  AO22X1_HVT U1815 ( .A1(n2660), .A2(sram_rdata_b6[14]), .A3(n2300), .A4(
        sram_rdata_a6[14]), .Y(N245) );
  AO22X1_HVT U1816 ( .A1(n2610), .A2(sram_rdata_b6[15]), .A3(n2280), .A4(
        sram_rdata_a6[15]), .Y(N246) );
  AO22X1_HVT U1817 ( .A1(n10600), .A2(sram_rdata_b6[16]), .A3(n2340), .A4(
        sram_rdata_a6[16]), .Y(N247) );
  AO22X1_HVT U1818 ( .A1(n2650), .A2(sram_rdata_b6[17]), .A3(n2330), .A4(
        sram_rdata_a6[17]), .Y(N248) );
  AO22X1_HVT U1819 ( .A1(n2650), .A2(sram_rdata_b6[18]), .A3(n2820), .A4(
        sram_rdata_a6[18]), .Y(N249) );
  AO22X1_HVT U1820 ( .A1(n2600), .A2(sram_rdata_b6[19]), .A3(n2280), .A4(
        sram_rdata_a6[19]), .Y(N250) );
  AO22X1_HVT U1821 ( .A1(n2600), .A2(sram_rdata_b6[20]), .A3(n2360), .A4(
        sram_rdata_a6[20]), .Y(N251) );
  AO22X1_HVT U1822 ( .A1(n14300), .A2(sram_rdata_b6[21]), .A3(n595), .A4(
        sram_rdata_a6[21]), .Y(N252) );
  AO22X1_HVT U1823 ( .A1(n2680), .A2(sram_rdata_b6[22]), .A3(n2340), .A4(
        sram_rdata_a6[22]), .Y(N253) );
  AO22X1_HVT U1824 ( .A1(n2630), .A2(sram_rdata_b6[23]), .A3(n2310), .A4(
        sram_rdata_a6[23]), .Y(N254) );
  AO22X1_HVT U1825 ( .A1(n1667), .A2(sram_rdata_b6[24]), .A3(n2310), .A4(
        sram_rdata_a6[24]), .Y(N255) );
  AO22X1_HVT U1826 ( .A1(n14200), .A2(sram_rdata_b6[25]), .A3(n2360), .A4(
        sram_rdata_a6[25]), .Y(N256) );
  AO22X1_HVT U1827 ( .A1(n14200), .A2(sram_rdata_b6[26]), .A3(n2330), .A4(
        sram_rdata_a6[26]), .Y(N257) );
  AO22X1_HVT U1828 ( .A1(n11900), .A2(sram_rdata_b6[27]), .A3(n2340), .A4(
        sram_rdata_a6[27]), .Y(N258) );
  AO22X1_HVT U1829 ( .A1(n1667), .A2(sram_rdata_b6[28]), .A3(n2280), .A4(
        sram_rdata_a6[28]), .Y(N259) );
  AO22X1_HVT U1830 ( .A1(n14300), .A2(sram_rdata_b6[29]), .A3(n2310), .A4(
        sram_rdata_a6[29]), .Y(N260) );
  AO22X1_HVT U1831 ( .A1(n2650), .A2(sram_rdata_b6[30]), .A3(n2350), .A4(
        sram_rdata_a6[30]), .Y(N261) );
  AO22X1_HVT U1832 ( .A1(n2600), .A2(sram_rdata_b6[31]), .A3(n2340), .A4(
        sram_rdata_a6[31]), .Y(N262) );
  AO22X1_HVT U1833 ( .A1(n11900), .A2(sram_rdata_b7[0]), .A3(n2330), .A4(
        sram_rdata_a7[0]), .Y(N263) );
  AO22X1_HVT U1834 ( .A1(n2660), .A2(sram_rdata_b7[1]), .A3(n2280), .A4(
        sram_rdata_a7[1]), .Y(N264) );
  AO22X1_HVT U1835 ( .A1(n14200), .A2(sram_rdata_b7[2]), .A3(n2280), .A4(
        sram_rdata_a7[2]), .Y(N265) );
  AO22X1_HVT U1836 ( .A1(n2620), .A2(sram_rdata_b7[3]), .A3(n1666), .A4(
        sram_rdata_a7[3]), .Y(N266) );
  AO22X1_HVT U1837 ( .A1(n2610), .A2(sram_rdata_b7[4]), .A3(n2320), .A4(
        sram_rdata_a7[4]), .Y(N267) );
  AO22X1_HVT U1838 ( .A1(n14200), .A2(sram_rdata_b7[5]), .A3(n2320), .A4(
        sram_rdata_a7[5]), .Y(N268) );
  AO22X1_HVT U1839 ( .A1(n2660), .A2(sram_rdata_b7[6]), .A3(n2820), .A4(
        sram_rdata_a7[6]), .Y(N269) );
  AO22X1_HVT U1840 ( .A1(n2610), .A2(sram_rdata_b7[7]), .A3(n14100), .A4(
        sram_rdata_a7[7]), .Y(N270) );
  AO22X1_HVT U1841 ( .A1(n2670), .A2(sram_rdata_b7[8]), .A3(n2350), .A4(
        sram_rdata_a7[8]), .Y(N271) );
  AO22X1_HVT U1842 ( .A1(n2650), .A2(sram_rdata_b7[9]), .A3(n2820), .A4(
        sram_rdata_a7[9]), .Y(N272) );
  AO22X1_HVT U1843 ( .A1(n10500), .A2(sram_rdata_b7[10]), .A3(n2290), .A4(
        sram_rdata_a7[10]), .Y(N273) );
  AO22X1_HVT U1844 ( .A1(n10600), .A2(sram_rdata_b7[11]), .A3(n2280), .A4(
        sram_rdata_a7[11]), .Y(N274) );
  AO22X1_HVT U1845 ( .A1(n2600), .A2(sram_rdata_b7[12]), .A3(n2300), .A4(
        sram_rdata_a7[12]), .Y(N275) );
  AO22X1_HVT U1846 ( .A1(n10500), .A2(sram_rdata_b7[13]), .A3(n2330), .A4(
        sram_rdata_a7[13]), .Y(N276) );
  AO22X1_HVT U1847 ( .A1(n14200), .A2(sram_rdata_b7[14]), .A3(n1666), .A4(
        sram_rdata_a7[14]), .Y(N277) );
  AO22X1_HVT U1848 ( .A1(n2670), .A2(sram_rdata_b7[15]), .A3(n2340), .A4(
        sram_rdata_a7[15]), .Y(N278) );
  AO22X1_HVT U1849 ( .A1(n10600), .A2(sram_rdata_b7[16]), .A3(n2350), .A4(
        sram_rdata_a7[16]), .Y(N279) );
  AO22X1_HVT U1850 ( .A1(n2680), .A2(sram_rdata_b7[17]), .A3(n2290), .A4(
        sram_rdata_a7[17]), .Y(N280) );
  AO22X1_HVT U1851 ( .A1(n14300), .A2(sram_rdata_b7[18]), .A3(n2280), .A4(
        sram_rdata_a7[18]), .Y(N281) );
  AO22X1_HVT U1852 ( .A1(n1667), .A2(sram_rdata_b7[19]), .A3(n2300), .A4(
        sram_rdata_a7[19]), .Y(N282) );
  AO22X1_HVT U1853 ( .A1(n2630), .A2(sram_rdata_b7[20]), .A3(n2320), .A4(
        sram_rdata_a7[20]), .Y(N283) );
  AO22X1_HVT U1854 ( .A1(n2650), .A2(sram_rdata_b7[21]), .A3(n2340), .A4(
        sram_rdata_a7[21]), .Y(N284) );
  AO22X1_HVT U1855 ( .A1(n2650), .A2(sram_rdata_b7[22]), .A3(n2820), .A4(
        sram_rdata_a7[22]), .Y(N285) );
  AO22X1_HVT U1856 ( .A1(n2600), .A2(sram_rdata_b7[23]), .A3(n2360), .A4(
        sram_rdata_a7[23]), .Y(N286) );
  AO22X1_HVT U1857 ( .A1(n2600), .A2(sram_rdata_b7[24]), .A3(n2360), .A4(
        sram_rdata_a7[24]), .Y(N287) );
  AO22X1_HVT U1858 ( .A1(n2660), .A2(sram_rdata_b7[25]), .A3(n2360), .A4(
        sram_rdata_a7[25]), .Y(N288) );
  AO22X1_HVT U1859 ( .A1(n2670), .A2(sram_rdata_b7[26]), .A3(n2330), .A4(
        sram_rdata_a7[26]), .Y(N289) );
  AO22X1_HVT U1860 ( .A1(n11900), .A2(sram_rdata_b7[27]), .A3(n2280), .A4(
        sram_rdata_a7[27]), .Y(N290) );
  AO22X1_HVT U1861 ( .A1(n2610), .A2(sram_rdata_b7[28]), .A3(n2290), .A4(
        sram_rdata_a7[28]), .Y(N291) );
  AO22X1_HVT U1862 ( .A1(n2670), .A2(sram_rdata_b7[29]), .A3(n2330), .A4(
        sram_rdata_a7[29]), .Y(N292) );
  AO22X1_HVT U1863 ( .A1(n14300), .A2(sram_rdata_b7[30]), .A3(n2350), .A4(
        sram_rdata_a7[30]), .Y(N293) );
  AO22X1_HVT U1864 ( .A1(n10500), .A2(sram_rdata_b7[31]), .A3(n2320), .A4(
        sram_rdata_a7[31]), .Y(N294) );
  AO22X1_HVT U1865 ( .A1(n11900), .A2(sram_rdata_b8[0]), .A3(n2290), .A4(
        sram_rdata_a8[0]), .Y(N295) );
  AO22X1_HVT U1866 ( .A1(n14300), .A2(sram_rdata_b8[1]), .A3(n2290), .A4(
        sram_rdata_a8[1]), .Y(N296) );
  AO22X1_HVT U1867 ( .A1(n2680), .A2(sram_rdata_b8[2]), .A3(n2360), .A4(
        sram_rdata_a8[2]), .Y(N297) );
  AO22X1_HVT U1868 ( .A1(n2630), .A2(sram_rdata_b8[3]), .A3(n2330), .A4(
        sram_rdata_a8[3]), .Y(N298) );
  AO22X1_HVT U1869 ( .A1(n1667), .A2(sram_rdata_b8[4]), .A3(n595), .A4(
        sram_rdata_a8[4]), .Y(N299) );
  AO22X1_HVT U1870 ( .A1(n2660), .A2(sram_rdata_b8[5]), .A3(n2310), .A4(
        sram_rdata_a8[5]), .Y(N300) );
  AO22X1_HVT U1871 ( .A1(n14200), .A2(sram_rdata_b8[6]), .A3(n2300), .A4(
        sram_rdata_a8[6]), .Y(N301) );
  AO22X1_HVT U1872 ( .A1(n2670), .A2(sram_rdata_b8[7]), .A3(n2350), .A4(
        sram_rdata_a8[7]), .Y(N302) );
  AO22X1_HVT U1873 ( .A1(n2610), .A2(sram_rdata_b8[8]), .A3(n2340), .A4(
        sram_rdata_a8[8]), .Y(N303) );
  AO22X1_HVT U1874 ( .A1(n2680), .A2(sram_rdata_b8[9]), .A3(n2320), .A4(
        sram_rdata_a8[9]), .Y(N304) );
  AO22X1_HVT U1875 ( .A1(n10500), .A2(sram_rdata_b8[10]), .A3(n2320), .A4(
        sram_rdata_a8[10]), .Y(N305) );
  AO22X1_HVT U1876 ( .A1(n10600), .A2(sram_rdata_b8[11]), .A3(n2820), .A4(
        sram_rdata_a8[11]), .Y(N306) );
  AO22X1_HVT U1877 ( .A1(n2630), .A2(sram_rdata_b8[12]), .A3(n2300), .A4(
        sram_rdata_a8[12]), .Y(N307) );
  AO22X1_HVT U1878 ( .A1(n10500), .A2(sram_rdata_b8[13]), .A3(n1666), .A4(
        sram_rdata_a8[13]), .Y(N308) );
  AO22X1_HVT U1879 ( .A1(n2680), .A2(sram_rdata_b8[14]), .A3(n2300), .A4(
        sram_rdata_a8[14]), .Y(N309) );
  AO22X1_HVT U1880 ( .A1(n2630), .A2(sram_rdata_b8[15]), .A3(n2290), .A4(
        sram_rdata_a8[15]), .Y(N310) );
  AO22X1_HVT U1881 ( .A1(n10600), .A2(sram_rdata_b8[16]), .A3(n2290), .A4(
        sram_rdata_a8[16]), .Y(N311) );
  AO22X1_HVT U1882 ( .A1(n14200), .A2(sram_rdata_b8[17]), .A3(n2320), .A4(
        sram_rdata_a8[17]), .Y(N312) );
  AO22X1_HVT U1883 ( .A1(n2660), .A2(sram_rdata_b8[18]), .A3(n2280), .A4(
        sram_rdata_a8[18]), .Y(N313) );
  AO22X1_HVT U1884 ( .A1(n2610), .A2(sram_rdata_b8[19]), .A3(n2340), .A4(
        sram_rdata_a8[19]), .Y(N314) );
  AO22X1_HVT U1885 ( .A1(n2670), .A2(sram_rdata_b8[20]), .A3(n14100), .A4(
        sram_rdata_a8[20]), .Y(N315) );
  AO22X1_HVT U1886 ( .A1(n2680), .A2(sram_rdata_b8[21]), .A3(n2310), .A4(
        sram_rdata_a8[21]), .Y(N316) );
  AO22X1_HVT U1887 ( .A1(n14300), .A2(sram_rdata_b8[22]), .A3(n2300), .A4(
        sram_rdata_a8[22]), .Y(N317) );
  AO22X1_HVT U1888 ( .A1(n1667), .A2(sram_rdata_b8[23]), .A3(n2280), .A4(
        sram_rdata_a8[23]), .Y(N318) );
  AO22X1_HVT U1889 ( .A1(n2630), .A2(sram_rdata_b8[24]), .A3(n2820), .A4(
        sram_rdata_a8[24]), .Y(N319) );
  AO22X1_HVT U1890 ( .A1(n14300), .A2(sram_rdata_b8[25]), .A3(n2340), .A4(
        sram_rdata_a8[25]), .Y(N320) );
  AO22X1_HVT U1891 ( .A1(n14300), .A2(sram_rdata_b8[26]), .A3(n2330), .A4(
        sram_rdata_a8[26]), .Y(N321) );
  AO22X1_HVT U1892 ( .A1(n11900), .A2(sram_rdata_b8[27]), .A3(n2320), .A4(
        sram_rdata_a8[27]), .Y(N322) );
  AO22X1_HVT U1893 ( .A1(n14200), .A2(sram_rdata_b8[28]), .A3(n1666), .A4(
        sram_rdata_a8[28]), .Y(N323) );
  AO22X1_HVT U1894 ( .A1(n14200), .A2(sram_rdata_b8[29]), .A3(n2350), .A4(
        sram_rdata_a8[29]), .Y(N324) );
  AO22X1_HVT U1895 ( .A1(n2660), .A2(sram_rdata_b8[30]), .A3(n2330), .A4(
        sram_rdata_a8[30]), .Y(N325) );
  AO22X1_HVT U1896 ( .A1(n2610), .A2(sram_rdata_b8[31]), .A3(n2310), .A4(
        sram_rdata_a8[31]), .Y(N326) );
  AO22X1_HVT U1897 ( .A1(n11900), .A2(sram_rdata_b0[0]), .A3(n2290), .A4(
        sram_rdata_a0[0]), .Y(N39) );
  AO22X1_HVT U1898 ( .A1(n2650), .A2(sram_rdata_b0[1]), .A3(n2350), .A4(
        sram_rdata_a0[1]), .Y(N40) );
  AO22X1_HVT U1899 ( .A1(n2650), .A2(sram_rdata_b0[2]), .A3(n2350), .A4(
        sram_rdata_a0[2]), .Y(N41) );
  AO22X1_HVT U1900 ( .A1(n2600), .A2(sram_rdata_b0[3]), .A3(n2820), .A4(
        sram_rdata_a0[3]), .Y(N42) );
  AO22X1_HVT U1901 ( .A1(n2600), .A2(sram_rdata_b0[4]), .A3(n2300), .A4(
        sram_rdata_a0[4]), .Y(N43) );
  AO22X1_HVT U1902 ( .A1(n14300), .A2(sram_rdata_b0[5]), .A3(n2310), .A4(
        sram_rdata_a0[5]), .Y(N44) );
  AO22X1_HVT U1903 ( .A1(n2680), .A2(sram_rdata_b0[6]), .A3(n2360), .A4(
        sram_rdata_a0[6]), .Y(N45) );
  AO22X1_HVT U1904 ( .A1(n2630), .A2(sram_rdata_b0[7]), .A3(n2340), .A4(
        sram_rdata_a0[7]), .Y(N46) );
  AO22X1_HVT U1905 ( .A1(n1667), .A2(sram_rdata_b0[8]), .A3(n2320), .A4(
        sram_rdata_a0[8]), .Y(N47) );
  AO22X1_HVT U1906 ( .A1(n14200), .A2(sram_rdata_b0[9]), .A3(n2310), .A4(
        sram_rdata_a0[9]), .Y(N48) );
  AO22X1_HVT U1907 ( .A1(n10500), .A2(sram_rdata_b0[10]), .A3(n2280), .A4(
        sram_rdata_a0[10]), .Y(N49) );
  AO22X1_HVT U1908 ( .A1(n10600), .A2(sram_rdata_b0[11]), .A3(n2360), .A4(
        sram_rdata_a0[11]), .Y(N50) );
  AO22X1_HVT U1909 ( .A1(n1667), .A2(sram_rdata_b0[12]), .A3(n2330), .A4(
        sram_rdata_a0[12]), .Y(N51) );
  AO22X1_HVT U1910 ( .A1(n10500), .A2(sram_rdata_b0[13]), .A3(n14100), .A4(
        sram_rdata_a0[13]), .Y(N52) );
  AO22X1_HVT U1911 ( .A1(n2650), .A2(sram_rdata_b0[14]), .A3(n2320), .A4(
        sram_rdata_a0[14]), .Y(N53) );
  AO22X1_HVT U1912 ( .A1(n2600), .A2(sram_rdata_b0[15]), .A3(n1666), .A4(
        sram_rdata_a0[15]), .Y(N54) );
  AO22X1_HVT U1913 ( .A1(n10600), .A2(sram_rdata_b0[16]), .A3(n1666), .A4(
        sram_rdata_a0[16]), .Y(N55) );
  AO22X1_HVT U1914 ( .A1(n2660), .A2(sram_rdata_b0[17]), .A3(n2360), .A4(
        sram_rdata_a0[17]), .Y(N56) );
  AO22X1_HVT U1915 ( .A1(n14200), .A2(sram_rdata_b0[18]), .A3(n2300), .A4(
        sram_rdata_a0[18]), .Y(N57) );
  AO22X1_HVT U1916 ( .A1(n2670), .A2(sram_rdata_b0[19]), .A3(n2310), .A4(
        sram_rdata_a0[19]), .Y(N58) );
  AO22X1_HVT U1917 ( .A1(n2610), .A2(sram_rdata_b0[20]), .A3(n2300), .A4(
        sram_rdata_a0[20]), .Y(N59) );
  AO22X1_HVT U1918 ( .A1(n14200), .A2(sram_rdata_b0[21]), .A3(n2340), .A4(
        sram_rdata_a0[21]), .Y(N60) );
  AO22X1_HVT U1919 ( .A1(n2660), .A2(sram_rdata_b0[22]), .A3(n2360), .A4(
        sram_rdata_a0[22]), .Y(N61) );
  AO22X1_HVT U1920 ( .A1(n2610), .A2(sram_rdata_b0[23]), .A3(n2330), .A4(
        sram_rdata_a0[23]), .Y(N62) );
  AO22X1_HVT U1921 ( .A1(n2620), .A2(sram_rdata_b0[24]), .A3(n2820), .A4(
        sram_rdata_a0[24]), .Y(N63) );
  AO22X1_HVT U1922 ( .A1(n2650), .A2(sram_rdata_b0[25]), .A3(n2290), .A4(
        sram_rdata_a0[25]), .Y(N64) );
  AO22X1_HVT U1923 ( .A1(n2670), .A2(sram_rdata_b0[26]), .A3(n2280), .A4(
        sram_rdata_a0[26]), .Y(N65) );
  AO22X1_HVT U1924 ( .A1(n11900), .A2(sram_rdata_b0[27]), .A3(n2310), .A4(
        sram_rdata_a0[27]), .Y(N66) );
  AO22X1_HVT U1925 ( .A1(n2600), .A2(sram_rdata_b0[28]), .A3(n2320), .A4(
        sram_rdata_a0[28]), .Y(N67) );
  AO22X1_HVT U1926 ( .A1(n2670), .A2(sram_rdata_b0[29]), .A3(n2330), .A4(
        sram_rdata_a0[29]), .Y(N68) );
  AO22X1_HVT U1927 ( .A1(n14200), .A2(sram_rdata_b0[30]), .A3(n14100), .A4(
        sram_rdata_a0[30]), .Y(N69) );
  AO22X1_HVT U1928 ( .A1(n2620), .A2(sram_rdata_b0[31]), .A3(n2350), .A4(
        sram_rdata_a0[31]), .Y(N70) );
  AO22X1_HVT U1929 ( .A1(n11900), .A2(sram_rdata_b1[0]), .A3(n2320), .A4(
        sram_rdata_a1[0]), .Y(N71) );
  AO22X1_HVT U1930 ( .A1(n2680), .A2(sram_rdata_b1[1]), .A3(n2340), .A4(
        sram_rdata_a1[1]), .Y(N72) );
  AO22X1_HVT U1931 ( .A1(n14300), .A2(sram_rdata_b1[2]), .A3(n2340), .A4(
        sram_rdata_a1[2]), .Y(N73) );
  AO22X1_HVT U1932 ( .A1(n1667), .A2(sram_rdata_b1[3]), .A3(n2310), .A4(
        sram_rdata_a1[3]), .Y(N74) );
  AO22X1_HVT U1933 ( .A1(n2630), .A2(sram_rdata_b1[4]), .A3(n2280), .A4(
        sram_rdata_a1[4]), .Y(N75) );
  AO22X1_HVT U1934 ( .A1(n2650), .A2(sram_rdata_b1[5]), .A3(n595), .A4(
        sram_rdata_a1[5]), .Y(N76) );
  AO22X1_HVT U1935 ( .A1(n2650), .A2(sram_rdata_b1[6]), .A3(n2820), .A4(
        sram_rdata_a1[6]), .Y(N77) );
  AO22X1_HVT U1936 ( .A1(n2600), .A2(sram_rdata_b1[7]), .A3(n2320), .A4(
        sram_rdata_a1[7]), .Y(N78) );
  AO22X1_HVT U1937 ( .A1(n2600), .A2(sram_rdata_b1[8]), .A3(n2280), .A4(
        sram_rdata_a1[8]), .Y(N79) );
  AO22X1_HVT U1938 ( .A1(n2660), .A2(sram_rdata_b1[9]), .A3(n2310), .A4(
        sram_rdata_a1[9]), .Y(N80) );
  AO22X1_HVT U1939 ( .A1(n10500), .A2(sram_rdata_b1[10]), .A3(n2350), .A4(
        sram_rdata_a1[10]), .Y(N81) );
  AO22X1_HVT U1940 ( .A1(n10600), .A2(sram_rdata_b1[11]), .A3(n2320), .A4(
        sram_rdata_a1[11]), .Y(N82) );
  AO22X1_HVT U1941 ( .A1(n2610), .A2(sram_rdata_b1[12]), .A3(n2320), .A4(
        sram_rdata_a1[12]), .Y(N83) );
  AO22X1_HVT U1942 ( .A1(n10500), .A2(sram_rdata_b1[13]), .A3(n2290), .A4(
        sram_rdata_a1[13]), .Y(N84) );
  AO22X1_HVT U1943 ( .A1(n14300), .A2(sram_rdata_b1[14]), .A3(n2300), .A4(
        sram_rdata_a1[14]), .Y(N85) );
  AO22X1_HVT U1944 ( .A1(n2620), .A2(sram_rdata_b1[15]), .A3(n2640), .A4(
        sram_rdata_a1[15]), .Y(N86) );
  AO22X1_HVT U1945 ( .A1(n10600), .A2(sram_rdata_b1[16]), .A3(n2320), .A4(
        sram_rdata_a1[16]), .Y(N87) );
  AO22X1_HVT U1946 ( .A1(n14300), .A2(sram_rdata_b1[17]), .A3(n2320), .A4(
        sram_rdata_a1[17]), .Y(N88) );
  AO22X1_HVT U1947 ( .A1(n2680), .A2(sram_rdata_b1[18]), .A3(n2820), .A4(
        sram_rdata_a1[18]), .Y(N89) );
  AO22X1_HVT U1948 ( .A1(n2630), .A2(sram_rdata_b1[19]), .A3(n2350), .A4(
        sram_rdata_a1[19]), .Y(N90) );
  AO22X1_HVT U1949 ( .A1(n1667), .A2(sram_rdata_b1[20]), .A3(n2350), .A4(
        sram_rdata_a1[20]), .Y(N91) );
  AO22X1_HVT U1950 ( .A1(n2660), .A2(sram_rdata_b1[21]), .A3(n2340), .A4(
        sram_rdata_a1[21]), .Y(N92) );
  AO22X1_HVT U1951 ( .A1(n14200), .A2(sram_rdata_b1[22]), .A3(n2300), .A4(
        sram_rdata_a1[22]), .Y(N93) );
  AO22X1_HVT U1952 ( .A1(n2620), .A2(sram_rdata_b1[23]), .A3(n2290), .A4(
        sram_rdata_a1[23]), .Y(N94) );
  AO22X1_HVT U1953 ( .A1(n2610), .A2(sram_rdata_b1[24]), .A3(n2280), .A4(
        sram_rdata_a1[24]), .Y(N95) );
  AO22X1_HVT U1954 ( .A1(n2680), .A2(sram_rdata_b1[25]), .A3(n2340), .A4(
        sram_rdata_a1[25]), .Y(N96) );
  AO22X1_HVT U1955 ( .A1(n2650), .A2(sram_rdata_b1[26]), .A3(n2300), .A4(
        sram_rdata_a1[26]), .Y(N97) );
  AO22X1_HVT U1956 ( .A1(n11900), .A2(sram_rdata_b1[27]), .A3(n2820), .A4(
        sram_rdata_a1[27]), .Y(N98) );
  AO22X1_HVT U1957 ( .A1(n2630), .A2(sram_rdata_b1[28]), .A3(n2310), .A4(
        sram_rdata_a1[28]), .Y(N99) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_0 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22041, n1;

  AND2X1_HVT main_gate ( .A1(net22041), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n1), .D(EN), .Q(net22041) );
  INVX0_HVT U1 ( .A(CLK), .Y(n1) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_20 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22041, n2;

  AND2X1_HVT main_gate ( .A1(net22041), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22041) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_19 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22041, n2;

  AND2X1_HVT main_gate ( .A1(net22041), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22041) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_18 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22041, n2;

  AND2X1_HVT main_gate ( .A1(net22041), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22041) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_17 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22041, n2;

  AND2X1_HVT main_gate ( .A1(net22041), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22041) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_16 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22041, n2;

  AND2X1_HVT main_gate ( .A1(net22041), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22041) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_15 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22041, n2;

  AND2X1_HVT main_gate ( .A1(net22041), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22041) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_14 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22041, n2;

  AND2X1_HVT main_gate ( .A1(net22041), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22041) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_13 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22041, n2;

  AND2X1_HVT main_gate ( .A1(net22041), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22041) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_12 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22041, n2;

  AND2X1_HVT main_gate ( .A1(net22041), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22041) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_11 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22041, n2;

  AND2X1_HVT main_gate ( .A1(net22041), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22041) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_10 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22041, n2;

  AND2X1_HVT main_gate ( .A1(net22041), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22041) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_9 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22041, n2;

  AND2X1_HVT main_gate ( .A1(net22041), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22041) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_8 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22041, n2;

  AND2X1_HVT main_gate ( .A1(net22041), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22041) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_7 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22041, n2;

  AND2X1_HVT main_gate ( .A1(net22041), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22041) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_6 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22041, n2;

  AND2X1_HVT main_gate ( .A1(net22041), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22041) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_5 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22041, n2;

  AND2X1_HVT main_gate ( .A1(net22041), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22041) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_4 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22041, n2;

  AND2X1_HVT main_gate ( .A1(net22041), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22041) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_3 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22041, n2;

  AND2X1_HVT main_gate ( .A1(net22041), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22041) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_2 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22041, n2;

  AND2X1_HVT main_gate ( .A1(net22041), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22041) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_1 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22041, n2;

  AND2X1_HVT main_gate ( .A1(net22041), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22041) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module bias_sel ( clk, srstn, mode, load_conv1_bias_enable, 
        load_conv2_bias0_enable, load_conv2_bias1_enable, sram_rdata_weight, 
        bias_data, conv1_bias_set_5_, conv1_bias_set_4_, conv1_bias_set_3_, 
        conv1_bias_set_2_, conv1_bias_set_1_, conv1_bias_set_0_, set_5_, 
        set_4_, set_3_, set_2_, set_1_, set_0_ );
  input [1:0] mode;
  input [99:0] sram_rdata_weight;
  output [3:0] bias_data;
  input clk, srstn, load_conv1_bias_enable, load_conv2_bias0_enable,
         load_conv2_bias1_enable, conv1_bias_set_5_, conv1_bias_set_4_,
         conv1_bias_set_3_, conv1_bias_set_2_, conv1_bias_set_1_,
         conv1_bias_set_0_, set_5_, set_4_, set_3_, set_2_, set_1_, set_0_;
  wire   net22070, net22073, net22074, net22075, net22076, net22077, net22078,
         net22079, net22080, net22081, net22084, net22089, net22090, net22091,
         net22092, net22093, net22094, net22095, net22096, net22097, net22098,
         net22101, net22106, net22107, net22108, net22109, net22110, net22111,
         net22112, net22113, net22114, net22115, net22118, net22123, net22124,
         net22125, net22126, net22127, net22128, net22129, net22130, net22131,
         net22132, net22135, net22140, net22141, net22142, net22143, net22144,
         net22145, net22146, net22147, net22148, net22149, net22152, net22157,
         net22158, net22159, net22160, net22161, net22162, net22163, net22164,
         net22165, net22166, net22169, net22174, net22175, net22176, net22177,
         net22178, net22179, net22180, net22181, net22182, net22183, net22186,
         net22191, net22192, net22193, net22194, net22195, net22196, net22197,
         net22198, net22199, net22200, net22203, net22208, net22209, net22210,
         net22211, net22212, net22213, net22214, net22215, net22216, net22217,
         net22220, net22224, net22225, net22226, net22227, net22228, net22229,
         net22230, net22231, net22232, net22233, net22234, net22237, net22250,
         net22251, net22252, net22253, net22254, net22255, net22256, net22257,
         net22258, net22259, net22262, net22267, net22268, net22269, net22270,
         net22271, net22272, net22273, net22274, net22275, net22276, net22279,
         net22284, net22285, net22286, net22287, net22288, net22289, net22290,
         net22291, net22292, net22293, net22296, net22301, net22302, net22303,
         net22304, net22305, net22306, net22307, net22308, net22309, net22310,
         net22313, net22318, net22319, net22320, net22321, net22322, net22323,
         net22324, net22325, net22326, net22327, net22330, net22335, net22336,
         net22337, net22338, net22339, net22340, net22341, net22342, net22343,
         net22344, net22347, net22352, net22353, net22354, net22355, net22356,
         net22357, net22358, net22359, net22360, net22361, net22364, net22369,
         net22370, net22371, net22372, net22373, net22374, net22375, net22376,
         net22377, net22378, net22381, net22386, net22387, net22388, net22389,
         net22390, net22391, net22392, net22393, net22394, net22395, net22398,
         net22402, net22403, net22404, net22405, net22406, net22407, net22408,
         net22409, net22410, net22411, net22412, net22415, net22426, net22432,
         net22436, net22440, net22444, net22447, n305, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403;
  wire   [199:0] conv_weight_box;
  wire   [99:0] delay_weight;

  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_0 clk_gate_conv_weight_box_reg_0_ ( 
        .CLK(clk), .EN(net22224), .ENCLK(net22084) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_20 clk_gate_conv_weight_box_reg_2_ ( 
        .CLK(clk), .EN(net22224), .ENCLK(net22101) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_19 clk_gate_conv_weight_box_reg_5_ ( 
        .CLK(clk), .EN(net22224), .ENCLK(net22118) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_18 clk_gate_conv_weight_box_reg_7_ ( 
        .CLK(clk), .EN(net22224), .ENCLK(net22135) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_17 clk_gate_conv_weight_box_reg_10_ ( 
        .CLK(clk), .EN(net22224), .ENCLK(net22152) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_16 clk_gate_conv_weight_box_reg_12_ ( 
        .CLK(clk), .EN(net22224), .ENCLK(net22169) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_15 clk_gate_conv_weight_box_reg_15_ ( 
        .CLK(clk), .EN(net22224), .ENCLK(net22186) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_14 clk_gate_conv_weight_box_reg_17_ ( 
        .CLK(clk), .EN(net22224), .ENCLK(net22203) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_13 clk_gate_conv_weight_box_reg_20_ ( 
        .CLK(clk), .EN(net22224), .ENCLK(net22220) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_12 clk_gate_conv_weight_box_reg_22_ ( 
        .CLK(clk), .EN(net22224), .ENCLK(net22237) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_11 clk_gate_conv_weight_box_reg_25_ ( 
        .CLK(clk), .EN(net22402), .ENCLK(net22262) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_10 clk_gate_conv_weight_box_reg_27_ ( 
        .CLK(clk), .EN(net22402), .ENCLK(net22279) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_9 clk_gate_conv_weight_box_reg_30_ ( 
        .CLK(clk), .EN(net22402), .ENCLK(net22296) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_8 clk_gate_conv_weight_box_reg_32_ ( 
        .CLK(clk), .EN(net22402), .ENCLK(net22313) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_7 clk_gate_conv_weight_box_reg_35_ ( 
        .CLK(clk), .EN(net22402), .ENCLK(net22330) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_6 clk_gate_conv_weight_box_reg_37_ ( 
        .CLK(clk), .EN(net22402), .ENCLK(net22347) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_5 clk_gate_conv_weight_box_reg_40_ ( 
        .CLK(clk), .EN(net22402), .ENCLK(net22364) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_4 clk_gate_conv_weight_box_reg_42_ ( 
        .CLK(clk), .EN(net22402), .ENCLK(net22381) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_3 clk_gate_conv_weight_box_reg_45_ ( 
        .CLK(clk), .EN(net22402), .ENCLK(net22398) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_2 clk_gate_conv_weight_box_reg_47_ ( 
        .CLK(clk), .EN(net22402), .ENCLK(net22415) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_1 clk_gate_bias_data_reg ( .CLK(clk), 
        .EN(net22426), .ENCLK(net22447) );
  DFFSSRX1_HVT delay_weight_reg_99_ ( .D(1'b0), .SETB(n117), .RSTB(
        sram_rdata_weight[99]), .CLK(clk), .Q(delay_weight[99]) );
  DFFSSRX1_HVT delay_weight_reg_98_ ( .D(1'b0), .SETB(n113), .RSTB(
        sram_rdata_weight[98]), .CLK(clk), .Q(delay_weight[98]) );
  DFFSSRX1_HVT delay_weight_reg_97_ ( .D(1'b0), .SETB(n108), .RSTB(
        sram_rdata_weight[97]), .CLK(clk), .Q(delay_weight[97]) );
  DFFSSRX1_HVT delay_weight_reg_96_ ( .D(1'b0), .SETB(n118), .RSTB(
        sram_rdata_weight[96]), .CLK(clk), .Q(delay_weight[96]) );
  DFFSSRX1_HVT delay_weight_reg_95_ ( .D(1'b0), .SETB(n114), .RSTB(
        sram_rdata_weight[95]), .CLK(clk), .Q(delay_weight[95]) );
  DFFSSRX1_HVT delay_weight_reg_94_ ( .D(1'b0), .SETB(n109), .RSTB(
        sram_rdata_weight[94]), .CLK(clk), .Q(delay_weight[94]) );
  DFFSSRX1_HVT delay_weight_reg_93_ ( .D(1'b0), .SETB(n119), .RSTB(
        sram_rdata_weight[93]), .CLK(clk), .Q(delay_weight[93]) );
  DFFSSRX1_HVT delay_weight_reg_92_ ( .D(1'b0), .SETB(n115), .RSTB(
        sram_rdata_weight[92]), .CLK(clk), .Q(delay_weight[92]) );
  DFFSSRX1_HVT delay_weight_reg_91_ ( .D(1'b0), .SETB(n110), .RSTB(
        sram_rdata_weight[91]), .CLK(clk), .Q(delay_weight[91]) );
  DFFSSRX1_HVT delay_weight_reg_90_ ( .D(1'b0), .SETB(n116), .RSTB(
        sram_rdata_weight[90]), .CLK(clk), .Q(delay_weight[90]) );
  DFFSSRX1_HVT delay_weight_reg_89_ ( .D(1'b0), .SETB(n112), .RSTB(
        sram_rdata_weight[89]), .CLK(clk), .Q(delay_weight[89]) );
  DFFSSRX1_HVT delay_weight_reg_88_ ( .D(1'b0), .SETB(n107), .RSTB(
        sram_rdata_weight[88]), .CLK(clk), .Q(delay_weight[88]) );
  DFFSSRX1_HVT delay_weight_reg_87_ ( .D(1'b0), .SETB(n117), .RSTB(
        sram_rdata_weight[87]), .CLK(clk), .Q(delay_weight[87]) );
  DFFSSRX1_HVT delay_weight_reg_86_ ( .D(1'b0), .SETB(n113), .RSTB(
        sram_rdata_weight[86]), .CLK(clk), .Q(delay_weight[86]) );
  DFFSSRX1_HVT delay_weight_reg_85_ ( .D(1'b0), .SETB(n108), .RSTB(
        sram_rdata_weight[85]), .CLK(clk), .Q(delay_weight[85]) );
  DFFSSRX1_HVT delay_weight_reg_84_ ( .D(1'b0), .SETB(n118), .RSTB(
        sram_rdata_weight[84]), .CLK(clk), .Q(delay_weight[84]) );
  DFFSSRX1_HVT delay_weight_reg_83_ ( .D(1'b0), .SETB(n114), .RSTB(
        sram_rdata_weight[83]), .CLK(clk), .Q(delay_weight[83]) );
  DFFSSRX1_HVT delay_weight_reg_82_ ( .D(1'b0), .SETB(n109), .RSTB(
        sram_rdata_weight[82]), .CLK(clk), .Q(delay_weight[82]) );
  DFFSSRX1_HVT delay_weight_reg_81_ ( .D(1'b0), .SETB(n119), .RSTB(
        sram_rdata_weight[81]), .CLK(clk), .Q(delay_weight[81]) );
  DFFSSRX1_HVT delay_weight_reg_80_ ( .D(1'b0), .SETB(n115), .RSTB(
        sram_rdata_weight[80]), .CLK(clk), .Q(delay_weight[80]) );
  DFFSSRX1_HVT delay_weight_reg_79_ ( .D(1'b0), .SETB(n110), .RSTB(
        sram_rdata_weight[79]), .CLK(clk), .Q(delay_weight[79]) );
  DFFSSRX1_HVT delay_weight_reg_78_ ( .D(1'b0), .SETB(n116), .RSTB(
        sram_rdata_weight[78]), .CLK(clk), .Q(delay_weight[78]) );
  DFFSSRX1_HVT delay_weight_reg_77_ ( .D(1'b0), .SETB(n112), .RSTB(
        sram_rdata_weight[77]), .CLK(clk), .Q(delay_weight[77]) );
  DFFSSRX1_HVT delay_weight_reg_76_ ( .D(1'b0), .SETB(n107), .RSTB(
        sram_rdata_weight[76]), .CLK(clk), .Q(delay_weight[76]) );
  DFFSSRX1_HVT delay_weight_reg_75_ ( .D(1'b0), .SETB(n117), .RSTB(
        sram_rdata_weight[75]), .CLK(clk), .Q(delay_weight[75]) );
  DFFSSRX1_HVT delay_weight_reg_74_ ( .D(1'b0), .SETB(n113), .RSTB(
        sram_rdata_weight[74]), .CLK(clk), .Q(delay_weight[74]) );
  DFFSSRX1_HVT delay_weight_reg_73_ ( .D(1'b0), .SETB(n108), .RSTB(
        sram_rdata_weight[73]), .CLK(clk), .Q(delay_weight[73]) );
  DFFSSRX1_HVT delay_weight_reg_72_ ( .D(1'b0), .SETB(n118), .RSTB(
        sram_rdata_weight[72]), .CLK(clk), .Q(delay_weight[72]) );
  DFFSSRX1_HVT delay_weight_reg_71_ ( .D(1'b0), .SETB(n114), .RSTB(
        sram_rdata_weight[71]), .CLK(clk), .Q(delay_weight[71]) );
  DFFSSRX1_HVT delay_weight_reg_70_ ( .D(1'b0), .SETB(n109), .RSTB(
        sram_rdata_weight[70]), .CLK(clk), .Q(delay_weight[70]) );
  DFFSSRX1_HVT delay_weight_reg_69_ ( .D(1'b0), .SETB(n119), .RSTB(
        sram_rdata_weight[69]), .CLK(clk), .Q(delay_weight[69]) );
  DFFSSRX1_HVT delay_weight_reg_68_ ( .D(1'b0), .SETB(n115), .RSTB(
        sram_rdata_weight[68]), .CLK(clk), .Q(delay_weight[68]) );
  DFFSSRX1_HVT delay_weight_reg_67_ ( .D(1'b0), .SETB(n110), .RSTB(
        sram_rdata_weight[67]), .CLK(clk), .Q(delay_weight[67]) );
  DFFSSRX1_HVT delay_weight_reg_66_ ( .D(1'b0), .SETB(n116), .RSTB(
        sram_rdata_weight[66]), .CLK(clk), .Q(delay_weight[66]) );
  DFFSSRX1_HVT delay_weight_reg_65_ ( .D(1'b0), .SETB(n112), .RSTB(
        sram_rdata_weight[65]), .CLK(clk), .Q(delay_weight[65]) );
  DFFSSRX1_HVT delay_weight_reg_64_ ( .D(1'b0), .SETB(n107), .RSTB(
        sram_rdata_weight[64]), .CLK(clk), .Q(delay_weight[64]) );
  DFFSSRX1_HVT delay_weight_reg_63_ ( .D(1'b0), .SETB(n117), .RSTB(
        sram_rdata_weight[63]), .CLK(clk), .Q(delay_weight[63]) );
  DFFSSRX1_HVT delay_weight_reg_62_ ( .D(1'b0), .SETB(n113), .RSTB(
        sram_rdata_weight[62]), .CLK(clk), .Q(delay_weight[62]) );
  DFFSSRX1_HVT delay_weight_reg_61_ ( .D(1'b0), .SETB(n108), .RSTB(
        sram_rdata_weight[61]), .CLK(clk), .Q(delay_weight[61]) );
  DFFSSRX1_HVT delay_weight_reg_60_ ( .D(1'b0), .SETB(n118), .RSTB(
        sram_rdata_weight[60]), .CLK(clk), .Q(delay_weight[60]) );
  DFFSSRX1_HVT delay_weight_reg_59_ ( .D(1'b0), .SETB(n114), .RSTB(
        sram_rdata_weight[59]), .CLK(clk), .Q(delay_weight[59]) );
  DFFSSRX1_HVT delay_weight_reg_58_ ( .D(1'b0), .SETB(n109), .RSTB(
        sram_rdata_weight[58]), .CLK(clk), .Q(delay_weight[58]) );
  DFFSSRX1_HVT delay_weight_reg_57_ ( .D(1'b0), .SETB(n119), .RSTB(
        sram_rdata_weight[57]), .CLK(clk), .Q(delay_weight[57]) );
  DFFSSRX1_HVT delay_weight_reg_56_ ( .D(1'b0), .SETB(n115), .RSTB(
        sram_rdata_weight[56]), .CLK(clk), .Q(delay_weight[56]) );
  DFFSSRX1_HVT delay_weight_reg_55_ ( .D(1'b0), .SETB(n110), .RSTB(
        sram_rdata_weight[55]), .CLK(clk), .Q(delay_weight[55]) );
  DFFSSRX1_HVT delay_weight_reg_54_ ( .D(1'b0), .SETB(n116), .RSTB(
        sram_rdata_weight[54]), .CLK(clk), .Q(delay_weight[54]) );
  DFFSSRX1_HVT delay_weight_reg_53_ ( .D(1'b0), .SETB(n112), .RSTB(
        sram_rdata_weight[53]), .CLK(clk), .Q(delay_weight[53]) );
  DFFSSRX1_HVT delay_weight_reg_52_ ( .D(1'b0), .SETB(n107), .RSTB(
        sram_rdata_weight[52]), .CLK(clk), .Q(delay_weight[52]) );
  DFFSSRX1_HVT delay_weight_reg_51_ ( .D(1'b0), .SETB(n117), .RSTB(
        sram_rdata_weight[51]), .CLK(clk), .Q(delay_weight[51]) );
  DFFSSRX1_HVT delay_weight_reg_50_ ( .D(1'b0), .SETB(n113), .RSTB(
        sram_rdata_weight[50]), .CLK(clk), .Q(delay_weight[50]) );
  DFFSSRX1_HVT delay_weight_reg_49_ ( .D(1'b0), .SETB(n108), .RSTB(
        sram_rdata_weight[49]), .CLK(clk), .Q(delay_weight[49]) );
  DFFSSRX1_HVT delay_weight_reg_48_ ( .D(1'b0), .SETB(n118), .RSTB(
        sram_rdata_weight[48]), .CLK(clk), .Q(delay_weight[48]) );
  DFFSSRX1_HVT delay_weight_reg_47_ ( .D(1'b0), .SETB(n114), .RSTB(
        sram_rdata_weight[47]), .CLK(clk), .Q(delay_weight[47]) );
  DFFSSRX1_HVT delay_weight_reg_46_ ( .D(1'b0), .SETB(n109), .RSTB(
        sram_rdata_weight[46]), .CLK(clk), .Q(delay_weight[46]) );
  DFFSSRX1_HVT delay_weight_reg_45_ ( .D(1'b0), .SETB(n119), .RSTB(
        sram_rdata_weight[45]), .CLK(clk), .Q(delay_weight[45]) );
  DFFSSRX1_HVT delay_weight_reg_44_ ( .D(1'b0), .SETB(n115), .RSTB(
        sram_rdata_weight[44]), .CLK(clk), .Q(delay_weight[44]) );
  DFFSSRX1_HVT delay_weight_reg_43_ ( .D(1'b0), .SETB(n110), .RSTB(
        sram_rdata_weight[43]), .CLK(clk), .Q(delay_weight[43]) );
  DFFSSRX1_HVT delay_weight_reg_42_ ( .D(1'b0), .SETB(n116), .RSTB(
        sram_rdata_weight[42]), .CLK(clk), .Q(delay_weight[42]) );
  DFFSSRX1_HVT delay_weight_reg_41_ ( .D(1'b0), .SETB(n112), .RSTB(
        sram_rdata_weight[41]), .CLK(clk), .Q(delay_weight[41]) );
  DFFSSRX1_HVT delay_weight_reg_40_ ( .D(1'b0), .SETB(n107), .RSTB(
        sram_rdata_weight[40]), .CLK(clk), .Q(delay_weight[40]) );
  DFFSSRX1_HVT delay_weight_reg_39_ ( .D(1'b0), .SETB(n117), .RSTB(
        sram_rdata_weight[39]), .CLK(clk), .Q(delay_weight[39]) );
  DFFSSRX1_HVT delay_weight_reg_38_ ( .D(1'b0), .SETB(n113), .RSTB(
        sram_rdata_weight[38]), .CLK(clk), .Q(delay_weight[38]) );
  DFFSSRX1_HVT delay_weight_reg_37_ ( .D(1'b0), .SETB(n108), .RSTB(
        sram_rdata_weight[37]), .CLK(clk), .Q(delay_weight[37]) );
  DFFSSRX1_HVT delay_weight_reg_36_ ( .D(1'b0), .SETB(n118), .RSTB(
        sram_rdata_weight[36]), .CLK(clk), .Q(delay_weight[36]) );
  DFFSSRX1_HVT delay_weight_reg_35_ ( .D(1'b0), .SETB(n114), .RSTB(
        sram_rdata_weight[35]), .CLK(clk), .Q(delay_weight[35]) );
  DFFSSRX1_HVT delay_weight_reg_34_ ( .D(1'b0), .SETB(n109), .RSTB(
        sram_rdata_weight[34]), .CLK(clk), .Q(delay_weight[34]) );
  DFFSSRX1_HVT delay_weight_reg_33_ ( .D(1'b0), .SETB(n119), .RSTB(
        sram_rdata_weight[33]), .CLK(clk), .Q(delay_weight[33]) );
  DFFSSRX1_HVT delay_weight_reg_32_ ( .D(1'b0), .SETB(n115), .RSTB(
        sram_rdata_weight[32]), .CLK(clk), .Q(delay_weight[32]) );
  DFFSSRX1_HVT delay_weight_reg_31_ ( .D(1'b0), .SETB(n110), .RSTB(
        sram_rdata_weight[31]), .CLK(clk), .Q(delay_weight[31]) );
  DFFSSRX1_HVT delay_weight_reg_30_ ( .D(1'b0), .SETB(n116), .RSTB(
        sram_rdata_weight[30]), .CLK(clk), .Q(delay_weight[30]) );
  DFFSSRX1_HVT delay_weight_reg_29_ ( .D(1'b0), .SETB(n112), .RSTB(
        sram_rdata_weight[29]), .CLK(clk), .Q(delay_weight[29]) );
  DFFSSRX1_HVT delay_weight_reg_28_ ( .D(1'b0), .SETB(n107), .RSTB(
        sram_rdata_weight[28]), .CLK(clk), .Q(delay_weight[28]) );
  DFFSSRX1_HVT delay_weight_reg_27_ ( .D(1'b0), .SETB(n117), .RSTB(
        sram_rdata_weight[27]), .CLK(clk), .Q(delay_weight[27]) );
  DFFSSRX1_HVT delay_weight_reg_26_ ( .D(1'b0), .SETB(n113), .RSTB(
        sram_rdata_weight[26]), .CLK(clk), .Q(delay_weight[26]) );
  DFFSSRX1_HVT delay_weight_reg_25_ ( .D(1'b0), .SETB(n108), .RSTB(
        sram_rdata_weight[25]), .CLK(clk), .Q(delay_weight[25]) );
  DFFSSRX1_HVT delay_weight_reg_24_ ( .D(1'b0), .SETB(n118), .RSTB(
        sram_rdata_weight[24]), .CLK(clk), .Q(delay_weight[24]) );
  DFFSSRX1_HVT delay_weight_reg_23_ ( .D(1'b0), .SETB(n114), .RSTB(
        sram_rdata_weight[23]), .CLK(clk), .Q(delay_weight[23]) );
  DFFSSRX1_HVT delay_weight_reg_22_ ( .D(1'b0), .SETB(n109), .RSTB(
        sram_rdata_weight[22]), .CLK(clk), .Q(delay_weight[22]) );
  DFFSSRX1_HVT delay_weight_reg_21_ ( .D(1'b0), .SETB(n119), .RSTB(
        sram_rdata_weight[21]), .CLK(clk), .Q(delay_weight[21]) );
  DFFSSRX1_HVT delay_weight_reg_20_ ( .D(1'b0), .SETB(n115), .RSTB(
        sram_rdata_weight[20]), .CLK(clk), .Q(delay_weight[20]) );
  DFFSSRX1_HVT delay_weight_reg_19_ ( .D(1'b0), .SETB(n110), .RSTB(
        sram_rdata_weight[19]), .CLK(clk), .Q(delay_weight[19]) );
  DFFSSRX1_HVT delay_weight_reg_18_ ( .D(1'b0), .SETB(n116), .RSTB(
        sram_rdata_weight[18]), .CLK(clk), .Q(delay_weight[18]) );
  DFFSSRX1_HVT delay_weight_reg_17_ ( .D(1'b0), .SETB(n112), .RSTB(
        sram_rdata_weight[17]), .CLK(clk), .Q(delay_weight[17]) );
  DFFSSRX1_HVT delay_weight_reg_16_ ( .D(1'b0), .SETB(n107), .RSTB(
        sram_rdata_weight[16]), .CLK(clk), .Q(delay_weight[16]) );
  DFFSSRX1_HVT delay_weight_reg_15_ ( .D(1'b0), .SETB(n117), .RSTB(
        sram_rdata_weight[15]), .CLK(clk), .Q(delay_weight[15]) );
  DFFSSRX1_HVT delay_weight_reg_14_ ( .D(1'b0), .SETB(n113), .RSTB(
        sram_rdata_weight[14]), .CLK(clk), .Q(delay_weight[14]) );
  DFFSSRX1_HVT delay_weight_reg_13_ ( .D(1'b0), .SETB(n108), .RSTB(
        sram_rdata_weight[13]), .CLK(clk), .Q(delay_weight[13]) );
  DFFSSRX1_HVT delay_weight_reg_12_ ( .D(1'b0), .SETB(n118), .RSTB(
        sram_rdata_weight[12]), .CLK(clk), .Q(delay_weight[12]) );
  DFFSSRX1_HVT delay_weight_reg_11_ ( .D(1'b0), .SETB(n114), .RSTB(
        sram_rdata_weight[11]), .CLK(clk), .Q(delay_weight[11]) );
  DFFSSRX1_HVT delay_weight_reg_10_ ( .D(1'b0), .SETB(n109), .RSTB(
        sram_rdata_weight[10]), .CLK(clk), .Q(delay_weight[10]) );
  DFFSSRX1_HVT delay_weight_reg_9_ ( .D(1'b0), .SETB(n119), .RSTB(
        sram_rdata_weight[9]), .CLK(clk), .Q(delay_weight[9]) );
  DFFSSRX1_HVT delay_weight_reg_8_ ( .D(1'b0), .SETB(n115), .RSTB(
        sram_rdata_weight[8]), .CLK(clk), .Q(delay_weight[8]) );
  DFFSSRX1_HVT delay_weight_reg_7_ ( .D(1'b0), .SETB(n110), .RSTB(
        sram_rdata_weight[7]), .CLK(clk), .Q(delay_weight[7]) );
  DFFSSRX1_HVT delay_weight_reg_6_ ( .D(1'b0), .SETB(n116), .RSTB(
        sram_rdata_weight[6]), .CLK(clk), .Q(delay_weight[6]) );
  DFFSSRX1_HVT delay_weight_reg_5_ ( .D(1'b0), .SETB(n112), .RSTB(
        sram_rdata_weight[5]), .CLK(clk), .Q(delay_weight[5]) );
  DFFSSRX1_HVT delay_weight_reg_4_ ( .D(1'b0), .SETB(n107), .RSTB(
        sram_rdata_weight[4]), .CLK(clk), .Q(delay_weight[4]) );
  DFFSSRX1_HVT delay_weight_reg_3_ ( .D(1'b0), .SETB(n117), .RSTB(
        sram_rdata_weight[3]), .CLK(clk), .Q(delay_weight[3]) );
  DFFSSRX1_HVT delay_weight_reg_2_ ( .D(1'b0), .SETB(n113), .RSTB(
        sram_rdata_weight[2]), .CLK(clk), .Q(delay_weight[2]) );
  DFFSSRX1_HVT delay_weight_reg_1_ ( .D(1'b0), .SETB(n108), .RSTB(
        sram_rdata_weight[1]), .CLK(clk), .Q(delay_weight[1]) );
  DFFSSRX1_HVT delay_weight_reg_0_ ( .D(1'b0), .SETB(n118), .RSTB(
        sram_rdata_weight[0]), .CLK(clk), .Q(delay_weight[0]) );
  DFFSSRX1_HVT conv_weight_box_reg_0__3_ ( .D(1'b0), .SETB(n114), .RSTB(
        net22070), .CLK(net22084), .Q(conv_weight_box[199]) );
  DFFSSRX1_HVT conv_weight_box_reg_0__2_ ( .D(1'b0), .SETB(n109), .RSTB(
        net22073), .CLK(net22084), .Q(conv_weight_box[198]) );
  DFFSSRX1_HVT conv_weight_box_reg_0__1_ ( .D(1'b0), .SETB(n119), .RSTB(
        net22074), .CLK(net22084), .Q(conv_weight_box[197]) );
  DFFSSRX1_HVT conv_weight_box_reg_0__0_ ( .D(1'b0), .SETB(n115), .RSTB(
        net22075), .CLK(net22084), .Q(conv_weight_box[196]) );
  DFFSSRX1_HVT conv_weight_box_reg_1__3_ ( .D(1'b0), .SETB(n110), .RSTB(
        net22076), .CLK(net22084), .Q(conv_weight_box[195]) );
  DFFSSRX1_HVT conv_weight_box_reg_1__2_ ( .D(1'b0), .SETB(n116), .RSTB(
        net22077), .CLK(net22084), .Q(conv_weight_box[194]) );
  DFFSSRX1_HVT conv_weight_box_reg_1__1_ ( .D(1'b0), .SETB(n112), .RSTB(
        net22078), .CLK(net22084), .Q(conv_weight_box[193]) );
  DFFSSRX1_HVT conv_weight_box_reg_1__0_ ( .D(1'b0), .SETB(n107), .RSTB(
        net22079), .CLK(net22084), .Q(conv_weight_box[192]) );
  DFFSSRX1_HVT conv_weight_box_reg_2__3_ ( .D(1'b0), .SETB(n117), .RSTB(
        net22080), .CLK(net22084), .Q(conv_weight_box[191]) );
  DFFSSRX1_HVT conv_weight_box_reg_2__2_ ( .D(1'b0), .SETB(n113), .RSTB(
        net22081), .CLK(net22084), .Q(conv_weight_box[190]) );
  DFFSSRX1_HVT conv_weight_box_reg_2__1_ ( .D(1'b0), .SETB(n108), .RSTB(
        net22089), .CLK(net22101), .Q(conv_weight_box[189]) );
  DFFSSRX1_HVT conv_weight_box_reg_2__0_ ( .D(1'b0), .SETB(n118), .RSTB(
        net22090), .CLK(net22101), .Q(conv_weight_box[188]) );
  DFFSSRX1_HVT conv_weight_box_reg_3__3_ ( .D(1'b0), .SETB(n114), .RSTB(
        net22091), .CLK(net22101), .Q(conv_weight_box[187]) );
  DFFSSRX1_HVT conv_weight_box_reg_3__2_ ( .D(1'b0), .SETB(n109), .RSTB(
        net22092), .CLK(net22101), .Q(conv_weight_box[186]) );
  DFFSSRX1_HVT conv_weight_box_reg_3__1_ ( .D(1'b0), .SETB(n119), .RSTB(
        net22093), .CLK(net22101), .Q(conv_weight_box[185]) );
  DFFSSRX1_HVT conv_weight_box_reg_3__0_ ( .D(1'b0), .SETB(n115), .RSTB(
        net22094), .CLK(net22101), .Q(conv_weight_box[184]) );
  DFFSSRX1_HVT conv_weight_box_reg_4__3_ ( .D(1'b0), .SETB(n110), .RSTB(
        net22095), .CLK(net22101), .Q(conv_weight_box[183]) );
  DFFSSRX1_HVT conv_weight_box_reg_4__2_ ( .D(1'b0), .SETB(n116), .RSTB(
        net22096), .CLK(net22101), .Q(conv_weight_box[182]) );
  DFFSSRX1_HVT conv_weight_box_reg_4__1_ ( .D(1'b0), .SETB(n112), .RSTB(
        net22097), .CLK(net22101), .Q(conv_weight_box[181]) );
  DFFSSRX1_HVT conv_weight_box_reg_4__0_ ( .D(1'b0), .SETB(n107), .RSTB(
        net22098), .CLK(net22101), .Q(conv_weight_box[180]) );
  DFFSSRX1_HVT conv_weight_box_reg_5__3_ ( .D(1'b0), .SETB(n117), .RSTB(
        net22106), .CLK(net22118), .Q(conv_weight_box[179]) );
  DFFSSRX1_HVT conv_weight_box_reg_5__2_ ( .D(1'b0), .SETB(n113), .RSTB(
        net22107), .CLK(net22118), .Q(conv_weight_box[178]) );
  DFFSSRX1_HVT conv_weight_box_reg_5__1_ ( .D(1'b0), .SETB(n108), .RSTB(
        net22108), .CLK(net22118), .Q(conv_weight_box[177]) );
  DFFSSRX1_HVT conv_weight_box_reg_5__0_ ( .D(1'b0), .SETB(n118), .RSTB(
        net22109), .CLK(net22118), .Q(conv_weight_box[176]) );
  DFFSSRX1_HVT conv_weight_box_reg_6__3_ ( .D(1'b0), .SETB(n114), .RSTB(
        net22110), .CLK(net22118), .Q(conv_weight_box[175]) );
  DFFSSRX1_HVT conv_weight_box_reg_6__2_ ( .D(1'b0), .SETB(n109), .RSTB(
        net22111), .CLK(net22118), .Q(conv_weight_box[174]) );
  DFFSSRX1_HVT conv_weight_box_reg_6__1_ ( .D(1'b0), .SETB(n119), .RSTB(
        net22112), .CLK(net22118), .Q(conv_weight_box[173]) );
  DFFSSRX1_HVT conv_weight_box_reg_6__0_ ( .D(1'b0), .SETB(n115), .RSTB(
        net22113), .CLK(net22118), .Q(conv_weight_box[172]) );
  DFFSSRX1_HVT conv_weight_box_reg_7__3_ ( .D(1'b0), .SETB(n110), .RSTB(
        net22114), .CLK(net22118), .Q(conv_weight_box[171]) );
  DFFSSRX1_HVT conv_weight_box_reg_7__2_ ( .D(1'b0), .SETB(n116), .RSTB(
        net22115), .CLK(net22118), .Q(conv_weight_box[170]) );
  DFFSSRX1_HVT conv_weight_box_reg_7__1_ ( .D(1'b0), .SETB(n112), .RSTB(
        net22123), .CLK(net22135), .Q(conv_weight_box[169]) );
  DFFSSRX1_HVT conv_weight_box_reg_7__0_ ( .D(1'b0), .SETB(n107), .RSTB(
        net22124), .CLK(net22135), .Q(conv_weight_box[168]) );
  DFFSSRX1_HVT conv_weight_box_reg_8__3_ ( .D(1'b0), .SETB(n117), .RSTB(
        net22125), .CLK(net22135), .Q(conv_weight_box[167]) );
  DFFSSRX1_HVT conv_weight_box_reg_8__2_ ( .D(1'b0), .SETB(n113), .RSTB(
        net22126), .CLK(net22135), .Q(conv_weight_box[166]) );
  DFFSSRX1_HVT conv_weight_box_reg_8__1_ ( .D(1'b0), .SETB(n108), .RSTB(
        net22127), .CLK(net22135), .Q(conv_weight_box[165]) );
  DFFSSRX1_HVT conv_weight_box_reg_8__0_ ( .D(1'b0), .SETB(n118), .RSTB(
        net22128), .CLK(net22135), .Q(conv_weight_box[164]) );
  DFFSSRX1_HVT conv_weight_box_reg_9__3_ ( .D(1'b0), .SETB(n114), .RSTB(
        net22129), .CLK(net22135), .Q(conv_weight_box[163]) );
  DFFSSRX1_HVT conv_weight_box_reg_9__2_ ( .D(1'b0), .SETB(n109), .RSTB(
        net22130), .CLK(net22135), .Q(conv_weight_box[162]) );
  DFFSSRX1_HVT conv_weight_box_reg_9__1_ ( .D(1'b0), .SETB(n119), .RSTB(
        net22131), .CLK(net22135), .Q(conv_weight_box[161]) );
  DFFSSRX1_HVT conv_weight_box_reg_9__0_ ( .D(1'b0), .SETB(n115), .RSTB(
        net22132), .CLK(net22135), .Q(conv_weight_box[160]) );
  DFFSSRX1_HVT conv_weight_box_reg_10__3_ ( .D(1'b0), .SETB(n110), .RSTB(
        net22140), .CLK(net22152), .Q(conv_weight_box[159]) );
  DFFSSRX1_HVT conv_weight_box_reg_10__2_ ( .D(1'b0), .SETB(n116), .RSTB(
        net22141), .CLK(net22152), .Q(conv_weight_box[158]) );
  DFFSSRX1_HVT conv_weight_box_reg_10__1_ ( .D(1'b0), .SETB(n112), .RSTB(
        net22142), .CLK(net22152), .Q(conv_weight_box[157]) );
  DFFSSRX1_HVT conv_weight_box_reg_10__0_ ( .D(1'b0), .SETB(n107), .RSTB(
        net22143), .CLK(net22152), .Q(conv_weight_box[156]) );
  DFFSSRX1_HVT conv_weight_box_reg_11__3_ ( .D(1'b0), .SETB(n117), .RSTB(
        net22144), .CLK(net22152), .Q(conv_weight_box[155]) );
  DFFSSRX1_HVT conv_weight_box_reg_11__2_ ( .D(1'b0), .SETB(n113), .RSTB(
        net22145), .CLK(net22152), .Q(conv_weight_box[154]) );
  DFFSSRX1_HVT conv_weight_box_reg_11__1_ ( .D(1'b0), .SETB(n108), .RSTB(
        net22146), .CLK(net22152), .Q(conv_weight_box[153]) );
  DFFSSRX1_HVT conv_weight_box_reg_11__0_ ( .D(1'b0), .SETB(n118), .RSTB(
        net22147), .CLK(net22152), .Q(conv_weight_box[152]) );
  DFFSSRX1_HVT conv_weight_box_reg_12__3_ ( .D(1'b0), .SETB(n114), .RSTB(
        net22148), .CLK(net22152), .Q(conv_weight_box[151]) );
  DFFSSRX1_HVT conv_weight_box_reg_12__2_ ( .D(1'b0), .SETB(n109), .RSTB(
        net22149), .CLK(net22152), .Q(conv_weight_box[150]) );
  DFFSSRX1_HVT conv_weight_box_reg_12__1_ ( .D(1'b0), .SETB(n119), .RSTB(
        net22157), .CLK(net22169), .Q(conv_weight_box[149]) );
  DFFSSRX1_HVT conv_weight_box_reg_12__0_ ( .D(1'b0), .SETB(n115), .RSTB(
        net22158), .CLK(net22169), .Q(conv_weight_box[148]) );
  DFFSSRX1_HVT conv_weight_box_reg_13__3_ ( .D(1'b0), .SETB(n110), .RSTB(
        net22159), .CLK(net22169), .Q(conv_weight_box[147]) );
  DFFSSRX1_HVT conv_weight_box_reg_13__2_ ( .D(1'b0), .SETB(n116), .RSTB(
        net22160), .CLK(net22169), .Q(conv_weight_box[146]) );
  DFFSSRX1_HVT conv_weight_box_reg_13__1_ ( .D(1'b0), .SETB(n112), .RSTB(
        net22161), .CLK(net22169), .Q(conv_weight_box[145]) );
  DFFSSRX1_HVT conv_weight_box_reg_13__0_ ( .D(1'b0), .SETB(n107), .RSTB(
        net22162), .CLK(net22169), .Q(conv_weight_box[144]) );
  DFFSSRX1_HVT conv_weight_box_reg_14__3_ ( .D(1'b0), .SETB(n117), .RSTB(
        net22163), .CLK(net22169), .Q(conv_weight_box[143]) );
  DFFSSRX1_HVT conv_weight_box_reg_14__2_ ( .D(1'b0), .SETB(n113), .RSTB(
        net22164), .CLK(net22169), .Q(conv_weight_box[142]) );
  DFFSSRX1_HVT conv_weight_box_reg_14__1_ ( .D(1'b0), .SETB(n108), .RSTB(
        net22165), .CLK(net22169), .Q(conv_weight_box[141]) );
  DFFSSRX1_HVT conv_weight_box_reg_14__0_ ( .D(1'b0), .SETB(n118), .RSTB(
        net22166), .CLK(net22169), .Q(conv_weight_box[140]) );
  DFFSSRX1_HVT conv_weight_box_reg_15__3_ ( .D(1'b0), .SETB(n114), .RSTB(
        net22174), .CLK(net22186), .Q(conv_weight_box[139]) );
  DFFSSRX1_HVT conv_weight_box_reg_15__2_ ( .D(1'b0), .SETB(n109), .RSTB(
        net22175), .CLK(net22186), .Q(conv_weight_box[138]) );
  DFFSSRX1_HVT conv_weight_box_reg_15__1_ ( .D(1'b0), .SETB(n119), .RSTB(
        net22176), .CLK(net22186), .Q(conv_weight_box[137]) );
  DFFSSRX1_HVT conv_weight_box_reg_15__0_ ( .D(1'b0), .SETB(n115), .RSTB(
        net22177), .CLK(net22186), .Q(conv_weight_box[136]) );
  DFFSSRX1_HVT conv_weight_box_reg_16__3_ ( .D(1'b0), .SETB(n110), .RSTB(
        net22178), .CLK(net22186), .Q(conv_weight_box[135]) );
  DFFSSRX1_HVT conv_weight_box_reg_16__2_ ( .D(1'b0), .SETB(n116), .RSTB(
        net22179), .CLK(net22186), .Q(conv_weight_box[134]) );
  DFFSSRX1_HVT conv_weight_box_reg_16__1_ ( .D(1'b0), .SETB(n112), .RSTB(
        net22180), .CLK(net22186), .Q(conv_weight_box[133]) );
  DFFSSRX1_HVT conv_weight_box_reg_16__0_ ( .D(1'b0), .SETB(n107), .RSTB(
        net22181), .CLK(net22186), .Q(conv_weight_box[132]) );
  DFFSSRX1_HVT conv_weight_box_reg_17__3_ ( .D(1'b0), .SETB(n117), .RSTB(
        net22182), .CLK(net22186), .Q(conv_weight_box[131]) );
  DFFSSRX1_HVT conv_weight_box_reg_17__2_ ( .D(1'b0), .SETB(n113), .RSTB(
        net22183), .CLK(net22186), .Q(conv_weight_box[130]) );
  DFFSSRX1_HVT conv_weight_box_reg_17__1_ ( .D(1'b0), .SETB(n108), .RSTB(
        net22191), .CLK(net22203), .Q(conv_weight_box[129]) );
  DFFSSRX1_HVT conv_weight_box_reg_17__0_ ( .D(1'b0), .SETB(n118), .RSTB(
        net22192), .CLK(net22203), .Q(conv_weight_box[128]) );
  DFFSSRX1_HVT conv_weight_box_reg_18__3_ ( .D(1'b0), .SETB(n114), .RSTB(
        net22193), .CLK(net22203), .Q(conv_weight_box[127]) );
  DFFSSRX1_HVT conv_weight_box_reg_18__2_ ( .D(1'b0), .SETB(n109), .RSTB(
        net22194), .CLK(net22203), .Q(conv_weight_box[126]) );
  DFFSSRX1_HVT conv_weight_box_reg_18__1_ ( .D(1'b0), .SETB(n119), .RSTB(
        net22195), .CLK(net22203), .Q(conv_weight_box[125]) );
  DFFSSRX1_HVT conv_weight_box_reg_18__0_ ( .D(1'b0), .SETB(n115), .RSTB(
        net22196), .CLK(net22203), .Q(conv_weight_box[124]) );
  DFFSSRX1_HVT conv_weight_box_reg_19__3_ ( .D(1'b0), .SETB(n110), .RSTB(
        net22197), .CLK(net22203), .Q(conv_weight_box[123]) );
  DFFSSRX1_HVT conv_weight_box_reg_19__2_ ( .D(1'b0), .SETB(n116), .RSTB(
        net22198), .CLK(net22203), .Q(conv_weight_box[122]) );
  DFFSSRX1_HVT conv_weight_box_reg_19__1_ ( .D(1'b0), .SETB(n112), .RSTB(
        net22199), .CLK(net22203), .Q(conv_weight_box[121]) );
  DFFSSRX1_HVT conv_weight_box_reg_19__0_ ( .D(1'b0), .SETB(n107), .RSTB(
        net22200), .CLK(net22203), .Q(conv_weight_box[120]) );
  DFFSSRX1_HVT conv_weight_box_reg_20__3_ ( .D(1'b0), .SETB(n117), .RSTB(
        net22208), .CLK(net22220), .Q(conv_weight_box[119]) );
  DFFSSRX1_HVT conv_weight_box_reg_20__2_ ( .D(1'b0), .SETB(n113), .RSTB(
        net22209), .CLK(net22220), .Q(conv_weight_box[118]) );
  DFFSSRX1_HVT conv_weight_box_reg_20__1_ ( .D(1'b0), .SETB(n108), .RSTB(
        net22210), .CLK(net22220), .Q(conv_weight_box[117]) );
  DFFSSRX1_HVT conv_weight_box_reg_20__0_ ( .D(1'b0), .SETB(n118), .RSTB(
        net22211), .CLK(net22220), .Q(conv_weight_box[116]) );
  DFFSSRX1_HVT conv_weight_box_reg_21__3_ ( .D(1'b0), .SETB(n114), .RSTB(
        net22212), .CLK(net22220), .Q(conv_weight_box[115]) );
  DFFSSRX1_HVT conv_weight_box_reg_21__2_ ( .D(1'b0), .SETB(n109), .RSTB(
        net22213), .CLK(net22220), .Q(conv_weight_box[114]) );
  DFFSSRX1_HVT conv_weight_box_reg_21__1_ ( .D(1'b0), .SETB(n119), .RSTB(
        net22214), .CLK(net22220), .Q(conv_weight_box[113]) );
  DFFSSRX1_HVT conv_weight_box_reg_21__0_ ( .D(1'b0), .SETB(n115), .RSTB(
        net22215), .CLK(net22220), .Q(conv_weight_box[112]) );
  DFFSSRX1_HVT conv_weight_box_reg_22__3_ ( .D(1'b0), .SETB(n110), .RSTB(
        net22216), .CLK(net22220), .Q(conv_weight_box[111]) );
  DFFSSRX1_HVT conv_weight_box_reg_22__2_ ( .D(1'b0), .SETB(n116), .RSTB(
        net22217), .CLK(net22220), .Q(conv_weight_box[110]) );
  DFFSSRX1_HVT conv_weight_box_reg_22__1_ ( .D(1'b0), .SETB(n112), .RSTB(
        net22225), .CLK(net22237), .Q(conv_weight_box[109]) );
  DFFSSRX1_HVT conv_weight_box_reg_22__0_ ( .D(1'b0), .SETB(n107), .RSTB(
        net22226), .CLK(net22237), .Q(conv_weight_box[108]) );
  DFFSSRX1_HVT conv_weight_box_reg_23__3_ ( .D(1'b0), .SETB(n117), .RSTB(
        net22227), .CLK(net22237), .Q(conv_weight_box[107]) );
  DFFSSRX1_HVT conv_weight_box_reg_23__2_ ( .D(1'b0), .SETB(n113), .RSTB(
        net22228), .CLK(net22237), .Q(conv_weight_box[106]) );
  DFFSSRX1_HVT conv_weight_box_reg_23__1_ ( .D(1'b0), .SETB(n108), .RSTB(
        net22229), .CLK(net22237), .Q(conv_weight_box[105]) );
  DFFSSRX1_HVT conv_weight_box_reg_23__0_ ( .D(1'b0), .SETB(n118), .RSTB(
        net22230), .CLK(net22237), .Q(conv_weight_box[104]) );
  DFFSSRX1_HVT conv_weight_box_reg_24__3_ ( .D(1'b0), .SETB(n114), .RSTB(
        net22231), .CLK(net22237), .Q(conv_weight_box[103]) );
  DFFSSRX1_HVT conv_weight_box_reg_24__2_ ( .D(1'b0), .SETB(n109), .RSTB(
        net22232), .CLK(net22237), .Q(conv_weight_box[102]) );
  DFFSSRX1_HVT conv_weight_box_reg_24__1_ ( .D(1'b0), .SETB(n119), .RSTB(
        net22233), .CLK(net22237), .Q(conv_weight_box[101]) );
  DFFSSRX1_HVT conv_weight_box_reg_24__0_ ( .D(1'b0), .SETB(n115), .RSTB(
        net22234), .CLK(net22237), .Q(conv_weight_box[100]) );
  DFFSSRX1_HVT conv_weight_box_reg_25__3_ ( .D(1'b0), .SETB(n110), .RSTB(
        net22250), .CLK(net22262), .Q(conv_weight_box[99]) );
  DFFSSRX1_HVT conv_weight_box_reg_25__2_ ( .D(1'b0), .SETB(n116), .RSTB(
        net22251), .CLK(net22262), .Q(conv_weight_box[98]) );
  DFFSSRX1_HVT conv_weight_box_reg_25__1_ ( .D(1'b0), .SETB(n112), .RSTB(
        net22252), .CLK(net22262), .Q(conv_weight_box[97]) );
  DFFSSRX1_HVT conv_weight_box_reg_25__0_ ( .D(1'b0), .SETB(n107), .RSTB(
        net22253), .CLK(net22262), .Q(conv_weight_box[96]) );
  DFFSSRX1_HVT conv_weight_box_reg_26__3_ ( .D(1'b0), .SETB(n117), .RSTB(
        net22254), .CLK(net22262), .Q(conv_weight_box[95]) );
  DFFSSRX1_HVT conv_weight_box_reg_26__2_ ( .D(1'b0), .SETB(n113), .RSTB(
        net22255), .CLK(net22262), .Q(conv_weight_box[94]) );
  DFFSSRX1_HVT conv_weight_box_reg_26__1_ ( .D(1'b0), .SETB(n108), .RSTB(
        net22256), .CLK(net22262), .Q(conv_weight_box[93]) );
  DFFSSRX1_HVT conv_weight_box_reg_26__0_ ( .D(1'b0), .SETB(n118), .RSTB(
        net22257), .CLK(net22262), .Q(conv_weight_box[92]) );
  DFFSSRX1_HVT conv_weight_box_reg_27__3_ ( .D(1'b0), .SETB(n114), .RSTB(
        net22258), .CLK(net22262), .Q(conv_weight_box[91]) );
  DFFSSRX1_HVT conv_weight_box_reg_27__2_ ( .D(1'b0), .SETB(n109), .RSTB(
        net22259), .CLK(net22262), .Q(conv_weight_box[90]) );
  DFFSSRX1_HVT conv_weight_box_reg_27__1_ ( .D(1'b0), .SETB(n119), .RSTB(
        net22267), .CLK(net22279), .Q(conv_weight_box[89]) );
  DFFSSRX1_HVT conv_weight_box_reg_27__0_ ( .D(1'b0), .SETB(n115), .RSTB(
        net22268), .CLK(net22279), .Q(conv_weight_box[88]) );
  DFFSSRX1_HVT conv_weight_box_reg_28__3_ ( .D(1'b0), .SETB(n110), .RSTB(
        net22269), .CLK(net22279), .Q(conv_weight_box[87]) );
  DFFSSRX1_HVT conv_weight_box_reg_28__2_ ( .D(1'b0), .SETB(n116), .RSTB(
        net22270), .CLK(net22279), .Q(conv_weight_box[86]) );
  DFFSSRX1_HVT conv_weight_box_reg_28__1_ ( .D(1'b0), .SETB(n112), .RSTB(
        net22271), .CLK(net22279), .Q(conv_weight_box[85]) );
  DFFSSRX1_HVT conv_weight_box_reg_28__0_ ( .D(1'b0), .SETB(n107), .RSTB(
        net22272), .CLK(net22279), .Q(conv_weight_box[84]) );
  DFFSSRX1_HVT conv_weight_box_reg_29__3_ ( .D(1'b0), .SETB(n117), .RSTB(
        net22273), .CLK(net22279), .Q(conv_weight_box[83]) );
  DFFSSRX1_HVT conv_weight_box_reg_29__2_ ( .D(1'b0), .SETB(n113), .RSTB(
        net22274), .CLK(net22279), .Q(conv_weight_box[82]) );
  DFFSSRX1_HVT conv_weight_box_reg_29__1_ ( .D(1'b0), .SETB(n108), .RSTB(
        net22275), .CLK(net22279), .Q(conv_weight_box[81]) );
  DFFSSRX1_HVT conv_weight_box_reg_29__0_ ( .D(1'b0), .SETB(n118), .RSTB(
        net22276), .CLK(net22279), .Q(conv_weight_box[80]) );
  DFFSSRX1_HVT conv_weight_box_reg_30__3_ ( .D(1'b0), .SETB(n114), .RSTB(
        net22284), .CLK(net22296), .Q(conv_weight_box[79]) );
  DFFSSRX1_HVT conv_weight_box_reg_30__2_ ( .D(1'b0), .SETB(n109), .RSTB(
        net22285), .CLK(net22296), .Q(conv_weight_box[78]) );
  DFFSSRX1_HVT conv_weight_box_reg_30__1_ ( .D(1'b0), .SETB(n119), .RSTB(
        net22286), .CLK(net22296), .Q(conv_weight_box[77]) );
  DFFSSRX1_HVT conv_weight_box_reg_30__0_ ( .D(1'b0), .SETB(n115), .RSTB(
        net22287), .CLK(net22296), .Q(conv_weight_box[76]) );
  DFFSSRX1_HVT conv_weight_box_reg_31__3_ ( .D(1'b0), .SETB(n110), .RSTB(
        net22288), .CLK(net22296), .Q(conv_weight_box[75]) );
  DFFSSRX1_HVT conv_weight_box_reg_31__2_ ( .D(1'b0), .SETB(n116), .RSTB(
        net22289), .CLK(net22296), .Q(conv_weight_box[74]) );
  DFFSSRX1_HVT conv_weight_box_reg_31__1_ ( .D(1'b0), .SETB(n112), .RSTB(
        net22290), .CLK(net22296), .Q(conv_weight_box[73]) );
  DFFSSRX1_HVT conv_weight_box_reg_31__0_ ( .D(1'b0), .SETB(n107), .RSTB(
        net22291), .CLK(net22296), .Q(conv_weight_box[72]) );
  DFFSSRX1_HVT conv_weight_box_reg_32__3_ ( .D(1'b0), .SETB(n117), .RSTB(
        net22292), .CLK(net22296), .Q(conv_weight_box[71]) );
  DFFSSRX1_HVT conv_weight_box_reg_32__2_ ( .D(1'b0), .SETB(n113), .RSTB(
        net22293), .CLK(net22296), .Q(conv_weight_box[70]) );
  DFFSSRX1_HVT conv_weight_box_reg_32__1_ ( .D(1'b0), .SETB(n108), .RSTB(
        net22301), .CLK(net22313), .Q(conv_weight_box[69]) );
  DFFSSRX1_HVT conv_weight_box_reg_32__0_ ( .D(1'b0), .SETB(n118), .RSTB(
        net22302), .CLK(net22313), .Q(conv_weight_box[68]) );
  DFFSSRX1_HVT conv_weight_box_reg_33__3_ ( .D(1'b0), .SETB(n114), .RSTB(
        net22303), .CLK(net22313), .Q(conv_weight_box[67]) );
  DFFSSRX1_HVT conv_weight_box_reg_33__2_ ( .D(1'b0), .SETB(n109), .RSTB(
        net22304), .CLK(net22313), .Q(conv_weight_box[66]) );
  DFFSSRX1_HVT conv_weight_box_reg_33__1_ ( .D(1'b0), .SETB(n119), .RSTB(
        net22305), .CLK(net22313), .Q(conv_weight_box[65]) );
  DFFSSRX1_HVT conv_weight_box_reg_33__0_ ( .D(1'b0), .SETB(n115), .RSTB(
        net22306), .CLK(net22313), .Q(conv_weight_box[64]) );
  DFFSSRX1_HVT conv_weight_box_reg_34__3_ ( .D(1'b0), .SETB(n110), .RSTB(
        net22307), .CLK(net22313), .Q(conv_weight_box[63]) );
  DFFSSRX1_HVT conv_weight_box_reg_34__2_ ( .D(1'b0), .SETB(n116), .RSTB(
        net22308), .CLK(net22313), .Q(conv_weight_box[62]) );
  DFFSSRX1_HVT conv_weight_box_reg_34__1_ ( .D(1'b0), .SETB(n112), .RSTB(
        net22309), .CLK(net22313), .Q(conv_weight_box[61]) );
  DFFSSRX1_HVT conv_weight_box_reg_34__0_ ( .D(1'b0), .SETB(n107), .RSTB(
        net22310), .CLK(net22313), .Q(conv_weight_box[60]) );
  DFFSSRX1_HVT conv_weight_box_reg_35__3_ ( .D(1'b0), .SETB(n117), .RSTB(
        net22318), .CLK(net22330), .Q(conv_weight_box[59]) );
  DFFSSRX1_HVT conv_weight_box_reg_35__2_ ( .D(1'b0), .SETB(n113), .RSTB(
        net22319), .CLK(net22330), .Q(conv_weight_box[58]) );
  DFFSSRX1_HVT conv_weight_box_reg_35__1_ ( .D(1'b0), .SETB(n108), .RSTB(
        net22320), .CLK(net22330), .Q(conv_weight_box[57]) );
  DFFSSRX1_HVT conv_weight_box_reg_35__0_ ( .D(1'b0), .SETB(n118), .RSTB(
        net22321), .CLK(net22330), .Q(conv_weight_box[56]) );
  DFFSSRX1_HVT conv_weight_box_reg_36__3_ ( .D(1'b0), .SETB(n114), .RSTB(
        net22322), .CLK(net22330), .Q(conv_weight_box[55]) );
  DFFSSRX1_HVT conv_weight_box_reg_36__2_ ( .D(1'b0), .SETB(n109), .RSTB(
        net22323), .CLK(net22330), .Q(conv_weight_box[54]) );
  DFFSSRX1_HVT conv_weight_box_reg_36__1_ ( .D(1'b0), .SETB(n119), .RSTB(
        net22324), .CLK(net22330), .Q(conv_weight_box[53]) );
  DFFSSRX1_HVT conv_weight_box_reg_36__0_ ( .D(1'b0), .SETB(n115), .RSTB(
        net22325), .CLK(net22330), .Q(conv_weight_box[52]) );
  DFFSSRX1_HVT conv_weight_box_reg_37__3_ ( .D(1'b0), .SETB(n110), .RSTB(
        net22326), .CLK(net22330), .Q(conv_weight_box[51]) );
  DFFSSRX1_HVT conv_weight_box_reg_37__2_ ( .D(1'b0), .SETB(n116), .RSTB(
        net22327), .CLK(net22330), .Q(conv_weight_box[50]) );
  DFFSSRX1_HVT conv_weight_box_reg_37__1_ ( .D(1'b0), .SETB(n112), .RSTB(
        net22335), .CLK(net22347), .Q(conv_weight_box[49]) );
  DFFSSRX1_HVT conv_weight_box_reg_37__0_ ( .D(1'b0), .SETB(n107), .RSTB(
        net22336), .CLK(net22347), .Q(conv_weight_box[48]) );
  DFFSSRX1_HVT conv_weight_box_reg_38__3_ ( .D(1'b0), .SETB(n117), .RSTB(
        net22337), .CLK(net22347), .Q(conv_weight_box[47]) );
  DFFSSRX1_HVT conv_weight_box_reg_38__2_ ( .D(1'b0), .SETB(n113), .RSTB(
        net22338), .CLK(net22347), .Q(conv_weight_box[46]) );
  DFFSSRX1_HVT conv_weight_box_reg_38__1_ ( .D(1'b0), .SETB(n108), .RSTB(
        net22339), .CLK(net22347), .Q(conv_weight_box[45]) );
  DFFSSRX1_HVT conv_weight_box_reg_38__0_ ( .D(1'b0), .SETB(n118), .RSTB(
        net22340), .CLK(net22347), .Q(conv_weight_box[44]) );
  DFFSSRX1_HVT conv_weight_box_reg_39__3_ ( .D(1'b0), .SETB(n114), .RSTB(
        net22341), .CLK(net22347), .Q(conv_weight_box[43]) );
  DFFSSRX1_HVT conv_weight_box_reg_39__2_ ( .D(1'b0), .SETB(n109), .RSTB(
        net22342), .CLK(net22347), .Q(conv_weight_box[42]) );
  DFFSSRX1_HVT conv_weight_box_reg_39__1_ ( .D(1'b0), .SETB(n119), .RSTB(
        net22343), .CLK(net22347), .Q(conv_weight_box[41]) );
  DFFSSRX1_HVT conv_weight_box_reg_39__0_ ( .D(1'b0), .SETB(n115), .RSTB(
        net22344), .CLK(net22347), .Q(conv_weight_box[40]) );
  DFFSSRX1_HVT conv_weight_box_reg_40__3_ ( .D(1'b0), .SETB(n110), .RSTB(
        net22352), .CLK(net22364), .Q(conv_weight_box[39]) );
  DFFSSRX1_HVT conv_weight_box_reg_40__2_ ( .D(1'b0), .SETB(n116), .RSTB(
        net22353), .CLK(net22364), .Q(conv_weight_box[38]) );
  DFFSSRX1_HVT conv_weight_box_reg_40__1_ ( .D(1'b0), .SETB(n112), .RSTB(
        net22354), .CLK(net22364), .Q(conv_weight_box[37]) );
  DFFSSRX1_HVT conv_weight_box_reg_40__0_ ( .D(1'b0), .SETB(n107), .RSTB(
        net22355), .CLK(net22364), .Q(conv_weight_box[36]) );
  DFFSSRX1_HVT conv_weight_box_reg_41__3_ ( .D(1'b0), .SETB(n117), .RSTB(
        net22356), .CLK(net22364), .Q(conv_weight_box[35]) );
  DFFSSRX1_HVT conv_weight_box_reg_41__2_ ( .D(1'b0), .SETB(n113), .RSTB(
        net22357), .CLK(net22364), .Q(conv_weight_box[34]) );
  DFFSSRX1_HVT conv_weight_box_reg_41__1_ ( .D(1'b0), .SETB(n108), .RSTB(
        net22358), .CLK(net22364), .Q(conv_weight_box[33]) );
  DFFSSRX1_HVT conv_weight_box_reg_41__0_ ( .D(1'b0), .SETB(n118), .RSTB(
        net22359), .CLK(net22364), .Q(conv_weight_box[32]) );
  DFFSSRX1_HVT conv_weight_box_reg_42__3_ ( .D(1'b0), .SETB(n114), .RSTB(
        net22360), .CLK(net22364), .Q(conv_weight_box[31]) );
  DFFSSRX1_HVT conv_weight_box_reg_42__2_ ( .D(1'b0), .SETB(n109), .RSTB(
        net22361), .CLK(net22364), .Q(conv_weight_box[30]) );
  DFFSSRX1_HVT conv_weight_box_reg_42__1_ ( .D(1'b0), .SETB(n119), .RSTB(
        net22369), .CLK(net22381), .Q(conv_weight_box[29]) );
  DFFSSRX1_HVT conv_weight_box_reg_42__0_ ( .D(1'b0), .SETB(n115), .RSTB(
        net22370), .CLK(net22381), .Q(conv_weight_box[28]) );
  DFFSSRX1_HVT conv_weight_box_reg_43__3_ ( .D(1'b0), .SETB(n110), .RSTB(
        net22371), .CLK(net22381), .Q(conv_weight_box[27]) );
  DFFSSRX1_HVT conv_weight_box_reg_43__2_ ( .D(1'b0), .SETB(n116), .RSTB(
        net22372), .CLK(net22381), .Q(conv_weight_box[26]) );
  DFFSSRX1_HVT conv_weight_box_reg_43__1_ ( .D(1'b0), .SETB(n112), .RSTB(
        net22373), .CLK(net22381), .Q(conv_weight_box[25]) );
  DFFSSRX1_HVT conv_weight_box_reg_43__0_ ( .D(1'b0), .SETB(n107), .RSTB(
        net22374), .CLK(net22381), .Q(conv_weight_box[24]) );
  DFFSSRX1_HVT conv_weight_box_reg_44__3_ ( .D(1'b0), .SETB(n117), .RSTB(
        net22375), .CLK(net22381), .Q(conv_weight_box[23]) );
  DFFSSRX1_HVT conv_weight_box_reg_44__2_ ( .D(1'b0), .SETB(n113), .RSTB(
        net22376), .CLK(net22381), .Q(conv_weight_box[22]) );
  DFFSSRX1_HVT conv_weight_box_reg_44__1_ ( .D(1'b0), .SETB(n108), .RSTB(
        net22377), .CLK(net22381), .Q(conv_weight_box[21]) );
  DFFSSRX1_HVT conv_weight_box_reg_44__0_ ( .D(1'b0), .SETB(n118), .RSTB(
        net22378), .CLK(net22381), .Q(conv_weight_box[20]) );
  DFFSSRX1_HVT conv_weight_box_reg_45__3_ ( .D(1'b0), .SETB(n114), .RSTB(
        net22386), .CLK(net22398), .Q(conv_weight_box[19]) );
  DFFSSRX1_HVT conv_weight_box_reg_45__2_ ( .D(1'b0), .SETB(n109), .RSTB(
        net22387), .CLK(net22398), .Q(conv_weight_box[18]) );
  DFFSSRX1_HVT conv_weight_box_reg_45__1_ ( .D(1'b0), .SETB(n119), .RSTB(
        net22388), .CLK(net22398), .Q(conv_weight_box[17]) );
  DFFSSRX1_HVT conv_weight_box_reg_45__0_ ( .D(1'b0), .SETB(n115), .RSTB(
        net22389), .CLK(net22398), .Q(conv_weight_box[16]) );
  DFFSSRX1_HVT conv_weight_box_reg_46__3_ ( .D(1'b0), .SETB(n110), .RSTB(
        net22390), .CLK(net22398), .Q(conv_weight_box[15]) );
  DFFSSRX1_HVT conv_weight_box_reg_46__2_ ( .D(1'b0), .SETB(n116), .RSTB(
        net22391), .CLK(net22398), .Q(conv_weight_box[14]) );
  DFFSSRX1_HVT conv_weight_box_reg_46__1_ ( .D(1'b0), .SETB(n112), .RSTB(
        net22392), .CLK(net22398), .Q(conv_weight_box[13]) );
  DFFSSRX1_HVT conv_weight_box_reg_46__0_ ( .D(1'b0), .SETB(n107), .RSTB(
        net22393), .CLK(net22398), .Q(conv_weight_box[12]) );
  DFFSSRX1_HVT conv_weight_box_reg_47__3_ ( .D(1'b0), .SETB(n117), .RSTB(
        net22394), .CLK(net22398), .Q(conv_weight_box[11]) );
  DFFSSRX1_HVT conv_weight_box_reg_47__2_ ( .D(1'b0), .SETB(n113), .RSTB(
        net22395), .CLK(net22398), .Q(conv_weight_box[10]) );
  DFFSSRX1_HVT conv_weight_box_reg_47__1_ ( .D(1'b0), .SETB(n108), .RSTB(
        net22403), .CLK(net22415), .Q(conv_weight_box[9]) );
  DFFSSRX1_HVT conv_weight_box_reg_47__0_ ( .D(1'b0), .SETB(n118), .RSTB(
        net22404), .CLK(net22415), .Q(conv_weight_box[8]) );
  DFFSSRX1_HVT conv_weight_box_reg_48__3_ ( .D(1'b0), .SETB(n114), .RSTB(
        net22405), .CLK(net22415), .Q(conv_weight_box[7]) );
  DFFSSRX1_HVT conv_weight_box_reg_48__2_ ( .D(1'b0), .SETB(n109), .RSTB(
        net22406), .CLK(net22415), .Q(conv_weight_box[6]) );
  DFFSSRX1_HVT conv_weight_box_reg_48__1_ ( .D(1'b0), .SETB(n119), .RSTB(
        net22407), .CLK(net22415), .Q(conv_weight_box[5]) );
  DFFSSRX1_HVT conv_weight_box_reg_48__0_ ( .D(1'b0), .SETB(n115), .RSTB(
        net22408), .CLK(net22415), .Q(conv_weight_box[4]) );
  DFFSSRX1_HVT conv_weight_box_reg_49__3_ ( .D(1'b0), .SETB(n110), .RSTB(
        net22409), .CLK(net22415), .Q(conv_weight_box[3]) );
  DFFSSRX1_HVT conv_weight_box_reg_49__2_ ( .D(1'b0), .SETB(n116), .RSTB(
        net22410), .CLK(net22415), .Q(conv_weight_box[2]) );
  DFFSSRX1_HVT conv_weight_box_reg_49__1_ ( .D(1'b0), .SETB(n112), .RSTB(
        net22411), .CLK(net22415), .Q(conv_weight_box[1]) );
  DFFSSRX1_HVT conv_weight_box_reg_49__0_ ( .D(1'b0), .SETB(n107), .RSTB(
        net22412), .CLK(net22415), .Q(conv_weight_box[0]) );
  DFFSSRX1_HVT bias_data_reg_3_ ( .D(1'b0), .SETB(n117), .RSTB(net22432), 
        .CLK(net22447), .Q(bias_data[3]) );
  DFFSSRX1_HVT bias_data_reg_2_ ( .D(1'b0), .SETB(n113), .RSTB(net22436), 
        .CLK(net22447), .Q(bias_data[2]) );
  DFFSSRX1_HVT bias_data_reg_1_ ( .D(1'b0), .SETB(n108), .RSTB(net22440), 
        .CLK(net22447), .Q(bias_data[1]) );
  DFFSSRX1_HVT bias_data_reg_0_ ( .D(1'b0), .SETB(n118), .RSTB(net22444), 
        .CLK(net22447), .Q(bias_data[0]) );
  OR2X1_HVT U3 ( .A1(n135), .A2(mode[0]), .Y(n158) );
  AO22X1_HVT U4 ( .A1(n137), .A2(load_conv2_bias0_enable), .A3(mode[0]), .A4(
        n135), .Y(n136) );
  NOR3X0_HVT U5 ( .A1(n158), .A2(load_conv2_bias1_enable), .A3(
        load_conv2_bias0_enable), .Y(n129) );
  AO22X1_HVT U6 ( .A1(conv_weight_box[10]), .A2(n288), .A3(conv_weight_box[14]), .A4(n289), .Y(n1) );
  AO22X1_HVT U7 ( .A1(conv_weight_box[86]), .A2(n290), .A3(conv_weight_box[82]), .A4(n291), .Y(n2) );
  AO22X1_HVT U8 ( .A1(conv_weight_box[22]), .A2(n292), .A3(conv_weight_box[74]), .A4(n293), .Y(n3) );
  AO22X1_HVT U9 ( .A1(conv_weight_box[70]), .A2(n294), .A3(conv_weight_box[66]), .A4(n295), .Y(n4) );
  NOR4X0_HVT U10 ( .A1(n1), .A2(n2), .A3(n3), .A4(n4), .Y(n5) );
  AO22X1_HVT U11 ( .A1(n326), .A2(conv_weight_box[98]), .A3(n324), .A4(
        conv_weight_box[114]), .Y(n6) );
  AO22X1_HVT U12 ( .A1(n320), .A2(conv_weight_box[34]), .A3(n318), .A4(
        conv_weight_box[50]), .Y(n7) );
  AO22X1_HVT U13 ( .A1(n319), .A2(conv_weight_box[194]), .A3(n317), .A4(
        conv_weight_box[178]), .Y(n8) );
  AO22X1_HVT U14 ( .A1(n322), .A2(conv_weight_box[146]), .A3(n321), .A4(
        conv_weight_box[162]), .Y(n9) );
  NOR4X0_HVT U15 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .Y(n10) );
  AO22X1_HVT U16 ( .A1(n320), .A2(conv_weight_box[38]), .A3(n318), .A4(
        conv_weight_box[54]), .Y(n11) );
  NOR4X0_HVT U17 ( .A1(n186), .A2(n187), .A3(n185), .A4(n11), .Y(n12) );
  OA22X1_HVT U18 ( .A1(n10), .A2(n284), .A3(n12), .A4(n286), .Y(n13) );
  AO22X1_HVT U19 ( .A1(conv_weight_box[78]), .A2(n306), .A3(
        conv_weight_box[130]), .A4(n307), .Y(n14) );
  AO22X1_HVT U20 ( .A1(conv_weight_box[134]), .A2(n300), .A3(
        conv_weight_box[18]), .A4(n301), .Y(n15) );
  AO22X1_HVT U21 ( .A1(conv_weight_box[6]), .A2(n302), .A3(conv_weight_box[2]), 
        .A4(n303), .Y(n16) );
  OR3X1_HVT U22 ( .A1(n193), .A2(n192), .A3(n191), .Y(n17) );
  OR3X1_HVT U23 ( .A1(n199), .A2(n198), .A3(n197), .Y(n18) );
  AO22X1_HVT U24 ( .A1(n336), .A2(n17), .A3(n334), .A4(n18), .Y(n19) );
  NOR4X0_HVT U25 ( .A1(n14), .A2(n15), .A3(n16), .A4(n19), .Y(n20) );
  NAND3X0_HVT U26 ( .A1(n5), .A2(n13), .A3(n20), .Y(n21) );
  AO22X1_HVT U27 ( .A1(conv_weight_box[10]), .A2(n353), .A3(
        conv_weight_box[14]), .A4(n354), .Y(n22) );
  AO22X1_HVT U28 ( .A1(conv_weight_box[86]), .A2(n355), .A3(
        conv_weight_box[82]), .A4(n356), .Y(n23) );
  AO22X1_HVT U29 ( .A1(conv_weight_box[22]), .A2(n357), .A3(
        conv_weight_box[74]), .A4(n358), .Y(n24) );
  AO22X1_HVT U30 ( .A1(conv_weight_box[70]), .A2(n359), .A3(
        conv_weight_box[66]), .A4(n360), .Y(n25) );
  NOR4X0_HVT U31 ( .A1(n22), .A2(n23), .A3(n24), .A4(n25), .Y(n26) );
  AO22X1_HVT U32 ( .A1(n389), .A2(conv_weight_box[98]), .A3(n387), .A4(
        conv_weight_box[114]), .Y(n27) );
  AO22X1_HVT U33 ( .A1(conv_weight_box[34]), .A2(n383), .A3(
        conv_weight_box[50]), .A4(n381), .Y(n28) );
  AO22X1_HVT U34 ( .A1(conv_weight_box[194]), .A2(n382), .A3(
        conv_weight_box[178]), .A4(n380), .Y(n29) );
  AO22X1_HVT U35 ( .A1(n385), .A2(conv_weight_box[146]), .A3(n384), .A4(
        conv_weight_box[162]), .Y(n30) );
  NOR4X0_HVT U36 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .Y(n31) );
  AO22X1_HVT U37 ( .A1(n389), .A2(conv_weight_box[102]), .A3(n387), .A4(
        conv_weight_box[118]), .Y(n32) );
  AO22X1_HVT U38 ( .A1(n383), .A2(conv_weight_box[38]), .A3(n381), .A4(
        conv_weight_box[54]), .Y(n33) );
  AO22X1_HVT U39 ( .A1(conv_weight_box[182]), .A2(n380), .A3(
        conv_weight_box[198]), .A4(n382), .Y(n34) );
  AO22X1_HVT U40 ( .A1(n385), .A2(conv_weight_box[150]), .A3(n384), .A4(
        conv_weight_box[166]), .Y(n35) );
  NOR4X0_HVT U41 ( .A1(n32), .A2(n33), .A3(n34), .A4(n35), .Y(n36) );
  OA22X1_HVT U42 ( .A1(n31), .A2(n349), .A3(n36), .A4(n351), .Y(n37) );
  AO22X1_HVT U43 ( .A1(conv_weight_box[78]), .A2(n369), .A3(
        conv_weight_box[130]), .A4(n370), .Y(n38) );
  AO22X1_HVT U44 ( .A1(conv_weight_box[134]), .A2(n365), .A3(
        conv_weight_box[18]), .A4(n366), .Y(n39) );
  AO22X1_HVT U45 ( .A1(conv_weight_box[6]), .A2(n367), .A3(conv_weight_box[2]), 
        .A4(n368), .Y(n40) );
  OR3X1_HVT U46 ( .A1(n202), .A2(n201), .A3(n200), .Y(n41) );
  AO22X1_HVT U47 ( .A1(conv_weight_box[30]), .A2(n383), .A3(
        conv_weight_box[190]), .A4(n382), .Y(n42) );
  AO22X1_HVT U48 ( .A1(conv_weight_box[46]), .A2(n381), .A3(
        conv_weight_box[174]), .A4(n380), .Y(n43) );
  OR3X1_HVT U49 ( .A1(n41), .A2(n42), .A3(n43), .Y(n44) );
  OR3X1_HVT U50 ( .A1(n205), .A2(n204), .A3(n203), .Y(n45) );
  AO22X1_HVT U51 ( .A1(conv_weight_box[26]), .A2(n383), .A3(
        conv_weight_box[186]), .A4(n382), .Y(n46) );
  AO22X1_HVT U52 ( .A1(conv_weight_box[42]), .A2(n381), .A3(
        conv_weight_box[170]), .A4(n380), .Y(n47) );
  OR3X1_HVT U53 ( .A1(n45), .A2(n46), .A3(n47), .Y(n48) );
  AO22X1_HVT U54 ( .A1(n399), .A2(n44), .A3(n397), .A4(n48), .Y(n49) );
  NOR4X0_HVT U55 ( .A1(n38), .A2(n39), .A3(n40), .A4(n49), .Y(n50) );
  NAND3X0_HVT U56 ( .A1(n26), .A2(n37), .A3(n50), .Y(n51) );
  AO22X1_HVT U57 ( .A1(n128), .A2(n21), .A3(n129), .A4(n51), .Y(net22436) );
  AO22X1_HVT U58 ( .A1(conv_weight_box[11]), .A2(n288), .A3(
        conv_weight_box[15]), .A4(n289), .Y(n52) );
  AO22X1_HVT U59 ( .A1(conv_weight_box[87]), .A2(n290), .A3(
        conv_weight_box[83]), .A4(n291), .Y(n53) );
  AO22X1_HVT U60 ( .A1(conv_weight_box[23]), .A2(n292), .A3(
        conv_weight_box[75]), .A4(n293), .Y(n54) );
  AO22X1_HVT U61 ( .A1(conv_weight_box[71]), .A2(n294), .A3(
        conv_weight_box[67]), .A4(n295), .Y(n55) );
  NOR4X0_HVT U62 ( .A1(n52), .A2(n53), .A3(n54), .A4(n55), .Y(n56) );
  AO22X1_HVT U63 ( .A1(n326), .A2(conv_weight_box[99]), .A3(n324), .A4(
        conv_weight_box[115]), .Y(n57) );
  AO22X1_HVT U64 ( .A1(conv_weight_box[35]), .A2(n320), .A3(
        conv_weight_box[51]), .A4(n318), .Y(n58) );
  AO22X1_HVT U65 ( .A1(conv_weight_box[179]), .A2(n317), .A3(
        conv_weight_box[195]), .A4(n319), .Y(n59) );
  AO22X1_HVT U66 ( .A1(n322), .A2(conv_weight_box[147]), .A3(n321), .A4(
        conv_weight_box[163]), .Y(n60) );
  NOR4X0_HVT U67 ( .A1(n57), .A2(n58), .A3(n59), .A4(n60), .Y(n61) );
  AO22X1_HVT U68 ( .A1(n326), .A2(conv_weight_box[103]), .A3(n324), .A4(
        conv_weight_box[119]), .Y(n62) );
  AO22X1_HVT U69 ( .A1(conv_weight_box[39]), .A2(n320), .A3(
        conv_weight_box[55]), .A4(n318), .Y(n63) );
  AO22X1_HVT U70 ( .A1(conv_weight_box[199]), .A2(n319), .A3(
        conv_weight_box[183]), .A4(n317), .Y(n64) );
  AO22X1_HVT U71 ( .A1(n322), .A2(conv_weight_box[151]), .A3(n321), .A4(
        conv_weight_box[167]), .Y(n65) );
  NOR4X0_HVT U72 ( .A1(n62), .A2(n63), .A3(n64), .A4(n65), .Y(n66) );
  OA22X1_HVT U73 ( .A1(n61), .A2(n284), .A3(n66), .A4(n286), .Y(n67) );
  AO22X1_HVT U74 ( .A1(conv_weight_box[79]), .A2(n306), .A3(
        conv_weight_box[131]), .A4(n307), .Y(n68) );
  AO22X1_HVT U75 ( .A1(conv_weight_box[135]), .A2(n300), .A3(
        conv_weight_box[19]), .A4(n301), .Y(n69) );
  AO22X1_HVT U76 ( .A1(conv_weight_box[7]), .A2(n302), .A3(conv_weight_box[3]), 
        .A4(n303), .Y(n70) );
  OR3X1_HVT U77 ( .A1(n154), .A2(n153), .A3(n152), .Y(n71) );
  AO22X1_HVT U78 ( .A1(conv_weight_box[31]), .A2(n320), .A3(
        conv_weight_box[191]), .A4(n319), .Y(n72) );
  AO22X1_HVT U79 ( .A1(conv_weight_box[47]), .A2(n318), .A3(
        conv_weight_box[175]), .A4(n317), .Y(n73) );
  OR3X1_HVT U80 ( .A1(n71), .A2(n72), .A3(n73), .Y(n74) );
  OR3X1_HVT U81 ( .A1(n157), .A2(n156), .A3(n155), .Y(n75) );
  AO22X1_HVT U82 ( .A1(conv_weight_box[27]), .A2(n320), .A3(
        conv_weight_box[187]), .A4(n319), .Y(n76) );
  AO22X1_HVT U83 ( .A1(conv_weight_box[43]), .A2(n318), .A3(
        conv_weight_box[171]), .A4(n317), .Y(n77) );
  OR3X1_HVT U84 ( .A1(n75), .A2(n76), .A3(n77), .Y(n78) );
  AO22X1_HVT U85 ( .A1(n336), .A2(n74), .A3(n334), .A4(n78), .Y(n79) );
  NOR4X0_HVT U86 ( .A1(n68), .A2(n69), .A3(n70), .A4(n79), .Y(n80) );
  NAND3X0_HVT U87 ( .A1(n56), .A2(n67), .A3(n80), .Y(n81) );
  AO22X1_HVT U88 ( .A1(conv_weight_box[11]), .A2(n353), .A3(
        conv_weight_box[15]), .A4(n354), .Y(n82) );
  AO22X1_HVT U89 ( .A1(conv_weight_box[87]), .A2(n355), .A3(
        conv_weight_box[83]), .A4(n356), .Y(n83) );
  AO22X1_HVT U90 ( .A1(conv_weight_box[23]), .A2(n357), .A3(
        conv_weight_box[75]), .A4(n358), .Y(n84) );
  AO22X1_HVT U91 ( .A1(conv_weight_box[71]), .A2(n359), .A3(
        conv_weight_box[67]), .A4(n360), .Y(n85) );
  NOR4X0_HVT U92 ( .A1(n82), .A2(n83), .A3(n84), .A4(n85), .Y(n86) );
  AO22X1_HVT U93 ( .A1(n387), .A2(conv_weight_box[115]), .A3(n389), .A4(
        conv_weight_box[99]), .Y(n87) );
  AO22X1_HVT U94 ( .A1(n383), .A2(conv_weight_box[35]), .A3(n381), .A4(
        conv_weight_box[51]), .Y(n88) );
  AO22X1_HVT U95 ( .A1(n382), .A2(conv_weight_box[195]), .A3(n380), .A4(
        conv_weight_box[179]), .Y(n89) );
  AO22X1_HVT U96 ( .A1(n385), .A2(conv_weight_box[147]), .A3(n384), .A4(
        conv_weight_box[163]), .Y(n90) );
  NOR4X0_HVT U97 ( .A1(n87), .A2(n88), .A3(n89), .A4(n90), .Y(n91) );
  AO22X1_HVT U98 ( .A1(n383), .A2(conv_weight_box[39]), .A3(n381), .A4(
        conv_weight_box[55]), .Y(n92) );
  NOR4X0_HVT U99 ( .A1(n160), .A2(n161), .A3(n159), .A4(n92), .Y(n93) );
  OA22X1_HVT U100 ( .A1(n91), .A2(n349), .A3(n93), .A4(n351), .Y(n94) );
  AO22X1_HVT U101 ( .A1(conv_weight_box[79]), .A2(n369), .A3(
        conv_weight_box[131]), .A4(n370), .Y(n95) );
  AO22X1_HVT U102 ( .A1(conv_weight_box[135]), .A2(n365), .A3(
        conv_weight_box[19]), .A4(n366), .Y(n96) );
  AO22X1_HVT U103 ( .A1(conv_weight_box[7]), .A2(n367), .A3(conv_weight_box[3]), .A4(n368), .Y(n97) );
  OR3X1_HVT U104 ( .A1(n178), .A2(n177), .A3(n176), .Y(n98) );
  OR3X1_HVT U105 ( .A1(n184), .A2(n183), .A3(n182), .Y(n99) );
  AO22X1_HVT U106 ( .A1(n399), .A2(n98), .A3(n397), .A4(n99), .Y(n100) );
  NOR4X0_HVT U107 ( .A1(n95), .A2(n96), .A3(n97), .A4(n100), .Y(n101) );
  NAND3X0_HVT U108 ( .A1(n86), .A2(n94), .A3(n101), .Y(n102) );
  AO22X1_HVT U109 ( .A1(n128), .A2(n81), .A3(n129), .A4(n102), .Y(net22432) );
  INVX1_HVT U110 ( .A(srstn), .Y(n305) );
  INVX1_HVT U111 ( .A(n124), .Y(n103) );
  INVX0_HVT U112 ( .A(n139), .Y(n121) );
  NAND2X0_HVT U113 ( .A1(load_conv2_bias1_enable), .A2(n137), .Y(n139) );
  INVX1_HVT U114 ( .A(n284), .Y(n151) );
  INVX1_HVT U115 ( .A(n349), .Y(n172) );
  INVX1_HVT U116 ( .A(set_0_), .Y(n170) );
  INVX1_HVT U117 ( .A(n124), .Y(n104) );
  INVX1_HVT U118 ( .A(n305), .Y(n111) );
  INVX1_HVT U119 ( .A(n305), .Y(n106) );
  NOR2X1_HVT U120 ( .A1(load_conv1_bias_enable), .A2(n140), .Y(n128) );
  INVX0_HVT U121 ( .A(n351), .Y(n169) );
  INVX0_HVT U122 ( .A(n286), .Y(n148) );
  INVX0_HVT U123 ( .A(set_1_), .Y(n162) );
  INVX0_HVT U124 ( .A(mode[1]), .Y(n135) );
  INVX1_HVT U125 ( .A(n124), .Y(n127) );
  INVX1_HVT U126 ( .A(n139), .Y(n105) );
  INVX2_HVT U127 ( .A(n106), .Y(n107) );
  INVX2_HVT U128 ( .A(n106), .Y(n108) );
  INVX2_HVT U129 ( .A(n106), .Y(n109) );
  INVX2_HVT U130 ( .A(n106), .Y(n110) );
  INVX2_HVT U131 ( .A(n111), .Y(n112) );
  INVX2_HVT U132 ( .A(n111), .Y(n113) );
  INVX2_HVT U133 ( .A(n111), .Y(n114) );
  INVX2_HVT U134 ( .A(n111), .Y(n115) );
  INVX2_HVT U135 ( .A(n106), .Y(n116) );
  INVX2_HVT U136 ( .A(n106), .Y(n117) );
  INVX2_HVT U137 ( .A(n111), .Y(n118) );
  INVX2_HVT U138 ( .A(n111), .Y(n119) );
  INVX2_HVT U139 ( .A(n139), .Y(n120) );
  INVX2_HVT U140 ( .A(n139), .Y(n122) );
  INVX2_HVT U141 ( .A(n139), .Y(n123) );
  INVX1_HVT U142 ( .A(n136), .Y(n124) );
  INVX2_HVT U143 ( .A(n124), .Y(n125) );
  INVX2_HVT U144 ( .A(n124), .Y(n126) );
  INVX1_HVT U145 ( .A(n158), .Y(n137) );
  NOR4X1_HVT U146 ( .A1(n254), .A2(n253), .A3(n252), .A4(n251), .Y(n274) );
  NOR4X1_HVT U147 ( .A1(n248), .A2(n247), .A3(n246), .A4(n245), .Y(n249) );
  NOR4X1_HVT U148 ( .A1(n244), .A2(n243), .A3(n242), .A4(n241), .Y(n250) );
  NOR4X1_HVT U149 ( .A1(n219), .A2(n218), .A3(n217), .A4(n216), .Y(n239) );
  NOR4X1_HVT U150 ( .A1(n213), .A2(n212), .A3(n211), .A4(n210), .Y(n214) );
  NOR4X1_HVT U151 ( .A1(n209), .A2(n208), .A3(n207), .A4(n206), .Y(n215) );
  NOR4X1_HVT U152 ( .A1(n364), .A2(n363), .A3(n362), .A4(n361), .Y(n402) );
  NOR4X1_HVT U153 ( .A1(n348), .A2(n347), .A3(n346), .A4(n345), .Y(n350) );
  NOR4X1_HVT U154 ( .A1(n344), .A2(n343), .A3(n342), .A4(n341), .Y(n352) );
  NOR4X1_HVT U155 ( .A1(n299), .A2(n298), .A3(n297), .A4(n296), .Y(n339) );
  NOR4X1_HVT U156 ( .A1(n283), .A2(n282), .A3(n281), .A4(n280), .Y(n285) );
  NOR4X1_HVT U157 ( .A1(n279), .A2(n278), .A3(n277), .A4(n276), .Y(n287) );
  AND2X1_HVT U158 ( .A1(set_4_), .A2(n168), .Y(n388) );
  AND2X1_HVT U159 ( .A1(set_5_), .A2(n168), .Y(n386) );
  INVX1_HVT U160 ( .A(set_4_), .Y(n167) );
  INVX1_HVT U161 ( .A(set_5_), .Y(n171) );
  AND3X1_HVT U162 ( .A1(set_5_), .A2(set_3_), .A3(n166), .Y(n383) );
  AND3X1_HVT U163 ( .A1(set_2_), .A2(set_5_), .A3(n165), .Y(n381) );
  AND3X1_HVT U164 ( .A1(set_3_), .A2(set_4_), .A3(n166), .Y(n389) );
  INVX1_HVT U165 ( .A(set_2_), .Y(n166) );
  AND3X1_HVT U166 ( .A1(set_2_), .A2(set_4_), .A3(n165), .Y(n387) );
  INVX1_HVT U167 ( .A(set_3_), .Y(n165) );
  AND2X1_HVT U168 ( .A1(conv1_bias_set_4_), .A2(n147), .Y(n325) );
  AND2X1_HVT U169 ( .A1(conv1_bias_set_5_), .A2(n147), .Y(n323) );
  INVX1_HVT U170 ( .A(conv1_bias_set_0_), .Y(n149) );
  INVX1_HVT U171 ( .A(conv1_bias_set_1_), .Y(n141) );
  INVX1_HVT U172 ( .A(conv1_bias_set_4_), .Y(n146) );
  INVX1_HVT U173 ( .A(conv1_bias_set_5_), .Y(n150) );
  AND3X1_HVT U174 ( .A1(conv1_bias_set_5_), .A2(conv1_bias_set_3_), .A3(n145), 
        .Y(n320) );
  AND3X1_HVT U175 ( .A1(conv1_bias_set_2_), .A2(conv1_bias_set_5_), .A3(n144), 
        .Y(n318) );
  AND3X1_HVT U176 ( .A1(conv1_bias_set_2_), .A2(conv1_bias_set_4_), .A3(n144), 
        .Y(n324) );
  INVX1_HVT U177 ( .A(conv1_bias_set_3_), .Y(n144) );
  AND3X1_HVT U178 ( .A1(conv1_bias_set_3_), .A2(conv1_bias_set_4_), .A3(n145), 
        .Y(n326) );
  INVX1_HVT U179 ( .A(conv1_bias_set_2_), .Y(n145) );
  NAND2X0_HVT U180 ( .A1(srstn), .A2(n134), .Y(net22224) );
  INVX1_HVT U181 ( .A(load_conv2_bias0_enable), .Y(n138) );
  NAND4X0_HVT U182 ( .A1(n337), .A2(n340), .A3(n339), .A4(n338), .Y(n131) );
  NAND4X0_HVT U183 ( .A1(n400), .A2(n403), .A3(n402), .A4(n401), .Y(n130) );
  AO22X1_HVT U184 ( .A1(n131), .A2(n128), .A3(n129), .A4(n130), .Y(net22444)
         );
  NAND4X0_HVT U185 ( .A1(n237), .A2(n240), .A3(n239), .A4(n238), .Y(n133) );
  NAND4X0_HVT U186 ( .A1(n272), .A2(n275), .A3(n274), .A4(n273), .Y(n132) );
  AO22X1_HVT U187 ( .A1(n133), .A2(n128), .A3(n129), .A4(n132), .Y(net22440)
         );
  NAND2X0_HVT U188 ( .A1(mode[0]), .A2(n135), .Y(n140) );
  AO221X1_HVT U189 ( .A1(n137), .A2(n138), .A3(n158), .A4(n140), .A5(n128), 
        .Y(n134) );
  AND2X1_HVT U190 ( .A1(delay_weight[99]), .A2(n126), .Y(net22070) );
  AND2X1_HVT U191 ( .A1(delay_weight[98]), .A2(n103), .Y(net22073) );
  AND2X1_HVT U192 ( .A1(delay_weight[97]), .A2(n126), .Y(net22074) );
  AND2X1_HVT U193 ( .A1(delay_weight[96]), .A2(n125), .Y(net22075) );
  AND2X1_HVT U194 ( .A1(delay_weight[95]), .A2(n136), .Y(net22076) );
  AND2X1_HVT U195 ( .A1(delay_weight[94]), .A2(n125), .Y(net22077) );
  AND2X1_HVT U196 ( .A1(delay_weight[93]), .A2(n104), .Y(net22078) );
  AND2X1_HVT U197 ( .A1(delay_weight[92]), .A2(n125), .Y(net22079) );
  AND2X1_HVT U198 ( .A1(delay_weight[91]), .A2(n104), .Y(net22080) );
  AND2X1_HVT U199 ( .A1(delay_weight[90]), .A2(n136), .Y(net22081) );
  AND2X1_HVT U200 ( .A1(delay_weight[89]), .A2(n125), .Y(net22089) );
  AND2X1_HVT U201 ( .A1(delay_weight[88]), .A2(n126), .Y(net22090) );
  AND2X1_HVT U202 ( .A1(delay_weight[87]), .A2(n125), .Y(net22091) );
  AND2X1_HVT U203 ( .A1(delay_weight[86]), .A2(n126), .Y(net22092) );
  AND2X1_HVT U204 ( .A1(delay_weight[85]), .A2(n103), .Y(net22093) );
  AND2X1_HVT U205 ( .A1(delay_weight[84]), .A2(n136), .Y(net22094) );
  AND2X1_HVT U206 ( .A1(delay_weight[83]), .A2(n127), .Y(net22095) );
  AND2X1_HVT U207 ( .A1(delay_weight[82]), .A2(n136), .Y(net22096) );
  AND2X1_HVT U208 ( .A1(delay_weight[81]), .A2(n103), .Y(net22097) );
  AND2X1_HVT U209 ( .A1(delay_weight[80]), .A2(n125), .Y(net22098) );
  AND2X1_HVT U210 ( .A1(delay_weight[79]), .A2(n126), .Y(net22106) );
  AND2X1_HVT U211 ( .A1(delay_weight[78]), .A2(n126), .Y(net22107) );
  AND2X1_HVT U212 ( .A1(delay_weight[77]), .A2(n103), .Y(net22108) );
  AND2X1_HVT U213 ( .A1(delay_weight[76]), .A2(n125), .Y(net22109) );
  AND2X1_HVT U214 ( .A1(delay_weight[75]), .A2(n104), .Y(net22110) );
  AND2X1_HVT U215 ( .A1(delay_weight[74]), .A2(n104), .Y(net22111) );
  AND2X1_HVT U216 ( .A1(delay_weight[73]), .A2(n104), .Y(net22112) );
  AND2X1_HVT U217 ( .A1(delay_weight[72]), .A2(n126), .Y(net22113) );
  AND2X1_HVT U218 ( .A1(delay_weight[71]), .A2(n126), .Y(net22114) );
  AND2X1_HVT U219 ( .A1(delay_weight[70]), .A2(n126), .Y(net22115) );
  AND2X1_HVT U220 ( .A1(delay_weight[69]), .A2(n103), .Y(net22123) );
  AND2X1_HVT U221 ( .A1(delay_weight[68]), .A2(n136), .Y(net22124) );
  AND2X1_HVT U222 ( .A1(delay_weight[67]), .A2(n127), .Y(net22125) );
  AND2X1_HVT U223 ( .A1(delay_weight[66]), .A2(n125), .Y(net22126) );
  AND2X1_HVT U224 ( .A1(delay_weight[65]), .A2(n104), .Y(net22127) );
  AND2X1_HVT U225 ( .A1(delay_weight[64]), .A2(n104), .Y(net22128) );
  AND2X1_HVT U226 ( .A1(delay_weight[63]), .A2(n126), .Y(net22129) );
  AND2X1_HVT U227 ( .A1(delay_weight[62]), .A2(n125), .Y(net22130) );
  AND2X1_HVT U228 ( .A1(delay_weight[61]), .A2(n103), .Y(net22131) );
  AND2X1_HVT U229 ( .A1(delay_weight[60]), .A2(n125), .Y(net22132) );
  AND2X1_HVT U230 ( .A1(delay_weight[59]), .A2(n126), .Y(net22140) );
  AND2X1_HVT U231 ( .A1(delay_weight[58]), .A2(n125), .Y(net22141) );
  AND2X1_HVT U232 ( .A1(delay_weight[57]), .A2(n104), .Y(net22142) );
  AND2X1_HVT U233 ( .A1(delay_weight[56]), .A2(n136), .Y(net22143) );
  AND2X1_HVT U234 ( .A1(delay_weight[55]), .A2(n127), .Y(net22144) );
  AND2X1_HVT U235 ( .A1(delay_weight[54]), .A2(n136), .Y(net22145) );
  AND2X1_HVT U236 ( .A1(delay_weight[53]), .A2(n103), .Y(net22146) );
  AND2X1_HVT U237 ( .A1(delay_weight[52]), .A2(n126), .Y(net22147) );
  AND2X1_HVT U238 ( .A1(delay_weight[51]), .A2(n125), .Y(net22148) );
  AND2X1_HVT U239 ( .A1(delay_weight[50]), .A2(n103), .Y(net22149) );
  AND2X1_HVT U240 ( .A1(delay_weight[49]), .A2(n103), .Y(net22157) );
  AND2X1_HVT U241 ( .A1(delay_weight[48]), .A2(n136), .Y(net22158) );
  AND2X1_HVT U242 ( .A1(delay_weight[47]), .A2(n125), .Y(net22159) );
  AND2X1_HVT U243 ( .A1(delay_weight[46]), .A2(n136), .Y(net22160) );
  AND2X1_HVT U244 ( .A1(delay_weight[45]), .A2(n103), .Y(net22161) );
  AND2X1_HVT U245 ( .A1(delay_weight[44]), .A2(n126), .Y(net22162) );
  AND2X1_HVT U246 ( .A1(delay_weight[43]), .A2(n127), .Y(net22163) );
  AND2X1_HVT U247 ( .A1(delay_weight[42]), .A2(n126), .Y(net22164) );
  AND2X1_HVT U248 ( .A1(delay_weight[41]), .A2(n126), .Y(net22165) );
  AND2X1_HVT U249 ( .A1(delay_weight[40]), .A2(n125), .Y(net22166) );
  AND2X1_HVT U250 ( .A1(delay_weight[39]), .A2(n104), .Y(net22174) );
  AND2X1_HVT U251 ( .A1(delay_weight[38]), .A2(n104), .Y(net22175) );
  AND2X1_HVT U252 ( .A1(delay_weight[37]), .A2(n104), .Y(net22176) );
  AND2X1_HVT U253 ( .A1(delay_weight[36]), .A2(n126), .Y(net22177) );
  AND2X1_HVT U254 ( .A1(delay_weight[35]), .A2(n125), .Y(net22178) );
  AND2X1_HVT U255 ( .A1(delay_weight[34]), .A2(n126), .Y(net22179) );
  AND2X1_HVT U256 ( .A1(delay_weight[33]), .A2(n103), .Y(net22180) );
  AND2X1_HVT U257 ( .A1(delay_weight[32]), .A2(n126), .Y(net22181) );
  AND2X1_HVT U258 ( .A1(delay_weight[31]), .A2(n127), .Y(net22182) );
  AND2X1_HVT U259 ( .A1(delay_weight[30]), .A2(n125), .Y(net22183) );
  AND2X1_HVT U260 ( .A1(delay_weight[29]), .A2(n104), .Y(net22191) );
  AND2X1_HVT U261 ( .A1(delay_weight[28]), .A2(n104), .Y(net22192) );
  AND2X1_HVT U262 ( .A1(delay_weight[27]), .A2(n126), .Y(net22193) );
  AND2X1_HVT U263 ( .A1(delay_weight[26]), .A2(n103), .Y(net22194) );
  AND2X1_HVT U264 ( .A1(delay_weight[25]), .A2(n103), .Y(net22195) );
  AND2X1_HVT U265 ( .A1(delay_weight[24]), .A2(n125), .Y(net22196) );
  AND2X1_HVT U266 ( .A1(delay_weight[23]), .A2(n136), .Y(net22197) );
  AND2X1_HVT U267 ( .A1(delay_weight[22]), .A2(n125), .Y(net22198) );
  AND2X1_HVT U268 ( .A1(delay_weight[21]), .A2(n104), .Y(net22199) );
  AND2X1_HVT U269 ( .A1(delay_weight[20]), .A2(n125), .Y(net22200) );
  AND2X1_HVT U270 ( .A1(delay_weight[19]), .A2(n127), .Y(net22208) );
  AND2X1_HVT U271 ( .A1(delay_weight[18]), .A2(n136), .Y(net22209) );
  AND2X1_HVT U272 ( .A1(delay_weight[17]), .A2(n125), .Y(net22210) );
  AND2X1_HVT U273 ( .A1(delay_weight[16]), .A2(n126), .Y(net22211) );
  AND2X1_HVT U274 ( .A1(delay_weight[15]), .A2(n125), .Y(net22212) );
  AND2X1_HVT U275 ( .A1(delay_weight[14]), .A2(n126), .Y(net22213) );
  AND2X1_HVT U276 ( .A1(delay_weight[13]), .A2(n103), .Y(net22214) );
  AND2X1_HVT U277 ( .A1(delay_weight[12]), .A2(n136), .Y(net22215) );
  AND2X1_HVT U278 ( .A1(delay_weight[11]), .A2(n103), .Y(net22216) );
  AND2X1_HVT U279 ( .A1(delay_weight[10]), .A2(n136), .Y(net22217) );
  AND2X1_HVT U280 ( .A1(delay_weight[9]), .A2(n103), .Y(net22225) );
  AND2X1_HVT U281 ( .A1(delay_weight[8]), .A2(n125), .Y(net22226) );
  AND2X1_HVT U282 ( .A1(delay_weight[7]), .A2(n127), .Y(net22227) );
  AND2X1_HVT U283 ( .A1(delay_weight[6]), .A2(n126), .Y(net22228) );
  AND2X1_HVT U284 ( .A1(delay_weight[5]), .A2(n103), .Y(net22229) );
  AND2X1_HVT U285 ( .A1(delay_weight[4]), .A2(n125), .Y(net22230) );
  AND2X1_HVT U286 ( .A1(delay_weight[3]), .A2(n104), .Y(net22231) );
  AND2X1_HVT U287 ( .A1(delay_weight[2]), .A2(n104), .Y(net22232) );
  AND2X1_HVT U288 ( .A1(delay_weight[1]), .A2(n104), .Y(net22233) );
  AND2X1_HVT U289 ( .A1(delay_weight[0]), .A2(n126), .Y(net22234) );
  AO21X1_HVT U290 ( .A1(n105), .A2(n138), .A3(n305), .Y(net22402) );
  AND2X1_HVT U291 ( .A1(delay_weight[99]), .A2(n122), .Y(net22250) );
  AND2X1_HVT U292 ( .A1(delay_weight[98]), .A2(n122), .Y(net22251) );
  AND2X1_HVT U293 ( .A1(delay_weight[97]), .A2(n121), .Y(net22252) );
  AND2X1_HVT U294 ( .A1(delay_weight[96]), .A2(n123), .Y(net22253) );
  AND2X1_HVT U295 ( .A1(delay_weight[95]), .A2(n105), .Y(net22254) );
  AND2X1_HVT U296 ( .A1(delay_weight[94]), .A2(n120), .Y(net22255) );
  AND2X1_HVT U297 ( .A1(delay_weight[93]), .A2(n123), .Y(net22256) );
  AND2X1_HVT U298 ( .A1(delay_weight[92]), .A2(n120), .Y(net22257) );
  AND2X1_HVT U299 ( .A1(delay_weight[91]), .A2(n123), .Y(net22258) );
  AND2X1_HVT U300 ( .A1(delay_weight[90]), .A2(n123), .Y(net22259) );
  AND2X1_HVT U301 ( .A1(delay_weight[89]), .A2(n123), .Y(net22267) );
  AND2X1_HVT U302 ( .A1(delay_weight[88]), .A2(n120), .Y(net22268) );
  AND2X1_HVT U303 ( .A1(delay_weight[87]), .A2(n120), .Y(net22269) );
  AND2X1_HVT U304 ( .A1(delay_weight[86]), .A2(n105), .Y(net22270) );
  AND2X1_HVT U305 ( .A1(delay_weight[85]), .A2(n122), .Y(net22271) );
  AND2X1_HVT U306 ( .A1(delay_weight[84]), .A2(n120), .Y(net22272) );
  AND2X1_HVT U307 ( .A1(delay_weight[83]), .A2(n122), .Y(net22273) );
  AND2X1_HVT U308 ( .A1(delay_weight[82]), .A2(n122), .Y(net22274) );
  AND2X1_HVT U309 ( .A1(delay_weight[81]), .A2(n120), .Y(net22275) );
  AND2X1_HVT U310 ( .A1(delay_weight[80]), .A2(n120), .Y(net22276) );
  AND2X1_HVT U311 ( .A1(delay_weight[79]), .A2(n122), .Y(net22284) );
  AND2X1_HVT U312 ( .A1(delay_weight[78]), .A2(n121), .Y(net22285) );
  AND2X1_HVT U313 ( .A1(delay_weight[77]), .A2(n105), .Y(net22286) );
  AND2X1_HVT U314 ( .A1(delay_weight[76]), .A2(n121), .Y(net22287) );
  AND2X1_HVT U315 ( .A1(delay_weight[75]), .A2(n121), .Y(net22288) );
  AND2X1_HVT U316 ( .A1(delay_weight[74]), .A2(n123), .Y(net22289) );
  AND2X1_HVT U317 ( .A1(delay_weight[73]), .A2(n120), .Y(net22290) );
  AND2X1_HVT U318 ( .A1(delay_weight[72]), .A2(n121), .Y(net22291) );
  AND2X1_HVT U319 ( .A1(delay_weight[71]), .A2(n122), .Y(net22292) );
  AND2X1_HVT U320 ( .A1(delay_weight[70]), .A2(n121), .Y(net22293) );
  AND2X1_HVT U321 ( .A1(delay_weight[69]), .A2(n121), .Y(net22301) );
  AND2X1_HVT U322 ( .A1(delay_weight[68]), .A2(n105), .Y(net22302) );
  AND2X1_HVT U323 ( .A1(delay_weight[67]), .A2(n123), .Y(net22303) );
  AND2X1_HVT U324 ( .A1(delay_weight[66]), .A2(n122), .Y(net22304) );
  AND2X1_HVT U325 ( .A1(delay_weight[65]), .A2(n120), .Y(net22305) );
  AND2X1_HVT U326 ( .A1(delay_weight[64]), .A2(n123), .Y(net22306) );
  AND2X1_HVT U327 ( .A1(delay_weight[63]), .A2(n122), .Y(net22307) );
  AND2X1_HVT U328 ( .A1(delay_weight[62]), .A2(n123), .Y(net22308) );
  AND2X1_HVT U329 ( .A1(delay_weight[61]), .A2(n123), .Y(net22309) );
  AND2X1_HVT U330 ( .A1(delay_weight[60]), .A2(n121), .Y(net22310) );
  AND2X1_HVT U331 ( .A1(delay_weight[59]), .A2(n105), .Y(net22318) );
  AND2X1_HVT U332 ( .A1(delay_weight[58]), .A2(n122), .Y(net22319) );
  AND2X1_HVT U333 ( .A1(delay_weight[57]), .A2(n123), .Y(net22320) );
  AND2X1_HVT U334 ( .A1(delay_weight[56]), .A2(n121), .Y(net22321) );
  AND2X1_HVT U335 ( .A1(delay_weight[55]), .A2(n121), .Y(net22322) );
  AND2X1_HVT U336 ( .A1(delay_weight[54]), .A2(n123), .Y(net22323) );
  AND2X1_HVT U337 ( .A1(delay_weight[53]), .A2(n120), .Y(net22324) );
  AND2X1_HVT U338 ( .A1(delay_weight[52]), .A2(n122), .Y(net22325) );
  AND2X1_HVT U339 ( .A1(delay_weight[51]), .A2(n121), .Y(net22326) );
  AND2X1_HVT U340 ( .A1(delay_weight[50]), .A2(n105), .Y(net22327) );
  AND2X1_HVT U341 ( .A1(delay_weight[49]), .A2(n120), .Y(net22335) );
  AND2X1_HVT U342 ( .A1(delay_weight[48]), .A2(n120), .Y(net22336) );
  AND2X1_HVT U343 ( .A1(delay_weight[47]), .A2(n122), .Y(net22337) );
  AND2X1_HVT U344 ( .A1(delay_weight[46]), .A2(n120), .Y(net22338) );
  AND2X1_HVT U345 ( .A1(delay_weight[45]), .A2(n122), .Y(net22339) );
  AND2X1_HVT U346 ( .A1(delay_weight[44]), .A2(n121), .Y(net22340) );
  AND2X1_HVT U347 ( .A1(delay_weight[43]), .A2(n120), .Y(net22341) );
  AND2X1_HVT U348 ( .A1(delay_weight[42]), .A2(n120), .Y(net22342) );
  AND2X1_HVT U349 ( .A1(delay_weight[41]), .A2(n105), .Y(net22343) );
  AND2X1_HVT U350 ( .A1(delay_weight[40]), .A2(n123), .Y(net22344) );
  AND2X1_HVT U351 ( .A1(delay_weight[39]), .A2(n121), .Y(net22352) );
  AND2X1_HVT U352 ( .A1(delay_weight[38]), .A2(n123), .Y(net22353) );
  AND2X1_HVT U353 ( .A1(delay_weight[37]), .A2(n122), .Y(net22354) );
  AND2X1_HVT U354 ( .A1(delay_weight[36]), .A2(n123), .Y(net22355) );
  AND2X1_HVT U355 ( .A1(delay_weight[35]), .A2(n122), .Y(net22356) );
  AND2X1_HVT U356 ( .A1(delay_weight[34]), .A2(n123), .Y(net22357) );
  AND2X1_HVT U357 ( .A1(delay_weight[33]), .A2(n122), .Y(net22358) );
  AND2X1_HVT U358 ( .A1(delay_weight[32]), .A2(n105), .Y(net22359) );
  AND2X1_HVT U359 ( .A1(delay_weight[31]), .A2(n122), .Y(net22360) );
  AND2X1_HVT U360 ( .A1(delay_weight[30]), .A2(n121), .Y(net22361) );
  AND2X1_HVT U361 ( .A1(delay_weight[29]), .A2(n120), .Y(net22369) );
  AND2X1_HVT U362 ( .A1(delay_weight[28]), .A2(n121), .Y(net22370) );
  AND2X1_HVT U363 ( .A1(delay_weight[27]), .A2(n120), .Y(net22371) );
  AND2X1_HVT U364 ( .A1(delay_weight[26]), .A2(n123), .Y(net22372) );
  AND2X1_HVT U365 ( .A1(delay_weight[25]), .A2(n122), .Y(net22373) );
  AND2X1_HVT U366 ( .A1(delay_weight[24]), .A2(n123), .Y(net22374) );
  AND2X1_HVT U367 ( .A1(delay_weight[23]), .A2(n105), .Y(net22375) );
  AND2X1_HVT U368 ( .A1(delay_weight[22]), .A2(n120), .Y(net22376) );
  AND2X1_HVT U369 ( .A1(delay_weight[21]), .A2(n105), .Y(net22377) );
  AND2X1_HVT U370 ( .A1(delay_weight[20]), .A2(n122), .Y(net22378) );
  AND2X1_HVT U371 ( .A1(delay_weight[19]), .A2(n123), .Y(net22386) );
  AND2X1_HVT U372 ( .A1(delay_weight[18]), .A2(n121), .Y(net22387) );
  AND2X1_HVT U373 ( .A1(delay_weight[17]), .A2(n120), .Y(net22388) );
  AND2X1_HVT U374 ( .A1(delay_weight[16]), .A2(n120), .Y(net22389) );
  AND2X1_HVT U375 ( .A1(delay_weight[15]), .A2(n120), .Y(net22390) );
  AND2X1_HVT U376 ( .A1(delay_weight[14]), .A2(n105), .Y(net22391) );
  AND2X1_HVT U377 ( .A1(delay_weight[13]), .A2(n123), .Y(net22392) );
  AND2X1_HVT U378 ( .A1(delay_weight[12]), .A2(n105), .Y(net22393) );
  AND2X1_HVT U379 ( .A1(delay_weight[11]), .A2(n123), .Y(net22394) );
  AND2X1_HVT U380 ( .A1(delay_weight[10]), .A2(n122), .Y(net22395) );
  AND2X1_HVT U381 ( .A1(delay_weight[9]), .A2(n122), .Y(net22403) );
  AND2X1_HVT U382 ( .A1(delay_weight[8]), .A2(n122), .Y(net22404) );
  AND2X1_HVT U383 ( .A1(delay_weight[7]), .A2(n123), .Y(net22405) );
  AND2X1_HVT U384 ( .A1(delay_weight[6]), .A2(n121), .Y(net22406) );
  AND2X1_HVT U385 ( .A1(delay_weight[5]), .A2(n105), .Y(net22407) );
  AND2X1_HVT U386 ( .A1(delay_weight[4]), .A2(n122), .Y(net22408) );
  AND2X1_HVT U387 ( .A1(delay_weight[3]), .A2(n105), .Y(net22409) );
  AND2X1_HVT U388 ( .A1(delay_weight[2]), .A2(n120), .Y(net22410) );
  AND2X1_HVT U389 ( .A1(delay_weight[1]), .A2(n120), .Y(net22411) );
  AND2X1_HVT U390 ( .A1(delay_weight[0]), .A2(n123), .Y(net22412) );
  NAND3X0_HVT U391 ( .A1(srstn), .A2(n140), .A3(n158), .Y(net22426) );
  AND4X1_HVT U392 ( .A1(conv1_bias_set_2_), .A2(n150), .A3(n144), .A4(n146), 
        .Y(n317) );
  AND4X1_HVT U393 ( .A1(n150), .A2(n145), .A3(n144), .A4(n146), .Y(n319) );
  AND4X1_HVT U394 ( .A1(conv1_bias_set_2_), .A2(conv1_bias_set_3_), .A3(n150), 
        .A4(n146), .Y(n322) );
  AND4X1_HVT U395 ( .A1(conv1_bias_set_3_), .A2(n150), .A3(n145), .A4(n146), 
        .Y(n321) );
  NAND2X0_HVT U396 ( .A1(n141), .A2(n149), .Y(n286) );
  NAND2X0_HVT U397 ( .A1(conv1_bias_set_0_), .A2(n141), .Y(n284) );
  AND2X1_HVT U398 ( .A1(conv1_bias_set_1_), .A2(n149), .Y(n336) );
  AND4X1_HVT U399 ( .A1(n336), .A2(conv1_bias_set_5_), .A3(conv1_bias_set_2_), 
        .A4(conv1_bias_set_3_), .Y(n289) );
  AND3X1_HVT U400 ( .A1(conv1_bias_set_5_), .A2(conv1_bias_set_2_), .A3(
        conv1_bias_set_3_), .Y(n142) );
  AND3X1_HVT U401 ( .A1(conv1_bias_set_1_), .A2(conv1_bias_set_0_), .A3(n142), 
        .Y(n288) );
  AND4X1_HVT U402 ( .A1(conv1_bias_set_2_), .A2(conv1_bias_set_3_), .A3(
        conv1_bias_set_4_), .A4(n151), .Y(n291) );
  AND4X1_HVT U403 ( .A1(conv1_bias_set_2_), .A2(conv1_bias_set_3_), .A3(
        conv1_bias_set_4_), .A4(n148), .Y(n290) );
  AND3X1_HVT U404 ( .A1(conv1_bias_set_2_), .A2(conv1_bias_set_3_), .A3(
        conv1_bias_set_4_), .Y(n143) );
  AND3X1_HVT U405 ( .A1(conv1_bias_set_1_), .A2(conv1_bias_set_0_), .A3(n143), 
        .Y(n293) );
  AND4X1_HVT U406 ( .A1(conv1_bias_set_5_), .A2(conv1_bias_set_2_), .A3(
        conv1_bias_set_3_), .A4(n148), .Y(n292) );
  AND2X1_HVT U407 ( .A1(n145), .A2(n144), .Y(n147) );
  AND3X1_HVT U408 ( .A1(n323), .A2(n151), .A3(n146), .Y(n295) );
  AND3X1_HVT U409 ( .A1(n323), .A2(n148), .A3(n146), .Y(n294) );
  AND4X1_HVT U410 ( .A1(conv1_bias_set_5_), .A2(conv1_bias_set_2_), .A3(
        conv1_bias_set_3_), .A4(n151), .Y(n301) );
  AND3X1_HVT U411 ( .A1(n325), .A2(n148), .A3(n150), .Y(n300) );
  AND3X1_HVT U412 ( .A1(conv1_bias_set_0_), .A2(conv1_bias_set_5_), .A3(
        conv1_bias_set_4_), .Y(n303) );
  AND3X1_HVT U413 ( .A1(conv1_bias_set_5_), .A2(conv1_bias_set_4_), .A3(n149), 
        .Y(n302) );
  AND3X1_HVT U414 ( .A1(n325), .A2(n151), .A3(n150), .Y(n307) );
  AND4X1_HVT U415 ( .A1(n336), .A2(conv1_bias_set_2_), .A3(conv1_bias_set_3_), 
        .A4(conv1_bias_set_4_), .Y(n306) );
  AO22X1_HVT U416 ( .A1(n322), .A2(conv_weight_box[143]), .A3(n321), .A4(
        conv_weight_box[159]), .Y(n154) );
  AO22X1_HVT U417 ( .A1(n324), .A2(conv_weight_box[111]), .A3(n323), .A4(
        conv_weight_box[63]), .Y(n153) );
  AO22X1_HVT U418 ( .A1(n326), .A2(conv_weight_box[95]), .A3(n325), .A4(
        conv_weight_box[127]), .Y(n152) );
  AND2X1_HVT U419 ( .A1(conv1_bias_set_1_), .A2(conv1_bias_set_0_), .Y(n334)
         );
  AO22X1_HVT U420 ( .A1(n322), .A2(conv_weight_box[139]), .A3(n321), .A4(
        conv_weight_box[155]), .Y(n157) );
  AO22X1_HVT U421 ( .A1(n324), .A2(conv_weight_box[107]), .A3(n323), .A4(
        conv_weight_box[59]), .Y(n156) );
  AO22X1_HVT U422 ( .A1(n326), .A2(conv_weight_box[91]), .A3(n325), .A4(
        conv_weight_box[123]), .Y(n155) );
  AO22X1_HVT U423 ( .A1(conv_weight_box[119]), .A2(n387), .A3(
        conv_weight_box[103]), .A4(n389), .Y(n161) );
  AND4X1_HVT U424 ( .A1(n171), .A2(n166), .A3(n165), .A4(n167), .Y(n382) );
  AND4X1_HVT U425 ( .A1(set_2_), .A2(n171), .A3(n165), .A4(n167), .Y(n380) );
  AO22X1_HVT U426 ( .A1(conv_weight_box[199]), .A2(n382), .A3(
        conv_weight_box[183]), .A4(n380), .Y(n160) );
  AND4X1_HVT U427 ( .A1(set_2_), .A2(set_3_), .A3(n171), .A4(n167), .Y(n385)
         );
  AND4X1_HVT U428 ( .A1(set_3_), .A2(n171), .A3(n166), .A4(n167), .Y(n384) );
  AO22X1_HVT U429 ( .A1(conv_weight_box[151]), .A2(n385), .A3(
        conv_weight_box[167]), .A4(n384), .Y(n159) );
  NAND2X0_HVT U430 ( .A1(n162), .A2(n170), .Y(n351) );
  NAND2X0_HVT U431 ( .A1(set_0_), .A2(n162), .Y(n349) );
  AND2X1_HVT U432 ( .A1(set_1_), .A2(n170), .Y(n399) );
  AND4X1_HVT U433 ( .A1(n399), .A2(set_5_), .A3(set_2_), .A4(set_3_), .Y(n354)
         );
  AND3X1_HVT U434 ( .A1(set_5_), .A2(set_2_), .A3(set_3_), .Y(n163) );
  AND3X1_HVT U435 ( .A1(set_1_), .A2(set_0_), .A3(n163), .Y(n353) );
  AND4X1_HVT U436 ( .A1(set_2_), .A2(set_3_), .A3(set_4_), .A4(n172), .Y(n356)
         );
  AND4X1_HVT U437 ( .A1(set_2_), .A2(set_3_), .A3(set_4_), .A4(n169), .Y(n355)
         );
  AND3X1_HVT U438 ( .A1(set_2_), .A2(set_3_), .A3(set_4_), .Y(n164) );
  AND3X1_HVT U439 ( .A1(set_1_), .A2(set_0_), .A3(n164), .Y(n358) );
  AND4X1_HVT U440 ( .A1(set_5_), .A2(set_2_), .A3(set_3_), .A4(n169), .Y(n357)
         );
  AND2X1_HVT U441 ( .A1(n166), .A2(n165), .Y(n168) );
  AND3X1_HVT U442 ( .A1(n386), .A2(n172), .A3(n167), .Y(n360) );
  AND3X1_HVT U443 ( .A1(n386), .A2(n169), .A3(n167), .Y(n359) );
  AND4X1_HVT U444 ( .A1(set_5_), .A2(set_2_), .A3(set_3_), .A4(n172), .Y(n366)
         );
  AND3X1_HVT U445 ( .A1(n388), .A2(n169), .A3(n171), .Y(n365) );
  AND3X1_HVT U446 ( .A1(set_0_), .A2(set_5_), .A3(set_4_), .Y(n368) );
  AND3X1_HVT U447 ( .A1(set_5_), .A2(set_4_), .A3(n170), .Y(n367) );
  AND3X1_HVT U448 ( .A1(n388), .A2(n172), .A3(n171), .Y(n370) );
  AND4X1_HVT U449 ( .A1(n399), .A2(set_2_), .A3(set_3_), .A4(set_4_), .Y(n369)
         );
  AO22X1_HVT U450 ( .A1(conv_weight_box[47]), .A2(n381), .A3(
        conv_weight_box[175]), .A4(n380), .Y(n178) );
  AO22X1_HVT U451 ( .A1(conv_weight_box[31]), .A2(n383), .A3(
        conv_weight_box[191]), .A4(n382), .Y(n177) );
  AO22X1_HVT U452 ( .A1(conv_weight_box[143]), .A2(n385), .A3(
        conv_weight_box[159]), .A4(n384), .Y(n175) );
  AO22X1_HVT U453 ( .A1(conv_weight_box[111]), .A2(n387), .A3(
        conv_weight_box[63]), .A4(n386), .Y(n174) );
  AO22X1_HVT U454 ( .A1(conv_weight_box[95]), .A2(n389), .A3(
        conv_weight_box[127]), .A4(n388), .Y(n173) );
  OR3X1_HVT U455 ( .A1(n175), .A2(n174), .A3(n173), .Y(n176) );
  AND2X1_HVT U456 ( .A1(set_1_), .A2(set_0_), .Y(n397) );
  AO22X1_HVT U457 ( .A1(conv_weight_box[43]), .A2(n381), .A3(
        conv_weight_box[171]), .A4(n380), .Y(n184) );
  AO22X1_HVT U458 ( .A1(conv_weight_box[27]), .A2(n383), .A3(
        conv_weight_box[187]), .A4(n382), .Y(n183) );
  AO22X1_HVT U459 ( .A1(conv_weight_box[139]), .A2(n385), .A3(
        conv_weight_box[155]), .A4(n384), .Y(n181) );
  AO22X1_HVT U460 ( .A1(conv_weight_box[107]), .A2(n387), .A3(
        conv_weight_box[59]), .A4(n386), .Y(n180) );
  AO22X1_HVT U461 ( .A1(conv_weight_box[91]), .A2(n389), .A3(
        conv_weight_box[123]), .A4(n388), .Y(n179) );
  OR3X1_HVT U462 ( .A1(n181), .A2(n180), .A3(n179), .Y(n182) );
  AO22X1_HVT U463 ( .A1(n326), .A2(conv_weight_box[102]), .A3(n324), .A4(
        conv_weight_box[118]), .Y(n187) );
  AO22X1_HVT U464 ( .A1(n317), .A2(conv_weight_box[182]), .A3(n319), .A4(
        conv_weight_box[198]), .Y(n186) );
  AO22X1_HVT U465 ( .A1(n322), .A2(conv_weight_box[150]), .A3(n321), .A4(
        conv_weight_box[166]), .Y(n185) );
  AO22X1_HVT U466 ( .A1(n318), .A2(conv_weight_box[46]), .A3(n317), .A4(
        conv_weight_box[174]), .Y(n193) );
  AO22X1_HVT U467 ( .A1(n320), .A2(conv_weight_box[30]), .A3(n319), .A4(
        conv_weight_box[190]), .Y(n192) );
  AO22X1_HVT U468 ( .A1(n322), .A2(conv_weight_box[142]), .A3(n321), .A4(
        conv_weight_box[158]), .Y(n190) );
  AO22X1_HVT U469 ( .A1(n324), .A2(conv_weight_box[110]), .A3(n323), .A4(
        conv_weight_box[62]), .Y(n189) );
  AO22X1_HVT U470 ( .A1(n326), .A2(conv_weight_box[94]), .A3(n325), .A4(
        conv_weight_box[126]), .Y(n188) );
  OR3X1_HVT U471 ( .A1(n190), .A2(n189), .A3(n188), .Y(n191) );
  AO22X1_HVT U472 ( .A1(n318), .A2(conv_weight_box[42]), .A3(n317), .A4(
        conv_weight_box[170]), .Y(n199) );
  AO22X1_HVT U473 ( .A1(n320), .A2(conv_weight_box[26]), .A3(n319), .A4(
        conv_weight_box[186]), .Y(n198) );
  AO22X1_HVT U474 ( .A1(n322), .A2(conv_weight_box[138]), .A3(n321), .A4(
        conv_weight_box[154]), .Y(n196) );
  AO22X1_HVT U475 ( .A1(n324), .A2(conv_weight_box[106]), .A3(n323), .A4(
        conv_weight_box[58]), .Y(n195) );
  AO22X1_HVT U476 ( .A1(n326), .A2(conv_weight_box[90]), .A3(n325), .A4(
        conv_weight_box[122]), .Y(n194) );
  OR3X1_HVT U477 ( .A1(n196), .A2(n195), .A3(n194), .Y(n197) );
  AO22X1_HVT U478 ( .A1(n385), .A2(conv_weight_box[142]), .A3(n384), .A4(
        conv_weight_box[158]), .Y(n202) );
  AO22X1_HVT U479 ( .A1(n387), .A2(conv_weight_box[110]), .A3(n386), .A4(
        conv_weight_box[62]), .Y(n201) );
  AO22X1_HVT U480 ( .A1(n389), .A2(conv_weight_box[94]), .A3(n388), .A4(
        conv_weight_box[126]), .Y(n200) );
  AO22X1_HVT U481 ( .A1(n385), .A2(conv_weight_box[138]), .A3(n384), .A4(
        conv_weight_box[154]), .Y(n205) );
  AO22X1_HVT U482 ( .A1(n387), .A2(conv_weight_box[106]), .A3(n386), .A4(
        conv_weight_box[58]), .Y(n204) );
  AO22X1_HVT U483 ( .A1(n389), .A2(conv_weight_box[90]), .A3(n388), .A4(
        conv_weight_box[122]), .Y(n203) );
  AO22X1_HVT U484 ( .A1(n326), .A2(conv_weight_box[101]), .A3(n324), .A4(
        conv_weight_box[117]), .Y(n209) );
  AO22X1_HVT U485 ( .A1(n318), .A2(conv_weight_box[53]), .A3(n320), .A4(
        conv_weight_box[37]), .Y(n208) );
  AO22X1_HVT U486 ( .A1(n317), .A2(conv_weight_box[181]), .A3(n319), .A4(
        conv_weight_box[197]), .Y(n207) );
  AO22X1_HVT U487 ( .A1(n322), .A2(conv_weight_box[149]), .A3(n321), .A4(
        conv_weight_box[165]), .Y(n206) );
  AO22X1_HVT U488 ( .A1(n326), .A2(conv_weight_box[97]), .A3(n324), .A4(
        conv_weight_box[113]), .Y(n213) );
  AO22X1_HVT U489 ( .A1(n318), .A2(conv_weight_box[49]), .A3(n320), .A4(
        conv_weight_box[33]), .Y(n212) );
  AO22X1_HVT U490 ( .A1(n317), .A2(conv_weight_box[177]), .A3(n319), .A4(
        conv_weight_box[193]), .Y(n211) );
  AO22X1_HVT U491 ( .A1(n322), .A2(conv_weight_box[145]), .A3(n321), .A4(
        conv_weight_box[161]), .Y(n210) );
  OA22X1_HVT U492 ( .A1(n215), .A2(n286), .A3(n214), .A4(n284), .Y(n240) );
  AO22X1_HVT U493 ( .A1(n289), .A2(conv_weight_box[13]), .A3(n288), .A4(
        conv_weight_box[9]), .Y(n219) );
  AO22X1_HVT U494 ( .A1(n291), .A2(conv_weight_box[81]), .A3(n290), .A4(
        conv_weight_box[85]), .Y(n218) );
  AO22X1_HVT U495 ( .A1(n293), .A2(conv_weight_box[73]), .A3(n292), .A4(
        conv_weight_box[21]), .Y(n217) );
  AO22X1_HVT U496 ( .A1(n295), .A2(conv_weight_box[65]), .A3(n294), .A4(
        conv_weight_box[69]), .Y(n216) );
  AO22X1_HVT U497 ( .A1(n301), .A2(conv_weight_box[17]), .A3(n300), .A4(
        conv_weight_box[133]), .Y(n222) );
  AO22X1_HVT U498 ( .A1(n303), .A2(conv_weight_box[1]), .A3(n302), .A4(
        conv_weight_box[5]), .Y(n221) );
  AO22X1_HVT U499 ( .A1(n307), .A2(conv_weight_box[129]), .A3(n306), .A4(
        conv_weight_box[77]), .Y(n220) );
  NOR3X0_HVT U500 ( .A1(n222), .A2(n221), .A3(n220), .Y(n238) );
  AO22X1_HVT U501 ( .A1(n318), .A2(conv_weight_box[45]), .A3(n317), .A4(
        conv_weight_box[173]), .Y(n228) );
  AO22X1_HVT U502 ( .A1(n320), .A2(conv_weight_box[29]), .A3(n319), .A4(
        conv_weight_box[189]), .Y(n227) );
  AO22X1_HVT U503 ( .A1(n322), .A2(conv_weight_box[141]), .A3(n321), .A4(
        conv_weight_box[157]), .Y(n225) );
  AO22X1_HVT U504 ( .A1(n324), .A2(conv_weight_box[109]), .A3(n323), .A4(
        conv_weight_box[61]), .Y(n224) );
  AO22X1_HVT U505 ( .A1(n326), .A2(conv_weight_box[93]), .A3(n325), .A4(
        conv_weight_box[125]), .Y(n223) );
  OR3X1_HVT U506 ( .A1(n225), .A2(n224), .A3(n223), .Y(n226) );
  OR3X1_HVT U507 ( .A1(n228), .A2(n227), .A3(n226), .Y(n236) );
  AO22X1_HVT U508 ( .A1(n318), .A2(conv_weight_box[41]), .A3(n317), .A4(
        conv_weight_box[169]), .Y(n234) );
  AO22X1_HVT U509 ( .A1(n320), .A2(conv_weight_box[25]), .A3(n319), .A4(
        conv_weight_box[185]), .Y(n233) );
  AO22X1_HVT U510 ( .A1(n322), .A2(conv_weight_box[137]), .A3(n321), .A4(
        conv_weight_box[153]), .Y(n231) );
  AO22X1_HVT U511 ( .A1(n324), .A2(conv_weight_box[105]), .A3(n323), .A4(
        conv_weight_box[57]), .Y(n230) );
  AO22X1_HVT U512 ( .A1(n326), .A2(conv_weight_box[89]), .A3(n325), .A4(
        conv_weight_box[121]), .Y(n229) );
  OR3X1_HVT U513 ( .A1(n231), .A2(n230), .A3(n229), .Y(n232) );
  OR3X1_HVT U514 ( .A1(n234), .A2(n233), .A3(n232), .Y(n235) );
  AOI22X1_HVT U515 ( .A1(n336), .A2(n236), .A3(n334), .A4(n235), .Y(n237) );
  AO22X1_HVT U516 ( .A1(n389), .A2(conv_weight_box[101]), .A3(n387), .A4(
        conv_weight_box[117]), .Y(n244) );
  AO22X1_HVT U517 ( .A1(n381), .A2(conv_weight_box[53]), .A3(n383), .A4(
        conv_weight_box[37]), .Y(n243) );
  AO22X1_HVT U518 ( .A1(n380), .A2(conv_weight_box[181]), .A3(n382), .A4(
        conv_weight_box[197]), .Y(n242) );
  AO22X1_HVT U519 ( .A1(n385), .A2(conv_weight_box[149]), .A3(n384), .A4(
        conv_weight_box[165]), .Y(n241) );
  AO22X1_HVT U520 ( .A1(n389), .A2(conv_weight_box[97]), .A3(n387), .A4(
        conv_weight_box[113]), .Y(n248) );
  AO22X1_HVT U521 ( .A1(n381), .A2(conv_weight_box[49]), .A3(n383), .A4(
        conv_weight_box[33]), .Y(n247) );
  AO22X1_HVT U522 ( .A1(n380), .A2(conv_weight_box[177]), .A3(n382), .A4(
        conv_weight_box[193]), .Y(n246) );
  AO22X1_HVT U523 ( .A1(n385), .A2(conv_weight_box[145]), .A3(n384), .A4(
        conv_weight_box[161]), .Y(n245) );
  OA22X1_HVT U524 ( .A1(n250), .A2(n351), .A3(n249), .A4(n349), .Y(n275) );
  AO22X1_HVT U525 ( .A1(n354), .A2(conv_weight_box[13]), .A3(n353), .A4(
        conv_weight_box[9]), .Y(n254) );
  AO22X1_HVT U526 ( .A1(n356), .A2(conv_weight_box[81]), .A3(n355), .A4(
        conv_weight_box[85]), .Y(n253) );
  AO22X1_HVT U527 ( .A1(n358), .A2(conv_weight_box[73]), .A3(n357), .A4(
        conv_weight_box[21]), .Y(n252) );
  AO22X1_HVT U528 ( .A1(n360), .A2(conv_weight_box[65]), .A3(n359), .A4(
        conv_weight_box[69]), .Y(n251) );
  AO22X1_HVT U529 ( .A1(n366), .A2(conv_weight_box[17]), .A3(n365), .A4(
        conv_weight_box[133]), .Y(n257) );
  AO22X1_HVT U530 ( .A1(n368), .A2(conv_weight_box[1]), .A3(n367), .A4(
        conv_weight_box[5]), .Y(n256) );
  AO22X1_HVT U531 ( .A1(n370), .A2(conv_weight_box[129]), .A3(n369), .A4(
        conv_weight_box[77]), .Y(n255) );
  NOR3X0_HVT U532 ( .A1(n257), .A2(n256), .A3(n255), .Y(n273) );
  AO22X1_HVT U533 ( .A1(n381), .A2(conv_weight_box[45]), .A3(n380), .A4(
        conv_weight_box[173]), .Y(n263) );
  AO22X1_HVT U534 ( .A1(n383), .A2(conv_weight_box[29]), .A3(n382), .A4(
        conv_weight_box[189]), .Y(n262) );
  AO22X1_HVT U535 ( .A1(n385), .A2(conv_weight_box[141]), .A3(n384), .A4(
        conv_weight_box[157]), .Y(n260) );
  AO22X1_HVT U536 ( .A1(n387), .A2(conv_weight_box[109]), .A3(n386), .A4(
        conv_weight_box[61]), .Y(n259) );
  AO22X1_HVT U537 ( .A1(n389), .A2(conv_weight_box[93]), .A3(n388), .A4(
        conv_weight_box[125]), .Y(n258) );
  OR3X1_HVT U538 ( .A1(n260), .A2(n259), .A3(n258), .Y(n261) );
  OR3X1_HVT U539 ( .A1(n263), .A2(n262), .A3(n261), .Y(n271) );
  AO22X1_HVT U540 ( .A1(n381), .A2(conv_weight_box[41]), .A3(n380), .A4(
        conv_weight_box[169]), .Y(n269) );
  AO22X1_HVT U541 ( .A1(n383), .A2(conv_weight_box[25]), .A3(n382), .A4(
        conv_weight_box[185]), .Y(n268) );
  AO22X1_HVT U542 ( .A1(n385), .A2(conv_weight_box[137]), .A3(n384), .A4(
        conv_weight_box[153]), .Y(n266) );
  AO22X1_HVT U543 ( .A1(n387), .A2(conv_weight_box[105]), .A3(n386), .A4(
        conv_weight_box[57]), .Y(n265) );
  AO22X1_HVT U544 ( .A1(n389), .A2(conv_weight_box[89]), .A3(n388), .A4(
        conv_weight_box[121]), .Y(n264) );
  OR3X1_HVT U545 ( .A1(n266), .A2(n265), .A3(n264), .Y(n267) );
  OR3X1_HVT U546 ( .A1(n269), .A2(n268), .A3(n267), .Y(n270) );
  AOI22X1_HVT U547 ( .A1(n399), .A2(n271), .A3(n397), .A4(n270), .Y(n272) );
  AO22X1_HVT U548 ( .A1(n326), .A2(conv_weight_box[100]), .A3(n324), .A4(
        conv_weight_box[116]), .Y(n279) );
  AO22X1_HVT U549 ( .A1(n318), .A2(conv_weight_box[52]), .A3(n320), .A4(
        conv_weight_box[36]), .Y(n278) );
  AO22X1_HVT U550 ( .A1(n317), .A2(conv_weight_box[180]), .A3(n319), .A4(
        conv_weight_box[196]), .Y(n277) );
  AO22X1_HVT U551 ( .A1(n322), .A2(conv_weight_box[148]), .A3(n321), .A4(
        conv_weight_box[164]), .Y(n276) );
  AO22X1_HVT U552 ( .A1(n326), .A2(conv_weight_box[96]), .A3(n324), .A4(
        conv_weight_box[112]), .Y(n283) );
  AO22X1_HVT U553 ( .A1(n318), .A2(conv_weight_box[48]), .A3(n320), .A4(
        conv_weight_box[32]), .Y(n282) );
  AO22X1_HVT U554 ( .A1(n317), .A2(conv_weight_box[176]), .A3(n319), .A4(
        conv_weight_box[192]), .Y(n281) );
  AO22X1_HVT U555 ( .A1(n322), .A2(conv_weight_box[144]), .A3(n321), .A4(
        conv_weight_box[160]), .Y(n280) );
  OA22X1_HVT U556 ( .A1(n287), .A2(n286), .A3(n285), .A4(n284), .Y(n340) );
  AO22X1_HVT U557 ( .A1(n289), .A2(conv_weight_box[12]), .A3(n288), .A4(
        conv_weight_box[8]), .Y(n299) );
  AO22X1_HVT U558 ( .A1(n291), .A2(conv_weight_box[80]), .A3(n290), .A4(
        conv_weight_box[84]), .Y(n298) );
  AO22X1_HVT U559 ( .A1(n293), .A2(conv_weight_box[72]), .A3(n292), .A4(
        conv_weight_box[20]), .Y(n297) );
  AO22X1_HVT U560 ( .A1(n295), .A2(conv_weight_box[64]), .A3(n294), .A4(
        conv_weight_box[68]), .Y(n296) );
  AO22X1_HVT U561 ( .A1(n301), .A2(conv_weight_box[16]), .A3(n300), .A4(
        conv_weight_box[132]), .Y(n310) );
  AO22X1_HVT U562 ( .A1(n303), .A2(conv_weight_box[0]), .A3(n302), .A4(
        conv_weight_box[4]), .Y(n309) );
  AO22X1_HVT U563 ( .A1(n307), .A2(conv_weight_box[128]), .A3(n306), .A4(
        conv_weight_box[76]), .Y(n308) );
  NOR3X0_HVT U564 ( .A1(n310), .A2(n309), .A3(n308), .Y(n338) );
  AO22X1_HVT U565 ( .A1(n318), .A2(conv_weight_box[44]), .A3(n317), .A4(
        conv_weight_box[172]), .Y(n316) );
  AO22X1_HVT U566 ( .A1(n320), .A2(conv_weight_box[28]), .A3(n319), .A4(
        conv_weight_box[188]), .Y(n315) );
  AO22X1_HVT U567 ( .A1(n322), .A2(conv_weight_box[140]), .A3(n321), .A4(
        conv_weight_box[156]), .Y(n313) );
  AO22X1_HVT U568 ( .A1(n324), .A2(conv_weight_box[108]), .A3(n323), .A4(
        conv_weight_box[60]), .Y(n312) );
  AO22X1_HVT U569 ( .A1(n326), .A2(conv_weight_box[92]), .A3(n325), .A4(
        conv_weight_box[124]), .Y(n311) );
  OR3X1_HVT U570 ( .A1(n313), .A2(n312), .A3(n311), .Y(n314) );
  OR3X1_HVT U571 ( .A1(n316), .A2(n315), .A3(n314), .Y(n335) );
  AO22X1_HVT U572 ( .A1(n318), .A2(conv_weight_box[40]), .A3(n317), .A4(
        conv_weight_box[168]), .Y(n332) );
  AO22X1_HVT U573 ( .A1(n320), .A2(conv_weight_box[24]), .A3(n319), .A4(
        conv_weight_box[184]), .Y(n331) );
  AO22X1_HVT U574 ( .A1(n322), .A2(conv_weight_box[136]), .A3(n321), .A4(
        conv_weight_box[152]), .Y(n329) );
  AO22X1_HVT U575 ( .A1(n324), .A2(conv_weight_box[104]), .A3(n323), .A4(
        conv_weight_box[56]), .Y(n328) );
  AO22X1_HVT U576 ( .A1(n326), .A2(conv_weight_box[88]), .A3(n325), .A4(
        conv_weight_box[120]), .Y(n327) );
  OR3X1_HVT U577 ( .A1(n329), .A2(n328), .A3(n327), .Y(n330) );
  OR3X1_HVT U578 ( .A1(n332), .A2(n331), .A3(n330), .Y(n333) );
  AOI22X1_HVT U579 ( .A1(n336), .A2(n335), .A3(n334), .A4(n333), .Y(n337) );
  AO22X1_HVT U580 ( .A1(n389), .A2(conv_weight_box[100]), .A3(n387), .A4(
        conv_weight_box[116]), .Y(n344) );
  AO22X1_HVT U581 ( .A1(n381), .A2(conv_weight_box[52]), .A3(n383), .A4(
        conv_weight_box[36]), .Y(n343) );
  AO22X1_HVT U582 ( .A1(n380), .A2(conv_weight_box[180]), .A3(n382), .A4(
        conv_weight_box[196]), .Y(n342) );
  AO22X1_HVT U583 ( .A1(n385), .A2(conv_weight_box[148]), .A3(n384), .A4(
        conv_weight_box[164]), .Y(n341) );
  AO22X1_HVT U584 ( .A1(n389), .A2(conv_weight_box[96]), .A3(n387), .A4(
        conv_weight_box[112]), .Y(n348) );
  AO22X1_HVT U585 ( .A1(n381), .A2(conv_weight_box[48]), .A3(n383), .A4(
        conv_weight_box[32]), .Y(n347) );
  AO22X1_HVT U586 ( .A1(n380), .A2(conv_weight_box[176]), .A3(n382), .A4(
        conv_weight_box[192]), .Y(n346) );
  AO22X1_HVT U587 ( .A1(n385), .A2(conv_weight_box[144]), .A3(n384), .A4(
        conv_weight_box[160]), .Y(n345) );
  OA22X1_HVT U588 ( .A1(n352), .A2(n351), .A3(n350), .A4(n349), .Y(n403) );
  AO22X1_HVT U589 ( .A1(n354), .A2(conv_weight_box[12]), .A3(n353), .A4(
        conv_weight_box[8]), .Y(n364) );
  AO22X1_HVT U590 ( .A1(n356), .A2(conv_weight_box[80]), .A3(n355), .A4(
        conv_weight_box[84]), .Y(n363) );
  AO22X1_HVT U591 ( .A1(n358), .A2(conv_weight_box[72]), .A3(n357), .A4(
        conv_weight_box[20]), .Y(n362) );
  AO22X1_HVT U592 ( .A1(n360), .A2(conv_weight_box[64]), .A3(n359), .A4(
        conv_weight_box[68]), .Y(n361) );
  AO22X1_HVT U593 ( .A1(n366), .A2(conv_weight_box[16]), .A3(n365), .A4(
        conv_weight_box[132]), .Y(n373) );
  AO22X1_HVT U594 ( .A1(n368), .A2(conv_weight_box[0]), .A3(n367), .A4(
        conv_weight_box[4]), .Y(n372) );
  AO22X1_HVT U595 ( .A1(n370), .A2(conv_weight_box[128]), .A3(n369), .A4(
        conv_weight_box[76]), .Y(n371) );
  NOR3X0_HVT U596 ( .A1(n373), .A2(n372), .A3(n371), .Y(n401) );
  AO22X1_HVT U597 ( .A1(n381), .A2(conv_weight_box[44]), .A3(n380), .A4(
        conv_weight_box[172]), .Y(n379) );
  AO22X1_HVT U598 ( .A1(n383), .A2(conv_weight_box[28]), .A3(n382), .A4(
        conv_weight_box[188]), .Y(n378) );
  AO22X1_HVT U599 ( .A1(n385), .A2(conv_weight_box[140]), .A3(n384), .A4(
        conv_weight_box[156]), .Y(n376) );
  AO22X1_HVT U600 ( .A1(n387), .A2(conv_weight_box[108]), .A3(n386), .A4(
        conv_weight_box[60]), .Y(n375) );
  AO22X1_HVT U601 ( .A1(n389), .A2(conv_weight_box[92]), .A3(n388), .A4(
        conv_weight_box[124]), .Y(n374) );
  OR3X1_HVT U602 ( .A1(n376), .A2(n375), .A3(n374), .Y(n377) );
  OR3X1_HVT U603 ( .A1(n379), .A2(n378), .A3(n377), .Y(n398) );
  AO22X1_HVT U604 ( .A1(n381), .A2(conv_weight_box[40]), .A3(n380), .A4(
        conv_weight_box[168]), .Y(n395) );
  AO22X1_HVT U605 ( .A1(n383), .A2(conv_weight_box[24]), .A3(n382), .A4(
        conv_weight_box[184]), .Y(n394) );
  AO22X1_HVT U606 ( .A1(n385), .A2(conv_weight_box[136]), .A3(n384), .A4(
        conv_weight_box[152]), .Y(n392) );
  AO22X1_HVT U607 ( .A1(n387), .A2(conv_weight_box[104]), .A3(n386), .A4(
        conv_weight_box[56]), .Y(n391) );
  AO22X1_HVT U608 ( .A1(n389), .A2(conv_weight_box[88]), .A3(n388), .A4(
        conv_weight_box[120]), .Y(n390) );
  OR3X1_HVT U609 ( .A1(n392), .A2(n391), .A3(n390), .Y(n393) );
  OR3X1_HVT U610 ( .A1(n395), .A2(n394), .A3(n393), .Y(n396) );
  AOI22X1_HVT U611 ( .A1(n399), .A2(n398), .A3(n397), .A4(n396), .Y(n400) );
endmodule


module multiply_compare ( clk, srstn, mode, channel, conv1_sram_rdata_weight, 
        conv2_sram_rdata_weight, src_window, data_out );
  input [1:0] mode;
  input [4:0] channel;
  input [99:0] conv1_sram_rdata_weight;
  input [99:0] conv2_sram_rdata_weight;
  input [287:0] src_window;
  output [31:0] data_out;
  input clk, srstn;
  wire   N5, N7, DP_OP_425J2_127_3477_n3054, DP_OP_425J2_127_3477_n3017,
         DP_OP_425J2_127_3477_n3015, DP_OP_425J2_127_3477_n3014,
         DP_OP_425J2_127_3477_n3013, DP_OP_425J2_127_3477_n3012,
         DP_OP_425J2_127_3477_n3011, DP_OP_425J2_127_3477_n3010,
         DP_OP_425J2_127_3477_n3009, DP_OP_425J2_127_3477_n3008,
         DP_OP_425J2_127_3477_n3007, DP_OP_425J2_127_3477_n3006,
         DP_OP_425J2_127_3477_n3005, DP_OP_425J2_127_3477_n3004,
         DP_OP_425J2_127_3477_n3003, DP_OP_425J2_127_3477_n3002,
         DP_OP_425J2_127_3477_n3001, DP_OP_425J2_127_3477_n3000,
         DP_OP_425J2_127_3477_n2999, DP_OP_425J2_127_3477_n2998,
         DP_OP_425J2_127_3477_n2997, DP_OP_425J2_127_3477_n2996,
         DP_OP_425J2_127_3477_n2995, DP_OP_425J2_127_3477_n2994,
         DP_OP_425J2_127_3477_n2993, DP_OP_425J2_127_3477_n2992,
         DP_OP_425J2_127_3477_n2991, DP_OP_425J2_127_3477_n2990,
         DP_OP_425J2_127_3477_n2989, DP_OP_425J2_127_3477_n2988,
         DP_OP_425J2_127_3477_n2987, DP_OP_425J2_127_3477_n2986,
         DP_OP_425J2_127_3477_n2985, DP_OP_425J2_127_3477_n2984,
         DP_OP_425J2_127_3477_n2983, DP_OP_425J2_127_3477_n2982,
         DP_OP_425J2_127_3477_n2981, DP_OP_425J2_127_3477_n2980,
         DP_OP_425J2_127_3477_n2979, DP_OP_425J2_127_3477_n2978,
         DP_OP_425J2_127_3477_n2977, DP_OP_425J2_127_3477_n2976,
         DP_OP_425J2_127_3477_n2975, DP_OP_425J2_127_3477_n2974,
         DP_OP_425J2_127_3477_n2973, DP_OP_425J2_127_3477_n2972,
         DP_OP_425J2_127_3477_n2971, DP_OP_425J2_127_3477_n2967,
         DP_OP_425J2_127_3477_n2965, DP_OP_425J2_127_3477_n2964,
         DP_OP_425J2_127_3477_n2963, DP_OP_425J2_127_3477_n2962,
         DP_OP_425J2_127_3477_n2961, DP_OP_425J2_127_3477_n2960,
         DP_OP_425J2_127_3477_n2959, DP_OP_425J2_127_3477_n2958,
         DP_OP_425J2_127_3477_n2957, DP_OP_425J2_127_3477_n2956,
         DP_OP_425J2_127_3477_n2955, DP_OP_425J2_127_3477_n2954,
         DP_OP_425J2_127_3477_n2953, DP_OP_425J2_127_3477_n2952,
         DP_OP_425J2_127_3477_n2951, DP_OP_425J2_127_3477_n2950,
         DP_OP_425J2_127_3477_n2949, DP_OP_425J2_127_3477_n2948,
         DP_OP_425J2_127_3477_n2947, DP_OP_425J2_127_3477_n2946,
         DP_OP_425J2_127_3477_n2945, DP_OP_425J2_127_3477_n2944,
         DP_OP_425J2_127_3477_n2943, DP_OP_425J2_127_3477_n2942,
         DP_OP_425J2_127_3477_n2941, DP_OP_425J2_127_3477_n2940,
         DP_OP_425J2_127_3477_n2939, DP_OP_425J2_127_3477_n2938,
         DP_OP_425J2_127_3477_n2937, DP_OP_425J2_127_3477_n2936,
         DP_OP_425J2_127_3477_n2935, DP_OP_425J2_127_3477_n2934,
         DP_OP_425J2_127_3477_n2933, DP_OP_425J2_127_3477_n2932,
         DP_OP_425J2_127_3477_n2931, DP_OP_425J2_127_3477_n2930,
         DP_OP_425J2_127_3477_n2929, DP_OP_425J2_127_3477_n2928,
         DP_OP_425J2_127_3477_n2927, DP_OP_425J2_127_3477_n2926,
         DP_OP_425J2_127_3477_n2924, DP_OP_425J2_127_3477_n2923,
         DP_OP_425J2_127_3477_n2922, DP_OP_425J2_127_3477_n2921,
         DP_OP_425J2_127_3477_n2920, DP_OP_425J2_127_3477_n2919,
         DP_OP_425J2_127_3477_n2918, DP_OP_425J2_127_3477_n2917,
         DP_OP_425J2_127_3477_n2916, DP_OP_425J2_127_3477_n2915,
         DP_OP_425J2_127_3477_n2914, DP_OP_425J2_127_3477_n2913,
         DP_OP_425J2_127_3477_n2912, DP_OP_425J2_127_3477_n2911,
         DP_OP_425J2_127_3477_n2910, DP_OP_425J2_127_3477_n2909,
         DP_OP_425J2_127_3477_n2908, DP_OP_425J2_127_3477_n2907,
         DP_OP_425J2_127_3477_n2906, DP_OP_425J2_127_3477_n2905,
         DP_OP_425J2_127_3477_n2904, DP_OP_425J2_127_3477_n2903,
         DP_OP_425J2_127_3477_n2902, DP_OP_425J2_127_3477_n2901,
         DP_OP_425J2_127_3477_n2900, DP_OP_425J2_127_3477_n2899,
         DP_OP_425J2_127_3477_n2898, DP_OP_425J2_127_3477_n2897,
         DP_OP_425J2_127_3477_n2896, DP_OP_425J2_127_3477_n2895,
         DP_OP_425J2_127_3477_n2894, DP_OP_425J2_127_3477_n2893,
         DP_OP_425J2_127_3477_n2892, DP_OP_425J2_127_3477_n2891,
         DP_OP_425J2_127_3477_n2890, DP_OP_425J2_127_3477_n2889,
         DP_OP_425J2_127_3477_n2888, DP_OP_425J2_127_3477_n2887,
         DP_OP_425J2_127_3477_n2884, DP_OP_425J2_127_3477_n2879,
         DP_OP_425J2_127_3477_n2878, DP_OP_425J2_127_3477_n2877,
         DP_OP_425J2_127_3477_n2875, DP_OP_425J2_127_3477_n2874,
         DP_OP_425J2_127_3477_n2873, DP_OP_425J2_127_3477_n2872,
         DP_OP_425J2_127_3477_n2871, DP_OP_425J2_127_3477_n2870,
         DP_OP_425J2_127_3477_n2869, DP_OP_425J2_127_3477_n2868,
         DP_OP_425J2_127_3477_n2867, DP_OP_425J2_127_3477_n2866,
         DP_OP_425J2_127_3477_n2865, DP_OP_425J2_127_3477_n2864,
         DP_OP_425J2_127_3477_n2863, DP_OP_425J2_127_3477_n2862,
         DP_OP_425J2_127_3477_n2861, DP_OP_425J2_127_3477_n2860,
         DP_OP_425J2_127_3477_n2859, DP_OP_425J2_127_3477_n2858,
         DP_OP_425J2_127_3477_n2857, DP_OP_425J2_127_3477_n2856,
         DP_OP_425J2_127_3477_n2855, DP_OP_425J2_127_3477_n2854,
         DP_OP_425J2_127_3477_n2853, DP_OP_425J2_127_3477_n2852,
         DP_OP_425J2_127_3477_n2851, DP_OP_425J2_127_3477_n2850,
         DP_OP_425J2_127_3477_n2849, DP_OP_425J2_127_3477_n2848,
         DP_OP_425J2_127_3477_n2847, DP_OP_425J2_127_3477_n2846,
         DP_OP_425J2_127_3477_n2845, DP_OP_425J2_127_3477_n2844,
         DP_OP_425J2_127_3477_n2843, DP_OP_425J2_127_3477_n2842,
         DP_OP_425J2_127_3477_n2841, DP_OP_425J2_127_3477_n2840,
         DP_OP_425J2_127_3477_n2837, DP_OP_425J2_127_3477_n2835,
         DP_OP_425J2_127_3477_n2834, DP_OP_425J2_127_3477_n2833,
         DP_OP_425J2_127_3477_n2831, DP_OP_425J2_127_3477_n2830,
         DP_OP_425J2_127_3477_n2829, DP_OP_425J2_127_3477_n2828,
         DP_OP_425J2_127_3477_n2827, DP_OP_425J2_127_3477_n2826,
         DP_OP_425J2_127_3477_n2825, DP_OP_425J2_127_3477_n2824,
         DP_OP_425J2_127_3477_n2823, DP_OP_425J2_127_3477_n2822,
         DP_OP_425J2_127_3477_n2821, DP_OP_425J2_127_3477_n2820,
         DP_OP_425J2_127_3477_n2819, DP_OP_425J2_127_3477_n2818,
         DP_OP_425J2_127_3477_n2817, DP_OP_425J2_127_3477_n2816,
         DP_OP_425J2_127_3477_n2815, DP_OP_425J2_127_3477_n2814,
         DP_OP_425J2_127_3477_n2813, DP_OP_425J2_127_3477_n2812,
         DP_OP_425J2_127_3477_n2811, DP_OP_425J2_127_3477_n2810,
         DP_OP_425J2_127_3477_n2809, DP_OP_425J2_127_3477_n2808,
         DP_OP_425J2_127_3477_n2807, DP_OP_425J2_127_3477_n2806,
         DP_OP_425J2_127_3477_n2805, DP_OP_425J2_127_3477_n2804,
         DP_OP_425J2_127_3477_n2803, DP_OP_425J2_127_3477_n2802,
         DP_OP_425J2_127_3477_n2801, DP_OP_425J2_127_3477_n2800,
         DP_OP_425J2_127_3477_n2799, DP_OP_425J2_127_3477_n2798,
         DP_OP_425J2_127_3477_n2797, DP_OP_425J2_127_3477_n2796,
         DP_OP_425J2_127_3477_n2795, DP_OP_425J2_127_3477_n2794,
         DP_OP_425J2_127_3477_n2793, DP_OP_425J2_127_3477_n2791,
         DP_OP_425J2_127_3477_n2790, DP_OP_425J2_127_3477_n2789,
         DP_OP_425J2_127_3477_n2787, DP_OP_425J2_127_3477_n2786,
         DP_OP_425J2_127_3477_n2785, DP_OP_425J2_127_3477_n2784,
         DP_OP_425J2_127_3477_n2783, DP_OP_425J2_127_3477_n2782,
         DP_OP_425J2_127_3477_n2781, DP_OP_425J2_127_3477_n2780,
         DP_OP_425J2_127_3477_n2779, DP_OP_425J2_127_3477_n2778,
         DP_OP_425J2_127_3477_n2777, DP_OP_425J2_127_3477_n2776,
         DP_OP_425J2_127_3477_n2775, DP_OP_425J2_127_3477_n2774,
         DP_OP_425J2_127_3477_n2773, DP_OP_425J2_127_3477_n2772,
         DP_OP_425J2_127_3477_n2771, DP_OP_425J2_127_3477_n2770,
         DP_OP_425J2_127_3477_n2769, DP_OP_425J2_127_3477_n2768,
         DP_OP_425J2_127_3477_n2767, DP_OP_425J2_127_3477_n2766,
         DP_OP_425J2_127_3477_n2765, DP_OP_425J2_127_3477_n2764,
         DP_OP_425J2_127_3477_n2763, DP_OP_425J2_127_3477_n2762,
         DP_OP_425J2_127_3477_n2761, DP_OP_425J2_127_3477_n2760,
         DP_OP_425J2_127_3477_n2759, DP_OP_425J2_127_3477_n2758,
         DP_OP_425J2_127_3477_n2757, DP_OP_425J2_127_3477_n2756,
         DP_OP_425J2_127_3477_n2755, DP_OP_425J2_127_3477_n2754,
         DP_OP_425J2_127_3477_n2752, DP_OP_425J2_127_3477_n2750,
         DP_OP_425J2_127_3477_n2749, DP_OP_425J2_127_3477_n2747,
         DP_OP_425J2_127_3477_n2745, DP_OP_425J2_127_3477_n2743,
         DP_OP_425J2_127_3477_n2742, DP_OP_425J2_127_3477_n2741,
         DP_OP_425J2_127_3477_n2740, DP_OP_425J2_127_3477_n2739,
         DP_OP_425J2_127_3477_n2738, DP_OP_425J2_127_3477_n2737,
         DP_OP_425J2_127_3477_n2736, DP_OP_425J2_127_3477_n2735,
         DP_OP_425J2_127_3477_n2734, DP_OP_425J2_127_3477_n2733,
         DP_OP_425J2_127_3477_n2732, DP_OP_425J2_127_3477_n2731,
         DP_OP_425J2_127_3477_n2730, DP_OP_425J2_127_3477_n2729,
         DP_OP_425J2_127_3477_n2728, DP_OP_425J2_127_3477_n2727,
         DP_OP_425J2_127_3477_n2726, DP_OP_425J2_127_3477_n2725,
         DP_OP_425J2_127_3477_n2724, DP_OP_425J2_127_3477_n2723,
         DP_OP_425J2_127_3477_n2722, DP_OP_425J2_127_3477_n2721,
         DP_OP_425J2_127_3477_n2720, DP_OP_425J2_127_3477_n2719,
         DP_OP_425J2_127_3477_n2718, DP_OP_425J2_127_3477_n2717,
         DP_OP_425J2_127_3477_n2716, DP_OP_425J2_127_3477_n2715,
         DP_OP_425J2_127_3477_n2714, DP_OP_425J2_127_3477_n2713,
         DP_OP_425J2_127_3477_n2712, DP_OP_425J2_127_3477_n2711,
         DP_OP_425J2_127_3477_n2710, DP_OP_425J2_127_3477_n2709,
         DP_OP_425J2_127_3477_n2708, DP_OP_425J2_127_3477_n2707,
         DP_OP_425J2_127_3477_n2705, DP_OP_425J2_127_3477_n2704,
         DP_OP_425J2_127_3477_n2700, DP_OP_425J2_127_3477_n2699,
         DP_OP_425J2_127_3477_n2698, DP_OP_425J2_127_3477_n2697,
         DP_OP_425J2_127_3477_n2696, DP_OP_425J2_127_3477_n2695,
         DP_OP_425J2_127_3477_n2694, DP_OP_425J2_127_3477_n2693,
         DP_OP_425J2_127_3477_n2692, DP_OP_425J2_127_3477_n2691,
         DP_OP_425J2_127_3477_n2690, DP_OP_425J2_127_3477_n2689,
         DP_OP_425J2_127_3477_n2688, DP_OP_425J2_127_3477_n2687,
         DP_OP_425J2_127_3477_n2686, DP_OP_425J2_127_3477_n2685,
         DP_OP_425J2_127_3477_n2684, DP_OP_425J2_127_3477_n2683,
         DP_OP_425J2_127_3477_n2682, DP_OP_425J2_127_3477_n2681,
         DP_OP_425J2_127_3477_n2680, DP_OP_425J2_127_3477_n2679,
         DP_OP_425J2_127_3477_n2678, DP_OP_425J2_127_3477_n2677,
         DP_OP_425J2_127_3477_n2676, DP_OP_425J2_127_3477_n2675,
         DP_OP_425J2_127_3477_n2674, DP_OP_425J2_127_3477_n2673,
         DP_OP_425J2_127_3477_n2672, DP_OP_425J2_127_3477_n2671,
         DP_OP_425J2_127_3477_n2670, DP_OP_425J2_127_3477_n2669,
         DP_OP_425J2_127_3477_n2668, DP_OP_425J2_127_3477_n2667,
         DP_OP_425J2_127_3477_n2666, DP_OP_425J2_127_3477_n2665,
         DP_OP_425J2_127_3477_n2664, DP_OP_425J2_127_3477_n2663,
         DP_OP_425J2_127_3477_n2662, DP_OP_425J2_127_3477_n2658,
         DP_OP_425J2_127_3477_n2655, DP_OP_425J2_127_3477_n2654,
         DP_OP_425J2_127_3477_n2653, DP_OP_425J2_127_3477_n2652,
         DP_OP_425J2_127_3477_n2651, DP_OP_425J2_127_3477_n2650,
         DP_OP_425J2_127_3477_n2649, DP_OP_425J2_127_3477_n2648,
         DP_OP_425J2_127_3477_n2647, DP_OP_425J2_127_3477_n2646,
         DP_OP_425J2_127_3477_n2645, DP_OP_425J2_127_3477_n2644,
         DP_OP_425J2_127_3477_n2643, DP_OP_425J2_127_3477_n2642,
         DP_OP_425J2_127_3477_n2641, DP_OP_425J2_127_3477_n2640,
         DP_OP_425J2_127_3477_n2639, DP_OP_425J2_127_3477_n2638,
         DP_OP_425J2_127_3477_n2637, DP_OP_425J2_127_3477_n2636,
         DP_OP_425J2_127_3477_n2635, DP_OP_425J2_127_3477_n2634,
         DP_OP_425J2_127_3477_n2633, DP_OP_425J2_127_3477_n2632,
         DP_OP_425J2_127_3477_n2631, DP_OP_425J2_127_3477_n2630,
         DP_OP_425J2_127_3477_n2629, DP_OP_425J2_127_3477_n2628,
         DP_OP_425J2_127_3477_n2627, DP_OP_425J2_127_3477_n2626,
         DP_OP_425J2_127_3477_n2625, DP_OP_425J2_127_3477_n2624,
         DP_OP_425J2_127_3477_n2623, DP_OP_425J2_127_3477_n2622,
         DP_OP_425J2_127_3477_n2621, DP_OP_425J2_127_3477_n2620,
         DP_OP_425J2_127_3477_n2619, DP_OP_425J2_127_3477_n2617,
         DP_OP_425J2_127_3477_n2616, DP_OP_425J2_127_3477_n2612,
         DP_OP_425J2_127_3477_n2611, DP_OP_425J2_127_3477_n2610,
         DP_OP_425J2_127_3477_n2609, DP_OP_425J2_127_3477_n2608,
         DP_OP_425J2_127_3477_n2607, DP_OP_425J2_127_3477_n2606,
         DP_OP_425J2_127_3477_n2605, DP_OP_425J2_127_3477_n2604,
         DP_OP_425J2_127_3477_n2603, DP_OP_425J2_127_3477_n2602,
         DP_OP_425J2_127_3477_n2601, DP_OP_425J2_127_3477_n2600,
         DP_OP_425J2_127_3477_n2599, DP_OP_425J2_127_3477_n2598,
         DP_OP_425J2_127_3477_n2597, DP_OP_425J2_127_3477_n2596,
         DP_OP_425J2_127_3477_n2595, DP_OP_425J2_127_3477_n2594,
         DP_OP_425J2_127_3477_n2593, DP_OP_425J2_127_3477_n2592,
         DP_OP_425J2_127_3477_n2591, DP_OP_425J2_127_3477_n2590,
         DP_OP_425J2_127_3477_n2589, DP_OP_425J2_127_3477_n2588,
         DP_OP_425J2_127_3477_n2587, DP_OP_425J2_127_3477_n2586,
         DP_OP_425J2_127_3477_n2585, DP_OP_425J2_127_3477_n2584,
         DP_OP_425J2_127_3477_n2583, DP_OP_425J2_127_3477_n2582,
         DP_OP_425J2_127_3477_n2581, DP_OP_425J2_127_3477_n2580,
         DP_OP_425J2_127_3477_n2579, DP_OP_425J2_127_3477_n2578,
         DP_OP_425J2_127_3477_n2577, DP_OP_425J2_127_3477_n2576,
         DP_OP_425J2_127_3477_n2572, DP_OP_425J2_127_3477_n2567,
         DP_OP_425J2_127_3477_n2566, DP_OP_425J2_127_3477_n2565,
         DP_OP_425J2_127_3477_n2564, DP_OP_425J2_127_3477_n2563,
         DP_OP_425J2_127_3477_n2562, DP_OP_425J2_127_3477_n2561,
         DP_OP_425J2_127_3477_n2560, DP_OP_425J2_127_3477_n2559,
         DP_OP_425J2_127_3477_n2558, DP_OP_425J2_127_3477_n2557,
         DP_OP_425J2_127_3477_n2556, DP_OP_425J2_127_3477_n2555,
         DP_OP_425J2_127_3477_n2554, DP_OP_425J2_127_3477_n2553,
         DP_OP_425J2_127_3477_n2552, DP_OP_425J2_127_3477_n2551,
         DP_OP_425J2_127_3477_n2550, DP_OP_425J2_127_3477_n2549,
         DP_OP_425J2_127_3477_n2548, DP_OP_425J2_127_3477_n2547,
         DP_OP_425J2_127_3477_n2546, DP_OP_425J2_127_3477_n2545,
         DP_OP_425J2_127_3477_n2544, DP_OP_425J2_127_3477_n2543,
         DP_OP_425J2_127_3477_n2542, DP_OP_425J2_127_3477_n2541,
         DP_OP_425J2_127_3477_n2540, DP_OP_425J2_127_3477_n2539,
         DP_OP_425J2_127_3477_n2538, DP_OP_425J2_127_3477_n2537,
         DP_OP_425J2_127_3477_n2536, DP_OP_425J2_127_3477_n2535,
         DP_OP_425J2_127_3477_n2534, DP_OP_425J2_127_3477_n2530,
         DP_OP_425J2_127_3477_n2529, DP_OP_425J2_127_3477_n2528,
         DP_OP_425J2_127_3477_n2526, DP_OP_425J2_127_3477_n2525,
         DP_OP_425J2_127_3477_n2523, DP_OP_425J2_127_3477_n2522,
         DP_OP_425J2_127_3477_n2521, DP_OP_425J2_127_3477_n2520,
         DP_OP_425J2_127_3477_n2519, DP_OP_425J2_127_3477_n2518,
         DP_OP_425J2_127_3477_n2517, DP_OP_425J2_127_3477_n2516,
         DP_OP_425J2_127_3477_n2515, DP_OP_425J2_127_3477_n2514,
         DP_OP_425J2_127_3477_n2513, DP_OP_425J2_127_3477_n2512,
         DP_OP_425J2_127_3477_n2511, DP_OP_425J2_127_3477_n2510,
         DP_OP_425J2_127_3477_n2509, DP_OP_425J2_127_3477_n2508,
         DP_OP_425J2_127_3477_n2507, DP_OP_425J2_127_3477_n2506,
         DP_OP_425J2_127_3477_n2505, DP_OP_425J2_127_3477_n2504,
         DP_OP_425J2_127_3477_n2503, DP_OP_425J2_127_3477_n2502,
         DP_OP_425J2_127_3477_n2501, DP_OP_425J2_127_3477_n2500,
         DP_OP_425J2_127_3477_n2499, DP_OP_425J2_127_3477_n2498,
         DP_OP_425J2_127_3477_n2497, DP_OP_425J2_127_3477_n2496,
         DP_OP_425J2_127_3477_n2495, DP_OP_425J2_127_3477_n2494,
         DP_OP_425J2_127_3477_n2493, DP_OP_425J2_127_3477_n2492,
         DP_OP_425J2_127_3477_n2491, DP_OP_425J2_127_3477_n2490,
         DP_OP_425J2_127_3477_n2489, DP_OP_425J2_127_3477_n2488,
         DP_OP_425J2_127_3477_n2484, DP_OP_425J2_127_3477_n2482,
         DP_OP_425J2_127_3477_n2481, DP_OP_425J2_127_3477_n2479,
         DP_OP_425J2_127_3477_n2478, DP_OP_425J2_127_3477_n2477,
         DP_OP_425J2_127_3477_n2476, DP_OP_425J2_127_3477_n2475,
         DP_OP_425J2_127_3477_n2474, DP_OP_425J2_127_3477_n2473,
         DP_OP_425J2_127_3477_n2472, DP_OP_425J2_127_3477_n2471,
         DP_OP_425J2_127_3477_n2470, DP_OP_425J2_127_3477_n2469,
         DP_OP_425J2_127_3477_n2468, DP_OP_425J2_127_3477_n2467,
         DP_OP_425J2_127_3477_n2466, DP_OP_425J2_127_3477_n2465,
         DP_OP_425J2_127_3477_n2464, DP_OP_425J2_127_3477_n2463,
         DP_OP_425J2_127_3477_n2462, DP_OP_425J2_127_3477_n2461,
         DP_OP_425J2_127_3477_n2460, DP_OP_425J2_127_3477_n2459,
         DP_OP_425J2_127_3477_n2458, DP_OP_425J2_127_3477_n2457,
         DP_OP_425J2_127_3477_n2456, DP_OP_425J2_127_3477_n2455,
         DP_OP_425J2_127_3477_n2454, DP_OP_425J2_127_3477_n2453,
         DP_OP_425J2_127_3477_n2452, DP_OP_425J2_127_3477_n2451,
         DP_OP_425J2_127_3477_n2450, DP_OP_425J2_127_3477_n2449,
         DP_OP_425J2_127_3477_n2448, DP_OP_425J2_127_3477_n2447,
         DP_OP_425J2_127_3477_n2446, DP_OP_425J2_127_3477_n2445,
         DP_OP_425J2_127_3477_n2442, DP_OP_425J2_127_3477_n2441,
         DP_OP_425J2_127_3477_n2439, DP_OP_425J2_127_3477_n2438,
         DP_OP_425J2_127_3477_n2435, DP_OP_425J2_127_3477_n2434,
         DP_OP_425J2_127_3477_n2433, DP_OP_425J2_127_3477_n2432,
         DP_OP_425J2_127_3477_n2431, DP_OP_425J2_127_3477_n2430,
         DP_OP_425J2_127_3477_n2429, DP_OP_425J2_127_3477_n2428,
         DP_OP_425J2_127_3477_n2427, DP_OP_425J2_127_3477_n2426,
         DP_OP_425J2_127_3477_n2425, DP_OP_425J2_127_3477_n2424,
         DP_OP_425J2_127_3477_n2423, DP_OP_425J2_127_3477_n2422,
         DP_OP_425J2_127_3477_n2421, DP_OP_425J2_127_3477_n2420,
         DP_OP_425J2_127_3477_n2419, DP_OP_425J2_127_3477_n2418,
         DP_OP_425J2_127_3477_n2417, DP_OP_425J2_127_3477_n2416,
         DP_OP_425J2_127_3477_n2415, DP_OP_425J2_127_3477_n2414,
         DP_OP_425J2_127_3477_n2413, DP_OP_425J2_127_3477_n2412,
         DP_OP_425J2_127_3477_n2411, DP_OP_425J2_127_3477_n2410,
         DP_OP_425J2_127_3477_n2409, DP_OP_425J2_127_3477_n2408,
         DP_OP_425J2_127_3477_n2407, DP_OP_425J2_127_3477_n2406,
         DP_OP_425J2_127_3477_n2405, DP_OP_425J2_127_3477_n2404,
         DP_OP_425J2_127_3477_n2403, DP_OP_425J2_127_3477_n2402,
         DP_OP_425J2_127_3477_n2401, DP_OP_425J2_127_3477_n2400,
         DP_OP_425J2_127_3477_n2398, DP_OP_425J2_127_3477_n2397,
         DP_OP_425J2_127_3477_n2396, DP_OP_425J2_127_3477_n2391,
         DP_OP_425J2_127_3477_n2390, DP_OP_425J2_127_3477_n2389,
         DP_OP_425J2_127_3477_n2388, DP_OP_425J2_127_3477_n2387,
         DP_OP_425J2_127_3477_n2386, DP_OP_425J2_127_3477_n2385,
         DP_OP_425J2_127_3477_n2384, DP_OP_425J2_127_3477_n2383,
         DP_OP_425J2_127_3477_n2382, DP_OP_425J2_127_3477_n2381,
         DP_OP_425J2_127_3477_n2380, DP_OP_425J2_127_3477_n2379,
         DP_OP_425J2_127_3477_n2378, DP_OP_425J2_127_3477_n2377,
         DP_OP_425J2_127_3477_n2376, DP_OP_425J2_127_3477_n2375,
         DP_OP_425J2_127_3477_n2374, DP_OP_425J2_127_3477_n2373,
         DP_OP_425J2_127_3477_n2372, DP_OP_425J2_127_3477_n2371,
         DP_OP_425J2_127_3477_n2370, DP_OP_425J2_127_3477_n2369,
         DP_OP_425J2_127_3477_n2368, DP_OP_425J2_127_3477_n2367,
         DP_OP_425J2_127_3477_n2366, DP_OP_425J2_127_3477_n2365,
         DP_OP_425J2_127_3477_n2364, DP_OP_425J2_127_3477_n2363,
         DP_OP_425J2_127_3477_n2362, DP_OP_425J2_127_3477_n2361,
         DP_OP_425J2_127_3477_n2360, DP_OP_425J2_127_3477_n2359,
         DP_OP_425J2_127_3477_n2358, DP_OP_425J2_127_3477_n2357,
         DP_OP_425J2_127_3477_n2356, DP_OP_425J2_127_3477_n2355,
         DP_OP_425J2_127_3477_n2354, DP_OP_425J2_127_3477_n2353,
         DP_OP_425J2_127_3477_n2351, DP_OP_425J2_127_3477_n2347,
         DP_OP_425J2_127_3477_n2346, DP_OP_425J2_127_3477_n2345,
         DP_OP_425J2_127_3477_n2344, DP_OP_425J2_127_3477_n2343,
         DP_OP_425J2_127_3477_n2342, DP_OP_425J2_127_3477_n2341,
         DP_OP_425J2_127_3477_n2340, DP_OP_425J2_127_3477_n2339,
         DP_OP_425J2_127_3477_n2338, DP_OP_425J2_127_3477_n2337,
         DP_OP_425J2_127_3477_n2336, DP_OP_425J2_127_3477_n2335,
         DP_OP_425J2_127_3477_n2334, DP_OP_425J2_127_3477_n2333,
         DP_OP_425J2_127_3477_n2332, DP_OP_425J2_127_3477_n2331,
         DP_OP_425J2_127_3477_n2330, DP_OP_425J2_127_3477_n2329,
         DP_OP_425J2_127_3477_n2328, DP_OP_425J2_127_3477_n2327,
         DP_OP_425J2_127_3477_n2326, DP_OP_425J2_127_3477_n2325,
         DP_OP_425J2_127_3477_n2324, DP_OP_425J2_127_3477_n2323,
         DP_OP_425J2_127_3477_n2322, DP_OP_425J2_127_3477_n2321,
         DP_OP_425J2_127_3477_n2320, DP_OP_425J2_127_3477_n2319,
         DP_OP_425J2_127_3477_n2318, DP_OP_425J2_127_3477_n2317,
         DP_OP_425J2_127_3477_n2316, DP_OP_425J2_127_3477_n2315,
         DP_OP_425J2_127_3477_n2314, DP_OP_425J2_127_3477_n2313,
         DP_OP_425J2_127_3477_n2312, DP_OP_425J2_127_3477_n2308,
         DP_OP_425J2_127_3477_n2307, DP_OP_425J2_127_3477_n2305,
         DP_OP_425J2_127_3477_n2304, DP_OP_425J2_127_3477_n2303,
         DP_OP_425J2_127_3477_n2302, DP_OP_425J2_127_3477_n2301,
         DP_OP_425J2_127_3477_n2300, DP_OP_425J2_127_3477_n2299,
         DP_OP_425J2_127_3477_n2298, DP_OP_425J2_127_3477_n2297,
         DP_OP_425J2_127_3477_n2296, DP_OP_425J2_127_3477_n2295,
         DP_OP_425J2_127_3477_n2294, DP_OP_425J2_127_3477_n2293,
         DP_OP_425J2_127_3477_n2292, DP_OP_425J2_127_3477_n2291,
         DP_OP_425J2_127_3477_n2290, DP_OP_425J2_127_3477_n2289,
         DP_OP_425J2_127_3477_n2288, DP_OP_425J2_127_3477_n2287,
         DP_OP_425J2_127_3477_n2286, DP_OP_425J2_127_3477_n2285,
         DP_OP_425J2_127_3477_n2284, DP_OP_425J2_127_3477_n2283,
         DP_OP_425J2_127_3477_n2282, DP_OP_425J2_127_3477_n2281,
         DP_OP_425J2_127_3477_n2280, DP_OP_425J2_127_3477_n2279,
         DP_OP_425J2_127_3477_n2278, DP_OP_425J2_127_3477_n2277,
         DP_OP_425J2_127_3477_n2276, DP_OP_425J2_127_3477_n2275,
         DP_OP_425J2_127_3477_n2274, DP_OP_425J2_127_3477_n2273,
         DP_OP_425J2_127_3477_n2272, DP_OP_425J2_127_3477_n2271,
         DP_OP_425J2_127_3477_n2270, DP_OP_425J2_127_3477_n2269,
         DP_OP_425J2_127_3477_n2268, DP_OP_425J2_127_3477_n2264,
         DP_OP_425J2_127_3477_n2261, DP_OP_425J2_127_3477_n2260,
         DP_OP_425J2_127_3477_n2259, DP_OP_425J2_127_3477_n2258,
         DP_OP_425J2_127_3477_n2257, DP_OP_425J2_127_3477_n2256,
         DP_OP_425J2_127_3477_n2255, DP_OP_425J2_127_3477_n2254,
         DP_OP_425J2_127_3477_n2253, DP_OP_425J2_127_3477_n2252,
         DP_OP_425J2_127_3477_n2251, DP_OP_425J2_127_3477_n2250,
         DP_OP_425J2_127_3477_n2249, DP_OP_425J2_127_3477_n2248,
         DP_OP_425J2_127_3477_n2247, DP_OP_425J2_127_3477_n2246,
         DP_OP_425J2_127_3477_n2245, DP_OP_425J2_127_3477_n2244,
         DP_OP_425J2_127_3477_n2243, DP_OP_425J2_127_3477_n2242,
         DP_OP_425J2_127_3477_n2241, DP_OP_425J2_127_3477_n2240,
         DP_OP_425J2_127_3477_n2239, DP_OP_425J2_127_3477_n2238,
         DP_OP_425J2_127_3477_n2237, DP_OP_425J2_127_3477_n2236,
         DP_OP_425J2_127_3477_n2235, DP_OP_425J2_127_3477_n2234,
         DP_OP_425J2_127_3477_n2233, DP_OP_425J2_127_3477_n2232,
         DP_OP_425J2_127_3477_n2231, DP_OP_425J2_127_3477_n2230,
         DP_OP_425J2_127_3477_n2229, DP_OP_425J2_127_3477_n2228,
         DP_OP_425J2_127_3477_n2227, DP_OP_425J2_127_3477_n2226,
         DP_OP_425J2_127_3477_n2224, DP_OP_425J2_127_3477_n2220,
         DP_OP_425J2_127_3477_n2219, DP_OP_425J2_127_3477_n2218,
         DP_OP_425J2_127_3477_n2217, DP_OP_425J2_127_3477_n2216,
         DP_OP_425J2_127_3477_n2215, DP_OP_425J2_127_3477_n2214,
         DP_OP_425J2_127_3477_n2213, DP_OP_425J2_127_3477_n2212,
         DP_OP_425J2_127_3477_n2211, DP_OP_425J2_127_3477_n2210,
         DP_OP_425J2_127_3477_n2209, DP_OP_425J2_127_3477_n2208,
         DP_OP_425J2_127_3477_n2207, DP_OP_425J2_127_3477_n2206,
         DP_OP_425J2_127_3477_n2205, DP_OP_425J2_127_3477_n2204,
         DP_OP_425J2_127_3477_n2203, DP_OP_425J2_127_3477_n2202,
         DP_OP_425J2_127_3477_n2201, DP_OP_425J2_127_3477_n2200,
         DP_OP_425J2_127_3477_n2199, DP_OP_425J2_127_3477_n2198,
         DP_OP_425J2_127_3477_n2197, DP_OP_425J2_127_3477_n2196,
         DP_OP_425J2_127_3477_n2195, DP_OP_425J2_127_3477_n2194,
         DP_OP_425J2_127_3477_n2193, DP_OP_425J2_127_3477_n2192,
         DP_OP_425J2_127_3477_n2191, DP_OP_425J2_127_3477_n2190,
         DP_OP_425J2_127_3477_n2189, DP_OP_425J2_127_3477_n2188,
         DP_OP_425J2_127_3477_n2187, DP_OP_425J2_127_3477_n2186,
         DP_OP_425J2_127_3477_n2185, DP_OP_425J2_127_3477_n2184,
         DP_OP_425J2_127_3477_n2182, DP_OP_425J2_127_3477_n2181,
         DP_OP_425J2_127_3477_n2180, DP_OP_425J2_127_3477_n2178,
         DP_OP_425J2_127_3477_n2175, DP_OP_425J2_127_3477_n2172,
         DP_OP_425J2_127_3477_n2171, DP_OP_425J2_127_3477_n2170,
         DP_OP_425J2_127_3477_n2169, DP_OP_425J2_127_3477_n2168,
         DP_OP_425J2_127_3477_n2167, DP_OP_425J2_127_3477_n2166,
         DP_OP_425J2_127_3477_n2165, DP_OP_425J2_127_3477_n2164,
         DP_OP_425J2_127_3477_n2163, DP_OP_425J2_127_3477_n2162,
         DP_OP_425J2_127_3477_n2161, DP_OP_425J2_127_3477_n2160,
         DP_OP_425J2_127_3477_n2159, DP_OP_425J2_127_3477_n2158,
         DP_OP_425J2_127_3477_n2157, DP_OP_425J2_127_3477_n2156,
         DP_OP_425J2_127_3477_n2155, DP_OP_425J2_127_3477_n2154,
         DP_OP_425J2_127_3477_n2153, DP_OP_425J2_127_3477_n2152,
         DP_OP_425J2_127_3477_n2151, DP_OP_425J2_127_3477_n2150,
         DP_OP_425J2_127_3477_n2149, DP_OP_425J2_127_3477_n2148,
         DP_OP_425J2_127_3477_n2147, DP_OP_425J2_127_3477_n2146,
         DP_OP_425J2_127_3477_n2145, DP_OP_425J2_127_3477_n2144,
         DP_OP_425J2_127_3477_n2143, DP_OP_425J2_127_3477_n2142,
         DP_OP_425J2_127_3477_n2141, DP_OP_425J2_127_3477_n2140,
         DP_OP_425J2_127_3477_n2139, DP_OP_425J2_127_3477_n2138,
         DP_OP_425J2_127_3477_n2137, DP_OP_425J2_127_3477_n2136,
         DP_OP_425J2_127_3477_n2135, DP_OP_425J2_127_3477_n2134,
         DP_OP_425J2_127_3477_n2133, DP_OP_425J2_127_3477_n2128,
         DP_OP_425J2_127_3477_n2127, DP_OP_425J2_127_3477_n2126,
         DP_OP_425J2_127_3477_n2125, DP_OP_425J2_127_3477_n2124,
         DP_OP_425J2_127_3477_n2123, DP_OP_425J2_127_3477_n2122,
         DP_OP_425J2_127_3477_n2121, DP_OP_425J2_127_3477_n2120,
         DP_OP_425J2_127_3477_n2119, DP_OP_425J2_127_3477_n2118,
         DP_OP_425J2_127_3477_n2117, DP_OP_425J2_127_3477_n2116,
         DP_OP_425J2_127_3477_n2115, DP_OP_425J2_127_3477_n2114,
         DP_OP_425J2_127_3477_n2113, DP_OP_425J2_127_3477_n2112,
         DP_OP_425J2_127_3477_n2111, DP_OP_425J2_127_3477_n2110,
         DP_OP_425J2_127_3477_n2109, DP_OP_425J2_127_3477_n2108,
         DP_OP_425J2_127_3477_n2107, DP_OP_425J2_127_3477_n2106,
         DP_OP_425J2_127_3477_n2105, DP_OP_425J2_127_3477_n2104,
         DP_OP_425J2_127_3477_n2103, DP_OP_425J2_127_3477_n2102,
         DP_OP_425J2_127_3477_n2101, DP_OP_425J2_127_3477_n2100,
         DP_OP_425J2_127_3477_n2099, DP_OP_425J2_127_3477_n2098,
         DP_OP_425J2_127_3477_n2097, DP_OP_425J2_127_3477_n2096,
         DP_OP_425J2_127_3477_n2095, DP_OP_425J2_127_3477_n2094,
         DP_OP_425J2_127_3477_n2093, DP_OP_425J2_127_3477_n2092,
         DP_OP_425J2_127_3477_n2088, DP_OP_425J2_127_3477_n2087,
         DP_OP_425J2_127_3477_n2086, DP_OP_425J2_127_3477_n2085,
         DP_OP_425J2_127_3477_n2084, DP_OP_425J2_127_3477_n2083,
         DP_OP_425J2_127_3477_n2082, DP_OP_425J2_127_3477_n2081,
         DP_OP_425J2_127_3477_n2080, DP_OP_425J2_127_3477_n2079,
         DP_OP_425J2_127_3477_n2078, DP_OP_425J2_127_3477_n2077,
         DP_OP_425J2_127_3477_n2076, DP_OP_425J2_127_3477_n2075,
         DP_OP_425J2_127_3477_n2074, DP_OP_425J2_127_3477_n2073,
         DP_OP_425J2_127_3477_n2072, DP_OP_425J2_127_3477_n2071,
         DP_OP_425J2_127_3477_n2070, DP_OP_425J2_127_3477_n2069,
         DP_OP_425J2_127_3477_n2068, DP_OP_425J2_127_3477_n2067,
         DP_OP_425J2_127_3477_n2066, DP_OP_425J2_127_3477_n2065,
         DP_OP_425J2_127_3477_n2064, DP_OP_425J2_127_3477_n2063,
         DP_OP_425J2_127_3477_n2062, DP_OP_425J2_127_3477_n2061,
         DP_OP_425J2_127_3477_n2060, DP_OP_425J2_127_3477_n2059,
         DP_OP_425J2_127_3477_n2058, DP_OP_425J2_127_3477_n2057,
         DP_OP_425J2_127_3477_n2056, DP_OP_425J2_127_3477_n2055,
         DP_OP_425J2_127_3477_n2054, DP_OP_425J2_127_3477_n2053,
         DP_OP_425J2_127_3477_n2052, DP_OP_425J2_127_3477_n2051,
         DP_OP_425J2_127_3477_n2050, DP_OP_425J2_127_3477_n2049,
         DP_OP_425J2_127_3477_n2048, DP_OP_425J2_127_3477_n2047,
         DP_OP_425J2_127_3477_n2039, DP_OP_425J2_127_3477_n2038,
         DP_OP_425J2_127_3477_n2037, DP_OP_425J2_127_3477_n2036,
         DP_OP_425J2_127_3477_n2035, DP_OP_425J2_127_3477_n2034,
         DP_OP_425J2_127_3477_n2033, DP_OP_425J2_127_3477_n2032,
         DP_OP_425J2_127_3477_n2031, DP_OP_425J2_127_3477_n2030,
         DP_OP_425J2_127_3477_n2029, DP_OP_425J2_127_3477_n2028,
         DP_OP_425J2_127_3477_n2027, DP_OP_425J2_127_3477_n2026,
         DP_OP_425J2_127_3477_n2025, DP_OP_425J2_127_3477_n2024,
         DP_OP_425J2_127_3477_n2023, DP_OP_425J2_127_3477_n2022,
         DP_OP_425J2_127_3477_n2021, DP_OP_425J2_127_3477_n2020,
         DP_OP_425J2_127_3477_n2019, DP_OP_425J2_127_3477_n2018,
         DP_OP_425J2_127_3477_n2017, DP_OP_425J2_127_3477_n2016,
         DP_OP_425J2_127_3477_n2015, DP_OP_425J2_127_3477_n2014,
         DP_OP_425J2_127_3477_n2013, DP_OP_425J2_127_3477_n2012,
         DP_OP_425J2_127_3477_n2011, DP_OP_425J2_127_3477_n2010,
         DP_OP_425J2_127_3477_n2009, DP_OP_425J2_127_3477_n2008,
         DP_OP_425J2_127_3477_n2007, DP_OP_425J2_127_3477_n2006,
         DP_OP_425J2_127_3477_n2005, DP_OP_425J2_127_3477_n2004,
         DP_OP_425J2_127_3477_n2003, DP_OP_425J2_127_3477_n2000,
         DP_OP_425J2_127_3477_n1998, DP_OP_425J2_127_3477_n1997,
         DP_OP_425J2_127_3477_n1995, DP_OP_425J2_127_3477_n1994,
         DP_OP_425J2_127_3477_n1993, DP_OP_425J2_127_3477_n1992,
         DP_OP_425J2_127_3477_n1991, DP_OP_425J2_127_3477_n1990,
         DP_OP_425J2_127_3477_n1989, DP_OP_425J2_127_3477_n1988,
         DP_OP_425J2_127_3477_n1987, DP_OP_425J2_127_3477_n1986,
         DP_OP_425J2_127_3477_n1985, DP_OP_425J2_127_3477_n1984,
         DP_OP_425J2_127_3477_n1983, DP_OP_425J2_127_3477_n1982,
         DP_OP_425J2_127_3477_n1981, DP_OP_425J2_127_3477_n1980,
         DP_OP_425J2_127_3477_n1979, DP_OP_425J2_127_3477_n1978,
         DP_OP_425J2_127_3477_n1977, DP_OP_425J2_127_3477_n1976,
         DP_OP_425J2_127_3477_n1975, DP_OP_425J2_127_3477_n1974,
         DP_OP_425J2_127_3477_n1973, DP_OP_425J2_127_3477_n1972,
         DP_OP_425J2_127_3477_n1971, DP_OP_425J2_127_3477_n1970,
         DP_OP_425J2_127_3477_n1969, DP_OP_425J2_127_3477_n1968,
         DP_OP_425J2_127_3477_n1967, DP_OP_425J2_127_3477_n1966,
         DP_OP_425J2_127_3477_n1965, DP_OP_425J2_127_3477_n1964,
         DP_OP_425J2_127_3477_n1963, DP_OP_425J2_127_3477_n1961,
         DP_OP_425J2_127_3477_n1960, DP_OP_425J2_127_3477_n1951,
         DP_OP_425J2_127_3477_n1950, DP_OP_425J2_127_3477_n1949,
         DP_OP_425J2_127_3477_n1948, DP_OP_425J2_127_3477_n1947,
         DP_OP_425J2_127_3477_n1946, DP_OP_425J2_127_3477_n1945,
         DP_OP_425J2_127_3477_n1944, DP_OP_425J2_127_3477_n1943,
         DP_OP_425J2_127_3477_n1942, DP_OP_425J2_127_3477_n1941,
         DP_OP_425J2_127_3477_n1940, DP_OP_425J2_127_3477_n1939,
         DP_OP_425J2_127_3477_n1938, DP_OP_425J2_127_3477_n1937,
         DP_OP_425J2_127_3477_n1936, DP_OP_425J2_127_3477_n1935,
         DP_OP_425J2_127_3477_n1934, DP_OP_425J2_127_3477_n1933,
         DP_OP_425J2_127_3477_n1932, DP_OP_425J2_127_3477_n1931,
         DP_OP_425J2_127_3477_n1930, DP_OP_425J2_127_3477_n1929,
         DP_OP_425J2_127_3477_n1928, DP_OP_425J2_127_3477_n1927,
         DP_OP_425J2_127_3477_n1926, DP_OP_425J2_127_3477_n1925,
         DP_OP_425J2_127_3477_n1924, DP_OP_425J2_127_3477_n1923,
         DP_OP_425J2_127_3477_n1922, DP_OP_425J2_127_3477_n1921,
         DP_OP_425J2_127_3477_n1920, DP_OP_425J2_127_3477_n1886,
         DP_OP_425J2_127_3477_n1885, DP_OP_425J2_127_3477_n1884,
         DP_OP_425J2_127_3477_n1883, DP_OP_425J2_127_3477_n1882,
         DP_OP_425J2_127_3477_n1881, DP_OP_425J2_127_3477_n1880,
         DP_OP_425J2_127_3477_n1879, DP_OP_425J2_127_3477_n1878,
         DP_OP_425J2_127_3477_n1877, DP_OP_425J2_127_3477_n1876,
         DP_OP_425J2_127_3477_n1875, DP_OP_425J2_127_3477_n1874,
         DP_OP_425J2_127_3477_n1873, DP_OP_425J2_127_3477_n1871,
         DP_OP_425J2_127_3477_n1870, DP_OP_425J2_127_3477_n1869,
         DP_OP_425J2_127_3477_n1868, DP_OP_425J2_127_3477_n1867,
         DP_OP_425J2_127_3477_n1866, DP_OP_425J2_127_3477_n1865,
         DP_OP_425J2_127_3477_n1864, DP_OP_425J2_127_3477_n1863,
         DP_OP_425J2_127_3477_n1862, DP_OP_425J2_127_3477_n1861,
         DP_OP_425J2_127_3477_n1860, DP_OP_425J2_127_3477_n1859,
         DP_OP_425J2_127_3477_n1858, DP_OP_425J2_127_3477_n1857,
         DP_OP_425J2_127_3477_n1856, DP_OP_425J2_127_3477_n1855,
         DP_OP_425J2_127_3477_n1854, DP_OP_425J2_127_3477_n1853,
         DP_OP_425J2_127_3477_n1852, DP_OP_425J2_127_3477_n1851,
         DP_OP_425J2_127_3477_n1850, DP_OP_425J2_127_3477_n1849,
         DP_OP_425J2_127_3477_n1848, DP_OP_425J2_127_3477_n1847,
         DP_OP_425J2_127_3477_n1846, DP_OP_425J2_127_3477_n1845,
         DP_OP_425J2_127_3477_n1844, DP_OP_425J2_127_3477_n1843,
         DP_OP_425J2_127_3477_n1842, DP_OP_425J2_127_3477_n1841,
         DP_OP_425J2_127_3477_n1840, DP_OP_425J2_127_3477_n1839,
         DP_OP_425J2_127_3477_n1838, DP_OP_425J2_127_3477_n1837,
         DP_OP_425J2_127_3477_n1836, DP_OP_425J2_127_3477_n1835,
         DP_OP_425J2_127_3477_n1834, DP_OP_425J2_127_3477_n1833,
         DP_OP_425J2_127_3477_n1832, DP_OP_425J2_127_3477_n1831,
         DP_OP_425J2_127_3477_n1830, DP_OP_425J2_127_3477_n1829,
         DP_OP_425J2_127_3477_n1828, DP_OP_425J2_127_3477_n1827,
         DP_OP_425J2_127_3477_n1826, DP_OP_425J2_127_3477_n1825,
         DP_OP_425J2_127_3477_n1824, DP_OP_425J2_127_3477_n1823,
         DP_OP_425J2_127_3477_n1822, DP_OP_425J2_127_3477_n1821,
         DP_OP_425J2_127_3477_n1820, DP_OP_425J2_127_3477_n1819,
         DP_OP_425J2_127_3477_n1818, DP_OP_425J2_127_3477_n1817,
         DP_OP_425J2_127_3477_n1816, DP_OP_425J2_127_3477_n1815,
         DP_OP_425J2_127_3477_n1814, DP_OP_425J2_127_3477_n1813,
         DP_OP_425J2_127_3477_n1812, DP_OP_425J2_127_3477_n1811,
         DP_OP_425J2_127_3477_n1810, DP_OP_425J2_127_3477_n1809,
         DP_OP_425J2_127_3477_n1808, DP_OP_425J2_127_3477_n1807,
         DP_OP_425J2_127_3477_n1806, DP_OP_425J2_127_3477_n1805,
         DP_OP_425J2_127_3477_n1804, DP_OP_425J2_127_3477_n1803,
         DP_OP_425J2_127_3477_n1802, DP_OP_425J2_127_3477_n1801,
         DP_OP_425J2_127_3477_n1800, DP_OP_425J2_127_3477_n1799,
         DP_OP_425J2_127_3477_n1798, DP_OP_425J2_127_3477_n1797,
         DP_OP_425J2_127_3477_n1796, DP_OP_425J2_127_3477_n1795,
         DP_OP_425J2_127_3477_n1794, DP_OP_425J2_127_3477_n1793,
         DP_OP_425J2_127_3477_n1792, DP_OP_425J2_127_3477_n1791,
         DP_OP_425J2_127_3477_n1790, DP_OP_425J2_127_3477_n1789,
         DP_OP_425J2_127_3477_n1788, DP_OP_425J2_127_3477_n1787,
         DP_OP_425J2_127_3477_n1786, DP_OP_425J2_127_3477_n1785,
         DP_OP_425J2_127_3477_n1784, DP_OP_425J2_127_3477_n1783,
         DP_OP_425J2_127_3477_n1782, DP_OP_425J2_127_3477_n1781,
         DP_OP_425J2_127_3477_n1780, DP_OP_425J2_127_3477_n1779,
         DP_OP_425J2_127_3477_n1778, DP_OP_425J2_127_3477_n1777,
         DP_OP_425J2_127_3477_n1776, DP_OP_425J2_127_3477_n1775,
         DP_OP_425J2_127_3477_n1774, DP_OP_425J2_127_3477_n1773,
         DP_OP_425J2_127_3477_n1772, DP_OP_425J2_127_3477_n1771,
         DP_OP_425J2_127_3477_n1770, DP_OP_425J2_127_3477_n1769,
         DP_OP_425J2_127_3477_n1768, DP_OP_425J2_127_3477_n1767,
         DP_OP_425J2_127_3477_n1766, DP_OP_425J2_127_3477_n1765,
         DP_OP_425J2_127_3477_n1764, DP_OP_425J2_127_3477_n1763,
         DP_OP_425J2_127_3477_n1762, DP_OP_425J2_127_3477_n1761,
         DP_OP_425J2_127_3477_n1760, DP_OP_425J2_127_3477_n1759,
         DP_OP_425J2_127_3477_n1758, DP_OP_425J2_127_3477_n1757,
         DP_OP_425J2_127_3477_n1756, DP_OP_425J2_127_3477_n1755,
         DP_OP_425J2_127_3477_n1754, DP_OP_425J2_127_3477_n1753,
         DP_OP_425J2_127_3477_n1752, DP_OP_425J2_127_3477_n1751,
         DP_OP_425J2_127_3477_n1750, DP_OP_425J2_127_3477_n1749,
         DP_OP_425J2_127_3477_n1748, DP_OP_425J2_127_3477_n1747,
         DP_OP_425J2_127_3477_n1746, DP_OP_425J2_127_3477_n1745,
         DP_OP_425J2_127_3477_n1744, DP_OP_425J2_127_3477_n1743,
         DP_OP_425J2_127_3477_n1742, DP_OP_425J2_127_3477_n1741,
         DP_OP_425J2_127_3477_n1740, DP_OP_425J2_127_3477_n1739,
         DP_OP_425J2_127_3477_n1738, DP_OP_425J2_127_3477_n1737,
         DP_OP_425J2_127_3477_n1736, DP_OP_425J2_127_3477_n1735,
         DP_OP_425J2_127_3477_n1734, DP_OP_425J2_127_3477_n1733,
         DP_OP_425J2_127_3477_n1732, DP_OP_425J2_127_3477_n1731,
         DP_OP_425J2_127_3477_n1730, DP_OP_425J2_127_3477_n1729,
         DP_OP_425J2_127_3477_n1728, DP_OP_425J2_127_3477_n1727,
         DP_OP_425J2_127_3477_n1726, DP_OP_425J2_127_3477_n1725,
         DP_OP_425J2_127_3477_n1724, DP_OP_425J2_127_3477_n1723,
         DP_OP_425J2_127_3477_n1722, DP_OP_425J2_127_3477_n1721,
         DP_OP_425J2_127_3477_n1720, DP_OP_425J2_127_3477_n1719,
         DP_OP_425J2_127_3477_n1718, DP_OP_425J2_127_3477_n1717,
         DP_OP_425J2_127_3477_n1716, DP_OP_425J2_127_3477_n1715,
         DP_OP_425J2_127_3477_n1714, DP_OP_425J2_127_3477_n1713,
         DP_OP_425J2_127_3477_n1712, DP_OP_425J2_127_3477_n1711,
         DP_OP_425J2_127_3477_n1710, DP_OP_425J2_127_3477_n1709,
         DP_OP_425J2_127_3477_n1708, DP_OP_425J2_127_3477_n1707,
         DP_OP_425J2_127_3477_n1706, DP_OP_425J2_127_3477_n1705,
         DP_OP_425J2_127_3477_n1704, DP_OP_425J2_127_3477_n1703,
         DP_OP_425J2_127_3477_n1702, DP_OP_425J2_127_3477_n1701,
         DP_OP_425J2_127_3477_n1700, DP_OP_425J2_127_3477_n1699,
         DP_OP_425J2_127_3477_n1698, DP_OP_425J2_127_3477_n1697,
         DP_OP_425J2_127_3477_n1696, DP_OP_425J2_127_3477_n1695,
         DP_OP_425J2_127_3477_n1694, DP_OP_425J2_127_3477_n1693,
         DP_OP_425J2_127_3477_n1692, DP_OP_425J2_127_3477_n1691,
         DP_OP_425J2_127_3477_n1690, DP_OP_425J2_127_3477_n1689,
         DP_OP_425J2_127_3477_n1688, DP_OP_425J2_127_3477_n1687,
         DP_OP_425J2_127_3477_n1686, DP_OP_425J2_127_3477_n1685,
         DP_OP_425J2_127_3477_n1684, DP_OP_425J2_127_3477_n1683,
         DP_OP_425J2_127_3477_n1682, DP_OP_425J2_127_3477_n1681,
         DP_OP_425J2_127_3477_n1680, DP_OP_425J2_127_3477_n1679,
         DP_OP_425J2_127_3477_n1678, DP_OP_425J2_127_3477_n1677,
         DP_OP_425J2_127_3477_n1676, DP_OP_425J2_127_3477_n1675,
         DP_OP_425J2_127_3477_n1674, DP_OP_425J2_127_3477_n1673,
         DP_OP_425J2_127_3477_n1672, DP_OP_425J2_127_3477_n1671,
         DP_OP_425J2_127_3477_n1670, DP_OP_425J2_127_3477_n1669,
         DP_OP_425J2_127_3477_n1668, DP_OP_425J2_127_3477_n1667,
         DP_OP_425J2_127_3477_n1666, DP_OP_425J2_127_3477_n1665,
         DP_OP_425J2_127_3477_n1664, DP_OP_425J2_127_3477_n1663,
         DP_OP_425J2_127_3477_n1662, DP_OP_425J2_127_3477_n1661,
         DP_OP_425J2_127_3477_n1660, DP_OP_425J2_127_3477_n1659,
         DP_OP_425J2_127_3477_n1658, DP_OP_425J2_127_3477_n1657,
         DP_OP_425J2_127_3477_n1656, DP_OP_425J2_127_3477_n1655,
         DP_OP_425J2_127_3477_n1654, DP_OP_425J2_127_3477_n1653,
         DP_OP_425J2_127_3477_n1652, DP_OP_425J2_127_3477_n1651,
         DP_OP_425J2_127_3477_n1650, DP_OP_425J2_127_3477_n1649,
         DP_OP_425J2_127_3477_n1648, DP_OP_425J2_127_3477_n1647,
         DP_OP_425J2_127_3477_n1646, DP_OP_425J2_127_3477_n1645,
         DP_OP_425J2_127_3477_n1644, DP_OP_425J2_127_3477_n1643,
         DP_OP_425J2_127_3477_n1642, DP_OP_425J2_127_3477_n1641,
         DP_OP_425J2_127_3477_n1640, DP_OP_425J2_127_3477_n1639,
         DP_OP_425J2_127_3477_n1638, DP_OP_425J2_127_3477_n1637,
         DP_OP_425J2_127_3477_n1636, DP_OP_425J2_127_3477_n1635,
         DP_OP_425J2_127_3477_n1634, DP_OP_425J2_127_3477_n1633,
         DP_OP_425J2_127_3477_n1632, DP_OP_425J2_127_3477_n1631,
         DP_OP_425J2_127_3477_n1630, DP_OP_425J2_127_3477_n1629,
         DP_OP_425J2_127_3477_n1628, DP_OP_425J2_127_3477_n1627,
         DP_OP_425J2_127_3477_n1626, DP_OP_425J2_127_3477_n1625,
         DP_OP_425J2_127_3477_n1624, DP_OP_425J2_127_3477_n1623,
         DP_OP_425J2_127_3477_n1622, DP_OP_425J2_127_3477_n1621,
         DP_OP_425J2_127_3477_n1620, DP_OP_425J2_127_3477_n1619,
         DP_OP_425J2_127_3477_n1618, DP_OP_425J2_127_3477_n1617,
         DP_OP_425J2_127_3477_n1616, DP_OP_425J2_127_3477_n1615,
         DP_OP_425J2_127_3477_n1614, DP_OP_425J2_127_3477_n1613,
         DP_OP_425J2_127_3477_n1612, DP_OP_425J2_127_3477_n1611,
         DP_OP_425J2_127_3477_n1610, DP_OP_425J2_127_3477_n1609,
         DP_OP_425J2_127_3477_n1608, DP_OP_425J2_127_3477_n1607,
         DP_OP_425J2_127_3477_n1606, DP_OP_425J2_127_3477_n1605,
         DP_OP_425J2_127_3477_n1604, DP_OP_425J2_127_3477_n1603,
         DP_OP_425J2_127_3477_n1602, DP_OP_425J2_127_3477_n1601,
         DP_OP_425J2_127_3477_n1600, DP_OP_425J2_127_3477_n1599,
         DP_OP_425J2_127_3477_n1598, DP_OP_425J2_127_3477_n1597,
         DP_OP_425J2_127_3477_n1596, DP_OP_425J2_127_3477_n1595,
         DP_OP_425J2_127_3477_n1594, DP_OP_425J2_127_3477_n1593,
         DP_OP_425J2_127_3477_n1592, DP_OP_425J2_127_3477_n1591,
         DP_OP_425J2_127_3477_n1590, DP_OP_425J2_127_3477_n1589,
         DP_OP_425J2_127_3477_n1588, DP_OP_425J2_127_3477_n1587,
         DP_OP_425J2_127_3477_n1586, DP_OP_425J2_127_3477_n1585,
         DP_OP_425J2_127_3477_n1584, DP_OP_425J2_127_3477_n1583,
         DP_OP_425J2_127_3477_n1582, DP_OP_425J2_127_3477_n1581,
         DP_OP_425J2_127_3477_n1580, DP_OP_425J2_127_3477_n1579,
         DP_OP_425J2_127_3477_n1578, DP_OP_425J2_127_3477_n1577,
         DP_OP_425J2_127_3477_n1576, DP_OP_425J2_127_3477_n1575,
         DP_OP_425J2_127_3477_n1574, DP_OP_425J2_127_3477_n1573,
         DP_OP_425J2_127_3477_n1572, DP_OP_425J2_127_3477_n1571,
         DP_OP_425J2_127_3477_n1570, DP_OP_425J2_127_3477_n1569,
         DP_OP_425J2_127_3477_n1568, DP_OP_425J2_127_3477_n1567,
         DP_OP_425J2_127_3477_n1566, DP_OP_425J2_127_3477_n1565,
         DP_OP_425J2_127_3477_n1564, DP_OP_425J2_127_3477_n1563,
         DP_OP_425J2_127_3477_n1562, DP_OP_425J2_127_3477_n1561,
         DP_OP_425J2_127_3477_n1560, DP_OP_425J2_127_3477_n1559,
         DP_OP_425J2_127_3477_n1558, DP_OP_425J2_127_3477_n1557,
         DP_OP_425J2_127_3477_n1556, DP_OP_425J2_127_3477_n1555,
         DP_OP_425J2_127_3477_n1554, DP_OP_425J2_127_3477_n1553,
         DP_OP_425J2_127_3477_n1552, DP_OP_425J2_127_3477_n1551,
         DP_OP_425J2_127_3477_n1550, DP_OP_425J2_127_3477_n1549,
         DP_OP_425J2_127_3477_n1548, DP_OP_425J2_127_3477_n1547,
         DP_OP_425J2_127_3477_n1546, DP_OP_425J2_127_3477_n1545,
         DP_OP_425J2_127_3477_n1544, DP_OP_425J2_127_3477_n1543,
         DP_OP_425J2_127_3477_n1542, DP_OP_425J2_127_3477_n1541,
         DP_OP_425J2_127_3477_n1540, DP_OP_425J2_127_3477_n1539,
         DP_OP_425J2_127_3477_n1538, DP_OP_425J2_127_3477_n1537,
         DP_OP_425J2_127_3477_n1536, DP_OP_425J2_127_3477_n1535,
         DP_OP_425J2_127_3477_n1534, DP_OP_425J2_127_3477_n1533,
         DP_OP_425J2_127_3477_n1532, DP_OP_425J2_127_3477_n1531,
         DP_OP_425J2_127_3477_n1530, DP_OP_425J2_127_3477_n1529,
         DP_OP_425J2_127_3477_n1528, DP_OP_425J2_127_3477_n1527,
         DP_OP_425J2_127_3477_n1526, DP_OP_425J2_127_3477_n1525,
         DP_OP_425J2_127_3477_n1524, DP_OP_425J2_127_3477_n1523,
         DP_OP_425J2_127_3477_n1522, DP_OP_425J2_127_3477_n1521,
         DP_OP_425J2_127_3477_n1520, DP_OP_425J2_127_3477_n1519,
         DP_OP_425J2_127_3477_n1518, DP_OP_425J2_127_3477_n1517,
         DP_OP_425J2_127_3477_n1516, DP_OP_425J2_127_3477_n1515,
         DP_OP_425J2_127_3477_n1514, DP_OP_425J2_127_3477_n1513,
         DP_OP_425J2_127_3477_n1512, DP_OP_425J2_127_3477_n1511,
         DP_OP_425J2_127_3477_n1510, DP_OP_425J2_127_3477_n1509,
         DP_OP_425J2_127_3477_n1508, DP_OP_425J2_127_3477_n1507,
         DP_OP_425J2_127_3477_n1506, DP_OP_425J2_127_3477_n1505,
         DP_OP_425J2_127_3477_n1504, DP_OP_425J2_127_3477_n1503,
         DP_OP_425J2_127_3477_n1502, DP_OP_425J2_127_3477_n1501,
         DP_OP_425J2_127_3477_n1500, DP_OP_425J2_127_3477_n1499,
         DP_OP_425J2_127_3477_n1498, DP_OP_425J2_127_3477_n1497,
         DP_OP_425J2_127_3477_n1496, DP_OP_425J2_127_3477_n1495,
         DP_OP_425J2_127_3477_n1494, DP_OP_425J2_127_3477_n1493,
         DP_OP_425J2_127_3477_n1492, DP_OP_425J2_127_3477_n1491,
         DP_OP_425J2_127_3477_n1490, DP_OP_425J2_127_3477_n1489,
         DP_OP_425J2_127_3477_n1488, DP_OP_425J2_127_3477_n1487,
         DP_OP_425J2_127_3477_n1486, DP_OP_425J2_127_3477_n1485,
         DP_OP_425J2_127_3477_n1484, DP_OP_425J2_127_3477_n1483,
         DP_OP_425J2_127_3477_n1482, DP_OP_425J2_127_3477_n1481,
         DP_OP_425J2_127_3477_n1480, DP_OP_425J2_127_3477_n1479,
         DP_OP_425J2_127_3477_n1478, DP_OP_425J2_127_3477_n1477,
         DP_OP_425J2_127_3477_n1476, DP_OP_425J2_127_3477_n1475,
         DP_OP_425J2_127_3477_n1474, DP_OP_425J2_127_3477_n1473,
         DP_OP_425J2_127_3477_n1472, DP_OP_425J2_127_3477_n1471,
         DP_OP_425J2_127_3477_n1470, DP_OP_425J2_127_3477_n1469,
         DP_OP_425J2_127_3477_n1468, DP_OP_425J2_127_3477_n1467,
         DP_OP_425J2_127_3477_n1466, DP_OP_425J2_127_3477_n1465,
         DP_OP_425J2_127_3477_n1464, DP_OP_425J2_127_3477_n1463,
         DP_OP_425J2_127_3477_n1462, DP_OP_425J2_127_3477_n1461,
         DP_OP_425J2_127_3477_n1460, DP_OP_425J2_127_3477_n1459,
         DP_OP_425J2_127_3477_n1458, DP_OP_425J2_127_3477_n1457,
         DP_OP_425J2_127_3477_n1456, DP_OP_425J2_127_3477_n1455,
         DP_OP_425J2_127_3477_n1454, DP_OP_425J2_127_3477_n1453,
         DP_OP_425J2_127_3477_n1452, DP_OP_425J2_127_3477_n1451,
         DP_OP_425J2_127_3477_n1450, DP_OP_425J2_127_3477_n1449,
         DP_OP_425J2_127_3477_n1448, DP_OP_425J2_127_3477_n1447,
         DP_OP_425J2_127_3477_n1446, DP_OP_425J2_127_3477_n1445,
         DP_OP_425J2_127_3477_n1444, DP_OP_425J2_127_3477_n1443,
         DP_OP_425J2_127_3477_n1442, DP_OP_425J2_127_3477_n1441,
         DP_OP_425J2_127_3477_n1440, DP_OP_425J2_127_3477_n1439,
         DP_OP_425J2_127_3477_n1438, DP_OP_425J2_127_3477_n1437,
         DP_OP_425J2_127_3477_n1436, DP_OP_425J2_127_3477_n1435,
         DP_OP_425J2_127_3477_n1434, DP_OP_425J2_127_3477_n1433,
         DP_OP_425J2_127_3477_n1432, DP_OP_425J2_127_3477_n1431,
         DP_OP_425J2_127_3477_n1430, DP_OP_425J2_127_3477_n1429,
         DP_OP_425J2_127_3477_n1428, DP_OP_425J2_127_3477_n1427,
         DP_OP_425J2_127_3477_n1426, DP_OP_425J2_127_3477_n1425,
         DP_OP_425J2_127_3477_n1424, DP_OP_425J2_127_3477_n1423,
         DP_OP_425J2_127_3477_n1422, DP_OP_425J2_127_3477_n1421,
         DP_OP_425J2_127_3477_n1420, DP_OP_425J2_127_3477_n1419,
         DP_OP_425J2_127_3477_n1418, DP_OP_425J2_127_3477_n1417,
         DP_OP_425J2_127_3477_n1416, DP_OP_425J2_127_3477_n1415,
         DP_OP_425J2_127_3477_n1414, DP_OP_425J2_127_3477_n1413,
         DP_OP_425J2_127_3477_n1412, DP_OP_425J2_127_3477_n1411,
         DP_OP_425J2_127_3477_n1410, DP_OP_425J2_127_3477_n1409,
         DP_OP_425J2_127_3477_n1408, DP_OP_425J2_127_3477_n1407,
         DP_OP_425J2_127_3477_n1406, DP_OP_425J2_127_3477_n1405,
         DP_OP_425J2_127_3477_n1404, DP_OP_425J2_127_3477_n1403,
         DP_OP_425J2_127_3477_n1402, DP_OP_425J2_127_3477_n1401,
         DP_OP_425J2_127_3477_n1400, DP_OP_425J2_127_3477_n1399,
         DP_OP_425J2_127_3477_n1398, DP_OP_425J2_127_3477_n1397,
         DP_OP_425J2_127_3477_n1396, DP_OP_425J2_127_3477_n1395,
         DP_OP_425J2_127_3477_n1394, DP_OP_425J2_127_3477_n1393,
         DP_OP_425J2_127_3477_n1392, DP_OP_425J2_127_3477_n1391,
         DP_OP_425J2_127_3477_n1390, DP_OP_425J2_127_3477_n1389,
         DP_OP_425J2_127_3477_n1388, DP_OP_425J2_127_3477_n1387,
         DP_OP_425J2_127_3477_n1386, DP_OP_425J2_127_3477_n1385,
         DP_OP_425J2_127_3477_n1384, DP_OP_425J2_127_3477_n1383,
         DP_OP_425J2_127_3477_n1382, DP_OP_425J2_127_3477_n1381,
         DP_OP_425J2_127_3477_n1380, DP_OP_425J2_127_3477_n1379,
         DP_OP_425J2_127_3477_n1378, DP_OP_425J2_127_3477_n1377,
         DP_OP_425J2_127_3477_n1376, DP_OP_425J2_127_3477_n1375,
         DP_OP_425J2_127_3477_n1374, DP_OP_425J2_127_3477_n1373,
         DP_OP_425J2_127_3477_n1372, DP_OP_425J2_127_3477_n1371,
         DP_OP_425J2_127_3477_n1370, DP_OP_425J2_127_3477_n1369,
         DP_OP_425J2_127_3477_n1368, DP_OP_425J2_127_3477_n1367,
         DP_OP_425J2_127_3477_n1366, DP_OP_425J2_127_3477_n1365,
         DP_OP_425J2_127_3477_n1364, DP_OP_425J2_127_3477_n1363,
         DP_OP_425J2_127_3477_n1362, DP_OP_425J2_127_3477_n1361,
         DP_OP_425J2_127_3477_n1360, DP_OP_425J2_127_3477_n1359,
         DP_OP_425J2_127_3477_n1358, DP_OP_425J2_127_3477_n1357,
         DP_OP_425J2_127_3477_n1356, DP_OP_425J2_127_3477_n1355,
         DP_OP_425J2_127_3477_n1354, DP_OP_425J2_127_3477_n1353,
         DP_OP_425J2_127_3477_n1352, DP_OP_425J2_127_3477_n1351,
         DP_OP_425J2_127_3477_n1350, DP_OP_425J2_127_3477_n1349,
         DP_OP_425J2_127_3477_n1348, DP_OP_425J2_127_3477_n1347,
         DP_OP_425J2_127_3477_n1346, DP_OP_425J2_127_3477_n1345,
         DP_OP_425J2_127_3477_n1344, DP_OP_425J2_127_3477_n1343,
         DP_OP_425J2_127_3477_n1342, DP_OP_425J2_127_3477_n1341,
         DP_OP_425J2_127_3477_n1340, DP_OP_425J2_127_3477_n1339,
         DP_OP_425J2_127_3477_n1338, DP_OP_425J2_127_3477_n1337,
         DP_OP_425J2_127_3477_n1336, DP_OP_425J2_127_3477_n1335,
         DP_OP_425J2_127_3477_n1334, DP_OP_425J2_127_3477_n1333,
         DP_OP_425J2_127_3477_n1332, DP_OP_425J2_127_3477_n1331,
         DP_OP_425J2_127_3477_n1330, DP_OP_425J2_127_3477_n1329,
         DP_OP_425J2_127_3477_n1328, DP_OP_425J2_127_3477_n1327,
         DP_OP_425J2_127_3477_n1326, DP_OP_425J2_127_3477_n1325,
         DP_OP_425J2_127_3477_n1324, DP_OP_425J2_127_3477_n1323,
         DP_OP_425J2_127_3477_n1322, DP_OP_425J2_127_3477_n1321,
         DP_OP_425J2_127_3477_n1320, DP_OP_425J2_127_3477_n1319,
         DP_OP_425J2_127_3477_n1318, DP_OP_425J2_127_3477_n1317,
         DP_OP_425J2_127_3477_n1316, DP_OP_425J2_127_3477_n1315,
         DP_OP_425J2_127_3477_n1314, DP_OP_425J2_127_3477_n1313,
         DP_OP_425J2_127_3477_n1312, DP_OP_425J2_127_3477_n1311,
         DP_OP_425J2_127_3477_n1310, DP_OP_425J2_127_3477_n1309,
         DP_OP_425J2_127_3477_n1308, DP_OP_425J2_127_3477_n1307,
         DP_OP_425J2_127_3477_n1306, DP_OP_425J2_127_3477_n1305,
         DP_OP_425J2_127_3477_n1304, DP_OP_425J2_127_3477_n1303,
         DP_OP_425J2_127_3477_n1302, DP_OP_425J2_127_3477_n1301,
         DP_OP_425J2_127_3477_n1300, DP_OP_425J2_127_3477_n1299,
         DP_OP_425J2_127_3477_n1298, DP_OP_425J2_127_3477_n1297,
         DP_OP_425J2_127_3477_n1296, DP_OP_425J2_127_3477_n1295,
         DP_OP_425J2_127_3477_n1294, DP_OP_425J2_127_3477_n1293,
         DP_OP_425J2_127_3477_n1292, DP_OP_425J2_127_3477_n1291,
         DP_OP_425J2_127_3477_n1290, DP_OP_425J2_127_3477_n1289,
         DP_OP_425J2_127_3477_n1288, DP_OP_425J2_127_3477_n1287,
         DP_OP_425J2_127_3477_n1286, DP_OP_425J2_127_3477_n1285,
         DP_OP_425J2_127_3477_n1284, DP_OP_425J2_127_3477_n1283,
         DP_OP_425J2_127_3477_n1282, DP_OP_425J2_127_3477_n1281,
         DP_OP_425J2_127_3477_n1280, DP_OP_425J2_127_3477_n1279,
         DP_OP_425J2_127_3477_n1278, DP_OP_425J2_127_3477_n1277,
         DP_OP_425J2_127_3477_n1276, DP_OP_425J2_127_3477_n1275,
         DP_OP_425J2_127_3477_n1274, DP_OP_425J2_127_3477_n1273,
         DP_OP_425J2_127_3477_n1272, DP_OP_425J2_127_3477_n1271,
         DP_OP_425J2_127_3477_n1270, DP_OP_425J2_127_3477_n1269,
         DP_OP_425J2_127_3477_n1268, DP_OP_425J2_127_3477_n1267,
         DP_OP_425J2_127_3477_n1266, DP_OP_425J2_127_3477_n1265,
         DP_OP_425J2_127_3477_n1264, DP_OP_425J2_127_3477_n1263,
         DP_OP_425J2_127_3477_n1262, DP_OP_425J2_127_3477_n1261,
         DP_OP_425J2_127_3477_n1260, DP_OP_425J2_127_3477_n1259,
         DP_OP_425J2_127_3477_n1258, DP_OP_425J2_127_3477_n1257,
         DP_OP_425J2_127_3477_n1256, DP_OP_425J2_127_3477_n1255,
         DP_OP_425J2_127_3477_n1254, DP_OP_425J2_127_3477_n1253,
         DP_OP_425J2_127_3477_n1252, DP_OP_425J2_127_3477_n1251,
         DP_OP_425J2_127_3477_n1250, DP_OP_425J2_127_3477_n1249,
         DP_OP_425J2_127_3477_n1248, DP_OP_425J2_127_3477_n1247,
         DP_OP_425J2_127_3477_n1246, DP_OP_425J2_127_3477_n1245,
         DP_OP_425J2_127_3477_n1244, DP_OP_425J2_127_3477_n1243,
         DP_OP_425J2_127_3477_n1242, DP_OP_425J2_127_3477_n1241,
         DP_OP_425J2_127_3477_n1240, DP_OP_425J2_127_3477_n1239,
         DP_OP_425J2_127_3477_n1238, DP_OP_425J2_127_3477_n1237,
         DP_OP_425J2_127_3477_n1236, DP_OP_425J2_127_3477_n1235,
         DP_OP_425J2_127_3477_n1234, DP_OP_425J2_127_3477_n1233,
         DP_OP_425J2_127_3477_n1232, DP_OP_425J2_127_3477_n1231,
         DP_OP_425J2_127_3477_n1230, DP_OP_425J2_127_3477_n1229,
         DP_OP_425J2_127_3477_n1228, DP_OP_425J2_127_3477_n1227,
         DP_OP_425J2_127_3477_n1226, DP_OP_425J2_127_3477_n1225,
         DP_OP_425J2_127_3477_n1224, DP_OP_425J2_127_3477_n1223,
         DP_OP_425J2_127_3477_n1222, DP_OP_425J2_127_3477_n1221,
         DP_OP_425J2_127_3477_n1220, DP_OP_425J2_127_3477_n1219,
         DP_OP_425J2_127_3477_n1218, DP_OP_425J2_127_3477_n1217,
         DP_OP_425J2_127_3477_n1216, DP_OP_425J2_127_3477_n1215,
         DP_OP_425J2_127_3477_n1214, DP_OP_425J2_127_3477_n1213,
         DP_OP_425J2_127_3477_n1212, DP_OP_425J2_127_3477_n1211,
         DP_OP_425J2_127_3477_n1210, DP_OP_425J2_127_3477_n1209,
         DP_OP_425J2_127_3477_n1208, DP_OP_425J2_127_3477_n1207,
         DP_OP_425J2_127_3477_n1206, DP_OP_425J2_127_3477_n1205,
         DP_OP_425J2_127_3477_n1204, DP_OP_425J2_127_3477_n1203,
         DP_OP_425J2_127_3477_n1202, DP_OP_425J2_127_3477_n1201,
         DP_OP_425J2_127_3477_n1200, DP_OP_425J2_127_3477_n1199,
         DP_OP_425J2_127_3477_n1198, DP_OP_425J2_127_3477_n1197,
         DP_OP_425J2_127_3477_n1196, DP_OP_425J2_127_3477_n1195,
         DP_OP_425J2_127_3477_n1194, DP_OP_425J2_127_3477_n1193,
         DP_OP_425J2_127_3477_n1192, DP_OP_425J2_127_3477_n1191,
         DP_OP_425J2_127_3477_n1190, DP_OP_425J2_127_3477_n1189,
         DP_OP_425J2_127_3477_n1188, DP_OP_425J2_127_3477_n1187,
         DP_OP_425J2_127_3477_n1186, DP_OP_425J2_127_3477_n1185,
         DP_OP_425J2_127_3477_n1184, DP_OP_425J2_127_3477_n1183,
         DP_OP_425J2_127_3477_n1182, DP_OP_425J2_127_3477_n1181,
         DP_OP_425J2_127_3477_n1180, DP_OP_425J2_127_3477_n1179,
         DP_OP_425J2_127_3477_n1178, DP_OP_425J2_127_3477_n1177,
         DP_OP_425J2_127_3477_n1176, DP_OP_425J2_127_3477_n1175,
         DP_OP_425J2_127_3477_n1174, DP_OP_425J2_127_3477_n1173,
         DP_OP_425J2_127_3477_n1172, DP_OP_425J2_127_3477_n1171,
         DP_OP_425J2_127_3477_n1170, DP_OP_425J2_127_3477_n1169,
         DP_OP_425J2_127_3477_n1168, DP_OP_425J2_127_3477_n1167,
         DP_OP_425J2_127_3477_n1166, DP_OP_425J2_127_3477_n1165,
         DP_OP_425J2_127_3477_n1164, DP_OP_425J2_127_3477_n1163,
         DP_OP_425J2_127_3477_n1162, DP_OP_425J2_127_3477_n1161,
         DP_OP_425J2_127_3477_n1160, DP_OP_425J2_127_3477_n1159,
         DP_OP_425J2_127_3477_n1158, DP_OP_425J2_127_3477_n1157,
         DP_OP_425J2_127_3477_n1156, DP_OP_425J2_127_3477_n1155,
         DP_OP_425J2_127_3477_n1154, DP_OP_425J2_127_3477_n1153,
         DP_OP_425J2_127_3477_n1152, DP_OP_425J2_127_3477_n1151,
         DP_OP_425J2_127_3477_n1150, DP_OP_425J2_127_3477_n1149,
         DP_OP_425J2_127_3477_n1148, DP_OP_425J2_127_3477_n1147,
         DP_OP_425J2_127_3477_n1146, DP_OP_425J2_127_3477_n1145,
         DP_OP_425J2_127_3477_n1144, DP_OP_425J2_127_3477_n1143,
         DP_OP_425J2_127_3477_n1142, DP_OP_425J2_127_3477_n1141,
         DP_OP_425J2_127_3477_n1140, DP_OP_425J2_127_3477_n1139,
         DP_OP_425J2_127_3477_n1138, DP_OP_425J2_127_3477_n1137,
         DP_OP_425J2_127_3477_n1136, DP_OP_425J2_127_3477_n1135,
         DP_OP_425J2_127_3477_n1134, DP_OP_425J2_127_3477_n1133,
         DP_OP_425J2_127_3477_n1132, DP_OP_425J2_127_3477_n1131,
         DP_OP_425J2_127_3477_n1130, DP_OP_425J2_127_3477_n1129,
         DP_OP_425J2_127_3477_n1128, DP_OP_425J2_127_3477_n1127,
         DP_OP_425J2_127_3477_n1126, DP_OP_425J2_127_3477_n1125,
         DP_OP_425J2_127_3477_n1124, DP_OP_425J2_127_3477_n1123,
         DP_OP_425J2_127_3477_n1122, DP_OP_425J2_127_3477_n1121,
         DP_OP_425J2_127_3477_n1120, DP_OP_425J2_127_3477_n1119,
         DP_OP_425J2_127_3477_n1118, DP_OP_425J2_127_3477_n1117,
         DP_OP_425J2_127_3477_n1116, DP_OP_425J2_127_3477_n1115,
         DP_OP_425J2_127_3477_n1114, DP_OP_425J2_127_3477_n1113,
         DP_OP_425J2_127_3477_n1112, DP_OP_425J2_127_3477_n1111,
         DP_OP_425J2_127_3477_n1110, DP_OP_425J2_127_3477_n1109,
         DP_OP_425J2_127_3477_n1108, DP_OP_425J2_127_3477_n1107,
         DP_OP_425J2_127_3477_n1106, DP_OP_425J2_127_3477_n1105,
         DP_OP_425J2_127_3477_n1104, DP_OP_425J2_127_3477_n1103,
         DP_OP_425J2_127_3477_n1102, DP_OP_425J2_127_3477_n1101,
         DP_OP_425J2_127_3477_n1100, DP_OP_425J2_127_3477_n1099,
         DP_OP_425J2_127_3477_n1098, DP_OP_425J2_127_3477_n1097,
         DP_OP_425J2_127_3477_n1096, DP_OP_425J2_127_3477_n1095,
         DP_OP_425J2_127_3477_n1094, DP_OP_425J2_127_3477_n1093,
         DP_OP_425J2_127_3477_n1092, DP_OP_425J2_127_3477_n1091,
         DP_OP_425J2_127_3477_n1090, DP_OP_425J2_127_3477_n1089,
         DP_OP_425J2_127_3477_n1088, DP_OP_425J2_127_3477_n1087,
         DP_OP_425J2_127_3477_n1086, DP_OP_425J2_127_3477_n1085,
         DP_OP_425J2_127_3477_n1084, DP_OP_425J2_127_3477_n1083,
         DP_OP_425J2_127_3477_n1082, DP_OP_425J2_127_3477_n1081,
         DP_OP_425J2_127_3477_n1080, DP_OP_425J2_127_3477_n1079,
         DP_OP_425J2_127_3477_n1078, DP_OP_425J2_127_3477_n1077,
         DP_OP_425J2_127_3477_n1076, DP_OP_425J2_127_3477_n1075,
         DP_OP_425J2_127_3477_n1074, DP_OP_425J2_127_3477_n1073,
         DP_OP_425J2_127_3477_n1072, DP_OP_425J2_127_3477_n1071,
         DP_OP_425J2_127_3477_n1070, DP_OP_425J2_127_3477_n1069,
         DP_OP_425J2_127_3477_n1068, DP_OP_425J2_127_3477_n1067,
         DP_OP_425J2_127_3477_n1066, DP_OP_425J2_127_3477_n1065,
         DP_OP_425J2_127_3477_n1064, DP_OP_425J2_127_3477_n1063,
         DP_OP_425J2_127_3477_n1062, DP_OP_425J2_127_3477_n1061,
         DP_OP_425J2_127_3477_n1060, DP_OP_425J2_127_3477_n1059,
         DP_OP_425J2_127_3477_n1058, DP_OP_425J2_127_3477_n1057,
         DP_OP_425J2_127_3477_n1056, DP_OP_425J2_127_3477_n1055,
         DP_OP_425J2_127_3477_n1054, DP_OP_425J2_127_3477_n1053,
         DP_OP_425J2_127_3477_n1052, DP_OP_425J2_127_3477_n1051,
         DP_OP_425J2_127_3477_n1050, DP_OP_425J2_127_3477_n1049,
         DP_OP_425J2_127_3477_n1048, DP_OP_425J2_127_3477_n1047,
         DP_OP_425J2_127_3477_n1046, DP_OP_425J2_127_3477_n1045,
         DP_OP_425J2_127_3477_n1044, DP_OP_425J2_127_3477_n1043,
         DP_OP_425J2_127_3477_n1042, DP_OP_425J2_127_3477_n1041,
         DP_OP_425J2_127_3477_n1040, DP_OP_425J2_127_3477_n1039,
         DP_OP_425J2_127_3477_n1038, DP_OP_425J2_127_3477_n1037,
         DP_OP_425J2_127_3477_n1036, DP_OP_425J2_127_3477_n1035,
         DP_OP_425J2_127_3477_n1034, DP_OP_425J2_127_3477_n1033,
         DP_OP_425J2_127_3477_n1032, DP_OP_425J2_127_3477_n1031,
         DP_OP_425J2_127_3477_n1030, DP_OP_425J2_127_3477_n1029,
         DP_OP_425J2_127_3477_n1028, DP_OP_425J2_127_3477_n1027,
         DP_OP_425J2_127_3477_n1026, DP_OP_425J2_127_3477_n1025,
         DP_OP_425J2_127_3477_n1024, DP_OP_425J2_127_3477_n1023,
         DP_OP_425J2_127_3477_n1022, DP_OP_425J2_127_3477_n1021,
         DP_OP_425J2_127_3477_n1020, DP_OP_425J2_127_3477_n1019,
         DP_OP_425J2_127_3477_n1018, DP_OP_425J2_127_3477_n1017,
         DP_OP_425J2_127_3477_n1016, DP_OP_425J2_127_3477_n1015,
         DP_OP_425J2_127_3477_n1014, DP_OP_425J2_127_3477_n1013,
         DP_OP_425J2_127_3477_n1012, DP_OP_425J2_127_3477_n1011,
         DP_OP_425J2_127_3477_n1010, DP_OP_425J2_127_3477_n1009,
         DP_OP_425J2_127_3477_n1008, DP_OP_425J2_127_3477_n1007,
         DP_OP_425J2_127_3477_n1006, DP_OP_425J2_127_3477_n1005,
         DP_OP_425J2_127_3477_n1004, DP_OP_425J2_127_3477_n1003,
         DP_OP_425J2_127_3477_n1002, DP_OP_425J2_127_3477_n1001,
         DP_OP_425J2_127_3477_n1000, DP_OP_425J2_127_3477_n999,
         DP_OP_425J2_127_3477_n998, DP_OP_425J2_127_3477_n997,
         DP_OP_425J2_127_3477_n996, DP_OP_425J2_127_3477_n995,
         DP_OP_425J2_127_3477_n994, DP_OP_425J2_127_3477_n993,
         DP_OP_425J2_127_3477_n992, DP_OP_425J2_127_3477_n991,
         DP_OP_425J2_127_3477_n990, DP_OP_425J2_127_3477_n989,
         DP_OP_425J2_127_3477_n988, DP_OP_425J2_127_3477_n987,
         DP_OP_425J2_127_3477_n986, DP_OP_425J2_127_3477_n985,
         DP_OP_425J2_127_3477_n984, DP_OP_425J2_127_3477_n983,
         DP_OP_425J2_127_3477_n982, DP_OP_425J2_127_3477_n981,
         DP_OP_425J2_127_3477_n980, DP_OP_425J2_127_3477_n979,
         DP_OP_425J2_127_3477_n978, DP_OP_425J2_127_3477_n977,
         DP_OP_425J2_127_3477_n976, DP_OP_425J2_127_3477_n975,
         DP_OP_425J2_127_3477_n974, DP_OP_425J2_127_3477_n973,
         DP_OP_425J2_127_3477_n972, DP_OP_425J2_127_3477_n971,
         DP_OP_425J2_127_3477_n970, DP_OP_425J2_127_3477_n969,
         DP_OP_425J2_127_3477_n968, DP_OP_425J2_127_3477_n967,
         DP_OP_425J2_127_3477_n966, DP_OP_425J2_127_3477_n965,
         DP_OP_425J2_127_3477_n964, DP_OP_425J2_127_3477_n963,
         DP_OP_425J2_127_3477_n962, DP_OP_425J2_127_3477_n961,
         DP_OP_425J2_127_3477_n960, DP_OP_425J2_127_3477_n959,
         DP_OP_425J2_127_3477_n958, DP_OP_425J2_127_3477_n957,
         DP_OP_425J2_127_3477_n956, DP_OP_425J2_127_3477_n955,
         DP_OP_425J2_127_3477_n954, DP_OP_425J2_127_3477_n953,
         DP_OP_425J2_127_3477_n952, DP_OP_425J2_127_3477_n951,
         DP_OP_425J2_127_3477_n950, DP_OP_425J2_127_3477_n949,
         DP_OP_425J2_127_3477_n948, DP_OP_425J2_127_3477_n947,
         DP_OP_425J2_127_3477_n946, DP_OP_425J2_127_3477_n945,
         DP_OP_425J2_127_3477_n944, DP_OP_425J2_127_3477_n943,
         DP_OP_425J2_127_3477_n942, DP_OP_425J2_127_3477_n941,
         DP_OP_425J2_127_3477_n940, DP_OP_425J2_127_3477_n939,
         DP_OP_425J2_127_3477_n938, DP_OP_425J2_127_3477_n937,
         DP_OP_425J2_127_3477_n936, DP_OP_425J2_127_3477_n935,
         DP_OP_425J2_127_3477_n934, DP_OP_425J2_127_3477_n933,
         DP_OP_425J2_127_3477_n932, DP_OP_425J2_127_3477_n931,
         DP_OP_425J2_127_3477_n930, DP_OP_425J2_127_3477_n929,
         DP_OP_425J2_127_3477_n928, DP_OP_425J2_127_3477_n927,
         DP_OP_425J2_127_3477_n926, DP_OP_425J2_127_3477_n925,
         DP_OP_425J2_127_3477_n924, DP_OP_425J2_127_3477_n923,
         DP_OP_425J2_127_3477_n922, DP_OP_425J2_127_3477_n921,
         DP_OP_425J2_127_3477_n920, DP_OP_425J2_127_3477_n919,
         DP_OP_425J2_127_3477_n918, DP_OP_425J2_127_3477_n917,
         DP_OP_425J2_127_3477_n916, DP_OP_425J2_127_3477_n915,
         DP_OP_425J2_127_3477_n914, DP_OP_425J2_127_3477_n913,
         DP_OP_425J2_127_3477_n912, DP_OP_425J2_127_3477_n911,
         DP_OP_425J2_127_3477_n910, DP_OP_425J2_127_3477_n909,
         DP_OP_425J2_127_3477_n908, DP_OP_425J2_127_3477_n907,
         DP_OP_425J2_127_3477_n906, DP_OP_425J2_127_3477_n905,
         DP_OP_425J2_127_3477_n904, DP_OP_425J2_127_3477_n903,
         DP_OP_425J2_127_3477_n902, DP_OP_425J2_127_3477_n901,
         DP_OP_425J2_127_3477_n900, DP_OP_425J2_127_3477_n899,
         DP_OP_425J2_127_3477_n898, DP_OP_425J2_127_3477_n897,
         DP_OP_425J2_127_3477_n896, DP_OP_425J2_127_3477_n895,
         DP_OP_425J2_127_3477_n894, DP_OP_425J2_127_3477_n893,
         DP_OP_425J2_127_3477_n892, DP_OP_425J2_127_3477_n891,
         DP_OP_425J2_127_3477_n890, DP_OP_425J2_127_3477_n889,
         DP_OP_425J2_127_3477_n888, DP_OP_425J2_127_3477_n887,
         DP_OP_425J2_127_3477_n886, DP_OP_425J2_127_3477_n885,
         DP_OP_425J2_127_3477_n884, DP_OP_425J2_127_3477_n883,
         DP_OP_425J2_127_3477_n882, DP_OP_425J2_127_3477_n881,
         DP_OP_425J2_127_3477_n880, DP_OP_425J2_127_3477_n879,
         DP_OP_425J2_127_3477_n878, DP_OP_425J2_127_3477_n877,
         DP_OP_425J2_127_3477_n876, DP_OP_425J2_127_3477_n875,
         DP_OP_425J2_127_3477_n874, DP_OP_425J2_127_3477_n873,
         DP_OP_425J2_127_3477_n872, DP_OP_425J2_127_3477_n871,
         DP_OP_425J2_127_3477_n870, DP_OP_425J2_127_3477_n869,
         DP_OP_425J2_127_3477_n868, DP_OP_425J2_127_3477_n867,
         DP_OP_425J2_127_3477_n866, DP_OP_425J2_127_3477_n865,
         DP_OP_425J2_127_3477_n864, DP_OP_425J2_127_3477_n863,
         DP_OP_425J2_127_3477_n862, DP_OP_425J2_127_3477_n861,
         DP_OP_425J2_127_3477_n860, DP_OP_425J2_127_3477_n859,
         DP_OP_425J2_127_3477_n858, DP_OP_425J2_127_3477_n857,
         DP_OP_425J2_127_3477_n856, DP_OP_425J2_127_3477_n855,
         DP_OP_425J2_127_3477_n854, DP_OP_425J2_127_3477_n853,
         DP_OP_425J2_127_3477_n852, DP_OP_425J2_127_3477_n851,
         DP_OP_425J2_127_3477_n850, DP_OP_425J2_127_3477_n849,
         DP_OP_425J2_127_3477_n848, DP_OP_425J2_127_3477_n847,
         DP_OP_425J2_127_3477_n846, DP_OP_425J2_127_3477_n845,
         DP_OP_425J2_127_3477_n844, DP_OP_425J2_127_3477_n843,
         DP_OP_425J2_127_3477_n842, DP_OP_425J2_127_3477_n841,
         DP_OP_425J2_127_3477_n840, DP_OP_425J2_127_3477_n839,
         DP_OP_425J2_127_3477_n838, DP_OP_425J2_127_3477_n837,
         DP_OP_425J2_127_3477_n836, DP_OP_425J2_127_3477_n835,
         DP_OP_425J2_127_3477_n834, DP_OP_425J2_127_3477_n833,
         DP_OP_425J2_127_3477_n832, DP_OP_425J2_127_3477_n831,
         DP_OP_425J2_127_3477_n830, DP_OP_425J2_127_3477_n829,
         DP_OP_425J2_127_3477_n828, DP_OP_425J2_127_3477_n827,
         DP_OP_425J2_127_3477_n826, DP_OP_425J2_127_3477_n825,
         DP_OP_425J2_127_3477_n824, DP_OP_425J2_127_3477_n823,
         DP_OP_425J2_127_3477_n822, DP_OP_425J2_127_3477_n821,
         DP_OP_425J2_127_3477_n820, DP_OP_425J2_127_3477_n819,
         DP_OP_425J2_127_3477_n818, DP_OP_425J2_127_3477_n817,
         DP_OP_425J2_127_3477_n816, DP_OP_425J2_127_3477_n815,
         DP_OP_425J2_127_3477_n814, DP_OP_425J2_127_3477_n813,
         DP_OP_425J2_127_3477_n812, DP_OP_425J2_127_3477_n811,
         DP_OP_425J2_127_3477_n810, DP_OP_425J2_127_3477_n809,
         DP_OP_425J2_127_3477_n808, DP_OP_425J2_127_3477_n807,
         DP_OP_425J2_127_3477_n806, DP_OP_425J2_127_3477_n805,
         DP_OP_425J2_127_3477_n804, DP_OP_425J2_127_3477_n803,
         DP_OP_425J2_127_3477_n802, DP_OP_425J2_127_3477_n801,
         DP_OP_425J2_127_3477_n800, DP_OP_425J2_127_3477_n799,
         DP_OP_425J2_127_3477_n798, DP_OP_425J2_127_3477_n797,
         DP_OP_425J2_127_3477_n796, DP_OP_425J2_127_3477_n795,
         DP_OP_425J2_127_3477_n794, DP_OP_425J2_127_3477_n793,
         DP_OP_425J2_127_3477_n792, DP_OP_425J2_127_3477_n791,
         DP_OP_425J2_127_3477_n790, DP_OP_425J2_127_3477_n789,
         DP_OP_425J2_127_3477_n788, DP_OP_425J2_127_3477_n787,
         DP_OP_425J2_127_3477_n786, DP_OP_425J2_127_3477_n785,
         DP_OP_425J2_127_3477_n784, DP_OP_425J2_127_3477_n783,
         DP_OP_425J2_127_3477_n782, DP_OP_425J2_127_3477_n781,
         DP_OP_425J2_127_3477_n780, DP_OP_425J2_127_3477_n779,
         DP_OP_425J2_127_3477_n778, DP_OP_425J2_127_3477_n777,
         DP_OP_425J2_127_3477_n776, DP_OP_425J2_127_3477_n775,
         DP_OP_425J2_127_3477_n774, DP_OP_425J2_127_3477_n773,
         DP_OP_425J2_127_3477_n772, DP_OP_425J2_127_3477_n771,
         DP_OP_425J2_127_3477_n770, DP_OP_425J2_127_3477_n769,
         DP_OP_425J2_127_3477_n768, DP_OP_425J2_127_3477_n767,
         DP_OP_425J2_127_3477_n766, DP_OP_425J2_127_3477_n765,
         DP_OP_425J2_127_3477_n764, DP_OP_425J2_127_3477_n763,
         DP_OP_425J2_127_3477_n762, DP_OP_425J2_127_3477_n761,
         DP_OP_425J2_127_3477_n760, DP_OP_425J2_127_3477_n759,
         DP_OP_425J2_127_3477_n758, DP_OP_425J2_127_3477_n757,
         DP_OP_425J2_127_3477_n756, DP_OP_425J2_127_3477_n755,
         DP_OP_425J2_127_3477_n754, DP_OP_425J2_127_3477_n753,
         DP_OP_425J2_127_3477_n752, DP_OP_425J2_127_3477_n751,
         DP_OP_425J2_127_3477_n750, DP_OP_425J2_127_3477_n749,
         DP_OP_425J2_127_3477_n748, DP_OP_425J2_127_3477_n747,
         DP_OP_425J2_127_3477_n746, DP_OP_425J2_127_3477_n745,
         DP_OP_425J2_127_3477_n744, DP_OP_425J2_127_3477_n743,
         DP_OP_425J2_127_3477_n742, DP_OP_425J2_127_3477_n741,
         DP_OP_425J2_127_3477_n740, DP_OP_425J2_127_3477_n739,
         DP_OP_425J2_127_3477_n738, DP_OP_425J2_127_3477_n737,
         DP_OP_425J2_127_3477_n736, DP_OP_425J2_127_3477_n735,
         DP_OP_425J2_127_3477_n734, DP_OP_425J2_127_3477_n733,
         DP_OP_425J2_127_3477_n732, DP_OP_425J2_127_3477_n731,
         DP_OP_425J2_127_3477_n730, DP_OP_425J2_127_3477_n729,
         DP_OP_425J2_127_3477_n728, DP_OP_425J2_127_3477_n727,
         DP_OP_425J2_127_3477_n726, DP_OP_425J2_127_3477_n725,
         DP_OP_425J2_127_3477_n724, DP_OP_425J2_127_3477_n723,
         DP_OP_425J2_127_3477_n722, DP_OP_425J2_127_3477_n721,
         DP_OP_425J2_127_3477_n720, DP_OP_425J2_127_3477_n719,
         DP_OP_425J2_127_3477_n718, DP_OP_425J2_127_3477_n717,
         DP_OP_425J2_127_3477_n716, DP_OP_425J2_127_3477_n715,
         DP_OP_425J2_127_3477_n714, DP_OP_425J2_127_3477_n713,
         DP_OP_425J2_127_3477_n712, DP_OP_425J2_127_3477_n711,
         DP_OP_425J2_127_3477_n710, DP_OP_425J2_127_3477_n709,
         DP_OP_425J2_127_3477_n708, DP_OP_425J2_127_3477_n707,
         DP_OP_425J2_127_3477_n706, DP_OP_425J2_127_3477_n705,
         DP_OP_425J2_127_3477_n704, DP_OP_425J2_127_3477_n703,
         DP_OP_425J2_127_3477_n702, DP_OP_425J2_127_3477_n701,
         DP_OP_425J2_127_3477_n700, DP_OP_425J2_127_3477_n699,
         DP_OP_425J2_127_3477_n698, DP_OP_425J2_127_3477_n697,
         DP_OP_425J2_127_3477_n696, DP_OP_425J2_127_3477_n695,
         DP_OP_425J2_127_3477_n694, DP_OP_425J2_127_3477_n693,
         DP_OP_425J2_127_3477_n692, DP_OP_425J2_127_3477_n691,
         DP_OP_425J2_127_3477_n690, DP_OP_425J2_127_3477_n689,
         DP_OP_425J2_127_3477_n688, DP_OP_425J2_127_3477_n687,
         DP_OP_425J2_127_3477_n686, DP_OP_425J2_127_3477_n685,
         DP_OP_425J2_127_3477_n684, DP_OP_425J2_127_3477_n683,
         DP_OP_425J2_127_3477_n682, DP_OP_425J2_127_3477_n681,
         DP_OP_425J2_127_3477_n680, DP_OP_425J2_127_3477_n679,
         DP_OP_425J2_127_3477_n678, DP_OP_425J2_127_3477_n677,
         DP_OP_425J2_127_3477_n676, DP_OP_425J2_127_3477_n675,
         DP_OP_425J2_127_3477_n674, DP_OP_425J2_127_3477_n673,
         DP_OP_425J2_127_3477_n672, DP_OP_425J2_127_3477_n671,
         DP_OP_425J2_127_3477_n670, DP_OP_425J2_127_3477_n669,
         DP_OP_425J2_127_3477_n668, DP_OP_425J2_127_3477_n667,
         DP_OP_425J2_127_3477_n666, DP_OP_425J2_127_3477_n665,
         DP_OP_425J2_127_3477_n664, DP_OP_425J2_127_3477_n663,
         DP_OP_425J2_127_3477_n662, DP_OP_425J2_127_3477_n661,
         DP_OP_425J2_127_3477_n660, DP_OP_425J2_127_3477_n659,
         DP_OP_425J2_127_3477_n658, DP_OP_425J2_127_3477_n657,
         DP_OP_425J2_127_3477_n656, DP_OP_425J2_127_3477_n655,
         DP_OP_425J2_127_3477_n654, DP_OP_425J2_127_3477_n653,
         DP_OP_425J2_127_3477_n652, DP_OP_425J2_127_3477_n651,
         DP_OP_425J2_127_3477_n650, DP_OP_425J2_127_3477_n649,
         DP_OP_425J2_127_3477_n648, DP_OP_425J2_127_3477_n647,
         DP_OP_425J2_127_3477_n646, DP_OP_425J2_127_3477_n645,
         DP_OP_425J2_127_3477_n644, DP_OP_425J2_127_3477_n643,
         DP_OP_425J2_127_3477_n642, DP_OP_425J2_127_3477_n641,
         DP_OP_425J2_127_3477_n640, DP_OP_425J2_127_3477_n639,
         DP_OP_425J2_127_3477_n638, DP_OP_425J2_127_3477_n637,
         DP_OP_425J2_127_3477_n636, DP_OP_425J2_127_3477_n635,
         DP_OP_425J2_127_3477_n634, DP_OP_425J2_127_3477_n633,
         DP_OP_425J2_127_3477_n632, DP_OP_425J2_127_3477_n631,
         DP_OP_425J2_127_3477_n630, DP_OP_425J2_127_3477_n629,
         DP_OP_425J2_127_3477_n628, DP_OP_425J2_127_3477_n627,
         DP_OP_425J2_127_3477_n626, DP_OP_425J2_127_3477_n625,
         DP_OP_425J2_127_3477_n624, DP_OP_425J2_127_3477_n623,
         DP_OP_425J2_127_3477_n622, DP_OP_425J2_127_3477_n621,
         DP_OP_425J2_127_3477_n620, DP_OP_425J2_127_3477_n619,
         DP_OP_425J2_127_3477_n618, DP_OP_425J2_127_3477_n617,
         DP_OP_425J2_127_3477_n616, DP_OP_425J2_127_3477_n615,
         DP_OP_425J2_127_3477_n614, DP_OP_425J2_127_3477_n613,
         DP_OP_425J2_127_3477_n612, DP_OP_425J2_127_3477_n611,
         DP_OP_425J2_127_3477_n610, DP_OP_425J2_127_3477_n609,
         DP_OP_425J2_127_3477_n608, DP_OP_425J2_127_3477_n607,
         DP_OP_425J2_127_3477_n606, DP_OP_425J2_127_3477_n605,
         DP_OP_425J2_127_3477_n604, DP_OP_425J2_127_3477_n603,
         DP_OP_425J2_127_3477_n602, DP_OP_425J2_127_3477_n601,
         DP_OP_425J2_127_3477_n600, DP_OP_425J2_127_3477_n599,
         DP_OP_425J2_127_3477_n598, DP_OP_425J2_127_3477_n597,
         DP_OP_425J2_127_3477_n596, DP_OP_425J2_127_3477_n595,
         DP_OP_425J2_127_3477_n594, DP_OP_425J2_127_3477_n593,
         DP_OP_425J2_127_3477_n592, DP_OP_425J2_127_3477_n591,
         DP_OP_425J2_127_3477_n590, DP_OP_425J2_127_3477_n589,
         DP_OP_425J2_127_3477_n588, DP_OP_425J2_127_3477_n587,
         DP_OP_425J2_127_3477_n586, DP_OP_425J2_127_3477_n585,
         DP_OP_425J2_127_3477_n584, DP_OP_425J2_127_3477_n583,
         DP_OP_425J2_127_3477_n582, DP_OP_425J2_127_3477_n581,
         DP_OP_425J2_127_3477_n580, DP_OP_425J2_127_3477_n579,
         DP_OP_425J2_127_3477_n578, DP_OP_425J2_127_3477_n577,
         DP_OP_425J2_127_3477_n576, DP_OP_425J2_127_3477_n575,
         DP_OP_425J2_127_3477_n574, DP_OP_425J2_127_3477_n573,
         DP_OP_425J2_127_3477_n572, DP_OP_425J2_127_3477_n571,
         DP_OP_425J2_127_3477_n570, DP_OP_425J2_127_3477_n569,
         DP_OP_425J2_127_3477_n568, DP_OP_425J2_127_3477_n567,
         DP_OP_425J2_127_3477_n566, DP_OP_425J2_127_3477_n565,
         DP_OP_425J2_127_3477_n564, DP_OP_425J2_127_3477_n563,
         DP_OP_425J2_127_3477_n562, DP_OP_425J2_127_3477_n561,
         DP_OP_425J2_127_3477_n560, DP_OP_425J2_127_3477_n559,
         DP_OP_425J2_127_3477_n558, DP_OP_425J2_127_3477_n557,
         DP_OP_425J2_127_3477_n556, DP_OP_425J2_127_3477_n555,
         DP_OP_425J2_127_3477_n554, DP_OP_425J2_127_3477_n553,
         DP_OP_425J2_127_3477_n552, DP_OP_425J2_127_3477_n551,
         DP_OP_425J2_127_3477_n550, DP_OP_425J2_127_3477_n549,
         DP_OP_425J2_127_3477_n548, DP_OP_425J2_127_3477_n547,
         DP_OP_425J2_127_3477_n546, DP_OP_425J2_127_3477_n545,
         DP_OP_425J2_127_3477_n544, DP_OP_425J2_127_3477_n543,
         DP_OP_425J2_127_3477_n542, DP_OP_425J2_127_3477_n541,
         DP_OP_425J2_127_3477_n540, DP_OP_425J2_127_3477_n539,
         DP_OP_425J2_127_3477_n538, DP_OP_425J2_127_3477_n537,
         DP_OP_425J2_127_3477_n536, DP_OP_425J2_127_3477_n535,
         DP_OP_425J2_127_3477_n534, DP_OP_425J2_127_3477_n533,
         DP_OP_425J2_127_3477_n532, DP_OP_425J2_127_3477_n531,
         DP_OP_425J2_127_3477_n530, DP_OP_425J2_127_3477_n529,
         DP_OP_425J2_127_3477_n528, DP_OP_425J2_127_3477_n527,
         DP_OP_425J2_127_3477_n526, DP_OP_425J2_127_3477_n525,
         DP_OP_425J2_127_3477_n524, DP_OP_425J2_127_3477_n523,
         DP_OP_425J2_127_3477_n522, DP_OP_425J2_127_3477_n521,
         DP_OP_425J2_127_3477_n520, DP_OP_425J2_127_3477_n519,
         DP_OP_425J2_127_3477_n518, DP_OP_425J2_127_3477_n517,
         DP_OP_425J2_127_3477_n516, DP_OP_425J2_127_3477_n515,
         DP_OP_425J2_127_3477_n514, DP_OP_425J2_127_3477_n513,
         DP_OP_425J2_127_3477_n512, DP_OP_425J2_127_3477_n511,
         DP_OP_425J2_127_3477_n510, DP_OP_425J2_127_3477_n509,
         DP_OP_425J2_127_3477_n508, DP_OP_425J2_127_3477_n507,
         DP_OP_425J2_127_3477_n506, DP_OP_425J2_127_3477_n505,
         DP_OP_425J2_127_3477_n504, DP_OP_425J2_127_3477_n503,
         DP_OP_425J2_127_3477_n502, DP_OP_425J2_127_3477_n501,
         DP_OP_425J2_127_3477_n500, DP_OP_425J2_127_3477_n499,
         DP_OP_425J2_127_3477_n498, DP_OP_425J2_127_3477_n497,
         DP_OP_425J2_127_3477_n496, DP_OP_425J2_127_3477_n495,
         DP_OP_425J2_127_3477_n494, DP_OP_425J2_127_3477_n493,
         DP_OP_425J2_127_3477_n492, DP_OP_425J2_127_3477_n491,
         DP_OP_425J2_127_3477_n490, DP_OP_425J2_127_3477_n489,
         DP_OP_425J2_127_3477_n488, DP_OP_425J2_127_3477_n487,
         DP_OP_425J2_127_3477_n486, DP_OP_425J2_127_3477_n485,
         DP_OP_425J2_127_3477_n484, DP_OP_425J2_127_3477_n483,
         DP_OP_425J2_127_3477_n482, DP_OP_425J2_127_3477_n481,
         DP_OP_425J2_127_3477_n480, DP_OP_425J2_127_3477_n479,
         DP_OP_425J2_127_3477_n478, DP_OP_425J2_127_3477_n477,
         DP_OP_425J2_127_3477_n476, DP_OP_425J2_127_3477_n475,
         DP_OP_425J2_127_3477_n474, DP_OP_425J2_127_3477_n473,
         DP_OP_425J2_127_3477_n472, DP_OP_425J2_127_3477_n471,
         DP_OP_425J2_127_3477_n470, DP_OP_425J2_127_3477_n469,
         DP_OP_425J2_127_3477_n468, DP_OP_425J2_127_3477_n467,
         DP_OP_425J2_127_3477_n466, DP_OP_425J2_127_3477_n465,
         DP_OP_425J2_127_3477_n464, DP_OP_425J2_127_3477_n463,
         DP_OP_425J2_127_3477_n462, DP_OP_425J2_127_3477_n461,
         DP_OP_425J2_127_3477_n460, DP_OP_425J2_127_3477_n459,
         DP_OP_425J2_127_3477_n458, DP_OP_425J2_127_3477_n457,
         DP_OP_425J2_127_3477_n456, DP_OP_425J2_127_3477_n455,
         DP_OP_425J2_127_3477_n454, DP_OP_425J2_127_3477_n453,
         DP_OP_425J2_127_3477_n452, DP_OP_425J2_127_3477_n451,
         DP_OP_425J2_127_3477_n450, DP_OP_425J2_127_3477_n449,
         DP_OP_425J2_127_3477_n448, DP_OP_425J2_127_3477_n447,
         DP_OP_425J2_127_3477_n446, DP_OP_425J2_127_3477_n445,
         DP_OP_425J2_127_3477_n444, DP_OP_425J2_127_3477_n443,
         DP_OP_425J2_127_3477_n442, DP_OP_425J2_127_3477_n441,
         DP_OP_425J2_127_3477_n440, DP_OP_425J2_127_3477_n439,
         DP_OP_425J2_127_3477_n438, DP_OP_425J2_127_3477_n437,
         DP_OP_425J2_127_3477_n436, DP_OP_425J2_127_3477_n435,
         DP_OP_425J2_127_3477_n434, DP_OP_425J2_127_3477_n433,
         DP_OP_425J2_127_3477_n432, DP_OP_425J2_127_3477_n431,
         DP_OP_425J2_127_3477_n430, DP_OP_425J2_127_3477_n429,
         DP_OP_425J2_127_3477_n428, DP_OP_425J2_127_3477_n427,
         DP_OP_425J2_127_3477_n426, DP_OP_425J2_127_3477_n425,
         DP_OP_425J2_127_3477_n424, DP_OP_425J2_127_3477_n423,
         DP_OP_425J2_127_3477_n422, DP_OP_425J2_127_3477_n421,
         DP_OP_425J2_127_3477_n420, DP_OP_425J2_127_3477_n419,
         DP_OP_425J2_127_3477_n418, DP_OP_425J2_127_3477_n417,
         DP_OP_425J2_127_3477_n416, DP_OP_425J2_127_3477_n415,
         DP_OP_425J2_127_3477_n414, DP_OP_425J2_127_3477_n413,
         DP_OP_425J2_127_3477_n412, DP_OP_425J2_127_3477_n411,
         DP_OP_425J2_127_3477_n410, DP_OP_425J2_127_3477_n409,
         DP_OP_425J2_127_3477_n408, DP_OP_425J2_127_3477_n407,
         DP_OP_425J2_127_3477_n406, DP_OP_425J2_127_3477_n405,
         DP_OP_425J2_127_3477_n404, DP_OP_425J2_127_3477_n403,
         DP_OP_425J2_127_3477_n402, DP_OP_425J2_127_3477_n401,
         DP_OP_425J2_127_3477_n400, DP_OP_425J2_127_3477_n399,
         DP_OP_425J2_127_3477_n398, DP_OP_425J2_127_3477_n397,
         DP_OP_425J2_127_3477_n396, DP_OP_425J2_127_3477_n395,
         DP_OP_425J2_127_3477_n394, DP_OP_425J2_127_3477_n393,
         DP_OP_425J2_127_3477_n392, DP_OP_425J2_127_3477_n391,
         DP_OP_425J2_127_3477_n390, DP_OP_425J2_127_3477_n389,
         DP_OP_425J2_127_3477_n388, DP_OP_425J2_127_3477_n387,
         DP_OP_425J2_127_3477_n386, DP_OP_425J2_127_3477_n385,
         DP_OP_425J2_127_3477_n384, DP_OP_425J2_127_3477_n383,
         DP_OP_425J2_127_3477_n382, DP_OP_425J2_127_3477_n381,
         DP_OP_425J2_127_3477_n380, DP_OP_425J2_127_3477_n379,
         DP_OP_425J2_127_3477_n378, DP_OP_425J2_127_3477_n377,
         DP_OP_425J2_127_3477_n376, DP_OP_425J2_127_3477_n375,
         DP_OP_425J2_127_3477_n374, DP_OP_425J2_127_3477_n373,
         DP_OP_425J2_127_3477_n372, DP_OP_425J2_127_3477_n371,
         DP_OP_425J2_127_3477_n370, DP_OP_425J2_127_3477_n369,
         DP_OP_425J2_127_3477_n368, DP_OP_425J2_127_3477_n367,
         DP_OP_425J2_127_3477_n366, DP_OP_425J2_127_3477_n365,
         DP_OP_425J2_127_3477_n364, DP_OP_425J2_127_3477_n363,
         DP_OP_425J2_127_3477_n362, DP_OP_425J2_127_3477_n361,
         DP_OP_425J2_127_3477_n360, DP_OP_425J2_127_3477_n359,
         DP_OP_425J2_127_3477_n358, DP_OP_425J2_127_3477_n357,
         DP_OP_425J2_127_3477_n356, DP_OP_425J2_127_3477_n355,
         DP_OP_425J2_127_3477_n354, DP_OP_425J2_127_3477_n353,
         DP_OP_425J2_127_3477_n352, DP_OP_425J2_127_3477_n351,
         DP_OP_425J2_127_3477_n350, DP_OP_425J2_127_3477_n349,
         DP_OP_425J2_127_3477_n348, DP_OP_425J2_127_3477_n347,
         DP_OP_425J2_127_3477_n346, DP_OP_425J2_127_3477_n345,
         DP_OP_425J2_127_3477_n344, DP_OP_425J2_127_3477_n343,
         DP_OP_425J2_127_3477_n342, DP_OP_425J2_127_3477_n341,
         DP_OP_425J2_127_3477_n340, DP_OP_425J2_127_3477_n339,
         DP_OP_425J2_127_3477_n338, DP_OP_425J2_127_3477_n337,
         DP_OP_425J2_127_3477_n336, DP_OP_425J2_127_3477_n335,
         DP_OP_425J2_127_3477_n334, DP_OP_425J2_127_3477_n333,
         DP_OP_425J2_127_3477_n332, DP_OP_425J2_127_3477_n331,
         DP_OP_425J2_127_3477_n330, DP_OP_425J2_127_3477_n329,
         DP_OP_425J2_127_3477_n328, DP_OP_425J2_127_3477_n327,
         DP_OP_425J2_127_3477_n326, DP_OP_425J2_127_3477_n325,
         DP_OP_425J2_127_3477_n324, DP_OP_425J2_127_3477_n323,
         DP_OP_425J2_127_3477_n322, DP_OP_425J2_127_3477_n321,
         DP_OP_425J2_127_3477_n320, DP_OP_425J2_127_3477_n319,
         DP_OP_425J2_127_3477_n318, DP_OP_425J2_127_3477_n317,
         DP_OP_425J2_127_3477_n316, DP_OP_425J2_127_3477_n315,
         DP_OP_425J2_127_3477_n314, DP_OP_425J2_127_3477_n313,
         DP_OP_425J2_127_3477_n312, DP_OP_425J2_127_3477_n311,
         DP_OP_425J2_127_3477_n310, DP_OP_425J2_127_3477_n309,
         DP_OP_425J2_127_3477_n308, DP_OP_425J2_127_3477_n307,
         DP_OP_425J2_127_3477_n306, DP_OP_425J2_127_3477_n305,
         DP_OP_425J2_127_3477_n304, DP_OP_425J2_127_3477_n303,
         DP_OP_425J2_127_3477_n302, DP_OP_425J2_127_3477_n301,
         DP_OP_425J2_127_3477_n300, DP_OP_425J2_127_3477_n299,
         DP_OP_425J2_127_3477_n298, DP_OP_425J2_127_3477_n297,
         DP_OP_425J2_127_3477_n296, DP_OP_425J2_127_3477_n295,
         DP_OP_425J2_127_3477_n294, DP_OP_425J2_127_3477_n293,
         DP_OP_425J2_127_3477_n292, DP_OP_425J2_127_3477_n291,
         DP_OP_425J2_127_3477_n290, DP_OP_425J2_127_3477_n289,
         DP_OP_425J2_127_3477_n288, DP_OP_425J2_127_3477_n287,
         DP_OP_425J2_127_3477_n286, DP_OP_425J2_127_3477_n285,
         DP_OP_425J2_127_3477_n284, DP_OP_425J2_127_3477_n283,
         DP_OP_425J2_127_3477_n282, DP_OP_425J2_127_3477_n281,
         DP_OP_425J2_127_3477_n280, DP_OP_425J2_127_3477_n279,
         DP_OP_425J2_127_3477_n278, DP_OP_425J2_127_3477_n277,
         DP_OP_425J2_127_3477_n276, DP_OP_425J2_127_3477_n275,
         DP_OP_425J2_127_3477_n274, DP_OP_425J2_127_3477_n273,
         DP_OP_425J2_127_3477_n272, DP_OP_425J2_127_3477_n271,
         DP_OP_425J2_127_3477_n270, DP_OP_425J2_127_3477_n269,
         DP_OP_425J2_127_3477_n268, DP_OP_425J2_127_3477_n267,
         DP_OP_425J2_127_3477_n266, DP_OP_425J2_127_3477_n265,
         DP_OP_425J2_127_3477_n264, DP_OP_425J2_127_3477_n263,
         DP_OP_425J2_127_3477_n262, DP_OP_425J2_127_3477_n261,
         DP_OP_425J2_127_3477_n260, DP_OP_425J2_127_3477_n259,
         DP_OP_425J2_127_3477_n258, DP_OP_425J2_127_3477_n257,
         DP_OP_425J2_127_3477_n256, DP_OP_425J2_127_3477_n255,
         DP_OP_425J2_127_3477_n254, DP_OP_425J2_127_3477_n253,
         DP_OP_425J2_127_3477_n252, DP_OP_425J2_127_3477_n241,
         DP_OP_425J2_127_3477_n240, DP_OP_425J2_127_3477_n237,
         DP_OP_425J2_127_3477_n236, DP_OP_425J2_127_3477_n235,
         DP_OP_425J2_127_3477_n234, DP_OP_425J2_127_3477_n233,
         DP_OP_425J2_127_3477_n231, DP_OP_425J2_127_3477_n229,
         DP_OP_425J2_127_3477_n227, DP_OP_425J2_127_3477_n219,
         DP_OP_425J2_127_3477_n218, DP_OP_425J2_127_3477_n217,
         DP_OP_425J2_127_3477_n216, DP_OP_425J2_127_3477_n215,
         DP_OP_425J2_127_3477_n211, DP_OP_425J2_127_3477_n210,
         DP_OP_425J2_127_3477_n209, DP_OP_425J2_127_3477_n208,
         DP_OP_425J2_127_3477_n207, DP_OP_425J2_127_3477_n203,
         DP_OP_425J2_127_3477_n202, DP_OP_425J2_127_3477_n201,
         DP_OP_425J2_127_3477_n200, DP_OP_425J2_127_3477_n199,
         DP_OP_425J2_127_3477_n195, DP_OP_425J2_127_3477_n194,
         DP_OP_425J2_127_3477_n193, DP_OP_425J2_127_3477_n192,
         DP_OP_425J2_127_3477_n191, DP_OP_425J2_127_3477_n190,
         DP_OP_425J2_127_3477_n189, DP_OP_425J2_127_3477_n187,
         DP_OP_425J2_127_3477_n186, DP_OP_425J2_127_3477_n185,
         DP_OP_425J2_127_3477_n184, DP_OP_425J2_127_3477_n183,
         DP_OP_425J2_127_3477_n182, DP_OP_425J2_127_3477_n181,
         DP_OP_425J2_127_3477_n180, DP_OP_425J2_127_3477_n179,
         DP_OP_425J2_127_3477_n177, DP_OP_425J2_127_3477_n176,
         DP_OP_425J2_127_3477_n175, DP_OP_425J2_127_3477_n174,
         DP_OP_425J2_127_3477_n173, DP_OP_425J2_127_3477_n172,
         DP_OP_425J2_127_3477_n171, DP_OP_425J2_127_3477_n170,
         DP_OP_425J2_127_3477_n168, DP_OP_425J2_127_3477_n167,
         DP_OP_425J2_127_3477_n166, DP_OP_425J2_127_3477_n165,
         DP_OP_425J2_127_3477_n164, DP_OP_425J2_127_3477_n163,
         DP_OP_425J2_127_3477_n162, DP_OP_425J2_127_3477_n161,
         DP_OP_425J2_127_3477_n158, DP_OP_425J2_127_3477_n152,
         DP_OP_425J2_127_3477_n151, DP_OP_425J2_127_3477_n149,
         DP_OP_425J2_127_3477_n148, DP_OP_425J2_127_3477_n145,
         DP_OP_425J2_127_3477_n144, DP_OP_425J2_127_3477_n141,
         DP_OP_425J2_127_3477_n140, DP_OP_425J2_127_3477_n137,
         DP_OP_425J2_127_3477_n136, DP_OP_425J2_127_3477_n135,
         DP_OP_425J2_127_3477_n133, DP_OP_425J2_127_3477_n132,
         DP_OP_425J2_127_3477_n131, DP_OP_425J2_127_3477_n130,
         DP_OP_425J2_127_3477_n129, DP_OP_425J2_127_3477_n128,
         DP_OP_425J2_127_3477_n127, DP_OP_425J2_127_3477_n126,
         DP_OP_425J2_127_3477_n125, DP_OP_425J2_127_3477_n124,
         DP_OP_425J2_127_3477_n123, DP_OP_425J2_127_3477_n119,
         DP_OP_425J2_127_3477_n118, DP_OP_425J2_127_3477_n116,
         DP_OP_425J2_127_3477_n115, DP_OP_425J2_127_3477_n114,
         DP_OP_425J2_127_3477_n113, DP_OP_425J2_127_3477_n112,
         DP_OP_425J2_127_3477_n111, DP_OP_425J2_127_3477_n109,
         DP_OP_425J2_127_3477_n105, DP_OP_425J2_127_3477_n104,
         DP_OP_425J2_127_3477_n102, DP_OP_425J2_127_3477_n101,
         DP_OP_425J2_127_3477_n100, DP_OP_425J2_127_3477_n99,
         DP_OP_425J2_127_3477_n98, DP_OP_425J2_127_3477_n97,
         DP_OP_425J2_127_3477_n95, DP_OP_425J2_127_3477_n91,
         DP_OP_425J2_127_3477_n90, DP_OP_425J2_127_3477_n88,
         DP_OP_425J2_127_3477_n87, DP_OP_425J2_127_3477_n86,
         DP_OP_425J2_127_3477_n85, DP_OP_425J2_127_3477_n84,
         DP_OP_425J2_127_3477_n83, DP_OP_425J2_127_3477_n81,
         DP_OP_425J2_127_3477_n76, DP_OP_425J2_127_3477_n75,
         DP_OP_425J2_127_3477_n74, DP_OP_425J2_127_3477_n73,
         DP_OP_425J2_127_3477_n72, DP_OP_425J2_127_3477_n70,
         DP_OP_425J2_127_3477_n65, DP_OP_425J2_127_3477_n63,
         DP_OP_425J2_127_3477_n62, DP_OP_425J2_127_3477_n61,
         DP_OP_425J2_127_3477_n59, DP_OP_425J2_127_3477_n58,
         DP_OP_425J2_127_3477_n57, DP_OP_425J2_127_3477_n56,
         DP_OP_425J2_127_3477_n55, DP_OP_425J2_127_3477_n52,
         DP_OP_425J2_127_3477_n48, DP_OP_425J2_127_3477_n47,
         DP_OP_425J2_127_3477_n45, DP_OP_425J2_127_3477_n44,
         DP_OP_425J2_127_3477_n43, DP_OP_425J2_127_3477_n42,
         DP_OP_425J2_127_3477_n41, DP_OP_425J2_127_3477_n40,
         DP_OP_425J2_127_3477_n39, DP_OP_425J2_127_3477_n37,
         DP_OP_425J2_127_3477_n25, DP_OP_425J2_127_3477_n20,
         DP_OP_425J2_127_3477_n19, DP_OP_425J2_127_3477_n18,
         DP_OP_425J2_127_3477_n17, DP_OP_425J2_127_3477_n4,
         DP_OP_425J2_127_3477_n3, DP_OP_425J2_127_3477_n2,
         DP_OP_424J2_126_3477_n3016, DP_OP_424J2_126_3477_n3015,
         DP_OP_424J2_126_3477_n3013, DP_OP_424J2_126_3477_n3012,
         DP_OP_424J2_126_3477_n3011, DP_OP_424J2_126_3477_n3010,
         DP_OP_424J2_126_3477_n3009, DP_OP_424J2_126_3477_n3008,
         DP_OP_424J2_126_3477_n3007, DP_OP_424J2_126_3477_n3006,
         DP_OP_424J2_126_3477_n3005, DP_OP_424J2_126_3477_n3004,
         DP_OP_424J2_126_3477_n3003, DP_OP_424J2_126_3477_n3002,
         DP_OP_424J2_126_3477_n3001, DP_OP_424J2_126_3477_n3000,
         DP_OP_424J2_126_3477_n2999, DP_OP_424J2_126_3477_n2998,
         DP_OP_424J2_126_3477_n2997, DP_OP_424J2_126_3477_n2996,
         DP_OP_424J2_126_3477_n2995, DP_OP_424J2_126_3477_n2994,
         DP_OP_424J2_126_3477_n2993, DP_OP_424J2_126_3477_n2992,
         DP_OP_424J2_126_3477_n2991, DP_OP_424J2_126_3477_n2990,
         DP_OP_424J2_126_3477_n2989, DP_OP_424J2_126_3477_n2988,
         DP_OP_424J2_126_3477_n2987, DP_OP_424J2_126_3477_n2986,
         DP_OP_424J2_126_3477_n2985, DP_OP_424J2_126_3477_n2984,
         DP_OP_424J2_126_3477_n2983, DP_OP_424J2_126_3477_n2982,
         DP_OP_424J2_126_3477_n2981, DP_OP_424J2_126_3477_n2980,
         DP_OP_424J2_126_3477_n2979, DP_OP_424J2_126_3477_n2978,
         DP_OP_424J2_126_3477_n2977, DP_OP_424J2_126_3477_n2976,
         DP_OP_424J2_126_3477_n2975, DP_OP_424J2_126_3477_n2970,
         DP_OP_424J2_126_3477_n2969, DP_OP_424J2_126_3477_n2967,
         DP_OP_424J2_126_3477_n2964, DP_OP_424J2_126_3477_n2963,
         DP_OP_424J2_126_3477_n2962, DP_OP_424J2_126_3477_n2961,
         DP_OP_424J2_126_3477_n2960, DP_OP_424J2_126_3477_n2959,
         DP_OP_424J2_126_3477_n2958, DP_OP_424J2_126_3477_n2957,
         DP_OP_424J2_126_3477_n2956, DP_OP_424J2_126_3477_n2955,
         DP_OP_424J2_126_3477_n2954, DP_OP_424J2_126_3477_n2953,
         DP_OP_424J2_126_3477_n2952, DP_OP_424J2_126_3477_n2951,
         DP_OP_424J2_126_3477_n2950, DP_OP_424J2_126_3477_n2949,
         DP_OP_424J2_126_3477_n2948, DP_OP_424J2_126_3477_n2947,
         DP_OP_424J2_126_3477_n2946, DP_OP_424J2_126_3477_n2945,
         DP_OP_424J2_126_3477_n2944, DP_OP_424J2_126_3477_n2943,
         DP_OP_424J2_126_3477_n2942, DP_OP_424J2_126_3477_n2941,
         DP_OP_424J2_126_3477_n2940, DP_OP_424J2_126_3477_n2939,
         DP_OP_424J2_126_3477_n2938, DP_OP_424J2_126_3477_n2937,
         DP_OP_424J2_126_3477_n2936, DP_OP_424J2_126_3477_n2935,
         DP_OP_424J2_126_3477_n2934, DP_OP_424J2_126_3477_n2933,
         DP_OP_424J2_126_3477_n2932, DP_OP_424J2_126_3477_n2929,
         DP_OP_424J2_126_3477_n2927, DP_OP_424J2_126_3477_n2926,
         DP_OP_424J2_126_3477_n2925, DP_OP_424J2_126_3477_n2924,
         DP_OP_424J2_126_3477_n2923, DP_OP_424J2_126_3477_n2922,
         DP_OP_424J2_126_3477_n2921, DP_OP_424J2_126_3477_n2920,
         DP_OP_424J2_126_3477_n2919, DP_OP_424J2_126_3477_n2918,
         DP_OP_424J2_126_3477_n2917, DP_OP_424J2_126_3477_n2916,
         DP_OP_424J2_126_3477_n2915, DP_OP_424J2_126_3477_n2914,
         DP_OP_424J2_126_3477_n2913, DP_OP_424J2_126_3477_n2912,
         DP_OP_424J2_126_3477_n2911, DP_OP_424J2_126_3477_n2910,
         DP_OP_424J2_126_3477_n2909, DP_OP_424J2_126_3477_n2908,
         DP_OP_424J2_126_3477_n2907, DP_OP_424J2_126_3477_n2906,
         DP_OP_424J2_126_3477_n2905, DP_OP_424J2_126_3477_n2904,
         DP_OP_424J2_126_3477_n2903, DP_OP_424J2_126_3477_n2902,
         DP_OP_424J2_126_3477_n2901, DP_OP_424J2_126_3477_n2900,
         DP_OP_424J2_126_3477_n2899, DP_OP_424J2_126_3477_n2898,
         DP_OP_424J2_126_3477_n2897, DP_OP_424J2_126_3477_n2896,
         DP_OP_424J2_126_3477_n2895, DP_OP_424J2_126_3477_n2894,
         DP_OP_424J2_126_3477_n2893, DP_OP_424J2_126_3477_n2892,
         DP_OP_424J2_126_3477_n2891, DP_OP_424J2_126_3477_n2890,
         DP_OP_424J2_126_3477_n2889, DP_OP_424J2_126_3477_n2888,
         DP_OP_424J2_126_3477_n2887, DP_OP_424J2_126_3477_n2886,
         DP_OP_424J2_126_3477_n2885, DP_OP_424J2_126_3477_n2883,
         DP_OP_424J2_126_3477_n2880, DP_OP_424J2_126_3477_n2878,
         DP_OP_424J2_126_3477_n2877, DP_OP_424J2_126_3477_n2875,
         DP_OP_424J2_126_3477_n2874, DP_OP_424J2_126_3477_n2873,
         DP_OP_424J2_126_3477_n2872, DP_OP_424J2_126_3477_n2871,
         DP_OP_424J2_126_3477_n2870, DP_OP_424J2_126_3477_n2869,
         DP_OP_424J2_126_3477_n2868, DP_OP_424J2_126_3477_n2867,
         DP_OP_424J2_126_3477_n2866, DP_OP_424J2_126_3477_n2865,
         DP_OP_424J2_126_3477_n2864, DP_OP_424J2_126_3477_n2863,
         DP_OP_424J2_126_3477_n2862, DP_OP_424J2_126_3477_n2861,
         DP_OP_424J2_126_3477_n2860, DP_OP_424J2_126_3477_n2859,
         DP_OP_424J2_126_3477_n2858, DP_OP_424J2_126_3477_n2857,
         DP_OP_424J2_126_3477_n2856, DP_OP_424J2_126_3477_n2855,
         DP_OP_424J2_126_3477_n2854, DP_OP_424J2_126_3477_n2853,
         DP_OP_424J2_126_3477_n2852, DP_OP_424J2_126_3477_n2851,
         DP_OP_424J2_126_3477_n2850, DP_OP_424J2_126_3477_n2849,
         DP_OP_424J2_126_3477_n2848, DP_OP_424J2_126_3477_n2847,
         DP_OP_424J2_126_3477_n2846, DP_OP_424J2_126_3477_n2845,
         DP_OP_424J2_126_3477_n2844, DP_OP_424J2_126_3477_n2841,
         DP_OP_424J2_126_3477_n2837, DP_OP_424J2_126_3477_n2835,
         DP_OP_424J2_126_3477_n2834, DP_OP_424J2_126_3477_n2833,
         DP_OP_424J2_126_3477_n2831, DP_OP_424J2_126_3477_n2830,
         DP_OP_424J2_126_3477_n2829, DP_OP_424J2_126_3477_n2828,
         DP_OP_424J2_126_3477_n2827, DP_OP_424J2_126_3477_n2826,
         DP_OP_424J2_126_3477_n2825, DP_OP_424J2_126_3477_n2824,
         DP_OP_424J2_126_3477_n2823, DP_OP_424J2_126_3477_n2822,
         DP_OP_424J2_126_3477_n2821, DP_OP_424J2_126_3477_n2820,
         DP_OP_424J2_126_3477_n2819, DP_OP_424J2_126_3477_n2818,
         DP_OP_424J2_126_3477_n2817, DP_OP_424J2_126_3477_n2816,
         DP_OP_424J2_126_3477_n2815, DP_OP_424J2_126_3477_n2814,
         DP_OP_424J2_126_3477_n2813, DP_OP_424J2_126_3477_n2812,
         DP_OP_424J2_126_3477_n2811, DP_OP_424J2_126_3477_n2810,
         DP_OP_424J2_126_3477_n2809, DP_OP_424J2_126_3477_n2808,
         DP_OP_424J2_126_3477_n2807, DP_OP_424J2_126_3477_n2806,
         DP_OP_424J2_126_3477_n2805, DP_OP_424J2_126_3477_n2804,
         DP_OP_424J2_126_3477_n2803, DP_OP_424J2_126_3477_n2802,
         DP_OP_424J2_126_3477_n2801, DP_OP_424J2_126_3477_n2800,
         DP_OP_424J2_126_3477_n2799, DP_OP_424J2_126_3477_n2797,
         DP_OP_424J2_126_3477_n2795, DP_OP_424J2_126_3477_n2794,
         DP_OP_424J2_126_3477_n2793, DP_OP_424J2_126_3477_n2791,
         DP_OP_424J2_126_3477_n2790, DP_OP_424J2_126_3477_n2789,
         DP_OP_424J2_126_3477_n2787, DP_OP_424J2_126_3477_n2786,
         DP_OP_424J2_126_3477_n2785, DP_OP_424J2_126_3477_n2784,
         DP_OP_424J2_126_3477_n2783, DP_OP_424J2_126_3477_n2782,
         DP_OP_424J2_126_3477_n2781, DP_OP_424J2_126_3477_n2780,
         DP_OP_424J2_126_3477_n2779, DP_OP_424J2_126_3477_n2778,
         DP_OP_424J2_126_3477_n2777, DP_OP_424J2_126_3477_n2776,
         DP_OP_424J2_126_3477_n2775, DP_OP_424J2_126_3477_n2774,
         DP_OP_424J2_126_3477_n2773, DP_OP_424J2_126_3477_n2772,
         DP_OP_424J2_126_3477_n2771, DP_OP_424J2_126_3477_n2770,
         DP_OP_424J2_126_3477_n2769, DP_OP_424J2_126_3477_n2768,
         DP_OP_424J2_126_3477_n2767, DP_OP_424J2_126_3477_n2766,
         DP_OP_424J2_126_3477_n2765, DP_OP_424J2_126_3477_n2764,
         DP_OP_424J2_126_3477_n2763, DP_OP_424J2_126_3477_n2762,
         DP_OP_424J2_126_3477_n2761, DP_OP_424J2_126_3477_n2760,
         DP_OP_424J2_126_3477_n2759, DP_OP_424J2_126_3477_n2758,
         DP_OP_424J2_126_3477_n2757, DP_OP_424J2_126_3477_n2756,
         DP_OP_424J2_126_3477_n2755, DP_OP_424J2_126_3477_n2753,
         DP_OP_424J2_126_3477_n2751, DP_OP_424J2_126_3477_n2750,
         DP_OP_424J2_126_3477_n2749, DP_OP_424J2_126_3477_n2747,
         DP_OP_424J2_126_3477_n2745, DP_OP_424J2_126_3477_n2743,
         DP_OP_424J2_126_3477_n2742, DP_OP_424J2_126_3477_n2741,
         DP_OP_424J2_126_3477_n2740, DP_OP_424J2_126_3477_n2739,
         DP_OP_424J2_126_3477_n2738, DP_OP_424J2_126_3477_n2737,
         DP_OP_424J2_126_3477_n2736, DP_OP_424J2_126_3477_n2735,
         DP_OP_424J2_126_3477_n2734, DP_OP_424J2_126_3477_n2733,
         DP_OP_424J2_126_3477_n2732, DP_OP_424J2_126_3477_n2731,
         DP_OP_424J2_126_3477_n2730, DP_OP_424J2_126_3477_n2729,
         DP_OP_424J2_126_3477_n2728, DP_OP_424J2_126_3477_n2727,
         DP_OP_424J2_126_3477_n2726, DP_OP_424J2_126_3477_n2725,
         DP_OP_424J2_126_3477_n2724, DP_OP_424J2_126_3477_n2723,
         DP_OP_424J2_126_3477_n2722, DP_OP_424J2_126_3477_n2721,
         DP_OP_424J2_126_3477_n2720, DP_OP_424J2_126_3477_n2719,
         DP_OP_424J2_126_3477_n2718, DP_OP_424J2_126_3477_n2717,
         DP_OP_424J2_126_3477_n2716, DP_OP_424J2_126_3477_n2715,
         DP_OP_424J2_126_3477_n2714, DP_OP_424J2_126_3477_n2713,
         DP_OP_424J2_126_3477_n2712, DP_OP_424J2_126_3477_n2711,
         DP_OP_424J2_126_3477_n2705, DP_OP_424J2_126_3477_n2703,
         DP_OP_424J2_126_3477_n2700, DP_OP_424J2_126_3477_n2699,
         DP_OP_424J2_126_3477_n2698, DP_OP_424J2_126_3477_n2697,
         DP_OP_424J2_126_3477_n2696, DP_OP_424J2_126_3477_n2695,
         DP_OP_424J2_126_3477_n2694, DP_OP_424J2_126_3477_n2693,
         DP_OP_424J2_126_3477_n2692, DP_OP_424J2_126_3477_n2691,
         DP_OP_424J2_126_3477_n2690, DP_OP_424J2_126_3477_n2689,
         DP_OP_424J2_126_3477_n2688, DP_OP_424J2_126_3477_n2687,
         DP_OP_424J2_126_3477_n2686, DP_OP_424J2_126_3477_n2685,
         DP_OP_424J2_126_3477_n2684, DP_OP_424J2_126_3477_n2683,
         DP_OP_424J2_126_3477_n2682, DP_OP_424J2_126_3477_n2681,
         DP_OP_424J2_126_3477_n2680, DP_OP_424J2_126_3477_n2679,
         DP_OP_424J2_126_3477_n2678, DP_OP_424J2_126_3477_n2677,
         DP_OP_424J2_126_3477_n2676, DP_OP_424J2_126_3477_n2675,
         DP_OP_424J2_126_3477_n2674, DP_OP_424J2_126_3477_n2673,
         DP_OP_424J2_126_3477_n2672, DP_OP_424J2_126_3477_n2671,
         DP_OP_424J2_126_3477_n2670, DP_OP_424J2_126_3477_n2669,
         DP_OP_424J2_126_3477_n2668, DP_OP_424J2_126_3477_n2666,
         DP_OP_424J2_126_3477_n2665, DP_OP_424J2_126_3477_n2663,
         DP_OP_424J2_126_3477_n2658, DP_OP_424J2_126_3477_n2655,
         DP_OP_424J2_126_3477_n2654, DP_OP_424J2_126_3477_n2653,
         DP_OP_424J2_126_3477_n2652, DP_OP_424J2_126_3477_n2651,
         DP_OP_424J2_126_3477_n2650, DP_OP_424J2_126_3477_n2649,
         DP_OP_424J2_126_3477_n2648, DP_OP_424J2_126_3477_n2647,
         DP_OP_424J2_126_3477_n2646, DP_OP_424J2_126_3477_n2645,
         DP_OP_424J2_126_3477_n2644, DP_OP_424J2_126_3477_n2643,
         DP_OP_424J2_126_3477_n2642, DP_OP_424J2_126_3477_n2641,
         DP_OP_424J2_126_3477_n2640, DP_OP_424J2_126_3477_n2639,
         DP_OP_424J2_126_3477_n2638, DP_OP_424J2_126_3477_n2637,
         DP_OP_424J2_126_3477_n2636, DP_OP_424J2_126_3477_n2635,
         DP_OP_424J2_126_3477_n2634, DP_OP_424J2_126_3477_n2633,
         DP_OP_424J2_126_3477_n2632, DP_OP_424J2_126_3477_n2631,
         DP_OP_424J2_126_3477_n2630, DP_OP_424J2_126_3477_n2629,
         DP_OP_424J2_126_3477_n2628, DP_OP_424J2_126_3477_n2627,
         DP_OP_424J2_126_3477_n2626, DP_OP_424J2_126_3477_n2625,
         DP_OP_424J2_126_3477_n2624, DP_OP_424J2_126_3477_n2623,
         DP_OP_424J2_126_3477_n2622, DP_OP_424J2_126_3477_n2620,
         DP_OP_424J2_126_3477_n2618, DP_OP_424J2_126_3477_n2616,
         DP_OP_424J2_126_3477_n2613, DP_OP_424J2_126_3477_n2612,
         DP_OP_424J2_126_3477_n2611, DP_OP_424J2_126_3477_n2610,
         DP_OP_424J2_126_3477_n2609, DP_OP_424J2_126_3477_n2608,
         DP_OP_424J2_126_3477_n2607, DP_OP_424J2_126_3477_n2606,
         DP_OP_424J2_126_3477_n2605, DP_OP_424J2_126_3477_n2604,
         DP_OP_424J2_126_3477_n2603, DP_OP_424J2_126_3477_n2602,
         DP_OP_424J2_126_3477_n2601, DP_OP_424J2_126_3477_n2600,
         DP_OP_424J2_126_3477_n2599, DP_OP_424J2_126_3477_n2598,
         DP_OP_424J2_126_3477_n2597, DP_OP_424J2_126_3477_n2596,
         DP_OP_424J2_126_3477_n2595, DP_OP_424J2_126_3477_n2594,
         DP_OP_424J2_126_3477_n2593, DP_OP_424J2_126_3477_n2592,
         DP_OP_424J2_126_3477_n2591, DP_OP_424J2_126_3477_n2590,
         DP_OP_424J2_126_3477_n2589, DP_OP_424J2_126_3477_n2588,
         DP_OP_424J2_126_3477_n2587, DP_OP_424J2_126_3477_n2586,
         DP_OP_424J2_126_3477_n2585, DP_OP_424J2_126_3477_n2584,
         DP_OP_424J2_126_3477_n2583, DP_OP_424J2_126_3477_n2582,
         DP_OP_424J2_126_3477_n2581, DP_OP_424J2_126_3477_n2580,
         DP_OP_424J2_126_3477_n2578, DP_OP_424J2_126_3477_n2572,
         DP_OP_424J2_126_3477_n2569, DP_OP_424J2_126_3477_n2567,
         DP_OP_424J2_126_3477_n2566, DP_OP_424J2_126_3477_n2565,
         DP_OP_424J2_126_3477_n2564, DP_OP_424J2_126_3477_n2563,
         DP_OP_424J2_126_3477_n2562, DP_OP_424J2_126_3477_n2561,
         DP_OP_424J2_126_3477_n2560, DP_OP_424J2_126_3477_n2559,
         DP_OP_424J2_126_3477_n2558, DP_OP_424J2_126_3477_n2557,
         DP_OP_424J2_126_3477_n2556, DP_OP_424J2_126_3477_n2555,
         DP_OP_424J2_126_3477_n2554, DP_OP_424J2_126_3477_n2553,
         DP_OP_424J2_126_3477_n2552, DP_OP_424J2_126_3477_n2551,
         DP_OP_424J2_126_3477_n2550, DP_OP_424J2_126_3477_n2549,
         DP_OP_424J2_126_3477_n2548, DP_OP_424J2_126_3477_n2547,
         DP_OP_424J2_126_3477_n2546, DP_OP_424J2_126_3477_n2545,
         DP_OP_424J2_126_3477_n2544, DP_OP_424J2_126_3477_n2543,
         DP_OP_424J2_126_3477_n2542, DP_OP_424J2_126_3477_n2541,
         DP_OP_424J2_126_3477_n2540, DP_OP_424J2_126_3477_n2539,
         DP_OP_424J2_126_3477_n2538, DP_OP_424J2_126_3477_n2537,
         DP_OP_424J2_126_3477_n2536, DP_OP_424J2_126_3477_n2533,
         DP_OP_424J2_126_3477_n2532, DP_OP_424J2_126_3477_n2530,
         DP_OP_424J2_126_3477_n2528, DP_OP_424J2_126_3477_n2526,
         DP_OP_424J2_126_3477_n2523, DP_OP_424J2_126_3477_n2522,
         DP_OP_424J2_126_3477_n2521, DP_OP_424J2_126_3477_n2520,
         DP_OP_424J2_126_3477_n2519, DP_OP_424J2_126_3477_n2518,
         DP_OP_424J2_126_3477_n2517, DP_OP_424J2_126_3477_n2516,
         DP_OP_424J2_126_3477_n2515, DP_OP_424J2_126_3477_n2514,
         DP_OP_424J2_126_3477_n2513, DP_OP_424J2_126_3477_n2512,
         DP_OP_424J2_126_3477_n2511, DP_OP_424J2_126_3477_n2510,
         DP_OP_424J2_126_3477_n2509, DP_OP_424J2_126_3477_n2508,
         DP_OP_424J2_126_3477_n2507, DP_OP_424J2_126_3477_n2506,
         DP_OP_424J2_126_3477_n2505, DP_OP_424J2_126_3477_n2504,
         DP_OP_424J2_126_3477_n2503, DP_OP_424J2_126_3477_n2502,
         DP_OP_424J2_126_3477_n2501, DP_OP_424J2_126_3477_n2500,
         DP_OP_424J2_126_3477_n2499, DP_OP_424J2_126_3477_n2498,
         DP_OP_424J2_126_3477_n2497, DP_OP_424J2_126_3477_n2496,
         DP_OP_424J2_126_3477_n2495, DP_OP_424J2_126_3477_n2494,
         DP_OP_424J2_126_3477_n2493, DP_OP_424J2_126_3477_n2492,
         DP_OP_424J2_126_3477_n2489, DP_OP_424J2_126_3477_n2488,
         DP_OP_424J2_126_3477_n2484, DP_OP_424J2_126_3477_n2482,
         DP_OP_424J2_126_3477_n2481, DP_OP_424J2_126_3477_n2479,
         DP_OP_424J2_126_3477_n2478, DP_OP_424J2_126_3477_n2477,
         DP_OP_424J2_126_3477_n2476, DP_OP_424J2_126_3477_n2475,
         DP_OP_424J2_126_3477_n2474, DP_OP_424J2_126_3477_n2473,
         DP_OP_424J2_126_3477_n2472, DP_OP_424J2_126_3477_n2471,
         DP_OP_424J2_126_3477_n2470, DP_OP_424J2_126_3477_n2469,
         DP_OP_424J2_126_3477_n2468, DP_OP_424J2_126_3477_n2467,
         DP_OP_424J2_126_3477_n2466, DP_OP_424J2_126_3477_n2465,
         DP_OP_424J2_126_3477_n2464, DP_OP_424J2_126_3477_n2463,
         DP_OP_424J2_126_3477_n2462, DP_OP_424J2_126_3477_n2461,
         DP_OP_424J2_126_3477_n2460, DP_OP_424J2_126_3477_n2459,
         DP_OP_424J2_126_3477_n2458, DP_OP_424J2_126_3477_n2457,
         DP_OP_424J2_126_3477_n2456, DP_OP_424J2_126_3477_n2455,
         DP_OP_424J2_126_3477_n2454, DP_OP_424J2_126_3477_n2453,
         DP_OP_424J2_126_3477_n2452, DP_OP_424J2_126_3477_n2451,
         DP_OP_424J2_126_3477_n2450, DP_OP_424J2_126_3477_n2449,
         DP_OP_424J2_126_3477_n2448, DP_OP_424J2_126_3477_n2447,
         DP_OP_424J2_126_3477_n2446, DP_OP_424J2_126_3477_n2445,
         DP_OP_424J2_126_3477_n2444, DP_OP_424J2_126_3477_n2442,
         DP_OP_424J2_126_3477_n2439, DP_OP_424J2_126_3477_n2435,
         DP_OP_424J2_126_3477_n2434, DP_OP_424J2_126_3477_n2433,
         DP_OP_424J2_126_3477_n2432, DP_OP_424J2_126_3477_n2431,
         DP_OP_424J2_126_3477_n2430, DP_OP_424J2_126_3477_n2429,
         DP_OP_424J2_126_3477_n2428, DP_OP_424J2_126_3477_n2427,
         DP_OP_424J2_126_3477_n2426, DP_OP_424J2_126_3477_n2425,
         DP_OP_424J2_126_3477_n2424, DP_OP_424J2_126_3477_n2423,
         DP_OP_424J2_126_3477_n2422, DP_OP_424J2_126_3477_n2421,
         DP_OP_424J2_126_3477_n2420, DP_OP_424J2_126_3477_n2419,
         DP_OP_424J2_126_3477_n2418, DP_OP_424J2_126_3477_n2417,
         DP_OP_424J2_126_3477_n2416, DP_OP_424J2_126_3477_n2415,
         DP_OP_424J2_126_3477_n2414, DP_OP_424J2_126_3477_n2413,
         DP_OP_424J2_126_3477_n2412, DP_OP_424J2_126_3477_n2411,
         DP_OP_424J2_126_3477_n2410, DP_OP_424J2_126_3477_n2409,
         DP_OP_424J2_126_3477_n2408, DP_OP_424J2_126_3477_n2407,
         DP_OP_424J2_126_3477_n2406, DP_OP_424J2_126_3477_n2405,
         DP_OP_424J2_126_3477_n2404, DP_OP_424J2_126_3477_n2402,
         DP_OP_424J2_126_3477_n2401, DP_OP_424J2_126_3477_n2397,
         DP_OP_424J2_126_3477_n2391, DP_OP_424J2_126_3477_n2390,
         DP_OP_424J2_126_3477_n2389, DP_OP_424J2_126_3477_n2388,
         DP_OP_424J2_126_3477_n2387, DP_OP_424J2_126_3477_n2386,
         DP_OP_424J2_126_3477_n2385, DP_OP_424J2_126_3477_n2384,
         DP_OP_424J2_126_3477_n2383, DP_OP_424J2_126_3477_n2382,
         DP_OP_424J2_126_3477_n2381, DP_OP_424J2_126_3477_n2380,
         DP_OP_424J2_126_3477_n2379, DP_OP_424J2_126_3477_n2378,
         DP_OP_424J2_126_3477_n2377, DP_OP_424J2_126_3477_n2376,
         DP_OP_424J2_126_3477_n2375, DP_OP_424J2_126_3477_n2374,
         DP_OP_424J2_126_3477_n2373, DP_OP_424J2_126_3477_n2372,
         DP_OP_424J2_126_3477_n2371, DP_OP_424J2_126_3477_n2370,
         DP_OP_424J2_126_3477_n2369, DP_OP_424J2_126_3477_n2368,
         DP_OP_424J2_126_3477_n2367, DP_OP_424J2_126_3477_n2366,
         DP_OP_424J2_126_3477_n2365, DP_OP_424J2_126_3477_n2364,
         DP_OP_424J2_126_3477_n2363, DP_OP_424J2_126_3477_n2362,
         DP_OP_424J2_126_3477_n2361, DP_OP_424J2_126_3477_n2360,
         DP_OP_424J2_126_3477_n2358, DP_OP_424J2_126_3477_n2357,
         DP_OP_424J2_126_3477_n2354, DP_OP_424J2_126_3477_n2353,
         DP_OP_424J2_126_3477_n2351, DP_OP_424J2_126_3477_n2347,
         DP_OP_424J2_126_3477_n2346, DP_OP_424J2_126_3477_n2345,
         DP_OP_424J2_126_3477_n2344, DP_OP_424J2_126_3477_n2343,
         DP_OP_424J2_126_3477_n2342, DP_OP_424J2_126_3477_n2341,
         DP_OP_424J2_126_3477_n2340, DP_OP_424J2_126_3477_n2339,
         DP_OP_424J2_126_3477_n2338, DP_OP_424J2_126_3477_n2337,
         DP_OP_424J2_126_3477_n2336, DP_OP_424J2_126_3477_n2335,
         DP_OP_424J2_126_3477_n2334, DP_OP_424J2_126_3477_n2333,
         DP_OP_424J2_126_3477_n2332, DP_OP_424J2_126_3477_n2331,
         DP_OP_424J2_126_3477_n2330, DP_OP_424J2_126_3477_n2329,
         DP_OP_424J2_126_3477_n2328, DP_OP_424J2_126_3477_n2327,
         DP_OP_424J2_126_3477_n2326, DP_OP_424J2_126_3477_n2325,
         DP_OP_424J2_126_3477_n2324, DP_OP_424J2_126_3477_n2323,
         DP_OP_424J2_126_3477_n2322, DP_OP_424J2_126_3477_n2321,
         DP_OP_424J2_126_3477_n2320, DP_OP_424J2_126_3477_n2319,
         DP_OP_424J2_126_3477_n2318, DP_OP_424J2_126_3477_n2317,
         DP_OP_424J2_126_3477_n2316, DP_OP_424J2_126_3477_n2315,
         DP_OP_424J2_126_3477_n2314, DP_OP_424J2_126_3477_n2310,
         DP_OP_424J2_126_3477_n2308, DP_OP_424J2_126_3477_n2304,
         DP_OP_424J2_126_3477_n2303, DP_OP_424J2_126_3477_n2302,
         DP_OP_424J2_126_3477_n2301, DP_OP_424J2_126_3477_n2300,
         DP_OP_424J2_126_3477_n2299, DP_OP_424J2_126_3477_n2298,
         DP_OP_424J2_126_3477_n2297, DP_OP_424J2_126_3477_n2296,
         DP_OP_424J2_126_3477_n2295, DP_OP_424J2_126_3477_n2294,
         DP_OP_424J2_126_3477_n2293, DP_OP_424J2_126_3477_n2292,
         DP_OP_424J2_126_3477_n2291, DP_OP_424J2_126_3477_n2290,
         DP_OP_424J2_126_3477_n2289, DP_OP_424J2_126_3477_n2288,
         DP_OP_424J2_126_3477_n2287, DP_OP_424J2_126_3477_n2286,
         DP_OP_424J2_126_3477_n2285, DP_OP_424J2_126_3477_n2284,
         DP_OP_424J2_126_3477_n2283, DP_OP_424J2_126_3477_n2282,
         DP_OP_424J2_126_3477_n2281, DP_OP_424J2_126_3477_n2280,
         DP_OP_424J2_126_3477_n2279, DP_OP_424J2_126_3477_n2278,
         DP_OP_424J2_126_3477_n2277, DP_OP_424J2_126_3477_n2276,
         DP_OP_424J2_126_3477_n2275, DP_OP_424J2_126_3477_n2274,
         DP_OP_424J2_126_3477_n2273, DP_OP_424J2_126_3477_n2272,
         DP_OP_424J2_126_3477_n2271, DP_OP_424J2_126_3477_n2270,
         DP_OP_424J2_126_3477_n2269, DP_OP_424J2_126_3477_n2265,
         DP_OP_424J2_126_3477_n2264, DP_OP_424J2_126_3477_n2261,
         DP_OP_424J2_126_3477_n2260, DP_OP_424J2_126_3477_n2259,
         DP_OP_424J2_126_3477_n2258, DP_OP_424J2_126_3477_n2257,
         DP_OP_424J2_126_3477_n2256, DP_OP_424J2_126_3477_n2255,
         DP_OP_424J2_126_3477_n2254, DP_OP_424J2_126_3477_n2253,
         DP_OP_424J2_126_3477_n2252, DP_OP_424J2_126_3477_n2251,
         DP_OP_424J2_126_3477_n2250, DP_OP_424J2_126_3477_n2249,
         DP_OP_424J2_126_3477_n2248, DP_OP_424J2_126_3477_n2247,
         DP_OP_424J2_126_3477_n2246, DP_OP_424J2_126_3477_n2245,
         DP_OP_424J2_126_3477_n2244, DP_OP_424J2_126_3477_n2243,
         DP_OP_424J2_126_3477_n2242, DP_OP_424J2_126_3477_n2241,
         DP_OP_424J2_126_3477_n2240, DP_OP_424J2_126_3477_n2239,
         DP_OP_424J2_126_3477_n2238, DP_OP_424J2_126_3477_n2237,
         DP_OP_424J2_126_3477_n2236, DP_OP_424J2_126_3477_n2235,
         DP_OP_424J2_126_3477_n2234, DP_OP_424J2_126_3477_n2233,
         DP_OP_424J2_126_3477_n2232, DP_OP_424J2_126_3477_n2231,
         DP_OP_424J2_126_3477_n2230, DP_OP_424J2_126_3477_n2229,
         DP_OP_424J2_126_3477_n2228, DP_OP_424J2_126_3477_n2227,
         DP_OP_424J2_126_3477_n2226, DP_OP_424J2_126_3477_n2225,
         DP_OP_424J2_126_3477_n2220, DP_OP_424J2_126_3477_n2219,
         DP_OP_424J2_126_3477_n2218, DP_OP_424J2_126_3477_n2217,
         DP_OP_424J2_126_3477_n2215, DP_OP_424J2_126_3477_n2214,
         DP_OP_424J2_126_3477_n2213, DP_OP_424J2_126_3477_n2212,
         DP_OP_424J2_126_3477_n2211, DP_OP_424J2_126_3477_n2210,
         DP_OP_424J2_126_3477_n2209, DP_OP_424J2_126_3477_n2208,
         DP_OP_424J2_126_3477_n2207, DP_OP_424J2_126_3477_n2206,
         DP_OP_424J2_126_3477_n2205, DP_OP_424J2_126_3477_n2204,
         DP_OP_424J2_126_3477_n2203, DP_OP_424J2_126_3477_n2202,
         DP_OP_424J2_126_3477_n2201, DP_OP_424J2_126_3477_n2200,
         DP_OP_424J2_126_3477_n2199, DP_OP_424J2_126_3477_n2198,
         DP_OP_424J2_126_3477_n2197, DP_OP_424J2_126_3477_n2196,
         DP_OP_424J2_126_3477_n2195, DP_OP_424J2_126_3477_n2194,
         DP_OP_424J2_126_3477_n2193, DP_OP_424J2_126_3477_n2192,
         DP_OP_424J2_126_3477_n2191, DP_OP_424J2_126_3477_n2190,
         DP_OP_424J2_126_3477_n2189, DP_OP_424J2_126_3477_n2188,
         DP_OP_424J2_126_3477_n2187, DP_OP_424J2_126_3477_n2186,
         DP_OP_424J2_126_3477_n2185, DP_OP_424J2_126_3477_n2184,
         DP_OP_424J2_126_3477_n2183, DP_OP_424J2_126_3477_n2182,
         DP_OP_424J2_126_3477_n2179, DP_OP_424J2_126_3477_n2178,
         DP_OP_424J2_126_3477_n2177, DP_OP_424J2_126_3477_n2172,
         DP_OP_424J2_126_3477_n2171, DP_OP_424J2_126_3477_n2170,
         DP_OP_424J2_126_3477_n2169, DP_OP_424J2_126_3477_n2168,
         DP_OP_424J2_126_3477_n2167, DP_OP_424J2_126_3477_n2166,
         DP_OP_424J2_126_3477_n2165, DP_OP_424J2_126_3477_n2164,
         DP_OP_424J2_126_3477_n2163, DP_OP_424J2_126_3477_n2162,
         DP_OP_424J2_126_3477_n2161, DP_OP_424J2_126_3477_n2160,
         DP_OP_424J2_126_3477_n2159, DP_OP_424J2_126_3477_n2158,
         DP_OP_424J2_126_3477_n2157, DP_OP_424J2_126_3477_n2156,
         DP_OP_424J2_126_3477_n2155, DP_OP_424J2_126_3477_n2154,
         DP_OP_424J2_126_3477_n2153, DP_OP_424J2_126_3477_n2152,
         DP_OP_424J2_126_3477_n2151, DP_OP_424J2_126_3477_n2150,
         DP_OP_424J2_126_3477_n2149, DP_OP_424J2_126_3477_n2148,
         DP_OP_424J2_126_3477_n2147, DP_OP_424J2_126_3477_n2146,
         DP_OP_424J2_126_3477_n2145, DP_OP_424J2_126_3477_n2144,
         DP_OP_424J2_126_3477_n2143, DP_OP_424J2_126_3477_n2142,
         DP_OP_424J2_126_3477_n2141, DP_OP_424J2_126_3477_n2140,
         DP_OP_424J2_126_3477_n2137, DP_OP_424J2_126_3477_n2133,
         DP_OP_424J2_126_3477_n2128, DP_OP_424J2_126_3477_n2127,
         DP_OP_424J2_126_3477_n2126, DP_OP_424J2_126_3477_n2125,
         DP_OP_424J2_126_3477_n2124, DP_OP_424J2_126_3477_n2123,
         DP_OP_424J2_126_3477_n2122, DP_OP_424J2_126_3477_n2121,
         DP_OP_424J2_126_3477_n2120, DP_OP_424J2_126_3477_n2119,
         DP_OP_424J2_126_3477_n2118, DP_OP_424J2_126_3477_n2117,
         DP_OP_424J2_126_3477_n2116, DP_OP_424J2_126_3477_n2115,
         DP_OP_424J2_126_3477_n2114, DP_OP_424J2_126_3477_n2113,
         DP_OP_424J2_126_3477_n2112, DP_OP_424J2_126_3477_n2111,
         DP_OP_424J2_126_3477_n2110, DP_OP_424J2_126_3477_n2109,
         DP_OP_424J2_126_3477_n2108, DP_OP_424J2_126_3477_n2107,
         DP_OP_424J2_126_3477_n2106, DP_OP_424J2_126_3477_n2105,
         DP_OP_424J2_126_3477_n2104, DP_OP_424J2_126_3477_n2103,
         DP_OP_424J2_126_3477_n2102, DP_OP_424J2_126_3477_n2101,
         DP_OP_424J2_126_3477_n2100, DP_OP_424J2_126_3477_n2099,
         DP_OP_424J2_126_3477_n2098, DP_OP_424J2_126_3477_n2097,
         DP_OP_424J2_126_3477_n2096, DP_OP_424J2_126_3477_n2095,
         DP_OP_424J2_126_3477_n2094, DP_OP_424J2_126_3477_n2090,
         DP_OP_424J2_126_3477_n2088, DP_OP_424J2_126_3477_n2087,
         DP_OP_424J2_126_3477_n2084, DP_OP_424J2_126_3477_n2083,
         DP_OP_424J2_126_3477_n2082, DP_OP_424J2_126_3477_n2081,
         DP_OP_424J2_126_3477_n2080, DP_OP_424J2_126_3477_n2079,
         DP_OP_424J2_126_3477_n2078, DP_OP_424J2_126_3477_n2077,
         DP_OP_424J2_126_3477_n2076, DP_OP_424J2_126_3477_n2075,
         DP_OP_424J2_126_3477_n2074, DP_OP_424J2_126_3477_n2073,
         DP_OP_424J2_126_3477_n2072, DP_OP_424J2_126_3477_n2071,
         DP_OP_424J2_126_3477_n2070, DP_OP_424J2_126_3477_n2069,
         DP_OP_424J2_126_3477_n2068, DP_OP_424J2_126_3477_n2067,
         DP_OP_424J2_126_3477_n2066, DP_OP_424J2_126_3477_n2065,
         DP_OP_424J2_126_3477_n2064, DP_OP_424J2_126_3477_n2063,
         DP_OP_424J2_126_3477_n2062, DP_OP_424J2_126_3477_n2061,
         DP_OP_424J2_126_3477_n2060, DP_OP_424J2_126_3477_n2059,
         DP_OP_424J2_126_3477_n2058, DP_OP_424J2_126_3477_n2057,
         DP_OP_424J2_126_3477_n2056, DP_OP_424J2_126_3477_n2055,
         DP_OP_424J2_126_3477_n2054, DP_OP_424J2_126_3477_n2053,
         DP_OP_424J2_126_3477_n2052, DP_OP_424J2_126_3477_n2051,
         DP_OP_424J2_126_3477_n2049, DP_OP_424J2_126_3477_n2047,
         DP_OP_424J2_126_3477_n2044, DP_OP_424J2_126_3477_n2039,
         DP_OP_424J2_126_3477_n2038, DP_OP_424J2_126_3477_n2037,
         DP_OP_424J2_126_3477_n2036, DP_OP_424J2_126_3477_n2035,
         DP_OP_424J2_126_3477_n2034, DP_OP_424J2_126_3477_n2033,
         DP_OP_424J2_126_3477_n2032, DP_OP_424J2_126_3477_n2031,
         DP_OP_424J2_126_3477_n2030, DP_OP_424J2_126_3477_n2029,
         DP_OP_424J2_126_3477_n2028, DP_OP_424J2_126_3477_n2027,
         DP_OP_424J2_126_3477_n2026, DP_OP_424J2_126_3477_n2025,
         DP_OP_424J2_126_3477_n2024, DP_OP_424J2_126_3477_n2023,
         DP_OP_424J2_126_3477_n2022, DP_OP_424J2_126_3477_n2021,
         DP_OP_424J2_126_3477_n2020, DP_OP_424J2_126_3477_n2019,
         DP_OP_424J2_126_3477_n2018, DP_OP_424J2_126_3477_n2017,
         DP_OP_424J2_126_3477_n2016, DP_OP_424J2_126_3477_n2015,
         DP_OP_424J2_126_3477_n2014, DP_OP_424J2_126_3477_n2013,
         DP_OP_424J2_126_3477_n2012, DP_OP_424J2_126_3477_n2011,
         DP_OP_424J2_126_3477_n2010, DP_OP_424J2_126_3477_n2009,
         DP_OP_424J2_126_3477_n2008, DP_OP_424J2_126_3477_n2001,
         DP_OP_424J2_126_3477_n1995, DP_OP_424J2_126_3477_n1994,
         DP_OP_424J2_126_3477_n1993, DP_OP_424J2_126_3477_n1992,
         DP_OP_424J2_126_3477_n1991, DP_OP_424J2_126_3477_n1990,
         DP_OP_424J2_126_3477_n1989, DP_OP_424J2_126_3477_n1988,
         DP_OP_424J2_126_3477_n1987, DP_OP_424J2_126_3477_n1986,
         DP_OP_424J2_126_3477_n1985, DP_OP_424J2_126_3477_n1984,
         DP_OP_424J2_126_3477_n1983, DP_OP_424J2_126_3477_n1982,
         DP_OP_424J2_126_3477_n1981, DP_OP_424J2_126_3477_n1980,
         DP_OP_424J2_126_3477_n1979, DP_OP_424J2_126_3477_n1978,
         DP_OP_424J2_126_3477_n1977, DP_OP_424J2_126_3477_n1976,
         DP_OP_424J2_126_3477_n1975, DP_OP_424J2_126_3477_n1974,
         DP_OP_424J2_126_3477_n1973, DP_OP_424J2_126_3477_n1972,
         DP_OP_424J2_126_3477_n1971, DP_OP_424J2_126_3477_n1970,
         DP_OP_424J2_126_3477_n1969, DP_OP_424J2_126_3477_n1968,
         DP_OP_424J2_126_3477_n1967, DP_OP_424J2_126_3477_n1966,
         DP_OP_424J2_126_3477_n1965, DP_OP_424J2_126_3477_n1964,
         DP_OP_424J2_126_3477_n1962, DP_OP_424J2_126_3477_n1961,
         DP_OP_424J2_126_3477_n1958, DP_OP_424J2_126_3477_n1957,
         DP_OP_424J2_126_3477_n1956, DP_OP_424J2_126_3477_n1954,
         DP_OP_424J2_126_3477_n1951, DP_OP_424J2_126_3477_n1950,
         DP_OP_424J2_126_3477_n1949, DP_OP_424J2_126_3477_n1948,
         DP_OP_424J2_126_3477_n1947, DP_OP_424J2_126_3477_n1946,
         DP_OP_424J2_126_3477_n1945, DP_OP_424J2_126_3477_n1944,
         DP_OP_424J2_126_3477_n1943, DP_OP_424J2_126_3477_n1942,
         DP_OP_424J2_126_3477_n1941, DP_OP_424J2_126_3477_n1940,
         DP_OP_424J2_126_3477_n1939, DP_OP_424J2_126_3477_n1938,
         DP_OP_424J2_126_3477_n1937, DP_OP_424J2_126_3477_n1936,
         DP_OP_424J2_126_3477_n1935, DP_OP_424J2_126_3477_n1934,
         DP_OP_424J2_126_3477_n1933, DP_OP_424J2_126_3477_n1932,
         DP_OP_424J2_126_3477_n1931, DP_OP_424J2_126_3477_n1930,
         DP_OP_424J2_126_3477_n1929, DP_OP_424J2_126_3477_n1928,
         DP_OP_424J2_126_3477_n1927, DP_OP_424J2_126_3477_n1926,
         DP_OP_424J2_126_3477_n1925, DP_OP_424J2_126_3477_n1924,
         DP_OP_424J2_126_3477_n1923, DP_OP_424J2_126_3477_n1922,
         DP_OP_424J2_126_3477_n1921, DP_OP_424J2_126_3477_n1920,
         DP_OP_424J2_126_3477_n1886, DP_OP_424J2_126_3477_n1885,
         DP_OP_424J2_126_3477_n1884, DP_OP_424J2_126_3477_n1883,
         DP_OP_424J2_126_3477_n1882, DP_OP_424J2_126_3477_n1881,
         DP_OP_424J2_126_3477_n1880, DP_OP_424J2_126_3477_n1879,
         DP_OP_424J2_126_3477_n1878, DP_OP_424J2_126_3477_n1877,
         DP_OP_424J2_126_3477_n1876, DP_OP_424J2_126_3477_n1875,
         DP_OP_424J2_126_3477_n1874, DP_OP_424J2_126_3477_n1873,
         DP_OP_424J2_126_3477_n1871, DP_OP_424J2_126_3477_n1870,
         DP_OP_424J2_126_3477_n1869, DP_OP_424J2_126_3477_n1868,
         DP_OP_424J2_126_3477_n1867, DP_OP_424J2_126_3477_n1866,
         DP_OP_424J2_126_3477_n1865, DP_OP_424J2_126_3477_n1864,
         DP_OP_424J2_126_3477_n1863, DP_OP_424J2_126_3477_n1862,
         DP_OP_424J2_126_3477_n1861, DP_OP_424J2_126_3477_n1860,
         DP_OP_424J2_126_3477_n1859, DP_OP_424J2_126_3477_n1858,
         DP_OP_424J2_126_3477_n1857, DP_OP_424J2_126_3477_n1856,
         DP_OP_424J2_126_3477_n1855, DP_OP_424J2_126_3477_n1854,
         DP_OP_424J2_126_3477_n1853, DP_OP_424J2_126_3477_n1852,
         DP_OP_424J2_126_3477_n1851, DP_OP_424J2_126_3477_n1850,
         DP_OP_424J2_126_3477_n1849, DP_OP_424J2_126_3477_n1848,
         DP_OP_424J2_126_3477_n1847, DP_OP_424J2_126_3477_n1846,
         DP_OP_424J2_126_3477_n1845, DP_OP_424J2_126_3477_n1844,
         DP_OP_424J2_126_3477_n1843, DP_OP_424J2_126_3477_n1842,
         DP_OP_424J2_126_3477_n1841, DP_OP_424J2_126_3477_n1840,
         DP_OP_424J2_126_3477_n1839, DP_OP_424J2_126_3477_n1838,
         DP_OP_424J2_126_3477_n1837, DP_OP_424J2_126_3477_n1836,
         DP_OP_424J2_126_3477_n1835, DP_OP_424J2_126_3477_n1834,
         DP_OP_424J2_126_3477_n1833, DP_OP_424J2_126_3477_n1832,
         DP_OP_424J2_126_3477_n1831, DP_OP_424J2_126_3477_n1830,
         DP_OP_424J2_126_3477_n1829, DP_OP_424J2_126_3477_n1828,
         DP_OP_424J2_126_3477_n1827, DP_OP_424J2_126_3477_n1826,
         DP_OP_424J2_126_3477_n1825, DP_OP_424J2_126_3477_n1824,
         DP_OP_424J2_126_3477_n1823, DP_OP_424J2_126_3477_n1822,
         DP_OP_424J2_126_3477_n1821, DP_OP_424J2_126_3477_n1820,
         DP_OP_424J2_126_3477_n1819, DP_OP_424J2_126_3477_n1818,
         DP_OP_424J2_126_3477_n1817, DP_OP_424J2_126_3477_n1816,
         DP_OP_424J2_126_3477_n1815, DP_OP_424J2_126_3477_n1814,
         DP_OP_424J2_126_3477_n1813, DP_OP_424J2_126_3477_n1812,
         DP_OP_424J2_126_3477_n1811, DP_OP_424J2_126_3477_n1810,
         DP_OP_424J2_126_3477_n1809, DP_OP_424J2_126_3477_n1808,
         DP_OP_424J2_126_3477_n1807, DP_OP_424J2_126_3477_n1806,
         DP_OP_424J2_126_3477_n1805, DP_OP_424J2_126_3477_n1804,
         DP_OP_424J2_126_3477_n1803, DP_OP_424J2_126_3477_n1802,
         DP_OP_424J2_126_3477_n1801, DP_OP_424J2_126_3477_n1800,
         DP_OP_424J2_126_3477_n1799, DP_OP_424J2_126_3477_n1798,
         DP_OP_424J2_126_3477_n1797, DP_OP_424J2_126_3477_n1796,
         DP_OP_424J2_126_3477_n1795, DP_OP_424J2_126_3477_n1794,
         DP_OP_424J2_126_3477_n1793, DP_OP_424J2_126_3477_n1792,
         DP_OP_424J2_126_3477_n1791, DP_OP_424J2_126_3477_n1790,
         DP_OP_424J2_126_3477_n1789, DP_OP_424J2_126_3477_n1788,
         DP_OP_424J2_126_3477_n1787, DP_OP_424J2_126_3477_n1786,
         DP_OP_424J2_126_3477_n1785, DP_OP_424J2_126_3477_n1784,
         DP_OP_424J2_126_3477_n1783, DP_OP_424J2_126_3477_n1782,
         DP_OP_424J2_126_3477_n1781, DP_OP_424J2_126_3477_n1780,
         DP_OP_424J2_126_3477_n1779, DP_OP_424J2_126_3477_n1778,
         DP_OP_424J2_126_3477_n1777, DP_OP_424J2_126_3477_n1776,
         DP_OP_424J2_126_3477_n1775, DP_OP_424J2_126_3477_n1774,
         DP_OP_424J2_126_3477_n1773, DP_OP_424J2_126_3477_n1772,
         DP_OP_424J2_126_3477_n1771, DP_OP_424J2_126_3477_n1770,
         DP_OP_424J2_126_3477_n1769, DP_OP_424J2_126_3477_n1768,
         DP_OP_424J2_126_3477_n1767, DP_OP_424J2_126_3477_n1766,
         DP_OP_424J2_126_3477_n1765, DP_OP_424J2_126_3477_n1764,
         DP_OP_424J2_126_3477_n1763, DP_OP_424J2_126_3477_n1762,
         DP_OP_424J2_126_3477_n1761, DP_OP_424J2_126_3477_n1760,
         DP_OP_424J2_126_3477_n1759, DP_OP_424J2_126_3477_n1758,
         DP_OP_424J2_126_3477_n1757, DP_OP_424J2_126_3477_n1756,
         DP_OP_424J2_126_3477_n1755, DP_OP_424J2_126_3477_n1754,
         DP_OP_424J2_126_3477_n1753, DP_OP_424J2_126_3477_n1752,
         DP_OP_424J2_126_3477_n1751, DP_OP_424J2_126_3477_n1750,
         DP_OP_424J2_126_3477_n1749, DP_OP_424J2_126_3477_n1748,
         DP_OP_424J2_126_3477_n1747, DP_OP_424J2_126_3477_n1746,
         DP_OP_424J2_126_3477_n1745, DP_OP_424J2_126_3477_n1744,
         DP_OP_424J2_126_3477_n1743, DP_OP_424J2_126_3477_n1742,
         DP_OP_424J2_126_3477_n1741, DP_OP_424J2_126_3477_n1740,
         DP_OP_424J2_126_3477_n1739, DP_OP_424J2_126_3477_n1738,
         DP_OP_424J2_126_3477_n1737, DP_OP_424J2_126_3477_n1736,
         DP_OP_424J2_126_3477_n1735, DP_OP_424J2_126_3477_n1734,
         DP_OP_424J2_126_3477_n1733, DP_OP_424J2_126_3477_n1732,
         DP_OP_424J2_126_3477_n1731, DP_OP_424J2_126_3477_n1730,
         DP_OP_424J2_126_3477_n1729, DP_OP_424J2_126_3477_n1728,
         DP_OP_424J2_126_3477_n1727, DP_OP_424J2_126_3477_n1726,
         DP_OP_424J2_126_3477_n1725, DP_OP_424J2_126_3477_n1724,
         DP_OP_424J2_126_3477_n1723, DP_OP_424J2_126_3477_n1722,
         DP_OP_424J2_126_3477_n1721, DP_OP_424J2_126_3477_n1720,
         DP_OP_424J2_126_3477_n1719, DP_OP_424J2_126_3477_n1718,
         DP_OP_424J2_126_3477_n1717, DP_OP_424J2_126_3477_n1716,
         DP_OP_424J2_126_3477_n1715, DP_OP_424J2_126_3477_n1714,
         DP_OP_424J2_126_3477_n1713, DP_OP_424J2_126_3477_n1712,
         DP_OP_424J2_126_3477_n1711, DP_OP_424J2_126_3477_n1710,
         DP_OP_424J2_126_3477_n1709, DP_OP_424J2_126_3477_n1708,
         DP_OP_424J2_126_3477_n1707, DP_OP_424J2_126_3477_n1706,
         DP_OP_424J2_126_3477_n1705, DP_OP_424J2_126_3477_n1704,
         DP_OP_424J2_126_3477_n1703, DP_OP_424J2_126_3477_n1702,
         DP_OP_424J2_126_3477_n1701, DP_OP_424J2_126_3477_n1700,
         DP_OP_424J2_126_3477_n1699, DP_OP_424J2_126_3477_n1698,
         DP_OP_424J2_126_3477_n1697, DP_OP_424J2_126_3477_n1696,
         DP_OP_424J2_126_3477_n1695, DP_OP_424J2_126_3477_n1694,
         DP_OP_424J2_126_3477_n1693, DP_OP_424J2_126_3477_n1692,
         DP_OP_424J2_126_3477_n1691, DP_OP_424J2_126_3477_n1690,
         DP_OP_424J2_126_3477_n1689, DP_OP_424J2_126_3477_n1688,
         DP_OP_424J2_126_3477_n1687, DP_OP_424J2_126_3477_n1686,
         DP_OP_424J2_126_3477_n1685, DP_OP_424J2_126_3477_n1684,
         DP_OP_424J2_126_3477_n1683, DP_OP_424J2_126_3477_n1682,
         DP_OP_424J2_126_3477_n1681, DP_OP_424J2_126_3477_n1680,
         DP_OP_424J2_126_3477_n1679, DP_OP_424J2_126_3477_n1678,
         DP_OP_424J2_126_3477_n1677, DP_OP_424J2_126_3477_n1676,
         DP_OP_424J2_126_3477_n1675, DP_OP_424J2_126_3477_n1674,
         DP_OP_424J2_126_3477_n1673, DP_OP_424J2_126_3477_n1672,
         DP_OP_424J2_126_3477_n1671, DP_OP_424J2_126_3477_n1670,
         DP_OP_424J2_126_3477_n1669, DP_OP_424J2_126_3477_n1668,
         DP_OP_424J2_126_3477_n1667, DP_OP_424J2_126_3477_n1666,
         DP_OP_424J2_126_3477_n1665, DP_OP_424J2_126_3477_n1664,
         DP_OP_424J2_126_3477_n1663, DP_OP_424J2_126_3477_n1662,
         DP_OP_424J2_126_3477_n1661, DP_OP_424J2_126_3477_n1660,
         DP_OP_424J2_126_3477_n1659, DP_OP_424J2_126_3477_n1658,
         DP_OP_424J2_126_3477_n1657, DP_OP_424J2_126_3477_n1656,
         DP_OP_424J2_126_3477_n1655, DP_OP_424J2_126_3477_n1654,
         DP_OP_424J2_126_3477_n1653, DP_OP_424J2_126_3477_n1652,
         DP_OP_424J2_126_3477_n1651, DP_OP_424J2_126_3477_n1650,
         DP_OP_424J2_126_3477_n1649, DP_OP_424J2_126_3477_n1648,
         DP_OP_424J2_126_3477_n1647, DP_OP_424J2_126_3477_n1646,
         DP_OP_424J2_126_3477_n1645, DP_OP_424J2_126_3477_n1644,
         DP_OP_424J2_126_3477_n1643, DP_OP_424J2_126_3477_n1642,
         DP_OP_424J2_126_3477_n1641, DP_OP_424J2_126_3477_n1640,
         DP_OP_424J2_126_3477_n1639, DP_OP_424J2_126_3477_n1638,
         DP_OP_424J2_126_3477_n1637, DP_OP_424J2_126_3477_n1636,
         DP_OP_424J2_126_3477_n1635, DP_OP_424J2_126_3477_n1634,
         DP_OP_424J2_126_3477_n1633, DP_OP_424J2_126_3477_n1632,
         DP_OP_424J2_126_3477_n1631, DP_OP_424J2_126_3477_n1630,
         DP_OP_424J2_126_3477_n1629, DP_OP_424J2_126_3477_n1628,
         DP_OP_424J2_126_3477_n1627, DP_OP_424J2_126_3477_n1626,
         DP_OP_424J2_126_3477_n1625, DP_OP_424J2_126_3477_n1624,
         DP_OP_424J2_126_3477_n1623, DP_OP_424J2_126_3477_n1622,
         DP_OP_424J2_126_3477_n1621, DP_OP_424J2_126_3477_n1620,
         DP_OP_424J2_126_3477_n1619, DP_OP_424J2_126_3477_n1618,
         DP_OP_424J2_126_3477_n1617, DP_OP_424J2_126_3477_n1616,
         DP_OP_424J2_126_3477_n1615, DP_OP_424J2_126_3477_n1614,
         DP_OP_424J2_126_3477_n1613, DP_OP_424J2_126_3477_n1612,
         DP_OP_424J2_126_3477_n1611, DP_OP_424J2_126_3477_n1610,
         DP_OP_424J2_126_3477_n1609, DP_OP_424J2_126_3477_n1608,
         DP_OP_424J2_126_3477_n1607, DP_OP_424J2_126_3477_n1606,
         DP_OP_424J2_126_3477_n1605, DP_OP_424J2_126_3477_n1604,
         DP_OP_424J2_126_3477_n1603, DP_OP_424J2_126_3477_n1602,
         DP_OP_424J2_126_3477_n1601, DP_OP_424J2_126_3477_n1600,
         DP_OP_424J2_126_3477_n1599, DP_OP_424J2_126_3477_n1598,
         DP_OP_424J2_126_3477_n1597, DP_OP_424J2_126_3477_n1596,
         DP_OP_424J2_126_3477_n1595, DP_OP_424J2_126_3477_n1594,
         DP_OP_424J2_126_3477_n1593, DP_OP_424J2_126_3477_n1592,
         DP_OP_424J2_126_3477_n1591, DP_OP_424J2_126_3477_n1590,
         DP_OP_424J2_126_3477_n1589, DP_OP_424J2_126_3477_n1588,
         DP_OP_424J2_126_3477_n1587, DP_OP_424J2_126_3477_n1586,
         DP_OP_424J2_126_3477_n1585, DP_OP_424J2_126_3477_n1584,
         DP_OP_424J2_126_3477_n1583, DP_OP_424J2_126_3477_n1582,
         DP_OP_424J2_126_3477_n1581, DP_OP_424J2_126_3477_n1580,
         DP_OP_424J2_126_3477_n1579, DP_OP_424J2_126_3477_n1578,
         DP_OP_424J2_126_3477_n1577, DP_OP_424J2_126_3477_n1576,
         DP_OP_424J2_126_3477_n1575, DP_OP_424J2_126_3477_n1574,
         DP_OP_424J2_126_3477_n1573, DP_OP_424J2_126_3477_n1572,
         DP_OP_424J2_126_3477_n1571, DP_OP_424J2_126_3477_n1570,
         DP_OP_424J2_126_3477_n1569, DP_OP_424J2_126_3477_n1568,
         DP_OP_424J2_126_3477_n1567, DP_OP_424J2_126_3477_n1566,
         DP_OP_424J2_126_3477_n1565, DP_OP_424J2_126_3477_n1564,
         DP_OP_424J2_126_3477_n1563, DP_OP_424J2_126_3477_n1562,
         DP_OP_424J2_126_3477_n1561, DP_OP_424J2_126_3477_n1560,
         DP_OP_424J2_126_3477_n1559, DP_OP_424J2_126_3477_n1558,
         DP_OP_424J2_126_3477_n1557, DP_OP_424J2_126_3477_n1556,
         DP_OP_424J2_126_3477_n1555, DP_OP_424J2_126_3477_n1554,
         DP_OP_424J2_126_3477_n1553, DP_OP_424J2_126_3477_n1552,
         DP_OP_424J2_126_3477_n1551, DP_OP_424J2_126_3477_n1550,
         DP_OP_424J2_126_3477_n1549, DP_OP_424J2_126_3477_n1548,
         DP_OP_424J2_126_3477_n1547, DP_OP_424J2_126_3477_n1546,
         DP_OP_424J2_126_3477_n1545, DP_OP_424J2_126_3477_n1544,
         DP_OP_424J2_126_3477_n1543, DP_OP_424J2_126_3477_n1542,
         DP_OP_424J2_126_3477_n1541, DP_OP_424J2_126_3477_n1540,
         DP_OP_424J2_126_3477_n1539, DP_OP_424J2_126_3477_n1538,
         DP_OP_424J2_126_3477_n1537, DP_OP_424J2_126_3477_n1536,
         DP_OP_424J2_126_3477_n1535, DP_OP_424J2_126_3477_n1534,
         DP_OP_424J2_126_3477_n1533, DP_OP_424J2_126_3477_n1532,
         DP_OP_424J2_126_3477_n1531, DP_OP_424J2_126_3477_n1530,
         DP_OP_424J2_126_3477_n1529, DP_OP_424J2_126_3477_n1528,
         DP_OP_424J2_126_3477_n1527, DP_OP_424J2_126_3477_n1526,
         DP_OP_424J2_126_3477_n1525, DP_OP_424J2_126_3477_n1524,
         DP_OP_424J2_126_3477_n1523, DP_OP_424J2_126_3477_n1522,
         DP_OP_424J2_126_3477_n1521, DP_OP_424J2_126_3477_n1520,
         DP_OP_424J2_126_3477_n1519, DP_OP_424J2_126_3477_n1518,
         DP_OP_424J2_126_3477_n1517, DP_OP_424J2_126_3477_n1516,
         DP_OP_424J2_126_3477_n1515, DP_OP_424J2_126_3477_n1514,
         DP_OP_424J2_126_3477_n1513, DP_OP_424J2_126_3477_n1512,
         DP_OP_424J2_126_3477_n1511, DP_OP_424J2_126_3477_n1510,
         DP_OP_424J2_126_3477_n1509, DP_OP_424J2_126_3477_n1508,
         DP_OP_424J2_126_3477_n1507, DP_OP_424J2_126_3477_n1506,
         DP_OP_424J2_126_3477_n1505, DP_OP_424J2_126_3477_n1504,
         DP_OP_424J2_126_3477_n1503, DP_OP_424J2_126_3477_n1502,
         DP_OP_424J2_126_3477_n1501, DP_OP_424J2_126_3477_n1500,
         DP_OP_424J2_126_3477_n1499, DP_OP_424J2_126_3477_n1498,
         DP_OP_424J2_126_3477_n1497, DP_OP_424J2_126_3477_n1496,
         DP_OP_424J2_126_3477_n1495, DP_OP_424J2_126_3477_n1494,
         DP_OP_424J2_126_3477_n1493, DP_OP_424J2_126_3477_n1492,
         DP_OP_424J2_126_3477_n1491, DP_OP_424J2_126_3477_n1490,
         DP_OP_424J2_126_3477_n1489, DP_OP_424J2_126_3477_n1488,
         DP_OP_424J2_126_3477_n1487, DP_OP_424J2_126_3477_n1486,
         DP_OP_424J2_126_3477_n1485, DP_OP_424J2_126_3477_n1484,
         DP_OP_424J2_126_3477_n1483, DP_OP_424J2_126_3477_n1482,
         DP_OP_424J2_126_3477_n1481, DP_OP_424J2_126_3477_n1480,
         DP_OP_424J2_126_3477_n1479, DP_OP_424J2_126_3477_n1478,
         DP_OP_424J2_126_3477_n1477, DP_OP_424J2_126_3477_n1476,
         DP_OP_424J2_126_3477_n1475, DP_OP_424J2_126_3477_n1474,
         DP_OP_424J2_126_3477_n1473, DP_OP_424J2_126_3477_n1472,
         DP_OP_424J2_126_3477_n1471, DP_OP_424J2_126_3477_n1470,
         DP_OP_424J2_126_3477_n1469, DP_OP_424J2_126_3477_n1468,
         DP_OP_424J2_126_3477_n1467, DP_OP_424J2_126_3477_n1466,
         DP_OP_424J2_126_3477_n1465, DP_OP_424J2_126_3477_n1464,
         DP_OP_424J2_126_3477_n1463, DP_OP_424J2_126_3477_n1462,
         DP_OP_424J2_126_3477_n1461, DP_OP_424J2_126_3477_n1460,
         DP_OP_424J2_126_3477_n1459, DP_OP_424J2_126_3477_n1458,
         DP_OP_424J2_126_3477_n1457, DP_OP_424J2_126_3477_n1456,
         DP_OP_424J2_126_3477_n1455, DP_OP_424J2_126_3477_n1454,
         DP_OP_424J2_126_3477_n1453, DP_OP_424J2_126_3477_n1452,
         DP_OP_424J2_126_3477_n1451, DP_OP_424J2_126_3477_n1450,
         DP_OP_424J2_126_3477_n1449, DP_OP_424J2_126_3477_n1448,
         DP_OP_424J2_126_3477_n1447, DP_OP_424J2_126_3477_n1446,
         DP_OP_424J2_126_3477_n1445, DP_OP_424J2_126_3477_n1444,
         DP_OP_424J2_126_3477_n1443, DP_OP_424J2_126_3477_n1442,
         DP_OP_424J2_126_3477_n1441, DP_OP_424J2_126_3477_n1440,
         DP_OP_424J2_126_3477_n1439, DP_OP_424J2_126_3477_n1438,
         DP_OP_424J2_126_3477_n1437, DP_OP_424J2_126_3477_n1436,
         DP_OP_424J2_126_3477_n1435, DP_OP_424J2_126_3477_n1434,
         DP_OP_424J2_126_3477_n1433, DP_OP_424J2_126_3477_n1432,
         DP_OP_424J2_126_3477_n1431, DP_OP_424J2_126_3477_n1430,
         DP_OP_424J2_126_3477_n1429, DP_OP_424J2_126_3477_n1428,
         DP_OP_424J2_126_3477_n1427, DP_OP_424J2_126_3477_n1426,
         DP_OP_424J2_126_3477_n1425, DP_OP_424J2_126_3477_n1424,
         DP_OP_424J2_126_3477_n1423, DP_OP_424J2_126_3477_n1422,
         DP_OP_424J2_126_3477_n1421, DP_OP_424J2_126_3477_n1420,
         DP_OP_424J2_126_3477_n1419, DP_OP_424J2_126_3477_n1418,
         DP_OP_424J2_126_3477_n1417, DP_OP_424J2_126_3477_n1416,
         DP_OP_424J2_126_3477_n1415, DP_OP_424J2_126_3477_n1414,
         DP_OP_424J2_126_3477_n1413, DP_OP_424J2_126_3477_n1412,
         DP_OP_424J2_126_3477_n1411, DP_OP_424J2_126_3477_n1410,
         DP_OP_424J2_126_3477_n1409, DP_OP_424J2_126_3477_n1408,
         DP_OP_424J2_126_3477_n1407, DP_OP_424J2_126_3477_n1406,
         DP_OP_424J2_126_3477_n1405, DP_OP_424J2_126_3477_n1404,
         DP_OP_424J2_126_3477_n1403, DP_OP_424J2_126_3477_n1402,
         DP_OP_424J2_126_3477_n1401, DP_OP_424J2_126_3477_n1400,
         DP_OP_424J2_126_3477_n1399, DP_OP_424J2_126_3477_n1398,
         DP_OP_424J2_126_3477_n1397, DP_OP_424J2_126_3477_n1396,
         DP_OP_424J2_126_3477_n1395, DP_OP_424J2_126_3477_n1394,
         DP_OP_424J2_126_3477_n1393, DP_OP_424J2_126_3477_n1392,
         DP_OP_424J2_126_3477_n1391, DP_OP_424J2_126_3477_n1390,
         DP_OP_424J2_126_3477_n1389, DP_OP_424J2_126_3477_n1388,
         DP_OP_424J2_126_3477_n1387, DP_OP_424J2_126_3477_n1386,
         DP_OP_424J2_126_3477_n1385, DP_OP_424J2_126_3477_n1384,
         DP_OP_424J2_126_3477_n1383, DP_OP_424J2_126_3477_n1382,
         DP_OP_424J2_126_3477_n1381, DP_OP_424J2_126_3477_n1380,
         DP_OP_424J2_126_3477_n1379, DP_OP_424J2_126_3477_n1378,
         DP_OP_424J2_126_3477_n1377, DP_OP_424J2_126_3477_n1376,
         DP_OP_424J2_126_3477_n1375, DP_OP_424J2_126_3477_n1374,
         DP_OP_424J2_126_3477_n1373, DP_OP_424J2_126_3477_n1372,
         DP_OP_424J2_126_3477_n1371, DP_OP_424J2_126_3477_n1370,
         DP_OP_424J2_126_3477_n1369, DP_OP_424J2_126_3477_n1368,
         DP_OP_424J2_126_3477_n1367, DP_OP_424J2_126_3477_n1366,
         DP_OP_424J2_126_3477_n1365, DP_OP_424J2_126_3477_n1364,
         DP_OP_424J2_126_3477_n1363, DP_OP_424J2_126_3477_n1362,
         DP_OP_424J2_126_3477_n1361, DP_OP_424J2_126_3477_n1360,
         DP_OP_424J2_126_3477_n1359, DP_OP_424J2_126_3477_n1358,
         DP_OP_424J2_126_3477_n1357, DP_OP_424J2_126_3477_n1356,
         DP_OP_424J2_126_3477_n1355, DP_OP_424J2_126_3477_n1354,
         DP_OP_424J2_126_3477_n1353, DP_OP_424J2_126_3477_n1352,
         DP_OP_424J2_126_3477_n1351, DP_OP_424J2_126_3477_n1350,
         DP_OP_424J2_126_3477_n1349, DP_OP_424J2_126_3477_n1348,
         DP_OP_424J2_126_3477_n1347, DP_OP_424J2_126_3477_n1346,
         DP_OP_424J2_126_3477_n1345, DP_OP_424J2_126_3477_n1344,
         DP_OP_424J2_126_3477_n1343, DP_OP_424J2_126_3477_n1342,
         DP_OP_424J2_126_3477_n1341, DP_OP_424J2_126_3477_n1340,
         DP_OP_424J2_126_3477_n1339, DP_OP_424J2_126_3477_n1338,
         DP_OP_424J2_126_3477_n1337, DP_OP_424J2_126_3477_n1336,
         DP_OP_424J2_126_3477_n1335, DP_OP_424J2_126_3477_n1334,
         DP_OP_424J2_126_3477_n1333, DP_OP_424J2_126_3477_n1332,
         DP_OP_424J2_126_3477_n1331, DP_OP_424J2_126_3477_n1330,
         DP_OP_424J2_126_3477_n1329, DP_OP_424J2_126_3477_n1328,
         DP_OP_424J2_126_3477_n1327, DP_OP_424J2_126_3477_n1326,
         DP_OP_424J2_126_3477_n1325, DP_OP_424J2_126_3477_n1324,
         DP_OP_424J2_126_3477_n1323, DP_OP_424J2_126_3477_n1322,
         DP_OP_424J2_126_3477_n1321, DP_OP_424J2_126_3477_n1320,
         DP_OP_424J2_126_3477_n1319, DP_OP_424J2_126_3477_n1318,
         DP_OP_424J2_126_3477_n1317, DP_OP_424J2_126_3477_n1316,
         DP_OP_424J2_126_3477_n1315, DP_OP_424J2_126_3477_n1314,
         DP_OP_424J2_126_3477_n1313, DP_OP_424J2_126_3477_n1312,
         DP_OP_424J2_126_3477_n1311, DP_OP_424J2_126_3477_n1310,
         DP_OP_424J2_126_3477_n1309, DP_OP_424J2_126_3477_n1308,
         DP_OP_424J2_126_3477_n1307, DP_OP_424J2_126_3477_n1306,
         DP_OP_424J2_126_3477_n1305, DP_OP_424J2_126_3477_n1304,
         DP_OP_424J2_126_3477_n1303, DP_OP_424J2_126_3477_n1302,
         DP_OP_424J2_126_3477_n1301, DP_OP_424J2_126_3477_n1300,
         DP_OP_424J2_126_3477_n1299, DP_OP_424J2_126_3477_n1298,
         DP_OP_424J2_126_3477_n1297, DP_OP_424J2_126_3477_n1296,
         DP_OP_424J2_126_3477_n1295, DP_OP_424J2_126_3477_n1294,
         DP_OP_424J2_126_3477_n1293, DP_OP_424J2_126_3477_n1292,
         DP_OP_424J2_126_3477_n1291, DP_OP_424J2_126_3477_n1290,
         DP_OP_424J2_126_3477_n1289, DP_OP_424J2_126_3477_n1288,
         DP_OP_424J2_126_3477_n1287, DP_OP_424J2_126_3477_n1286,
         DP_OP_424J2_126_3477_n1285, DP_OP_424J2_126_3477_n1284,
         DP_OP_424J2_126_3477_n1283, DP_OP_424J2_126_3477_n1282,
         DP_OP_424J2_126_3477_n1281, DP_OP_424J2_126_3477_n1280,
         DP_OP_424J2_126_3477_n1279, DP_OP_424J2_126_3477_n1278,
         DP_OP_424J2_126_3477_n1277, DP_OP_424J2_126_3477_n1276,
         DP_OP_424J2_126_3477_n1275, DP_OP_424J2_126_3477_n1274,
         DP_OP_424J2_126_3477_n1273, DP_OP_424J2_126_3477_n1272,
         DP_OP_424J2_126_3477_n1271, DP_OP_424J2_126_3477_n1270,
         DP_OP_424J2_126_3477_n1269, DP_OP_424J2_126_3477_n1268,
         DP_OP_424J2_126_3477_n1267, DP_OP_424J2_126_3477_n1266,
         DP_OP_424J2_126_3477_n1265, DP_OP_424J2_126_3477_n1264,
         DP_OP_424J2_126_3477_n1263, DP_OP_424J2_126_3477_n1262,
         DP_OP_424J2_126_3477_n1261, DP_OP_424J2_126_3477_n1260,
         DP_OP_424J2_126_3477_n1259, DP_OP_424J2_126_3477_n1258,
         DP_OP_424J2_126_3477_n1257, DP_OP_424J2_126_3477_n1256,
         DP_OP_424J2_126_3477_n1255, DP_OP_424J2_126_3477_n1254,
         DP_OP_424J2_126_3477_n1253, DP_OP_424J2_126_3477_n1252,
         DP_OP_424J2_126_3477_n1251, DP_OP_424J2_126_3477_n1250,
         DP_OP_424J2_126_3477_n1249, DP_OP_424J2_126_3477_n1248,
         DP_OP_424J2_126_3477_n1247, DP_OP_424J2_126_3477_n1246,
         DP_OP_424J2_126_3477_n1245, DP_OP_424J2_126_3477_n1244,
         DP_OP_424J2_126_3477_n1243, DP_OP_424J2_126_3477_n1242,
         DP_OP_424J2_126_3477_n1241, DP_OP_424J2_126_3477_n1240,
         DP_OP_424J2_126_3477_n1239, DP_OP_424J2_126_3477_n1238,
         DP_OP_424J2_126_3477_n1237, DP_OP_424J2_126_3477_n1236,
         DP_OP_424J2_126_3477_n1235, DP_OP_424J2_126_3477_n1234,
         DP_OP_424J2_126_3477_n1233, DP_OP_424J2_126_3477_n1232,
         DP_OP_424J2_126_3477_n1231, DP_OP_424J2_126_3477_n1230,
         DP_OP_424J2_126_3477_n1229, DP_OP_424J2_126_3477_n1228,
         DP_OP_424J2_126_3477_n1227, DP_OP_424J2_126_3477_n1226,
         DP_OP_424J2_126_3477_n1225, DP_OP_424J2_126_3477_n1224,
         DP_OP_424J2_126_3477_n1223, DP_OP_424J2_126_3477_n1222,
         DP_OP_424J2_126_3477_n1221, DP_OP_424J2_126_3477_n1220,
         DP_OP_424J2_126_3477_n1219, DP_OP_424J2_126_3477_n1218,
         DP_OP_424J2_126_3477_n1217, DP_OP_424J2_126_3477_n1216,
         DP_OP_424J2_126_3477_n1215, DP_OP_424J2_126_3477_n1214,
         DP_OP_424J2_126_3477_n1213, DP_OP_424J2_126_3477_n1212,
         DP_OP_424J2_126_3477_n1211, DP_OP_424J2_126_3477_n1210,
         DP_OP_424J2_126_3477_n1209, DP_OP_424J2_126_3477_n1208,
         DP_OP_424J2_126_3477_n1207, DP_OP_424J2_126_3477_n1206,
         DP_OP_424J2_126_3477_n1205, DP_OP_424J2_126_3477_n1204,
         DP_OP_424J2_126_3477_n1203, DP_OP_424J2_126_3477_n1202,
         DP_OP_424J2_126_3477_n1201, DP_OP_424J2_126_3477_n1200,
         DP_OP_424J2_126_3477_n1199, DP_OP_424J2_126_3477_n1198,
         DP_OP_424J2_126_3477_n1197, DP_OP_424J2_126_3477_n1196,
         DP_OP_424J2_126_3477_n1195, DP_OP_424J2_126_3477_n1194,
         DP_OP_424J2_126_3477_n1193, DP_OP_424J2_126_3477_n1192,
         DP_OP_424J2_126_3477_n1191, DP_OP_424J2_126_3477_n1190,
         DP_OP_424J2_126_3477_n1189, DP_OP_424J2_126_3477_n1188,
         DP_OP_424J2_126_3477_n1187, DP_OP_424J2_126_3477_n1186,
         DP_OP_424J2_126_3477_n1185, DP_OP_424J2_126_3477_n1184,
         DP_OP_424J2_126_3477_n1183, DP_OP_424J2_126_3477_n1182,
         DP_OP_424J2_126_3477_n1181, DP_OP_424J2_126_3477_n1180,
         DP_OP_424J2_126_3477_n1179, DP_OP_424J2_126_3477_n1178,
         DP_OP_424J2_126_3477_n1177, DP_OP_424J2_126_3477_n1176,
         DP_OP_424J2_126_3477_n1175, DP_OP_424J2_126_3477_n1174,
         DP_OP_424J2_126_3477_n1173, DP_OP_424J2_126_3477_n1172,
         DP_OP_424J2_126_3477_n1171, DP_OP_424J2_126_3477_n1170,
         DP_OP_424J2_126_3477_n1169, DP_OP_424J2_126_3477_n1168,
         DP_OP_424J2_126_3477_n1167, DP_OP_424J2_126_3477_n1166,
         DP_OP_424J2_126_3477_n1165, DP_OP_424J2_126_3477_n1164,
         DP_OP_424J2_126_3477_n1163, DP_OP_424J2_126_3477_n1162,
         DP_OP_424J2_126_3477_n1161, DP_OP_424J2_126_3477_n1160,
         DP_OP_424J2_126_3477_n1159, DP_OP_424J2_126_3477_n1158,
         DP_OP_424J2_126_3477_n1157, DP_OP_424J2_126_3477_n1156,
         DP_OP_424J2_126_3477_n1155, DP_OP_424J2_126_3477_n1154,
         DP_OP_424J2_126_3477_n1153, DP_OP_424J2_126_3477_n1152,
         DP_OP_424J2_126_3477_n1151, DP_OP_424J2_126_3477_n1150,
         DP_OP_424J2_126_3477_n1149, DP_OP_424J2_126_3477_n1148,
         DP_OP_424J2_126_3477_n1147, DP_OP_424J2_126_3477_n1146,
         DP_OP_424J2_126_3477_n1145, DP_OP_424J2_126_3477_n1144,
         DP_OP_424J2_126_3477_n1143, DP_OP_424J2_126_3477_n1142,
         DP_OP_424J2_126_3477_n1141, DP_OP_424J2_126_3477_n1140,
         DP_OP_424J2_126_3477_n1139, DP_OP_424J2_126_3477_n1138,
         DP_OP_424J2_126_3477_n1137, DP_OP_424J2_126_3477_n1136,
         DP_OP_424J2_126_3477_n1135, DP_OP_424J2_126_3477_n1134,
         DP_OP_424J2_126_3477_n1133, DP_OP_424J2_126_3477_n1132,
         DP_OP_424J2_126_3477_n1131, DP_OP_424J2_126_3477_n1130,
         DP_OP_424J2_126_3477_n1129, DP_OP_424J2_126_3477_n1128,
         DP_OP_424J2_126_3477_n1127, DP_OP_424J2_126_3477_n1126,
         DP_OP_424J2_126_3477_n1125, DP_OP_424J2_126_3477_n1124,
         DP_OP_424J2_126_3477_n1123, DP_OP_424J2_126_3477_n1122,
         DP_OP_424J2_126_3477_n1121, DP_OP_424J2_126_3477_n1120,
         DP_OP_424J2_126_3477_n1119, DP_OP_424J2_126_3477_n1118,
         DP_OP_424J2_126_3477_n1117, DP_OP_424J2_126_3477_n1116,
         DP_OP_424J2_126_3477_n1115, DP_OP_424J2_126_3477_n1114,
         DP_OP_424J2_126_3477_n1113, DP_OP_424J2_126_3477_n1112,
         DP_OP_424J2_126_3477_n1111, DP_OP_424J2_126_3477_n1110,
         DP_OP_424J2_126_3477_n1109, DP_OP_424J2_126_3477_n1108,
         DP_OP_424J2_126_3477_n1107, DP_OP_424J2_126_3477_n1106,
         DP_OP_424J2_126_3477_n1105, DP_OP_424J2_126_3477_n1104,
         DP_OP_424J2_126_3477_n1103, DP_OP_424J2_126_3477_n1102,
         DP_OP_424J2_126_3477_n1101, DP_OP_424J2_126_3477_n1100,
         DP_OP_424J2_126_3477_n1099, DP_OP_424J2_126_3477_n1098,
         DP_OP_424J2_126_3477_n1097, DP_OP_424J2_126_3477_n1096,
         DP_OP_424J2_126_3477_n1095, DP_OP_424J2_126_3477_n1094,
         DP_OP_424J2_126_3477_n1093, DP_OP_424J2_126_3477_n1092,
         DP_OP_424J2_126_3477_n1091, DP_OP_424J2_126_3477_n1090,
         DP_OP_424J2_126_3477_n1089, DP_OP_424J2_126_3477_n1088,
         DP_OP_424J2_126_3477_n1087, DP_OP_424J2_126_3477_n1086,
         DP_OP_424J2_126_3477_n1085, DP_OP_424J2_126_3477_n1084,
         DP_OP_424J2_126_3477_n1083, DP_OP_424J2_126_3477_n1082,
         DP_OP_424J2_126_3477_n1081, DP_OP_424J2_126_3477_n1080,
         DP_OP_424J2_126_3477_n1079, DP_OP_424J2_126_3477_n1078,
         DP_OP_424J2_126_3477_n1077, DP_OP_424J2_126_3477_n1076,
         DP_OP_424J2_126_3477_n1075, DP_OP_424J2_126_3477_n1074,
         DP_OP_424J2_126_3477_n1073, DP_OP_424J2_126_3477_n1072,
         DP_OP_424J2_126_3477_n1071, DP_OP_424J2_126_3477_n1070,
         DP_OP_424J2_126_3477_n1069, DP_OP_424J2_126_3477_n1068,
         DP_OP_424J2_126_3477_n1067, DP_OP_424J2_126_3477_n1066,
         DP_OP_424J2_126_3477_n1065, DP_OP_424J2_126_3477_n1064,
         DP_OP_424J2_126_3477_n1063, DP_OP_424J2_126_3477_n1062,
         DP_OP_424J2_126_3477_n1061, DP_OP_424J2_126_3477_n1060,
         DP_OP_424J2_126_3477_n1059, DP_OP_424J2_126_3477_n1058,
         DP_OP_424J2_126_3477_n1057, DP_OP_424J2_126_3477_n1056,
         DP_OP_424J2_126_3477_n1055, DP_OP_424J2_126_3477_n1054,
         DP_OP_424J2_126_3477_n1053, DP_OP_424J2_126_3477_n1052,
         DP_OP_424J2_126_3477_n1051, DP_OP_424J2_126_3477_n1050,
         DP_OP_424J2_126_3477_n1049, DP_OP_424J2_126_3477_n1048,
         DP_OP_424J2_126_3477_n1047, DP_OP_424J2_126_3477_n1046,
         DP_OP_424J2_126_3477_n1045, DP_OP_424J2_126_3477_n1044,
         DP_OP_424J2_126_3477_n1043, DP_OP_424J2_126_3477_n1042,
         DP_OP_424J2_126_3477_n1041, DP_OP_424J2_126_3477_n1040,
         DP_OP_424J2_126_3477_n1039, DP_OP_424J2_126_3477_n1038,
         DP_OP_424J2_126_3477_n1037, DP_OP_424J2_126_3477_n1036,
         DP_OP_424J2_126_3477_n1035, DP_OP_424J2_126_3477_n1034,
         DP_OP_424J2_126_3477_n1033, DP_OP_424J2_126_3477_n1032,
         DP_OP_424J2_126_3477_n1031, DP_OP_424J2_126_3477_n1030,
         DP_OP_424J2_126_3477_n1029, DP_OP_424J2_126_3477_n1028,
         DP_OP_424J2_126_3477_n1027, DP_OP_424J2_126_3477_n1026,
         DP_OP_424J2_126_3477_n1025, DP_OP_424J2_126_3477_n1024,
         DP_OP_424J2_126_3477_n1023, DP_OP_424J2_126_3477_n1022,
         DP_OP_424J2_126_3477_n1021, DP_OP_424J2_126_3477_n1020,
         DP_OP_424J2_126_3477_n1019, DP_OP_424J2_126_3477_n1018,
         DP_OP_424J2_126_3477_n1017, DP_OP_424J2_126_3477_n1016,
         DP_OP_424J2_126_3477_n1015, DP_OP_424J2_126_3477_n1014,
         DP_OP_424J2_126_3477_n1013, DP_OP_424J2_126_3477_n1012,
         DP_OP_424J2_126_3477_n1011, DP_OP_424J2_126_3477_n1010,
         DP_OP_424J2_126_3477_n1009, DP_OP_424J2_126_3477_n1008,
         DP_OP_424J2_126_3477_n1007, DP_OP_424J2_126_3477_n1006,
         DP_OP_424J2_126_3477_n1005, DP_OP_424J2_126_3477_n1004,
         DP_OP_424J2_126_3477_n1003, DP_OP_424J2_126_3477_n1002,
         DP_OP_424J2_126_3477_n1001, DP_OP_424J2_126_3477_n1000,
         DP_OP_424J2_126_3477_n999, DP_OP_424J2_126_3477_n998,
         DP_OP_424J2_126_3477_n997, DP_OP_424J2_126_3477_n996,
         DP_OP_424J2_126_3477_n995, DP_OP_424J2_126_3477_n994,
         DP_OP_424J2_126_3477_n993, DP_OP_424J2_126_3477_n992,
         DP_OP_424J2_126_3477_n991, DP_OP_424J2_126_3477_n990,
         DP_OP_424J2_126_3477_n989, DP_OP_424J2_126_3477_n988,
         DP_OP_424J2_126_3477_n987, DP_OP_424J2_126_3477_n986,
         DP_OP_424J2_126_3477_n985, DP_OP_424J2_126_3477_n984,
         DP_OP_424J2_126_3477_n983, DP_OP_424J2_126_3477_n982,
         DP_OP_424J2_126_3477_n981, DP_OP_424J2_126_3477_n980,
         DP_OP_424J2_126_3477_n979, DP_OP_424J2_126_3477_n978,
         DP_OP_424J2_126_3477_n977, DP_OP_424J2_126_3477_n976,
         DP_OP_424J2_126_3477_n975, DP_OP_424J2_126_3477_n974,
         DP_OP_424J2_126_3477_n973, DP_OP_424J2_126_3477_n972,
         DP_OP_424J2_126_3477_n971, DP_OP_424J2_126_3477_n970,
         DP_OP_424J2_126_3477_n969, DP_OP_424J2_126_3477_n968,
         DP_OP_424J2_126_3477_n967, DP_OP_424J2_126_3477_n966,
         DP_OP_424J2_126_3477_n965, DP_OP_424J2_126_3477_n964,
         DP_OP_424J2_126_3477_n963, DP_OP_424J2_126_3477_n962,
         DP_OP_424J2_126_3477_n961, DP_OP_424J2_126_3477_n960,
         DP_OP_424J2_126_3477_n959, DP_OP_424J2_126_3477_n958,
         DP_OP_424J2_126_3477_n957, DP_OP_424J2_126_3477_n956,
         DP_OP_424J2_126_3477_n955, DP_OP_424J2_126_3477_n954,
         DP_OP_424J2_126_3477_n953, DP_OP_424J2_126_3477_n952,
         DP_OP_424J2_126_3477_n951, DP_OP_424J2_126_3477_n950,
         DP_OP_424J2_126_3477_n949, DP_OP_424J2_126_3477_n948,
         DP_OP_424J2_126_3477_n947, DP_OP_424J2_126_3477_n946,
         DP_OP_424J2_126_3477_n945, DP_OP_424J2_126_3477_n944,
         DP_OP_424J2_126_3477_n943, DP_OP_424J2_126_3477_n942,
         DP_OP_424J2_126_3477_n941, DP_OP_424J2_126_3477_n940,
         DP_OP_424J2_126_3477_n939, DP_OP_424J2_126_3477_n938,
         DP_OP_424J2_126_3477_n937, DP_OP_424J2_126_3477_n936,
         DP_OP_424J2_126_3477_n935, DP_OP_424J2_126_3477_n934,
         DP_OP_424J2_126_3477_n933, DP_OP_424J2_126_3477_n932,
         DP_OP_424J2_126_3477_n931, DP_OP_424J2_126_3477_n930,
         DP_OP_424J2_126_3477_n929, DP_OP_424J2_126_3477_n928,
         DP_OP_424J2_126_3477_n927, DP_OP_424J2_126_3477_n926,
         DP_OP_424J2_126_3477_n925, DP_OP_424J2_126_3477_n924,
         DP_OP_424J2_126_3477_n923, DP_OP_424J2_126_3477_n922,
         DP_OP_424J2_126_3477_n921, DP_OP_424J2_126_3477_n920,
         DP_OP_424J2_126_3477_n919, DP_OP_424J2_126_3477_n918,
         DP_OP_424J2_126_3477_n917, DP_OP_424J2_126_3477_n916,
         DP_OP_424J2_126_3477_n915, DP_OP_424J2_126_3477_n914,
         DP_OP_424J2_126_3477_n913, DP_OP_424J2_126_3477_n912,
         DP_OP_424J2_126_3477_n911, DP_OP_424J2_126_3477_n910,
         DP_OP_424J2_126_3477_n909, DP_OP_424J2_126_3477_n908,
         DP_OP_424J2_126_3477_n907, DP_OP_424J2_126_3477_n906,
         DP_OP_424J2_126_3477_n905, DP_OP_424J2_126_3477_n904,
         DP_OP_424J2_126_3477_n903, DP_OP_424J2_126_3477_n902,
         DP_OP_424J2_126_3477_n901, DP_OP_424J2_126_3477_n900,
         DP_OP_424J2_126_3477_n899, DP_OP_424J2_126_3477_n898,
         DP_OP_424J2_126_3477_n897, DP_OP_424J2_126_3477_n896,
         DP_OP_424J2_126_3477_n895, DP_OP_424J2_126_3477_n894,
         DP_OP_424J2_126_3477_n893, DP_OP_424J2_126_3477_n892,
         DP_OP_424J2_126_3477_n891, DP_OP_424J2_126_3477_n890,
         DP_OP_424J2_126_3477_n889, DP_OP_424J2_126_3477_n888,
         DP_OP_424J2_126_3477_n887, DP_OP_424J2_126_3477_n886,
         DP_OP_424J2_126_3477_n885, DP_OP_424J2_126_3477_n884,
         DP_OP_424J2_126_3477_n883, DP_OP_424J2_126_3477_n882,
         DP_OP_424J2_126_3477_n881, DP_OP_424J2_126_3477_n880,
         DP_OP_424J2_126_3477_n879, DP_OP_424J2_126_3477_n878,
         DP_OP_424J2_126_3477_n877, DP_OP_424J2_126_3477_n876,
         DP_OP_424J2_126_3477_n875, DP_OP_424J2_126_3477_n874,
         DP_OP_424J2_126_3477_n873, DP_OP_424J2_126_3477_n872,
         DP_OP_424J2_126_3477_n871, DP_OP_424J2_126_3477_n870,
         DP_OP_424J2_126_3477_n869, DP_OP_424J2_126_3477_n868,
         DP_OP_424J2_126_3477_n867, DP_OP_424J2_126_3477_n866,
         DP_OP_424J2_126_3477_n865, DP_OP_424J2_126_3477_n864,
         DP_OP_424J2_126_3477_n863, DP_OP_424J2_126_3477_n862,
         DP_OP_424J2_126_3477_n861, DP_OP_424J2_126_3477_n860,
         DP_OP_424J2_126_3477_n859, DP_OP_424J2_126_3477_n858,
         DP_OP_424J2_126_3477_n857, DP_OP_424J2_126_3477_n856,
         DP_OP_424J2_126_3477_n855, DP_OP_424J2_126_3477_n854,
         DP_OP_424J2_126_3477_n853, DP_OP_424J2_126_3477_n852,
         DP_OP_424J2_126_3477_n851, DP_OP_424J2_126_3477_n850,
         DP_OP_424J2_126_3477_n849, DP_OP_424J2_126_3477_n848,
         DP_OP_424J2_126_3477_n847, DP_OP_424J2_126_3477_n846,
         DP_OP_424J2_126_3477_n845, DP_OP_424J2_126_3477_n844,
         DP_OP_424J2_126_3477_n843, DP_OP_424J2_126_3477_n842,
         DP_OP_424J2_126_3477_n841, DP_OP_424J2_126_3477_n840,
         DP_OP_424J2_126_3477_n839, DP_OP_424J2_126_3477_n838,
         DP_OP_424J2_126_3477_n837, DP_OP_424J2_126_3477_n836,
         DP_OP_424J2_126_3477_n835, DP_OP_424J2_126_3477_n834,
         DP_OP_424J2_126_3477_n833, DP_OP_424J2_126_3477_n832,
         DP_OP_424J2_126_3477_n831, DP_OP_424J2_126_3477_n830,
         DP_OP_424J2_126_3477_n829, DP_OP_424J2_126_3477_n828,
         DP_OP_424J2_126_3477_n827, DP_OP_424J2_126_3477_n826,
         DP_OP_424J2_126_3477_n825, DP_OP_424J2_126_3477_n824,
         DP_OP_424J2_126_3477_n823, DP_OP_424J2_126_3477_n822,
         DP_OP_424J2_126_3477_n821, DP_OP_424J2_126_3477_n820,
         DP_OP_424J2_126_3477_n819, DP_OP_424J2_126_3477_n818,
         DP_OP_424J2_126_3477_n817, DP_OP_424J2_126_3477_n816,
         DP_OP_424J2_126_3477_n815, DP_OP_424J2_126_3477_n814,
         DP_OP_424J2_126_3477_n813, DP_OP_424J2_126_3477_n812,
         DP_OP_424J2_126_3477_n811, DP_OP_424J2_126_3477_n810,
         DP_OP_424J2_126_3477_n809, DP_OP_424J2_126_3477_n808,
         DP_OP_424J2_126_3477_n807, DP_OP_424J2_126_3477_n806,
         DP_OP_424J2_126_3477_n805, DP_OP_424J2_126_3477_n804,
         DP_OP_424J2_126_3477_n803, DP_OP_424J2_126_3477_n802,
         DP_OP_424J2_126_3477_n801, DP_OP_424J2_126_3477_n800,
         DP_OP_424J2_126_3477_n799, DP_OP_424J2_126_3477_n798,
         DP_OP_424J2_126_3477_n797, DP_OP_424J2_126_3477_n796,
         DP_OP_424J2_126_3477_n795, DP_OP_424J2_126_3477_n794,
         DP_OP_424J2_126_3477_n793, DP_OP_424J2_126_3477_n792,
         DP_OP_424J2_126_3477_n791, DP_OP_424J2_126_3477_n790,
         DP_OP_424J2_126_3477_n789, DP_OP_424J2_126_3477_n788,
         DP_OP_424J2_126_3477_n787, DP_OP_424J2_126_3477_n786,
         DP_OP_424J2_126_3477_n785, DP_OP_424J2_126_3477_n784,
         DP_OP_424J2_126_3477_n783, DP_OP_424J2_126_3477_n782,
         DP_OP_424J2_126_3477_n781, DP_OP_424J2_126_3477_n780,
         DP_OP_424J2_126_3477_n779, DP_OP_424J2_126_3477_n778,
         DP_OP_424J2_126_3477_n777, DP_OP_424J2_126_3477_n776,
         DP_OP_424J2_126_3477_n775, DP_OP_424J2_126_3477_n774,
         DP_OP_424J2_126_3477_n773, DP_OP_424J2_126_3477_n772,
         DP_OP_424J2_126_3477_n771, DP_OP_424J2_126_3477_n770,
         DP_OP_424J2_126_3477_n769, DP_OP_424J2_126_3477_n768,
         DP_OP_424J2_126_3477_n767, DP_OP_424J2_126_3477_n766,
         DP_OP_424J2_126_3477_n765, DP_OP_424J2_126_3477_n764,
         DP_OP_424J2_126_3477_n763, DP_OP_424J2_126_3477_n762,
         DP_OP_424J2_126_3477_n761, DP_OP_424J2_126_3477_n760,
         DP_OP_424J2_126_3477_n759, DP_OP_424J2_126_3477_n758,
         DP_OP_424J2_126_3477_n757, DP_OP_424J2_126_3477_n756,
         DP_OP_424J2_126_3477_n755, DP_OP_424J2_126_3477_n754,
         DP_OP_424J2_126_3477_n753, DP_OP_424J2_126_3477_n752,
         DP_OP_424J2_126_3477_n751, DP_OP_424J2_126_3477_n750,
         DP_OP_424J2_126_3477_n749, DP_OP_424J2_126_3477_n748,
         DP_OP_424J2_126_3477_n747, DP_OP_424J2_126_3477_n746,
         DP_OP_424J2_126_3477_n745, DP_OP_424J2_126_3477_n744,
         DP_OP_424J2_126_3477_n743, DP_OP_424J2_126_3477_n742,
         DP_OP_424J2_126_3477_n741, DP_OP_424J2_126_3477_n740,
         DP_OP_424J2_126_3477_n739, DP_OP_424J2_126_3477_n738,
         DP_OP_424J2_126_3477_n737, DP_OP_424J2_126_3477_n736,
         DP_OP_424J2_126_3477_n735, DP_OP_424J2_126_3477_n734,
         DP_OP_424J2_126_3477_n733, DP_OP_424J2_126_3477_n732,
         DP_OP_424J2_126_3477_n731, DP_OP_424J2_126_3477_n730,
         DP_OP_424J2_126_3477_n729, DP_OP_424J2_126_3477_n728,
         DP_OP_424J2_126_3477_n727, DP_OP_424J2_126_3477_n726,
         DP_OP_424J2_126_3477_n725, DP_OP_424J2_126_3477_n724,
         DP_OP_424J2_126_3477_n723, DP_OP_424J2_126_3477_n722,
         DP_OP_424J2_126_3477_n721, DP_OP_424J2_126_3477_n720,
         DP_OP_424J2_126_3477_n719, DP_OP_424J2_126_3477_n718,
         DP_OP_424J2_126_3477_n717, DP_OP_424J2_126_3477_n716,
         DP_OP_424J2_126_3477_n715, DP_OP_424J2_126_3477_n714,
         DP_OP_424J2_126_3477_n713, DP_OP_424J2_126_3477_n712,
         DP_OP_424J2_126_3477_n711, DP_OP_424J2_126_3477_n710,
         DP_OP_424J2_126_3477_n709, DP_OP_424J2_126_3477_n708,
         DP_OP_424J2_126_3477_n707, DP_OP_424J2_126_3477_n706,
         DP_OP_424J2_126_3477_n705, DP_OP_424J2_126_3477_n704,
         DP_OP_424J2_126_3477_n703, DP_OP_424J2_126_3477_n702,
         DP_OP_424J2_126_3477_n701, DP_OP_424J2_126_3477_n700,
         DP_OP_424J2_126_3477_n699, DP_OP_424J2_126_3477_n698,
         DP_OP_424J2_126_3477_n697, DP_OP_424J2_126_3477_n696,
         DP_OP_424J2_126_3477_n695, DP_OP_424J2_126_3477_n694,
         DP_OP_424J2_126_3477_n693, DP_OP_424J2_126_3477_n692,
         DP_OP_424J2_126_3477_n691, DP_OP_424J2_126_3477_n690,
         DP_OP_424J2_126_3477_n689, DP_OP_424J2_126_3477_n688,
         DP_OP_424J2_126_3477_n687, DP_OP_424J2_126_3477_n686,
         DP_OP_424J2_126_3477_n685, DP_OP_424J2_126_3477_n684,
         DP_OP_424J2_126_3477_n683, DP_OP_424J2_126_3477_n682,
         DP_OP_424J2_126_3477_n681, DP_OP_424J2_126_3477_n680,
         DP_OP_424J2_126_3477_n679, DP_OP_424J2_126_3477_n678,
         DP_OP_424J2_126_3477_n677, DP_OP_424J2_126_3477_n676,
         DP_OP_424J2_126_3477_n675, DP_OP_424J2_126_3477_n674,
         DP_OP_424J2_126_3477_n673, DP_OP_424J2_126_3477_n672,
         DP_OP_424J2_126_3477_n671, DP_OP_424J2_126_3477_n670,
         DP_OP_424J2_126_3477_n669, DP_OP_424J2_126_3477_n668,
         DP_OP_424J2_126_3477_n667, DP_OP_424J2_126_3477_n666,
         DP_OP_424J2_126_3477_n665, DP_OP_424J2_126_3477_n664,
         DP_OP_424J2_126_3477_n663, DP_OP_424J2_126_3477_n662,
         DP_OP_424J2_126_3477_n661, DP_OP_424J2_126_3477_n660,
         DP_OP_424J2_126_3477_n659, DP_OP_424J2_126_3477_n658,
         DP_OP_424J2_126_3477_n657, DP_OP_424J2_126_3477_n656,
         DP_OP_424J2_126_3477_n655, DP_OP_424J2_126_3477_n654,
         DP_OP_424J2_126_3477_n653, DP_OP_424J2_126_3477_n652,
         DP_OP_424J2_126_3477_n651, DP_OP_424J2_126_3477_n650,
         DP_OP_424J2_126_3477_n649, DP_OP_424J2_126_3477_n648,
         DP_OP_424J2_126_3477_n647, DP_OP_424J2_126_3477_n646,
         DP_OP_424J2_126_3477_n645, DP_OP_424J2_126_3477_n644,
         DP_OP_424J2_126_3477_n643, DP_OP_424J2_126_3477_n642,
         DP_OP_424J2_126_3477_n641, DP_OP_424J2_126_3477_n640,
         DP_OP_424J2_126_3477_n639, DP_OP_424J2_126_3477_n638,
         DP_OP_424J2_126_3477_n637, DP_OP_424J2_126_3477_n636,
         DP_OP_424J2_126_3477_n635, DP_OP_424J2_126_3477_n634,
         DP_OP_424J2_126_3477_n633, DP_OP_424J2_126_3477_n632,
         DP_OP_424J2_126_3477_n631, DP_OP_424J2_126_3477_n630,
         DP_OP_424J2_126_3477_n629, DP_OP_424J2_126_3477_n628,
         DP_OP_424J2_126_3477_n627, DP_OP_424J2_126_3477_n626,
         DP_OP_424J2_126_3477_n625, DP_OP_424J2_126_3477_n624,
         DP_OP_424J2_126_3477_n623, DP_OP_424J2_126_3477_n622,
         DP_OP_424J2_126_3477_n621, DP_OP_424J2_126_3477_n620,
         DP_OP_424J2_126_3477_n619, DP_OP_424J2_126_3477_n618,
         DP_OP_424J2_126_3477_n617, DP_OP_424J2_126_3477_n616,
         DP_OP_424J2_126_3477_n615, DP_OP_424J2_126_3477_n614,
         DP_OP_424J2_126_3477_n613, DP_OP_424J2_126_3477_n612,
         DP_OP_424J2_126_3477_n611, DP_OP_424J2_126_3477_n610,
         DP_OP_424J2_126_3477_n609, DP_OP_424J2_126_3477_n608,
         DP_OP_424J2_126_3477_n607, DP_OP_424J2_126_3477_n606,
         DP_OP_424J2_126_3477_n605, DP_OP_424J2_126_3477_n604,
         DP_OP_424J2_126_3477_n603, DP_OP_424J2_126_3477_n602,
         DP_OP_424J2_126_3477_n601, DP_OP_424J2_126_3477_n600,
         DP_OP_424J2_126_3477_n599, DP_OP_424J2_126_3477_n598,
         DP_OP_424J2_126_3477_n597, DP_OP_424J2_126_3477_n596,
         DP_OP_424J2_126_3477_n595, DP_OP_424J2_126_3477_n594,
         DP_OP_424J2_126_3477_n593, DP_OP_424J2_126_3477_n592,
         DP_OP_424J2_126_3477_n591, DP_OP_424J2_126_3477_n590,
         DP_OP_424J2_126_3477_n589, DP_OP_424J2_126_3477_n588,
         DP_OP_424J2_126_3477_n587, DP_OP_424J2_126_3477_n586,
         DP_OP_424J2_126_3477_n585, DP_OP_424J2_126_3477_n584,
         DP_OP_424J2_126_3477_n583, DP_OP_424J2_126_3477_n582,
         DP_OP_424J2_126_3477_n581, DP_OP_424J2_126_3477_n580,
         DP_OP_424J2_126_3477_n579, DP_OP_424J2_126_3477_n578,
         DP_OP_424J2_126_3477_n577, DP_OP_424J2_126_3477_n576,
         DP_OP_424J2_126_3477_n575, DP_OP_424J2_126_3477_n574,
         DP_OP_424J2_126_3477_n573, DP_OP_424J2_126_3477_n572,
         DP_OP_424J2_126_3477_n571, DP_OP_424J2_126_3477_n570,
         DP_OP_424J2_126_3477_n569, DP_OP_424J2_126_3477_n568,
         DP_OP_424J2_126_3477_n567, DP_OP_424J2_126_3477_n566,
         DP_OP_424J2_126_3477_n565, DP_OP_424J2_126_3477_n564,
         DP_OP_424J2_126_3477_n563, DP_OP_424J2_126_3477_n562,
         DP_OP_424J2_126_3477_n561, DP_OP_424J2_126_3477_n560,
         DP_OP_424J2_126_3477_n559, DP_OP_424J2_126_3477_n558,
         DP_OP_424J2_126_3477_n557, DP_OP_424J2_126_3477_n556,
         DP_OP_424J2_126_3477_n555, DP_OP_424J2_126_3477_n554,
         DP_OP_424J2_126_3477_n553, DP_OP_424J2_126_3477_n552,
         DP_OP_424J2_126_3477_n551, DP_OP_424J2_126_3477_n550,
         DP_OP_424J2_126_3477_n549, DP_OP_424J2_126_3477_n548,
         DP_OP_424J2_126_3477_n547, DP_OP_424J2_126_3477_n546,
         DP_OP_424J2_126_3477_n545, DP_OP_424J2_126_3477_n544,
         DP_OP_424J2_126_3477_n543, DP_OP_424J2_126_3477_n542,
         DP_OP_424J2_126_3477_n541, DP_OP_424J2_126_3477_n540,
         DP_OP_424J2_126_3477_n539, DP_OP_424J2_126_3477_n538,
         DP_OP_424J2_126_3477_n537, DP_OP_424J2_126_3477_n536,
         DP_OP_424J2_126_3477_n535, DP_OP_424J2_126_3477_n534,
         DP_OP_424J2_126_3477_n533, DP_OP_424J2_126_3477_n532,
         DP_OP_424J2_126_3477_n531, DP_OP_424J2_126_3477_n530,
         DP_OP_424J2_126_3477_n529, DP_OP_424J2_126_3477_n528,
         DP_OP_424J2_126_3477_n527, DP_OP_424J2_126_3477_n526,
         DP_OP_424J2_126_3477_n525, DP_OP_424J2_126_3477_n524,
         DP_OP_424J2_126_3477_n523, DP_OP_424J2_126_3477_n522,
         DP_OP_424J2_126_3477_n521, DP_OP_424J2_126_3477_n520,
         DP_OP_424J2_126_3477_n519, DP_OP_424J2_126_3477_n518,
         DP_OP_424J2_126_3477_n517, DP_OP_424J2_126_3477_n516,
         DP_OP_424J2_126_3477_n515, DP_OP_424J2_126_3477_n514,
         DP_OP_424J2_126_3477_n513, DP_OP_424J2_126_3477_n512,
         DP_OP_424J2_126_3477_n511, DP_OP_424J2_126_3477_n510,
         DP_OP_424J2_126_3477_n509, DP_OP_424J2_126_3477_n508,
         DP_OP_424J2_126_3477_n507, DP_OP_424J2_126_3477_n506,
         DP_OP_424J2_126_3477_n505, DP_OP_424J2_126_3477_n504,
         DP_OP_424J2_126_3477_n503, DP_OP_424J2_126_3477_n502,
         DP_OP_424J2_126_3477_n501, DP_OP_424J2_126_3477_n500,
         DP_OP_424J2_126_3477_n499, DP_OP_424J2_126_3477_n498,
         DP_OP_424J2_126_3477_n497, DP_OP_424J2_126_3477_n496,
         DP_OP_424J2_126_3477_n495, DP_OP_424J2_126_3477_n494,
         DP_OP_424J2_126_3477_n493, DP_OP_424J2_126_3477_n492,
         DP_OP_424J2_126_3477_n491, DP_OP_424J2_126_3477_n490,
         DP_OP_424J2_126_3477_n489, DP_OP_424J2_126_3477_n488,
         DP_OP_424J2_126_3477_n487, DP_OP_424J2_126_3477_n486,
         DP_OP_424J2_126_3477_n485, DP_OP_424J2_126_3477_n484,
         DP_OP_424J2_126_3477_n483, DP_OP_424J2_126_3477_n482,
         DP_OP_424J2_126_3477_n481, DP_OP_424J2_126_3477_n480,
         DP_OP_424J2_126_3477_n479, DP_OP_424J2_126_3477_n478,
         DP_OP_424J2_126_3477_n477, DP_OP_424J2_126_3477_n476,
         DP_OP_424J2_126_3477_n475, DP_OP_424J2_126_3477_n474,
         DP_OP_424J2_126_3477_n473, DP_OP_424J2_126_3477_n472,
         DP_OP_424J2_126_3477_n471, DP_OP_424J2_126_3477_n470,
         DP_OP_424J2_126_3477_n469, DP_OP_424J2_126_3477_n468,
         DP_OP_424J2_126_3477_n467, DP_OP_424J2_126_3477_n466,
         DP_OP_424J2_126_3477_n465, DP_OP_424J2_126_3477_n464,
         DP_OP_424J2_126_3477_n463, DP_OP_424J2_126_3477_n462,
         DP_OP_424J2_126_3477_n461, DP_OP_424J2_126_3477_n460,
         DP_OP_424J2_126_3477_n459, DP_OP_424J2_126_3477_n458,
         DP_OP_424J2_126_3477_n457, DP_OP_424J2_126_3477_n456,
         DP_OP_424J2_126_3477_n455, DP_OP_424J2_126_3477_n454,
         DP_OP_424J2_126_3477_n453, DP_OP_424J2_126_3477_n452,
         DP_OP_424J2_126_3477_n451, DP_OP_424J2_126_3477_n450,
         DP_OP_424J2_126_3477_n449, DP_OP_424J2_126_3477_n448,
         DP_OP_424J2_126_3477_n447, DP_OP_424J2_126_3477_n446,
         DP_OP_424J2_126_3477_n445, DP_OP_424J2_126_3477_n444,
         DP_OP_424J2_126_3477_n443, DP_OP_424J2_126_3477_n442,
         DP_OP_424J2_126_3477_n441, DP_OP_424J2_126_3477_n440,
         DP_OP_424J2_126_3477_n439, DP_OP_424J2_126_3477_n438,
         DP_OP_424J2_126_3477_n437, DP_OP_424J2_126_3477_n436,
         DP_OP_424J2_126_3477_n435, DP_OP_424J2_126_3477_n434,
         DP_OP_424J2_126_3477_n433, DP_OP_424J2_126_3477_n432,
         DP_OP_424J2_126_3477_n431, DP_OP_424J2_126_3477_n430,
         DP_OP_424J2_126_3477_n429, DP_OP_424J2_126_3477_n428,
         DP_OP_424J2_126_3477_n427, DP_OP_424J2_126_3477_n426,
         DP_OP_424J2_126_3477_n425, DP_OP_424J2_126_3477_n424,
         DP_OP_424J2_126_3477_n423, DP_OP_424J2_126_3477_n422,
         DP_OP_424J2_126_3477_n421, DP_OP_424J2_126_3477_n420,
         DP_OP_424J2_126_3477_n419, DP_OP_424J2_126_3477_n418,
         DP_OP_424J2_126_3477_n417, DP_OP_424J2_126_3477_n416,
         DP_OP_424J2_126_3477_n415, DP_OP_424J2_126_3477_n414,
         DP_OP_424J2_126_3477_n413, DP_OP_424J2_126_3477_n412,
         DP_OP_424J2_126_3477_n411, DP_OP_424J2_126_3477_n410,
         DP_OP_424J2_126_3477_n409, DP_OP_424J2_126_3477_n408,
         DP_OP_424J2_126_3477_n407, DP_OP_424J2_126_3477_n406,
         DP_OP_424J2_126_3477_n405, DP_OP_424J2_126_3477_n404,
         DP_OP_424J2_126_3477_n403, DP_OP_424J2_126_3477_n402,
         DP_OP_424J2_126_3477_n401, DP_OP_424J2_126_3477_n400,
         DP_OP_424J2_126_3477_n399, DP_OP_424J2_126_3477_n398,
         DP_OP_424J2_126_3477_n397, DP_OP_424J2_126_3477_n396,
         DP_OP_424J2_126_3477_n395, DP_OP_424J2_126_3477_n394,
         DP_OP_424J2_126_3477_n393, DP_OP_424J2_126_3477_n392,
         DP_OP_424J2_126_3477_n391, DP_OP_424J2_126_3477_n390,
         DP_OP_424J2_126_3477_n389, DP_OP_424J2_126_3477_n388,
         DP_OP_424J2_126_3477_n387, DP_OP_424J2_126_3477_n386,
         DP_OP_424J2_126_3477_n385, DP_OP_424J2_126_3477_n384,
         DP_OP_424J2_126_3477_n383, DP_OP_424J2_126_3477_n382,
         DP_OP_424J2_126_3477_n381, DP_OP_424J2_126_3477_n380,
         DP_OP_424J2_126_3477_n379, DP_OP_424J2_126_3477_n378,
         DP_OP_424J2_126_3477_n377, DP_OP_424J2_126_3477_n376,
         DP_OP_424J2_126_3477_n375, DP_OP_424J2_126_3477_n374,
         DP_OP_424J2_126_3477_n373, DP_OP_424J2_126_3477_n372,
         DP_OP_424J2_126_3477_n371, DP_OP_424J2_126_3477_n370,
         DP_OP_424J2_126_3477_n369, DP_OP_424J2_126_3477_n368,
         DP_OP_424J2_126_3477_n367, DP_OP_424J2_126_3477_n366,
         DP_OP_424J2_126_3477_n365, DP_OP_424J2_126_3477_n364,
         DP_OP_424J2_126_3477_n363, DP_OP_424J2_126_3477_n362,
         DP_OP_424J2_126_3477_n361, DP_OP_424J2_126_3477_n360,
         DP_OP_424J2_126_3477_n359, DP_OP_424J2_126_3477_n358,
         DP_OP_424J2_126_3477_n357, DP_OP_424J2_126_3477_n356,
         DP_OP_424J2_126_3477_n355, DP_OP_424J2_126_3477_n354,
         DP_OP_424J2_126_3477_n353, DP_OP_424J2_126_3477_n352,
         DP_OP_424J2_126_3477_n351, DP_OP_424J2_126_3477_n350,
         DP_OP_424J2_126_3477_n349, DP_OP_424J2_126_3477_n348,
         DP_OP_424J2_126_3477_n347, DP_OP_424J2_126_3477_n346,
         DP_OP_424J2_126_3477_n345, DP_OP_424J2_126_3477_n344,
         DP_OP_424J2_126_3477_n343, DP_OP_424J2_126_3477_n342,
         DP_OP_424J2_126_3477_n341, DP_OP_424J2_126_3477_n340,
         DP_OP_424J2_126_3477_n339, DP_OP_424J2_126_3477_n338,
         DP_OP_424J2_126_3477_n337, DP_OP_424J2_126_3477_n336,
         DP_OP_424J2_126_3477_n335, DP_OP_424J2_126_3477_n334,
         DP_OP_424J2_126_3477_n333, DP_OP_424J2_126_3477_n332,
         DP_OP_424J2_126_3477_n331, DP_OP_424J2_126_3477_n330,
         DP_OP_424J2_126_3477_n329, DP_OP_424J2_126_3477_n328,
         DP_OP_424J2_126_3477_n327, DP_OP_424J2_126_3477_n326,
         DP_OP_424J2_126_3477_n325, DP_OP_424J2_126_3477_n324,
         DP_OP_424J2_126_3477_n323, DP_OP_424J2_126_3477_n322,
         DP_OP_424J2_126_3477_n321, DP_OP_424J2_126_3477_n320,
         DP_OP_424J2_126_3477_n319, DP_OP_424J2_126_3477_n318,
         DP_OP_424J2_126_3477_n317, DP_OP_424J2_126_3477_n316,
         DP_OP_424J2_126_3477_n315, DP_OP_424J2_126_3477_n314,
         DP_OP_424J2_126_3477_n313, DP_OP_424J2_126_3477_n312,
         DP_OP_424J2_126_3477_n311, DP_OP_424J2_126_3477_n310,
         DP_OP_424J2_126_3477_n309, DP_OP_424J2_126_3477_n308,
         DP_OP_424J2_126_3477_n307, DP_OP_424J2_126_3477_n306,
         DP_OP_424J2_126_3477_n305, DP_OP_424J2_126_3477_n304,
         DP_OP_424J2_126_3477_n303, DP_OP_424J2_126_3477_n302,
         DP_OP_424J2_126_3477_n301, DP_OP_424J2_126_3477_n300,
         DP_OP_424J2_126_3477_n299, DP_OP_424J2_126_3477_n298,
         DP_OP_424J2_126_3477_n297, DP_OP_424J2_126_3477_n296,
         DP_OP_424J2_126_3477_n295, DP_OP_424J2_126_3477_n294,
         DP_OP_424J2_126_3477_n293, DP_OP_424J2_126_3477_n292,
         DP_OP_424J2_126_3477_n291, DP_OP_424J2_126_3477_n290,
         DP_OP_424J2_126_3477_n289, DP_OP_424J2_126_3477_n288,
         DP_OP_424J2_126_3477_n287, DP_OP_424J2_126_3477_n286,
         DP_OP_424J2_126_3477_n285, DP_OP_424J2_126_3477_n284,
         DP_OP_424J2_126_3477_n283, DP_OP_424J2_126_3477_n282,
         DP_OP_424J2_126_3477_n281, DP_OP_424J2_126_3477_n280,
         DP_OP_424J2_126_3477_n279, DP_OP_424J2_126_3477_n278,
         DP_OP_424J2_126_3477_n277, DP_OP_424J2_126_3477_n276,
         DP_OP_424J2_126_3477_n275, DP_OP_424J2_126_3477_n274,
         DP_OP_424J2_126_3477_n273, DP_OP_424J2_126_3477_n272,
         DP_OP_424J2_126_3477_n271, DP_OP_424J2_126_3477_n270,
         DP_OP_424J2_126_3477_n269, DP_OP_424J2_126_3477_n268,
         DP_OP_424J2_126_3477_n267, DP_OP_424J2_126_3477_n266,
         DP_OP_424J2_126_3477_n265, DP_OP_424J2_126_3477_n264,
         DP_OP_424J2_126_3477_n263, DP_OP_424J2_126_3477_n262,
         DP_OP_424J2_126_3477_n261, DP_OP_424J2_126_3477_n260,
         DP_OP_424J2_126_3477_n259, DP_OP_424J2_126_3477_n258,
         DP_OP_424J2_126_3477_n257, DP_OP_424J2_126_3477_n256,
         DP_OP_424J2_126_3477_n255, DP_OP_424J2_126_3477_n254,
         DP_OP_424J2_126_3477_n253, DP_OP_424J2_126_3477_n252,
         DP_OP_424J2_126_3477_n241, DP_OP_424J2_126_3477_n240,
         DP_OP_424J2_126_3477_n237, DP_OP_424J2_126_3477_n236,
         DP_OP_424J2_126_3477_n233, DP_OP_424J2_126_3477_n231,
         DP_OP_424J2_126_3477_n229, DP_OP_424J2_126_3477_n227,
         DP_OP_424J2_126_3477_n219, DP_OP_424J2_126_3477_n218,
         DP_OP_424J2_126_3477_n217, DP_OP_424J2_126_3477_n216,
         DP_OP_424J2_126_3477_n215, DP_OP_424J2_126_3477_n211,
         DP_OP_424J2_126_3477_n210, DP_OP_424J2_126_3477_n209,
         DP_OP_424J2_126_3477_n208, DP_OP_424J2_126_3477_n207,
         DP_OP_424J2_126_3477_n203, DP_OP_424J2_126_3477_n202,
         DP_OP_424J2_126_3477_n201, DP_OP_424J2_126_3477_n200,
         DP_OP_424J2_126_3477_n199, DP_OP_424J2_126_3477_n195,
         DP_OP_424J2_126_3477_n194, DP_OP_424J2_126_3477_n193,
         DP_OP_424J2_126_3477_n192, DP_OP_424J2_126_3477_n191,
         DP_OP_424J2_126_3477_n190, DP_OP_424J2_126_3477_n189,
         DP_OP_424J2_126_3477_n187, DP_OP_424J2_126_3477_n186,
         DP_OP_424J2_126_3477_n185, DP_OP_424J2_126_3477_n184,
         DP_OP_424J2_126_3477_n183, DP_OP_424J2_126_3477_n182,
         DP_OP_424J2_126_3477_n181, DP_OP_424J2_126_3477_n180,
         DP_OP_424J2_126_3477_n179, DP_OP_424J2_126_3477_n177,
         DP_OP_424J2_126_3477_n176, DP_OP_424J2_126_3477_n175,
         DP_OP_424J2_126_3477_n174, DP_OP_424J2_126_3477_n173,
         DP_OP_424J2_126_3477_n172, DP_OP_424J2_126_3477_n171,
         DP_OP_424J2_126_3477_n170, DP_OP_424J2_126_3477_n168,
         DP_OP_424J2_126_3477_n167, DP_OP_424J2_126_3477_n166,
         DP_OP_424J2_126_3477_n165, DP_OP_424J2_126_3477_n164,
         DP_OP_424J2_126_3477_n163, DP_OP_424J2_126_3477_n162,
         DP_OP_424J2_126_3477_n161, DP_OP_424J2_126_3477_n158,
         DP_OP_424J2_126_3477_n152, DP_OP_424J2_126_3477_n151,
         DP_OP_424J2_126_3477_n150, DP_OP_424J2_126_3477_n149,
         DP_OP_424J2_126_3477_n148, DP_OP_424J2_126_3477_n145,
         DP_OP_424J2_126_3477_n144, DP_OP_424J2_126_3477_n143,
         DP_OP_424J2_126_3477_n142, DP_OP_424J2_126_3477_n141,
         DP_OP_424J2_126_3477_n140, DP_OP_424J2_126_3477_n137,
         DP_OP_424J2_126_3477_n136, DP_OP_424J2_126_3477_n135,
         DP_OP_424J2_126_3477_n133, DP_OP_424J2_126_3477_n132,
         DP_OP_424J2_126_3477_n130, DP_OP_424J2_126_3477_n129,
         DP_OP_424J2_126_3477_n128, DP_OP_424J2_126_3477_n127,
         DP_OP_424J2_126_3477_n126, DP_OP_424J2_126_3477_n125,
         DP_OP_424J2_126_3477_n123, DP_OP_424J2_126_3477_n119,
         DP_OP_424J2_126_3477_n118, DP_OP_424J2_126_3477_n116,
         DP_OP_424J2_126_3477_n115, DP_OP_424J2_126_3477_n114,
         DP_OP_424J2_126_3477_n113, DP_OP_424J2_126_3477_n112,
         DP_OP_424J2_126_3477_n111, DP_OP_424J2_126_3477_n109,
         DP_OP_424J2_126_3477_n105, DP_OP_424J2_126_3477_n104,
         DP_OP_424J2_126_3477_n102, DP_OP_424J2_126_3477_n101,
         DP_OP_424J2_126_3477_n100, DP_OP_424J2_126_3477_n99,
         DP_OP_424J2_126_3477_n98, DP_OP_424J2_126_3477_n97,
         DP_OP_424J2_126_3477_n95, DP_OP_424J2_126_3477_n91,
         DP_OP_424J2_126_3477_n90, DP_OP_424J2_126_3477_n88,
         DP_OP_424J2_126_3477_n87, DP_OP_424J2_126_3477_n86,
         DP_OP_424J2_126_3477_n85, DP_OP_424J2_126_3477_n84,
         DP_OP_424J2_126_3477_n83, DP_OP_424J2_126_3477_n81,
         DP_OP_424J2_126_3477_n76, DP_OP_424J2_126_3477_n75,
         DP_OP_424J2_126_3477_n74, DP_OP_424J2_126_3477_n73,
         DP_OP_424J2_126_3477_n72, DP_OP_424J2_126_3477_n70,
         DP_OP_424J2_126_3477_n65, DP_OP_424J2_126_3477_n63,
         DP_OP_424J2_126_3477_n62, DP_OP_424J2_126_3477_n61,
         DP_OP_424J2_126_3477_n59, DP_OP_424J2_126_3477_n58,
         DP_OP_424J2_126_3477_n57, DP_OP_424J2_126_3477_n56,
         DP_OP_424J2_126_3477_n55, DP_OP_424J2_126_3477_n52,
         DP_OP_424J2_126_3477_n48, DP_OP_424J2_126_3477_n47,
         DP_OP_424J2_126_3477_n45, DP_OP_424J2_126_3477_n44,
         DP_OP_424J2_126_3477_n43, DP_OP_424J2_126_3477_n42,
         DP_OP_424J2_126_3477_n41, DP_OP_424J2_126_3477_n40,
         DP_OP_424J2_126_3477_n39, DP_OP_424J2_126_3477_n37,
         DP_OP_424J2_126_3477_n26, DP_OP_424J2_126_3477_n25,
         DP_OP_424J2_126_3477_n22, DP_OP_424J2_126_3477_n21,
         DP_OP_424J2_126_3477_n4, DP_OP_424J2_126_3477_n3,
         DP_OP_424J2_126_3477_n2, DP_OP_423J2_125_3477_n3017,
         DP_OP_423J2_125_3477_n3016, DP_OP_423J2_125_3477_n3014,
         DP_OP_423J2_125_3477_n3012, DP_OP_423J2_125_3477_n3011,
         DP_OP_423J2_125_3477_n3010, DP_OP_423J2_125_3477_n3009,
         DP_OP_423J2_125_3477_n3008, DP_OP_423J2_125_3477_n3007,
         DP_OP_423J2_125_3477_n3006, DP_OP_423J2_125_3477_n3005,
         DP_OP_423J2_125_3477_n3004, DP_OP_423J2_125_3477_n3003,
         DP_OP_423J2_125_3477_n3002, DP_OP_423J2_125_3477_n3001,
         DP_OP_423J2_125_3477_n3000, DP_OP_423J2_125_3477_n2999,
         DP_OP_423J2_125_3477_n2998, DP_OP_423J2_125_3477_n2997,
         DP_OP_423J2_125_3477_n2996, DP_OP_423J2_125_3477_n2995,
         DP_OP_423J2_125_3477_n2994, DP_OP_423J2_125_3477_n2993,
         DP_OP_423J2_125_3477_n2992, DP_OP_423J2_125_3477_n2991,
         DP_OP_423J2_125_3477_n2990, DP_OP_423J2_125_3477_n2989,
         DP_OP_423J2_125_3477_n2988, DP_OP_423J2_125_3477_n2987,
         DP_OP_423J2_125_3477_n2986, DP_OP_423J2_125_3477_n2985,
         DP_OP_423J2_125_3477_n2984, DP_OP_423J2_125_3477_n2983,
         DP_OP_423J2_125_3477_n2982, DP_OP_423J2_125_3477_n2981,
         DP_OP_423J2_125_3477_n2980, DP_OP_423J2_125_3477_n2979,
         DP_OP_423J2_125_3477_n2978, DP_OP_423J2_125_3477_n2977,
         DP_OP_423J2_125_3477_n2976, DP_OP_423J2_125_3477_n2974,
         DP_OP_423J2_125_3477_n2973, DP_OP_423J2_125_3477_n2972,
         DP_OP_423J2_125_3477_n2971, DP_OP_423J2_125_3477_n2970,
         DP_OP_423J2_125_3477_n2969, DP_OP_423J2_125_3477_n2967,
         DP_OP_423J2_125_3477_n2964, DP_OP_423J2_125_3477_n2963,
         DP_OP_423J2_125_3477_n2962, DP_OP_423J2_125_3477_n2961,
         DP_OP_423J2_125_3477_n2960, DP_OP_423J2_125_3477_n2959,
         DP_OP_423J2_125_3477_n2958, DP_OP_423J2_125_3477_n2957,
         DP_OP_423J2_125_3477_n2956, DP_OP_423J2_125_3477_n2955,
         DP_OP_423J2_125_3477_n2954, DP_OP_423J2_125_3477_n2953,
         DP_OP_423J2_125_3477_n2952, DP_OP_423J2_125_3477_n2951,
         DP_OP_423J2_125_3477_n2950, DP_OP_423J2_125_3477_n2949,
         DP_OP_423J2_125_3477_n2948, DP_OP_423J2_125_3477_n2947,
         DP_OP_423J2_125_3477_n2946, DP_OP_423J2_125_3477_n2945,
         DP_OP_423J2_125_3477_n2944, DP_OP_423J2_125_3477_n2943,
         DP_OP_423J2_125_3477_n2942, DP_OP_423J2_125_3477_n2941,
         DP_OP_423J2_125_3477_n2940, DP_OP_423J2_125_3477_n2939,
         DP_OP_423J2_125_3477_n2938, DP_OP_423J2_125_3477_n2937,
         DP_OP_423J2_125_3477_n2936, DP_OP_423J2_125_3477_n2935,
         DP_OP_423J2_125_3477_n2934, DP_OP_423J2_125_3477_n2933,
         DP_OP_423J2_125_3477_n2932, DP_OP_423J2_125_3477_n2931,
         DP_OP_423J2_125_3477_n2930, DP_OP_423J2_125_3477_n2929,
         DP_OP_423J2_125_3477_n2928, DP_OP_423J2_125_3477_n2927,
         DP_OP_423J2_125_3477_n2926, DP_OP_423J2_125_3477_n2924,
         DP_OP_423J2_125_3477_n2923, DP_OP_423J2_125_3477_n2922,
         DP_OP_423J2_125_3477_n2921, DP_OP_423J2_125_3477_n2920,
         DP_OP_423J2_125_3477_n2919, DP_OP_423J2_125_3477_n2918,
         DP_OP_423J2_125_3477_n2917, DP_OP_423J2_125_3477_n2916,
         DP_OP_423J2_125_3477_n2915, DP_OP_423J2_125_3477_n2914,
         DP_OP_423J2_125_3477_n2913, DP_OP_423J2_125_3477_n2912,
         DP_OP_423J2_125_3477_n2911, DP_OP_423J2_125_3477_n2910,
         DP_OP_423J2_125_3477_n2909, DP_OP_423J2_125_3477_n2908,
         DP_OP_423J2_125_3477_n2907, DP_OP_423J2_125_3477_n2906,
         DP_OP_423J2_125_3477_n2905, DP_OP_423J2_125_3477_n2904,
         DP_OP_423J2_125_3477_n2903, DP_OP_423J2_125_3477_n2902,
         DP_OP_423J2_125_3477_n2901, DP_OP_423J2_125_3477_n2900,
         DP_OP_423J2_125_3477_n2899, DP_OP_423J2_125_3477_n2898,
         DP_OP_423J2_125_3477_n2897, DP_OP_423J2_125_3477_n2896,
         DP_OP_423J2_125_3477_n2895, DP_OP_423J2_125_3477_n2894,
         DP_OP_423J2_125_3477_n2893, DP_OP_423J2_125_3477_n2892,
         DP_OP_423J2_125_3477_n2891, DP_OP_423J2_125_3477_n2890,
         DP_OP_423J2_125_3477_n2889, DP_OP_423J2_125_3477_n2888,
         DP_OP_423J2_125_3477_n2886, DP_OP_423J2_125_3477_n2885,
         DP_OP_423J2_125_3477_n2884, DP_OP_423J2_125_3477_n2880,
         DP_OP_423J2_125_3477_n2878, DP_OP_423J2_125_3477_n2877,
         DP_OP_423J2_125_3477_n2875, DP_OP_423J2_125_3477_n2874,
         DP_OP_423J2_125_3477_n2873, DP_OP_423J2_125_3477_n2872,
         DP_OP_423J2_125_3477_n2871, DP_OP_423J2_125_3477_n2870,
         DP_OP_423J2_125_3477_n2869, DP_OP_423J2_125_3477_n2868,
         DP_OP_423J2_125_3477_n2867, DP_OP_423J2_125_3477_n2866,
         DP_OP_423J2_125_3477_n2865, DP_OP_423J2_125_3477_n2864,
         DP_OP_423J2_125_3477_n2863, DP_OP_423J2_125_3477_n2862,
         DP_OP_423J2_125_3477_n2861, DP_OP_423J2_125_3477_n2860,
         DP_OP_423J2_125_3477_n2859, DP_OP_423J2_125_3477_n2858,
         DP_OP_423J2_125_3477_n2857, DP_OP_423J2_125_3477_n2856,
         DP_OP_423J2_125_3477_n2855, DP_OP_423J2_125_3477_n2854,
         DP_OP_423J2_125_3477_n2853, DP_OP_423J2_125_3477_n2852,
         DP_OP_423J2_125_3477_n2851, DP_OP_423J2_125_3477_n2850,
         DP_OP_423J2_125_3477_n2849, DP_OP_423J2_125_3477_n2848,
         DP_OP_423J2_125_3477_n2847, DP_OP_423J2_125_3477_n2846,
         DP_OP_423J2_125_3477_n2845, DP_OP_423J2_125_3477_n2844,
         DP_OP_423J2_125_3477_n2843, DP_OP_423J2_125_3477_n2842,
         DP_OP_423J2_125_3477_n2841, DP_OP_423J2_125_3477_n2840,
         DP_OP_423J2_125_3477_n2837, DP_OP_423J2_125_3477_n2834,
         DP_OP_423J2_125_3477_n2831, DP_OP_423J2_125_3477_n2830,
         DP_OP_423J2_125_3477_n2829, DP_OP_423J2_125_3477_n2828,
         DP_OP_423J2_125_3477_n2827, DP_OP_423J2_125_3477_n2826,
         DP_OP_423J2_125_3477_n2825, DP_OP_423J2_125_3477_n2824,
         DP_OP_423J2_125_3477_n2823, DP_OP_423J2_125_3477_n2822,
         DP_OP_423J2_125_3477_n2821, DP_OP_423J2_125_3477_n2820,
         DP_OP_423J2_125_3477_n2819, DP_OP_423J2_125_3477_n2818,
         DP_OP_423J2_125_3477_n2817, DP_OP_423J2_125_3477_n2816,
         DP_OP_423J2_125_3477_n2815, DP_OP_423J2_125_3477_n2814,
         DP_OP_423J2_125_3477_n2813, DP_OP_423J2_125_3477_n2812,
         DP_OP_423J2_125_3477_n2811, DP_OP_423J2_125_3477_n2810,
         DP_OP_423J2_125_3477_n2809, DP_OP_423J2_125_3477_n2808,
         DP_OP_423J2_125_3477_n2807, DP_OP_423J2_125_3477_n2806,
         DP_OP_423J2_125_3477_n2805, DP_OP_423J2_125_3477_n2804,
         DP_OP_423J2_125_3477_n2803, DP_OP_423J2_125_3477_n2802,
         DP_OP_423J2_125_3477_n2801, DP_OP_423J2_125_3477_n2800,
         DP_OP_423J2_125_3477_n2798, DP_OP_423J2_125_3477_n2796,
         DP_OP_423J2_125_3477_n2795, DP_OP_423J2_125_3477_n2794,
         DP_OP_423J2_125_3477_n2793, DP_OP_423J2_125_3477_n2791,
         DP_OP_423J2_125_3477_n2790, DP_OP_423J2_125_3477_n2787,
         DP_OP_423J2_125_3477_n2786, DP_OP_423J2_125_3477_n2785,
         DP_OP_423J2_125_3477_n2784, DP_OP_423J2_125_3477_n2783,
         DP_OP_423J2_125_3477_n2782, DP_OP_423J2_125_3477_n2781,
         DP_OP_423J2_125_3477_n2780, DP_OP_423J2_125_3477_n2779,
         DP_OP_423J2_125_3477_n2778, DP_OP_423J2_125_3477_n2777,
         DP_OP_423J2_125_3477_n2776, DP_OP_423J2_125_3477_n2775,
         DP_OP_423J2_125_3477_n2774, DP_OP_423J2_125_3477_n2773,
         DP_OP_423J2_125_3477_n2772, DP_OP_423J2_125_3477_n2771,
         DP_OP_423J2_125_3477_n2770, DP_OP_423J2_125_3477_n2769,
         DP_OP_423J2_125_3477_n2768, DP_OP_423J2_125_3477_n2767,
         DP_OP_423J2_125_3477_n2766, DP_OP_423J2_125_3477_n2765,
         DP_OP_423J2_125_3477_n2764, DP_OP_423J2_125_3477_n2763,
         DP_OP_423J2_125_3477_n2762, DP_OP_423J2_125_3477_n2761,
         DP_OP_423J2_125_3477_n2760, DP_OP_423J2_125_3477_n2759,
         DP_OP_423J2_125_3477_n2758, DP_OP_423J2_125_3477_n2757,
         DP_OP_423J2_125_3477_n2756, DP_OP_423J2_125_3477_n2755,
         DP_OP_423J2_125_3477_n2754, DP_OP_423J2_125_3477_n2753,
         DP_OP_423J2_125_3477_n2752, DP_OP_423J2_125_3477_n2750,
         DP_OP_423J2_125_3477_n2749, DP_OP_423J2_125_3477_n2748,
         DP_OP_423J2_125_3477_n2747, DP_OP_423J2_125_3477_n2746,
         DP_OP_423J2_125_3477_n2745, DP_OP_423J2_125_3477_n2743,
         DP_OP_423J2_125_3477_n2742, DP_OP_423J2_125_3477_n2741,
         DP_OP_423J2_125_3477_n2740, DP_OP_423J2_125_3477_n2739,
         DP_OP_423J2_125_3477_n2738, DP_OP_423J2_125_3477_n2737,
         DP_OP_423J2_125_3477_n2736, DP_OP_423J2_125_3477_n2735,
         DP_OP_423J2_125_3477_n2734, DP_OP_423J2_125_3477_n2733,
         DP_OP_423J2_125_3477_n2732, DP_OP_423J2_125_3477_n2731,
         DP_OP_423J2_125_3477_n2730, DP_OP_423J2_125_3477_n2729,
         DP_OP_423J2_125_3477_n2728, DP_OP_423J2_125_3477_n2727,
         DP_OP_423J2_125_3477_n2726, DP_OP_423J2_125_3477_n2725,
         DP_OP_423J2_125_3477_n2724, DP_OP_423J2_125_3477_n2723,
         DP_OP_423J2_125_3477_n2722, DP_OP_423J2_125_3477_n2721,
         DP_OP_423J2_125_3477_n2720, DP_OP_423J2_125_3477_n2719,
         DP_OP_423J2_125_3477_n2718, DP_OP_423J2_125_3477_n2717,
         DP_OP_423J2_125_3477_n2716, DP_OP_423J2_125_3477_n2715,
         DP_OP_423J2_125_3477_n2714, DP_OP_423J2_125_3477_n2713,
         DP_OP_423J2_125_3477_n2712, DP_OP_423J2_125_3477_n2710,
         DP_OP_423J2_125_3477_n2709, DP_OP_423J2_125_3477_n2708,
         DP_OP_423J2_125_3477_n2707, DP_OP_423J2_125_3477_n2705,
         DP_OP_423J2_125_3477_n2702, DP_OP_423J2_125_3477_n2700,
         DP_OP_423J2_125_3477_n2699, DP_OP_423J2_125_3477_n2698,
         DP_OP_423J2_125_3477_n2697, DP_OP_423J2_125_3477_n2696,
         DP_OP_423J2_125_3477_n2695, DP_OP_423J2_125_3477_n2694,
         DP_OP_423J2_125_3477_n2693, DP_OP_423J2_125_3477_n2692,
         DP_OP_423J2_125_3477_n2691, DP_OP_423J2_125_3477_n2690,
         DP_OP_423J2_125_3477_n2689, DP_OP_423J2_125_3477_n2688,
         DP_OP_423J2_125_3477_n2687, DP_OP_423J2_125_3477_n2686,
         DP_OP_423J2_125_3477_n2685, DP_OP_423J2_125_3477_n2684,
         DP_OP_423J2_125_3477_n2683, DP_OP_423J2_125_3477_n2682,
         DP_OP_423J2_125_3477_n2681, DP_OP_423J2_125_3477_n2680,
         DP_OP_423J2_125_3477_n2679, DP_OP_423J2_125_3477_n2678,
         DP_OP_423J2_125_3477_n2677, DP_OP_423J2_125_3477_n2676,
         DP_OP_423J2_125_3477_n2675, DP_OP_423J2_125_3477_n2674,
         DP_OP_423J2_125_3477_n2673, DP_OP_423J2_125_3477_n2672,
         DP_OP_423J2_125_3477_n2671, DP_OP_423J2_125_3477_n2670,
         DP_OP_423J2_125_3477_n2669, DP_OP_423J2_125_3477_n2668,
         DP_OP_423J2_125_3477_n2667, DP_OP_423J2_125_3477_n2665,
         DP_OP_423J2_125_3477_n2664, DP_OP_423J2_125_3477_n2663,
         DP_OP_423J2_125_3477_n2662, DP_OP_423J2_125_3477_n2659,
         DP_OP_423J2_125_3477_n2658, DP_OP_423J2_125_3477_n2656,
         DP_OP_423J2_125_3477_n2655, DP_OP_423J2_125_3477_n2654,
         DP_OP_423J2_125_3477_n2653, DP_OP_423J2_125_3477_n2652,
         DP_OP_423J2_125_3477_n2651, DP_OP_423J2_125_3477_n2650,
         DP_OP_423J2_125_3477_n2649, DP_OP_423J2_125_3477_n2648,
         DP_OP_423J2_125_3477_n2647, DP_OP_423J2_125_3477_n2646,
         DP_OP_423J2_125_3477_n2645, DP_OP_423J2_125_3477_n2644,
         DP_OP_423J2_125_3477_n2643, DP_OP_423J2_125_3477_n2642,
         DP_OP_423J2_125_3477_n2641, DP_OP_423J2_125_3477_n2640,
         DP_OP_423J2_125_3477_n2639, DP_OP_423J2_125_3477_n2638,
         DP_OP_423J2_125_3477_n2637, DP_OP_423J2_125_3477_n2636,
         DP_OP_423J2_125_3477_n2635, DP_OP_423J2_125_3477_n2634,
         DP_OP_423J2_125_3477_n2633, DP_OP_423J2_125_3477_n2632,
         DP_OP_423J2_125_3477_n2631, DP_OP_423J2_125_3477_n2630,
         DP_OP_423J2_125_3477_n2629, DP_OP_423J2_125_3477_n2628,
         DP_OP_423J2_125_3477_n2627, DP_OP_423J2_125_3477_n2626,
         DP_OP_423J2_125_3477_n2625, DP_OP_423J2_125_3477_n2624,
         DP_OP_423J2_125_3477_n2623, DP_OP_423J2_125_3477_n2621,
         DP_OP_423J2_125_3477_n2619, DP_OP_423J2_125_3477_n2617,
         DP_OP_423J2_125_3477_n2613, DP_OP_423J2_125_3477_n2612,
         DP_OP_423J2_125_3477_n2611, DP_OP_423J2_125_3477_n2610,
         DP_OP_423J2_125_3477_n2609, DP_OP_423J2_125_3477_n2608,
         DP_OP_423J2_125_3477_n2607, DP_OP_423J2_125_3477_n2606,
         DP_OP_423J2_125_3477_n2605, DP_OP_423J2_125_3477_n2604,
         DP_OP_423J2_125_3477_n2603, DP_OP_423J2_125_3477_n2602,
         DP_OP_423J2_125_3477_n2601, DP_OP_423J2_125_3477_n2600,
         DP_OP_423J2_125_3477_n2599, DP_OP_423J2_125_3477_n2598,
         DP_OP_423J2_125_3477_n2597, DP_OP_423J2_125_3477_n2596,
         DP_OP_423J2_125_3477_n2595, DP_OP_423J2_125_3477_n2594,
         DP_OP_423J2_125_3477_n2593, DP_OP_423J2_125_3477_n2592,
         DP_OP_423J2_125_3477_n2591, DP_OP_423J2_125_3477_n2590,
         DP_OP_423J2_125_3477_n2589, DP_OP_423J2_125_3477_n2588,
         DP_OP_423J2_125_3477_n2587, DP_OP_423J2_125_3477_n2586,
         DP_OP_423J2_125_3477_n2585, DP_OP_423J2_125_3477_n2584,
         DP_OP_423J2_125_3477_n2583, DP_OP_423J2_125_3477_n2582,
         DP_OP_423J2_125_3477_n2581, DP_OP_423J2_125_3477_n2580,
         DP_OP_423J2_125_3477_n2579, DP_OP_423J2_125_3477_n2577,
         DP_OP_423J2_125_3477_n2576, DP_OP_423J2_125_3477_n2575,
         DP_OP_423J2_125_3477_n2574, DP_OP_423J2_125_3477_n2573,
         DP_OP_423J2_125_3477_n2572, DP_OP_423J2_125_3477_n2571,
         DP_OP_423J2_125_3477_n2570, DP_OP_423J2_125_3477_n2569,
         DP_OP_423J2_125_3477_n2568, DP_OP_423J2_125_3477_n2567,
         DP_OP_423J2_125_3477_n2566, DP_OP_423J2_125_3477_n2565,
         DP_OP_423J2_125_3477_n2564, DP_OP_423J2_125_3477_n2563,
         DP_OP_423J2_125_3477_n2562, DP_OP_423J2_125_3477_n2561,
         DP_OP_423J2_125_3477_n2560, DP_OP_423J2_125_3477_n2559,
         DP_OP_423J2_125_3477_n2558, DP_OP_423J2_125_3477_n2557,
         DP_OP_423J2_125_3477_n2556, DP_OP_423J2_125_3477_n2555,
         DP_OP_423J2_125_3477_n2554, DP_OP_423J2_125_3477_n2553,
         DP_OP_423J2_125_3477_n2552, DP_OP_423J2_125_3477_n2551,
         DP_OP_423J2_125_3477_n2550, DP_OP_423J2_125_3477_n2549,
         DP_OP_423J2_125_3477_n2548, DP_OP_423J2_125_3477_n2547,
         DP_OP_423J2_125_3477_n2546, DP_OP_423J2_125_3477_n2545,
         DP_OP_423J2_125_3477_n2544, DP_OP_423J2_125_3477_n2543,
         DP_OP_423J2_125_3477_n2542, DP_OP_423J2_125_3477_n2541,
         DP_OP_423J2_125_3477_n2540, DP_OP_423J2_125_3477_n2539,
         DP_OP_423J2_125_3477_n2538, DP_OP_423J2_125_3477_n2537,
         DP_OP_423J2_125_3477_n2536, DP_OP_423J2_125_3477_n2535,
         DP_OP_423J2_125_3477_n2534, DP_OP_423J2_125_3477_n2533,
         DP_OP_423J2_125_3477_n2532, DP_OP_423J2_125_3477_n2531,
         DP_OP_423J2_125_3477_n2530, DP_OP_423J2_125_3477_n2529,
         DP_OP_423J2_125_3477_n2528, DP_OP_423J2_125_3477_n2527,
         DP_OP_423J2_125_3477_n2526, DP_OP_423J2_125_3477_n2525,
         DP_OP_423J2_125_3477_n2523, DP_OP_423J2_125_3477_n2522,
         DP_OP_423J2_125_3477_n2521, DP_OP_423J2_125_3477_n2520,
         DP_OP_423J2_125_3477_n2519, DP_OP_423J2_125_3477_n2518,
         DP_OP_423J2_125_3477_n2517, DP_OP_423J2_125_3477_n2516,
         DP_OP_423J2_125_3477_n2515, DP_OP_423J2_125_3477_n2514,
         DP_OP_423J2_125_3477_n2513, DP_OP_423J2_125_3477_n2512,
         DP_OP_423J2_125_3477_n2511, DP_OP_423J2_125_3477_n2510,
         DP_OP_423J2_125_3477_n2509, DP_OP_423J2_125_3477_n2508,
         DP_OP_423J2_125_3477_n2507, DP_OP_423J2_125_3477_n2506,
         DP_OP_423J2_125_3477_n2505, DP_OP_423J2_125_3477_n2504,
         DP_OP_423J2_125_3477_n2503, DP_OP_423J2_125_3477_n2502,
         DP_OP_423J2_125_3477_n2501, DP_OP_423J2_125_3477_n2500,
         DP_OP_423J2_125_3477_n2499, DP_OP_423J2_125_3477_n2498,
         DP_OP_423J2_125_3477_n2497, DP_OP_423J2_125_3477_n2496,
         DP_OP_423J2_125_3477_n2495, DP_OP_423J2_125_3477_n2494,
         DP_OP_423J2_125_3477_n2493, DP_OP_423J2_125_3477_n2492,
         DP_OP_423J2_125_3477_n2491, DP_OP_423J2_125_3477_n2490,
         DP_OP_423J2_125_3477_n2489, DP_OP_423J2_125_3477_n2488,
         DP_OP_423J2_125_3477_n2487, DP_OP_423J2_125_3477_n2484,
         DP_OP_423J2_125_3477_n2482, DP_OP_423J2_125_3477_n2481,
         DP_OP_423J2_125_3477_n2479, DP_OP_423J2_125_3477_n2478,
         DP_OP_423J2_125_3477_n2477, DP_OP_423J2_125_3477_n2476,
         DP_OP_423J2_125_3477_n2475, DP_OP_423J2_125_3477_n2474,
         DP_OP_423J2_125_3477_n2473, DP_OP_423J2_125_3477_n2472,
         DP_OP_423J2_125_3477_n2471, DP_OP_423J2_125_3477_n2470,
         DP_OP_423J2_125_3477_n2469, DP_OP_423J2_125_3477_n2468,
         DP_OP_423J2_125_3477_n2467, DP_OP_423J2_125_3477_n2466,
         DP_OP_423J2_125_3477_n2465, DP_OP_423J2_125_3477_n2464,
         DP_OP_423J2_125_3477_n2463, DP_OP_423J2_125_3477_n2462,
         DP_OP_423J2_125_3477_n2461, DP_OP_423J2_125_3477_n2460,
         DP_OP_423J2_125_3477_n2459, DP_OP_423J2_125_3477_n2458,
         DP_OP_423J2_125_3477_n2457, DP_OP_423J2_125_3477_n2456,
         DP_OP_423J2_125_3477_n2455, DP_OP_423J2_125_3477_n2454,
         DP_OP_423J2_125_3477_n2453, DP_OP_423J2_125_3477_n2452,
         DP_OP_423J2_125_3477_n2451, DP_OP_423J2_125_3477_n2450,
         DP_OP_423J2_125_3477_n2449, DP_OP_423J2_125_3477_n2448,
         DP_OP_423J2_125_3477_n2446, DP_OP_423J2_125_3477_n2445,
         DP_OP_423J2_125_3477_n2444, DP_OP_423J2_125_3477_n2442,
         DP_OP_423J2_125_3477_n2441, DP_OP_423J2_125_3477_n2439,
         DP_OP_423J2_125_3477_n2437, DP_OP_423J2_125_3477_n2436,
         DP_OP_423J2_125_3477_n2435, DP_OP_423J2_125_3477_n2434,
         DP_OP_423J2_125_3477_n2433, DP_OP_423J2_125_3477_n2432,
         DP_OP_423J2_125_3477_n2431, DP_OP_423J2_125_3477_n2430,
         DP_OP_423J2_125_3477_n2429, DP_OP_423J2_125_3477_n2428,
         DP_OP_423J2_125_3477_n2427, DP_OP_423J2_125_3477_n2426,
         DP_OP_423J2_125_3477_n2425, DP_OP_423J2_125_3477_n2424,
         DP_OP_423J2_125_3477_n2423, DP_OP_423J2_125_3477_n2422,
         DP_OP_423J2_125_3477_n2421, DP_OP_423J2_125_3477_n2420,
         DP_OP_423J2_125_3477_n2419, DP_OP_423J2_125_3477_n2418,
         DP_OP_423J2_125_3477_n2417, DP_OP_423J2_125_3477_n2416,
         DP_OP_423J2_125_3477_n2415, DP_OP_423J2_125_3477_n2414,
         DP_OP_423J2_125_3477_n2413, DP_OP_423J2_125_3477_n2412,
         DP_OP_423J2_125_3477_n2411, DP_OP_423J2_125_3477_n2410,
         DP_OP_423J2_125_3477_n2409, DP_OP_423J2_125_3477_n2408,
         DP_OP_423J2_125_3477_n2407, DP_OP_423J2_125_3477_n2406,
         DP_OP_423J2_125_3477_n2405, DP_OP_423J2_125_3477_n2404,
         DP_OP_423J2_125_3477_n2403, DP_OP_423J2_125_3477_n2402,
         DP_OP_423J2_125_3477_n2401, DP_OP_423J2_125_3477_n2400,
         DP_OP_423J2_125_3477_n2398, DP_OP_423J2_125_3477_n2397,
         DP_OP_423J2_125_3477_n2396, DP_OP_423J2_125_3477_n2391,
         DP_OP_423J2_125_3477_n2390, DP_OP_423J2_125_3477_n2389,
         DP_OP_423J2_125_3477_n2388, DP_OP_423J2_125_3477_n2387,
         DP_OP_423J2_125_3477_n2386, DP_OP_423J2_125_3477_n2385,
         DP_OP_423J2_125_3477_n2384, DP_OP_423J2_125_3477_n2383,
         DP_OP_423J2_125_3477_n2382, DP_OP_423J2_125_3477_n2381,
         DP_OP_423J2_125_3477_n2380, DP_OP_423J2_125_3477_n2379,
         DP_OP_423J2_125_3477_n2378, DP_OP_423J2_125_3477_n2377,
         DP_OP_423J2_125_3477_n2376, DP_OP_423J2_125_3477_n2375,
         DP_OP_423J2_125_3477_n2374, DP_OP_423J2_125_3477_n2373,
         DP_OP_423J2_125_3477_n2372, DP_OP_423J2_125_3477_n2371,
         DP_OP_423J2_125_3477_n2370, DP_OP_423J2_125_3477_n2369,
         DP_OP_423J2_125_3477_n2368, DP_OP_423J2_125_3477_n2367,
         DP_OP_423J2_125_3477_n2366, DP_OP_423J2_125_3477_n2365,
         DP_OP_423J2_125_3477_n2364, DP_OP_423J2_125_3477_n2363,
         DP_OP_423J2_125_3477_n2362, DP_OP_423J2_125_3477_n2361,
         DP_OP_423J2_125_3477_n2360, DP_OP_423J2_125_3477_n2359,
         DP_OP_423J2_125_3477_n2358, DP_OP_423J2_125_3477_n2357,
         DP_OP_423J2_125_3477_n2356, DP_OP_423J2_125_3477_n2355,
         DP_OP_423J2_125_3477_n2354, DP_OP_423J2_125_3477_n2353,
         DP_OP_423J2_125_3477_n2351, DP_OP_423J2_125_3477_n2350,
         DP_OP_423J2_125_3477_n2348, DP_OP_423J2_125_3477_n2347,
         DP_OP_423J2_125_3477_n2346, DP_OP_423J2_125_3477_n2345,
         DP_OP_423J2_125_3477_n2344, DP_OP_423J2_125_3477_n2343,
         DP_OP_423J2_125_3477_n2342, DP_OP_423J2_125_3477_n2341,
         DP_OP_423J2_125_3477_n2340, DP_OP_423J2_125_3477_n2339,
         DP_OP_423J2_125_3477_n2338, DP_OP_423J2_125_3477_n2337,
         DP_OP_423J2_125_3477_n2336, DP_OP_423J2_125_3477_n2335,
         DP_OP_423J2_125_3477_n2334, DP_OP_423J2_125_3477_n2333,
         DP_OP_423J2_125_3477_n2332, DP_OP_423J2_125_3477_n2331,
         DP_OP_423J2_125_3477_n2330, DP_OP_423J2_125_3477_n2329,
         DP_OP_423J2_125_3477_n2328, DP_OP_423J2_125_3477_n2327,
         DP_OP_423J2_125_3477_n2326, DP_OP_423J2_125_3477_n2325,
         DP_OP_423J2_125_3477_n2324, DP_OP_423J2_125_3477_n2323,
         DP_OP_423J2_125_3477_n2322, DP_OP_423J2_125_3477_n2321,
         DP_OP_423J2_125_3477_n2320, DP_OP_423J2_125_3477_n2319,
         DP_OP_423J2_125_3477_n2318, DP_OP_423J2_125_3477_n2317,
         DP_OP_423J2_125_3477_n2316, DP_OP_423J2_125_3477_n2315,
         DP_OP_423J2_125_3477_n2314, DP_OP_423J2_125_3477_n2313,
         DP_OP_423J2_125_3477_n2312, DP_OP_423J2_125_3477_n2311,
         DP_OP_423J2_125_3477_n2308, DP_OP_423J2_125_3477_n2307,
         DP_OP_423J2_125_3477_n2305, DP_OP_423J2_125_3477_n2304,
         DP_OP_423J2_125_3477_n2303, DP_OP_423J2_125_3477_n2302,
         DP_OP_423J2_125_3477_n2301, DP_OP_423J2_125_3477_n2300,
         DP_OP_423J2_125_3477_n2299, DP_OP_423J2_125_3477_n2298,
         DP_OP_423J2_125_3477_n2297, DP_OP_423J2_125_3477_n2296,
         DP_OP_423J2_125_3477_n2295, DP_OP_423J2_125_3477_n2294,
         DP_OP_423J2_125_3477_n2293, DP_OP_423J2_125_3477_n2292,
         DP_OP_423J2_125_3477_n2291, DP_OP_423J2_125_3477_n2290,
         DP_OP_423J2_125_3477_n2289, DP_OP_423J2_125_3477_n2288,
         DP_OP_423J2_125_3477_n2287, DP_OP_423J2_125_3477_n2286,
         DP_OP_423J2_125_3477_n2285, DP_OP_423J2_125_3477_n2284,
         DP_OP_423J2_125_3477_n2283, DP_OP_423J2_125_3477_n2282,
         DP_OP_423J2_125_3477_n2281, DP_OP_423J2_125_3477_n2280,
         DP_OP_423J2_125_3477_n2279, DP_OP_423J2_125_3477_n2278,
         DP_OP_423J2_125_3477_n2277, DP_OP_423J2_125_3477_n2276,
         DP_OP_423J2_125_3477_n2275, DP_OP_423J2_125_3477_n2274,
         DP_OP_423J2_125_3477_n2273, DP_OP_423J2_125_3477_n2272,
         DP_OP_423J2_125_3477_n2270, DP_OP_423J2_125_3477_n2268,
         DP_OP_423J2_125_3477_n2267, DP_OP_423J2_125_3477_n2266,
         DP_OP_423J2_125_3477_n2265, DP_OP_423J2_125_3477_n2263,
         DP_OP_423J2_125_3477_n2262, DP_OP_423J2_125_3477_n2261,
         DP_OP_423J2_125_3477_n2260, DP_OP_423J2_125_3477_n2259,
         DP_OP_423J2_125_3477_n2258, DP_OP_423J2_125_3477_n2257,
         DP_OP_423J2_125_3477_n2256, DP_OP_423J2_125_3477_n2255,
         DP_OP_423J2_125_3477_n2254, DP_OP_423J2_125_3477_n2253,
         DP_OP_423J2_125_3477_n2252, DP_OP_423J2_125_3477_n2251,
         DP_OP_423J2_125_3477_n2250, DP_OP_423J2_125_3477_n2249,
         DP_OP_423J2_125_3477_n2248, DP_OP_423J2_125_3477_n2247,
         DP_OP_423J2_125_3477_n2246, DP_OP_423J2_125_3477_n2245,
         DP_OP_423J2_125_3477_n2244, DP_OP_423J2_125_3477_n2243,
         DP_OP_423J2_125_3477_n2242, DP_OP_423J2_125_3477_n2241,
         DP_OP_423J2_125_3477_n2240, DP_OP_423J2_125_3477_n2239,
         DP_OP_423J2_125_3477_n2238, DP_OP_423J2_125_3477_n2237,
         DP_OP_423J2_125_3477_n2236, DP_OP_423J2_125_3477_n2235,
         DP_OP_423J2_125_3477_n2234, DP_OP_423J2_125_3477_n2233,
         DP_OP_423J2_125_3477_n2232, DP_OP_423J2_125_3477_n2231,
         DP_OP_423J2_125_3477_n2230, DP_OP_423J2_125_3477_n2229,
         DP_OP_423J2_125_3477_n2228, DP_OP_423J2_125_3477_n2226,
         DP_OP_423J2_125_3477_n2225, DP_OP_423J2_125_3477_n2224,
         DP_OP_423J2_125_3477_n2219, DP_OP_423J2_125_3477_n2218,
         DP_OP_423J2_125_3477_n2217, DP_OP_423J2_125_3477_n2215,
         DP_OP_423J2_125_3477_n2214, DP_OP_423J2_125_3477_n2213,
         DP_OP_423J2_125_3477_n2212, DP_OP_423J2_125_3477_n2211,
         DP_OP_423J2_125_3477_n2210, DP_OP_423J2_125_3477_n2209,
         DP_OP_423J2_125_3477_n2208, DP_OP_423J2_125_3477_n2207,
         DP_OP_423J2_125_3477_n2206, DP_OP_423J2_125_3477_n2205,
         DP_OP_423J2_125_3477_n2204, DP_OP_423J2_125_3477_n2203,
         DP_OP_423J2_125_3477_n2202, DP_OP_423J2_125_3477_n2201,
         DP_OP_423J2_125_3477_n2200, DP_OP_423J2_125_3477_n2199,
         DP_OP_423J2_125_3477_n2198, DP_OP_423J2_125_3477_n2197,
         DP_OP_423J2_125_3477_n2196, DP_OP_423J2_125_3477_n2195,
         DP_OP_423J2_125_3477_n2194, DP_OP_423J2_125_3477_n2193,
         DP_OP_423J2_125_3477_n2192, DP_OP_423J2_125_3477_n2191,
         DP_OP_423J2_125_3477_n2190, DP_OP_423J2_125_3477_n2189,
         DP_OP_423J2_125_3477_n2188, DP_OP_423J2_125_3477_n2187,
         DP_OP_423J2_125_3477_n2186, DP_OP_423J2_125_3477_n2185,
         DP_OP_423J2_125_3477_n2184, DP_OP_423J2_125_3477_n2183,
         DP_OP_423J2_125_3477_n2181, DP_OP_423J2_125_3477_n2180,
         DP_OP_423J2_125_3477_n2178, DP_OP_423J2_125_3477_n2175,
         DP_OP_423J2_125_3477_n2172, DP_OP_423J2_125_3477_n2171,
         DP_OP_423J2_125_3477_n2170, DP_OP_423J2_125_3477_n2169,
         DP_OP_423J2_125_3477_n2168, DP_OP_423J2_125_3477_n2167,
         DP_OP_423J2_125_3477_n2166, DP_OP_423J2_125_3477_n2165,
         DP_OP_423J2_125_3477_n2164, DP_OP_423J2_125_3477_n2163,
         DP_OP_423J2_125_3477_n2162, DP_OP_423J2_125_3477_n2161,
         DP_OP_423J2_125_3477_n2160, DP_OP_423J2_125_3477_n2159,
         DP_OP_423J2_125_3477_n2158, DP_OP_423J2_125_3477_n2157,
         DP_OP_423J2_125_3477_n2156, DP_OP_423J2_125_3477_n2155,
         DP_OP_423J2_125_3477_n2154, DP_OP_423J2_125_3477_n2153,
         DP_OP_423J2_125_3477_n2152, DP_OP_423J2_125_3477_n2151,
         DP_OP_423J2_125_3477_n2150, DP_OP_423J2_125_3477_n2149,
         DP_OP_423J2_125_3477_n2148, DP_OP_423J2_125_3477_n2147,
         DP_OP_423J2_125_3477_n2146, DP_OP_423J2_125_3477_n2145,
         DP_OP_423J2_125_3477_n2144, DP_OP_423J2_125_3477_n2143,
         DP_OP_423J2_125_3477_n2142, DP_OP_423J2_125_3477_n2141,
         DP_OP_423J2_125_3477_n2140, DP_OP_423J2_125_3477_n2139,
         DP_OP_423J2_125_3477_n2138, DP_OP_423J2_125_3477_n2136,
         DP_OP_423J2_125_3477_n2135, DP_OP_423J2_125_3477_n2134,
         DP_OP_423J2_125_3477_n2128, DP_OP_423J2_125_3477_n2127,
         DP_OP_423J2_125_3477_n2126, DP_OP_423J2_125_3477_n2125,
         DP_OP_423J2_125_3477_n2124, DP_OP_423J2_125_3477_n2123,
         DP_OP_423J2_125_3477_n2122, DP_OP_423J2_125_3477_n2121,
         DP_OP_423J2_125_3477_n2120, DP_OP_423J2_125_3477_n2119,
         DP_OP_423J2_125_3477_n2118, DP_OP_423J2_125_3477_n2117,
         DP_OP_423J2_125_3477_n2116, DP_OP_423J2_125_3477_n2115,
         DP_OP_423J2_125_3477_n2114, DP_OP_423J2_125_3477_n2113,
         DP_OP_423J2_125_3477_n2112, DP_OP_423J2_125_3477_n2111,
         DP_OP_423J2_125_3477_n2110, DP_OP_423J2_125_3477_n2109,
         DP_OP_423J2_125_3477_n2108, DP_OP_423J2_125_3477_n2107,
         DP_OP_423J2_125_3477_n2106, DP_OP_423J2_125_3477_n2105,
         DP_OP_423J2_125_3477_n2104, DP_OP_423J2_125_3477_n2103,
         DP_OP_423J2_125_3477_n2102, DP_OP_423J2_125_3477_n2101,
         DP_OP_423J2_125_3477_n2100, DP_OP_423J2_125_3477_n2099,
         DP_OP_423J2_125_3477_n2098, DP_OP_423J2_125_3477_n2097,
         DP_OP_423J2_125_3477_n2096, DP_OP_423J2_125_3477_n2093,
         DP_OP_423J2_125_3477_n2092, DP_OP_423J2_125_3477_n2088,
         DP_OP_423J2_125_3477_n2087, DP_OP_423J2_125_3477_n2086,
         DP_OP_423J2_125_3477_n2084, DP_OP_423J2_125_3477_n2083,
         DP_OP_423J2_125_3477_n2082, DP_OP_423J2_125_3477_n2081,
         DP_OP_423J2_125_3477_n2080, DP_OP_423J2_125_3477_n2079,
         DP_OP_423J2_125_3477_n2078, DP_OP_423J2_125_3477_n2077,
         DP_OP_423J2_125_3477_n2076, DP_OP_423J2_125_3477_n2075,
         DP_OP_423J2_125_3477_n2074, DP_OP_423J2_125_3477_n2073,
         DP_OP_423J2_125_3477_n2072, DP_OP_423J2_125_3477_n2071,
         DP_OP_423J2_125_3477_n2070, DP_OP_423J2_125_3477_n2069,
         DP_OP_423J2_125_3477_n2068, DP_OP_423J2_125_3477_n2067,
         DP_OP_423J2_125_3477_n2066, DP_OP_423J2_125_3477_n2065,
         DP_OP_423J2_125_3477_n2064, DP_OP_423J2_125_3477_n2063,
         DP_OP_423J2_125_3477_n2062, DP_OP_423J2_125_3477_n2061,
         DP_OP_423J2_125_3477_n2060, DP_OP_423J2_125_3477_n2059,
         DP_OP_423J2_125_3477_n2058, DP_OP_423J2_125_3477_n2057,
         DP_OP_423J2_125_3477_n2056, DP_OP_423J2_125_3477_n2055,
         DP_OP_423J2_125_3477_n2054, DP_OP_423J2_125_3477_n2053,
         DP_OP_423J2_125_3477_n2052, DP_OP_423J2_125_3477_n2050,
         DP_OP_423J2_125_3477_n2048, DP_OP_423J2_125_3477_n2044,
         DP_OP_423J2_125_3477_n2040, DP_OP_423J2_125_3477_n2039,
         DP_OP_423J2_125_3477_n2038, DP_OP_423J2_125_3477_n2037,
         DP_OP_423J2_125_3477_n2036, DP_OP_423J2_125_3477_n2035,
         DP_OP_423J2_125_3477_n2034, DP_OP_423J2_125_3477_n2033,
         DP_OP_423J2_125_3477_n2032, DP_OP_423J2_125_3477_n2031,
         DP_OP_423J2_125_3477_n2030, DP_OP_423J2_125_3477_n2029,
         DP_OP_423J2_125_3477_n2028, DP_OP_423J2_125_3477_n2027,
         DP_OP_423J2_125_3477_n2026, DP_OP_423J2_125_3477_n2025,
         DP_OP_423J2_125_3477_n2024, DP_OP_423J2_125_3477_n2023,
         DP_OP_423J2_125_3477_n2022, DP_OP_423J2_125_3477_n2021,
         DP_OP_423J2_125_3477_n2020, DP_OP_423J2_125_3477_n2019,
         DP_OP_423J2_125_3477_n2018, DP_OP_423J2_125_3477_n2017,
         DP_OP_423J2_125_3477_n2016, DP_OP_423J2_125_3477_n2015,
         DP_OP_423J2_125_3477_n2014, DP_OP_423J2_125_3477_n2013,
         DP_OP_423J2_125_3477_n2012, DP_OP_423J2_125_3477_n2011,
         DP_OP_423J2_125_3477_n2010, DP_OP_423J2_125_3477_n2009,
         DP_OP_423J2_125_3477_n2008, DP_OP_423J2_125_3477_n2007,
         DP_OP_423J2_125_3477_n2006, DP_OP_423J2_125_3477_n2005,
         DP_OP_423J2_125_3477_n2004, DP_OP_423J2_125_3477_n2003,
         DP_OP_423J2_125_3477_n2000, DP_OP_423J2_125_3477_n1998,
         DP_OP_423J2_125_3477_n1997, DP_OP_423J2_125_3477_n1995,
         DP_OP_423J2_125_3477_n1994, DP_OP_423J2_125_3477_n1993,
         DP_OP_423J2_125_3477_n1992, DP_OP_423J2_125_3477_n1991,
         DP_OP_423J2_125_3477_n1990, DP_OP_423J2_125_3477_n1989,
         DP_OP_423J2_125_3477_n1988, DP_OP_423J2_125_3477_n1987,
         DP_OP_423J2_125_3477_n1986, DP_OP_423J2_125_3477_n1985,
         DP_OP_423J2_125_3477_n1984, DP_OP_423J2_125_3477_n1983,
         DP_OP_423J2_125_3477_n1982, DP_OP_423J2_125_3477_n1981,
         DP_OP_423J2_125_3477_n1980, DP_OP_423J2_125_3477_n1979,
         DP_OP_423J2_125_3477_n1978, DP_OP_423J2_125_3477_n1977,
         DP_OP_423J2_125_3477_n1976, DP_OP_423J2_125_3477_n1975,
         DP_OP_423J2_125_3477_n1974, DP_OP_423J2_125_3477_n1973,
         DP_OP_423J2_125_3477_n1972, DP_OP_423J2_125_3477_n1971,
         DP_OP_423J2_125_3477_n1970, DP_OP_423J2_125_3477_n1969,
         DP_OP_423J2_125_3477_n1968, DP_OP_423J2_125_3477_n1967,
         DP_OP_423J2_125_3477_n1966, DP_OP_423J2_125_3477_n1965,
         DP_OP_423J2_125_3477_n1964, DP_OP_423J2_125_3477_n1963,
         DP_OP_423J2_125_3477_n1962, DP_OP_423J2_125_3477_n1960,
         DP_OP_423J2_125_3477_n1958, DP_OP_423J2_125_3477_n1957,
         DP_OP_423J2_125_3477_n1952, DP_OP_423J2_125_3477_n1951,
         DP_OP_423J2_125_3477_n1950, DP_OP_423J2_125_3477_n1949,
         DP_OP_423J2_125_3477_n1948, DP_OP_423J2_125_3477_n1947,
         DP_OP_423J2_125_3477_n1946, DP_OP_423J2_125_3477_n1945,
         DP_OP_423J2_125_3477_n1944, DP_OP_423J2_125_3477_n1943,
         DP_OP_423J2_125_3477_n1942, DP_OP_423J2_125_3477_n1941,
         DP_OP_423J2_125_3477_n1940, DP_OP_423J2_125_3477_n1939,
         DP_OP_423J2_125_3477_n1938, DP_OP_423J2_125_3477_n1937,
         DP_OP_423J2_125_3477_n1936, DP_OP_423J2_125_3477_n1935,
         DP_OP_423J2_125_3477_n1934, DP_OP_423J2_125_3477_n1933,
         DP_OP_423J2_125_3477_n1932, DP_OP_423J2_125_3477_n1931,
         DP_OP_423J2_125_3477_n1930, DP_OP_423J2_125_3477_n1929,
         DP_OP_423J2_125_3477_n1928, DP_OP_423J2_125_3477_n1927,
         DP_OP_423J2_125_3477_n1926, DP_OP_423J2_125_3477_n1925,
         DP_OP_423J2_125_3477_n1924, DP_OP_423J2_125_3477_n1923,
         DP_OP_423J2_125_3477_n1922, DP_OP_423J2_125_3477_n1921,
         DP_OP_423J2_125_3477_n1920, DP_OP_423J2_125_3477_n1886,
         DP_OP_423J2_125_3477_n1885, DP_OP_423J2_125_3477_n1884,
         DP_OP_423J2_125_3477_n1883, DP_OP_423J2_125_3477_n1882,
         DP_OP_423J2_125_3477_n1881, DP_OP_423J2_125_3477_n1880,
         DP_OP_423J2_125_3477_n1879, DP_OP_423J2_125_3477_n1878,
         DP_OP_423J2_125_3477_n1877, DP_OP_423J2_125_3477_n1876,
         DP_OP_423J2_125_3477_n1875, DP_OP_423J2_125_3477_n1874,
         DP_OP_423J2_125_3477_n1873, DP_OP_423J2_125_3477_n1871,
         DP_OP_423J2_125_3477_n1870, DP_OP_423J2_125_3477_n1869,
         DP_OP_423J2_125_3477_n1868, DP_OP_423J2_125_3477_n1867,
         DP_OP_423J2_125_3477_n1866, DP_OP_423J2_125_3477_n1865,
         DP_OP_423J2_125_3477_n1864, DP_OP_423J2_125_3477_n1863,
         DP_OP_423J2_125_3477_n1862, DP_OP_423J2_125_3477_n1861,
         DP_OP_423J2_125_3477_n1860, DP_OP_423J2_125_3477_n1859,
         DP_OP_423J2_125_3477_n1858, DP_OP_423J2_125_3477_n1857,
         DP_OP_423J2_125_3477_n1856, DP_OP_423J2_125_3477_n1855,
         DP_OP_423J2_125_3477_n1854, DP_OP_423J2_125_3477_n1853,
         DP_OP_423J2_125_3477_n1852, DP_OP_423J2_125_3477_n1851,
         DP_OP_423J2_125_3477_n1850, DP_OP_423J2_125_3477_n1849,
         DP_OP_423J2_125_3477_n1848, DP_OP_423J2_125_3477_n1847,
         DP_OP_423J2_125_3477_n1846, DP_OP_423J2_125_3477_n1845,
         DP_OP_423J2_125_3477_n1844, DP_OP_423J2_125_3477_n1843,
         DP_OP_423J2_125_3477_n1842, DP_OP_423J2_125_3477_n1841,
         DP_OP_423J2_125_3477_n1840, DP_OP_423J2_125_3477_n1839,
         DP_OP_423J2_125_3477_n1838, DP_OP_423J2_125_3477_n1837,
         DP_OP_423J2_125_3477_n1836, DP_OP_423J2_125_3477_n1835,
         DP_OP_423J2_125_3477_n1834, DP_OP_423J2_125_3477_n1833,
         DP_OP_423J2_125_3477_n1832, DP_OP_423J2_125_3477_n1831,
         DP_OP_423J2_125_3477_n1830, DP_OP_423J2_125_3477_n1829,
         DP_OP_423J2_125_3477_n1828, DP_OP_423J2_125_3477_n1827,
         DP_OP_423J2_125_3477_n1826, DP_OP_423J2_125_3477_n1825,
         DP_OP_423J2_125_3477_n1824, DP_OP_423J2_125_3477_n1823,
         DP_OP_423J2_125_3477_n1822, DP_OP_423J2_125_3477_n1821,
         DP_OP_423J2_125_3477_n1820, DP_OP_423J2_125_3477_n1819,
         DP_OP_423J2_125_3477_n1818, DP_OP_423J2_125_3477_n1817,
         DP_OP_423J2_125_3477_n1816, DP_OP_423J2_125_3477_n1815,
         DP_OP_423J2_125_3477_n1814, DP_OP_423J2_125_3477_n1813,
         DP_OP_423J2_125_3477_n1812, DP_OP_423J2_125_3477_n1811,
         DP_OP_423J2_125_3477_n1810, DP_OP_423J2_125_3477_n1809,
         DP_OP_423J2_125_3477_n1808, DP_OP_423J2_125_3477_n1807,
         DP_OP_423J2_125_3477_n1806, DP_OP_423J2_125_3477_n1805,
         DP_OP_423J2_125_3477_n1804, DP_OP_423J2_125_3477_n1803,
         DP_OP_423J2_125_3477_n1802, DP_OP_423J2_125_3477_n1801,
         DP_OP_423J2_125_3477_n1800, DP_OP_423J2_125_3477_n1799,
         DP_OP_423J2_125_3477_n1798, DP_OP_423J2_125_3477_n1797,
         DP_OP_423J2_125_3477_n1796, DP_OP_423J2_125_3477_n1795,
         DP_OP_423J2_125_3477_n1794, DP_OP_423J2_125_3477_n1793,
         DP_OP_423J2_125_3477_n1792, DP_OP_423J2_125_3477_n1791,
         DP_OP_423J2_125_3477_n1790, DP_OP_423J2_125_3477_n1789,
         DP_OP_423J2_125_3477_n1788, DP_OP_423J2_125_3477_n1787,
         DP_OP_423J2_125_3477_n1786, DP_OP_423J2_125_3477_n1785,
         DP_OP_423J2_125_3477_n1784, DP_OP_423J2_125_3477_n1783,
         DP_OP_423J2_125_3477_n1782, DP_OP_423J2_125_3477_n1781,
         DP_OP_423J2_125_3477_n1780, DP_OP_423J2_125_3477_n1779,
         DP_OP_423J2_125_3477_n1778, DP_OP_423J2_125_3477_n1777,
         DP_OP_423J2_125_3477_n1776, DP_OP_423J2_125_3477_n1775,
         DP_OP_423J2_125_3477_n1774, DP_OP_423J2_125_3477_n1773,
         DP_OP_423J2_125_3477_n1772, DP_OP_423J2_125_3477_n1771,
         DP_OP_423J2_125_3477_n1770, DP_OP_423J2_125_3477_n1769,
         DP_OP_423J2_125_3477_n1768, DP_OP_423J2_125_3477_n1767,
         DP_OP_423J2_125_3477_n1766, DP_OP_423J2_125_3477_n1765,
         DP_OP_423J2_125_3477_n1764, DP_OP_423J2_125_3477_n1763,
         DP_OP_423J2_125_3477_n1762, DP_OP_423J2_125_3477_n1761,
         DP_OP_423J2_125_3477_n1760, DP_OP_423J2_125_3477_n1759,
         DP_OP_423J2_125_3477_n1758, DP_OP_423J2_125_3477_n1757,
         DP_OP_423J2_125_3477_n1756, DP_OP_423J2_125_3477_n1755,
         DP_OP_423J2_125_3477_n1754, DP_OP_423J2_125_3477_n1753,
         DP_OP_423J2_125_3477_n1752, DP_OP_423J2_125_3477_n1751,
         DP_OP_423J2_125_3477_n1750, DP_OP_423J2_125_3477_n1749,
         DP_OP_423J2_125_3477_n1748, DP_OP_423J2_125_3477_n1747,
         DP_OP_423J2_125_3477_n1746, DP_OP_423J2_125_3477_n1745,
         DP_OP_423J2_125_3477_n1744, DP_OP_423J2_125_3477_n1743,
         DP_OP_423J2_125_3477_n1742, DP_OP_423J2_125_3477_n1741,
         DP_OP_423J2_125_3477_n1740, DP_OP_423J2_125_3477_n1739,
         DP_OP_423J2_125_3477_n1738, DP_OP_423J2_125_3477_n1737,
         DP_OP_423J2_125_3477_n1736, DP_OP_423J2_125_3477_n1735,
         DP_OP_423J2_125_3477_n1734, DP_OP_423J2_125_3477_n1733,
         DP_OP_423J2_125_3477_n1732, DP_OP_423J2_125_3477_n1731,
         DP_OP_423J2_125_3477_n1730, DP_OP_423J2_125_3477_n1729,
         DP_OP_423J2_125_3477_n1728, DP_OP_423J2_125_3477_n1727,
         DP_OP_423J2_125_3477_n1726, DP_OP_423J2_125_3477_n1725,
         DP_OP_423J2_125_3477_n1724, DP_OP_423J2_125_3477_n1723,
         DP_OP_423J2_125_3477_n1722, DP_OP_423J2_125_3477_n1721,
         DP_OP_423J2_125_3477_n1720, DP_OP_423J2_125_3477_n1719,
         DP_OP_423J2_125_3477_n1718, DP_OP_423J2_125_3477_n1717,
         DP_OP_423J2_125_3477_n1716, DP_OP_423J2_125_3477_n1715,
         DP_OP_423J2_125_3477_n1714, DP_OP_423J2_125_3477_n1713,
         DP_OP_423J2_125_3477_n1712, DP_OP_423J2_125_3477_n1711,
         DP_OP_423J2_125_3477_n1710, DP_OP_423J2_125_3477_n1709,
         DP_OP_423J2_125_3477_n1708, DP_OP_423J2_125_3477_n1707,
         DP_OP_423J2_125_3477_n1706, DP_OP_423J2_125_3477_n1705,
         DP_OP_423J2_125_3477_n1704, DP_OP_423J2_125_3477_n1703,
         DP_OP_423J2_125_3477_n1702, DP_OP_423J2_125_3477_n1701,
         DP_OP_423J2_125_3477_n1700, DP_OP_423J2_125_3477_n1699,
         DP_OP_423J2_125_3477_n1698, DP_OP_423J2_125_3477_n1697,
         DP_OP_423J2_125_3477_n1696, DP_OP_423J2_125_3477_n1695,
         DP_OP_423J2_125_3477_n1694, DP_OP_423J2_125_3477_n1693,
         DP_OP_423J2_125_3477_n1692, DP_OP_423J2_125_3477_n1691,
         DP_OP_423J2_125_3477_n1690, DP_OP_423J2_125_3477_n1689,
         DP_OP_423J2_125_3477_n1688, DP_OP_423J2_125_3477_n1687,
         DP_OP_423J2_125_3477_n1686, DP_OP_423J2_125_3477_n1685,
         DP_OP_423J2_125_3477_n1684, DP_OP_423J2_125_3477_n1683,
         DP_OP_423J2_125_3477_n1682, DP_OP_423J2_125_3477_n1681,
         DP_OP_423J2_125_3477_n1680, DP_OP_423J2_125_3477_n1679,
         DP_OP_423J2_125_3477_n1678, DP_OP_423J2_125_3477_n1677,
         DP_OP_423J2_125_3477_n1676, DP_OP_423J2_125_3477_n1675,
         DP_OP_423J2_125_3477_n1674, DP_OP_423J2_125_3477_n1673,
         DP_OP_423J2_125_3477_n1672, DP_OP_423J2_125_3477_n1671,
         DP_OP_423J2_125_3477_n1670, DP_OP_423J2_125_3477_n1669,
         DP_OP_423J2_125_3477_n1668, DP_OP_423J2_125_3477_n1667,
         DP_OP_423J2_125_3477_n1666, DP_OP_423J2_125_3477_n1665,
         DP_OP_423J2_125_3477_n1664, DP_OP_423J2_125_3477_n1663,
         DP_OP_423J2_125_3477_n1662, DP_OP_423J2_125_3477_n1661,
         DP_OP_423J2_125_3477_n1660, DP_OP_423J2_125_3477_n1659,
         DP_OP_423J2_125_3477_n1658, DP_OP_423J2_125_3477_n1657,
         DP_OP_423J2_125_3477_n1656, DP_OP_423J2_125_3477_n1655,
         DP_OP_423J2_125_3477_n1654, DP_OP_423J2_125_3477_n1653,
         DP_OP_423J2_125_3477_n1652, DP_OP_423J2_125_3477_n1651,
         DP_OP_423J2_125_3477_n1650, DP_OP_423J2_125_3477_n1649,
         DP_OP_423J2_125_3477_n1648, DP_OP_423J2_125_3477_n1647,
         DP_OP_423J2_125_3477_n1646, DP_OP_423J2_125_3477_n1645,
         DP_OP_423J2_125_3477_n1644, DP_OP_423J2_125_3477_n1643,
         DP_OP_423J2_125_3477_n1642, DP_OP_423J2_125_3477_n1641,
         DP_OP_423J2_125_3477_n1640, DP_OP_423J2_125_3477_n1639,
         DP_OP_423J2_125_3477_n1638, DP_OP_423J2_125_3477_n1637,
         DP_OP_423J2_125_3477_n1636, DP_OP_423J2_125_3477_n1635,
         DP_OP_423J2_125_3477_n1634, DP_OP_423J2_125_3477_n1633,
         DP_OP_423J2_125_3477_n1632, DP_OP_423J2_125_3477_n1631,
         DP_OP_423J2_125_3477_n1630, DP_OP_423J2_125_3477_n1629,
         DP_OP_423J2_125_3477_n1628, DP_OP_423J2_125_3477_n1627,
         DP_OP_423J2_125_3477_n1626, DP_OP_423J2_125_3477_n1625,
         DP_OP_423J2_125_3477_n1624, DP_OP_423J2_125_3477_n1623,
         DP_OP_423J2_125_3477_n1622, DP_OP_423J2_125_3477_n1621,
         DP_OP_423J2_125_3477_n1620, DP_OP_423J2_125_3477_n1619,
         DP_OP_423J2_125_3477_n1618, DP_OP_423J2_125_3477_n1617,
         DP_OP_423J2_125_3477_n1616, DP_OP_423J2_125_3477_n1615,
         DP_OP_423J2_125_3477_n1614, DP_OP_423J2_125_3477_n1613,
         DP_OP_423J2_125_3477_n1612, DP_OP_423J2_125_3477_n1611,
         DP_OP_423J2_125_3477_n1610, DP_OP_423J2_125_3477_n1609,
         DP_OP_423J2_125_3477_n1608, DP_OP_423J2_125_3477_n1607,
         DP_OP_423J2_125_3477_n1606, DP_OP_423J2_125_3477_n1605,
         DP_OP_423J2_125_3477_n1604, DP_OP_423J2_125_3477_n1603,
         DP_OP_423J2_125_3477_n1602, DP_OP_423J2_125_3477_n1601,
         DP_OP_423J2_125_3477_n1600, DP_OP_423J2_125_3477_n1599,
         DP_OP_423J2_125_3477_n1598, DP_OP_423J2_125_3477_n1597,
         DP_OP_423J2_125_3477_n1596, DP_OP_423J2_125_3477_n1595,
         DP_OP_423J2_125_3477_n1594, DP_OP_423J2_125_3477_n1593,
         DP_OP_423J2_125_3477_n1592, DP_OP_423J2_125_3477_n1591,
         DP_OP_423J2_125_3477_n1590, DP_OP_423J2_125_3477_n1589,
         DP_OP_423J2_125_3477_n1588, DP_OP_423J2_125_3477_n1587,
         DP_OP_423J2_125_3477_n1586, DP_OP_423J2_125_3477_n1585,
         DP_OP_423J2_125_3477_n1584, DP_OP_423J2_125_3477_n1583,
         DP_OP_423J2_125_3477_n1582, DP_OP_423J2_125_3477_n1581,
         DP_OP_423J2_125_3477_n1580, DP_OP_423J2_125_3477_n1579,
         DP_OP_423J2_125_3477_n1578, DP_OP_423J2_125_3477_n1577,
         DP_OP_423J2_125_3477_n1576, DP_OP_423J2_125_3477_n1575,
         DP_OP_423J2_125_3477_n1574, DP_OP_423J2_125_3477_n1573,
         DP_OP_423J2_125_3477_n1572, DP_OP_423J2_125_3477_n1571,
         DP_OP_423J2_125_3477_n1570, DP_OP_423J2_125_3477_n1569,
         DP_OP_423J2_125_3477_n1568, DP_OP_423J2_125_3477_n1567,
         DP_OP_423J2_125_3477_n1566, DP_OP_423J2_125_3477_n1565,
         DP_OP_423J2_125_3477_n1564, DP_OP_423J2_125_3477_n1563,
         DP_OP_423J2_125_3477_n1562, DP_OP_423J2_125_3477_n1561,
         DP_OP_423J2_125_3477_n1560, DP_OP_423J2_125_3477_n1559,
         DP_OP_423J2_125_3477_n1558, DP_OP_423J2_125_3477_n1557,
         DP_OP_423J2_125_3477_n1556, DP_OP_423J2_125_3477_n1555,
         DP_OP_423J2_125_3477_n1554, DP_OP_423J2_125_3477_n1553,
         DP_OP_423J2_125_3477_n1552, DP_OP_423J2_125_3477_n1551,
         DP_OP_423J2_125_3477_n1550, DP_OP_423J2_125_3477_n1549,
         DP_OP_423J2_125_3477_n1548, DP_OP_423J2_125_3477_n1547,
         DP_OP_423J2_125_3477_n1546, DP_OP_423J2_125_3477_n1545,
         DP_OP_423J2_125_3477_n1544, DP_OP_423J2_125_3477_n1543,
         DP_OP_423J2_125_3477_n1542, DP_OP_423J2_125_3477_n1541,
         DP_OP_423J2_125_3477_n1540, DP_OP_423J2_125_3477_n1539,
         DP_OP_423J2_125_3477_n1538, DP_OP_423J2_125_3477_n1537,
         DP_OP_423J2_125_3477_n1536, DP_OP_423J2_125_3477_n1535,
         DP_OP_423J2_125_3477_n1534, DP_OP_423J2_125_3477_n1533,
         DP_OP_423J2_125_3477_n1532, DP_OP_423J2_125_3477_n1531,
         DP_OP_423J2_125_3477_n1530, DP_OP_423J2_125_3477_n1529,
         DP_OP_423J2_125_3477_n1528, DP_OP_423J2_125_3477_n1527,
         DP_OP_423J2_125_3477_n1526, DP_OP_423J2_125_3477_n1525,
         DP_OP_423J2_125_3477_n1524, DP_OP_423J2_125_3477_n1523,
         DP_OP_423J2_125_3477_n1522, DP_OP_423J2_125_3477_n1521,
         DP_OP_423J2_125_3477_n1520, DP_OP_423J2_125_3477_n1519,
         DP_OP_423J2_125_3477_n1518, DP_OP_423J2_125_3477_n1517,
         DP_OP_423J2_125_3477_n1516, DP_OP_423J2_125_3477_n1515,
         DP_OP_423J2_125_3477_n1514, DP_OP_423J2_125_3477_n1513,
         DP_OP_423J2_125_3477_n1512, DP_OP_423J2_125_3477_n1511,
         DP_OP_423J2_125_3477_n1510, DP_OP_423J2_125_3477_n1509,
         DP_OP_423J2_125_3477_n1508, DP_OP_423J2_125_3477_n1507,
         DP_OP_423J2_125_3477_n1506, DP_OP_423J2_125_3477_n1505,
         DP_OP_423J2_125_3477_n1504, DP_OP_423J2_125_3477_n1503,
         DP_OP_423J2_125_3477_n1502, DP_OP_423J2_125_3477_n1501,
         DP_OP_423J2_125_3477_n1500, DP_OP_423J2_125_3477_n1499,
         DP_OP_423J2_125_3477_n1498, DP_OP_423J2_125_3477_n1497,
         DP_OP_423J2_125_3477_n1496, DP_OP_423J2_125_3477_n1495,
         DP_OP_423J2_125_3477_n1494, DP_OP_423J2_125_3477_n1493,
         DP_OP_423J2_125_3477_n1492, DP_OP_423J2_125_3477_n1491,
         DP_OP_423J2_125_3477_n1490, DP_OP_423J2_125_3477_n1489,
         DP_OP_423J2_125_3477_n1488, DP_OP_423J2_125_3477_n1487,
         DP_OP_423J2_125_3477_n1486, DP_OP_423J2_125_3477_n1485,
         DP_OP_423J2_125_3477_n1484, DP_OP_423J2_125_3477_n1483,
         DP_OP_423J2_125_3477_n1482, DP_OP_423J2_125_3477_n1481,
         DP_OP_423J2_125_3477_n1480, DP_OP_423J2_125_3477_n1479,
         DP_OP_423J2_125_3477_n1478, DP_OP_423J2_125_3477_n1477,
         DP_OP_423J2_125_3477_n1476, DP_OP_423J2_125_3477_n1475,
         DP_OP_423J2_125_3477_n1474, DP_OP_423J2_125_3477_n1473,
         DP_OP_423J2_125_3477_n1472, DP_OP_423J2_125_3477_n1471,
         DP_OP_423J2_125_3477_n1470, DP_OP_423J2_125_3477_n1469,
         DP_OP_423J2_125_3477_n1468, DP_OP_423J2_125_3477_n1467,
         DP_OP_423J2_125_3477_n1466, DP_OP_423J2_125_3477_n1465,
         DP_OP_423J2_125_3477_n1464, DP_OP_423J2_125_3477_n1463,
         DP_OP_423J2_125_3477_n1462, DP_OP_423J2_125_3477_n1461,
         DP_OP_423J2_125_3477_n1460, DP_OP_423J2_125_3477_n1459,
         DP_OP_423J2_125_3477_n1458, DP_OP_423J2_125_3477_n1457,
         DP_OP_423J2_125_3477_n1456, DP_OP_423J2_125_3477_n1455,
         DP_OP_423J2_125_3477_n1454, DP_OP_423J2_125_3477_n1453,
         DP_OP_423J2_125_3477_n1452, DP_OP_423J2_125_3477_n1451,
         DP_OP_423J2_125_3477_n1450, DP_OP_423J2_125_3477_n1449,
         DP_OP_423J2_125_3477_n1448, DP_OP_423J2_125_3477_n1447,
         DP_OP_423J2_125_3477_n1446, DP_OP_423J2_125_3477_n1445,
         DP_OP_423J2_125_3477_n1444, DP_OP_423J2_125_3477_n1443,
         DP_OP_423J2_125_3477_n1442, DP_OP_423J2_125_3477_n1441,
         DP_OP_423J2_125_3477_n1440, DP_OP_423J2_125_3477_n1439,
         DP_OP_423J2_125_3477_n1438, DP_OP_423J2_125_3477_n1437,
         DP_OP_423J2_125_3477_n1436, DP_OP_423J2_125_3477_n1435,
         DP_OP_423J2_125_3477_n1434, DP_OP_423J2_125_3477_n1433,
         DP_OP_423J2_125_3477_n1432, DP_OP_423J2_125_3477_n1431,
         DP_OP_423J2_125_3477_n1430, DP_OP_423J2_125_3477_n1429,
         DP_OP_423J2_125_3477_n1428, DP_OP_423J2_125_3477_n1427,
         DP_OP_423J2_125_3477_n1426, DP_OP_423J2_125_3477_n1425,
         DP_OP_423J2_125_3477_n1424, DP_OP_423J2_125_3477_n1423,
         DP_OP_423J2_125_3477_n1422, DP_OP_423J2_125_3477_n1421,
         DP_OP_423J2_125_3477_n1420, DP_OP_423J2_125_3477_n1419,
         DP_OP_423J2_125_3477_n1418, DP_OP_423J2_125_3477_n1417,
         DP_OP_423J2_125_3477_n1416, DP_OP_423J2_125_3477_n1415,
         DP_OP_423J2_125_3477_n1414, DP_OP_423J2_125_3477_n1413,
         DP_OP_423J2_125_3477_n1412, DP_OP_423J2_125_3477_n1411,
         DP_OP_423J2_125_3477_n1410, DP_OP_423J2_125_3477_n1409,
         DP_OP_423J2_125_3477_n1408, DP_OP_423J2_125_3477_n1407,
         DP_OP_423J2_125_3477_n1406, DP_OP_423J2_125_3477_n1405,
         DP_OP_423J2_125_3477_n1404, DP_OP_423J2_125_3477_n1403,
         DP_OP_423J2_125_3477_n1402, DP_OP_423J2_125_3477_n1401,
         DP_OP_423J2_125_3477_n1400, DP_OP_423J2_125_3477_n1399,
         DP_OP_423J2_125_3477_n1398, DP_OP_423J2_125_3477_n1397,
         DP_OP_423J2_125_3477_n1396, DP_OP_423J2_125_3477_n1395,
         DP_OP_423J2_125_3477_n1394, DP_OP_423J2_125_3477_n1393,
         DP_OP_423J2_125_3477_n1392, DP_OP_423J2_125_3477_n1391,
         DP_OP_423J2_125_3477_n1390, DP_OP_423J2_125_3477_n1389,
         DP_OP_423J2_125_3477_n1388, DP_OP_423J2_125_3477_n1387,
         DP_OP_423J2_125_3477_n1386, DP_OP_423J2_125_3477_n1385,
         DP_OP_423J2_125_3477_n1384, DP_OP_423J2_125_3477_n1383,
         DP_OP_423J2_125_3477_n1382, DP_OP_423J2_125_3477_n1381,
         DP_OP_423J2_125_3477_n1380, DP_OP_423J2_125_3477_n1379,
         DP_OP_423J2_125_3477_n1378, DP_OP_423J2_125_3477_n1377,
         DP_OP_423J2_125_3477_n1376, DP_OP_423J2_125_3477_n1375,
         DP_OP_423J2_125_3477_n1374, DP_OP_423J2_125_3477_n1373,
         DP_OP_423J2_125_3477_n1372, DP_OP_423J2_125_3477_n1371,
         DP_OP_423J2_125_3477_n1370, DP_OP_423J2_125_3477_n1369,
         DP_OP_423J2_125_3477_n1368, DP_OP_423J2_125_3477_n1367,
         DP_OP_423J2_125_3477_n1366, DP_OP_423J2_125_3477_n1365,
         DP_OP_423J2_125_3477_n1364, DP_OP_423J2_125_3477_n1363,
         DP_OP_423J2_125_3477_n1362, DP_OP_423J2_125_3477_n1361,
         DP_OP_423J2_125_3477_n1360, DP_OP_423J2_125_3477_n1359,
         DP_OP_423J2_125_3477_n1358, DP_OP_423J2_125_3477_n1357,
         DP_OP_423J2_125_3477_n1356, DP_OP_423J2_125_3477_n1355,
         DP_OP_423J2_125_3477_n1354, DP_OP_423J2_125_3477_n1353,
         DP_OP_423J2_125_3477_n1352, DP_OP_423J2_125_3477_n1351,
         DP_OP_423J2_125_3477_n1350, DP_OP_423J2_125_3477_n1349,
         DP_OP_423J2_125_3477_n1348, DP_OP_423J2_125_3477_n1347,
         DP_OP_423J2_125_3477_n1346, DP_OP_423J2_125_3477_n1345,
         DP_OP_423J2_125_3477_n1344, DP_OP_423J2_125_3477_n1343,
         DP_OP_423J2_125_3477_n1342, DP_OP_423J2_125_3477_n1341,
         DP_OP_423J2_125_3477_n1340, DP_OP_423J2_125_3477_n1339,
         DP_OP_423J2_125_3477_n1338, DP_OP_423J2_125_3477_n1337,
         DP_OP_423J2_125_3477_n1336, DP_OP_423J2_125_3477_n1335,
         DP_OP_423J2_125_3477_n1334, DP_OP_423J2_125_3477_n1333,
         DP_OP_423J2_125_3477_n1332, DP_OP_423J2_125_3477_n1331,
         DP_OP_423J2_125_3477_n1330, DP_OP_423J2_125_3477_n1329,
         DP_OP_423J2_125_3477_n1328, DP_OP_423J2_125_3477_n1327,
         DP_OP_423J2_125_3477_n1326, DP_OP_423J2_125_3477_n1325,
         DP_OP_423J2_125_3477_n1324, DP_OP_423J2_125_3477_n1323,
         DP_OP_423J2_125_3477_n1322, DP_OP_423J2_125_3477_n1321,
         DP_OP_423J2_125_3477_n1320, DP_OP_423J2_125_3477_n1319,
         DP_OP_423J2_125_3477_n1318, DP_OP_423J2_125_3477_n1317,
         DP_OP_423J2_125_3477_n1316, DP_OP_423J2_125_3477_n1315,
         DP_OP_423J2_125_3477_n1314, DP_OP_423J2_125_3477_n1313,
         DP_OP_423J2_125_3477_n1312, DP_OP_423J2_125_3477_n1311,
         DP_OP_423J2_125_3477_n1310, DP_OP_423J2_125_3477_n1309,
         DP_OP_423J2_125_3477_n1308, DP_OP_423J2_125_3477_n1307,
         DP_OP_423J2_125_3477_n1306, DP_OP_423J2_125_3477_n1305,
         DP_OP_423J2_125_3477_n1304, DP_OP_423J2_125_3477_n1303,
         DP_OP_423J2_125_3477_n1302, DP_OP_423J2_125_3477_n1301,
         DP_OP_423J2_125_3477_n1300, DP_OP_423J2_125_3477_n1299,
         DP_OP_423J2_125_3477_n1298, DP_OP_423J2_125_3477_n1297,
         DP_OP_423J2_125_3477_n1296, DP_OP_423J2_125_3477_n1295,
         DP_OP_423J2_125_3477_n1294, DP_OP_423J2_125_3477_n1293,
         DP_OP_423J2_125_3477_n1292, DP_OP_423J2_125_3477_n1291,
         DP_OP_423J2_125_3477_n1290, DP_OP_423J2_125_3477_n1289,
         DP_OP_423J2_125_3477_n1288, DP_OP_423J2_125_3477_n1287,
         DP_OP_423J2_125_3477_n1286, DP_OP_423J2_125_3477_n1285,
         DP_OP_423J2_125_3477_n1284, DP_OP_423J2_125_3477_n1283,
         DP_OP_423J2_125_3477_n1282, DP_OP_423J2_125_3477_n1281,
         DP_OP_423J2_125_3477_n1280, DP_OP_423J2_125_3477_n1279,
         DP_OP_423J2_125_3477_n1278, DP_OP_423J2_125_3477_n1277,
         DP_OP_423J2_125_3477_n1276, DP_OP_423J2_125_3477_n1275,
         DP_OP_423J2_125_3477_n1274, DP_OP_423J2_125_3477_n1273,
         DP_OP_423J2_125_3477_n1272, DP_OP_423J2_125_3477_n1271,
         DP_OP_423J2_125_3477_n1270, DP_OP_423J2_125_3477_n1269,
         DP_OP_423J2_125_3477_n1268, DP_OP_423J2_125_3477_n1267,
         DP_OP_423J2_125_3477_n1266, DP_OP_423J2_125_3477_n1265,
         DP_OP_423J2_125_3477_n1264, DP_OP_423J2_125_3477_n1263,
         DP_OP_423J2_125_3477_n1262, DP_OP_423J2_125_3477_n1261,
         DP_OP_423J2_125_3477_n1260, DP_OP_423J2_125_3477_n1259,
         DP_OP_423J2_125_3477_n1258, DP_OP_423J2_125_3477_n1257,
         DP_OP_423J2_125_3477_n1256, DP_OP_423J2_125_3477_n1255,
         DP_OP_423J2_125_3477_n1254, DP_OP_423J2_125_3477_n1253,
         DP_OP_423J2_125_3477_n1252, DP_OP_423J2_125_3477_n1251,
         DP_OP_423J2_125_3477_n1250, DP_OP_423J2_125_3477_n1249,
         DP_OP_423J2_125_3477_n1248, DP_OP_423J2_125_3477_n1247,
         DP_OP_423J2_125_3477_n1246, DP_OP_423J2_125_3477_n1245,
         DP_OP_423J2_125_3477_n1244, DP_OP_423J2_125_3477_n1243,
         DP_OP_423J2_125_3477_n1242, DP_OP_423J2_125_3477_n1241,
         DP_OP_423J2_125_3477_n1240, DP_OP_423J2_125_3477_n1239,
         DP_OP_423J2_125_3477_n1238, DP_OP_423J2_125_3477_n1237,
         DP_OP_423J2_125_3477_n1236, DP_OP_423J2_125_3477_n1235,
         DP_OP_423J2_125_3477_n1234, DP_OP_423J2_125_3477_n1233,
         DP_OP_423J2_125_3477_n1232, DP_OP_423J2_125_3477_n1231,
         DP_OP_423J2_125_3477_n1230, DP_OP_423J2_125_3477_n1229,
         DP_OP_423J2_125_3477_n1228, DP_OP_423J2_125_3477_n1227,
         DP_OP_423J2_125_3477_n1226, DP_OP_423J2_125_3477_n1225,
         DP_OP_423J2_125_3477_n1224, DP_OP_423J2_125_3477_n1223,
         DP_OP_423J2_125_3477_n1222, DP_OP_423J2_125_3477_n1221,
         DP_OP_423J2_125_3477_n1220, DP_OP_423J2_125_3477_n1219,
         DP_OP_423J2_125_3477_n1218, DP_OP_423J2_125_3477_n1217,
         DP_OP_423J2_125_3477_n1216, DP_OP_423J2_125_3477_n1215,
         DP_OP_423J2_125_3477_n1214, DP_OP_423J2_125_3477_n1213,
         DP_OP_423J2_125_3477_n1212, DP_OP_423J2_125_3477_n1211,
         DP_OP_423J2_125_3477_n1210, DP_OP_423J2_125_3477_n1209,
         DP_OP_423J2_125_3477_n1208, DP_OP_423J2_125_3477_n1207,
         DP_OP_423J2_125_3477_n1206, DP_OP_423J2_125_3477_n1205,
         DP_OP_423J2_125_3477_n1204, DP_OP_423J2_125_3477_n1203,
         DP_OP_423J2_125_3477_n1202, DP_OP_423J2_125_3477_n1201,
         DP_OP_423J2_125_3477_n1200, DP_OP_423J2_125_3477_n1199,
         DP_OP_423J2_125_3477_n1198, DP_OP_423J2_125_3477_n1197,
         DP_OP_423J2_125_3477_n1196, DP_OP_423J2_125_3477_n1195,
         DP_OP_423J2_125_3477_n1194, DP_OP_423J2_125_3477_n1193,
         DP_OP_423J2_125_3477_n1192, DP_OP_423J2_125_3477_n1191,
         DP_OP_423J2_125_3477_n1190, DP_OP_423J2_125_3477_n1189,
         DP_OP_423J2_125_3477_n1188, DP_OP_423J2_125_3477_n1187,
         DP_OP_423J2_125_3477_n1186, DP_OP_423J2_125_3477_n1185,
         DP_OP_423J2_125_3477_n1184, DP_OP_423J2_125_3477_n1183,
         DP_OP_423J2_125_3477_n1182, DP_OP_423J2_125_3477_n1181,
         DP_OP_423J2_125_3477_n1180, DP_OP_423J2_125_3477_n1179,
         DP_OP_423J2_125_3477_n1178, DP_OP_423J2_125_3477_n1177,
         DP_OP_423J2_125_3477_n1176, DP_OP_423J2_125_3477_n1175,
         DP_OP_423J2_125_3477_n1174, DP_OP_423J2_125_3477_n1173,
         DP_OP_423J2_125_3477_n1172, DP_OP_423J2_125_3477_n1171,
         DP_OP_423J2_125_3477_n1170, DP_OP_423J2_125_3477_n1169,
         DP_OP_423J2_125_3477_n1168, DP_OP_423J2_125_3477_n1167,
         DP_OP_423J2_125_3477_n1166, DP_OP_423J2_125_3477_n1165,
         DP_OP_423J2_125_3477_n1164, DP_OP_423J2_125_3477_n1163,
         DP_OP_423J2_125_3477_n1162, DP_OP_423J2_125_3477_n1161,
         DP_OP_423J2_125_3477_n1160, DP_OP_423J2_125_3477_n1159,
         DP_OP_423J2_125_3477_n1158, DP_OP_423J2_125_3477_n1157,
         DP_OP_423J2_125_3477_n1156, DP_OP_423J2_125_3477_n1155,
         DP_OP_423J2_125_3477_n1154, DP_OP_423J2_125_3477_n1153,
         DP_OP_423J2_125_3477_n1152, DP_OP_423J2_125_3477_n1151,
         DP_OP_423J2_125_3477_n1150, DP_OP_423J2_125_3477_n1149,
         DP_OP_423J2_125_3477_n1148, DP_OP_423J2_125_3477_n1147,
         DP_OP_423J2_125_3477_n1146, DP_OP_423J2_125_3477_n1145,
         DP_OP_423J2_125_3477_n1144, DP_OP_423J2_125_3477_n1143,
         DP_OP_423J2_125_3477_n1142, DP_OP_423J2_125_3477_n1141,
         DP_OP_423J2_125_3477_n1140, DP_OP_423J2_125_3477_n1139,
         DP_OP_423J2_125_3477_n1138, DP_OP_423J2_125_3477_n1137,
         DP_OP_423J2_125_3477_n1136, DP_OP_423J2_125_3477_n1135,
         DP_OP_423J2_125_3477_n1134, DP_OP_423J2_125_3477_n1133,
         DP_OP_423J2_125_3477_n1132, DP_OP_423J2_125_3477_n1131,
         DP_OP_423J2_125_3477_n1130, DP_OP_423J2_125_3477_n1129,
         DP_OP_423J2_125_3477_n1128, DP_OP_423J2_125_3477_n1127,
         DP_OP_423J2_125_3477_n1126, DP_OP_423J2_125_3477_n1125,
         DP_OP_423J2_125_3477_n1124, DP_OP_423J2_125_3477_n1123,
         DP_OP_423J2_125_3477_n1122, DP_OP_423J2_125_3477_n1121,
         DP_OP_423J2_125_3477_n1120, DP_OP_423J2_125_3477_n1119,
         DP_OP_423J2_125_3477_n1118, DP_OP_423J2_125_3477_n1117,
         DP_OP_423J2_125_3477_n1116, DP_OP_423J2_125_3477_n1115,
         DP_OP_423J2_125_3477_n1114, DP_OP_423J2_125_3477_n1113,
         DP_OP_423J2_125_3477_n1112, DP_OP_423J2_125_3477_n1111,
         DP_OP_423J2_125_3477_n1110, DP_OP_423J2_125_3477_n1109,
         DP_OP_423J2_125_3477_n1108, DP_OP_423J2_125_3477_n1107,
         DP_OP_423J2_125_3477_n1106, DP_OP_423J2_125_3477_n1105,
         DP_OP_423J2_125_3477_n1104, DP_OP_423J2_125_3477_n1103,
         DP_OP_423J2_125_3477_n1102, DP_OP_423J2_125_3477_n1101,
         DP_OP_423J2_125_3477_n1100, DP_OP_423J2_125_3477_n1099,
         DP_OP_423J2_125_3477_n1098, DP_OP_423J2_125_3477_n1097,
         DP_OP_423J2_125_3477_n1096, DP_OP_423J2_125_3477_n1095,
         DP_OP_423J2_125_3477_n1094, DP_OP_423J2_125_3477_n1093,
         DP_OP_423J2_125_3477_n1092, DP_OP_423J2_125_3477_n1091,
         DP_OP_423J2_125_3477_n1090, DP_OP_423J2_125_3477_n1089,
         DP_OP_423J2_125_3477_n1088, DP_OP_423J2_125_3477_n1087,
         DP_OP_423J2_125_3477_n1086, DP_OP_423J2_125_3477_n1085,
         DP_OP_423J2_125_3477_n1084, DP_OP_423J2_125_3477_n1083,
         DP_OP_423J2_125_3477_n1082, DP_OP_423J2_125_3477_n1081,
         DP_OP_423J2_125_3477_n1080, DP_OP_423J2_125_3477_n1079,
         DP_OP_423J2_125_3477_n1078, DP_OP_423J2_125_3477_n1077,
         DP_OP_423J2_125_3477_n1076, DP_OP_423J2_125_3477_n1075,
         DP_OP_423J2_125_3477_n1074, DP_OP_423J2_125_3477_n1073,
         DP_OP_423J2_125_3477_n1072, DP_OP_423J2_125_3477_n1071,
         DP_OP_423J2_125_3477_n1070, DP_OP_423J2_125_3477_n1069,
         DP_OP_423J2_125_3477_n1068, DP_OP_423J2_125_3477_n1067,
         DP_OP_423J2_125_3477_n1066, DP_OP_423J2_125_3477_n1065,
         DP_OP_423J2_125_3477_n1064, DP_OP_423J2_125_3477_n1063,
         DP_OP_423J2_125_3477_n1062, DP_OP_423J2_125_3477_n1061,
         DP_OP_423J2_125_3477_n1060, DP_OP_423J2_125_3477_n1059,
         DP_OP_423J2_125_3477_n1058, DP_OP_423J2_125_3477_n1057,
         DP_OP_423J2_125_3477_n1056, DP_OP_423J2_125_3477_n1055,
         DP_OP_423J2_125_3477_n1054, DP_OP_423J2_125_3477_n1053,
         DP_OP_423J2_125_3477_n1052, DP_OP_423J2_125_3477_n1051,
         DP_OP_423J2_125_3477_n1050, DP_OP_423J2_125_3477_n1049,
         DP_OP_423J2_125_3477_n1048, DP_OP_423J2_125_3477_n1047,
         DP_OP_423J2_125_3477_n1046, DP_OP_423J2_125_3477_n1045,
         DP_OP_423J2_125_3477_n1044, DP_OP_423J2_125_3477_n1043,
         DP_OP_423J2_125_3477_n1042, DP_OP_423J2_125_3477_n1041,
         DP_OP_423J2_125_3477_n1040, DP_OP_423J2_125_3477_n1039,
         DP_OP_423J2_125_3477_n1038, DP_OP_423J2_125_3477_n1037,
         DP_OP_423J2_125_3477_n1036, DP_OP_423J2_125_3477_n1035,
         DP_OP_423J2_125_3477_n1034, DP_OP_423J2_125_3477_n1033,
         DP_OP_423J2_125_3477_n1032, DP_OP_423J2_125_3477_n1031,
         DP_OP_423J2_125_3477_n1030, DP_OP_423J2_125_3477_n1029,
         DP_OP_423J2_125_3477_n1028, DP_OP_423J2_125_3477_n1027,
         DP_OP_423J2_125_3477_n1026, DP_OP_423J2_125_3477_n1025,
         DP_OP_423J2_125_3477_n1024, DP_OP_423J2_125_3477_n1023,
         DP_OP_423J2_125_3477_n1022, DP_OP_423J2_125_3477_n1021,
         DP_OP_423J2_125_3477_n1020, DP_OP_423J2_125_3477_n1019,
         DP_OP_423J2_125_3477_n1018, DP_OP_423J2_125_3477_n1017,
         DP_OP_423J2_125_3477_n1016, DP_OP_423J2_125_3477_n1015,
         DP_OP_423J2_125_3477_n1014, DP_OP_423J2_125_3477_n1013,
         DP_OP_423J2_125_3477_n1012, DP_OP_423J2_125_3477_n1011,
         DP_OP_423J2_125_3477_n1010, DP_OP_423J2_125_3477_n1009,
         DP_OP_423J2_125_3477_n1008, DP_OP_423J2_125_3477_n1007,
         DP_OP_423J2_125_3477_n1006, DP_OP_423J2_125_3477_n1005,
         DP_OP_423J2_125_3477_n1004, DP_OP_423J2_125_3477_n1003,
         DP_OP_423J2_125_3477_n1002, DP_OP_423J2_125_3477_n1001,
         DP_OP_423J2_125_3477_n1000, DP_OP_423J2_125_3477_n999,
         DP_OP_423J2_125_3477_n998, DP_OP_423J2_125_3477_n997,
         DP_OP_423J2_125_3477_n996, DP_OP_423J2_125_3477_n995,
         DP_OP_423J2_125_3477_n994, DP_OP_423J2_125_3477_n993,
         DP_OP_423J2_125_3477_n992, DP_OP_423J2_125_3477_n991,
         DP_OP_423J2_125_3477_n990, DP_OP_423J2_125_3477_n989,
         DP_OP_423J2_125_3477_n988, DP_OP_423J2_125_3477_n987,
         DP_OP_423J2_125_3477_n986, DP_OP_423J2_125_3477_n985,
         DP_OP_423J2_125_3477_n984, DP_OP_423J2_125_3477_n983,
         DP_OP_423J2_125_3477_n982, DP_OP_423J2_125_3477_n981,
         DP_OP_423J2_125_3477_n980, DP_OP_423J2_125_3477_n979,
         DP_OP_423J2_125_3477_n978, DP_OP_423J2_125_3477_n977,
         DP_OP_423J2_125_3477_n976, DP_OP_423J2_125_3477_n975,
         DP_OP_423J2_125_3477_n974, DP_OP_423J2_125_3477_n973,
         DP_OP_423J2_125_3477_n972, DP_OP_423J2_125_3477_n971,
         DP_OP_423J2_125_3477_n970, DP_OP_423J2_125_3477_n969,
         DP_OP_423J2_125_3477_n968, DP_OP_423J2_125_3477_n967,
         DP_OP_423J2_125_3477_n966, DP_OP_423J2_125_3477_n965,
         DP_OP_423J2_125_3477_n964, DP_OP_423J2_125_3477_n963,
         DP_OP_423J2_125_3477_n962, DP_OP_423J2_125_3477_n961,
         DP_OP_423J2_125_3477_n960, DP_OP_423J2_125_3477_n959,
         DP_OP_423J2_125_3477_n958, DP_OP_423J2_125_3477_n957,
         DP_OP_423J2_125_3477_n956, DP_OP_423J2_125_3477_n955,
         DP_OP_423J2_125_3477_n954, DP_OP_423J2_125_3477_n953,
         DP_OP_423J2_125_3477_n952, DP_OP_423J2_125_3477_n951,
         DP_OP_423J2_125_3477_n950, DP_OP_423J2_125_3477_n949,
         DP_OP_423J2_125_3477_n948, DP_OP_423J2_125_3477_n947,
         DP_OP_423J2_125_3477_n946, DP_OP_423J2_125_3477_n945,
         DP_OP_423J2_125_3477_n944, DP_OP_423J2_125_3477_n943,
         DP_OP_423J2_125_3477_n942, DP_OP_423J2_125_3477_n941,
         DP_OP_423J2_125_3477_n940, DP_OP_423J2_125_3477_n939,
         DP_OP_423J2_125_3477_n938, DP_OP_423J2_125_3477_n937,
         DP_OP_423J2_125_3477_n936, DP_OP_423J2_125_3477_n935,
         DP_OP_423J2_125_3477_n934, DP_OP_423J2_125_3477_n933,
         DP_OP_423J2_125_3477_n932, DP_OP_423J2_125_3477_n931,
         DP_OP_423J2_125_3477_n930, DP_OP_423J2_125_3477_n929,
         DP_OP_423J2_125_3477_n928, DP_OP_423J2_125_3477_n927,
         DP_OP_423J2_125_3477_n926, DP_OP_423J2_125_3477_n925,
         DP_OP_423J2_125_3477_n924, DP_OP_423J2_125_3477_n923,
         DP_OP_423J2_125_3477_n922, DP_OP_423J2_125_3477_n921,
         DP_OP_423J2_125_3477_n920, DP_OP_423J2_125_3477_n919,
         DP_OP_423J2_125_3477_n918, DP_OP_423J2_125_3477_n917,
         DP_OP_423J2_125_3477_n916, DP_OP_423J2_125_3477_n915,
         DP_OP_423J2_125_3477_n914, DP_OP_423J2_125_3477_n913,
         DP_OP_423J2_125_3477_n912, DP_OP_423J2_125_3477_n911,
         DP_OP_423J2_125_3477_n910, DP_OP_423J2_125_3477_n909,
         DP_OP_423J2_125_3477_n908, DP_OP_423J2_125_3477_n907,
         DP_OP_423J2_125_3477_n906, DP_OP_423J2_125_3477_n905,
         DP_OP_423J2_125_3477_n904, DP_OP_423J2_125_3477_n903,
         DP_OP_423J2_125_3477_n902, DP_OP_423J2_125_3477_n901,
         DP_OP_423J2_125_3477_n900, DP_OP_423J2_125_3477_n899,
         DP_OP_423J2_125_3477_n898, DP_OP_423J2_125_3477_n897,
         DP_OP_423J2_125_3477_n896, DP_OP_423J2_125_3477_n895,
         DP_OP_423J2_125_3477_n894, DP_OP_423J2_125_3477_n893,
         DP_OP_423J2_125_3477_n892, DP_OP_423J2_125_3477_n891,
         DP_OP_423J2_125_3477_n890, DP_OP_423J2_125_3477_n889,
         DP_OP_423J2_125_3477_n888, DP_OP_423J2_125_3477_n887,
         DP_OP_423J2_125_3477_n886, DP_OP_423J2_125_3477_n885,
         DP_OP_423J2_125_3477_n884, DP_OP_423J2_125_3477_n883,
         DP_OP_423J2_125_3477_n882, DP_OP_423J2_125_3477_n881,
         DP_OP_423J2_125_3477_n880, DP_OP_423J2_125_3477_n879,
         DP_OP_423J2_125_3477_n878, DP_OP_423J2_125_3477_n877,
         DP_OP_423J2_125_3477_n876, DP_OP_423J2_125_3477_n875,
         DP_OP_423J2_125_3477_n874, DP_OP_423J2_125_3477_n873,
         DP_OP_423J2_125_3477_n872, DP_OP_423J2_125_3477_n871,
         DP_OP_423J2_125_3477_n870, DP_OP_423J2_125_3477_n869,
         DP_OP_423J2_125_3477_n868, DP_OP_423J2_125_3477_n867,
         DP_OP_423J2_125_3477_n866, DP_OP_423J2_125_3477_n865,
         DP_OP_423J2_125_3477_n864, DP_OP_423J2_125_3477_n863,
         DP_OP_423J2_125_3477_n862, DP_OP_423J2_125_3477_n861,
         DP_OP_423J2_125_3477_n860, DP_OP_423J2_125_3477_n859,
         DP_OP_423J2_125_3477_n858, DP_OP_423J2_125_3477_n857,
         DP_OP_423J2_125_3477_n856, DP_OP_423J2_125_3477_n855,
         DP_OP_423J2_125_3477_n854, DP_OP_423J2_125_3477_n853,
         DP_OP_423J2_125_3477_n852, DP_OP_423J2_125_3477_n851,
         DP_OP_423J2_125_3477_n850, DP_OP_423J2_125_3477_n849,
         DP_OP_423J2_125_3477_n848, DP_OP_423J2_125_3477_n847,
         DP_OP_423J2_125_3477_n846, DP_OP_423J2_125_3477_n845,
         DP_OP_423J2_125_3477_n844, DP_OP_423J2_125_3477_n843,
         DP_OP_423J2_125_3477_n842, DP_OP_423J2_125_3477_n841,
         DP_OP_423J2_125_3477_n840, DP_OP_423J2_125_3477_n839,
         DP_OP_423J2_125_3477_n838, DP_OP_423J2_125_3477_n837,
         DP_OP_423J2_125_3477_n836, DP_OP_423J2_125_3477_n835,
         DP_OP_423J2_125_3477_n834, DP_OP_423J2_125_3477_n833,
         DP_OP_423J2_125_3477_n832, DP_OP_423J2_125_3477_n831,
         DP_OP_423J2_125_3477_n830, DP_OP_423J2_125_3477_n829,
         DP_OP_423J2_125_3477_n828, DP_OP_423J2_125_3477_n827,
         DP_OP_423J2_125_3477_n826, DP_OP_423J2_125_3477_n825,
         DP_OP_423J2_125_3477_n824, DP_OP_423J2_125_3477_n823,
         DP_OP_423J2_125_3477_n822, DP_OP_423J2_125_3477_n821,
         DP_OP_423J2_125_3477_n820, DP_OP_423J2_125_3477_n819,
         DP_OP_423J2_125_3477_n818, DP_OP_423J2_125_3477_n817,
         DP_OP_423J2_125_3477_n816, DP_OP_423J2_125_3477_n815,
         DP_OP_423J2_125_3477_n814, DP_OP_423J2_125_3477_n813,
         DP_OP_423J2_125_3477_n812, DP_OP_423J2_125_3477_n811,
         DP_OP_423J2_125_3477_n810, DP_OP_423J2_125_3477_n809,
         DP_OP_423J2_125_3477_n808, DP_OP_423J2_125_3477_n807,
         DP_OP_423J2_125_3477_n806, DP_OP_423J2_125_3477_n805,
         DP_OP_423J2_125_3477_n804, DP_OP_423J2_125_3477_n803,
         DP_OP_423J2_125_3477_n802, DP_OP_423J2_125_3477_n801,
         DP_OP_423J2_125_3477_n800, DP_OP_423J2_125_3477_n799,
         DP_OP_423J2_125_3477_n798, DP_OP_423J2_125_3477_n797,
         DP_OP_423J2_125_3477_n796, DP_OP_423J2_125_3477_n795,
         DP_OP_423J2_125_3477_n794, DP_OP_423J2_125_3477_n793,
         DP_OP_423J2_125_3477_n792, DP_OP_423J2_125_3477_n791,
         DP_OP_423J2_125_3477_n790, DP_OP_423J2_125_3477_n789,
         DP_OP_423J2_125_3477_n788, DP_OP_423J2_125_3477_n787,
         DP_OP_423J2_125_3477_n786, DP_OP_423J2_125_3477_n785,
         DP_OP_423J2_125_3477_n784, DP_OP_423J2_125_3477_n783,
         DP_OP_423J2_125_3477_n782, DP_OP_423J2_125_3477_n781,
         DP_OP_423J2_125_3477_n780, DP_OP_423J2_125_3477_n779,
         DP_OP_423J2_125_3477_n778, DP_OP_423J2_125_3477_n777,
         DP_OP_423J2_125_3477_n776, DP_OP_423J2_125_3477_n775,
         DP_OP_423J2_125_3477_n774, DP_OP_423J2_125_3477_n773,
         DP_OP_423J2_125_3477_n772, DP_OP_423J2_125_3477_n771,
         DP_OP_423J2_125_3477_n770, DP_OP_423J2_125_3477_n769,
         DP_OP_423J2_125_3477_n768, DP_OP_423J2_125_3477_n767,
         DP_OP_423J2_125_3477_n766, DP_OP_423J2_125_3477_n765,
         DP_OP_423J2_125_3477_n764, DP_OP_423J2_125_3477_n763,
         DP_OP_423J2_125_3477_n762, DP_OP_423J2_125_3477_n761,
         DP_OP_423J2_125_3477_n760, DP_OP_423J2_125_3477_n759,
         DP_OP_423J2_125_3477_n758, DP_OP_423J2_125_3477_n757,
         DP_OP_423J2_125_3477_n756, DP_OP_423J2_125_3477_n755,
         DP_OP_423J2_125_3477_n754, DP_OP_423J2_125_3477_n753,
         DP_OP_423J2_125_3477_n752, DP_OP_423J2_125_3477_n751,
         DP_OP_423J2_125_3477_n750, DP_OP_423J2_125_3477_n749,
         DP_OP_423J2_125_3477_n748, DP_OP_423J2_125_3477_n747,
         DP_OP_423J2_125_3477_n746, DP_OP_423J2_125_3477_n745,
         DP_OP_423J2_125_3477_n744, DP_OP_423J2_125_3477_n743,
         DP_OP_423J2_125_3477_n742, DP_OP_423J2_125_3477_n741,
         DP_OP_423J2_125_3477_n740, DP_OP_423J2_125_3477_n739,
         DP_OP_423J2_125_3477_n738, DP_OP_423J2_125_3477_n737,
         DP_OP_423J2_125_3477_n736, DP_OP_423J2_125_3477_n735,
         DP_OP_423J2_125_3477_n734, DP_OP_423J2_125_3477_n733,
         DP_OP_423J2_125_3477_n732, DP_OP_423J2_125_3477_n731,
         DP_OP_423J2_125_3477_n730, DP_OP_423J2_125_3477_n729,
         DP_OP_423J2_125_3477_n728, DP_OP_423J2_125_3477_n727,
         DP_OP_423J2_125_3477_n726, DP_OP_423J2_125_3477_n725,
         DP_OP_423J2_125_3477_n724, DP_OP_423J2_125_3477_n723,
         DP_OP_423J2_125_3477_n722, DP_OP_423J2_125_3477_n721,
         DP_OP_423J2_125_3477_n720, DP_OP_423J2_125_3477_n719,
         DP_OP_423J2_125_3477_n718, DP_OP_423J2_125_3477_n717,
         DP_OP_423J2_125_3477_n716, DP_OP_423J2_125_3477_n715,
         DP_OP_423J2_125_3477_n714, DP_OP_423J2_125_3477_n713,
         DP_OP_423J2_125_3477_n712, DP_OP_423J2_125_3477_n711,
         DP_OP_423J2_125_3477_n710, DP_OP_423J2_125_3477_n709,
         DP_OP_423J2_125_3477_n708, DP_OP_423J2_125_3477_n707,
         DP_OP_423J2_125_3477_n706, DP_OP_423J2_125_3477_n705,
         DP_OP_423J2_125_3477_n704, DP_OP_423J2_125_3477_n703,
         DP_OP_423J2_125_3477_n702, DP_OP_423J2_125_3477_n701,
         DP_OP_423J2_125_3477_n700, DP_OP_423J2_125_3477_n699,
         DP_OP_423J2_125_3477_n698, DP_OP_423J2_125_3477_n697,
         DP_OP_423J2_125_3477_n696, DP_OP_423J2_125_3477_n695,
         DP_OP_423J2_125_3477_n694, DP_OP_423J2_125_3477_n693,
         DP_OP_423J2_125_3477_n692, DP_OP_423J2_125_3477_n691,
         DP_OP_423J2_125_3477_n690, DP_OP_423J2_125_3477_n689,
         DP_OP_423J2_125_3477_n688, DP_OP_423J2_125_3477_n687,
         DP_OP_423J2_125_3477_n686, DP_OP_423J2_125_3477_n685,
         DP_OP_423J2_125_3477_n684, DP_OP_423J2_125_3477_n683,
         DP_OP_423J2_125_3477_n682, DP_OP_423J2_125_3477_n681,
         DP_OP_423J2_125_3477_n680, DP_OP_423J2_125_3477_n679,
         DP_OP_423J2_125_3477_n678, DP_OP_423J2_125_3477_n677,
         DP_OP_423J2_125_3477_n676, DP_OP_423J2_125_3477_n675,
         DP_OP_423J2_125_3477_n674, DP_OP_423J2_125_3477_n673,
         DP_OP_423J2_125_3477_n672, DP_OP_423J2_125_3477_n671,
         DP_OP_423J2_125_3477_n670, DP_OP_423J2_125_3477_n669,
         DP_OP_423J2_125_3477_n668, DP_OP_423J2_125_3477_n667,
         DP_OP_423J2_125_3477_n666, DP_OP_423J2_125_3477_n665,
         DP_OP_423J2_125_3477_n664, DP_OP_423J2_125_3477_n663,
         DP_OP_423J2_125_3477_n662, DP_OP_423J2_125_3477_n661,
         DP_OP_423J2_125_3477_n660, DP_OP_423J2_125_3477_n659,
         DP_OP_423J2_125_3477_n658, DP_OP_423J2_125_3477_n657,
         DP_OP_423J2_125_3477_n656, DP_OP_423J2_125_3477_n655,
         DP_OP_423J2_125_3477_n654, DP_OP_423J2_125_3477_n653,
         DP_OP_423J2_125_3477_n652, DP_OP_423J2_125_3477_n651,
         DP_OP_423J2_125_3477_n650, DP_OP_423J2_125_3477_n649,
         DP_OP_423J2_125_3477_n648, DP_OP_423J2_125_3477_n647,
         DP_OP_423J2_125_3477_n646, DP_OP_423J2_125_3477_n645,
         DP_OP_423J2_125_3477_n644, DP_OP_423J2_125_3477_n643,
         DP_OP_423J2_125_3477_n642, DP_OP_423J2_125_3477_n641,
         DP_OP_423J2_125_3477_n640, DP_OP_423J2_125_3477_n639,
         DP_OP_423J2_125_3477_n638, DP_OP_423J2_125_3477_n637,
         DP_OP_423J2_125_3477_n636, DP_OP_423J2_125_3477_n635,
         DP_OP_423J2_125_3477_n634, DP_OP_423J2_125_3477_n633,
         DP_OP_423J2_125_3477_n632, DP_OP_423J2_125_3477_n631,
         DP_OP_423J2_125_3477_n630, DP_OP_423J2_125_3477_n629,
         DP_OP_423J2_125_3477_n628, DP_OP_423J2_125_3477_n627,
         DP_OP_423J2_125_3477_n626, DP_OP_423J2_125_3477_n625,
         DP_OP_423J2_125_3477_n624, DP_OP_423J2_125_3477_n623,
         DP_OP_423J2_125_3477_n622, DP_OP_423J2_125_3477_n621,
         DP_OP_423J2_125_3477_n620, DP_OP_423J2_125_3477_n619,
         DP_OP_423J2_125_3477_n618, DP_OP_423J2_125_3477_n617,
         DP_OP_423J2_125_3477_n616, DP_OP_423J2_125_3477_n615,
         DP_OP_423J2_125_3477_n614, DP_OP_423J2_125_3477_n613,
         DP_OP_423J2_125_3477_n612, DP_OP_423J2_125_3477_n611,
         DP_OP_423J2_125_3477_n610, DP_OP_423J2_125_3477_n609,
         DP_OP_423J2_125_3477_n608, DP_OP_423J2_125_3477_n607,
         DP_OP_423J2_125_3477_n606, DP_OP_423J2_125_3477_n605,
         DP_OP_423J2_125_3477_n604, DP_OP_423J2_125_3477_n603,
         DP_OP_423J2_125_3477_n602, DP_OP_423J2_125_3477_n601,
         DP_OP_423J2_125_3477_n600, DP_OP_423J2_125_3477_n599,
         DP_OP_423J2_125_3477_n598, DP_OP_423J2_125_3477_n597,
         DP_OP_423J2_125_3477_n596, DP_OP_423J2_125_3477_n595,
         DP_OP_423J2_125_3477_n594, DP_OP_423J2_125_3477_n593,
         DP_OP_423J2_125_3477_n592, DP_OP_423J2_125_3477_n591,
         DP_OP_423J2_125_3477_n590, DP_OP_423J2_125_3477_n589,
         DP_OP_423J2_125_3477_n588, DP_OP_423J2_125_3477_n587,
         DP_OP_423J2_125_3477_n586, DP_OP_423J2_125_3477_n585,
         DP_OP_423J2_125_3477_n584, DP_OP_423J2_125_3477_n583,
         DP_OP_423J2_125_3477_n582, DP_OP_423J2_125_3477_n581,
         DP_OP_423J2_125_3477_n580, DP_OP_423J2_125_3477_n579,
         DP_OP_423J2_125_3477_n578, DP_OP_423J2_125_3477_n577,
         DP_OP_423J2_125_3477_n576, DP_OP_423J2_125_3477_n575,
         DP_OP_423J2_125_3477_n574, DP_OP_423J2_125_3477_n573,
         DP_OP_423J2_125_3477_n572, DP_OP_423J2_125_3477_n571,
         DP_OP_423J2_125_3477_n570, DP_OP_423J2_125_3477_n569,
         DP_OP_423J2_125_3477_n568, DP_OP_423J2_125_3477_n567,
         DP_OP_423J2_125_3477_n566, DP_OP_423J2_125_3477_n565,
         DP_OP_423J2_125_3477_n564, DP_OP_423J2_125_3477_n563,
         DP_OP_423J2_125_3477_n562, DP_OP_423J2_125_3477_n561,
         DP_OP_423J2_125_3477_n560, DP_OP_423J2_125_3477_n559,
         DP_OP_423J2_125_3477_n558, DP_OP_423J2_125_3477_n557,
         DP_OP_423J2_125_3477_n556, DP_OP_423J2_125_3477_n555,
         DP_OP_423J2_125_3477_n554, DP_OP_423J2_125_3477_n553,
         DP_OP_423J2_125_3477_n552, DP_OP_423J2_125_3477_n551,
         DP_OP_423J2_125_3477_n550, DP_OP_423J2_125_3477_n549,
         DP_OP_423J2_125_3477_n548, DP_OP_423J2_125_3477_n547,
         DP_OP_423J2_125_3477_n546, DP_OP_423J2_125_3477_n545,
         DP_OP_423J2_125_3477_n544, DP_OP_423J2_125_3477_n543,
         DP_OP_423J2_125_3477_n542, DP_OP_423J2_125_3477_n541,
         DP_OP_423J2_125_3477_n540, DP_OP_423J2_125_3477_n539,
         DP_OP_423J2_125_3477_n538, DP_OP_423J2_125_3477_n537,
         DP_OP_423J2_125_3477_n536, DP_OP_423J2_125_3477_n535,
         DP_OP_423J2_125_3477_n534, DP_OP_423J2_125_3477_n533,
         DP_OP_423J2_125_3477_n532, DP_OP_423J2_125_3477_n531,
         DP_OP_423J2_125_3477_n530, DP_OP_423J2_125_3477_n529,
         DP_OP_423J2_125_3477_n528, DP_OP_423J2_125_3477_n527,
         DP_OP_423J2_125_3477_n526, DP_OP_423J2_125_3477_n525,
         DP_OP_423J2_125_3477_n524, DP_OP_423J2_125_3477_n523,
         DP_OP_423J2_125_3477_n522, DP_OP_423J2_125_3477_n521,
         DP_OP_423J2_125_3477_n520, DP_OP_423J2_125_3477_n519,
         DP_OP_423J2_125_3477_n518, DP_OP_423J2_125_3477_n517,
         DP_OP_423J2_125_3477_n516, DP_OP_423J2_125_3477_n515,
         DP_OP_423J2_125_3477_n514, DP_OP_423J2_125_3477_n513,
         DP_OP_423J2_125_3477_n512, DP_OP_423J2_125_3477_n511,
         DP_OP_423J2_125_3477_n510, DP_OP_423J2_125_3477_n509,
         DP_OP_423J2_125_3477_n508, DP_OP_423J2_125_3477_n507,
         DP_OP_423J2_125_3477_n506, DP_OP_423J2_125_3477_n505,
         DP_OP_423J2_125_3477_n504, DP_OP_423J2_125_3477_n503,
         DP_OP_423J2_125_3477_n502, DP_OP_423J2_125_3477_n501,
         DP_OP_423J2_125_3477_n500, DP_OP_423J2_125_3477_n499,
         DP_OP_423J2_125_3477_n498, DP_OP_423J2_125_3477_n497,
         DP_OP_423J2_125_3477_n496, DP_OP_423J2_125_3477_n495,
         DP_OP_423J2_125_3477_n494, DP_OP_423J2_125_3477_n493,
         DP_OP_423J2_125_3477_n492, DP_OP_423J2_125_3477_n491,
         DP_OP_423J2_125_3477_n490, DP_OP_423J2_125_3477_n489,
         DP_OP_423J2_125_3477_n488, DP_OP_423J2_125_3477_n487,
         DP_OP_423J2_125_3477_n486, DP_OP_423J2_125_3477_n485,
         DP_OP_423J2_125_3477_n484, DP_OP_423J2_125_3477_n483,
         DP_OP_423J2_125_3477_n482, DP_OP_423J2_125_3477_n481,
         DP_OP_423J2_125_3477_n480, DP_OP_423J2_125_3477_n479,
         DP_OP_423J2_125_3477_n478, DP_OP_423J2_125_3477_n477,
         DP_OP_423J2_125_3477_n476, DP_OP_423J2_125_3477_n475,
         DP_OP_423J2_125_3477_n474, DP_OP_423J2_125_3477_n473,
         DP_OP_423J2_125_3477_n472, DP_OP_423J2_125_3477_n471,
         DP_OP_423J2_125_3477_n470, DP_OP_423J2_125_3477_n469,
         DP_OP_423J2_125_3477_n468, DP_OP_423J2_125_3477_n467,
         DP_OP_423J2_125_3477_n466, DP_OP_423J2_125_3477_n465,
         DP_OP_423J2_125_3477_n464, DP_OP_423J2_125_3477_n463,
         DP_OP_423J2_125_3477_n462, DP_OP_423J2_125_3477_n461,
         DP_OP_423J2_125_3477_n460, DP_OP_423J2_125_3477_n459,
         DP_OP_423J2_125_3477_n458, DP_OP_423J2_125_3477_n457,
         DP_OP_423J2_125_3477_n456, DP_OP_423J2_125_3477_n455,
         DP_OP_423J2_125_3477_n454, DP_OP_423J2_125_3477_n453,
         DP_OP_423J2_125_3477_n452, DP_OP_423J2_125_3477_n451,
         DP_OP_423J2_125_3477_n450, DP_OP_423J2_125_3477_n449,
         DP_OP_423J2_125_3477_n448, DP_OP_423J2_125_3477_n447,
         DP_OP_423J2_125_3477_n446, DP_OP_423J2_125_3477_n445,
         DP_OP_423J2_125_3477_n444, DP_OP_423J2_125_3477_n443,
         DP_OP_423J2_125_3477_n442, DP_OP_423J2_125_3477_n441,
         DP_OP_423J2_125_3477_n440, DP_OP_423J2_125_3477_n439,
         DP_OP_423J2_125_3477_n438, DP_OP_423J2_125_3477_n437,
         DP_OP_423J2_125_3477_n436, DP_OP_423J2_125_3477_n435,
         DP_OP_423J2_125_3477_n434, DP_OP_423J2_125_3477_n433,
         DP_OP_423J2_125_3477_n432, DP_OP_423J2_125_3477_n431,
         DP_OP_423J2_125_3477_n430, DP_OP_423J2_125_3477_n429,
         DP_OP_423J2_125_3477_n428, DP_OP_423J2_125_3477_n427,
         DP_OP_423J2_125_3477_n426, DP_OP_423J2_125_3477_n425,
         DP_OP_423J2_125_3477_n424, DP_OP_423J2_125_3477_n423,
         DP_OP_423J2_125_3477_n422, DP_OP_423J2_125_3477_n421,
         DP_OP_423J2_125_3477_n420, DP_OP_423J2_125_3477_n419,
         DP_OP_423J2_125_3477_n418, DP_OP_423J2_125_3477_n417,
         DP_OP_423J2_125_3477_n416, DP_OP_423J2_125_3477_n415,
         DP_OP_423J2_125_3477_n414, DP_OP_423J2_125_3477_n413,
         DP_OP_423J2_125_3477_n412, DP_OP_423J2_125_3477_n411,
         DP_OP_423J2_125_3477_n410, DP_OP_423J2_125_3477_n409,
         DP_OP_423J2_125_3477_n408, DP_OP_423J2_125_3477_n407,
         DP_OP_423J2_125_3477_n406, DP_OP_423J2_125_3477_n405,
         DP_OP_423J2_125_3477_n404, DP_OP_423J2_125_3477_n403,
         DP_OP_423J2_125_3477_n402, DP_OP_423J2_125_3477_n401,
         DP_OP_423J2_125_3477_n400, DP_OP_423J2_125_3477_n399,
         DP_OP_423J2_125_3477_n398, DP_OP_423J2_125_3477_n397,
         DP_OP_423J2_125_3477_n396, DP_OP_423J2_125_3477_n395,
         DP_OP_423J2_125_3477_n394, DP_OP_423J2_125_3477_n393,
         DP_OP_423J2_125_3477_n392, DP_OP_423J2_125_3477_n391,
         DP_OP_423J2_125_3477_n390, DP_OP_423J2_125_3477_n389,
         DP_OP_423J2_125_3477_n388, DP_OP_423J2_125_3477_n387,
         DP_OP_423J2_125_3477_n386, DP_OP_423J2_125_3477_n385,
         DP_OP_423J2_125_3477_n384, DP_OP_423J2_125_3477_n383,
         DP_OP_423J2_125_3477_n382, DP_OP_423J2_125_3477_n381,
         DP_OP_423J2_125_3477_n380, DP_OP_423J2_125_3477_n379,
         DP_OP_423J2_125_3477_n378, DP_OP_423J2_125_3477_n377,
         DP_OP_423J2_125_3477_n376, DP_OP_423J2_125_3477_n375,
         DP_OP_423J2_125_3477_n374, DP_OP_423J2_125_3477_n373,
         DP_OP_423J2_125_3477_n372, DP_OP_423J2_125_3477_n371,
         DP_OP_423J2_125_3477_n370, DP_OP_423J2_125_3477_n369,
         DP_OP_423J2_125_3477_n368, DP_OP_423J2_125_3477_n367,
         DP_OP_423J2_125_3477_n366, DP_OP_423J2_125_3477_n365,
         DP_OP_423J2_125_3477_n364, DP_OP_423J2_125_3477_n363,
         DP_OP_423J2_125_3477_n362, DP_OP_423J2_125_3477_n361,
         DP_OP_423J2_125_3477_n360, DP_OP_423J2_125_3477_n359,
         DP_OP_423J2_125_3477_n358, DP_OP_423J2_125_3477_n357,
         DP_OP_423J2_125_3477_n356, DP_OP_423J2_125_3477_n355,
         DP_OP_423J2_125_3477_n354, DP_OP_423J2_125_3477_n353,
         DP_OP_423J2_125_3477_n352, DP_OP_423J2_125_3477_n351,
         DP_OP_423J2_125_3477_n350, DP_OP_423J2_125_3477_n349,
         DP_OP_423J2_125_3477_n348, DP_OP_423J2_125_3477_n347,
         DP_OP_423J2_125_3477_n346, DP_OP_423J2_125_3477_n345,
         DP_OP_423J2_125_3477_n344, DP_OP_423J2_125_3477_n343,
         DP_OP_423J2_125_3477_n342, DP_OP_423J2_125_3477_n341,
         DP_OP_423J2_125_3477_n340, DP_OP_423J2_125_3477_n339,
         DP_OP_423J2_125_3477_n338, DP_OP_423J2_125_3477_n337,
         DP_OP_423J2_125_3477_n336, DP_OP_423J2_125_3477_n335,
         DP_OP_423J2_125_3477_n334, DP_OP_423J2_125_3477_n333,
         DP_OP_423J2_125_3477_n332, DP_OP_423J2_125_3477_n331,
         DP_OP_423J2_125_3477_n330, DP_OP_423J2_125_3477_n329,
         DP_OP_423J2_125_3477_n328, DP_OP_423J2_125_3477_n327,
         DP_OP_423J2_125_3477_n326, DP_OP_423J2_125_3477_n325,
         DP_OP_423J2_125_3477_n324, DP_OP_423J2_125_3477_n323,
         DP_OP_423J2_125_3477_n322, DP_OP_423J2_125_3477_n321,
         DP_OP_423J2_125_3477_n320, DP_OP_423J2_125_3477_n319,
         DP_OP_423J2_125_3477_n318, DP_OP_423J2_125_3477_n317,
         DP_OP_423J2_125_3477_n316, DP_OP_423J2_125_3477_n315,
         DP_OP_423J2_125_3477_n314, DP_OP_423J2_125_3477_n313,
         DP_OP_423J2_125_3477_n312, DP_OP_423J2_125_3477_n311,
         DP_OP_423J2_125_3477_n310, DP_OP_423J2_125_3477_n309,
         DP_OP_423J2_125_3477_n308, DP_OP_423J2_125_3477_n307,
         DP_OP_423J2_125_3477_n306, DP_OP_423J2_125_3477_n305,
         DP_OP_423J2_125_3477_n304, DP_OP_423J2_125_3477_n303,
         DP_OP_423J2_125_3477_n302, DP_OP_423J2_125_3477_n301,
         DP_OP_423J2_125_3477_n300, DP_OP_423J2_125_3477_n299,
         DP_OP_423J2_125_3477_n298, DP_OP_423J2_125_3477_n297,
         DP_OP_423J2_125_3477_n296, DP_OP_423J2_125_3477_n295,
         DP_OP_423J2_125_3477_n294, DP_OP_423J2_125_3477_n293,
         DP_OP_423J2_125_3477_n292, DP_OP_423J2_125_3477_n291,
         DP_OP_423J2_125_3477_n290, DP_OP_423J2_125_3477_n289,
         DP_OP_423J2_125_3477_n288, DP_OP_423J2_125_3477_n287,
         DP_OP_423J2_125_3477_n286, DP_OP_423J2_125_3477_n285,
         DP_OP_423J2_125_3477_n284, DP_OP_423J2_125_3477_n283,
         DP_OP_423J2_125_3477_n282, DP_OP_423J2_125_3477_n281,
         DP_OP_423J2_125_3477_n280, DP_OP_423J2_125_3477_n279,
         DP_OP_423J2_125_3477_n278, DP_OP_423J2_125_3477_n277,
         DP_OP_423J2_125_3477_n276, DP_OP_423J2_125_3477_n275,
         DP_OP_423J2_125_3477_n274, DP_OP_423J2_125_3477_n273,
         DP_OP_423J2_125_3477_n272, DP_OP_423J2_125_3477_n271,
         DP_OP_423J2_125_3477_n270, DP_OP_423J2_125_3477_n269,
         DP_OP_423J2_125_3477_n268, DP_OP_423J2_125_3477_n267,
         DP_OP_423J2_125_3477_n266, DP_OP_423J2_125_3477_n265,
         DP_OP_423J2_125_3477_n264, DP_OP_423J2_125_3477_n263,
         DP_OP_423J2_125_3477_n262, DP_OP_423J2_125_3477_n261,
         DP_OP_423J2_125_3477_n260, DP_OP_423J2_125_3477_n259,
         DP_OP_423J2_125_3477_n258, DP_OP_423J2_125_3477_n257,
         DP_OP_423J2_125_3477_n256, DP_OP_423J2_125_3477_n255,
         DP_OP_423J2_125_3477_n254, DP_OP_423J2_125_3477_n253,
         DP_OP_423J2_125_3477_n252, DP_OP_423J2_125_3477_n241,
         DP_OP_423J2_125_3477_n240, DP_OP_423J2_125_3477_n237,
         DP_OP_423J2_125_3477_n236, DP_OP_423J2_125_3477_n235,
         DP_OP_423J2_125_3477_n234, DP_OP_423J2_125_3477_n233,
         DP_OP_423J2_125_3477_n231, DP_OP_423J2_125_3477_n229,
         DP_OP_423J2_125_3477_n227, DP_OP_423J2_125_3477_n219,
         DP_OP_423J2_125_3477_n218, DP_OP_423J2_125_3477_n217,
         DP_OP_423J2_125_3477_n216, DP_OP_423J2_125_3477_n215,
         DP_OP_423J2_125_3477_n211, DP_OP_423J2_125_3477_n210,
         DP_OP_423J2_125_3477_n209, DP_OP_423J2_125_3477_n208,
         DP_OP_423J2_125_3477_n207, DP_OP_423J2_125_3477_n203,
         DP_OP_423J2_125_3477_n202, DP_OP_423J2_125_3477_n201,
         DP_OP_423J2_125_3477_n200, DP_OP_423J2_125_3477_n199,
         DP_OP_423J2_125_3477_n195, DP_OP_423J2_125_3477_n194,
         DP_OP_423J2_125_3477_n193, DP_OP_423J2_125_3477_n192,
         DP_OP_423J2_125_3477_n191, DP_OP_423J2_125_3477_n190,
         DP_OP_423J2_125_3477_n189, DP_OP_423J2_125_3477_n187,
         DP_OP_423J2_125_3477_n186, DP_OP_423J2_125_3477_n185,
         DP_OP_423J2_125_3477_n184, DP_OP_423J2_125_3477_n183,
         DP_OP_423J2_125_3477_n182, DP_OP_423J2_125_3477_n181,
         DP_OP_423J2_125_3477_n180, DP_OP_423J2_125_3477_n179,
         DP_OP_423J2_125_3477_n177, DP_OP_423J2_125_3477_n176,
         DP_OP_423J2_125_3477_n175, DP_OP_423J2_125_3477_n174,
         DP_OP_423J2_125_3477_n173, DP_OP_423J2_125_3477_n172,
         DP_OP_423J2_125_3477_n171, DP_OP_423J2_125_3477_n170,
         DP_OP_423J2_125_3477_n168, DP_OP_423J2_125_3477_n167,
         DP_OP_423J2_125_3477_n166, DP_OP_423J2_125_3477_n165,
         DP_OP_423J2_125_3477_n164, DP_OP_423J2_125_3477_n163,
         DP_OP_423J2_125_3477_n162, DP_OP_423J2_125_3477_n161,
         DP_OP_423J2_125_3477_n158, DP_OP_423J2_125_3477_n152,
         DP_OP_423J2_125_3477_n151, DP_OP_423J2_125_3477_n149,
         DP_OP_423J2_125_3477_n148, DP_OP_423J2_125_3477_n145,
         DP_OP_423J2_125_3477_n144, DP_OP_423J2_125_3477_n141,
         DP_OP_423J2_125_3477_n140, DP_OP_423J2_125_3477_n137,
         DP_OP_423J2_125_3477_n136, DP_OP_423J2_125_3477_n135,
         DP_OP_423J2_125_3477_n133, DP_OP_423J2_125_3477_n132,
         DP_OP_423J2_125_3477_n131, DP_OP_423J2_125_3477_n130,
         DP_OP_423J2_125_3477_n129, DP_OP_423J2_125_3477_n128,
         DP_OP_423J2_125_3477_n127, DP_OP_423J2_125_3477_n126,
         DP_OP_423J2_125_3477_n125, DP_OP_423J2_125_3477_n124,
         DP_OP_423J2_125_3477_n123, DP_OP_423J2_125_3477_n119,
         DP_OP_423J2_125_3477_n118, DP_OP_423J2_125_3477_n116,
         DP_OP_423J2_125_3477_n115, DP_OP_423J2_125_3477_n114,
         DP_OP_423J2_125_3477_n113, DP_OP_423J2_125_3477_n112,
         DP_OP_423J2_125_3477_n111, DP_OP_423J2_125_3477_n109,
         DP_OP_423J2_125_3477_n105, DP_OP_423J2_125_3477_n104,
         DP_OP_423J2_125_3477_n102, DP_OP_423J2_125_3477_n101,
         DP_OP_423J2_125_3477_n100, DP_OP_423J2_125_3477_n99,
         DP_OP_423J2_125_3477_n98, DP_OP_423J2_125_3477_n97,
         DP_OP_423J2_125_3477_n95, DP_OP_423J2_125_3477_n91,
         DP_OP_423J2_125_3477_n90, DP_OP_423J2_125_3477_n88,
         DP_OP_423J2_125_3477_n87, DP_OP_423J2_125_3477_n86,
         DP_OP_423J2_125_3477_n85, DP_OP_423J2_125_3477_n84,
         DP_OP_423J2_125_3477_n83, DP_OP_423J2_125_3477_n81,
         DP_OP_423J2_125_3477_n76, DP_OP_423J2_125_3477_n75,
         DP_OP_423J2_125_3477_n74, DP_OP_423J2_125_3477_n73,
         DP_OP_423J2_125_3477_n72, DP_OP_423J2_125_3477_n70,
         DP_OP_423J2_125_3477_n65, DP_OP_423J2_125_3477_n63,
         DP_OP_423J2_125_3477_n62, DP_OP_423J2_125_3477_n61,
         DP_OP_423J2_125_3477_n59, DP_OP_423J2_125_3477_n58,
         DP_OP_423J2_125_3477_n57, DP_OP_423J2_125_3477_n56,
         DP_OP_423J2_125_3477_n55, DP_OP_423J2_125_3477_n52,
         DP_OP_423J2_125_3477_n48, DP_OP_423J2_125_3477_n47,
         DP_OP_423J2_125_3477_n45, DP_OP_423J2_125_3477_n44,
         DP_OP_423J2_125_3477_n43, DP_OP_423J2_125_3477_n42,
         DP_OP_423J2_125_3477_n41, DP_OP_423J2_125_3477_n40,
         DP_OP_423J2_125_3477_n39, DP_OP_423J2_125_3477_n37,
         DP_OP_423J2_125_3477_n25, DP_OP_423J2_125_3477_n20,
         DP_OP_423J2_125_3477_n19, DP_OP_423J2_125_3477_n18,
         DP_OP_423J2_125_3477_n17, DP_OP_423J2_125_3477_n4,
         DP_OP_423J2_125_3477_n3, DP_OP_423J2_125_3477_n2,
         DP_OP_422J2_124_3477_n3017, DP_OP_422J2_124_3477_n3016,
         DP_OP_422J2_124_3477_n3015, DP_OP_422J2_124_3477_n3014,
         DP_OP_422J2_124_3477_n3013, DP_OP_422J2_124_3477_n3012,
         DP_OP_422J2_124_3477_n3011, DP_OP_422J2_124_3477_n3010,
         DP_OP_422J2_124_3477_n3009, DP_OP_422J2_124_3477_n3008,
         DP_OP_422J2_124_3477_n3007, DP_OP_422J2_124_3477_n3006,
         DP_OP_422J2_124_3477_n3005, DP_OP_422J2_124_3477_n3004,
         DP_OP_422J2_124_3477_n3003, DP_OP_422J2_124_3477_n3002,
         DP_OP_422J2_124_3477_n3001, DP_OP_422J2_124_3477_n3000,
         DP_OP_422J2_124_3477_n2999, DP_OP_422J2_124_3477_n2998,
         DP_OP_422J2_124_3477_n2997, DP_OP_422J2_124_3477_n2996,
         DP_OP_422J2_124_3477_n2995, DP_OP_422J2_124_3477_n2994,
         DP_OP_422J2_124_3477_n2993, DP_OP_422J2_124_3477_n2992,
         DP_OP_422J2_124_3477_n2991, DP_OP_422J2_124_3477_n2990,
         DP_OP_422J2_124_3477_n2989, DP_OP_422J2_124_3477_n2988,
         DP_OP_422J2_124_3477_n2987, DP_OP_422J2_124_3477_n2986,
         DP_OP_422J2_124_3477_n2985, DP_OP_422J2_124_3477_n2984,
         DP_OP_422J2_124_3477_n2983, DP_OP_422J2_124_3477_n2982,
         DP_OP_422J2_124_3477_n2981, DP_OP_422J2_124_3477_n2980,
         DP_OP_422J2_124_3477_n2979, DP_OP_422J2_124_3477_n2978,
         DP_OP_422J2_124_3477_n2977, DP_OP_422J2_124_3477_n2976,
         DP_OP_422J2_124_3477_n2975, DP_OP_422J2_124_3477_n2974,
         DP_OP_422J2_124_3477_n2973, DP_OP_422J2_124_3477_n2972,
         DP_OP_422J2_124_3477_n2971, DP_OP_422J2_124_3477_n2970,
         DP_OP_422J2_124_3477_n2969, DP_OP_422J2_124_3477_n2964,
         DP_OP_422J2_124_3477_n2963, DP_OP_422J2_124_3477_n2962,
         DP_OP_422J2_124_3477_n2961, DP_OP_422J2_124_3477_n2960,
         DP_OP_422J2_124_3477_n2959, DP_OP_422J2_124_3477_n2958,
         DP_OP_422J2_124_3477_n2957, DP_OP_422J2_124_3477_n2956,
         DP_OP_422J2_124_3477_n2955, DP_OP_422J2_124_3477_n2954,
         DP_OP_422J2_124_3477_n2953, DP_OP_422J2_124_3477_n2952,
         DP_OP_422J2_124_3477_n2951, DP_OP_422J2_124_3477_n2950,
         DP_OP_422J2_124_3477_n2949, DP_OP_422J2_124_3477_n2948,
         DP_OP_422J2_124_3477_n2947, DP_OP_422J2_124_3477_n2946,
         DP_OP_422J2_124_3477_n2945, DP_OP_422J2_124_3477_n2944,
         DP_OP_422J2_124_3477_n2943, DP_OP_422J2_124_3477_n2942,
         DP_OP_422J2_124_3477_n2941, DP_OP_422J2_124_3477_n2940,
         DP_OP_422J2_124_3477_n2939, DP_OP_422J2_124_3477_n2938,
         DP_OP_422J2_124_3477_n2937, DP_OP_422J2_124_3477_n2936,
         DP_OP_422J2_124_3477_n2935, DP_OP_422J2_124_3477_n2934,
         DP_OP_422J2_124_3477_n2933, DP_OP_422J2_124_3477_n2932,
         DP_OP_422J2_124_3477_n2931, DP_OP_422J2_124_3477_n2930,
         DP_OP_422J2_124_3477_n2929, DP_OP_422J2_124_3477_n2928,
         DP_OP_422J2_124_3477_n2927, DP_OP_422J2_124_3477_n2926,
         DP_OP_422J2_124_3477_n2924, DP_OP_422J2_124_3477_n2923,
         DP_OP_422J2_124_3477_n2922, DP_OP_422J2_124_3477_n2921,
         DP_OP_422J2_124_3477_n2919, DP_OP_422J2_124_3477_n2918,
         DP_OP_422J2_124_3477_n2917, DP_OP_422J2_124_3477_n2916,
         DP_OP_422J2_124_3477_n2915, DP_OP_422J2_124_3477_n2914,
         DP_OP_422J2_124_3477_n2913, DP_OP_422J2_124_3477_n2912,
         DP_OP_422J2_124_3477_n2911, DP_OP_422J2_124_3477_n2910,
         DP_OP_422J2_124_3477_n2909, DP_OP_422J2_124_3477_n2908,
         DP_OP_422J2_124_3477_n2907, DP_OP_422J2_124_3477_n2906,
         DP_OP_422J2_124_3477_n2905, DP_OP_422J2_124_3477_n2904,
         DP_OP_422J2_124_3477_n2903, DP_OP_422J2_124_3477_n2902,
         DP_OP_422J2_124_3477_n2901, DP_OP_422J2_124_3477_n2900,
         DP_OP_422J2_124_3477_n2899, DP_OP_422J2_124_3477_n2898,
         DP_OP_422J2_124_3477_n2897, DP_OP_422J2_124_3477_n2896,
         DP_OP_422J2_124_3477_n2895, DP_OP_422J2_124_3477_n2894,
         DP_OP_422J2_124_3477_n2893, DP_OP_422J2_124_3477_n2892,
         DP_OP_422J2_124_3477_n2891, DP_OP_422J2_124_3477_n2890,
         DP_OP_422J2_124_3477_n2889, DP_OP_422J2_124_3477_n2888,
         DP_OP_422J2_124_3477_n2887, DP_OP_422J2_124_3477_n2886,
         DP_OP_422J2_124_3477_n2885, DP_OP_422J2_124_3477_n2884,
         DP_OP_422J2_124_3477_n2883, DP_OP_422J2_124_3477_n2880,
         DP_OP_422J2_124_3477_n2878, DP_OP_422J2_124_3477_n2877,
         DP_OP_422J2_124_3477_n2875, DP_OP_422J2_124_3477_n2874,
         DP_OP_422J2_124_3477_n2873, DP_OP_422J2_124_3477_n2872,
         DP_OP_422J2_124_3477_n2871, DP_OP_422J2_124_3477_n2870,
         DP_OP_422J2_124_3477_n2869, DP_OP_422J2_124_3477_n2868,
         DP_OP_422J2_124_3477_n2867, DP_OP_422J2_124_3477_n2866,
         DP_OP_422J2_124_3477_n2865, DP_OP_422J2_124_3477_n2864,
         DP_OP_422J2_124_3477_n2863, DP_OP_422J2_124_3477_n2862,
         DP_OP_422J2_124_3477_n2861, DP_OP_422J2_124_3477_n2860,
         DP_OP_422J2_124_3477_n2859, DP_OP_422J2_124_3477_n2858,
         DP_OP_422J2_124_3477_n2857, DP_OP_422J2_124_3477_n2856,
         DP_OP_422J2_124_3477_n2855, DP_OP_422J2_124_3477_n2854,
         DP_OP_422J2_124_3477_n2853, DP_OP_422J2_124_3477_n2852,
         DP_OP_422J2_124_3477_n2851, DP_OP_422J2_124_3477_n2850,
         DP_OP_422J2_124_3477_n2849, DP_OP_422J2_124_3477_n2848,
         DP_OP_422J2_124_3477_n2847, DP_OP_422J2_124_3477_n2846,
         DP_OP_422J2_124_3477_n2845, DP_OP_422J2_124_3477_n2844,
         DP_OP_422J2_124_3477_n2843, DP_OP_422J2_124_3477_n2842,
         DP_OP_422J2_124_3477_n2841, DP_OP_422J2_124_3477_n2840,
         DP_OP_422J2_124_3477_n2838, DP_OP_422J2_124_3477_n2837,
         DP_OP_422J2_124_3477_n2835, DP_OP_422J2_124_3477_n2834,
         DP_OP_422J2_124_3477_n2833, DP_OP_422J2_124_3477_n2831,
         DP_OP_422J2_124_3477_n2830, DP_OP_422J2_124_3477_n2829,
         DP_OP_422J2_124_3477_n2828, DP_OP_422J2_124_3477_n2827,
         DP_OP_422J2_124_3477_n2826, DP_OP_422J2_124_3477_n2825,
         DP_OP_422J2_124_3477_n2824, DP_OP_422J2_124_3477_n2823,
         DP_OP_422J2_124_3477_n2822, DP_OP_422J2_124_3477_n2821,
         DP_OP_422J2_124_3477_n2820, DP_OP_422J2_124_3477_n2819,
         DP_OP_422J2_124_3477_n2818, DP_OP_422J2_124_3477_n2817,
         DP_OP_422J2_124_3477_n2816, DP_OP_422J2_124_3477_n2815,
         DP_OP_422J2_124_3477_n2814, DP_OP_422J2_124_3477_n2813,
         DP_OP_422J2_124_3477_n2812, DP_OP_422J2_124_3477_n2811,
         DP_OP_422J2_124_3477_n2810, DP_OP_422J2_124_3477_n2809,
         DP_OP_422J2_124_3477_n2808, DP_OP_422J2_124_3477_n2807,
         DP_OP_422J2_124_3477_n2806, DP_OP_422J2_124_3477_n2805,
         DP_OP_422J2_124_3477_n2804, DP_OP_422J2_124_3477_n2803,
         DP_OP_422J2_124_3477_n2802, DP_OP_422J2_124_3477_n2801,
         DP_OP_422J2_124_3477_n2800, DP_OP_422J2_124_3477_n2799,
         DP_OP_422J2_124_3477_n2798, DP_OP_422J2_124_3477_n2797,
         DP_OP_422J2_124_3477_n2796, DP_OP_422J2_124_3477_n2795,
         DP_OP_422J2_124_3477_n2793, DP_OP_422J2_124_3477_n2792,
         DP_OP_422J2_124_3477_n2791, DP_OP_422J2_124_3477_n2790,
         DP_OP_422J2_124_3477_n2789, DP_OP_422J2_124_3477_n2787,
         DP_OP_422J2_124_3477_n2786, DP_OP_422J2_124_3477_n2785,
         DP_OP_422J2_124_3477_n2784, DP_OP_422J2_124_3477_n2783,
         DP_OP_422J2_124_3477_n2782, DP_OP_422J2_124_3477_n2781,
         DP_OP_422J2_124_3477_n2780, DP_OP_422J2_124_3477_n2779,
         DP_OP_422J2_124_3477_n2778, DP_OP_422J2_124_3477_n2777,
         DP_OP_422J2_124_3477_n2776, DP_OP_422J2_124_3477_n2775,
         DP_OP_422J2_124_3477_n2774, DP_OP_422J2_124_3477_n2773,
         DP_OP_422J2_124_3477_n2772, DP_OP_422J2_124_3477_n2771,
         DP_OP_422J2_124_3477_n2770, DP_OP_422J2_124_3477_n2769,
         DP_OP_422J2_124_3477_n2768, DP_OP_422J2_124_3477_n2767,
         DP_OP_422J2_124_3477_n2766, DP_OP_422J2_124_3477_n2765,
         DP_OP_422J2_124_3477_n2764, DP_OP_422J2_124_3477_n2763,
         DP_OP_422J2_124_3477_n2762, DP_OP_422J2_124_3477_n2761,
         DP_OP_422J2_124_3477_n2760, DP_OP_422J2_124_3477_n2759,
         DP_OP_422J2_124_3477_n2758, DP_OP_422J2_124_3477_n2757,
         DP_OP_422J2_124_3477_n2756, DP_OP_422J2_124_3477_n2755,
         DP_OP_422J2_124_3477_n2754, DP_OP_422J2_124_3477_n2753,
         DP_OP_422J2_124_3477_n2752, DP_OP_422J2_124_3477_n2751,
         DP_OP_422J2_124_3477_n2750, DP_OP_422J2_124_3477_n2749,
         DP_OP_422J2_124_3477_n2747, DP_OP_422J2_124_3477_n2746,
         DP_OP_422J2_124_3477_n2745, DP_OP_422J2_124_3477_n2743,
         DP_OP_422J2_124_3477_n2742, DP_OP_422J2_124_3477_n2741,
         DP_OP_422J2_124_3477_n2740, DP_OP_422J2_124_3477_n2739,
         DP_OP_422J2_124_3477_n2738, DP_OP_422J2_124_3477_n2737,
         DP_OP_422J2_124_3477_n2736, DP_OP_422J2_124_3477_n2735,
         DP_OP_422J2_124_3477_n2734, DP_OP_422J2_124_3477_n2733,
         DP_OP_422J2_124_3477_n2732, DP_OP_422J2_124_3477_n2731,
         DP_OP_422J2_124_3477_n2730, DP_OP_422J2_124_3477_n2729,
         DP_OP_422J2_124_3477_n2728, DP_OP_422J2_124_3477_n2727,
         DP_OP_422J2_124_3477_n2726, DP_OP_422J2_124_3477_n2725,
         DP_OP_422J2_124_3477_n2724, DP_OP_422J2_124_3477_n2723,
         DP_OP_422J2_124_3477_n2722, DP_OP_422J2_124_3477_n2721,
         DP_OP_422J2_124_3477_n2720, DP_OP_422J2_124_3477_n2719,
         DP_OP_422J2_124_3477_n2718, DP_OP_422J2_124_3477_n2717,
         DP_OP_422J2_124_3477_n2716, DP_OP_422J2_124_3477_n2715,
         DP_OP_422J2_124_3477_n2714, DP_OP_422J2_124_3477_n2713,
         DP_OP_422J2_124_3477_n2712, DP_OP_422J2_124_3477_n2711,
         DP_OP_422J2_124_3477_n2710, DP_OP_422J2_124_3477_n2709,
         DP_OP_422J2_124_3477_n2708, DP_OP_422J2_124_3477_n2707,
         DP_OP_422J2_124_3477_n2704, DP_OP_422J2_124_3477_n2702,
         DP_OP_422J2_124_3477_n2701, DP_OP_422J2_124_3477_n2700,
         DP_OP_422J2_124_3477_n2699, DP_OP_422J2_124_3477_n2698,
         DP_OP_422J2_124_3477_n2697, DP_OP_422J2_124_3477_n2696,
         DP_OP_422J2_124_3477_n2695, DP_OP_422J2_124_3477_n2694,
         DP_OP_422J2_124_3477_n2693, DP_OP_422J2_124_3477_n2692,
         DP_OP_422J2_124_3477_n2691, DP_OP_422J2_124_3477_n2690,
         DP_OP_422J2_124_3477_n2689, DP_OP_422J2_124_3477_n2688,
         DP_OP_422J2_124_3477_n2687, DP_OP_422J2_124_3477_n2686,
         DP_OP_422J2_124_3477_n2685, DP_OP_422J2_124_3477_n2684,
         DP_OP_422J2_124_3477_n2683, DP_OP_422J2_124_3477_n2682,
         DP_OP_422J2_124_3477_n2681, DP_OP_422J2_124_3477_n2680,
         DP_OP_422J2_124_3477_n2679, DP_OP_422J2_124_3477_n2678,
         DP_OP_422J2_124_3477_n2677, DP_OP_422J2_124_3477_n2676,
         DP_OP_422J2_124_3477_n2675, DP_OP_422J2_124_3477_n2674,
         DP_OP_422J2_124_3477_n2673, DP_OP_422J2_124_3477_n2672,
         DP_OP_422J2_124_3477_n2671, DP_OP_422J2_124_3477_n2670,
         DP_OP_422J2_124_3477_n2669, DP_OP_422J2_124_3477_n2668,
         DP_OP_422J2_124_3477_n2667, DP_OP_422J2_124_3477_n2666,
         DP_OP_422J2_124_3477_n2664, DP_OP_422J2_124_3477_n2663,
         DP_OP_422J2_124_3477_n2662, DP_OP_422J2_124_3477_n2659,
         DP_OP_422J2_124_3477_n2658, DP_OP_422J2_124_3477_n2656,
         DP_OP_422J2_124_3477_n2655, DP_OP_422J2_124_3477_n2654,
         DP_OP_422J2_124_3477_n2653, DP_OP_422J2_124_3477_n2652,
         DP_OP_422J2_124_3477_n2651, DP_OP_422J2_124_3477_n2650,
         DP_OP_422J2_124_3477_n2649, DP_OP_422J2_124_3477_n2648,
         DP_OP_422J2_124_3477_n2647, DP_OP_422J2_124_3477_n2646,
         DP_OP_422J2_124_3477_n2645, DP_OP_422J2_124_3477_n2644,
         DP_OP_422J2_124_3477_n2643, DP_OP_422J2_124_3477_n2642,
         DP_OP_422J2_124_3477_n2641, DP_OP_422J2_124_3477_n2640,
         DP_OP_422J2_124_3477_n2639, DP_OP_422J2_124_3477_n2638,
         DP_OP_422J2_124_3477_n2637, DP_OP_422J2_124_3477_n2636,
         DP_OP_422J2_124_3477_n2635, DP_OP_422J2_124_3477_n2634,
         DP_OP_422J2_124_3477_n2633, DP_OP_422J2_124_3477_n2632,
         DP_OP_422J2_124_3477_n2631, DP_OP_422J2_124_3477_n2630,
         DP_OP_422J2_124_3477_n2629, DP_OP_422J2_124_3477_n2628,
         DP_OP_422J2_124_3477_n2627, DP_OP_422J2_124_3477_n2626,
         DP_OP_422J2_124_3477_n2625, DP_OP_422J2_124_3477_n2624,
         DP_OP_422J2_124_3477_n2623, DP_OP_422J2_124_3477_n2622,
         DP_OP_422J2_124_3477_n2621, DP_OP_422J2_124_3477_n2620,
         DP_OP_422J2_124_3477_n2619, DP_OP_422J2_124_3477_n2617,
         DP_OP_422J2_124_3477_n2616, DP_OP_422J2_124_3477_n2613,
         DP_OP_422J2_124_3477_n2612, DP_OP_422J2_124_3477_n2611,
         DP_OP_422J2_124_3477_n2610, DP_OP_422J2_124_3477_n2609,
         DP_OP_422J2_124_3477_n2608, DP_OP_422J2_124_3477_n2607,
         DP_OP_422J2_124_3477_n2606, DP_OP_422J2_124_3477_n2605,
         DP_OP_422J2_124_3477_n2604, DP_OP_422J2_124_3477_n2603,
         DP_OP_422J2_124_3477_n2602, DP_OP_422J2_124_3477_n2601,
         DP_OP_422J2_124_3477_n2600, DP_OP_422J2_124_3477_n2599,
         DP_OP_422J2_124_3477_n2598, DP_OP_422J2_124_3477_n2597,
         DP_OP_422J2_124_3477_n2596, DP_OP_422J2_124_3477_n2595,
         DP_OP_422J2_124_3477_n2594, DP_OP_422J2_124_3477_n2593,
         DP_OP_422J2_124_3477_n2592, DP_OP_422J2_124_3477_n2591,
         DP_OP_422J2_124_3477_n2590, DP_OP_422J2_124_3477_n2589,
         DP_OP_422J2_124_3477_n2588, DP_OP_422J2_124_3477_n2587,
         DP_OP_422J2_124_3477_n2586, DP_OP_422J2_124_3477_n2585,
         DP_OP_422J2_124_3477_n2584, DP_OP_422J2_124_3477_n2583,
         DP_OP_422J2_124_3477_n2582, DP_OP_422J2_124_3477_n2581,
         DP_OP_422J2_124_3477_n2580, DP_OP_422J2_124_3477_n2579,
         DP_OP_422J2_124_3477_n2578, DP_OP_422J2_124_3477_n2577,
         DP_OP_422J2_124_3477_n2576, DP_OP_422J2_124_3477_n2575,
         DP_OP_422J2_124_3477_n2571, DP_OP_422J2_124_3477_n2570,
         DP_OP_422J2_124_3477_n2569, DP_OP_422J2_124_3477_n2568,
         DP_OP_422J2_124_3477_n2567, DP_OP_422J2_124_3477_n2566,
         DP_OP_422J2_124_3477_n2565, DP_OP_422J2_124_3477_n2564,
         DP_OP_422J2_124_3477_n2563, DP_OP_422J2_124_3477_n2562,
         DP_OP_422J2_124_3477_n2561, DP_OP_422J2_124_3477_n2560,
         DP_OP_422J2_124_3477_n2559, DP_OP_422J2_124_3477_n2558,
         DP_OP_422J2_124_3477_n2557, DP_OP_422J2_124_3477_n2556,
         DP_OP_422J2_124_3477_n2555, DP_OP_422J2_124_3477_n2554,
         DP_OP_422J2_124_3477_n2553, DP_OP_422J2_124_3477_n2552,
         DP_OP_422J2_124_3477_n2551, DP_OP_422J2_124_3477_n2550,
         DP_OP_422J2_124_3477_n2549, DP_OP_422J2_124_3477_n2548,
         DP_OP_422J2_124_3477_n2547, DP_OP_422J2_124_3477_n2546,
         DP_OP_422J2_124_3477_n2545, DP_OP_422J2_124_3477_n2544,
         DP_OP_422J2_124_3477_n2543, DP_OP_422J2_124_3477_n2542,
         DP_OP_422J2_124_3477_n2541, DP_OP_422J2_124_3477_n2540,
         DP_OP_422J2_124_3477_n2539, DP_OP_422J2_124_3477_n2538,
         DP_OP_422J2_124_3477_n2537, DP_OP_422J2_124_3477_n2536,
         DP_OP_422J2_124_3477_n2535, DP_OP_422J2_124_3477_n2534,
         DP_OP_422J2_124_3477_n2533, DP_OP_422J2_124_3477_n2532,
         DP_OP_422J2_124_3477_n2531, DP_OP_422J2_124_3477_n2528,
         DP_OP_422J2_124_3477_n2526, DP_OP_422J2_124_3477_n2523,
         DP_OP_422J2_124_3477_n2522, DP_OP_422J2_124_3477_n2521,
         DP_OP_422J2_124_3477_n2520, DP_OP_422J2_124_3477_n2519,
         DP_OP_422J2_124_3477_n2518, DP_OP_422J2_124_3477_n2517,
         DP_OP_422J2_124_3477_n2516, DP_OP_422J2_124_3477_n2515,
         DP_OP_422J2_124_3477_n2514, DP_OP_422J2_124_3477_n2513,
         DP_OP_422J2_124_3477_n2512, DP_OP_422J2_124_3477_n2511,
         DP_OP_422J2_124_3477_n2510, DP_OP_422J2_124_3477_n2509,
         DP_OP_422J2_124_3477_n2508, DP_OP_422J2_124_3477_n2507,
         DP_OP_422J2_124_3477_n2506, DP_OP_422J2_124_3477_n2505,
         DP_OP_422J2_124_3477_n2504, DP_OP_422J2_124_3477_n2503,
         DP_OP_422J2_124_3477_n2502, DP_OP_422J2_124_3477_n2501,
         DP_OP_422J2_124_3477_n2500, DP_OP_422J2_124_3477_n2499,
         DP_OP_422J2_124_3477_n2498, DP_OP_422J2_124_3477_n2497,
         DP_OP_422J2_124_3477_n2496, DP_OP_422J2_124_3477_n2495,
         DP_OP_422J2_124_3477_n2494, DP_OP_422J2_124_3477_n2493,
         DP_OP_422J2_124_3477_n2492, DP_OP_422J2_124_3477_n2491,
         DP_OP_422J2_124_3477_n2490, DP_OP_422J2_124_3477_n2489,
         DP_OP_422J2_124_3477_n2488, DP_OP_422J2_124_3477_n2487,
         DP_OP_422J2_124_3477_n2486, DP_OP_422J2_124_3477_n2485,
         DP_OP_422J2_124_3477_n2484, DP_OP_422J2_124_3477_n2483,
         DP_OP_422J2_124_3477_n2482, DP_OP_422J2_124_3477_n2481,
         DP_OP_422J2_124_3477_n2480, DP_OP_422J2_124_3477_n2479,
         DP_OP_422J2_124_3477_n2478, DP_OP_422J2_124_3477_n2477,
         DP_OP_422J2_124_3477_n2476, DP_OP_422J2_124_3477_n2475,
         DP_OP_422J2_124_3477_n2474, DP_OP_422J2_124_3477_n2473,
         DP_OP_422J2_124_3477_n2472, DP_OP_422J2_124_3477_n2471,
         DP_OP_422J2_124_3477_n2470, DP_OP_422J2_124_3477_n2469,
         DP_OP_422J2_124_3477_n2468, DP_OP_422J2_124_3477_n2467,
         DP_OP_422J2_124_3477_n2466, DP_OP_422J2_124_3477_n2465,
         DP_OP_422J2_124_3477_n2464, DP_OP_422J2_124_3477_n2463,
         DP_OP_422J2_124_3477_n2462, DP_OP_422J2_124_3477_n2461,
         DP_OP_422J2_124_3477_n2460, DP_OP_422J2_124_3477_n2459,
         DP_OP_422J2_124_3477_n2458, DP_OP_422J2_124_3477_n2457,
         DP_OP_422J2_124_3477_n2456, DP_OP_422J2_124_3477_n2455,
         DP_OP_422J2_124_3477_n2454, DP_OP_422J2_124_3477_n2453,
         DP_OP_422J2_124_3477_n2452, DP_OP_422J2_124_3477_n2451,
         DP_OP_422J2_124_3477_n2450, DP_OP_422J2_124_3477_n2449,
         DP_OP_422J2_124_3477_n2448, DP_OP_422J2_124_3477_n2447,
         DP_OP_422J2_124_3477_n2446, DP_OP_422J2_124_3477_n2445,
         DP_OP_422J2_124_3477_n2444, DP_OP_422J2_124_3477_n2442,
         DP_OP_422J2_124_3477_n2441, DP_OP_422J2_124_3477_n2439,
         DP_OP_422J2_124_3477_n2436, DP_OP_422J2_124_3477_n2435,
         DP_OP_422J2_124_3477_n2434, DP_OP_422J2_124_3477_n2433,
         DP_OP_422J2_124_3477_n2432, DP_OP_422J2_124_3477_n2431,
         DP_OP_422J2_124_3477_n2430, DP_OP_422J2_124_3477_n2429,
         DP_OP_422J2_124_3477_n2428, DP_OP_422J2_124_3477_n2427,
         DP_OP_422J2_124_3477_n2426, DP_OP_422J2_124_3477_n2425,
         DP_OP_422J2_124_3477_n2424, DP_OP_422J2_124_3477_n2423,
         DP_OP_422J2_124_3477_n2422, DP_OP_422J2_124_3477_n2421,
         DP_OP_422J2_124_3477_n2420, DP_OP_422J2_124_3477_n2419,
         DP_OP_422J2_124_3477_n2418, DP_OP_422J2_124_3477_n2417,
         DP_OP_422J2_124_3477_n2416, DP_OP_422J2_124_3477_n2415,
         DP_OP_422J2_124_3477_n2414, DP_OP_422J2_124_3477_n2413,
         DP_OP_422J2_124_3477_n2412, DP_OP_422J2_124_3477_n2411,
         DP_OP_422J2_124_3477_n2410, DP_OP_422J2_124_3477_n2409,
         DP_OP_422J2_124_3477_n2408, DP_OP_422J2_124_3477_n2407,
         DP_OP_422J2_124_3477_n2406, DP_OP_422J2_124_3477_n2405,
         DP_OP_422J2_124_3477_n2404, DP_OP_422J2_124_3477_n2403,
         DP_OP_422J2_124_3477_n2401, DP_OP_422J2_124_3477_n2400,
         DP_OP_422J2_124_3477_n2392, DP_OP_422J2_124_3477_n2391,
         DP_OP_422J2_124_3477_n2390, DP_OP_422J2_124_3477_n2389,
         DP_OP_422J2_124_3477_n2388, DP_OP_422J2_124_3477_n2387,
         DP_OP_422J2_124_3477_n2386, DP_OP_422J2_124_3477_n2385,
         DP_OP_422J2_124_3477_n2384, DP_OP_422J2_124_3477_n2383,
         DP_OP_422J2_124_3477_n2382, DP_OP_422J2_124_3477_n2381,
         DP_OP_422J2_124_3477_n2380, DP_OP_422J2_124_3477_n2379,
         DP_OP_422J2_124_3477_n2378, DP_OP_422J2_124_3477_n2377,
         DP_OP_422J2_124_3477_n2376, DP_OP_422J2_124_3477_n2375,
         DP_OP_422J2_124_3477_n2374, DP_OP_422J2_124_3477_n2373,
         DP_OP_422J2_124_3477_n2372, DP_OP_422J2_124_3477_n2371,
         DP_OP_422J2_124_3477_n2370, DP_OP_422J2_124_3477_n2369,
         DP_OP_422J2_124_3477_n2368, DP_OP_422J2_124_3477_n2367,
         DP_OP_422J2_124_3477_n2366, DP_OP_422J2_124_3477_n2365,
         DP_OP_422J2_124_3477_n2364, DP_OP_422J2_124_3477_n2363,
         DP_OP_422J2_124_3477_n2362, DP_OP_422J2_124_3477_n2361,
         DP_OP_422J2_124_3477_n2360, DP_OP_422J2_124_3477_n2359,
         DP_OP_422J2_124_3477_n2358, DP_OP_422J2_124_3477_n2357,
         DP_OP_422J2_124_3477_n2356, DP_OP_422J2_124_3477_n2355,
         DP_OP_422J2_124_3477_n2354, DP_OP_422J2_124_3477_n2353,
         DP_OP_422J2_124_3477_n2351, DP_OP_422J2_124_3477_n2348,
         DP_OP_422J2_124_3477_n2347, DP_OP_422J2_124_3477_n2346,
         DP_OP_422J2_124_3477_n2345, DP_OP_422J2_124_3477_n2344,
         DP_OP_422J2_124_3477_n2343, DP_OP_422J2_124_3477_n2342,
         DP_OP_422J2_124_3477_n2341, DP_OP_422J2_124_3477_n2340,
         DP_OP_422J2_124_3477_n2339, DP_OP_422J2_124_3477_n2338,
         DP_OP_422J2_124_3477_n2337, DP_OP_422J2_124_3477_n2336,
         DP_OP_422J2_124_3477_n2335, DP_OP_422J2_124_3477_n2334,
         DP_OP_422J2_124_3477_n2333, DP_OP_422J2_124_3477_n2332,
         DP_OP_422J2_124_3477_n2331, DP_OP_422J2_124_3477_n2330,
         DP_OP_422J2_124_3477_n2329, DP_OP_422J2_124_3477_n2328,
         DP_OP_422J2_124_3477_n2327, DP_OP_422J2_124_3477_n2326,
         DP_OP_422J2_124_3477_n2325, DP_OP_422J2_124_3477_n2324,
         DP_OP_422J2_124_3477_n2323, DP_OP_422J2_124_3477_n2322,
         DP_OP_422J2_124_3477_n2321, DP_OP_422J2_124_3477_n2320,
         DP_OP_422J2_124_3477_n2319, DP_OP_422J2_124_3477_n2318,
         DP_OP_422J2_124_3477_n2317, DP_OP_422J2_124_3477_n2316,
         DP_OP_422J2_124_3477_n2315, DP_OP_422J2_124_3477_n2313,
         DP_OP_422J2_124_3477_n2312, DP_OP_422J2_124_3477_n2311,
         DP_OP_422J2_124_3477_n2308, DP_OP_422J2_124_3477_n2307,
         DP_OP_422J2_124_3477_n2305, DP_OP_422J2_124_3477_n2304,
         DP_OP_422J2_124_3477_n2303, DP_OP_422J2_124_3477_n2302,
         DP_OP_422J2_124_3477_n2301, DP_OP_422J2_124_3477_n2300,
         DP_OP_422J2_124_3477_n2299, DP_OP_422J2_124_3477_n2298,
         DP_OP_422J2_124_3477_n2297, DP_OP_422J2_124_3477_n2296,
         DP_OP_422J2_124_3477_n2295, DP_OP_422J2_124_3477_n2294,
         DP_OP_422J2_124_3477_n2293, DP_OP_422J2_124_3477_n2292,
         DP_OP_422J2_124_3477_n2291, DP_OP_422J2_124_3477_n2290,
         DP_OP_422J2_124_3477_n2289, DP_OP_422J2_124_3477_n2288,
         DP_OP_422J2_124_3477_n2287, DP_OP_422J2_124_3477_n2286,
         DP_OP_422J2_124_3477_n2285, DP_OP_422J2_124_3477_n2284,
         DP_OP_422J2_124_3477_n2283, DP_OP_422J2_124_3477_n2282,
         DP_OP_422J2_124_3477_n2281, DP_OP_422J2_124_3477_n2280,
         DP_OP_422J2_124_3477_n2279, DP_OP_422J2_124_3477_n2278,
         DP_OP_422J2_124_3477_n2277, DP_OP_422J2_124_3477_n2276,
         DP_OP_422J2_124_3477_n2275, DP_OP_422J2_124_3477_n2274,
         DP_OP_422J2_124_3477_n2273, DP_OP_422J2_124_3477_n2272,
         DP_OP_422J2_124_3477_n2271, DP_OP_422J2_124_3477_n2270,
         DP_OP_422J2_124_3477_n2269, DP_OP_422J2_124_3477_n2268,
         DP_OP_422J2_124_3477_n2267, DP_OP_422J2_124_3477_n2265,
         DP_OP_422J2_124_3477_n2263, DP_OP_422J2_124_3477_n2262,
         DP_OP_422J2_124_3477_n2261, DP_OP_422J2_124_3477_n2260,
         DP_OP_422J2_124_3477_n2259, DP_OP_422J2_124_3477_n2258,
         DP_OP_422J2_124_3477_n2257, DP_OP_422J2_124_3477_n2256,
         DP_OP_422J2_124_3477_n2255, DP_OP_422J2_124_3477_n2254,
         DP_OP_422J2_124_3477_n2253, DP_OP_422J2_124_3477_n2252,
         DP_OP_422J2_124_3477_n2251, DP_OP_422J2_124_3477_n2250,
         DP_OP_422J2_124_3477_n2249, DP_OP_422J2_124_3477_n2248,
         DP_OP_422J2_124_3477_n2247, DP_OP_422J2_124_3477_n2246,
         DP_OP_422J2_124_3477_n2245, DP_OP_422J2_124_3477_n2244,
         DP_OP_422J2_124_3477_n2243, DP_OP_422J2_124_3477_n2242,
         DP_OP_422J2_124_3477_n2241, DP_OP_422J2_124_3477_n2240,
         DP_OP_422J2_124_3477_n2239, DP_OP_422J2_124_3477_n2238,
         DP_OP_422J2_124_3477_n2237, DP_OP_422J2_124_3477_n2236,
         DP_OP_422J2_124_3477_n2235, DP_OP_422J2_124_3477_n2234,
         DP_OP_422J2_124_3477_n2233, DP_OP_422J2_124_3477_n2232,
         DP_OP_422J2_124_3477_n2231, DP_OP_422J2_124_3477_n2230,
         DP_OP_422J2_124_3477_n2229, DP_OP_422J2_124_3477_n2228,
         DP_OP_422J2_124_3477_n2227, DP_OP_422J2_124_3477_n2225,
         DP_OP_422J2_124_3477_n2224, DP_OP_422J2_124_3477_n2220,
         DP_OP_422J2_124_3477_n2219, DP_OP_422J2_124_3477_n2218,
         DP_OP_422J2_124_3477_n2217, DP_OP_422J2_124_3477_n2215,
         DP_OP_422J2_124_3477_n2214, DP_OP_422J2_124_3477_n2213,
         DP_OP_422J2_124_3477_n2212, DP_OP_422J2_124_3477_n2211,
         DP_OP_422J2_124_3477_n2210, DP_OP_422J2_124_3477_n2209,
         DP_OP_422J2_124_3477_n2208, DP_OP_422J2_124_3477_n2207,
         DP_OP_422J2_124_3477_n2206, DP_OP_422J2_124_3477_n2205,
         DP_OP_422J2_124_3477_n2204, DP_OP_422J2_124_3477_n2203,
         DP_OP_422J2_124_3477_n2202, DP_OP_422J2_124_3477_n2201,
         DP_OP_422J2_124_3477_n2200, DP_OP_422J2_124_3477_n2199,
         DP_OP_422J2_124_3477_n2198, DP_OP_422J2_124_3477_n2197,
         DP_OP_422J2_124_3477_n2196, DP_OP_422J2_124_3477_n2195,
         DP_OP_422J2_124_3477_n2194, DP_OP_422J2_124_3477_n2193,
         DP_OP_422J2_124_3477_n2192, DP_OP_422J2_124_3477_n2191,
         DP_OP_422J2_124_3477_n2190, DP_OP_422J2_124_3477_n2189,
         DP_OP_422J2_124_3477_n2188, DP_OP_422J2_124_3477_n2187,
         DP_OP_422J2_124_3477_n2186, DP_OP_422J2_124_3477_n2185,
         DP_OP_422J2_124_3477_n2184, DP_OP_422J2_124_3477_n2183,
         DP_OP_422J2_124_3477_n2182, DP_OP_422J2_124_3477_n2181,
         DP_OP_422J2_124_3477_n2180, DP_OP_422J2_124_3477_n2179,
         DP_OP_422J2_124_3477_n2178, DP_OP_422J2_124_3477_n2177,
         DP_OP_422J2_124_3477_n2172, DP_OP_422J2_124_3477_n2171,
         DP_OP_422J2_124_3477_n2170, DP_OP_422J2_124_3477_n2169,
         DP_OP_422J2_124_3477_n2168, DP_OP_422J2_124_3477_n2167,
         DP_OP_422J2_124_3477_n2166, DP_OP_422J2_124_3477_n2165,
         DP_OP_422J2_124_3477_n2164, DP_OP_422J2_124_3477_n2163,
         DP_OP_422J2_124_3477_n2162, DP_OP_422J2_124_3477_n2161,
         DP_OP_422J2_124_3477_n2160, DP_OP_422J2_124_3477_n2159,
         DP_OP_422J2_124_3477_n2158, DP_OP_422J2_124_3477_n2157,
         DP_OP_422J2_124_3477_n2156, DP_OP_422J2_124_3477_n2155,
         DP_OP_422J2_124_3477_n2154, DP_OP_422J2_124_3477_n2153,
         DP_OP_422J2_124_3477_n2152, DP_OP_422J2_124_3477_n2151,
         DP_OP_422J2_124_3477_n2150, DP_OP_422J2_124_3477_n2149,
         DP_OP_422J2_124_3477_n2148, DP_OP_422J2_124_3477_n2147,
         DP_OP_422J2_124_3477_n2146, DP_OP_422J2_124_3477_n2145,
         DP_OP_422J2_124_3477_n2144, DP_OP_422J2_124_3477_n2143,
         DP_OP_422J2_124_3477_n2142, DP_OP_422J2_124_3477_n2141,
         DP_OP_422J2_124_3477_n2140, DP_OP_422J2_124_3477_n2139,
         DP_OP_422J2_124_3477_n2138, DP_OP_422J2_124_3477_n2137,
         DP_OP_422J2_124_3477_n2136, DP_OP_422J2_124_3477_n2135,
         DP_OP_422J2_124_3477_n2134, DP_OP_422J2_124_3477_n2132,
         DP_OP_422J2_124_3477_n2130, DP_OP_422J2_124_3477_n2129,
         DP_OP_422J2_124_3477_n2127, DP_OP_422J2_124_3477_n2126,
         DP_OP_422J2_124_3477_n2125, DP_OP_422J2_124_3477_n2124,
         DP_OP_422J2_124_3477_n2123, DP_OP_422J2_124_3477_n2122,
         DP_OP_422J2_124_3477_n2121, DP_OP_422J2_124_3477_n2120,
         DP_OP_422J2_124_3477_n2119, DP_OP_422J2_124_3477_n2118,
         DP_OP_422J2_124_3477_n2117, DP_OP_422J2_124_3477_n2116,
         DP_OP_422J2_124_3477_n2115, DP_OP_422J2_124_3477_n2114,
         DP_OP_422J2_124_3477_n2113, DP_OP_422J2_124_3477_n2112,
         DP_OP_422J2_124_3477_n2111, DP_OP_422J2_124_3477_n2110,
         DP_OP_422J2_124_3477_n2109, DP_OP_422J2_124_3477_n2108,
         DP_OP_422J2_124_3477_n2107, DP_OP_422J2_124_3477_n2106,
         DP_OP_422J2_124_3477_n2105, DP_OP_422J2_124_3477_n2104,
         DP_OP_422J2_124_3477_n2103, DP_OP_422J2_124_3477_n2102,
         DP_OP_422J2_124_3477_n2101, DP_OP_422J2_124_3477_n2100,
         DP_OP_422J2_124_3477_n2099, DP_OP_422J2_124_3477_n2098,
         DP_OP_422J2_124_3477_n2097, DP_OP_422J2_124_3477_n2096,
         DP_OP_422J2_124_3477_n2095, DP_OP_422J2_124_3477_n2094,
         DP_OP_422J2_124_3477_n2093, DP_OP_422J2_124_3477_n2092,
         DP_OP_422J2_124_3477_n2091, DP_OP_422J2_124_3477_n2090,
         DP_OP_422J2_124_3477_n2088, DP_OP_422J2_124_3477_n2084,
         DP_OP_422J2_124_3477_n2083, DP_OP_422J2_124_3477_n2082,
         DP_OP_422J2_124_3477_n2081, DP_OP_422J2_124_3477_n2080,
         DP_OP_422J2_124_3477_n2079, DP_OP_422J2_124_3477_n2078,
         DP_OP_422J2_124_3477_n2077, DP_OP_422J2_124_3477_n2076,
         DP_OP_422J2_124_3477_n2075, DP_OP_422J2_124_3477_n2074,
         DP_OP_422J2_124_3477_n2073, DP_OP_422J2_124_3477_n2072,
         DP_OP_422J2_124_3477_n2071, DP_OP_422J2_124_3477_n2070,
         DP_OP_422J2_124_3477_n2069, DP_OP_422J2_124_3477_n2068,
         DP_OP_422J2_124_3477_n2067, DP_OP_422J2_124_3477_n2066,
         DP_OP_422J2_124_3477_n2065, DP_OP_422J2_124_3477_n2064,
         DP_OP_422J2_124_3477_n2063, DP_OP_422J2_124_3477_n2062,
         DP_OP_422J2_124_3477_n2061, DP_OP_422J2_124_3477_n2060,
         DP_OP_422J2_124_3477_n2059, DP_OP_422J2_124_3477_n2058,
         DP_OP_422J2_124_3477_n2057, DP_OP_422J2_124_3477_n2056,
         DP_OP_422J2_124_3477_n2055, DP_OP_422J2_124_3477_n2054,
         DP_OP_422J2_124_3477_n2053, DP_OP_422J2_124_3477_n2052,
         DP_OP_422J2_124_3477_n2051, DP_OP_422J2_124_3477_n2050,
         DP_OP_422J2_124_3477_n2049, DP_OP_422J2_124_3477_n2048,
         DP_OP_422J2_124_3477_n2047, DP_OP_422J2_124_3477_n2045,
         DP_OP_422J2_124_3477_n2044, DP_OP_422J2_124_3477_n2040,
         DP_OP_422J2_124_3477_n2039, DP_OP_422J2_124_3477_n2038,
         DP_OP_422J2_124_3477_n2037, DP_OP_422J2_124_3477_n2036,
         DP_OP_422J2_124_3477_n2035, DP_OP_422J2_124_3477_n2034,
         DP_OP_422J2_124_3477_n2033, DP_OP_422J2_124_3477_n2032,
         DP_OP_422J2_124_3477_n2031, DP_OP_422J2_124_3477_n2030,
         DP_OP_422J2_124_3477_n2029, DP_OP_422J2_124_3477_n2028,
         DP_OP_422J2_124_3477_n2027, DP_OP_422J2_124_3477_n2026,
         DP_OP_422J2_124_3477_n2025, DP_OP_422J2_124_3477_n2024,
         DP_OP_422J2_124_3477_n2023, DP_OP_422J2_124_3477_n2022,
         DP_OP_422J2_124_3477_n2021, DP_OP_422J2_124_3477_n2020,
         DP_OP_422J2_124_3477_n2019, DP_OP_422J2_124_3477_n2018,
         DP_OP_422J2_124_3477_n2017, DP_OP_422J2_124_3477_n2016,
         DP_OP_422J2_124_3477_n2015, DP_OP_422J2_124_3477_n2014,
         DP_OP_422J2_124_3477_n2013, DP_OP_422J2_124_3477_n2012,
         DP_OP_422J2_124_3477_n2011, DP_OP_422J2_124_3477_n2010,
         DP_OP_422J2_124_3477_n2009, DP_OP_422J2_124_3477_n2008,
         DP_OP_422J2_124_3477_n2007, DP_OP_422J2_124_3477_n2006,
         DP_OP_422J2_124_3477_n2005, DP_OP_422J2_124_3477_n2004,
         DP_OP_422J2_124_3477_n2000, DP_OP_422J2_124_3477_n1995,
         DP_OP_422J2_124_3477_n1994, DP_OP_422J2_124_3477_n1993,
         DP_OP_422J2_124_3477_n1992, DP_OP_422J2_124_3477_n1991,
         DP_OP_422J2_124_3477_n1990, DP_OP_422J2_124_3477_n1989,
         DP_OP_422J2_124_3477_n1988, DP_OP_422J2_124_3477_n1987,
         DP_OP_422J2_124_3477_n1986, DP_OP_422J2_124_3477_n1985,
         DP_OP_422J2_124_3477_n1984, DP_OP_422J2_124_3477_n1983,
         DP_OP_422J2_124_3477_n1982, DP_OP_422J2_124_3477_n1981,
         DP_OP_422J2_124_3477_n1980, DP_OP_422J2_124_3477_n1979,
         DP_OP_422J2_124_3477_n1978, DP_OP_422J2_124_3477_n1977,
         DP_OP_422J2_124_3477_n1976, DP_OP_422J2_124_3477_n1975,
         DP_OP_422J2_124_3477_n1974, DP_OP_422J2_124_3477_n1973,
         DP_OP_422J2_124_3477_n1972, DP_OP_422J2_124_3477_n1971,
         DP_OP_422J2_124_3477_n1970, DP_OP_422J2_124_3477_n1969,
         DP_OP_422J2_124_3477_n1968, DP_OP_422J2_124_3477_n1967,
         DP_OP_422J2_124_3477_n1966, DP_OP_422J2_124_3477_n1965,
         DP_OP_422J2_124_3477_n1964, DP_OP_422J2_124_3477_n1963,
         DP_OP_422J2_124_3477_n1962, DP_OP_422J2_124_3477_n1961,
         DP_OP_422J2_124_3477_n1960, DP_OP_422J2_124_3477_n1958,
         DP_OP_422J2_124_3477_n1957, DP_OP_422J2_124_3477_n1951,
         DP_OP_422J2_124_3477_n1950, DP_OP_422J2_124_3477_n1949,
         DP_OP_422J2_124_3477_n1948, DP_OP_422J2_124_3477_n1947,
         DP_OP_422J2_124_3477_n1946, DP_OP_422J2_124_3477_n1945,
         DP_OP_422J2_124_3477_n1944, DP_OP_422J2_124_3477_n1943,
         DP_OP_422J2_124_3477_n1942, DP_OP_422J2_124_3477_n1941,
         DP_OP_422J2_124_3477_n1940, DP_OP_422J2_124_3477_n1939,
         DP_OP_422J2_124_3477_n1938, DP_OP_422J2_124_3477_n1937,
         DP_OP_422J2_124_3477_n1936, DP_OP_422J2_124_3477_n1935,
         DP_OP_422J2_124_3477_n1934, DP_OP_422J2_124_3477_n1933,
         DP_OP_422J2_124_3477_n1932, DP_OP_422J2_124_3477_n1931,
         DP_OP_422J2_124_3477_n1930, DP_OP_422J2_124_3477_n1929,
         DP_OP_422J2_124_3477_n1928, DP_OP_422J2_124_3477_n1927,
         DP_OP_422J2_124_3477_n1926, DP_OP_422J2_124_3477_n1925,
         DP_OP_422J2_124_3477_n1924, DP_OP_422J2_124_3477_n1923,
         DP_OP_422J2_124_3477_n1922, DP_OP_422J2_124_3477_n1921,
         DP_OP_422J2_124_3477_n1920, DP_OP_422J2_124_3477_n1886,
         DP_OP_422J2_124_3477_n1885, DP_OP_422J2_124_3477_n1884,
         DP_OP_422J2_124_3477_n1883, DP_OP_422J2_124_3477_n1882,
         DP_OP_422J2_124_3477_n1881, DP_OP_422J2_124_3477_n1880,
         DP_OP_422J2_124_3477_n1879, DP_OP_422J2_124_3477_n1878,
         DP_OP_422J2_124_3477_n1877, DP_OP_422J2_124_3477_n1876,
         DP_OP_422J2_124_3477_n1875, DP_OP_422J2_124_3477_n1874,
         DP_OP_422J2_124_3477_n1873, DP_OP_422J2_124_3477_n1871,
         DP_OP_422J2_124_3477_n1870, DP_OP_422J2_124_3477_n1869,
         DP_OP_422J2_124_3477_n1868, DP_OP_422J2_124_3477_n1867,
         DP_OP_422J2_124_3477_n1866, DP_OP_422J2_124_3477_n1865,
         DP_OP_422J2_124_3477_n1864, DP_OP_422J2_124_3477_n1863,
         DP_OP_422J2_124_3477_n1862, DP_OP_422J2_124_3477_n1861,
         DP_OP_422J2_124_3477_n1860, DP_OP_422J2_124_3477_n1859,
         DP_OP_422J2_124_3477_n1858, DP_OP_422J2_124_3477_n1857,
         DP_OP_422J2_124_3477_n1856, DP_OP_422J2_124_3477_n1855,
         DP_OP_422J2_124_3477_n1854, DP_OP_422J2_124_3477_n1853,
         DP_OP_422J2_124_3477_n1852, DP_OP_422J2_124_3477_n1851,
         DP_OP_422J2_124_3477_n1850, DP_OP_422J2_124_3477_n1849,
         DP_OP_422J2_124_3477_n1848, DP_OP_422J2_124_3477_n1847,
         DP_OP_422J2_124_3477_n1846, DP_OP_422J2_124_3477_n1845,
         DP_OP_422J2_124_3477_n1844, DP_OP_422J2_124_3477_n1843,
         DP_OP_422J2_124_3477_n1842, DP_OP_422J2_124_3477_n1841,
         DP_OP_422J2_124_3477_n1840, DP_OP_422J2_124_3477_n1839,
         DP_OP_422J2_124_3477_n1838, DP_OP_422J2_124_3477_n1837,
         DP_OP_422J2_124_3477_n1836, DP_OP_422J2_124_3477_n1835,
         DP_OP_422J2_124_3477_n1834, DP_OP_422J2_124_3477_n1833,
         DP_OP_422J2_124_3477_n1832, DP_OP_422J2_124_3477_n1831,
         DP_OP_422J2_124_3477_n1830, DP_OP_422J2_124_3477_n1829,
         DP_OP_422J2_124_3477_n1828, DP_OP_422J2_124_3477_n1827,
         DP_OP_422J2_124_3477_n1826, DP_OP_422J2_124_3477_n1825,
         DP_OP_422J2_124_3477_n1824, DP_OP_422J2_124_3477_n1823,
         DP_OP_422J2_124_3477_n1822, DP_OP_422J2_124_3477_n1821,
         DP_OP_422J2_124_3477_n1820, DP_OP_422J2_124_3477_n1819,
         DP_OP_422J2_124_3477_n1818, DP_OP_422J2_124_3477_n1817,
         DP_OP_422J2_124_3477_n1816, DP_OP_422J2_124_3477_n1815,
         DP_OP_422J2_124_3477_n1814, DP_OP_422J2_124_3477_n1813,
         DP_OP_422J2_124_3477_n1812, DP_OP_422J2_124_3477_n1811,
         DP_OP_422J2_124_3477_n1810, DP_OP_422J2_124_3477_n1809,
         DP_OP_422J2_124_3477_n1808, DP_OP_422J2_124_3477_n1807,
         DP_OP_422J2_124_3477_n1806, DP_OP_422J2_124_3477_n1805,
         DP_OP_422J2_124_3477_n1804, DP_OP_422J2_124_3477_n1803,
         DP_OP_422J2_124_3477_n1802, DP_OP_422J2_124_3477_n1801,
         DP_OP_422J2_124_3477_n1800, DP_OP_422J2_124_3477_n1799,
         DP_OP_422J2_124_3477_n1798, DP_OP_422J2_124_3477_n1797,
         DP_OP_422J2_124_3477_n1796, DP_OP_422J2_124_3477_n1795,
         DP_OP_422J2_124_3477_n1794, DP_OP_422J2_124_3477_n1793,
         DP_OP_422J2_124_3477_n1792, DP_OP_422J2_124_3477_n1791,
         DP_OP_422J2_124_3477_n1790, DP_OP_422J2_124_3477_n1789,
         DP_OP_422J2_124_3477_n1788, DP_OP_422J2_124_3477_n1787,
         DP_OP_422J2_124_3477_n1786, DP_OP_422J2_124_3477_n1785,
         DP_OP_422J2_124_3477_n1784, DP_OP_422J2_124_3477_n1783,
         DP_OP_422J2_124_3477_n1782, DP_OP_422J2_124_3477_n1781,
         DP_OP_422J2_124_3477_n1780, DP_OP_422J2_124_3477_n1779,
         DP_OP_422J2_124_3477_n1778, DP_OP_422J2_124_3477_n1777,
         DP_OP_422J2_124_3477_n1776, DP_OP_422J2_124_3477_n1775,
         DP_OP_422J2_124_3477_n1774, DP_OP_422J2_124_3477_n1773,
         DP_OP_422J2_124_3477_n1772, DP_OP_422J2_124_3477_n1771,
         DP_OP_422J2_124_3477_n1770, DP_OP_422J2_124_3477_n1769,
         DP_OP_422J2_124_3477_n1768, DP_OP_422J2_124_3477_n1767,
         DP_OP_422J2_124_3477_n1766, DP_OP_422J2_124_3477_n1765,
         DP_OP_422J2_124_3477_n1764, DP_OP_422J2_124_3477_n1763,
         DP_OP_422J2_124_3477_n1762, DP_OP_422J2_124_3477_n1761,
         DP_OP_422J2_124_3477_n1760, DP_OP_422J2_124_3477_n1759,
         DP_OP_422J2_124_3477_n1758, DP_OP_422J2_124_3477_n1757,
         DP_OP_422J2_124_3477_n1756, DP_OP_422J2_124_3477_n1755,
         DP_OP_422J2_124_3477_n1754, DP_OP_422J2_124_3477_n1753,
         DP_OP_422J2_124_3477_n1752, DP_OP_422J2_124_3477_n1751,
         DP_OP_422J2_124_3477_n1750, DP_OP_422J2_124_3477_n1749,
         DP_OP_422J2_124_3477_n1748, DP_OP_422J2_124_3477_n1747,
         DP_OP_422J2_124_3477_n1746, DP_OP_422J2_124_3477_n1745,
         DP_OP_422J2_124_3477_n1744, DP_OP_422J2_124_3477_n1743,
         DP_OP_422J2_124_3477_n1742, DP_OP_422J2_124_3477_n1741,
         DP_OP_422J2_124_3477_n1740, DP_OP_422J2_124_3477_n1739,
         DP_OP_422J2_124_3477_n1738, DP_OP_422J2_124_3477_n1737,
         DP_OP_422J2_124_3477_n1736, DP_OP_422J2_124_3477_n1735,
         DP_OP_422J2_124_3477_n1734, DP_OP_422J2_124_3477_n1733,
         DP_OP_422J2_124_3477_n1732, DP_OP_422J2_124_3477_n1731,
         DP_OP_422J2_124_3477_n1730, DP_OP_422J2_124_3477_n1729,
         DP_OP_422J2_124_3477_n1728, DP_OP_422J2_124_3477_n1727,
         DP_OP_422J2_124_3477_n1726, DP_OP_422J2_124_3477_n1725,
         DP_OP_422J2_124_3477_n1724, DP_OP_422J2_124_3477_n1723,
         DP_OP_422J2_124_3477_n1722, DP_OP_422J2_124_3477_n1721,
         DP_OP_422J2_124_3477_n1720, DP_OP_422J2_124_3477_n1719,
         DP_OP_422J2_124_3477_n1718, DP_OP_422J2_124_3477_n1717,
         DP_OP_422J2_124_3477_n1716, DP_OP_422J2_124_3477_n1715,
         DP_OP_422J2_124_3477_n1714, DP_OP_422J2_124_3477_n1713,
         DP_OP_422J2_124_3477_n1712, DP_OP_422J2_124_3477_n1711,
         DP_OP_422J2_124_3477_n1710, DP_OP_422J2_124_3477_n1709,
         DP_OP_422J2_124_3477_n1708, DP_OP_422J2_124_3477_n1707,
         DP_OP_422J2_124_3477_n1706, DP_OP_422J2_124_3477_n1705,
         DP_OP_422J2_124_3477_n1704, DP_OP_422J2_124_3477_n1703,
         DP_OP_422J2_124_3477_n1702, DP_OP_422J2_124_3477_n1701,
         DP_OP_422J2_124_3477_n1700, DP_OP_422J2_124_3477_n1699,
         DP_OP_422J2_124_3477_n1698, DP_OP_422J2_124_3477_n1697,
         DP_OP_422J2_124_3477_n1696, DP_OP_422J2_124_3477_n1695,
         DP_OP_422J2_124_3477_n1694, DP_OP_422J2_124_3477_n1693,
         DP_OP_422J2_124_3477_n1692, DP_OP_422J2_124_3477_n1691,
         DP_OP_422J2_124_3477_n1690, DP_OP_422J2_124_3477_n1689,
         DP_OP_422J2_124_3477_n1688, DP_OP_422J2_124_3477_n1687,
         DP_OP_422J2_124_3477_n1686, DP_OP_422J2_124_3477_n1685,
         DP_OP_422J2_124_3477_n1684, DP_OP_422J2_124_3477_n1683,
         DP_OP_422J2_124_3477_n1682, DP_OP_422J2_124_3477_n1681,
         DP_OP_422J2_124_3477_n1680, DP_OP_422J2_124_3477_n1679,
         DP_OP_422J2_124_3477_n1678, DP_OP_422J2_124_3477_n1677,
         DP_OP_422J2_124_3477_n1676, DP_OP_422J2_124_3477_n1675,
         DP_OP_422J2_124_3477_n1674, DP_OP_422J2_124_3477_n1673,
         DP_OP_422J2_124_3477_n1672, DP_OP_422J2_124_3477_n1671,
         DP_OP_422J2_124_3477_n1670, DP_OP_422J2_124_3477_n1669,
         DP_OP_422J2_124_3477_n1668, DP_OP_422J2_124_3477_n1667,
         DP_OP_422J2_124_3477_n1666, DP_OP_422J2_124_3477_n1665,
         DP_OP_422J2_124_3477_n1664, DP_OP_422J2_124_3477_n1663,
         DP_OP_422J2_124_3477_n1662, DP_OP_422J2_124_3477_n1661,
         DP_OP_422J2_124_3477_n1660, DP_OP_422J2_124_3477_n1659,
         DP_OP_422J2_124_3477_n1658, DP_OP_422J2_124_3477_n1657,
         DP_OP_422J2_124_3477_n1656, DP_OP_422J2_124_3477_n1655,
         DP_OP_422J2_124_3477_n1654, DP_OP_422J2_124_3477_n1653,
         DP_OP_422J2_124_3477_n1652, DP_OP_422J2_124_3477_n1651,
         DP_OP_422J2_124_3477_n1650, DP_OP_422J2_124_3477_n1649,
         DP_OP_422J2_124_3477_n1648, DP_OP_422J2_124_3477_n1647,
         DP_OP_422J2_124_3477_n1646, DP_OP_422J2_124_3477_n1645,
         DP_OP_422J2_124_3477_n1644, DP_OP_422J2_124_3477_n1643,
         DP_OP_422J2_124_3477_n1642, DP_OP_422J2_124_3477_n1641,
         DP_OP_422J2_124_3477_n1640, DP_OP_422J2_124_3477_n1639,
         DP_OP_422J2_124_3477_n1638, DP_OP_422J2_124_3477_n1637,
         DP_OP_422J2_124_3477_n1636, DP_OP_422J2_124_3477_n1635,
         DP_OP_422J2_124_3477_n1634, DP_OP_422J2_124_3477_n1633,
         DP_OP_422J2_124_3477_n1632, DP_OP_422J2_124_3477_n1631,
         DP_OP_422J2_124_3477_n1630, DP_OP_422J2_124_3477_n1629,
         DP_OP_422J2_124_3477_n1628, DP_OP_422J2_124_3477_n1627,
         DP_OP_422J2_124_3477_n1626, DP_OP_422J2_124_3477_n1625,
         DP_OP_422J2_124_3477_n1624, DP_OP_422J2_124_3477_n1623,
         DP_OP_422J2_124_3477_n1622, DP_OP_422J2_124_3477_n1621,
         DP_OP_422J2_124_3477_n1620, DP_OP_422J2_124_3477_n1619,
         DP_OP_422J2_124_3477_n1618, DP_OP_422J2_124_3477_n1617,
         DP_OP_422J2_124_3477_n1616, DP_OP_422J2_124_3477_n1615,
         DP_OP_422J2_124_3477_n1614, DP_OP_422J2_124_3477_n1613,
         DP_OP_422J2_124_3477_n1612, DP_OP_422J2_124_3477_n1611,
         DP_OP_422J2_124_3477_n1610, DP_OP_422J2_124_3477_n1609,
         DP_OP_422J2_124_3477_n1608, DP_OP_422J2_124_3477_n1607,
         DP_OP_422J2_124_3477_n1606, DP_OP_422J2_124_3477_n1605,
         DP_OP_422J2_124_3477_n1604, DP_OP_422J2_124_3477_n1603,
         DP_OP_422J2_124_3477_n1602, DP_OP_422J2_124_3477_n1601,
         DP_OP_422J2_124_3477_n1600, DP_OP_422J2_124_3477_n1599,
         DP_OP_422J2_124_3477_n1598, DP_OP_422J2_124_3477_n1597,
         DP_OP_422J2_124_3477_n1596, DP_OP_422J2_124_3477_n1595,
         DP_OP_422J2_124_3477_n1594, DP_OP_422J2_124_3477_n1593,
         DP_OP_422J2_124_3477_n1592, DP_OP_422J2_124_3477_n1591,
         DP_OP_422J2_124_3477_n1590, DP_OP_422J2_124_3477_n1589,
         DP_OP_422J2_124_3477_n1588, DP_OP_422J2_124_3477_n1587,
         DP_OP_422J2_124_3477_n1586, DP_OP_422J2_124_3477_n1585,
         DP_OP_422J2_124_3477_n1584, DP_OP_422J2_124_3477_n1583,
         DP_OP_422J2_124_3477_n1582, DP_OP_422J2_124_3477_n1581,
         DP_OP_422J2_124_3477_n1580, DP_OP_422J2_124_3477_n1579,
         DP_OP_422J2_124_3477_n1578, DP_OP_422J2_124_3477_n1577,
         DP_OP_422J2_124_3477_n1576, DP_OP_422J2_124_3477_n1575,
         DP_OP_422J2_124_3477_n1574, DP_OP_422J2_124_3477_n1573,
         DP_OP_422J2_124_3477_n1572, DP_OP_422J2_124_3477_n1571,
         DP_OP_422J2_124_3477_n1570, DP_OP_422J2_124_3477_n1569,
         DP_OP_422J2_124_3477_n1568, DP_OP_422J2_124_3477_n1567,
         DP_OP_422J2_124_3477_n1566, DP_OP_422J2_124_3477_n1565,
         DP_OP_422J2_124_3477_n1564, DP_OP_422J2_124_3477_n1563,
         DP_OP_422J2_124_3477_n1562, DP_OP_422J2_124_3477_n1561,
         DP_OP_422J2_124_3477_n1560, DP_OP_422J2_124_3477_n1559,
         DP_OP_422J2_124_3477_n1558, DP_OP_422J2_124_3477_n1557,
         DP_OP_422J2_124_3477_n1556, DP_OP_422J2_124_3477_n1555,
         DP_OP_422J2_124_3477_n1554, DP_OP_422J2_124_3477_n1553,
         DP_OP_422J2_124_3477_n1552, DP_OP_422J2_124_3477_n1551,
         DP_OP_422J2_124_3477_n1550, DP_OP_422J2_124_3477_n1549,
         DP_OP_422J2_124_3477_n1548, DP_OP_422J2_124_3477_n1547,
         DP_OP_422J2_124_3477_n1546, DP_OP_422J2_124_3477_n1545,
         DP_OP_422J2_124_3477_n1544, DP_OP_422J2_124_3477_n1543,
         DP_OP_422J2_124_3477_n1542, DP_OP_422J2_124_3477_n1541,
         DP_OP_422J2_124_3477_n1540, DP_OP_422J2_124_3477_n1539,
         DP_OP_422J2_124_3477_n1538, DP_OP_422J2_124_3477_n1537,
         DP_OP_422J2_124_3477_n1536, DP_OP_422J2_124_3477_n1535,
         DP_OP_422J2_124_3477_n1534, DP_OP_422J2_124_3477_n1533,
         DP_OP_422J2_124_3477_n1532, DP_OP_422J2_124_3477_n1531,
         DP_OP_422J2_124_3477_n1530, DP_OP_422J2_124_3477_n1529,
         DP_OP_422J2_124_3477_n1528, DP_OP_422J2_124_3477_n1527,
         DP_OP_422J2_124_3477_n1526, DP_OP_422J2_124_3477_n1525,
         DP_OP_422J2_124_3477_n1524, DP_OP_422J2_124_3477_n1523,
         DP_OP_422J2_124_3477_n1522, DP_OP_422J2_124_3477_n1521,
         DP_OP_422J2_124_3477_n1520, DP_OP_422J2_124_3477_n1519,
         DP_OP_422J2_124_3477_n1518, DP_OP_422J2_124_3477_n1517,
         DP_OP_422J2_124_3477_n1516, DP_OP_422J2_124_3477_n1515,
         DP_OP_422J2_124_3477_n1514, DP_OP_422J2_124_3477_n1513,
         DP_OP_422J2_124_3477_n1512, DP_OP_422J2_124_3477_n1511,
         DP_OP_422J2_124_3477_n1510, DP_OP_422J2_124_3477_n1509,
         DP_OP_422J2_124_3477_n1508, DP_OP_422J2_124_3477_n1507,
         DP_OP_422J2_124_3477_n1506, DP_OP_422J2_124_3477_n1505,
         DP_OP_422J2_124_3477_n1504, DP_OP_422J2_124_3477_n1503,
         DP_OP_422J2_124_3477_n1502, DP_OP_422J2_124_3477_n1501,
         DP_OP_422J2_124_3477_n1500, DP_OP_422J2_124_3477_n1499,
         DP_OP_422J2_124_3477_n1498, DP_OP_422J2_124_3477_n1497,
         DP_OP_422J2_124_3477_n1496, DP_OP_422J2_124_3477_n1495,
         DP_OP_422J2_124_3477_n1494, DP_OP_422J2_124_3477_n1493,
         DP_OP_422J2_124_3477_n1492, DP_OP_422J2_124_3477_n1491,
         DP_OP_422J2_124_3477_n1490, DP_OP_422J2_124_3477_n1489,
         DP_OP_422J2_124_3477_n1488, DP_OP_422J2_124_3477_n1487,
         DP_OP_422J2_124_3477_n1486, DP_OP_422J2_124_3477_n1485,
         DP_OP_422J2_124_3477_n1484, DP_OP_422J2_124_3477_n1483,
         DP_OP_422J2_124_3477_n1482, DP_OP_422J2_124_3477_n1481,
         DP_OP_422J2_124_3477_n1480, DP_OP_422J2_124_3477_n1479,
         DP_OP_422J2_124_3477_n1478, DP_OP_422J2_124_3477_n1477,
         DP_OP_422J2_124_3477_n1476, DP_OP_422J2_124_3477_n1475,
         DP_OP_422J2_124_3477_n1474, DP_OP_422J2_124_3477_n1473,
         DP_OP_422J2_124_3477_n1472, DP_OP_422J2_124_3477_n1471,
         DP_OP_422J2_124_3477_n1470, DP_OP_422J2_124_3477_n1469,
         DP_OP_422J2_124_3477_n1468, DP_OP_422J2_124_3477_n1467,
         DP_OP_422J2_124_3477_n1466, DP_OP_422J2_124_3477_n1465,
         DP_OP_422J2_124_3477_n1464, DP_OP_422J2_124_3477_n1463,
         DP_OP_422J2_124_3477_n1462, DP_OP_422J2_124_3477_n1461,
         DP_OP_422J2_124_3477_n1460, DP_OP_422J2_124_3477_n1459,
         DP_OP_422J2_124_3477_n1458, DP_OP_422J2_124_3477_n1457,
         DP_OP_422J2_124_3477_n1456, DP_OP_422J2_124_3477_n1455,
         DP_OP_422J2_124_3477_n1454, DP_OP_422J2_124_3477_n1453,
         DP_OP_422J2_124_3477_n1452, DP_OP_422J2_124_3477_n1451,
         DP_OP_422J2_124_3477_n1450, DP_OP_422J2_124_3477_n1449,
         DP_OP_422J2_124_3477_n1448, DP_OP_422J2_124_3477_n1447,
         DP_OP_422J2_124_3477_n1446, DP_OP_422J2_124_3477_n1445,
         DP_OP_422J2_124_3477_n1444, DP_OP_422J2_124_3477_n1443,
         DP_OP_422J2_124_3477_n1442, DP_OP_422J2_124_3477_n1441,
         DP_OP_422J2_124_3477_n1440, DP_OP_422J2_124_3477_n1439,
         DP_OP_422J2_124_3477_n1438, DP_OP_422J2_124_3477_n1437,
         DP_OP_422J2_124_3477_n1436, DP_OP_422J2_124_3477_n1435,
         DP_OP_422J2_124_3477_n1434, DP_OP_422J2_124_3477_n1433,
         DP_OP_422J2_124_3477_n1432, DP_OP_422J2_124_3477_n1431,
         DP_OP_422J2_124_3477_n1430, DP_OP_422J2_124_3477_n1429,
         DP_OP_422J2_124_3477_n1428, DP_OP_422J2_124_3477_n1427,
         DP_OP_422J2_124_3477_n1426, DP_OP_422J2_124_3477_n1425,
         DP_OP_422J2_124_3477_n1424, DP_OP_422J2_124_3477_n1423,
         DP_OP_422J2_124_3477_n1422, DP_OP_422J2_124_3477_n1421,
         DP_OP_422J2_124_3477_n1420, DP_OP_422J2_124_3477_n1419,
         DP_OP_422J2_124_3477_n1418, DP_OP_422J2_124_3477_n1417,
         DP_OP_422J2_124_3477_n1416, DP_OP_422J2_124_3477_n1415,
         DP_OP_422J2_124_3477_n1414, DP_OP_422J2_124_3477_n1413,
         DP_OP_422J2_124_3477_n1412, DP_OP_422J2_124_3477_n1411,
         DP_OP_422J2_124_3477_n1410, DP_OP_422J2_124_3477_n1409,
         DP_OP_422J2_124_3477_n1408, DP_OP_422J2_124_3477_n1407,
         DP_OP_422J2_124_3477_n1406, DP_OP_422J2_124_3477_n1405,
         DP_OP_422J2_124_3477_n1404, DP_OP_422J2_124_3477_n1403,
         DP_OP_422J2_124_3477_n1402, DP_OP_422J2_124_3477_n1401,
         DP_OP_422J2_124_3477_n1400, DP_OP_422J2_124_3477_n1399,
         DP_OP_422J2_124_3477_n1398, DP_OP_422J2_124_3477_n1397,
         DP_OP_422J2_124_3477_n1396, DP_OP_422J2_124_3477_n1395,
         DP_OP_422J2_124_3477_n1394, DP_OP_422J2_124_3477_n1393,
         DP_OP_422J2_124_3477_n1392, DP_OP_422J2_124_3477_n1391,
         DP_OP_422J2_124_3477_n1390, DP_OP_422J2_124_3477_n1389,
         DP_OP_422J2_124_3477_n1388, DP_OP_422J2_124_3477_n1387,
         DP_OP_422J2_124_3477_n1386, DP_OP_422J2_124_3477_n1385,
         DP_OP_422J2_124_3477_n1384, DP_OP_422J2_124_3477_n1383,
         DP_OP_422J2_124_3477_n1382, DP_OP_422J2_124_3477_n1381,
         DP_OP_422J2_124_3477_n1380, DP_OP_422J2_124_3477_n1379,
         DP_OP_422J2_124_3477_n1378, DP_OP_422J2_124_3477_n1377,
         DP_OP_422J2_124_3477_n1376, DP_OP_422J2_124_3477_n1375,
         DP_OP_422J2_124_3477_n1374, DP_OP_422J2_124_3477_n1373,
         DP_OP_422J2_124_3477_n1372, DP_OP_422J2_124_3477_n1371,
         DP_OP_422J2_124_3477_n1370, DP_OP_422J2_124_3477_n1369,
         DP_OP_422J2_124_3477_n1368, DP_OP_422J2_124_3477_n1367,
         DP_OP_422J2_124_3477_n1366, DP_OP_422J2_124_3477_n1365,
         DP_OP_422J2_124_3477_n1364, DP_OP_422J2_124_3477_n1363,
         DP_OP_422J2_124_3477_n1362, DP_OP_422J2_124_3477_n1361,
         DP_OP_422J2_124_3477_n1360, DP_OP_422J2_124_3477_n1359,
         DP_OP_422J2_124_3477_n1358, DP_OP_422J2_124_3477_n1357,
         DP_OP_422J2_124_3477_n1356, DP_OP_422J2_124_3477_n1355,
         DP_OP_422J2_124_3477_n1354, DP_OP_422J2_124_3477_n1353,
         DP_OP_422J2_124_3477_n1352, DP_OP_422J2_124_3477_n1351,
         DP_OP_422J2_124_3477_n1350, DP_OP_422J2_124_3477_n1349,
         DP_OP_422J2_124_3477_n1348, DP_OP_422J2_124_3477_n1347,
         DP_OP_422J2_124_3477_n1346, DP_OP_422J2_124_3477_n1345,
         DP_OP_422J2_124_3477_n1344, DP_OP_422J2_124_3477_n1343,
         DP_OP_422J2_124_3477_n1342, DP_OP_422J2_124_3477_n1341,
         DP_OP_422J2_124_3477_n1340, DP_OP_422J2_124_3477_n1339,
         DP_OP_422J2_124_3477_n1338, DP_OP_422J2_124_3477_n1337,
         DP_OP_422J2_124_3477_n1336, DP_OP_422J2_124_3477_n1335,
         DP_OP_422J2_124_3477_n1334, DP_OP_422J2_124_3477_n1333,
         DP_OP_422J2_124_3477_n1332, DP_OP_422J2_124_3477_n1331,
         DP_OP_422J2_124_3477_n1330, DP_OP_422J2_124_3477_n1329,
         DP_OP_422J2_124_3477_n1328, DP_OP_422J2_124_3477_n1327,
         DP_OP_422J2_124_3477_n1326, DP_OP_422J2_124_3477_n1325,
         DP_OP_422J2_124_3477_n1324, DP_OP_422J2_124_3477_n1323,
         DP_OP_422J2_124_3477_n1322, DP_OP_422J2_124_3477_n1321,
         DP_OP_422J2_124_3477_n1320, DP_OP_422J2_124_3477_n1319,
         DP_OP_422J2_124_3477_n1318, DP_OP_422J2_124_3477_n1317,
         DP_OP_422J2_124_3477_n1316, DP_OP_422J2_124_3477_n1315,
         DP_OP_422J2_124_3477_n1314, DP_OP_422J2_124_3477_n1313,
         DP_OP_422J2_124_3477_n1312, DP_OP_422J2_124_3477_n1311,
         DP_OP_422J2_124_3477_n1310, DP_OP_422J2_124_3477_n1309,
         DP_OP_422J2_124_3477_n1308, DP_OP_422J2_124_3477_n1307,
         DP_OP_422J2_124_3477_n1306, DP_OP_422J2_124_3477_n1305,
         DP_OP_422J2_124_3477_n1304, DP_OP_422J2_124_3477_n1303,
         DP_OP_422J2_124_3477_n1302, DP_OP_422J2_124_3477_n1301,
         DP_OP_422J2_124_3477_n1300, DP_OP_422J2_124_3477_n1299,
         DP_OP_422J2_124_3477_n1298, DP_OP_422J2_124_3477_n1297,
         DP_OP_422J2_124_3477_n1296, DP_OP_422J2_124_3477_n1295,
         DP_OP_422J2_124_3477_n1294, DP_OP_422J2_124_3477_n1293,
         DP_OP_422J2_124_3477_n1292, DP_OP_422J2_124_3477_n1291,
         DP_OP_422J2_124_3477_n1290, DP_OP_422J2_124_3477_n1289,
         DP_OP_422J2_124_3477_n1288, DP_OP_422J2_124_3477_n1287,
         DP_OP_422J2_124_3477_n1286, DP_OP_422J2_124_3477_n1285,
         DP_OP_422J2_124_3477_n1284, DP_OP_422J2_124_3477_n1283,
         DP_OP_422J2_124_3477_n1282, DP_OP_422J2_124_3477_n1281,
         DP_OP_422J2_124_3477_n1280, DP_OP_422J2_124_3477_n1279,
         DP_OP_422J2_124_3477_n1278, DP_OP_422J2_124_3477_n1277,
         DP_OP_422J2_124_3477_n1276, DP_OP_422J2_124_3477_n1275,
         DP_OP_422J2_124_3477_n1274, DP_OP_422J2_124_3477_n1273,
         DP_OP_422J2_124_3477_n1272, DP_OP_422J2_124_3477_n1271,
         DP_OP_422J2_124_3477_n1270, DP_OP_422J2_124_3477_n1269,
         DP_OP_422J2_124_3477_n1268, DP_OP_422J2_124_3477_n1267,
         DP_OP_422J2_124_3477_n1266, DP_OP_422J2_124_3477_n1265,
         DP_OP_422J2_124_3477_n1264, DP_OP_422J2_124_3477_n1263,
         DP_OP_422J2_124_3477_n1262, DP_OP_422J2_124_3477_n1261,
         DP_OP_422J2_124_3477_n1260, DP_OP_422J2_124_3477_n1259,
         DP_OP_422J2_124_3477_n1258, DP_OP_422J2_124_3477_n1257,
         DP_OP_422J2_124_3477_n1256, DP_OP_422J2_124_3477_n1255,
         DP_OP_422J2_124_3477_n1254, DP_OP_422J2_124_3477_n1253,
         DP_OP_422J2_124_3477_n1252, DP_OP_422J2_124_3477_n1251,
         DP_OP_422J2_124_3477_n1250, DP_OP_422J2_124_3477_n1249,
         DP_OP_422J2_124_3477_n1248, DP_OP_422J2_124_3477_n1247,
         DP_OP_422J2_124_3477_n1246, DP_OP_422J2_124_3477_n1245,
         DP_OP_422J2_124_3477_n1244, DP_OP_422J2_124_3477_n1243,
         DP_OP_422J2_124_3477_n1242, DP_OP_422J2_124_3477_n1241,
         DP_OP_422J2_124_3477_n1240, DP_OP_422J2_124_3477_n1239,
         DP_OP_422J2_124_3477_n1238, DP_OP_422J2_124_3477_n1237,
         DP_OP_422J2_124_3477_n1236, DP_OP_422J2_124_3477_n1235,
         DP_OP_422J2_124_3477_n1234, DP_OP_422J2_124_3477_n1233,
         DP_OP_422J2_124_3477_n1232, DP_OP_422J2_124_3477_n1231,
         DP_OP_422J2_124_3477_n1230, DP_OP_422J2_124_3477_n1229,
         DP_OP_422J2_124_3477_n1228, DP_OP_422J2_124_3477_n1227,
         DP_OP_422J2_124_3477_n1226, DP_OP_422J2_124_3477_n1225,
         DP_OP_422J2_124_3477_n1224, DP_OP_422J2_124_3477_n1223,
         DP_OP_422J2_124_3477_n1222, DP_OP_422J2_124_3477_n1221,
         DP_OP_422J2_124_3477_n1220, DP_OP_422J2_124_3477_n1219,
         DP_OP_422J2_124_3477_n1218, DP_OP_422J2_124_3477_n1217,
         DP_OP_422J2_124_3477_n1216, DP_OP_422J2_124_3477_n1215,
         DP_OP_422J2_124_3477_n1214, DP_OP_422J2_124_3477_n1213,
         DP_OP_422J2_124_3477_n1212, DP_OP_422J2_124_3477_n1211,
         DP_OP_422J2_124_3477_n1210, DP_OP_422J2_124_3477_n1209,
         DP_OP_422J2_124_3477_n1208, DP_OP_422J2_124_3477_n1207,
         DP_OP_422J2_124_3477_n1206, DP_OP_422J2_124_3477_n1205,
         DP_OP_422J2_124_3477_n1204, DP_OP_422J2_124_3477_n1203,
         DP_OP_422J2_124_3477_n1202, DP_OP_422J2_124_3477_n1201,
         DP_OP_422J2_124_3477_n1200, DP_OP_422J2_124_3477_n1199,
         DP_OP_422J2_124_3477_n1198, DP_OP_422J2_124_3477_n1197,
         DP_OP_422J2_124_3477_n1196, DP_OP_422J2_124_3477_n1195,
         DP_OP_422J2_124_3477_n1194, DP_OP_422J2_124_3477_n1193,
         DP_OP_422J2_124_3477_n1192, DP_OP_422J2_124_3477_n1191,
         DP_OP_422J2_124_3477_n1190, DP_OP_422J2_124_3477_n1189,
         DP_OP_422J2_124_3477_n1188, DP_OP_422J2_124_3477_n1187,
         DP_OP_422J2_124_3477_n1186, DP_OP_422J2_124_3477_n1185,
         DP_OP_422J2_124_3477_n1184, DP_OP_422J2_124_3477_n1183,
         DP_OP_422J2_124_3477_n1182, DP_OP_422J2_124_3477_n1181,
         DP_OP_422J2_124_3477_n1180, DP_OP_422J2_124_3477_n1179,
         DP_OP_422J2_124_3477_n1178, DP_OP_422J2_124_3477_n1177,
         DP_OP_422J2_124_3477_n1176, DP_OP_422J2_124_3477_n1175,
         DP_OP_422J2_124_3477_n1174, DP_OP_422J2_124_3477_n1173,
         DP_OP_422J2_124_3477_n1172, DP_OP_422J2_124_3477_n1171,
         DP_OP_422J2_124_3477_n1170, DP_OP_422J2_124_3477_n1169,
         DP_OP_422J2_124_3477_n1168, DP_OP_422J2_124_3477_n1167,
         DP_OP_422J2_124_3477_n1166, DP_OP_422J2_124_3477_n1165,
         DP_OP_422J2_124_3477_n1164, DP_OP_422J2_124_3477_n1163,
         DP_OP_422J2_124_3477_n1162, DP_OP_422J2_124_3477_n1161,
         DP_OP_422J2_124_3477_n1160, DP_OP_422J2_124_3477_n1159,
         DP_OP_422J2_124_3477_n1158, DP_OP_422J2_124_3477_n1157,
         DP_OP_422J2_124_3477_n1156, DP_OP_422J2_124_3477_n1155,
         DP_OP_422J2_124_3477_n1154, DP_OP_422J2_124_3477_n1153,
         DP_OP_422J2_124_3477_n1152, DP_OP_422J2_124_3477_n1151,
         DP_OP_422J2_124_3477_n1150, DP_OP_422J2_124_3477_n1149,
         DP_OP_422J2_124_3477_n1148, DP_OP_422J2_124_3477_n1147,
         DP_OP_422J2_124_3477_n1146, DP_OP_422J2_124_3477_n1145,
         DP_OP_422J2_124_3477_n1144, DP_OP_422J2_124_3477_n1143,
         DP_OP_422J2_124_3477_n1142, DP_OP_422J2_124_3477_n1141,
         DP_OP_422J2_124_3477_n1140, DP_OP_422J2_124_3477_n1139,
         DP_OP_422J2_124_3477_n1138, DP_OP_422J2_124_3477_n1137,
         DP_OP_422J2_124_3477_n1136, DP_OP_422J2_124_3477_n1135,
         DP_OP_422J2_124_3477_n1134, DP_OP_422J2_124_3477_n1133,
         DP_OP_422J2_124_3477_n1132, DP_OP_422J2_124_3477_n1131,
         DP_OP_422J2_124_3477_n1130, DP_OP_422J2_124_3477_n1129,
         DP_OP_422J2_124_3477_n1128, DP_OP_422J2_124_3477_n1127,
         DP_OP_422J2_124_3477_n1126, DP_OP_422J2_124_3477_n1125,
         DP_OP_422J2_124_3477_n1124, DP_OP_422J2_124_3477_n1123,
         DP_OP_422J2_124_3477_n1122, DP_OP_422J2_124_3477_n1121,
         DP_OP_422J2_124_3477_n1120, DP_OP_422J2_124_3477_n1119,
         DP_OP_422J2_124_3477_n1118, DP_OP_422J2_124_3477_n1117,
         DP_OP_422J2_124_3477_n1116, DP_OP_422J2_124_3477_n1115,
         DP_OP_422J2_124_3477_n1114, DP_OP_422J2_124_3477_n1113,
         DP_OP_422J2_124_3477_n1112, DP_OP_422J2_124_3477_n1111,
         DP_OP_422J2_124_3477_n1110, DP_OP_422J2_124_3477_n1109,
         DP_OP_422J2_124_3477_n1108, DP_OP_422J2_124_3477_n1107,
         DP_OP_422J2_124_3477_n1106, DP_OP_422J2_124_3477_n1105,
         DP_OP_422J2_124_3477_n1104, DP_OP_422J2_124_3477_n1103,
         DP_OP_422J2_124_3477_n1102, DP_OP_422J2_124_3477_n1101,
         DP_OP_422J2_124_3477_n1100, DP_OP_422J2_124_3477_n1099,
         DP_OP_422J2_124_3477_n1098, DP_OP_422J2_124_3477_n1097,
         DP_OP_422J2_124_3477_n1096, DP_OP_422J2_124_3477_n1095,
         DP_OP_422J2_124_3477_n1094, DP_OP_422J2_124_3477_n1093,
         DP_OP_422J2_124_3477_n1092, DP_OP_422J2_124_3477_n1091,
         DP_OP_422J2_124_3477_n1090, DP_OP_422J2_124_3477_n1089,
         DP_OP_422J2_124_3477_n1088, DP_OP_422J2_124_3477_n1087,
         DP_OP_422J2_124_3477_n1086, DP_OP_422J2_124_3477_n1085,
         DP_OP_422J2_124_3477_n1084, DP_OP_422J2_124_3477_n1083,
         DP_OP_422J2_124_3477_n1082, DP_OP_422J2_124_3477_n1081,
         DP_OP_422J2_124_3477_n1080, DP_OP_422J2_124_3477_n1079,
         DP_OP_422J2_124_3477_n1078, DP_OP_422J2_124_3477_n1077,
         DP_OP_422J2_124_3477_n1076, DP_OP_422J2_124_3477_n1075,
         DP_OP_422J2_124_3477_n1074, DP_OP_422J2_124_3477_n1073,
         DP_OP_422J2_124_3477_n1072, DP_OP_422J2_124_3477_n1071,
         DP_OP_422J2_124_3477_n1070, DP_OP_422J2_124_3477_n1069,
         DP_OP_422J2_124_3477_n1068, DP_OP_422J2_124_3477_n1067,
         DP_OP_422J2_124_3477_n1066, DP_OP_422J2_124_3477_n1065,
         DP_OP_422J2_124_3477_n1064, DP_OP_422J2_124_3477_n1063,
         DP_OP_422J2_124_3477_n1062, DP_OP_422J2_124_3477_n1061,
         DP_OP_422J2_124_3477_n1060, DP_OP_422J2_124_3477_n1059,
         DP_OP_422J2_124_3477_n1058, DP_OP_422J2_124_3477_n1057,
         DP_OP_422J2_124_3477_n1056, DP_OP_422J2_124_3477_n1055,
         DP_OP_422J2_124_3477_n1054, DP_OP_422J2_124_3477_n1053,
         DP_OP_422J2_124_3477_n1052, DP_OP_422J2_124_3477_n1051,
         DP_OP_422J2_124_3477_n1050, DP_OP_422J2_124_3477_n1049,
         DP_OP_422J2_124_3477_n1048, DP_OP_422J2_124_3477_n1047,
         DP_OP_422J2_124_3477_n1046, DP_OP_422J2_124_3477_n1045,
         DP_OP_422J2_124_3477_n1044, DP_OP_422J2_124_3477_n1043,
         DP_OP_422J2_124_3477_n1042, DP_OP_422J2_124_3477_n1041,
         DP_OP_422J2_124_3477_n1040, DP_OP_422J2_124_3477_n1039,
         DP_OP_422J2_124_3477_n1038, DP_OP_422J2_124_3477_n1037,
         DP_OP_422J2_124_3477_n1036, DP_OP_422J2_124_3477_n1035,
         DP_OP_422J2_124_3477_n1034, DP_OP_422J2_124_3477_n1033,
         DP_OP_422J2_124_3477_n1032, DP_OP_422J2_124_3477_n1031,
         DP_OP_422J2_124_3477_n1030, DP_OP_422J2_124_3477_n1029,
         DP_OP_422J2_124_3477_n1028, DP_OP_422J2_124_3477_n1027,
         DP_OP_422J2_124_3477_n1026, DP_OP_422J2_124_3477_n1025,
         DP_OP_422J2_124_3477_n1024, DP_OP_422J2_124_3477_n1023,
         DP_OP_422J2_124_3477_n1022, DP_OP_422J2_124_3477_n1021,
         DP_OP_422J2_124_3477_n1020, DP_OP_422J2_124_3477_n1019,
         DP_OP_422J2_124_3477_n1018, DP_OP_422J2_124_3477_n1017,
         DP_OP_422J2_124_3477_n1016, DP_OP_422J2_124_3477_n1015,
         DP_OP_422J2_124_3477_n1014, DP_OP_422J2_124_3477_n1013,
         DP_OP_422J2_124_3477_n1012, DP_OP_422J2_124_3477_n1011,
         DP_OP_422J2_124_3477_n1010, DP_OP_422J2_124_3477_n1009,
         DP_OP_422J2_124_3477_n1008, DP_OP_422J2_124_3477_n1007,
         DP_OP_422J2_124_3477_n1006, DP_OP_422J2_124_3477_n1005,
         DP_OP_422J2_124_3477_n1004, DP_OP_422J2_124_3477_n1003,
         DP_OP_422J2_124_3477_n1002, DP_OP_422J2_124_3477_n1001,
         DP_OP_422J2_124_3477_n1000, DP_OP_422J2_124_3477_n999,
         DP_OP_422J2_124_3477_n998, DP_OP_422J2_124_3477_n997,
         DP_OP_422J2_124_3477_n996, DP_OP_422J2_124_3477_n995,
         DP_OP_422J2_124_3477_n994, DP_OP_422J2_124_3477_n993,
         DP_OP_422J2_124_3477_n992, DP_OP_422J2_124_3477_n991,
         DP_OP_422J2_124_3477_n990, DP_OP_422J2_124_3477_n989,
         DP_OP_422J2_124_3477_n988, DP_OP_422J2_124_3477_n987,
         DP_OP_422J2_124_3477_n986, DP_OP_422J2_124_3477_n985,
         DP_OP_422J2_124_3477_n984, DP_OP_422J2_124_3477_n983,
         DP_OP_422J2_124_3477_n982, DP_OP_422J2_124_3477_n981,
         DP_OP_422J2_124_3477_n980, DP_OP_422J2_124_3477_n979,
         DP_OP_422J2_124_3477_n978, DP_OP_422J2_124_3477_n977,
         DP_OP_422J2_124_3477_n976, DP_OP_422J2_124_3477_n975,
         DP_OP_422J2_124_3477_n974, DP_OP_422J2_124_3477_n973,
         DP_OP_422J2_124_3477_n972, DP_OP_422J2_124_3477_n971,
         DP_OP_422J2_124_3477_n970, DP_OP_422J2_124_3477_n969,
         DP_OP_422J2_124_3477_n968, DP_OP_422J2_124_3477_n967,
         DP_OP_422J2_124_3477_n966, DP_OP_422J2_124_3477_n965,
         DP_OP_422J2_124_3477_n964, DP_OP_422J2_124_3477_n963,
         DP_OP_422J2_124_3477_n962, DP_OP_422J2_124_3477_n961,
         DP_OP_422J2_124_3477_n960, DP_OP_422J2_124_3477_n959,
         DP_OP_422J2_124_3477_n958, DP_OP_422J2_124_3477_n957,
         DP_OP_422J2_124_3477_n956, DP_OP_422J2_124_3477_n955,
         DP_OP_422J2_124_3477_n954, DP_OP_422J2_124_3477_n953,
         DP_OP_422J2_124_3477_n952, DP_OP_422J2_124_3477_n951,
         DP_OP_422J2_124_3477_n950, DP_OP_422J2_124_3477_n949,
         DP_OP_422J2_124_3477_n948, DP_OP_422J2_124_3477_n947,
         DP_OP_422J2_124_3477_n946, DP_OP_422J2_124_3477_n945,
         DP_OP_422J2_124_3477_n944, DP_OP_422J2_124_3477_n943,
         DP_OP_422J2_124_3477_n942, DP_OP_422J2_124_3477_n941,
         DP_OP_422J2_124_3477_n940, DP_OP_422J2_124_3477_n939,
         DP_OP_422J2_124_3477_n938, DP_OP_422J2_124_3477_n937,
         DP_OP_422J2_124_3477_n936, DP_OP_422J2_124_3477_n935,
         DP_OP_422J2_124_3477_n934, DP_OP_422J2_124_3477_n933,
         DP_OP_422J2_124_3477_n932, DP_OP_422J2_124_3477_n931,
         DP_OP_422J2_124_3477_n930, DP_OP_422J2_124_3477_n929,
         DP_OP_422J2_124_3477_n928, DP_OP_422J2_124_3477_n927,
         DP_OP_422J2_124_3477_n926, DP_OP_422J2_124_3477_n925,
         DP_OP_422J2_124_3477_n924, DP_OP_422J2_124_3477_n923,
         DP_OP_422J2_124_3477_n922, DP_OP_422J2_124_3477_n921,
         DP_OP_422J2_124_3477_n920, DP_OP_422J2_124_3477_n919,
         DP_OP_422J2_124_3477_n918, DP_OP_422J2_124_3477_n917,
         DP_OP_422J2_124_3477_n916, DP_OP_422J2_124_3477_n915,
         DP_OP_422J2_124_3477_n914, DP_OP_422J2_124_3477_n913,
         DP_OP_422J2_124_3477_n912, DP_OP_422J2_124_3477_n911,
         DP_OP_422J2_124_3477_n910, DP_OP_422J2_124_3477_n909,
         DP_OP_422J2_124_3477_n908, DP_OP_422J2_124_3477_n907,
         DP_OP_422J2_124_3477_n906, DP_OP_422J2_124_3477_n905,
         DP_OP_422J2_124_3477_n904, DP_OP_422J2_124_3477_n903,
         DP_OP_422J2_124_3477_n902, DP_OP_422J2_124_3477_n901,
         DP_OP_422J2_124_3477_n900, DP_OP_422J2_124_3477_n899,
         DP_OP_422J2_124_3477_n898, DP_OP_422J2_124_3477_n897,
         DP_OP_422J2_124_3477_n896, DP_OP_422J2_124_3477_n895,
         DP_OP_422J2_124_3477_n894, DP_OP_422J2_124_3477_n893,
         DP_OP_422J2_124_3477_n892, DP_OP_422J2_124_3477_n891,
         DP_OP_422J2_124_3477_n890, DP_OP_422J2_124_3477_n889,
         DP_OP_422J2_124_3477_n888, DP_OP_422J2_124_3477_n887,
         DP_OP_422J2_124_3477_n886, DP_OP_422J2_124_3477_n885,
         DP_OP_422J2_124_3477_n884, DP_OP_422J2_124_3477_n883,
         DP_OP_422J2_124_3477_n882, DP_OP_422J2_124_3477_n881,
         DP_OP_422J2_124_3477_n880, DP_OP_422J2_124_3477_n879,
         DP_OP_422J2_124_3477_n878, DP_OP_422J2_124_3477_n877,
         DP_OP_422J2_124_3477_n876, DP_OP_422J2_124_3477_n875,
         DP_OP_422J2_124_3477_n874, DP_OP_422J2_124_3477_n873,
         DP_OP_422J2_124_3477_n872, DP_OP_422J2_124_3477_n871,
         DP_OP_422J2_124_3477_n870, DP_OP_422J2_124_3477_n869,
         DP_OP_422J2_124_3477_n868, DP_OP_422J2_124_3477_n867,
         DP_OP_422J2_124_3477_n866, DP_OP_422J2_124_3477_n865,
         DP_OP_422J2_124_3477_n864, DP_OP_422J2_124_3477_n863,
         DP_OP_422J2_124_3477_n862, DP_OP_422J2_124_3477_n861,
         DP_OP_422J2_124_3477_n860, DP_OP_422J2_124_3477_n859,
         DP_OP_422J2_124_3477_n858, DP_OP_422J2_124_3477_n857,
         DP_OP_422J2_124_3477_n856, DP_OP_422J2_124_3477_n855,
         DP_OP_422J2_124_3477_n854, DP_OP_422J2_124_3477_n853,
         DP_OP_422J2_124_3477_n852, DP_OP_422J2_124_3477_n851,
         DP_OP_422J2_124_3477_n850, DP_OP_422J2_124_3477_n849,
         DP_OP_422J2_124_3477_n848, DP_OP_422J2_124_3477_n847,
         DP_OP_422J2_124_3477_n846, DP_OP_422J2_124_3477_n845,
         DP_OP_422J2_124_3477_n844, DP_OP_422J2_124_3477_n843,
         DP_OP_422J2_124_3477_n842, DP_OP_422J2_124_3477_n841,
         DP_OP_422J2_124_3477_n840, DP_OP_422J2_124_3477_n839,
         DP_OP_422J2_124_3477_n838, DP_OP_422J2_124_3477_n837,
         DP_OP_422J2_124_3477_n836, DP_OP_422J2_124_3477_n835,
         DP_OP_422J2_124_3477_n834, DP_OP_422J2_124_3477_n833,
         DP_OP_422J2_124_3477_n832, DP_OP_422J2_124_3477_n831,
         DP_OP_422J2_124_3477_n830, DP_OP_422J2_124_3477_n829,
         DP_OP_422J2_124_3477_n828, DP_OP_422J2_124_3477_n827,
         DP_OP_422J2_124_3477_n826, DP_OP_422J2_124_3477_n825,
         DP_OP_422J2_124_3477_n824, DP_OP_422J2_124_3477_n823,
         DP_OP_422J2_124_3477_n822, DP_OP_422J2_124_3477_n821,
         DP_OP_422J2_124_3477_n820, DP_OP_422J2_124_3477_n819,
         DP_OP_422J2_124_3477_n818, DP_OP_422J2_124_3477_n817,
         DP_OP_422J2_124_3477_n816, DP_OP_422J2_124_3477_n815,
         DP_OP_422J2_124_3477_n814, DP_OP_422J2_124_3477_n813,
         DP_OP_422J2_124_3477_n812, DP_OP_422J2_124_3477_n811,
         DP_OP_422J2_124_3477_n810, DP_OP_422J2_124_3477_n809,
         DP_OP_422J2_124_3477_n808, DP_OP_422J2_124_3477_n807,
         DP_OP_422J2_124_3477_n806, DP_OP_422J2_124_3477_n805,
         DP_OP_422J2_124_3477_n804, DP_OP_422J2_124_3477_n803,
         DP_OP_422J2_124_3477_n802, DP_OP_422J2_124_3477_n801,
         DP_OP_422J2_124_3477_n800, DP_OP_422J2_124_3477_n799,
         DP_OP_422J2_124_3477_n798, DP_OP_422J2_124_3477_n797,
         DP_OP_422J2_124_3477_n796, DP_OP_422J2_124_3477_n795,
         DP_OP_422J2_124_3477_n794, DP_OP_422J2_124_3477_n793,
         DP_OP_422J2_124_3477_n792, DP_OP_422J2_124_3477_n791,
         DP_OP_422J2_124_3477_n790, DP_OP_422J2_124_3477_n789,
         DP_OP_422J2_124_3477_n788, DP_OP_422J2_124_3477_n787,
         DP_OP_422J2_124_3477_n786, DP_OP_422J2_124_3477_n785,
         DP_OP_422J2_124_3477_n784, DP_OP_422J2_124_3477_n783,
         DP_OP_422J2_124_3477_n782, DP_OP_422J2_124_3477_n781,
         DP_OP_422J2_124_3477_n780, DP_OP_422J2_124_3477_n779,
         DP_OP_422J2_124_3477_n778, DP_OP_422J2_124_3477_n777,
         DP_OP_422J2_124_3477_n776, DP_OP_422J2_124_3477_n775,
         DP_OP_422J2_124_3477_n774, DP_OP_422J2_124_3477_n773,
         DP_OP_422J2_124_3477_n772, DP_OP_422J2_124_3477_n771,
         DP_OP_422J2_124_3477_n770, DP_OP_422J2_124_3477_n769,
         DP_OP_422J2_124_3477_n768, DP_OP_422J2_124_3477_n767,
         DP_OP_422J2_124_3477_n766, DP_OP_422J2_124_3477_n765,
         DP_OP_422J2_124_3477_n764, DP_OP_422J2_124_3477_n763,
         DP_OP_422J2_124_3477_n762, DP_OP_422J2_124_3477_n761,
         DP_OP_422J2_124_3477_n760, DP_OP_422J2_124_3477_n759,
         DP_OP_422J2_124_3477_n758, DP_OP_422J2_124_3477_n757,
         DP_OP_422J2_124_3477_n756, DP_OP_422J2_124_3477_n755,
         DP_OP_422J2_124_3477_n754, DP_OP_422J2_124_3477_n753,
         DP_OP_422J2_124_3477_n752, DP_OP_422J2_124_3477_n751,
         DP_OP_422J2_124_3477_n750, DP_OP_422J2_124_3477_n749,
         DP_OP_422J2_124_3477_n748, DP_OP_422J2_124_3477_n747,
         DP_OP_422J2_124_3477_n746, DP_OP_422J2_124_3477_n745,
         DP_OP_422J2_124_3477_n744, DP_OP_422J2_124_3477_n743,
         DP_OP_422J2_124_3477_n742, DP_OP_422J2_124_3477_n741,
         DP_OP_422J2_124_3477_n740, DP_OP_422J2_124_3477_n739,
         DP_OP_422J2_124_3477_n738, DP_OP_422J2_124_3477_n737,
         DP_OP_422J2_124_3477_n736, DP_OP_422J2_124_3477_n735,
         DP_OP_422J2_124_3477_n734, DP_OP_422J2_124_3477_n733,
         DP_OP_422J2_124_3477_n732, DP_OP_422J2_124_3477_n731,
         DP_OP_422J2_124_3477_n730, DP_OP_422J2_124_3477_n729,
         DP_OP_422J2_124_3477_n728, DP_OP_422J2_124_3477_n727,
         DP_OP_422J2_124_3477_n726, DP_OP_422J2_124_3477_n725,
         DP_OP_422J2_124_3477_n724, DP_OP_422J2_124_3477_n723,
         DP_OP_422J2_124_3477_n722, DP_OP_422J2_124_3477_n721,
         DP_OP_422J2_124_3477_n720, DP_OP_422J2_124_3477_n719,
         DP_OP_422J2_124_3477_n718, DP_OP_422J2_124_3477_n717,
         DP_OP_422J2_124_3477_n716, DP_OP_422J2_124_3477_n715,
         DP_OP_422J2_124_3477_n714, DP_OP_422J2_124_3477_n713,
         DP_OP_422J2_124_3477_n712, DP_OP_422J2_124_3477_n711,
         DP_OP_422J2_124_3477_n710, DP_OP_422J2_124_3477_n709,
         DP_OP_422J2_124_3477_n708, DP_OP_422J2_124_3477_n707,
         DP_OP_422J2_124_3477_n706, DP_OP_422J2_124_3477_n705,
         DP_OP_422J2_124_3477_n704, DP_OP_422J2_124_3477_n703,
         DP_OP_422J2_124_3477_n702, DP_OP_422J2_124_3477_n701,
         DP_OP_422J2_124_3477_n700, DP_OP_422J2_124_3477_n699,
         DP_OP_422J2_124_3477_n698, DP_OP_422J2_124_3477_n697,
         DP_OP_422J2_124_3477_n696, DP_OP_422J2_124_3477_n695,
         DP_OP_422J2_124_3477_n694, DP_OP_422J2_124_3477_n693,
         DP_OP_422J2_124_3477_n692, DP_OP_422J2_124_3477_n691,
         DP_OP_422J2_124_3477_n690, DP_OP_422J2_124_3477_n689,
         DP_OP_422J2_124_3477_n688, DP_OP_422J2_124_3477_n687,
         DP_OP_422J2_124_3477_n686, DP_OP_422J2_124_3477_n685,
         DP_OP_422J2_124_3477_n684, DP_OP_422J2_124_3477_n683,
         DP_OP_422J2_124_3477_n682, DP_OP_422J2_124_3477_n681,
         DP_OP_422J2_124_3477_n680, DP_OP_422J2_124_3477_n679,
         DP_OP_422J2_124_3477_n678, DP_OP_422J2_124_3477_n677,
         DP_OP_422J2_124_3477_n676, DP_OP_422J2_124_3477_n675,
         DP_OP_422J2_124_3477_n674, DP_OP_422J2_124_3477_n673,
         DP_OP_422J2_124_3477_n672, DP_OP_422J2_124_3477_n671,
         DP_OP_422J2_124_3477_n670, DP_OP_422J2_124_3477_n669,
         DP_OP_422J2_124_3477_n668, DP_OP_422J2_124_3477_n667,
         DP_OP_422J2_124_3477_n666, DP_OP_422J2_124_3477_n665,
         DP_OP_422J2_124_3477_n664, DP_OP_422J2_124_3477_n663,
         DP_OP_422J2_124_3477_n662, DP_OP_422J2_124_3477_n661,
         DP_OP_422J2_124_3477_n660, DP_OP_422J2_124_3477_n659,
         DP_OP_422J2_124_3477_n658, DP_OP_422J2_124_3477_n657,
         DP_OP_422J2_124_3477_n656, DP_OP_422J2_124_3477_n655,
         DP_OP_422J2_124_3477_n654, DP_OP_422J2_124_3477_n653,
         DP_OP_422J2_124_3477_n652, DP_OP_422J2_124_3477_n651,
         DP_OP_422J2_124_3477_n650, DP_OP_422J2_124_3477_n649,
         DP_OP_422J2_124_3477_n648, DP_OP_422J2_124_3477_n647,
         DP_OP_422J2_124_3477_n646, DP_OP_422J2_124_3477_n645,
         DP_OP_422J2_124_3477_n644, DP_OP_422J2_124_3477_n643,
         DP_OP_422J2_124_3477_n642, DP_OP_422J2_124_3477_n641,
         DP_OP_422J2_124_3477_n640, DP_OP_422J2_124_3477_n639,
         DP_OP_422J2_124_3477_n638, DP_OP_422J2_124_3477_n637,
         DP_OP_422J2_124_3477_n636, DP_OP_422J2_124_3477_n635,
         DP_OP_422J2_124_3477_n634, DP_OP_422J2_124_3477_n633,
         DP_OP_422J2_124_3477_n632, DP_OP_422J2_124_3477_n631,
         DP_OP_422J2_124_3477_n630, DP_OP_422J2_124_3477_n629,
         DP_OP_422J2_124_3477_n628, DP_OP_422J2_124_3477_n627,
         DP_OP_422J2_124_3477_n626, DP_OP_422J2_124_3477_n625,
         DP_OP_422J2_124_3477_n624, DP_OP_422J2_124_3477_n623,
         DP_OP_422J2_124_3477_n622, DP_OP_422J2_124_3477_n621,
         DP_OP_422J2_124_3477_n620, DP_OP_422J2_124_3477_n619,
         DP_OP_422J2_124_3477_n618, DP_OP_422J2_124_3477_n617,
         DP_OP_422J2_124_3477_n616, DP_OP_422J2_124_3477_n615,
         DP_OP_422J2_124_3477_n614, DP_OP_422J2_124_3477_n613,
         DP_OP_422J2_124_3477_n612, DP_OP_422J2_124_3477_n611,
         DP_OP_422J2_124_3477_n610, DP_OP_422J2_124_3477_n609,
         DP_OP_422J2_124_3477_n608, DP_OP_422J2_124_3477_n607,
         DP_OP_422J2_124_3477_n606, DP_OP_422J2_124_3477_n605,
         DP_OP_422J2_124_3477_n604, DP_OP_422J2_124_3477_n603,
         DP_OP_422J2_124_3477_n602, DP_OP_422J2_124_3477_n601,
         DP_OP_422J2_124_3477_n600, DP_OP_422J2_124_3477_n599,
         DP_OP_422J2_124_3477_n598, DP_OP_422J2_124_3477_n597,
         DP_OP_422J2_124_3477_n596, DP_OP_422J2_124_3477_n595,
         DP_OP_422J2_124_3477_n594, DP_OP_422J2_124_3477_n593,
         DP_OP_422J2_124_3477_n592, DP_OP_422J2_124_3477_n591,
         DP_OP_422J2_124_3477_n590, DP_OP_422J2_124_3477_n589,
         DP_OP_422J2_124_3477_n588, DP_OP_422J2_124_3477_n587,
         DP_OP_422J2_124_3477_n586, DP_OP_422J2_124_3477_n585,
         DP_OP_422J2_124_3477_n584, DP_OP_422J2_124_3477_n583,
         DP_OP_422J2_124_3477_n582, DP_OP_422J2_124_3477_n581,
         DP_OP_422J2_124_3477_n580, DP_OP_422J2_124_3477_n579,
         DP_OP_422J2_124_3477_n578, DP_OP_422J2_124_3477_n577,
         DP_OP_422J2_124_3477_n576, DP_OP_422J2_124_3477_n575,
         DP_OP_422J2_124_3477_n574, DP_OP_422J2_124_3477_n573,
         DP_OP_422J2_124_3477_n572, DP_OP_422J2_124_3477_n571,
         DP_OP_422J2_124_3477_n570, DP_OP_422J2_124_3477_n569,
         DP_OP_422J2_124_3477_n568, DP_OP_422J2_124_3477_n567,
         DP_OP_422J2_124_3477_n566, DP_OP_422J2_124_3477_n565,
         DP_OP_422J2_124_3477_n564, DP_OP_422J2_124_3477_n563,
         DP_OP_422J2_124_3477_n562, DP_OP_422J2_124_3477_n561,
         DP_OP_422J2_124_3477_n560, DP_OP_422J2_124_3477_n559,
         DP_OP_422J2_124_3477_n558, DP_OP_422J2_124_3477_n557,
         DP_OP_422J2_124_3477_n556, DP_OP_422J2_124_3477_n555,
         DP_OP_422J2_124_3477_n554, DP_OP_422J2_124_3477_n553,
         DP_OP_422J2_124_3477_n552, DP_OP_422J2_124_3477_n551,
         DP_OP_422J2_124_3477_n550, DP_OP_422J2_124_3477_n549,
         DP_OP_422J2_124_3477_n548, DP_OP_422J2_124_3477_n547,
         DP_OP_422J2_124_3477_n546, DP_OP_422J2_124_3477_n545,
         DP_OP_422J2_124_3477_n544, DP_OP_422J2_124_3477_n543,
         DP_OP_422J2_124_3477_n542, DP_OP_422J2_124_3477_n541,
         DP_OP_422J2_124_3477_n540, DP_OP_422J2_124_3477_n539,
         DP_OP_422J2_124_3477_n538, DP_OP_422J2_124_3477_n537,
         DP_OP_422J2_124_3477_n536, DP_OP_422J2_124_3477_n535,
         DP_OP_422J2_124_3477_n534, DP_OP_422J2_124_3477_n533,
         DP_OP_422J2_124_3477_n532, DP_OP_422J2_124_3477_n531,
         DP_OP_422J2_124_3477_n530, DP_OP_422J2_124_3477_n529,
         DP_OP_422J2_124_3477_n528, DP_OP_422J2_124_3477_n527,
         DP_OP_422J2_124_3477_n526, DP_OP_422J2_124_3477_n525,
         DP_OP_422J2_124_3477_n524, DP_OP_422J2_124_3477_n523,
         DP_OP_422J2_124_3477_n522, DP_OP_422J2_124_3477_n521,
         DP_OP_422J2_124_3477_n520, DP_OP_422J2_124_3477_n519,
         DP_OP_422J2_124_3477_n518, DP_OP_422J2_124_3477_n517,
         DP_OP_422J2_124_3477_n516, DP_OP_422J2_124_3477_n515,
         DP_OP_422J2_124_3477_n514, DP_OP_422J2_124_3477_n513,
         DP_OP_422J2_124_3477_n512, DP_OP_422J2_124_3477_n511,
         DP_OP_422J2_124_3477_n510, DP_OP_422J2_124_3477_n509,
         DP_OP_422J2_124_3477_n508, DP_OP_422J2_124_3477_n507,
         DP_OP_422J2_124_3477_n506, DP_OP_422J2_124_3477_n505,
         DP_OP_422J2_124_3477_n504, DP_OP_422J2_124_3477_n503,
         DP_OP_422J2_124_3477_n502, DP_OP_422J2_124_3477_n501,
         DP_OP_422J2_124_3477_n500, DP_OP_422J2_124_3477_n499,
         DP_OP_422J2_124_3477_n498, DP_OP_422J2_124_3477_n497,
         DP_OP_422J2_124_3477_n496, DP_OP_422J2_124_3477_n495,
         DP_OP_422J2_124_3477_n494, DP_OP_422J2_124_3477_n493,
         DP_OP_422J2_124_3477_n492, DP_OP_422J2_124_3477_n491,
         DP_OP_422J2_124_3477_n490, DP_OP_422J2_124_3477_n489,
         DP_OP_422J2_124_3477_n488, DP_OP_422J2_124_3477_n487,
         DP_OP_422J2_124_3477_n486, DP_OP_422J2_124_3477_n485,
         DP_OP_422J2_124_3477_n484, DP_OP_422J2_124_3477_n483,
         DP_OP_422J2_124_3477_n482, DP_OP_422J2_124_3477_n481,
         DP_OP_422J2_124_3477_n480, DP_OP_422J2_124_3477_n479,
         DP_OP_422J2_124_3477_n478, DP_OP_422J2_124_3477_n477,
         DP_OP_422J2_124_3477_n476, DP_OP_422J2_124_3477_n475,
         DP_OP_422J2_124_3477_n474, DP_OP_422J2_124_3477_n473,
         DP_OP_422J2_124_3477_n472, DP_OP_422J2_124_3477_n471,
         DP_OP_422J2_124_3477_n470, DP_OP_422J2_124_3477_n469,
         DP_OP_422J2_124_3477_n468, DP_OP_422J2_124_3477_n467,
         DP_OP_422J2_124_3477_n466, DP_OP_422J2_124_3477_n465,
         DP_OP_422J2_124_3477_n464, DP_OP_422J2_124_3477_n463,
         DP_OP_422J2_124_3477_n462, DP_OP_422J2_124_3477_n461,
         DP_OP_422J2_124_3477_n460, DP_OP_422J2_124_3477_n459,
         DP_OP_422J2_124_3477_n458, DP_OP_422J2_124_3477_n457,
         DP_OP_422J2_124_3477_n456, DP_OP_422J2_124_3477_n455,
         DP_OP_422J2_124_3477_n454, DP_OP_422J2_124_3477_n453,
         DP_OP_422J2_124_3477_n452, DP_OP_422J2_124_3477_n451,
         DP_OP_422J2_124_3477_n450, DP_OP_422J2_124_3477_n449,
         DP_OP_422J2_124_3477_n448, DP_OP_422J2_124_3477_n447,
         DP_OP_422J2_124_3477_n446, DP_OP_422J2_124_3477_n445,
         DP_OP_422J2_124_3477_n444, DP_OP_422J2_124_3477_n443,
         DP_OP_422J2_124_3477_n442, DP_OP_422J2_124_3477_n441,
         DP_OP_422J2_124_3477_n440, DP_OP_422J2_124_3477_n439,
         DP_OP_422J2_124_3477_n438, DP_OP_422J2_124_3477_n437,
         DP_OP_422J2_124_3477_n436, DP_OP_422J2_124_3477_n435,
         DP_OP_422J2_124_3477_n434, DP_OP_422J2_124_3477_n433,
         DP_OP_422J2_124_3477_n432, DP_OP_422J2_124_3477_n431,
         DP_OP_422J2_124_3477_n430, DP_OP_422J2_124_3477_n429,
         DP_OP_422J2_124_3477_n428, DP_OP_422J2_124_3477_n427,
         DP_OP_422J2_124_3477_n426, DP_OP_422J2_124_3477_n425,
         DP_OP_422J2_124_3477_n424, DP_OP_422J2_124_3477_n423,
         DP_OP_422J2_124_3477_n422, DP_OP_422J2_124_3477_n421,
         DP_OP_422J2_124_3477_n420, DP_OP_422J2_124_3477_n419,
         DP_OP_422J2_124_3477_n418, DP_OP_422J2_124_3477_n417,
         DP_OP_422J2_124_3477_n416, DP_OP_422J2_124_3477_n415,
         DP_OP_422J2_124_3477_n414, DP_OP_422J2_124_3477_n413,
         DP_OP_422J2_124_3477_n412, DP_OP_422J2_124_3477_n411,
         DP_OP_422J2_124_3477_n410, DP_OP_422J2_124_3477_n409,
         DP_OP_422J2_124_3477_n408, DP_OP_422J2_124_3477_n407,
         DP_OP_422J2_124_3477_n406, DP_OP_422J2_124_3477_n405,
         DP_OP_422J2_124_3477_n404, DP_OP_422J2_124_3477_n403,
         DP_OP_422J2_124_3477_n402, DP_OP_422J2_124_3477_n401,
         DP_OP_422J2_124_3477_n400, DP_OP_422J2_124_3477_n399,
         DP_OP_422J2_124_3477_n398, DP_OP_422J2_124_3477_n397,
         DP_OP_422J2_124_3477_n396, DP_OP_422J2_124_3477_n395,
         DP_OP_422J2_124_3477_n394, DP_OP_422J2_124_3477_n393,
         DP_OP_422J2_124_3477_n392, DP_OP_422J2_124_3477_n391,
         DP_OP_422J2_124_3477_n390, DP_OP_422J2_124_3477_n389,
         DP_OP_422J2_124_3477_n388, DP_OP_422J2_124_3477_n387,
         DP_OP_422J2_124_3477_n386, DP_OP_422J2_124_3477_n385,
         DP_OP_422J2_124_3477_n384, DP_OP_422J2_124_3477_n383,
         DP_OP_422J2_124_3477_n382, DP_OP_422J2_124_3477_n381,
         DP_OP_422J2_124_3477_n380, DP_OP_422J2_124_3477_n379,
         DP_OP_422J2_124_3477_n378, DP_OP_422J2_124_3477_n377,
         DP_OP_422J2_124_3477_n376, DP_OP_422J2_124_3477_n375,
         DP_OP_422J2_124_3477_n374, DP_OP_422J2_124_3477_n373,
         DP_OP_422J2_124_3477_n372, DP_OP_422J2_124_3477_n371,
         DP_OP_422J2_124_3477_n370, DP_OP_422J2_124_3477_n369,
         DP_OP_422J2_124_3477_n368, DP_OP_422J2_124_3477_n367,
         DP_OP_422J2_124_3477_n366, DP_OP_422J2_124_3477_n365,
         DP_OP_422J2_124_3477_n364, DP_OP_422J2_124_3477_n363,
         DP_OP_422J2_124_3477_n362, DP_OP_422J2_124_3477_n361,
         DP_OP_422J2_124_3477_n360, DP_OP_422J2_124_3477_n359,
         DP_OP_422J2_124_3477_n358, DP_OP_422J2_124_3477_n357,
         DP_OP_422J2_124_3477_n356, DP_OP_422J2_124_3477_n355,
         DP_OP_422J2_124_3477_n354, DP_OP_422J2_124_3477_n353,
         DP_OP_422J2_124_3477_n352, DP_OP_422J2_124_3477_n351,
         DP_OP_422J2_124_3477_n350, DP_OP_422J2_124_3477_n349,
         DP_OP_422J2_124_3477_n348, DP_OP_422J2_124_3477_n347,
         DP_OP_422J2_124_3477_n346, DP_OP_422J2_124_3477_n345,
         DP_OP_422J2_124_3477_n344, DP_OP_422J2_124_3477_n343,
         DP_OP_422J2_124_3477_n342, DP_OP_422J2_124_3477_n341,
         DP_OP_422J2_124_3477_n340, DP_OP_422J2_124_3477_n339,
         DP_OP_422J2_124_3477_n338, DP_OP_422J2_124_3477_n337,
         DP_OP_422J2_124_3477_n336, DP_OP_422J2_124_3477_n335,
         DP_OP_422J2_124_3477_n334, DP_OP_422J2_124_3477_n333,
         DP_OP_422J2_124_3477_n332, DP_OP_422J2_124_3477_n331,
         DP_OP_422J2_124_3477_n330, DP_OP_422J2_124_3477_n329,
         DP_OP_422J2_124_3477_n328, DP_OP_422J2_124_3477_n327,
         DP_OP_422J2_124_3477_n326, DP_OP_422J2_124_3477_n325,
         DP_OP_422J2_124_3477_n324, DP_OP_422J2_124_3477_n323,
         DP_OP_422J2_124_3477_n322, DP_OP_422J2_124_3477_n321,
         DP_OP_422J2_124_3477_n320, DP_OP_422J2_124_3477_n319,
         DP_OP_422J2_124_3477_n318, DP_OP_422J2_124_3477_n317,
         DP_OP_422J2_124_3477_n316, DP_OP_422J2_124_3477_n315,
         DP_OP_422J2_124_3477_n314, DP_OP_422J2_124_3477_n313,
         DP_OP_422J2_124_3477_n312, DP_OP_422J2_124_3477_n311,
         DP_OP_422J2_124_3477_n310, DP_OP_422J2_124_3477_n309,
         DP_OP_422J2_124_3477_n308, DP_OP_422J2_124_3477_n307,
         DP_OP_422J2_124_3477_n306, DP_OP_422J2_124_3477_n305,
         DP_OP_422J2_124_3477_n304, DP_OP_422J2_124_3477_n303,
         DP_OP_422J2_124_3477_n302, DP_OP_422J2_124_3477_n301,
         DP_OP_422J2_124_3477_n300, DP_OP_422J2_124_3477_n299,
         DP_OP_422J2_124_3477_n298, DP_OP_422J2_124_3477_n297,
         DP_OP_422J2_124_3477_n296, DP_OP_422J2_124_3477_n295,
         DP_OP_422J2_124_3477_n294, DP_OP_422J2_124_3477_n293,
         DP_OP_422J2_124_3477_n292, DP_OP_422J2_124_3477_n291,
         DP_OP_422J2_124_3477_n290, DP_OP_422J2_124_3477_n289,
         DP_OP_422J2_124_3477_n288, DP_OP_422J2_124_3477_n287,
         DP_OP_422J2_124_3477_n286, DP_OP_422J2_124_3477_n285,
         DP_OP_422J2_124_3477_n284, DP_OP_422J2_124_3477_n283,
         DP_OP_422J2_124_3477_n282, DP_OP_422J2_124_3477_n281,
         DP_OP_422J2_124_3477_n280, DP_OP_422J2_124_3477_n279,
         DP_OP_422J2_124_3477_n278, DP_OP_422J2_124_3477_n277,
         DP_OP_422J2_124_3477_n276, DP_OP_422J2_124_3477_n275,
         DP_OP_422J2_124_3477_n274, DP_OP_422J2_124_3477_n273,
         DP_OP_422J2_124_3477_n272, DP_OP_422J2_124_3477_n271,
         DP_OP_422J2_124_3477_n270, DP_OP_422J2_124_3477_n269,
         DP_OP_422J2_124_3477_n268, DP_OP_422J2_124_3477_n267,
         DP_OP_422J2_124_3477_n266, DP_OP_422J2_124_3477_n265,
         DP_OP_422J2_124_3477_n264, DP_OP_422J2_124_3477_n263,
         DP_OP_422J2_124_3477_n262, DP_OP_422J2_124_3477_n261,
         DP_OP_422J2_124_3477_n260, DP_OP_422J2_124_3477_n259,
         DP_OP_422J2_124_3477_n258, DP_OP_422J2_124_3477_n257,
         DP_OP_422J2_124_3477_n256, DP_OP_422J2_124_3477_n255,
         DP_OP_422J2_124_3477_n254, DP_OP_422J2_124_3477_n253,
         DP_OP_422J2_124_3477_n252, DP_OP_422J2_124_3477_n241,
         DP_OP_422J2_124_3477_n240, DP_OP_422J2_124_3477_n237,
         DP_OP_422J2_124_3477_n236, DP_OP_422J2_124_3477_n233,
         DP_OP_422J2_124_3477_n231, DP_OP_422J2_124_3477_n229,
         DP_OP_422J2_124_3477_n227, DP_OP_422J2_124_3477_n219,
         DP_OP_422J2_124_3477_n218, DP_OP_422J2_124_3477_n217,
         DP_OP_422J2_124_3477_n216, DP_OP_422J2_124_3477_n215,
         DP_OP_422J2_124_3477_n211, DP_OP_422J2_124_3477_n210,
         DP_OP_422J2_124_3477_n209, DP_OP_422J2_124_3477_n208,
         DP_OP_422J2_124_3477_n207, DP_OP_422J2_124_3477_n203,
         DP_OP_422J2_124_3477_n202, DP_OP_422J2_124_3477_n201,
         DP_OP_422J2_124_3477_n200, DP_OP_422J2_124_3477_n199,
         DP_OP_422J2_124_3477_n195, DP_OP_422J2_124_3477_n194,
         DP_OP_422J2_124_3477_n193, DP_OP_422J2_124_3477_n192,
         DP_OP_422J2_124_3477_n191, DP_OP_422J2_124_3477_n190,
         DP_OP_422J2_124_3477_n189, DP_OP_422J2_124_3477_n187,
         DP_OP_422J2_124_3477_n186, DP_OP_422J2_124_3477_n185,
         DP_OP_422J2_124_3477_n184, DP_OP_422J2_124_3477_n183,
         DP_OP_422J2_124_3477_n182, DP_OP_422J2_124_3477_n181,
         DP_OP_422J2_124_3477_n180, DP_OP_422J2_124_3477_n179,
         DP_OP_422J2_124_3477_n177, DP_OP_422J2_124_3477_n176,
         DP_OP_422J2_124_3477_n175, DP_OP_422J2_124_3477_n174,
         DP_OP_422J2_124_3477_n173, DP_OP_422J2_124_3477_n172,
         DP_OP_422J2_124_3477_n171, DP_OP_422J2_124_3477_n170,
         DP_OP_422J2_124_3477_n168, DP_OP_422J2_124_3477_n167,
         DP_OP_422J2_124_3477_n166, DP_OP_422J2_124_3477_n165,
         DP_OP_422J2_124_3477_n164, DP_OP_422J2_124_3477_n163,
         DP_OP_422J2_124_3477_n162, DP_OP_422J2_124_3477_n161,
         DP_OP_422J2_124_3477_n158, DP_OP_422J2_124_3477_n152,
         DP_OP_422J2_124_3477_n151, DP_OP_422J2_124_3477_n150,
         DP_OP_422J2_124_3477_n149, DP_OP_422J2_124_3477_n148,
         DP_OP_422J2_124_3477_n145, DP_OP_422J2_124_3477_n144,
         DP_OP_422J2_124_3477_n143, DP_OP_422J2_124_3477_n142,
         DP_OP_422J2_124_3477_n141, DP_OP_422J2_124_3477_n140,
         DP_OP_422J2_124_3477_n137, DP_OP_422J2_124_3477_n136,
         DP_OP_422J2_124_3477_n135, DP_OP_422J2_124_3477_n133,
         DP_OP_422J2_124_3477_n132, DP_OP_422J2_124_3477_n130,
         DP_OP_422J2_124_3477_n129, DP_OP_422J2_124_3477_n128,
         DP_OP_422J2_124_3477_n127, DP_OP_422J2_124_3477_n126,
         DP_OP_422J2_124_3477_n125, DP_OP_422J2_124_3477_n123,
         DP_OP_422J2_124_3477_n119, DP_OP_422J2_124_3477_n118,
         DP_OP_422J2_124_3477_n116, DP_OP_422J2_124_3477_n115,
         DP_OP_422J2_124_3477_n114, DP_OP_422J2_124_3477_n113,
         DP_OP_422J2_124_3477_n112, DP_OP_422J2_124_3477_n111,
         DP_OP_422J2_124_3477_n109, DP_OP_422J2_124_3477_n105,
         DP_OP_422J2_124_3477_n104, DP_OP_422J2_124_3477_n102,
         DP_OP_422J2_124_3477_n101, DP_OP_422J2_124_3477_n100,
         DP_OP_422J2_124_3477_n99, DP_OP_422J2_124_3477_n98,
         DP_OP_422J2_124_3477_n97, DP_OP_422J2_124_3477_n95,
         DP_OP_422J2_124_3477_n91, DP_OP_422J2_124_3477_n90,
         DP_OP_422J2_124_3477_n88, DP_OP_422J2_124_3477_n87,
         DP_OP_422J2_124_3477_n86, DP_OP_422J2_124_3477_n85,
         DP_OP_422J2_124_3477_n84, DP_OP_422J2_124_3477_n83,
         DP_OP_422J2_124_3477_n81, DP_OP_422J2_124_3477_n76,
         DP_OP_422J2_124_3477_n75, DP_OP_422J2_124_3477_n74,
         DP_OP_422J2_124_3477_n73, DP_OP_422J2_124_3477_n72,
         DP_OP_422J2_124_3477_n70, DP_OP_422J2_124_3477_n65,
         DP_OP_422J2_124_3477_n63, DP_OP_422J2_124_3477_n62,
         DP_OP_422J2_124_3477_n61, DP_OP_422J2_124_3477_n59,
         DP_OP_422J2_124_3477_n58, DP_OP_422J2_124_3477_n57,
         DP_OP_422J2_124_3477_n56, DP_OP_422J2_124_3477_n55,
         DP_OP_422J2_124_3477_n52, DP_OP_422J2_124_3477_n48,
         DP_OP_422J2_124_3477_n47, DP_OP_422J2_124_3477_n45,
         DP_OP_422J2_124_3477_n44, DP_OP_422J2_124_3477_n43,
         DP_OP_422J2_124_3477_n42, DP_OP_422J2_124_3477_n41,
         DP_OP_422J2_124_3477_n40, DP_OP_422J2_124_3477_n39,
         DP_OP_422J2_124_3477_n37, DP_OP_422J2_124_3477_n25,
         DP_OP_422J2_124_3477_n22, DP_OP_422J2_124_3477_n21,
         DP_OP_422J2_124_3477_n4, DP_OP_422J2_124_3477_n3,
         DP_OP_422J2_124_3477_n2, n1, n2, n3, n4, n5010, n6, n7010, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n5000,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n7000, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n115, n117, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n139, n141, n142, n143, n144,
         n145, n147, n148, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n216, n217, n218, n219, n220, n221, n223, n224, n225, n226,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n5001, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n7001, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765;
  wire   [31:0] conv2_sum_a;
  wire   [31:0] conv2_sum_b;
  wire   [31:0] tmp_big1;
  wire   [31:0] conv2_sum_c;
  wire   [31:0] conv2_sum_d;
  wire   [31:0] tmp_big2;
  wire   [99:0] conv_weight_box;
  wire   [31:0] n_conv2_sum_a;
  wire   [31:0] n_conv2_sum_b;
  wire   [31:0] n_conv2_sum_c;
  wire   [31:0] n_conv2_sum_d;

  DFFSSRX1_HVT conv2_sum_c_reg_31_ ( .D(1'b0), .SETB(n383), .RSTB(
        n_conv2_sum_c[31]), .CLK(clk), .Q(conv2_sum_c[31]), .QN(n378) );
  DFFSSRX1_HVT conv2_sum_c_reg_30_ ( .D(1'b0), .SETB(n408), .RSTB(
        n_conv2_sum_c[30]), .CLK(clk), .Q(conv2_sum_c[30]), .QN(n528) );
  DFFSSRX1_HVT conv2_sum_c_reg_29_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_c[29]), .CLK(clk), .Q(conv2_sum_c[29]), .QN(n526) );
  DFFSSRX1_HVT conv2_sum_c_reg_28_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_c[28]), .CLK(clk), .Q(conv2_sum_c[28]), .QN(n522) );
  DFFSSRX1_HVT conv2_sum_c_reg_27_ ( .D(1'b0), .SETB(n382), .RSTB(
        n_conv2_sum_c[27]), .CLK(clk), .Q(conv2_sum_c[27]), .QN(n525) );
  DFFSSRX1_HVT conv2_sum_c_reg_26_ ( .D(1'b0), .SETB(n408), .RSTB(
        n_conv2_sum_c[26]), .CLK(clk), .Q(conv2_sum_c[26]), .QN(n521) );
  DFFSSRX1_HVT conv2_sum_c_reg_25_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_c[25]), .CLK(clk), .Q(conv2_sum_c[25]), .QN(n518) );
  DFFSSRX1_HVT conv2_sum_c_reg_24_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_c[24]), .CLK(clk), .Q(conv2_sum_c[24]), .QN(n504) );
  DFFSSRX1_HVT conv2_sum_c_reg_23_ ( .D(1'b0), .SETB(n383), .RSTB(
        n_conv2_sum_c[23]), .CLK(clk), .Q(conv2_sum_c[23]), .QN(n517) );
  DFFSSRX1_HVT conv2_sum_c_reg_22_ ( .D(1'b0), .SETB(n408), .RSTB(
        n_conv2_sum_c[22]), .CLK(clk), .Q(conv2_sum_c[22]), .QN(n503) );
  DFFSSRX1_HVT conv2_sum_c_reg_21_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_c[21]), .CLK(clk), .Q(conv2_sum_c[21]), .QN(n516) );
  DFFSSRX1_HVT conv2_sum_c_reg_20_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_c[20]), .CLK(clk), .Q(conv2_sum_c[20]), .QN(n502) );
  DFFSSRX1_HVT conv2_sum_c_reg_19_ ( .D(1'b0), .SETB(n382), .RSTB(
        n_conv2_sum_c[19]), .CLK(clk), .Q(conv2_sum_c[19]), .QN(n515) );
  DFFSSRX1_HVT conv2_sum_c_reg_18_ ( .D(1'b0), .SETB(n408), .RSTB(
        n_conv2_sum_c[18]), .CLK(clk), .Q(conv2_sum_c[18]), .QN(n485) );
  DFFSSRX1_HVT conv2_sum_c_reg_17_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_c[17]), .CLK(clk), .Q(conv2_sum_c[17]), .QN(n514) );
  DFFSSRX1_HVT conv2_sum_c_reg_16_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_c[16]), .CLK(clk), .Q(conv2_sum_c[16]), .QN(n338) );
  DFFSSRX1_HVT conv2_sum_c_reg_15_ ( .D(1'b0), .SETB(n383), .RSTB(
        n_conv2_sum_c[15]), .CLK(clk), .Q(conv2_sum_c[15]), .QN(n513) );
  DFFSSRX1_HVT conv2_sum_c_reg_14_ ( .D(1'b0), .SETB(n408), .RSTB(
        n_conv2_sum_c[14]), .CLK(clk), .Q(conv2_sum_c[14]), .QN(n501) );
  DFFSSRX1_HVT conv2_sum_c_reg_13_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_c[13]), .CLK(clk), .Q(conv2_sum_c[13]), .QN(n512) );
  DFFSSRX1_HVT conv2_sum_c_reg_12_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_c[12]), .CLK(clk), .Q(conv2_sum_c[12]), .QN(n5001) );
  DFFSSRX1_HVT conv2_sum_c_reg_11_ ( .D(1'b0), .SETB(n382), .RSTB(
        n_conv2_sum_c[11]), .CLK(clk), .Q(conv2_sum_c[11]), .QN(n476) );
  DFFSSRX1_HVT conv2_sum_c_reg_10_ ( .D(1'b0), .SETB(n408), .RSTB(
        n_conv2_sum_c[10]), .CLK(clk), .Q(conv2_sum_c[10]), .QN(n486) );
  DFFSSRX1_HVT conv2_sum_c_reg_9_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_c[9]), .CLK(clk), .Q(conv2_sum_c[9]), .QN(n489) );
  DFFSSRX1_HVT conv2_sum_c_reg_8_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_c[8]), .CLK(clk), .Q(conv2_sum_c[8]), .QN(n332) );
  DFFSSRX1_HVT conv2_sum_c_reg_7_ ( .D(1'b0), .SETB(n383), .RSTB(
        n_conv2_sum_c[7]), .CLK(clk), .Q(conv2_sum_c[7]), .QN(n475) );
  DFFSSRX1_HVT conv2_sum_c_reg_6_ ( .D(1'b0), .SETB(n408), .RSTB(
        n_conv2_sum_c[6]), .CLK(clk), .Q(conv2_sum_c[6]), .QN(n487) );
  DFFSSRX1_HVT conv2_sum_c_reg_5_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_c[5]), .CLK(clk), .Q(conv2_sum_c[5]), .QN(n474) );
  DFFSSRX1_HVT conv2_sum_c_reg_4_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_c[4]), .CLK(clk), .Q(conv2_sum_c[4]), .QN(n480) );
  DFFSSRX1_HVT conv2_sum_c_reg_3_ ( .D(1'b0), .SETB(n382), .RSTB(
        n_conv2_sum_c[3]), .CLK(clk), .Q(conv2_sum_c[3]), .QN(n490) );
  DFFSSRX1_HVT conv2_sum_c_reg_2_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_c[2]), .CLK(clk), .Q(conv2_sum_c[2]), .QN(n481) );
  DFFSSRX1_HVT conv2_sum_c_reg_1_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_c[1]), .CLK(clk), .Q(conv2_sum_c[1]), .QN(n544) );
  DFFSSRX1_HVT conv2_sum_c_reg_0_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_c[0]), .CLK(clk), .Q(conv2_sum_c[0]), .QN(n342) );
  DFFSSRX1_HVT conv2_sum_d_reg_31_ ( .D(1'b0), .SETB(n383), .RSTB(
        n_conv2_sum_d[31]), .CLK(clk), .Q(conv2_sum_d[31]), .QN(n530) );
  DFFSSRX1_HVT conv2_sum_d_reg_30_ ( .D(1'b0), .SETB(n408), .RSTB(
        n_conv2_sum_d[30]), .CLK(clk), .Q(conv2_sum_d[30]), .QN(n380) );
  DFFSSRX1_HVT conv2_sum_d_reg_29_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_d[29]), .CLK(clk), .Q(conv2_sum_d[29]), .QN(n376) );
  DFFSSRX1_HVT conv2_sum_d_reg_28_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_d[28]), .CLK(clk), .Q(conv2_sum_d[28]), .QN(n374) );
  DFFSSRX1_HVT conv2_sum_d_reg_27_ ( .D(1'b0), .SETB(n382), .RSTB(
        n_conv2_sum_d[27]), .CLK(clk), .Q(conv2_sum_d[27]), .QN(n370) );
  DFFSSRX1_HVT conv2_sum_d_reg_26_ ( .D(1'b0), .SETB(n408), .RSTB(
        n_conv2_sum_d[26]), .CLK(clk), .Q(conv2_sum_d[26]), .QN(n372) );
  DFFSSRX1_HVT conv2_sum_d_reg_25_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_d[25]), .CLK(clk), .Q(conv2_sum_d[25]), .QN(n360) );
  DFFSSRX1_HVT conv2_sum_d_reg_24_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_d[24]), .CLK(clk), .Q(conv2_sum_d[24]), .QN(n356) );
  DFFSSRX1_HVT conv2_sum_d_reg_23_ ( .D(1'b0), .SETB(n383), .RSTB(
        n_conv2_sum_d[23]), .CLK(clk), .Q(conv2_sum_d[23]), .QN(n349) );
  DFFSSRX1_HVT conv2_sum_d_reg_22_ ( .D(1'b0), .SETB(n408), .RSTB(
        n_conv2_sum_d[22]), .CLK(clk), .Q(conv2_sum_d[22]), .QN(n353) );
  DFFSSRX1_HVT conv2_sum_d_reg_21_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_d[21]), .CLK(clk), .Q(conv2_sum_d[21]), .QN(n359) );
  DFFSSRX1_HVT conv2_sum_d_reg_20_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_d[20]), .CLK(clk), .Q(conv2_sum_d[20]), .QN(n355) );
  DFFSSRX1_HVT conv2_sum_d_reg_19_ ( .D(1'b0), .SETB(n382), .RSTB(
        n_conv2_sum_d[19]), .CLK(clk), .Q(conv2_sum_d[19]), .QN(n352) );
  DFFSSRX1_HVT conv2_sum_d_reg_18_ ( .D(1'b0), .SETB(n408), .RSTB(
        n_conv2_sum_d[18]), .CLK(clk), .Q(conv2_sum_d[18]), .QN(n324) );
  DFFSSRX1_HVT conv2_sum_d_reg_17_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_d[17]), .CLK(clk), .Q(conv2_sum_d[17]), .QN(n339) );
  DFFSSRX1_HVT conv2_sum_d_reg_16_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_d[16]), .CLK(clk), .Q(conv2_sum_d[16]), .QN(n494) );
  DFFSSRX1_HVT conv2_sum_d_reg_15_ ( .D(1'b0), .SETB(n383), .RSTB(
        n_conv2_sum_d[15]), .CLK(clk), .Q(conv2_sum_d[15]), .QN(n350) );
  DFFSSRX1_HVT conv2_sum_d_reg_14_ ( .D(1'b0), .SETB(n408), .RSTB(
        n_conv2_sum_d[14]), .CLK(clk), .Q(conv2_sum_d[14]), .QN(n364) );
  DFFSSRX1_HVT conv2_sum_d_reg_13_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_d[13]), .CLK(clk), .Q(conv2_sum_d[13]), .QN(n368) );
  DFFSSRX1_HVT conv2_sum_d_reg_12_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_d[12]), .CLK(clk), .Q(conv2_sum_d[12]), .QN(n365) );
  DFFSSRX1_HVT conv2_sum_d_reg_11_ ( .D(1'b0), .SETB(n382), .RSTB(
        n_conv2_sum_d[11]), .CLK(clk), .Q(conv2_sum_d[11]), .QN(n323) );
  DFFSSRX1_HVT conv2_sum_d_reg_10_ ( .D(1'b0), .SETB(n408), .RSTB(
        n_conv2_sum_d[10]), .CLK(clk), .Q(conv2_sum_d[10]), .QN(n334) );
  DFFSSRX1_HVT conv2_sum_d_reg_9_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_d[9]), .CLK(clk), .Q(conv2_sum_d[9]), .QN(n340) );
  DFFSSRX1_HVT conv2_sum_d_reg_8_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_d[8]), .CLK(clk), .Q(conv2_sum_d[8]), .QN(n478) );
  DFFSSRX1_HVT conv2_sum_d_reg_7_ ( .D(1'b0), .SETB(n383), .RSTB(
        n_conv2_sum_d[7]), .CLK(clk), .Q(conv2_sum_d[7]), .QN(n318) );
  DFFSSRX1_HVT conv2_sum_d_reg_6_ ( .D(1'b0), .SETB(n408), .RSTB(
        n_conv2_sum_d[6]), .CLK(clk), .Q(conv2_sum_d[6]), .QN(n330) );
  DFFSSRX1_HVT conv2_sum_d_reg_5_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_d[5]), .CLK(clk), .Q(conv2_sum_d[5]), .QN(n321) );
  DFFSSRX1_HVT conv2_sum_d_reg_4_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_d[4]), .CLK(clk), .Q(conv2_sum_d[4]), .QN(n328) );
  DFFSSRX1_HVT conv2_sum_d_reg_3_ ( .D(1'b0), .SETB(n382), .RSTB(
        n_conv2_sum_d[3]), .CLK(clk), .Q(conv2_sum_d[3]), .QN(n538) );
  DFFSSRX1_HVT conv2_sum_d_reg_2_ ( .D(1'b0), .SETB(n408), .RSTB(
        n_conv2_sum_d[2]), .CLK(clk), .Q(conv2_sum_d[2]), .QN(n335) );
  DFFSSRX1_HVT conv2_sum_d_reg_1_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_d[1]), .CLK(clk), .QN(n543) );
  DFFSSRX1_HVT conv2_sum_d_reg_0_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_d[0]), .CLK(clk), .Q(conv2_sum_d[0]), .QN(n343) );
  DFFSSRX1_HVT conv2_sum_a_reg_31_ ( .D(1'b0), .SETB(n383), .RSTB(
        n_conv2_sum_a[31]), .CLK(clk), .Q(conv2_sum_a[31]), .QN(n377) );
  DFFSSRX1_HVT conv2_sum_a_reg_30_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_a[30]), .CLK(clk), .Q(conv2_sum_a[30]), .QN(n527) );
  DFFSSRX1_HVT conv2_sum_a_reg_29_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_a[29]), .CLK(clk), .Q(conv2_sum_a[29]), .QN(n524) );
  DFFSSRX1_HVT conv2_sum_a_reg_28_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_a[28]), .CLK(clk), .Q(conv2_sum_a[28]), .QN(n520) );
  DFFSSRX1_HVT conv2_sum_a_reg_27_ ( .D(1'b0), .SETB(n382), .RSTB(
        n_conv2_sum_a[27]), .CLK(clk), .Q(conv2_sum_a[27]), .QN(n523) );
  DFFSSRX1_HVT conv2_sum_a_reg_26_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_a[26]), .CLK(clk), .Q(conv2_sum_a[26]), .QN(n519) );
  DFFSSRX1_HVT conv2_sum_a_reg_25_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_a[25]), .CLK(clk), .Q(conv2_sum_a[25]), .QN(n511) );
  DFFSSRX1_HVT conv2_sum_a_reg_24_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_a[24]), .CLK(clk), .Q(conv2_sum_a[24]), .QN(n499) );
  DFFSSRX1_HVT conv2_sum_a_reg_23_ ( .D(1'b0), .SETB(n383), .RSTB(
        n_conv2_sum_a[23]), .CLK(clk), .Q(conv2_sum_a[23]), .QN(n510) );
  DFFSSRX1_HVT conv2_sum_a_reg_22_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_a[22]), .CLK(clk), .Q(conv2_sum_a[22]), .QN(n498) );
  DFFSSRX1_HVT conv2_sum_a_reg_21_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_a[21]), .CLK(clk), .Q(conv2_sum_a[21]), .QN(n509) );
  DFFSSRX1_HVT conv2_sum_a_reg_20_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_a[20]), .CLK(clk), .Q(conv2_sum_a[20]), .QN(n497) );
  DFFSSRX1_HVT conv2_sum_a_reg_19_ ( .D(1'b0), .SETB(n382), .RSTB(
        n_conv2_sum_a[19]), .CLK(clk), .Q(conv2_sum_a[19]), .QN(n508) );
  DFFSSRX1_HVT conv2_sum_a_reg_18_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_a[18]), .CLK(clk), .Q(conv2_sum_a[18]), .QN(n482) );
  DFFSSRX1_HVT conv2_sum_a_reg_17_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_a[17]), .CLK(clk), .Q(conv2_sum_a[17]), .QN(n507) );
  DFFSSRX1_HVT conv2_sum_a_reg_16_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_a[16]), .CLK(clk), .Q(conv2_sum_a[16]), .QN(n337) );
  DFFSSRX1_HVT conv2_sum_a_reg_15_ ( .D(1'b0), .SETB(n383), .RSTB(
        n_conv2_sum_a[15]), .CLK(clk), .Q(conv2_sum_a[15]), .QN(n506) );
  DFFSSRX1_HVT conv2_sum_a_reg_14_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_a[14]), .CLK(clk), .Q(conv2_sum_a[14]), .QN(n496) );
  DFFSSRX1_HVT conv2_sum_a_reg_13_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_a[13]), .CLK(clk), .Q(conv2_sum_a[13]), .QN(n505) );
  DFFSSRX1_HVT conv2_sum_a_reg_12_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_a[12]), .CLK(clk), .Q(conv2_sum_a[12]), .QN(n495) );
  DFFSSRX1_HVT conv2_sum_a_reg_11_ ( .D(1'b0), .SETB(n382), .RSTB(
        n_conv2_sum_a[11]), .CLK(clk), .Q(conv2_sum_a[11]), .QN(n539) );
  DFFSSRX1_HVT conv2_sum_a_reg_10_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_a[10]), .CLK(clk), .Q(conv2_sum_a[10]), .QN(n483) );
  DFFSSRX1_HVT conv2_sum_a_reg_9_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_a[9]), .CLK(clk), .Q(conv2_sum_a[9]), .QN(n549) );
  DFFSSRX1_HVT conv2_sum_a_reg_8_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_a[8]), .CLK(clk), .Q(conv2_sum_a[8]), .QN(n331) );
  DFFSSRX1_HVT conv2_sum_a_reg_7_ ( .D(1'b0), .SETB(n383), .RSTB(
        n_conv2_sum_a[7]), .CLK(clk), .Q(conv2_sum_a[7]), .QN(n473) );
  DFFSSRX1_HVT conv2_sum_a_reg_6_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_a[6]), .CLK(clk), .Q(conv2_sum_a[6]), .QN(n484) );
  DFFSSRX1_HVT conv2_sum_a_reg_5_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_a[5]), .CLK(clk), .Q(conv2_sum_a[5]), .QN(n472) );
  DFFSSRX1_HVT conv2_sum_a_reg_4_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_a[4]), .CLK(clk), .Q(conv2_sum_a[4]), .QN(n479) );
  DFFSSRX1_HVT conv2_sum_a_reg_3_ ( .D(1'b0), .SETB(n382), .RSTB(
        n_conv2_sum_a[3]), .CLK(clk), .QN(n545) );
  DFFSSRX1_HVT conv2_sum_a_reg_2_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_a[2]), .CLK(clk), .Q(conv2_sum_a[2]), .QN(n488) );
  DFFSSRX1_HVT conv2_sum_a_reg_1_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_a[1]), .CLK(clk), .Q(conv2_sum_a[1]), .QN(n345) );
  DFFSSRX1_HVT conv2_sum_a_reg_0_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_a[0]), .CLK(clk), .Q(conv2_sum_a[0]), .QN(n341) );
  DFFSSRX1_HVT conv2_sum_b_reg_31_ ( .D(1'b0), .SETB(n383), .RSTB(
        n_conv2_sum_b[31]), .CLK(clk), .Q(conv2_sum_b[31]), .QN(n529) );
  DFFSSRX1_HVT conv2_sum_b_reg_30_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_b[30]), .CLK(clk), .Q(conv2_sum_b[30]), .QN(n379) );
  DFFSSRX1_HVT conv2_sum_b_reg_29_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_b[29]), .CLK(clk), .Q(conv2_sum_b[29]), .QN(n375) );
  DFFSSRX1_HVT conv2_sum_b_reg_28_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_b[28]), .CLK(clk), .Q(conv2_sum_b[28]), .QN(n373) );
  DFFSSRX1_HVT conv2_sum_b_reg_27_ ( .D(1'b0), .SETB(n382), .RSTB(
        n_conv2_sum_b[27]), .CLK(clk), .Q(conv2_sum_b[27]), .QN(n369) );
  DFFSSRX1_HVT conv2_sum_b_reg_26_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_b[26]), .CLK(clk), .Q(conv2_sum_b[26]), .QN(n371) );
  DFFSSRX1_HVT conv2_sum_b_reg_25_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_b[25]), .CLK(clk), .Q(conv2_sum_b[25]), .QN(n361) );
  DFFSSRX1_HVT conv2_sum_b_reg_24_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_b[24]), .CLK(clk), .Q(conv2_sum_b[24]), .QN(n357) );
  DFFSSRX1_HVT conv2_sum_b_reg_23_ ( .D(1'b0), .SETB(n383), .RSTB(
        n_conv2_sum_b[23]), .CLK(clk), .Q(conv2_sum_b[23]), .QN(n347) );
  DFFSSRX1_HVT conv2_sum_b_reg_22_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_b[22]), .CLK(clk), .Q(conv2_sum_b[22]), .QN(n354) );
  DFFSSRX1_HVT conv2_sum_b_reg_21_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_b[21]), .CLK(clk), .Q(conv2_sum_b[21]), .QN(n362) );
  DFFSSRX1_HVT conv2_sum_b_reg_20_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_b[20]), .CLK(clk), .Q(conv2_sum_b[20]), .QN(n358) );
  DFFSSRX1_HVT conv2_sum_b_reg_19_ ( .D(1'b0), .SETB(n382), .RSTB(
        n_conv2_sum_b[19]), .CLK(clk), .Q(conv2_sum_b[19]), .QN(n348) );
  DFFSSRX1_HVT conv2_sum_b_reg_18_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_b[18]), .CLK(clk), .Q(conv2_sum_b[18]), .QN(n325) );
  DFFSSRX1_HVT conv2_sum_b_reg_17_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_b[17]), .CLK(clk), .Q(conv2_sum_b[17]), .QN(n333) );
  DFFSSRX1_HVT conv2_sum_b_reg_16_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_b[16]), .CLK(clk), .Q(conv2_sum_b[16]), .QN(n493) );
  DFFSSRX1_HVT conv2_sum_b_reg_15_ ( .D(1'b0), .SETB(n383), .RSTB(
        n_conv2_sum_b[15]), .CLK(clk), .Q(conv2_sum_b[15]), .QN(n351) );
  DFFSSRX1_HVT conv2_sum_b_reg_14_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_b[14]), .CLK(clk), .Q(conv2_sum_b[14]), .QN(n363) );
  DFFSSRX1_HVT conv2_sum_b_reg_13_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_b[13]), .CLK(clk), .Q(conv2_sum_b[13]), .QN(n367) );
  DFFSSRX1_HVT conv2_sum_b_reg_12_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_b[12]), .CLK(clk), .Q(conv2_sum_b[12]), .QN(n366) );
  DFFSSRX1_HVT conv2_sum_b_reg_11_ ( .D(1'b0), .SETB(n382), .RSTB(
        n_conv2_sum_b[11]), .CLK(clk), .Q(conv2_sum_b[11]), .QN(n322) );
  DFFSSRX1_HVT conv2_sum_b_reg_10_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_b[10]), .CLK(clk), .Q(conv2_sum_b[10]), .QN(n336) );
  DFFSSRX1_HVT conv2_sum_b_reg_9_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_b[9]), .CLK(clk), .Q(conv2_sum_b[9]), .QN(n548) );
  DFFSSRX1_HVT conv2_sum_b_reg_8_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_b[8]), .CLK(clk), .Q(conv2_sum_b[8]), .QN(n477) );
  DFFSSRX1_HVT conv2_sum_b_reg_7_ ( .D(1'b0), .SETB(n383), .RSTB(
        n_conv2_sum_b[7]), .CLK(clk), .Q(conv2_sum_b[7]), .QN(n319) );
  DFFSSRX1_HVT conv2_sum_b_reg_6_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_b[6]), .CLK(clk), .Q(conv2_sum_b[6]), .QN(n329) );
  DFFSSRX1_HVT conv2_sum_b_reg_5_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_b[5]), .CLK(clk), .Q(conv2_sum_b[5]), .QN(n320) );
  DFFSSRX1_HVT conv2_sum_b_reg_4_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_b[4]), .CLK(clk), .Q(conv2_sum_b[4]), .QN(n327) );
  DFFSSRX1_HVT conv2_sum_b_reg_3_ ( .D(1'b0), .SETB(n382), .RSTB(
        n_conv2_sum_b[3]), .CLK(clk), .Q(conv2_sum_b[3]), .QN(n466) );
  DFFSSRX1_HVT conv2_sum_b_reg_2_ ( .D(1'b0), .SETB(n405), .RSTB(
        n_conv2_sum_b[2]), .CLK(clk), .Q(conv2_sum_b[2]), .QN(n326) );
  DFFSSRX1_HVT conv2_sum_b_reg_1_ ( .D(1'b0), .SETB(n407), .RSTB(
        n_conv2_sum_b[1]), .CLK(clk), .Q(conv2_sum_b[1]), .QN(n546) );
  DFFSSRX1_HVT conv2_sum_b_reg_0_ ( .D(1'b0), .SETB(n406), .RSTB(
        n_conv2_sum_b[0]), .CLK(clk), .Q(conv2_sum_b[0]), .QN(n344) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U96 ( .A1(DP_OP_425J2_127_3477_n101), .A2(
        DP_OP_425J2_127_3477_n105), .A3(DP_OP_425J2_127_3477_n102), .Y(
        DP_OP_425J2_127_3477_n100) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U261 ( .A1(DP_OP_425J2_127_3477_n211), .A2(
        DP_OP_425J2_127_3477_n209), .A3(DP_OP_425J2_127_3477_n210), .Y(
        DP_OP_425J2_127_3477_n208) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U76 ( .A1(DP_OP_425J2_127_3477_n87), .A2(
        DP_OP_425J2_127_3477_n91), .A3(DP_OP_425J2_127_3477_n88), .Y(
        DP_OP_425J2_127_3477_n86) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U116 ( .A1(DP_OP_425J2_127_3477_n115), .A2(
        DP_OP_425J2_127_3477_n119), .A3(DP_OP_425J2_127_3477_n116), .Y(
        DP_OP_425J2_127_3477_n114) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U136 ( .A1(DP_OP_425J2_127_3477_n133), .A2(
        DP_OP_425J2_127_3477_n129), .A3(DP_OP_425J2_127_3477_n130), .Y(
        DP_OP_425J2_127_3477_n128) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U275 ( .A1(DP_OP_425J2_127_3477_n4), .A2(
        DP_OP_425J2_127_3477_n217), .A3(DP_OP_425J2_127_3477_n218), .Y(
        DP_OP_425J2_127_3477_n216) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1111 ( .A1(n364), .A2(
        DP_OP_424J2_126_3477_n2), .Y(DP_OP_425J2_127_3477_n288) );
  XNOR2X1_HVT DP_OP_425J2_127_3477_U737 ( .A1(DP_OP_425J2_127_3477_n2452), 
        .A2(DP_OP_425J2_127_3477_n2979), .Y(DP_OP_425J2_127_3477_n1161) );
  XNOR2X2_HVT DP_OP_425J2_127_3477_U131 ( .A1(DP_OP_425J2_127_3477_n131), .A2(
        DP_OP_425J2_127_3477_n18), .Y(n_conv2_sum_d[18]) );
  OAI21X2_HVT DP_OP_425J2_127_3477_U142 ( .A1(DP_OP_425J2_127_3477_n132), .A2(
        DP_OP_425J2_127_3477_n3), .A3(DP_OP_425J2_127_3477_n133), .Y(
        DP_OP_425J2_127_3477_n131) );
  XNOR2X2_HVT DP_OP_425J2_127_3477_U121 ( .A1(DP_OP_425J2_127_3477_n124), .A2(
        DP_OP_425J2_127_3477_n17), .Y(n_conv2_sum_d[19]) );
  OAI21X2_HVT DP_OP_425J2_127_3477_U132 ( .A1(DP_OP_425J2_127_3477_n125), .A2(
        DP_OP_425J2_127_3477_n3), .A3(DP_OP_425J2_127_3477_n126), .Y(
        DP_OP_425J2_127_3477_n124) );
  OAI21X2_HVT DP_OP_425J2_127_3477_U185 ( .A1(DP_OP_425J2_127_3477_n163), .A2(
        DP_OP_425J2_127_3477_n183), .A3(DP_OP_425J2_127_3477_n164), .Y(
        DP_OP_425J2_127_3477_n162) );
  OAI21X2_HVT DP_OP_425J2_127_3477_U203 ( .A1(DP_OP_425J2_127_3477_n181), .A2(
        DP_OP_425J2_127_3477_n175), .A3(DP_OP_425J2_127_3477_n176), .Y(
        DP_OP_425J2_127_3477_n174) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1109 ( .A1(n494), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_425J2_127_3477_n280) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2239 ( .A1(DP_OP_425J2_127_3477_n3006), .A2(
        DP_OP_425J2_127_3477_n3017), .Y(DP_OP_425J2_127_3477_n2998) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2231 ( .A1(DP_OP_425J2_127_3477_n3006), .A2(
        DP_OP_422J2_124_3477_n3016), .Y(DP_OP_425J2_127_3477_n2990) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2223 ( .A1(DP_OP_425J2_127_3477_n3006), .A2(
        DP_OP_425J2_127_3477_n3015), .Y(DP_OP_425J2_127_3477_n2982) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2222 ( .A1(DP_OP_425J2_127_3477_n3013), .A2(
        DP_OP_425J2_127_3477_n3014), .Y(DP_OP_425J2_127_3477_n1678) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2221 ( .A1(DP_OP_425J2_127_3477_n3012), .A2(
        DP_OP_425J2_127_3477_n3014), .Y(DP_OP_425J2_127_3477_n2981) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2220 ( .A1(DP_OP_425J2_127_3477_n3011), .A2(
        DP_OP_425J2_127_3477_n3014), .Y(DP_OP_425J2_127_3477_n2980) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2219 ( .A1(DP_OP_425J2_127_3477_n3010), .A2(
        DP_OP_425J2_127_3477_n3014), .Y(DP_OP_425J2_127_3477_n2979) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2218 ( .A1(DP_OP_425J2_127_3477_n3009), .A2(
        DP_OP_425J2_127_3477_n3014), .Y(DP_OP_425J2_127_3477_n2978) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2217 ( .A1(DP_OP_425J2_127_3477_n3008), .A2(
        DP_OP_425J2_127_3477_n3014), .Y(DP_OP_425J2_127_3477_n770) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2216 ( .A1(DP_OP_425J2_127_3477_n3007), .A2(
        DP_OP_425J2_127_3477_n3014), .Y(DP_OP_425J2_127_3477_n2977) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2215 ( .A1(DP_OP_425J2_127_3477_n3006), 
        .A2(DP_OP_425J2_127_3477_n3014), .Y(DP_OP_425J2_127_3477_n2976) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2195 ( .A1(DP_OP_425J2_127_3477_n2964), .A2(
        DP_OP_425J2_127_3477_n2975), .Y(DP_OP_425J2_127_3477_n2956) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2187 ( .A1(DP_OP_425J2_127_3477_n2964), .A2(
        DP_OP_425J2_127_3477_n2974), .Y(DP_OP_425J2_127_3477_n2948) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2179 ( .A1(DP_OP_425J2_127_3477_n2964), .A2(
        DP_OP_425J2_127_3477_n2973), .Y(DP_OP_425J2_127_3477_n2940) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2178 ( .A1(DP_OP_425J2_127_3477_n2971), .A2(
        DP_OP_425J2_127_3477_n2972), .Y(DP_OP_425J2_127_3477_n2939) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2177 ( .A1(DP_OP_424J2_126_3477_n1958), .A2(
        DP_OP_425J2_127_3477_n2972), .Y(DP_OP_425J2_127_3477_n2938) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2176 ( .A1(DP_OP_424J2_126_3477_n1957), .A2(
        DP_OP_425J2_127_3477_n2972), .Y(DP_OP_425J2_127_3477_n2937) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2175 ( .A1(DP_OP_424J2_126_3477_n1956), .A2(
        DP_OP_425J2_127_3477_n2972), .Y(DP_OP_425J2_127_3477_n2936) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2174 ( .A1(DP_OP_425J2_127_3477_n2967), .A2(
        DP_OP_425J2_127_3477_n2972), .Y(DP_OP_425J2_127_3477_n2935) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2173 ( .A1(DP_OP_424J2_126_3477_n1954), .A2(
        DP_OP_425J2_127_3477_n2972), .Y(DP_OP_425J2_127_3477_n2934) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2172 ( .A1(DP_OP_425J2_127_3477_n2965), .A2(
        DP_OP_425J2_127_3477_n2972), .Y(DP_OP_425J2_127_3477_n2933) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2171 ( .A1(DP_OP_425J2_127_3477_n2964), 
        .A2(DP_OP_425J2_127_3477_n2972), .Y(DP_OP_425J2_127_3477_n2932) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2151 ( .A1(DP_OP_425J2_127_3477_n2920), .A2(
        DP_OP_425J2_127_3477_n2931), .Y(DP_OP_425J2_127_3477_n2912) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2143 ( .A1(DP_OP_425J2_127_3477_n2920), .A2(
        DP_OP_425J2_127_3477_n2930), .Y(DP_OP_425J2_127_3477_n2904) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2135 ( .A1(DP_OP_425J2_127_3477_n2920), .A2(
        DP_OP_425J2_127_3477_n2929), .Y(DP_OP_425J2_127_3477_n2896) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2134 ( .A1(DP_OP_425J2_127_3477_n2927), .A2(
        DP_OP_425J2_127_3477_n2928), .Y(DP_OP_425J2_127_3477_n2895) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2133 ( .A1(DP_OP_425J2_127_3477_n2926), .A2(
        DP_OP_425J2_127_3477_n2928), .Y(DP_OP_425J2_127_3477_n2894) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2132 ( .A1(DP_OP_424J2_126_3477_n2001), .A2(
        DP_OP_425J2_127_3477_n2928), .Y(DP_OP_425J2_127_3477_n2893) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2131 ( .A1(DP_OP_425J2_127_3477_n2924), .A2(
        DP_OP_425J2_127_3477_n2928), .Y(DP_OP_425J2_127_3477_n2892) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2130 ( .A1(DP_OP_425J2_127_3477_n2923), .A2(
        DP_OP_425J2_127_3477_n2928), .Y(DP_OP_425J2_127_3477_n2891) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2129 ( .A1(DP_OP_425J2_127_3477_n2922), .A2(
        DP_OP_425J2_127_3477_n2928), .Y(DP_OP_425J2_127_3477_n2890) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2128 ( .A1(DP_OP_425J2_127_3477_n2921), .A2(
        DP_OP_425J2_127_3477_n2928), .Y(DP_OP_425J2_127_3477_n2889) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2127 ( .A1(DP_OP_425J2_127_3477_n2920), 
        .A2(DP_OP_425J2_127_3477_n2928), .Y(DP_OP_425J2_127_3477_n2888) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2107 ( .A1(DP_OP_423J2_125_3477_n1952), .A2(
        DP_OP_425J2_127_3477_n2887), .Y(DP_OP_425J2_127_3477_n2868) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2099 ( .A1(DP_OP_422J2_124_3477_n3006), .A2(
        DP_OP_422J2_124_3477_n2886), .Y(DP_OP_425J2_127_3477_n2860) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2092 ( .A1(DP_OP_425J2_127_3477_n2877), 
        .A2(DP_OP_422J2_124_3477_n2885), .Y(DP_OP_425J2_127_3477_n2853) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2091 ( .A1(DP_OP_423J2_125_3477_n1952), .A2(
        DP_OP_423J2_125_3477_n2885), .Y(DP_OP_425J2_127_3477_n2852) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2090 ( .A1(DP_OP_424J2_126_3477_n2047), .A2(
        DP_OP_425J2_127_3477_n2884), .Y(DP_OP_425J2_127_3477_n2851) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2089 ( .A1(DP_OP_422J2_124_3477_n3012), .A2(
        DP_OP_425J2_127_3477_n2884), .Y(DP_OP_425J2_127_3477_n2850) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2088 ( .A1(DP_OP_422J2_124_3477_n3011), .A2(
        DP_OP_425J2_127_3477_n2884), .Y(DP_OP_425J2_127_3477_n2849) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2087 ( .A1(DP_OP_422J2_124_3477_n3010), .A2(
        DP_OP_425J2_127_3477_n2884), .Y(DP_OP_425J2_127_3477_n2848) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2086 ( .A1(DP_OP_425J2_127_3477_n2879), .A2(
        DP_OP_425J2_127_3477_n2884), .Y(DP_OP_425J2_127_3477_n2847) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2085 ( .A1(DP_OP_425J2_127_3477_n2878), .A2(
        DP_OP_425J2_127_3477_n2884), .Y(DP_OP_425J2_127_3477_n2846) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2084 ( .A1(DP_OP_425J2_127_3477_n2877), .A2(
        DP_OP_425J2_127_3477_n2884), .Y(DP_OP_425J2_127_3477_n2845) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2083 ( .A1(DP_OP_422J2_124_3477_n3006), 
        .A2(DP_OP_425J2_127_3477_n2884), .Y(DP_OP_425J2_127_3477_n2844) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2063 ( .A1(DP_OP_422J2_124_3477_n2964), .A2(
        DP_OP_425J2_127_3477_n2843), .Y(DP_OP_425J2_127_3477_n2824) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2055 ( .A1(DP_OP_424J2_126_3477_n2084), .A2(
        DP_OP_425J2_127_3477_n2842), .Y(DP_OP_425J2_127_3477_n2816) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2048 ( .A1(DP_OP_425J2_127_3477_n2833), 
        .A2(DP_OP_425J2_127_3477_n2841), .Y(DP_OP_425J2_127_3477_n2809) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2047 ( .A1(DP_OP_422J2_124_3477_n2964), .A2(
        DP_OP_424J2_126_3477_n2841), .Y(DP_OP_425J2_127_3477_n2808) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2046 ( .A1(DP_OP_422J2_124_3477_n2971), .A2(
        DP_OP_425J2_127_3477_n2840), .Y(DP_OP_425J2_127_3477_n2807) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2045 ( .A1(DP_OP_422J2_124_3477_n2970), .A2(
        DP_OP_425J2_127_3477_n2840), .Y(DP_OP_425J2_127_3477_n2806) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2044 ( .A1(DP_OP_425J2_127_3477_n2837), .A2(
        DP_OP_425J2_127_3477_n2840), .Y(DP_OP_425J2_127_3477_n2805) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2043 ( .A1(DP_OP_423J2_125_3477_n2000), .A2(
        DP_OP_425J2_127_3477_n2840), .Y(DP_OP_425J2_127_3477_n2804) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2042 ( .A1(DP_OP_425J2_127_3477_n2835), .A2(
        DP_OP_425J2_127_3477_n2840), .Y(DP_OP_425J2_127_3477_n2803) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2041 ( .A1(DP_OP_425J2_127_3477_n2834), .A2(
        DP_OP_425J2_127_3477_n2840), .Y(DP_OP_425J2_127_3477_n2802) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2040 ( .A1(DP_OP_425J2_127_3477_n2833), .A2(
        DP_OP_425J2_127_3477_n2840), .Y(DP_OP_425J2_127_3477_n2801) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2039 ( .A1(DP_OP_424J2_126_3477_n2084), 
        .A2(DP_OP_425J2_127_3477_n2840), .Y(DP_OP_425J2_127_3477_n2800) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2019 ( .A1(DP_OP_423J2_125_3477_n2040), .A2(
        DP_OP_425J2_127_3477_n2799), .Y(DP_OP_425J2_127_3477_n2780) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2011 ( .A1(DP_OP_423J2_125_3477_n2040), .A2(
        DP_OP_425J2_127_3477_n2798), .Y(DP_OP_425J2_127_3477_n2772) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2004 ( .A1(DP_OP_425J2_127_3477_n2789), 
        .A2(DP_OP_425J2_127_3477_n2797), .Y(DP_OP_425J2_127_3477_n2765) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2003 ( .A1(DP_OP_423J2_125_3477_n2040), .A2(
        DP_OP_425J2_127_3477_n2797), .Y(DP_OP_425J2_127_3477_n2764) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2002 ( .A1(DP_OP_425J2_127_3477_n2795), .A2(
        DP_OP_425J2_127_3477_n2796), .Y(DP_OP_425J2_127_3477_n2763) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2001 ( .A1(DP_OP_425J2_127_3477_n2794), .A2(
        DP_OP_425J2_127_3477_n2796), .Y(DP_OP_425J2_127_3477_n2762) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2000 ( .A1(DP_OP_425J2_127_3477_n2793), .A2(
        DP_OP_425J2_127_3477_n2796), .Y(DP_OP_425J2_127_3477_n2761) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1999 ( .A1(DP_OP_423J2_125_3477_n2044), .A2(
        DP_OP_425J2_127_3477_n2796), .Y(DP_OP_425J2_127_3477_n2760) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1998 ( .A1(DP_OP_425J2_127_3477_n2791), .A2(
        DP_OP_425J2_127_3477_n2796), .Y(DP_OP_425J2_127_3477_n2759) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1997 ( .A1(DP_OP_425J2_127_3477_n2790), .A2(
        DP_OP_425J2_127_3477_n2796), .Y(DP_OP_425J2_127_3477_n2758) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1996 ( .A1(DP_OP_425J2_127_3477_n2789), .A2(
        DP_OP_425J2_127_3477_n2796), .Y(DP_OP_425J2_127_3477_n2757) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1995 ( .A1(DP_OP_423J2_125_3477_n2040), 
        .A2(DP_OP_425J2_127_3477_n2796), .Y(DP_OP_425J2_127_3477_n2756) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1982 ( .A1(DP_OP_422J2_124_3477_n2883), 
        .A2(DP_OP_425J2_127_3477_n2755), .Y(DP_OP_425J2_127_3477_n2743) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1981 ( .A1(DP_OP_425J2_127_3477_n2750), 
        .A2(DP_OP_425J2_127_3477_n2755), .Y(DP_OP_425J2_127_3477_n2742) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1980 ( .A1(DP_OP_425J2_127_3477_n2749), 
        .A2(DP_OP_425J2_127_3477_n2755), .Y(DP_OP_425J2_127_3477_n2741) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1979 ( .A1(DP_OP_422J2_124_3477_n2880), 
        .A2(DP_OP_425J2_127_3477_n2755), .Y(DP_OP_425J2_127_3477_n2740) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1978 ( .A1(DP_OP_425J2_127_3477_n2747), 
        .A2(DP_OP_425J2_127_3477_n2755), .Y(DP_OP_425J2_127_3477_n2739) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1977 ( .A1(DP_OP_423J2_125_3477_n2086), 
        .A2(DP_OP_425J2_127_3477_n2755), .Y(DP_OP_425J2_127_3477_n2738) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1976 ( .A1(DP_OP_425J2_127_3477_n2745), 
        .A2(DP_OP_425J2_127_3477_n2755), .Y(DP_OP_425J2_127_3477_n2737) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1975 ( .A1(DP_OP_423J2_125_3477_n2084), .A2(
        DP_OP_425J2_127_3477_n2755), .Y(DP_OP_425J2_127_3477_n2736) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1967 ( .A1(DP_OP_423J2_125_3477_n2084), .A2(
        DP_OP_425J2_127_3477_n2754), .Y(DP_OP_425J2_127_3477_n2728) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1959 ( .A1(DP_OP_423J2_125_3477_n2084), .A2(
        DP_OP_423J2_125_3477_n2753), .Y(DP_OP_425J2_127_3477_n2720) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1958 ( .A1(DP_OP_422J2_124_3477_n2883), .A2(
        DP_OP_425J2_127_3477_n2752), .Y(DP_OP_425J2_127_3477_n2719) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1957 ( .A1(DP_OP_425J2_127_3477_n2750), .A2(
        DP_OP_425J2_127_3477_n2752), .Y(DP_OP_425J2_127_3477_n2718) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1956 ( .A1(DP_OP_425J2_127_3477_n2749), .A2(
        DP_OP_425J2_127_3477_n2752), .Y(DP_OP_425J2_127_3477_n2717) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1955 ( .A1(DP_OP_423J2_125_3477_n2088), .A2(
        DP_OP_425J2_127_3477_n2752), .Y(DP_OP_425J2_127_3477_n2716) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1954 ( .A1(DP_OP_425J2_127_3477_n2747), .A2(
        DP_OP_425J2_127_3477_n2752), .Y(DP_OP_425J2_127_3477_n2715) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1953 ( .A1(DP_OP_423J2_125_3477_n2086), .A2(
        DP_OP_425J2_127_3477_n2752), .Y(DP_OP_425J2_127_3477_n2714) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1952 ( .A1(DP_OP_425J2_127_3477_n2745), .A2(
        DP_OP_425J2_127_3477_n2752), .Y(DP_OP_425J2_127_3477_n2713) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1951 ( .A1(DP_OP_423J2_125_3477_n2084), 
        .A2(DP_OP_425J2_127_3477_n2752), .Y(DP_OP_425J2_127_3477_n2712) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1931 ( .A1(DP_OP_425J2_127_3477_n2700), .A2(
        DP_OP_425J2_127_3477_n2711), .Y(DP_OP_425J2_127_3477_n2692) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1923 ( .A1(DP_OP_425J2_127_3477_n2700), .A2(
        DP_OP_425J2_127_3477_n2710), .Y(DP_OP_425J2_127_3477_n2684) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1916 ( .A1(DP_OP_422J2_124_3477_n2833), 
        .A2(DP_OP_425J2_127_3477_n2709), .Y(DP_OP_425J2_127_3477_n2677) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1915 ( .A1(DP_OP_425J2_127_3477_n2700), .A2(
        DP_OP_425J2_127_3477_n2709), .Y(DP_OP_425J2_127_3477_n2676) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1914 ( .A1(DP_OP_425J2_127_3477_n2707), .A2(
        DP_OP_425J2_127_3477_n2708), .Y(DP_OP_425J2_127_3477_n2675) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1913 ( .A1(DP_OP_422J2_124_3477_n2838), .A2(
        DP_OP_425J2_127_3477_n2708), .Y(DP_OP_425J2_127_3477_n2674) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1912 ( .A1(DP_OP_425J2_127_3477_n2705), .A2(
        DP_OP_425J2_127_3477_n2708), .Y(DP_OP_425J2_127_3477_n2673) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1911 ( .A1(DP_OP_425J2_127_3477_n2704), .A2(
        DP_OP_425J2_127_3477_n2708), .Y(DP_OP_425J2_127_3477_n2672) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1910 ( .A1(DP_OP_424J2_126_3477_n2219), .A2(
        DP_OP_425J2_127_3477_n2708), .Y(DP_OP_425J2_127_3477_n2671) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1909 ( .A1(DP_OP_424J2_126_3477_n2218), .A2(
        DP_OP_425J2_127_3477_n2708), .Y(DP_OP_425J2_127_3477_n2670) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1908 ( .A1(DP_OP_422J2_124_3477_n2833), .A2(
        DP_OP_425J2_127_3477_n2708), .Y(DP_OP_425J2_127_3477_n2669) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1907 ( .A1(DP_OP_425J2_127_3477_n2700), 
        .A2(DP_OP_425J2_127_3477_n2708), .Y(DP_OP_425J2_127_3477_n2668) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1888 ( .A1(DP_OP_424J2_126_3477_n2261), 
        .A2(DP_OP_425J2_127_3477_n2667), .Y(DP_OP_425J2_127_3477_n2649) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1887 ( .A1(DP_OP_423J2_125_3477_n2172), .A2(
        DP_OP_425J2_127_3477_n2667), .Y(DP_OP_425J2_127_3477_n2648) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1879 ( .A1(DP_OP_424J2_126_3477_n2260), .A2(
        DP_OP_425J2_127_3477_n2666), .Y(DP_OP_425J2_127_3477_n2640) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1871 ( .A1(DP_OP_423J2_125_3477_n2172), .A2(
        DP_OP_425J2_127_3477_n2665), .Y(DP_OP_425J2_127_3477_n2632) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1870 ( .A1(DP_OP_425J2_127_3477_n2663), .A2(
        DP_OP_425J2_127_3477_n2664), .Y(DP_OP_425J2_127_3477_n2631) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1869 ( .A1(DP_OP_425J2_127_3477_n2662), .A2(
        DP_OP_425J2_127_3477_n2664), .Y(DP_OP_425J2_127_3477_n2630) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1868 ( .A1(DP_OP_424J2_126_3477_n2265), .A2(
        DP_OP_425J2_127_3477_n2664), .Y(DP_OP_425J2_127_3477_n2629) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1867 ( .A1(DP_OP_422J2_124_3477_n2792), .A2(
        DP_OP_425J2_127_3477_n2664), .Y(DP_OP_425J2_127_3477_n2628) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1866 ( .A1(DP_OP_423J2_125_3477_n2175), .A2(
        DP_OP_425J2_127_3477_n2664), .Y(DP_OP_425J2_127_3477_n2627) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1865 ( .A1(DP_OP_425J2_127_3477_n2658), .A2(
        DP_OP_425J2_127_3477_n2664), .Y(DP_OP_425J2_127_3477_n2626) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1864 ( .A1(DP_OP_422J2_124_3477_n2789), .A2(
        DP_OP_425J2_127_3477_n2664), .Y(DP_OP_425J2_127_3477_n2625) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1863 ( .A1(DP_OP_424J2_126_3477_n2260), 
        .A2(DP_OP_425J2_127_3477_n2664), .Y(DP_OP_425J2_127_3477_n2624) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1843 ( .A1(DP_OP_425J2_127_3477_n2612), .A2(
        DP_OP_425J2_127_3477_n2623), .Y(DP_OP_425J2_127_3477_n2604) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1842 ( .A1(DP_OP_425J2_127_3477_n2619), 
        .A2(DP_OP_425J2_127_3477_n2622), .Y(DP_OP_425J2_127_3477_n2603) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1841 ( .A1(DP_OP_424J2_126_3477_n2310), 
        .A2(DP_OP_425J2_127_3477_n2622), .Y(DP_OP_425J2_127_3477_n2602) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1840 ( .A1(DP_OP_425J2_127_3477_n2617), 
        .A2(DP_OP_425J2_127_3477_n2622), .Y(DP_OP_425J2_127_3477_n2601) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1839 ( .A1(DP_OP_425J2_127_3477_n2616), 
        .A2(DP_OP_425J2_127_3477_n2622), .Y(DP_OP_425J2_127_3477_n2600) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1838 ( .A1(DP_OP_423J2_125_3477_n2219), 
        .A2(DP_OP_425J2_127_3477_n2622), .Y(DP_OP_425J2_127_3477_n2599) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1837 ( .A1(DP_OP_422J2_124_3477_n2746), 
        .A2(DP_OP_425J2_127_3477_n2622), .Y(DP_OP_425J2_127_3477_n2598) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1836 ( .A1(DP_OP_422J2_124_3477_n2745), 
        .A2(DP_OP_425J2_127_3477_n2622), .Y(DP_OP_425J2_127_3477_n2597) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1835 ( .A1(DP_OP_425J2_127_3477_n2612), .A2(
        DP_OP_425J2_127_3477_n2622), .Y(DP_OP_425J2_127_3477_n2596) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1827 ( .A1(DP_OP_425J2_127_3477_n2612), .A2(
        DP_OP_425J2_127_3477_n2621), .Y(DP_OP_425J2_127_3477_n2588) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1826 ( .A1(DP_OP_425J2_127_3477_n2619), .A2(
        DP_OP_425J2_127_3477_n2620), .Y(DP_OP_425J2_127_3477_n2587) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1825 ( .A1(DP_OP_424J2_126_3477_n2310), .A2(
        DP_OP_425J2_127_3477_n2620), .Y(DP_OP_425J2_127_3477_n2586) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1824 ( .A1(DP_OP_425J2_127_3477_n2617), .A2(
        DP_OP_425J2_127_3477_n2620), .Y(DP_OP_425J2_127_3477_n2585) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1823 ( .A1(DP_OP_425J2_127_3477_n2616), .A2(
        DP_OP_425J2_127_3477_n2620), .Y(DP_OP_425J2_127_3477_n2584) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1822 ( .A1(DP_OP_423J2_125_3477_n2219), .A2(
        DP_OP_425J2_127_3477_n2620), .Y(DP_OP_425J2_127_3477_n2583) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1821 ( .A1(DP_OP_422J2_124_3477_n2746), .A2(
        DP_OP_425J2_127_3477_n2620), .Y(DP_OP_425J2_127_3477_n2582) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1820 ( .A1(DP_OP_422J2_124_3477_n2745), .A2(
        DP_OP_425J2_127_3477_n2620), .Y(DP_OP_425J2_127_3477_n2581) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1819 ( .A1(DP_OP_425J2_127_3477_n2612), 
        .A2(DP_OP_425J2_127_3477_n2620), .Y(DP_OP_425J2_127_3477_n2580) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1800 ( .A1(DP_OP_423J2_125_3477_n2261), 
        .A2(DP_OP_425J2_127_3477_n2579), .Y(DP_OP_425J2_127_3477_n2561) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1799 ( .A1(DP_OP_423J2_125_3477_n2260), .A2(
        DP_OP_425J2_127_3477_n2579), .Y(DP_OP_425J2_127_3477_n2560) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1791 ( .A1(DP_OP_423J2_125_3477_n2260), .A2(
        DP_OP_425J2_127_3477_n2578), .Y(DP_OP_425J2_127_3477_n2552) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1783 ( .A1(DP_OP_423J2_125_3477_n2260), .A2(
        DP_OP_425J2_127_3477_n2577), .Y(DP_OP_425J2_127_3477_n2544) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1782 ( .A1(DP_OP_423J2_125_3477_n2267), .A2(
        DP_OP_425J2_127_3477_n2576), .Y(DP_OP_425J2_127_3477_n2543) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1781 ( .A1(DP_OP_423J2_125_3477_n2266), .A2(
        DP_OP_425J2_127_3477_n2576), .Y(DP_OP_425J2_127_3477_n2542) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1780 ( .A1(DP_OP_423J2_125_3477_n2265), .A2(
        DP_OP_425J2_127_3477_n2576), .Y(DP_OP_425J2_127_3477_n2541) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1779 ( .A1(DP_OP_425J2_127_3477_n2572), .A2(
        DP_OP_425J2_127_3477_n2576), .Y(DP_OP_425J2_127_3477_n2540) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1778 ( .A1(DP_OP_423J2_125_3477_n2263), .A2(
        DP_OP_425J2_127_3477_n2576), .Y(DP_OP_425J2_127_3477_n2539) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1777 ( .A1(DP_OP_423J2_125_3477_n2262), .A2(
        DP_OP_425J2_127_3477_n2576), .Y(DP_OP_425J2_127_3477_n2538) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1776 ( .A1(DP_OP_423J2_125_3477_n2261), .A2(
        DP_OP_425J2_127_3477_n2576), .Y(DP_OP_425J2_127_3477_n2537) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1775 ( .A1(DP_OP_423J2_125_3477_n2260), 
        .A2(DP_OP_425J2_127_3477_n2576), .Y(DP_OP_425J2_127_3477_n2536) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1755 ( .A1(DP_OP_422J2_124_3477_n2656), .A2(
        DP_OP_425J2_127_3477_n2535), .Y(DP_OP_425J2_127_3477_n2516) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1747 ( .A1(DP_OP_422J2_124_3477_n2656), .A2(
        DP_OP_425J2_127_3477_n2534), .Y(DP_OP_425J2_127_3477_n2508) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1740 ( .A1(DP_OP_425J2_127_3477_n2525), 
        .A2(DP_OP_423J2_125_3477_n2533), .Y(DP_OP_425J2_127_3477_n2501) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1739 ( .A1(DP_OP_422J2_124_3477_n2656), .A2(
        DP_OP_423J2_125_3477_n2533), .Y(DP_OP_425J2_127_3477_n2500) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1738 ( .A1(DP_OP_423J2_125_3477_n2311), .A2(
        DP_OP_424J2_126_3477_n2532), .Y(DP_OP_425J2_127_3477_n2499) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1737 ( .A1(DP_OP_425J2_127_3477_n2530), .A2(
        DP_OP_422J2_124_3477_n2532), .Y(DP_OP_425J2_127_3477_n2498) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1736 ( .A1(DP_OP_425J2_127_3477_n2529), .A2(
        DP_OP_423J2_125_3477_n2532), .Y(DP_OP_425J2_127_3477_n2497) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1735 ( .A1(DP_OP_425J2_127_3477_n2528), .A2(
        DP_OP_423J2_125_3477_n2532), .Y(DP_OP_425J2_127_3477_n2496) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1734 ( .A1(DP_OP_422J2_124_3477_n2659), .A2(
        DP_OP_422J2_124_3477_n2532), .Y(DP_OP_425J2_127_3477_n2495) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1733 ( .A1(DP_OP_425J2_127_3477_n2526), .A2(
        DP_OP_424J2_126_3477_n2532), .Y(DP_OP_425J2_127_3477_n2494) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1732 ( .A1(DP_OP_425J2_127_3477_n2525), .A2(
        DP_OP_422J2_124_3477_n2532), .Y(DP_OP_425J2_127_3477_n2493) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1731 ( .A1(DP_OP_422J2_124_3477_n2656), 
        .A2(DP_OP_424J2_126_3477_n2532), .Y(DP_OP_425J2_127_3477_n2492) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1711 ( .A1(DP_OP_422J2_124_3477_n2612), .A2(
        DP_OP_425J2_127_3477_n2491), .Y(DP_OP_425J2_127_3477_n2472) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1703 ( .A1(DP_OP_423J2_125_3477_n2348), .A2(
        DP_OP_425J2_127_3477_n2490), .Y(DP_OP_425J2_127_3477_n2464) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1695 ( .A1(DP_OP_423J2_125_3477_n2348), .A2(
        DP_OP_425J2_127_3477_n2489), .Y(DP_OP_425J2_127_3477_n2456) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1694 ( .A1(DP_OP_423J2_125_3477_n2355), .A2(
        DP_OP_425J2_127_3477_n2488), .Y(DP_OP_425J2_127_3477_n2455) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1693 ( .A1(DP_OP_423J2_125_3477_n2354), .A2(
        DP_OP_425J2_127_3477_n2488), .Y(DP_OP_425J2_127_3477_n2454) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1692 ( .A1(DP_OP_423J2_125_3477_n2353), .A2(
        DP_OP_425J2_127_3477_n2488), .Y(DP_OP_425J2_127_3477_n2453) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1691 ( .A1(DP_OP_425J2_127_3477_n2484), .A2(
        DP_OP_425J2_127_3477_n2488), .Y(DP_OP_425J2_127_3477_n2452) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1690 ( .A1(DP_OP_424J2_126_3477_n2439), .A2(
        DP_OP_425J2_127_3477_n2488), .Y(DP_OP_425J2_127_3477_n2451) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1689 ( .A1(DP_OP_425J2_127_3477_n2482), .A2(
        DP_OP_425J2_127_3477_n2488), .Y(DP_OP_425J2_127_3477_n2450) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1688 ( .A1(DP_OP_425J2_127_3477_n2481), .A2(
        DP_OP_425J2_127_3477_n2488), .Y(DP_OP_425J2_127_3477_n2449) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1687 ( .A1(DP_OP_423J2_125_3477_n2348), 
        .A2(DP_OP_425J2_127_3477_n2488), .Y(DP_OP_425J2_127_3477_n2448) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1667 ( .A1(DP_OP_423J2_125_3477_n2612), .A2(
        DP_OP_425J2_127_3477_n2447), .Y(DP_OP_425J2_127_3477_n2428) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1659 ( .A1(DP_OP_423J2_125_3477_n2612), .A2(
        DP_OP_425J2_127_3477_n2446), .Y(DP_OP_425J2_127_3477_n2420) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1651 ( .A1(DP_OP_423J2_125_3477_n2612), .A2(
        DP_OP_425J2_127_3477_n2445), .Y(DP_OP_425J2_127_3477_n2412) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1650 ( .A1(DP_OP_422J2_124_3477_n2311), .A2(
        DP_OP_423J2_125_3477_n2444), .Y(DP_OP_425J2_127_3477_n2411) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1649 ( .A1(DP_OP_425J2_127_3477_n2442), .A2(
        DP_OP_424J2_126_3477_n2444), .Y(DP_OP_425J2_127_3477_n2410) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1648 ( .A1(DP_OP_425J2_127_3477_n2441), .A2(
        DP_OP_423J2_125_3477_n2444), .Y(DP_OP_425J2_127_3477_n2409) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1647 ( .A1(DP_OP_422J2_124_3477_n2308), .A2(
        DP_OP_422J2_124_3477_n2444), .Y(DP_OP_425J2_127_3477_n2408) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1646 ( .A1(DP_OP_425J2_127_3477_n2439), .A2(
        DP_OP_422J2_124_3477_n2444), .Y(DP_OP_425J2_127_3477_n2407) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1645 ( .A1(DP_OP_425J2_127_3477_n2438), .A2(
        DP_OP_424J2_126_3477_n2444), .Y(DP_OP_425J2_127_3477_n2406) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1644 ( .A1(DP_OP_422J2_124_3477_n2305), .A2(
        DP_OP_422J2_124_3477_n2444), .Y(DP_OP_425J2_127_3477_n2405) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1643 ( .A1(DP_OP_423J2_125_3477_n2612), 
        .A2(DP_OP_423J2_125_3477_n2444), .Y(DP_OP_425J2_127_3477_n2404) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1623 ( .A1(DP_OP_422J2_124_3477_n2260), .A2(
        DP_OP_425J2_127_3477_n2403), .Y(DP_OP_425J2_127_3477_n2384) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1615 ( .A1(DP_OP_422J2_124_3477_n2260), .A2(
        DP_OP_425J2_127_3477_n2402), .Y(DP_OP_425J2_127_3477_n2376) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1608 ( .A1(DP_OP_424J2_126_3477_n2569), 
        .A2(DP_OP_425J2_127_3477_n2401), .Y(DP_OP_425J2_127_3477_n2369) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1607 ( .A1(DP_OP_423J2_125_3477_n2656), .A2(
        DP_OP_425J2_127_3477_n2401), .Y(DP_OP_425J2_127_3477_n2368) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1606 ( .A1(DP_OP_423J2_125_3477_n2663), .A2(
        DP_OP_425J2_127_3477_n2400), .Y(DP_OP_425J2_127_3477_n2367) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1605 ( .A1(DP_OP_425J2_127_3477_n2398), .A2(
        DP_OP_425J2_127_3477_n2400), .Y(DP_OP_425J2_127_3477_n2366) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1604 ( .A1(DP_OP_425J2_127_3477_n2397), .A2(
        DP_OP_425J2_127_3477_n2400), .Y(DP_OP_425J2_127_3477_n2365) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1603 ( .A1(DP_OP_425J2_127_3477_n2396), .A2(
        DP_OP_425J2_127_3477_n2400), .Y(DP_OP_425J2_127_3477_n2364) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1602 ( .A1(DP_OP_423J2_125_3477_n2659), .A2(
        DP_OP_425J2_127_3477_n2400), .Y(DP_OP_425J2_127_3477_n2363) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1601 ( .A1(DP_OP_423J2_125_3477_n2658), .A2(
        DP_OP_425J2_127_3477_n2400), .Y(DP_OP_425J2_127_3477_n2362) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1600 ( .A1(DP_OP_422J2_124_3477_n2261), .A2(
        DP_OP_425J2_127_3477_n2400), .Y(DP_OP_425J2_127_3477_n2361) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1599 ( .A1(DP_OP_423J2_125_3477_n2656), 
        .A2(DP_OP_425J2_127_3477_n2400), .Y(DP_OP_425J2_127_3477_n2360) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1579 ( .A1(DP_OP_423J2_125_3477_n2700), .A2(
        DP_OP_425J2_127_3477_n2359), .Y(DP_OP_425J2_127_3477_n2340) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1571 ( .A1(DP_OP_423J2_125_3477_n2700), .A2(
        DP_OP_425J2_127_3477_n2358), .Y(DP_OP_425J2_127_3477_n2332) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1563 ( .A1(DP_OP_424J2_126_3477_n2612), .A2(
        DP_OP_425J2_127_3477_n2357), .Y(DP_OP_425J2_127_3477_n2324) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1562 ( .A1(DP_OP_425J2_127_3477_n2355), .A2(
        DP_OP_425J2_127_3477_n2356), .Y(DP_OP_425J2_127_3477_n2323) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1561 ( .A1(DP_OP_425J2_127_3477_n2354), .A2(
        DP_OP_425J2_127_3477_n2356), .Y(DP_OP_425J2_127_3477_n2322) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1560 ( .A1(DP_OP_425J2_127_3477_n2353), .A2(
        DP_OP_425J2_127_3477_n2356), .Y(DP_OP_425J2_127_3477_n2321) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1559 ( .A1(DP_OP_422J2_124_3477_n2220), .A2(
        DP_OP_425J2_127_3477_n2356), .Y(DP_OP_425J2_127_3477_n2320) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1558 ( .A1(DP_OP_425J2_127_3477_n2351), .A2(
        DP_OP_425J2_127_3477_n2356), .Y(DP_OP_425J2_127_3477_n2319) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1557 ( .A1(DP_OP_423J2_125_3477_n2702), .A2(
        DP_OP_425J2_127_3477_n2356), .Y(DP_OP_425J2_127_3477_n2318) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1556 ( .A1(DP_OP_424J2_126_3477_n2613), .A2(
        DP_OP_425J2_127_3477_n2356), .Y(DP_OP_425J2_127_3477_n2317) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1555 ( .A1(DP_OP_424J2_126_3477_n2612), 
        .A2(DP_OP_425J2_127_3477_n2356), .Y(DP_OP_425J2_127_3477_n2316) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1536 ( .A1(DP_OP_425J2_127_3477_n2305), 
        .A2(DP_OP_425J2_127_3477_n2315), .Y(DP_OP_425J2_127_3477_n2297) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1535 ( .A1(DP_OP_425J2_127_3477_n2304), .A2(
        DP_OP_425J2_127_3477_n2315), .Y(DP_OP_425J2_127_3477_n2296) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1527 ( .A1(DP_OP_425J2_127_3477_n2304), .A2(
        DP_OP_425J2_127_3477_n2314), .Y(DP_OP_425J2_127_3477_n2288) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1519 ( .A1(DP_OP_425J2_127_3477_n2304), .A2(
        DP_OP_425J2_127_3477_n2313), .Y(DP_OP_425J2_127_3477_n2280) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1518 ( .A1(DP_OP_424J2_126_3477_n2663), .A2(
        DP_OP_425J2_127_3477_n2312), .Y(DP_OP_425J2_127_3477_n2279) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1517 ( .A1(DP_OP_422J2_124_3477_n2178), .A2(
        DP_OP_425J2_127_3477_n2312), .Y(DP_OP_425J2_127_3477_n2278) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1516 ( .A1(DP_OP_422J2_124_3477_n2177), .A2(
        DP_OP_425J2_127_3477_n2312), .Y(DP_OP_425J2_127_3477_n2277) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1515 ( .A1(DP_OP_425J2_127_3477_n2308), .A2(
        DP_OP_425J2_127_3477_n2312), .Y(DP_OP_425J2_127_3477_n2276) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1514 ( .A1(DP_OP_425J2_127_3477_n2307), .A2(
        DP_OP_425J2_127_3477_n2312), .Y(DP_OP_425J2_127_3477_n2275) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1513 ( .A1(DP_OP_423J2_125_3477_n2746), .A2(
        DP_OP_425J2_127_3477_n2312), .Y(DP_OP_425J2_127_3477_n2274) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1512 ( .A1(DP_OP_425J2_127_3477_n2305), .A2(
        DP_OP_425J2_127_3477_n2312), .Y(DP_OP_425J2_127_3477_n2273) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1511 ( .A1(DP_OP_425J2_127_3477_n2304), 
        .A2(DP_OP_425J2_127_3477_n2312), .Y(DP_OP_425J2_127_3477_n2272) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1492 ( .A1(DP_OP_425J2_127_3477_n2261), 
        .A2(DP_OP_425J2_127_3477_n2271), .Y(DP_OP_425J2_127_3477_n2253) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1491 ( .A1(DP_OP_425J2_127_3477_n2260), .A2(
        DP_OP_425J2_127_3477_n2271), .Y(DP_OP_425J2_127_3477_n2252) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1483 ( .A1(DP_OP_425J2_127_3477_n2260), .A2(
        DP_OP_425J2_127_3477_n2270), .Y(DP_OP_425J2_127_3477_n2244) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1475 ( .A1(DP_OP_425J2_127_3477_n2260), .A2(
        DP_OP_425J2_127_3477_n2269), .Y(DP_OP_425J2_127_3477_n2236) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1474 ( .A1(DP_OP_423J2_125_3477_n2795), .A2(
        DP_OP_425J2_127_3477_n2268), .Y(DP_OP_425J2_127_3477_n2235) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1473 ( .A1(DP_OP_423J2_125_3477_n2794), .A2(
        DP_OP_425J2_127_3477_n2268), .Y(DP_OP_425J2_127_3477_n2234) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1472 ( .A1(DP_OP_423J2_125_3477_n2793), .A2(
        DP_OP_425J2_127_3477_n2268), .Y(DP_OP_425J2_127_3477_n2233) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1471 ( .A1(DP_OP_425J2_127_3477_n2264), .A2(
        DP_OP_425J2_127_3477_n2268), .Y(DP_OP_425J2_127_3477_n2232) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1470 ( .A1(DP_OP_423J2_125_3477_n2791), .A2(
        DP_OP_425J2_127_3477_n2268), .Y(DP_OP_425J2_127_3477_n2231) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1469 ( .A1(DP_OP_423J2_125_3477_n2790), .A2(
        DP_OP_425J2_127_3477_n2268), .Y(DP_OP_425J2_127_3477_n2230) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1468 ( .A1(DP_OP_425J2_127_3477_n2261), .A2(
        DP_OP_425J2_127_3477_n2268), .Y(DP_OP_425J2_127_3477_n2229) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1467 ( .A1(DP_OP_425J2_127_3477_n2260), 
        .A2(DP_OP_425J2_127_3477_n2268), .Y(DP_OP_425J2_127_3477_n2228) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1447 ( .A1(DP_OP_425J2_127_3477_n2216), .A2(
        DP_OP_425J2_127_3477_n2227), .Y(DP_OP_425J2_127_3477_n2208) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1440 ( .A1(DP_OP_425J2_127_3477_n2217), 
        .A2(DP_OP_425J2_127_3477_n2226), .Y(DP_OP_425J2_127_3477_n2201) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1439 ( .A1(DP_OP_425J2_127_3477_n2216), .A2(
        DP_OP_425J2_127_3477_n2226), .Y(DP_OP_425J2_127_3477_n2200) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1432 ( .A1(DP_OP_425J2_127_3477_n2217), 
        .A2(DP_OP_424J2_126_3477_n2225), .Y(DP_OP_425J2_127_3477_n2193) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1431 ( .A1(DP_OP_425J2_127_3477_n2216), .A2(
        DP_OP_424J2_126_3477_n2225), .Y(DP_OP_425J2_127_3477_n2192) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1430 ( .A1(DP_OP_424J2_126_3477_n2751), .A2(
        DP_OP_425J2_127_3477_n2224), .Y(DP_OP_425J2_127_3477_n2191) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1429 ( .A1(DP_OP_424J2_126_3477_n2750), .A2(
        DP_OP_425J2_127_3477_n2224), .Y(DP_OP_425J2_127_3477_n2190) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1428 ( .A1(DP_OP_423J2_125_3477_n2837), .A2(
        DP_OP_425J2_127_3477_n2224), .Y(DP_OP_425J2_127_3477_n2189) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1427 ( .A1(DP_OP_425J2_127_3477_n2220), .A2(
        DP_OP_425J2_127_3477_n2224), .Y(DP_OP_425J2_127_3477_n2188) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1426 ( .A1(DP_OP_425J2_127_3477_n2219), .A2(
        DP_OP_425J2_127_3477_n2224), .Y(DP_OP_425J2_127_3477_n2187) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1425 ( .A1(DP_OP_425J2_127_3477_n2218), .A2(
        DP_OP_425J2_127_3477_n2224), .Y(DP_OP_425J2_127_3477_n2186) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1424 ( .A1(DP_OP_425J2_127_3477_n2217), .A2(
        DP_OP_425J2_127_3477_n2224), .Y(DP_OP_425J2_127_3477_n2185) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1423 ( .A1(DP_OP_425J2_127_3477_n2216), 
        .A2(DP_OP_425J2_127_3477_n2224), .Y(DP_OP_425J2_127_3477_n2184) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1403 ( .A1(DP_OP_425J2_127_3477_n2172), .A2(
        DP_OP_422J2_124_3477_n2183), .Y(DP_OP_425J2_127_3477_n2164) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1395 ( .A1(DP_OP_425J2_127_3477_n2172), .A2(
        DP_OP_425J2_127_3477_n2182), .Y(DP_OP_425J2_127_3477_n2156) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1387 ( .A1(DP_OP_425J2_127_3477_n2172), .A2(
        DP_OP_425J2_127_3477_n2181), .Y(DP_OP_425J2_127_3477_n2148) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1386 ( .A1(DP_OP_422J2_124_3477_n2047), .A2(
        DP_OP_425J2_127_3477_n2180), .Y(DP_OP_425J2_127_3477_n2147) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1385 ( .A1(DP_OP_425J2_127_3477_n2178), .A2(
        DP_OP_425J2_127_3477_n2180), .Y(DP_OP_425J2_127_3477_n2146) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1384 ( .A1(DP_OP_422J2_124_3477_n2045), .A2(
        DP_OP_425J2_127_3477_n2180), .Y(DP_OP_425J2_127_3477_n2145) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1383 ( .A1(DP_OP_423J2_125_3477_n2880), .A2(
        DP_OP_425J2_127_3477_n2180), .Y(DP_OP_425J2_127_3477_n2144) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1382 ( .A1(DP_OP_425J2_127_3477_n2175), .A2(
        DP_OP_425J2_127_3477_n2180), .Y(DP_OP_425J2_127_3477_n2143) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1381 ( .A1(DP_OP_424J2_126_3477_n2790), .A2(
        DP_OP_425J2_127_3477_n2180), .Y(DP_OP_425J2_127_3477_n2142) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1380 ( .A1(DP_OP_424J2_126_3477_n2789), .A2(
        DP_OP_425J2_127_3477_n2180), .Y(DP_OP_425J2_127_3477_n2141) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1379 ( .A1(DP_OP_425J2_127_3477_n2172), 
        .A2(DP_OP_425J2_127_3477_n2180), .Y(DP_OP_425J2_127_3477_n2140) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1359 ( .A1(DP_OP_425J2_127_3477_n2128), .A2(
        DP_OP_425J2_127_3477_n2139), .Y(DP_OP_425J2_127_3477_n2120) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1351 ( .A1(DP_OP_425J2_127_3477_n2128), .A2(
        DP_OP_425J2_127_3477_n2138), .Y(DP_OP_425J2_127_3477_n2112) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1344 ( .A1(DP_OP_424J2_126_3477_n2833), 
        .A2(DP_OP_425J2_127_3477_n2137), .Y(DP_OP_425J2_127_3477_n2105) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1343 ( .A1(DP_OP_425J2_127_3477_n2128), .A2(
        DP_OP_425J2_127_3477_n2137), .Y(DP_OP_425J2_127_3477_n2104) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1342 ( .A1(DP_OP_425J2_127_3477_n2135), .A2(
        DP_OP_425J2_127_3477_n2136), .Y(DP_OP_425J2_127_3477_n2103) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1341 ( .A1(DP_OP_425J2_127_3477_n2134), .A2(
        DP_OP_425J2_127_3477_n2136), .Y(DP_OP_425J2_127_3477_n2102) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1340 ( .A1(DP_OP_425J2_127_3477_n2133), .A2(
        DP_OP_425J2_127_3477_n2136), .Y(DP_OP_425J2_127_3477_n2101) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1339 ( .A1(DP_OP_422J2_124_3477_n2000), .A2(
        DP_OP_425J2_127_3477_n2136), .Y(DP_OP_425J2_127_3477_n2100) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1338 ( .A1(DP_OP_424J2_126_3477_n2835), .A2(
        DP_OP_425J2_127_3477_n2136), .Y(DP_OP_425J2_127_3477_n2099) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1337 ( .A1(DP_OP_423J2_125_3477_n2922), .A2(
        DP_OP_425J2_127_3477_n2136), .Y(DP_OP_425J2_127_3477_n2098) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1336 ( .A1(DP_OP_424J2_126_3477_n2833), .A2(
        DP_OP_425J2_127_3477_n2136), .Y(DP_OP_425J2_127_3477_n2097) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1335 ( .A1(DP_OP_425J2_127_3477_n2128), 
        .A2(DP_OP_425J2_127_3477_n2136), .Y(DP_OP_425J2_127_3477_n2096) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1322 ( .A1(DP_OP_424J2_126_3477_n2883), 
        .A2(DP_OP_425J2_127_3477_n2095), .Y(DP_OP_425J2_127_3477_n2083) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1321 ( .A1(DP_OP_422J2_124_3477_n1958), 
        .A2(DP_OP_425J2_127_3477_n2095), .Y(DP_OP_425J2_127_3477_n2082) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1320 ( .A1(DP_OP_423J2_125_3477_n2969), 
        .A2(DP_OP_425J2_127_3477_n2095), .Y(DP_OP_425J2_127_3477_n2081) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1319 ( .A1(DP_OP_425J2_127_3477_n2088), 
        .A2(DP_OP_425J2_127_3477_n2095), .Y(DP_OP_425J2_127_3477_n2080) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1318 ( .A1(DP_OP_425J2_127_3477_n2087), 
        .A2(DP_OP_425J2_127_3477_n2095), .Y(DP_OP_425J2_127_3477_n2079) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1317 ( .A1(DP_OP_425J2_127_3477_n2086), 
        .A2(DP_OP_425J2_127_3477_n2095), .Y(DP_OP_425J2_127_3477_n2078) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1316 ( .A1(DP_OP_425J2_127_3477_n2085), 
        .A2(DP_OP_425J2_127_3477_n2095), .Y(DP_OP_425J2_127_3477_n2077) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1315 ( .A1(DP_OP_425J2_127_3477_n2084), .A2(
        DP_OP_425J2_127_3477_n2095), .Y(DP_OP_425J2_127_3477_n2076) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1314 ( .A1(DP_OP_424J2_126_3477_n2883), 
        .A2(DP_OP_425J2_127_3477_n2094), .Y(DP_OP_425J2_127_3477_n2075) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1313 ( .A1(DP_OP_422J2_124_3477_n1958), 
        .A2(DP_OP_425J2_127_3477_n2094), .Y(DP_OP_425J2_127_3477_n2074) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1312 ( .A1(DP_OP_423J2_125_3477_n2969), 
        .A2(DP_OP_425J2_127_3477_n2094), .Y(DP_OP_425J2_127_3477_n2073) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1311 ( .A1(DP_OP_425J2_127_3477_n2088), 
        .A2(DP_OP_425J2_127_3477_n2094), .Y(DP_OP_425J2_127_3477_n2072) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1310 ( .A1(DP_OP_425J2_127_3477_n2087), 
        .A2(DP_OP_425J2_127_3477_n2094), .Y(DP_OP_425J2_127_3477_n2071) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1309 ( .A1(DP_OP_425J2_127_3477_n2086), 
        .A2(DP_OP_425J2_127_3477_n2094), .Y(DP_OP_425J2_127_3477_n2070) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1308 ( .A1(DP_OP_425J2_127_3477_n2085), 
        .A2(DP_OP_425J2_127_3477_n2094), .Y(DP_OP_425J2_127_3477_n2069) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1307 ( .A1(DP_OP_425J2_127_3477_n2084), .A2(
        DP_OP_425J2_127_3477_n2094), .Y(DP_OP_425J2_127_3477_n2068) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1299 ( .A1(DP_OP_425J2_127_3477_n2084), .A2(
        DP_OP_425J2_127_3477_n2093), .Y(DP_OP_425J2_127_3477_n2060) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1298 ( .A1(DP_OP_423J2_125_3477_n2971), .A2(
        DP_OP_425J2_127_3477_n2092), .Y(DP_OP_425J2_127_3477_n2059) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1297 ( .A1(DP_OP_423J2_125_3477_n2970), .A2(
        DP_OP_425J2_127_3477_n2092), .Y(DP_OP_425J2_127_3477_n2058) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1296 ( .A1(DP_OP_423J2_125_3477_n2969), .A2(
        DP_OP_425J2_127_3477_n2092), .Y(DP_OP_425J2_127_3477_n2057) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1295 ( .A1(DP_OP_425J2_127_3477_n2088), .A2(
        DP_OP_425J2_127_3477_n2092), .Y(DP_OP_425J2_127_3477_n2056) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1294 ( .A1(DP_OP_425J2_127_3477_n2087), .A2(
        DP_OP_425J2_127_3477_n2092), .Y(DP_OP_425J2_127_3477_n2055) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1293 ( .A1(DP_OP_425J2_127_3477_n2086), .A2(
        DP_OP_425J2_127_3477_n2092), .Y(DP_OP_425J2_127_3477_n2054) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1292 ( .A1(DP_OP_425J2_127_3477_n2085), .A2(
        DP_OP_425J2_127_3477_n2092), .Y(DP_OP_425J2_127_3477_n2053) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1291 ( .A1(DP_OP_425J2_127_3477_n2084), 
        .A2(DP_OP_425J2_127_3477_n2092), .Y(DP_OP_425J2_127_3477_n2052) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1278 ( .A1(DP_OP_425J2_127_3477_n2047), 
        .A2(DP_OP_425J2_127_3477_n2051), .Y(DP_OP_425J2_127_3477_n2039) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1277 ( .A1(DP_OP_423J2_125_3477_n3012), 
        .A2(DP_OP_425J2_127_3477_n2051), .Y(DP_OP_425J2_127_3477_n2038) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1276 ( .A1(DP_OP_423J2_125_3477_n3011), 
        .A2(DP_OP_425J2_127_3477_n2051), .Y(DP_OP_425J2_127_3477_n2037) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1275 ( .A1(DP_OP_423J2_125_3477_n3010), 
        .A2(DP_OP_425J2_127_3477_n2051), .Y(DP_OP_425J2_127_3477_n2036) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1274 ( .A1(DP_OP_423J2_125_3477_n3009), 
        .A2(DP_OP_425J2_127_3477_n2051), .Y(DP_OP_425J2_127_3477_n2035) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1273 ( .A1(DP_OP_423J2_125_3477_n3008), 
        .A2(DP_OP_425J2_127_3477_n2051), .Y(DP_OP_425J2_127_3477_n2034) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1272 ( .A1(DP_OP_423J2_125_3477_n3007), 
        .A2(DP_OP_425J2_127_3477_n2051), .Y(DP_OP_425J2_127_3477_n2033) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1271 ( .A1(DP_OP_423J2_125_3477_n3006), .A2(
        DP_OP_425J2_127_3477_n2051), .Y(DP_OP_425J2_127_3477_n2032) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1263 ( .A1(DP_OP_423J2_125_3477_n3006), .A2(
        DP_OP_425J2_127_3477_n2050), .Y(DP_OP_425J2_127_3477_n2024) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1255 ( .A1(DP_OP_423J2_125_3477_n3006), .A2(
        DP_OP_425J2_127_3477_n2049), .Y(DP_OP_425J2_127_3477_n2016) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1254 ( .A1(DP_OP_425J2_127_3477_n2047), .A2(
        DP_OP_425J2_127_3477_n2048), .Y(DP_OP_425J2_127_3477_n2015) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1253 ( .A1(DP_OP_423J2_125_3477_n3012), .A2(
        DP_OP_425J2_127_3477_n2048), .Y(DP_OP_425J2_127_3477_n2014) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1252 ( .A1(DP_OP_423J2_125_3477_n3011), .A2(
        DP_OP_425J2_127_3477_n2048), .Y(DP_OP_425J2_127_3477_n2013) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1251 ( .A1(DP_OP_423J2_125_3477_n3010), .A2(
        DP_OP_425J2_127_3477_n2048), .Y(DP_OP_425J2_127_3477_n2012) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1250 ( .A1(DP_OP_423J2_125_3477_n3009), .A2(
        DP_OP_425J2_127_3477_n2048), .Y(DP_OP_425J2_127_3477_n2011) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1249 ( .A1(DP_OP_423J2_125_3477_n3008), .A2(
        DP_OP_425J2_127_3477_n2048), .Y(DP_OP_425J2_127_3477_n2010) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1248 ( .A1(DP_OP_423J2_125_3477_n3007), .A2(
        DP_OP_425J2_127_3477_n2048), .Y(DP_OP_425J2_127_3477_n2009) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1247 ( .A1(DP_OP_423J2_125_3477_n3006), 
        .A2(DP_OP_425J2_127_3477_n2048), .Y(DP_OP_425J2_127_3477_n2008) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1227 ( .A1(DP_OP_424J2_126_3477_n2964), .A2(
        DP_OP_425J2_127_3477_n2007), .Y(DP_OP_425J2_127_3477_n1988) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1219 ( .A1(DP_OP_424J2_126_3477_n2964), .A2(
        DP_OP_425J2_127_3477_n2006), .Y(DP_OP_425J2_127_3477_n1980) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1212 ( .A1(DP_OP_425J2_127_3477_n1997), 
        .A2(DP_OP_425J2_127_3477_n2005), .Y(DP_OP_425J2_127_3477_n1973) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1211 ( .A1(DP_OP_424J2_126_3477_n2964), .A2(
        DP_OP_425J2_127_3477_n2005), .Y(DP_OP_425J2_127_3477_n1972) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1210 ( .A1(DP_OP_425J2_127_3477_n2003), .A2(
        DP_OP_425J2_127_3477_n2004), .Y(DP_OP_425J2_127_3477_n1971) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1209 ( .A1(DP_OP_424J2_126_3477_n2970), .A2(
        DP_OP_425J2_127_3477_n2004), .Y(DP_OP_425J2_127_3477_n1970) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1208 ( .A1(DP_OP_424J2_126_3477_n2969), .A2(
        DP_OP_425J2_127_3477_n2004), .Y(DP_OP_425J2_127_3477_n1969) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1207 ( .A1(DP_OP_425J2_127_3477_n2000), .A2(
        DP_OP_425J2_127_3477_n2004), .Y(DP_OP_425J2_127_3477_n1968) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1206 ( .A1(DP_OP_424J2_126_3477_n2967), .A2(
        DP_OP_425J2_127_3477_n2004), .Y(DP_OP_425J2_127_3477_n1967) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1205 ( .A1(DP_OP_425J2_127_3477_n1998), .A2(
        DP_OP_425J2_127_3477_n2004), .Y(DP_OP_425J2_127_3477_n1966) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1204 ( .A1(DP_OP_425J2_127_3477_n1997), .A2(
        DP_OP_425J2_127_3477_n2004), .Y(DP_OP_425J2_127_3477_n1965) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1203 ( .A1(DP_OP_424J2_126_3477_n2964), 
        .A2(DP_OP_425J2_127_3477_n2004), .Y(DP_OP_425J2_127_3477_n1964) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1184 ( .A1(DP_OP_424J2_126_3477_n3007), 
        .A2(DP_OP_425J2_127_3477_n1963), .Y(DP_OP_425J2_127_3477_n1945) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1183 ( .A1(DP_OP_424J2_126_3477_n3006), .A2(
        DP_OP_425J2_127_3477_n1963), .Y(DP_OP_425J2_127_3477_n1944) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1175 ( .A1(DP_OP_424J2_126_3477_n3006), .A2(
        DP_OP_423J2_125_3477_n1962), .Y(DP_OP_425J2_127_3477_n1936) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1167 ( .A1(DP_OP_424J2_126_3477_n3006), .A2(
        DP_OP_425J2_127_3477_n1961), .Y(DP_OP_425J2_127_3477_n1928) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1166 ( .A1(DP_OP_424J2_126_3477_n3013), .A2(
        DP_OP_425J2_127_3477_n1960), .Y(DP_OP_425J2_127_3477_n1927) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1165 ( .A1(DP_OP_424J2_126_3477_n3012), .A2(
        DP_OP_425J2_127_3477_n1960), .Y(DP_OP_425J2_127_3477_n1926) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1164 ( .A1(DP_OP_424J2_126_3477_n3011), .A2(
        DP_OP_425J2_127_3477_n1960), .Y(DP_OP_425J2_127_3477_n1925) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1163 ( .A1(DP_OP_424J2_126_3477_n3010), .A2(
        DP_OP_425J2_127_3477_n1960), .Y(DP_OP_425J2_127_3477_n1924) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1162 ( .A1(DP_OP_424J2_126_3477_n3009), .A2(
        DP_OP_425J2_127_3477_n1960), .Y(DP_OP_425J2_127_3477_n1923) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1161 ( .A1(DP_OP_424J2_126_3477_n3008), .A2(
        DP_OP_425J2_127_3477_n1960), .Y(DP_OP_425J2_127_3477_n1922) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1160 ( .A1(DP_OP_424J2_126_3477_n3007), .A2(
        DP_OP_425J2_127_3477_n1960), .Y(DP_OP_425J2_127_3477_n1921) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1159 ( .A1(DP_OP_424J2_126_3477_n3006), 
        .A2(DP_OP_425J2_127_3477_n1960), .Y(DP_OP_425J2_127_3477_n1920) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1112 ( .A1(n368), .A2(n389), .Y(
        DP_OP_425J2_127_3477_n1874) );
  HADDX1_HVT DP_OP_425J2_127_3477_U1093 ( .A0(DP_OP_425J2_127_3477_n1886), 
        .B0(DP_OP_425J2_127_3477_n1995), .C1(DP_OP_425J2_127_3477_n1870), .SO(
        DP_OP_425J2_127_3477_n1871) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1092 ( .A(DP_OP_425J2_127_3477_n2039), .B(
        DP_OP_425J2_127_3477_n1951), .CI(DP_OP_425J2_127_3477_n2083), .CO(
        DP_OP_425J2_127_3477_n1868), .S(DP_OP_425J2_127_3477_n1869) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1091 ( .A(DP_OP_425J2_127_3477_n2171), .B(
        DP_OP_425J2_127_3477_n2127), .CI(DP_OP_425J2_127_3477_n2215), .CO(
        DP_OP_425J2_127_3477_n1866), .S(DP_OP_425J2_127_3477_n1867) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1090 ( .A(DP_OP_425J2_127_3477_n2303), .B(
        DP_OP_425J2_127_3477_n2259), .CI(DP_OP_425J2_127_3477_n2347), .CO(
        DP_OP_425J2_127_3477_n1864), .S(DP_OP_425J2_127_3477_n1865) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1089 ( .A(DP_OP_425J2_127_3477_n2435), .B(
        DP_OP_425J2_127_3477_n2391), .CI(DP_OP_425J2_127_3477_n2479), .CO(
        DP_OP_425J2_127_3477_n1862), .S(DP_OP_425J2_127_3477_n1863) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1088 ( .A(DP_OP_425J2_127_3477_n2567), .B(
        DP_OP_425J2_127_3477_n2523), .CI(DP_OP_425J2_127_3477_n2611), .CO(
        DP_OP_425J2_127_3477_n1860), .S(DP_OP_425J2_127_3477_n1861) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1087 ( .A(DP_OP_425J2_127_3477_n2699), .B(
        DP_OP_425J2_127_3477_n2655), .CI(DP_OP_425J2_127_3477_n2743), .CO(
        DP_OP_425J2_127_3477_n1858), .S(DP_OP_425J2_127_3477_n1859) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1086 ( .A(DP_OP_425J2_127_3477_n3005), .B(
        DP_OP_425J2_127_3477_n2787), .CI(DP_OP_425J2_127_3477_n2831), .CO(
        DP_OP_425J2_127_3477_n1856), .S(DP_OP_425J2_127_3477_n1857) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1085 ( .A(DP_OP_425J2_127_3477_n2963), .B(
        DP_OP_425J2_127_3477_n2875), .CI(DP_OP_425J2_127_3477_n2919), .CO(
        DP_OP_425J2_127_3477_n1854), .S(DP_OP_425J2_127_3477_n1855) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1084 ( .A(DP_OP_425J2_127_3477_n1871), .B(
        DP_OP_425J2_127_3477_n1857), .CI(DP_OP_425J2_127_3477_n1859), .CO(
        DP_OP_425J2_127_3477_n1852), .S(DP_OP_425J2_127_3477_n1853) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1083 ( .A(DP_OP_425J2_127_3477_n1861), .B(
        DP_OP_425J2_127_3477_n1855), .CI(DP_OP_425J2_127_3477_n1863), .CO(
        DP_OP_425J2_127_3477_n1850), .S(DP_OP_425J2_127_3477_n1851) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1082 ( .A(DP_OP_425J2_127_3477_n1869), .B(
        DP_OP_425J2_127_3477_n1865), .CI(DP_OP_425J2_127_3477_n1867), .CO(
        DP_OP_425J2_127_3477_n1848), .S(DP_OP_425J2_127_3477_n1849) );
  HADDX1_HVT DP_OP_425J2_127_3477_U1081 ( .A0(DP_OP_425J2_127_3477_n1885), 
        .B0(DP_OP_425J2_127_3477_n1950), .C1(DP_OP_425J2_127_3477_n1846), .SO(
        DP_OP_425J2_127_3477_n1847) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1080 ( .A(DP_OP_425J2_127_3477_n1987), .B(
        DP_OP_425J2_127_3477_n1943), .CI(DP_OP_425J2_127_3477_n1994), .CO(
        DP_OP_425J2_127_3477_n1844), .S(DP_OP_425J2_127_3477_n1845) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1079 ( .A(DP_OP_425J2_127_3477_n2038), .B(
        DP_OP_425J2_127_3477_n2031), .CI(DP_OP_425J2_127_3477_n2075), .CO(
        DP_OP_425J2_127_3477_n1842), .S(DP_OP_425J2_127_3477_n1843) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1078 ( .A(DP_OP_425J2_127_3477_n2119), .B(
        DP_OP_425J2_127_3477_n2082), .CI(DP_OP_425J2_127_3477_n2126), .CO(
        DP_OP_425J2_127_3477_n1840), .S(DP_OP_425J2_127_3477_n1841) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1077 ( .A(DP_OP_425J2_127_3477_n2170), .B(
        DP_OP_425J2_127_3477_n2163), .CI(DP_OP_425J2_127_3477_n2207), .CO(
        DP_OP_425J2_127_3477_n1838), .S(DP_OP_425J2_127_3477_n1839) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1076 ( .A(DP_OP_425J2_127_3477_n2251), .B(
        DP_OP_425J2_127_3477_n2214), .CI(DP_OP_425J2_127_3477_n2258), .CO(
        DP_OP_425J2_127_3477_n1836), .S(DP_OP_425J2_127_3477_n1837) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1075 ( .A(DP_OP_425J2_127_3477_n2302), .B(
        DP_OP_425J2_127_3477_n2295), .CI(DP_OP_425J2_127_3477_n2339), .CO(
        DP_OP_425J2_127_3477_n1834), .S(DP_OP_425J2_127_3477_n1835) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1074 ( .A(DP_OP_425J2_127_3477_n2383), .B(
        DP_OP_425J2_127_3477_n2346), .CI(DP_OP_425J2_127_3477_n2390), .CO(
        DP_OP_425J2_127_3477_n1832), .S(DP_OP_425J2_127_3477_n1833) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1073 ( .A(DP_OP_425J2_127_3477_n2434), .B(
        DP_OP_425J2_127_3477_n2427), .CI(DP_OP_425J2_127_3477_n2471), .CO(
        DP_OP_425J2_127_3477_n1830), .S(DP_OP_425J2_127_3477_n1831) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1072 ( .A(DP_OP_425J2_127_3477_n2515), .B(
        DP_OP_425J2_127_3477_n2478), .CI(DP_OP_425J2_127_3477_n2522), .CO(
        DP_OP_425J2_127_3477_n1828), .S(DP_OP_425J2_127_3477_n1829) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1071 ( .A(DP_OP_425J2_127_3477_n3004), .B(
        DP_OP_425J2_127_3477_n2559), .CI(DP_OP_425J2_127_3477_n2997), .CO(
        DP_OP_425J2_127_3477_n1826), .S(DP_OP_425J2_127_3477_n1827) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1070 ( .A(DP_OP_425J2_127_3477_n2742), .B(
        DP_OP_425J2_127_3477_n2566), .CI(DP_OP_425J2_127_3477_n2603), .CO(
        DP_OP_425J2_127_3477_n1824), .S(DP_OP_425J2_127_3477_n1825) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1069 ( .A(DP_OP_425J2_127_3477_n2779), .B(
        DP_OP_425J2_127_3477_n2962), .CI(DP_OP_425J2_127_3477_n2955), .CO(
        DP_OP_425J2_127_3477_n1822), .S(DP_OP_425J2_127_3477_n1823) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1068 ( .A(DP_OP_425J2_127_3477_n2698), .B(
        DP_OP_425J2_127_3477_n2918), .CI(DP_OP_425J2_127_3477_n2911), .CO(
        DP_OP_425J2_127_3477_n1820), .S(DP_OP_425J2_127_3477_n1821) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1067 ( .A(DP_OP_425J2_127_3477_n2691), .B(
        DP_OP_425J2_127_3477_n2874), .CI(DP_OP_425J2_127_3477_n2610), .CO(
        DP_OP_425J2_127_3477_n1818), .S(DP_OP_425J2_127_3477_n1819) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1066 ( .A(DP_OP_425J2_127_3477_n2867), .B(
        DP_OP_425J2_127_3477_n2647), .CI(DP_OP_425J2_127_3477_n2654), .CO(
        DP_OP_425J2_127_3477_n1816), .S(DP_OP_425J2_127_3477_n1817) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1065 ( .A(DP_OP_425J2_127_3477_n2823), .B(
        DP_OP_425J2_127_3477_n2735), .CI(DP_OP_425J2_127_3477_n2786), .CO(
        DP_OP_425J2_127_3477_n1814), .S(DP_OP_425J2_127_3477_n1815) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1064 ( .A(DP_OP_425J2_127_3477_n2830), .B(
        DP_OP_425J2_127_3477_n1870), .CI(DP_OP_425J2_127_3477_n1847), .CO(
        DP_OP_425J2_127_3477_n1812), .S(DP_OP_425J2_127_3477_n1813) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1063 ( .A(DP_OP_425J2_127_3477_n1854), .B(
        DP_OP_425J2_127_3477_n1868), .CI(DP_OP_425J2_127_3477_n1866), .CO(
        DP_OP_425J2_127_3477_n1810), .S(DP_OP_425J2_127_3477_n1811) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1062 ( .A(DP_OP_425J2_127_3477_n1860), .B(
        DP_OP_425J2_127_3477_n1856), .CI(DP_OP_425J2_127_3477_n1864), .CO(
        DP_OP_425J2_127_3477_n1808), .S(DP_OP_425J2_127_3477_n1809) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1061 ( .A(DP_OP_425J2_127_3477_n1862), .B(
        DP_OP_425J2_127_3477_n1858), .CI(DP_OP_425J2_127_3477_n1815), .CO(
        DP_OP_425J2_127_3477_n1806), .S(DP_OP_425J2_127_3477_n1807) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1060 ( .A(DP_OP_425J2_127_3477_n1837), .B(
        DP_OP_425J2_127_3477_n1823), .CI(DP_OP_425J2_127_3477_n1821), .CO(
        DP_OP_425J2_127_3477_n1804), .S(DP_OP_425J2_127_3477_n1805) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1059 ( .A(DP_OP_425J2_127_3477_n1841), .B(
        DP_OP_425J2_127_3477_n1825), .CI(DP_OP_425J2_127_3477_n1829), .CO(
        DP_OP_425J2_127_3477_n1802), .S(DP_OP_425J2_127_3477_n1803) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1058 ( .A(DP_OP_425J2_127_3477_n1843), .B(
        DP_OP_425J2_127_3477_n1831), .CI(DP_OP_425J2_127_3477_n1827), .CO(
        DP_OP_425J2_127_3477_n1800), .S(DP_OP_425J2_127_3477_n1801) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1057 ( .A(DP_OP_425J2_127_3477_n1845), .B(
        DP_OP_425J2_127_3477_n1835), .CI(DP_OP_425J2_127_3477_n1819), .CO(
        DP_OP_425J2_127_3477_n1798), .S(DP_OP_425J2_127_3477_n1799) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1056 ( .A(DP_OP_425J2_127_3477_n1839), .B(
        DP_OP_425J2_127_3477_n1833), .CI(DP_OP_425J2_127_3477_n1817), .CO(
        DP_OP_425J2_127_3477_n1796), .S(DP_OP_425J2_127_3477_n1797) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1055 ( .A(DP_OP_425J2_127_3477_n1813), .B(
        DP_OP_425J2_127_3477_n1852), .CI(DP_OP_425J2_127_3477_n1850), .CO(
        DP_OP_425J2_127_3477_n1794), .S(DP_OP_425J2_127_3477_n1795) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1054 ( .A(DP_OP_425J2_127_3477_n1848), .B(
        DP_OP_425J2_127_3477_n1809), .CI(DP_OP_425J2_127_3477_n1811), .CO(
        DP_OP_425J2_127_3477_n1792), .S(DP_OP_425J2_127_3477_n1793) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1053 ( .A(DP_OP_425J2_127_3477_n1807), .B(
        DP_OP_425J2_127_3477_n1799), .CI(DP_OP_425J2_127_3477_n1801), .CO(
        DP_OP_425J2_127_3477_n1790), .S(DP_OP_425J2_127_3477_n1791) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1052 ( .A(DP_OP_425J2_127_3477_n1805), .B(
        DP_OP_425J2_127_3477_n1797), .CI(DP_OP_425J2_127_3477_n1803), .CO(
        DP_OP_425J2_127_3477_n1788), .S(DP_OP_425J2_127_3477_n1789) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1051 ( .A(DP_OP_425J2_127_3477_n1795), .B(
        DP_OP_425J2_127_3477_n1793), .CI(DP_OP_425J2_127_3477_n1791), .CO(
        DP_OP_425J2_127_3477_n1786), .S(DP_OP_425J2_127_3477_n1787) );
  HADDX1_HVT DP_OP_425J2_127_3477_U1050 ( .A0(DP_OP_425J2_127_3477_n1884), 
        .B0(DP_OP_425J2_127_3477_n1949), .C1(DP_OP_425J2_127_3477_n1784), .SO(
        DP_OP_425J2_127_3477_n1785) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1049 ( .A(DP_OP_425J2_127_3477_n1979), .B(
        DP_OP_425J2_127_3477_n1942), .CI(DP_OP_425J2_127_3477_n1935), .CO(
        DP_OP_425J2_127_3477_n1782), .S(DP_OP_425J2_127_3477_n1783) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1048 ( .A(DP_OP_425J2_127_3477_n1993), .B(
        DP_OP_425J2_127_3477_n1986), .CI(DP_OP_425J2_127_3477_n2023), .CO(
        DP_OP_425J2_127_3477_n1780), .S(DP_OP_425J2_127_3477_n1781) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1047 ( .A(DP_OP_425J2_127_3477_n2037), .B(
        DP_OP_425J2_127_3477_n2030), .CI(DP_OP_425J2_127_3477_n2067), .CO(
        DP_OP_425J2_127_3477_n1778), .S(DP_OP_425J2_127_3477_n1779) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1046 ( .A(DP_OP_425J2_127_3477_n2081), .B(
        DP_OP_425J2_127_3477_n2074), .CI(DP_OP_425J2_127_3477_n2111), .CO(
        DP_OP_425J2_127_3477_n1776), .S(DP_OP_425J2_127_3477_n1777) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1045 ( .A(DP_OP_425J2_127_3477_n2125), .B(
        DP_OP_425J2_127_3477_n2118), .CI(DP_OP_425J2_127_3477_n2155), .CO(
        DP_OP_425J2_127_3477_n1774), .S(DP_OP_425J2_127_3477_n1775) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1044 ( .A(DP_OP_425J2_127_3477_n2169), .B(
        DP_OP_425J2_127_3477_n2162), .CI(DP_OP_425J2_127_3477_n2199), .CO(
        DP_OP_425J2_127_3477_n1772), .S(DP_OP_425J2_127_3477_n1773) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1043 ( .A(DP_OP_425J2_127_3477_n2213), .B(
        DP_OP_425J2_127_3477_n2206), .CI(DP_OP_425J2_127_3477_n2243), .CO(
        DP_OP_425J2_127_3477_n1770), .S(DP_OP_425J2_127_3477_n1771) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1042 ( .A(DP_OP_425J2_127_3477_n2257), .B(
        DP_OP_425J2_127_3477_n2250), .CI(DP_OP_425J2_127_3477_n2287), .CO(
        DP_OP_425J2_127_3477_n1768), .S(DP_OP_425J2_127_3477_n1769) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1041 ( .A(DP_OP_425J2_127_3477_n2301), .B(
        DP_OP_425J2_127_3477_n2294), .CI(DP_OP_425J2_127_3477_n2331), .CO(
        DP_OP_425J2_127_3477_n1766), .S(DP_OP_425J2_127_3477_n1767) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1040 ( .A(DP_OP_425J2_127_3477_n2345), .B(
        DP_OP_425J2_127_3477_n2338), .CI(DP_OP_425J2_127_3477_n2375), .CO(
        DP_OP_425J2_127_3477_n1764), .S(DP_OP_425J2_127_3477_n1765) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1039 ( .A(DP_OP_425J2_127_3477_n2389), .B(
        DP_OP_425J2_127_3477_n2382), .CI(DP_OP_425J2_127_3477_n2419), .CO(
        DP_OP_425J2_127_3477_n1762), .S(DP_OP_425J2_127_3477_n1763) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1038 ( .A(DP_OP_425J2_127_3477_n2690), .B(
        DP_OP_425J2_127_3477_n3003), .CI(DP_OP_425J2_127_3477_n2996), .CO(
        DP_OP_425J2_127_3477_n1760), .S(DP_OP_425J2_127_3477_n1761) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1037 ( .A(DP_OP_425J2_127_3477_n2653), .B(
        DP_OP_425J2_127_3477_n2426), .CI(DP_OP_425J2_127_3477_n2989), .CO(
        DP_OP_425J2_127_3477_n1758), .S(DP_OP_425J2_127_3477_n1759) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1036 ( .A(DP_OP_425J2_127_3477_n2646), .B(
        DP_OP_425J2_127_3477_n2961), .CI(DP_OP_425J2_127_3477_n2433), .CO(
        DP_OP_425J2_127_3477_n1756), .S(DP_OP_425J2_127_3477_n1757) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1035 ( .A(DP_OP_425J2_127_3477_n2683), .B(
        DP_OP_425J2_127_3477_n2463), .CI(DP_OP_425J2_127_3477_n2470), .CO(
        DP_OP_425J2_127_3477_n1754), .S(DP_OP_425J2_127_3477_n1755) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1034 ( .A(DP_OP_425J2_127_3477_n2697), .B(
        DP_OP_425J2_127_3477_n2477), .CI(DP_OP_425J2_127_3477_n2954), .CO(
        DP_OP_425J2_127_3477_n1752), .S(DP_OP_425J2_127_3477_n1753) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1033 ( .A(DP_OP_425J2_127_3477_n2727), .B(
        DP_OP_425J2_127_3477_n2507), .CI(DP_OP_425J2_127_3477_n2947), .CO(
        DP_OP_425J2_127_3477_n1750), .S(DP_OP_425J2_127_3477_n1751) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1032 ( .A(DP_OP_425J2_127_3477_n2639), .B(
        DP_OP_425J2_127_3477_n2514), .CI(DP_OP_425J2_127_3477_n2917), .CO(
        DP_OP_425J2_127_3477_n1748), .S(DP_OP_425J2_127_3477_n1749) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1031 ( .A(DP_OP_425J2_127_3477_n2609), .B(
        DP_OP_425J2_127_3477_n2521), .CI(DP_OP_425J2_127_3477_n2910), .CO(
        DP_OP_425J2_127_3477_n1746), .S(DP_OP_425J2_127_3477_n1747) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1030 ( .A(DP_OP_425J2_127_3477_n2903), .B(
        DP_OP_425J2_127_3477_n2551), .CI(DP_OP_425J2_127_3477_n2558), .CO(
        DP_OP_425J2_127_3477_n1744), .S(DP_OP_425J2_127_3477_n1745) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1029 ( .A(DP_OP_425J2_127_3477_n2873), .B(
        DP_OP_425J2_127_3477_n2565), .CI(DP_OP_425J2_127_3477_n2595), .CO(
        DP_OP_425J2_127_3477_n1742), .S(DP_OP_425J2_127_3477_n1743) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1028 ( .A(DP_OP_425J2_127_3477_n2866), .B(
        DP_OP_425J2_127_3477_n2602), .CI(DP_OP_425J2_127_3477_n2734), .CO(
        DP_OP_425J2_127_3477_n1740), .S(DP_OP_425J2_127_3477_n1741) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1027 ( .A(DP_OP_425J2_127_3477_n2859), .B(
        DP_OP_425J2_127_3477_n2741), .CI(DP_OP_425J2_127_3477_n2771), .CO(
        DP_OP_425J2_127_3477_n1738), .S(DP_OP_425J2_127_3477_n1739) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1026 ( .A(DP_OP_425J2_127_3477_n2829), .B(
        DP_OP_425J2_127_3477_n2778), .CI(DP_OP_425J2_127_3477_n2785), .CO(
        DP_OP_425J2_127_3477_n1736), .S(DP_OP_425J2_127_3477_n1737) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1025 ( .A(DP_OP_425J2_127_3477_n2822), .B(
        DP_OP_425J2_127_3477_n2815), .CI(DP_OP_425J2_127_3477_n1846), .CO(
        DP_OP_425J2_127_3477_n1734), .S(DP_OP_425J2_127_3477_n1735) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1024 ( .A(DP_OP_425J2_127_3477_n1785), .B(
        DP_OP_425J2_127_3477_n1814), .CI(DP_OP_425J2_127_3477_n1816), .CO(
        DP_OP_425J2_127_3477_n1732), .S(DP_OP_425J2_127_3477_n1733) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1023 ( .A(DP_OP_425J2_127_3477_n1832), .B(
        DP_OP_425J2_127_3477_n1844), .CI(DP_OP_425J2_127_3477_n1818), .CO(
        DP_OP_425J2_127_3477_n1730), .S(DP_OP_425J2_127_3477_n1731) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1022 ( .A(DP_OP_425J2_127_3477_n1830), .B(
        DP_OP_425J2_127_3477_n1842), .CI(DP_OP_425J2_127_3477_n1820), .CO(
        DP_OP_425J2_127_3477_n1728), .S(DP_OP_425J2_127_3477_n1729) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1021 ( .A(DP_OP_425J2_127_3477_n1826), .B(
        DP_OP_425J2_127_3477_n1840), .CI(DP_OP_425J2_127_3477_n1822), .CO(
        DP_OP_425J2_127_3477_n1726), .S(DP_OP_425J2_127_3477_n1727) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1020 ( .A(DP_OP_425J2_127_3477_n1838), .B(
        DP_OP_425J2_127_3477_n1836), .CI(DP_OP_425J2_127_3477_n1834), .CO(
        DP_OP_425J2_127_3477_n1724), .S(DP_OP_425J2_127_3477_n1725) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1019 ( .A(DP_OP_425J2_127_3477_n1828), .B(
        DP_OP_425J2_127_3477_n1824), .CI(DP_OP_425J2_127_3477_n1757), .CO(
        DP_OP_425J2_127_3477_n1722), .S(DP_OP_425J2_127_3477_n1723) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1018 ( .A(DP_OP_425J2_127_3477_n1751), .B(
        DP_OP_425J2_127_3477_n1765), .CI(DP_OP_425J2_127_3477_n1769), .CO(
        DP_OP_425J2_127_3477_n1720), .S(DP_OP_425J2_127_3477_n1721) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1017 ( .A(DP_OP_425J2_127_3477_n1747), .B(
        DP_OP_425J2_127_3477_n1775), .CI(DP_OP_425J2_127_3477_n1777), .CO(
        DP_OP_425J2_127_3477_n1718), .S(DP_OP_425J2_127_3477_n1719) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1016 ( .A(DP_OP_425J2_127_3477_n1745), .B(
        DP_OP_425J2_127_3477_n1767), .CI(DP_OP_425J2_127_3477_n1781), .CO(
        DP_OP_425J2_127_3477_n1716), .S(DP_OP_425J2_127_3477_n1717) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1015 ( .A(DP_OP_425J2_127_3477_n1743), .B(
        DP_OP_425J2_127_3477_n1761), .CI(DP_OP_425J2_127_3477_n1779), .CO(
        DP_OP_425J2_127_3477_n1714), .S(DP_OP_425J2_127_3477_n1715) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1014 ( .A(DP_OP_425J2_127_3477_n1741), .B(
        DP_OP_425J2_127_3477_n1771), .CI(DP_OP_425J2_127_3477_n1759), .CO(
        DP_OP_425J2_127_3477_n1712), .S(DP_OP_425J2_127_3477_n1713) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1013 ( .A(DP_OP_425J2_127_3477_n1739), .B(
        DP_OP_425J2_127_3477_n1773), .CI(DP_OP_425J2_127_3477_n1783), .CO(
        DP_OP_425J2_127_3477_n1710), .S(DP_OP_425J2_127_3477_n1711) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1012 ( .A(DP_OP_425J2_127_3477_n1737), .B(
        DP_OP_425J2_127_3477_n1763), .CI(DP_OP_425J2_127_3477_n1749), .CO(
        DP_OP_425J2_127_3477_n1708), .S(DP_OP_425J2_127_3477_n1709) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1011 ( .A(DP_OP_425J2_127_3477_n1755), .B(
        DP_OP_425J2_127_3477_n1753), .CI(DP_OP_425J2_127_3477_n1812), .CO(
        DP_OP_425J2_127_3477_n1706), .S(DP_OP_425J2_127_3477_n1707) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1010 ( .A(DP_OP_425J2_127_3477_n1735), .B(
        DP_OP_425J2_127_3477_n1810), .CI(DP_OP_425J2_127_3477_n1808), .CO(
        DP_OP_425J2_127_3477_n1704), .S(DP_OP_425J2_127_3477_n1705) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1009 ( .A(DP_OP_425J2_127_3477_n1806), .B(
        DP_OP_425J2_127_3477_n1733), .CI(DP_OP_425J2_127_3477_n1800), .CO(
        DP_OP_425J2_127_3477_n1702), .S(DP_OP_425J2_127_3477_n1703) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1008 ( .A(DP_OP_425J2_127_3477_n1804), .B(
        DP_OP_425J2_127_3477_n1725), .CI(DP_OP_425J2_127_3477_n1731), .CO(
        DP_OP_425J2_127_3477_n1700), .S(DP_OP_425J2_127_3477_n1701) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1007 ( .A(DP_OP_425J2_127_3477_n1802), .B(
        DP_OP_425J2_127_3477_n1729), .CI(DP_OP_425J2_127_3477_n1727), .CO(
        DP_OP_425J2_127_3477_n1698), .S(DP_OP_425J2_127_3477_n1699) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1006 ( .A(DP_OP_425J2_127_3477_n1798), .B(
        DP_OP_425J2_127_3477_n1796), .CI(DP_OP_425J2_127_3477_n1723), .CO(
        DP_OP_425J2_127_3477_n1696), .S(DP_OP_425J2_127_3477_n1697) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1005 ( .A(DP_OP_425J2_127_3477_n1721), .B(
        DP_OP_425J2_127_3477_n1709), .CI(DP_OP_425J2_127_3477_n1707), .CO(
        DP_OP_425J2_127_3477_n1694), .S(DP_OP_425J2_127_3477_n1695) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1004 ( .A(DP_OP_425J2_127_3477_n1711), .B(
        DP_OP_425J2_127_3477_n1719), .CI(DP_OP_425J2_127_3477_n1717), .CO(
        DP_OP_425J2_127_3477_n1692), .S(DP_OP_425J2_127_3477_n1693) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1003 ( .A(DP_OP_425J2_127_3477_n1713), .B(
        DP_OP_425J2_127_3477_n1715), .CI(DP_OP_425J2_127_3477_n1794), .CO(
        DP_OP_425J2_127_3477_n1690), .S(DP_OP_425J2_127_3477_n1691) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1002 ( .A(DP_OP_425J2_127_3477_n1705), .B(
        DP_OP_425J2_127_3477_n1792), .CI(DP_OP_425J2_127_3477_n1703), .CO(
        DP_OP_425J2_127_3477_n1688), .S(DP_OP_425J2_127_3477_n1689) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1001 ( .A(DP_OP_425J2_127_3477_n1790), .B(
        DP_OP_425J2_127_3477_n1788), .CI(DP_OP_425J2_127_3477_n1699), .CO(
        DP_OP_425J2_127_3477_n1686), .S(DP_OP_425J2_127_3477_n1687) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1000 ( .A(DP_OP_425J2_127_3477_n1701), .B(
        DP_OP_425J2_127_3477_n1697), .CI(DP_OP_425J2_127_3477_n1695), .CO(
        DP_OP_425J2_127_3477_n1684), .S(DP_OP_425J2_127_3477_n1685) );
  FADDX1_HVT DP_OP_425J2_127_3477_U999 ( .A(DP_OP_425J2_127_3477_n1693), .B(
        DP_OP_425J2_127_3477_n1691), .CI(DP_OP_425J2_127_3477_n1689), .CO(
        DP_OP_425J2_127_3477_n1682), .S(DP_OP_425J2_127_3477_n1683) );
  FADDX1_HVT DP_OP_425J2_127_3477_U998 ( .A(DP_OP_425J2_127_3477_n1786), .B(
        DP_OP_425J2_127_3477_n1687), .CI(DP_OP_425J2_127_3477_n1685), .CO(
        DP_OP_425J2_127_3477_n1680), .S(DP_OP_425J2_127_3477_n1681) );
  FADDX1_HVT DP_OP_425J2_127_3477_U996 ( .A(DP_OP_425J2_127_3477_n2455), .B(
        DP_OP_425J2_127_3477_n1927), .CI(DP_OP_425J2_127_3477_n1883), .CO(
        DP_OP_425J2_127_3477_n1676), .S(DP_OP_425J2_127_3477_n1677) );
  FADDX1_HVT DP_OP_425J2_127_3477_U995 ( .A(DP_OP_425J2_127_3477_n2147), .B(
        DP_OP_425J2_127_3477_n2587), .CI(DP_OP_425J2_127_3477_n2367), .CO(
        DP_OP_425J2_127_3477_n1674), .S(DP_OP_425J2_127_3477_n1675) );
  FADDX1_HVT DP_OP_425J2_127_3477_U994 ( .A(DP_OP_425J2_127_3477_n2895), .B(
        DP_OP_425J2_127_3477_n2103), .CI(DP_OP_425J2_127_3477_n2323), .CO(
        DP_OP_425J2_127_3477_n1672), .S(DP_OP_425J2_127_3477_n1673) );
  FADDX1_HVT DP_OP_425J2_127_3477_U993 ( .A(DP_OP_425J2_127_3477_n2499), .B(
        DP_OP_425J2_127_3477_n2807), .CI(DP_OP_425J2_127_3477_n2411), .CO(
        DP_OP_425J2_127_3477_n1670), .S(DP_OP_425J2_127_3477_n1671) );
  FADDX1_HVT DP_OP_425J2_127_3477_U992 ( .A(DP_OP_425J2_127_3477_n2235), .B(
        DP_OP_425J2_127_3477_n2279), .CI(DP_OP_425J2_127_3477_n2059), .CO(
        DP_OP_425J2_127_3477_n1668), .S(DP_OP_425J2_127_3477_n1669) );
  FADDX1_HVT DP_OP_425J2_127_3477_U991 ( .A(DP_OP_425J2_127_3477_n2763), .B(
        DP_OP_425J2_127_3477_n2631), .CI(DP_OP_425J2_127_3477_n2675), .CO(
        DP_OP_425J2_127_3477_n1666), .S(DP_OP_425J2_127_3477_n1667) );
  FADDX1_HVT DP_OP_425J2_127_3477_U990 ( .A(DP_OP_425J2_127_3477_n2015), .B(
        DP_OP_425J2_127_3477_n2851), .CI(DP_OP_425J2_127_3477_n2719), .CO(
        DP_OP_425J2_127_3477_n1664), .S(DP_OP_425J2_127_3477_n1665) );
  FADDX1_HVT DP_OP_425J2_127_3477_U989 ( .A(DP_OP_425J2_127_3477_n2543), .B(
        DP_OP_425J2_127_3477_n2939), .CI(DP_OP_425J2_127_3477_n2191), .CO(
        DP_OP_425J2_127_3477_n1662), .S(DP_OP_425J2_127_3477_n1663) );
  FADDX1_HVT DP_OP_425J2_127_3477_U988 ( .A(DP_OP_425J2_127_3477_n1971), .B(
        DP_OP_425J2_127_3477_n1679), .CI(DP_OP_425J2_127_3477_n1948), .CO(
        DP_OP_425J2_127_3477_n1660), .S(DP_OP_425J2_127_3477_n1661) );
  FADDX1_HVT DP_OP_425J2_127_3477_U987 ( .A(DP_OP_425J2_127_3477_n1978), .B(
        DP_OP_425J2_127_3477_n1941), .CI(DP_OP_425J2_127_3477_n1934), .CO(
        DP_OP_425J2_127_3477_n1658), .S(DP_OP_425J2_127_3477_n1659) );
  FADDX1_HVT DP_OP_425J2_127_3477_U986 ( .A(DP_OP_425J2_127_3477_n1992), .B(
        DP_OP_425J2_127_3477_n1985), .CI(DP_OP_425J2_127_3477_n2022), .CO(
        DP_OP_425J2_127_3477_n1656), .S(DP_OP_425J2_127_3477_n1657) );
  FADDX1_HVT DP_OP_425J2_127_3477_U985 ( .A(DP_OP_425J2_127_3477_n2036), .B(
        DP_OP_425J2_127_3477_n2029), .CI(DP_OP_425J2_127_3477_n2066), .CO(
        DP_OP_425J2_127_3477_n1654), .S(DP_OP_425J2_127_3477_n1655) );
  FADDX1_HVT DP_OP_425J2_127_3477_U984 ( .A(DP_OP_425J2_127_3477_n3002), .B(
        DP_OP_425J2_127_3477_n2073), .CI(DP_OP_425J2_127_3477_n2080), .CO(
        DP_OP_425J2_127_3477_n1652), .S(DP_OP_425J2_127_3477_n1653) );
  FADDX1_HVT DP_OP_425J2_127_3477_U983 ( .A(DP_OP_425J2_127_3477_n2513), .B(
        DP_OP_425J2_127_3477_n2995), .CI(DP_OP_425J2_127_3477_n2988), .CO(
        DP_OP_425J2_127_3477_n1650), .S(DP_OP_425J2_127_3477_n1651) );
  FADDX1_HVT DP_OP_425J2_127_3477_U982 ( .A(DP_OP_425J2_127_3477_n2476), .B(
        DP_OP_425J2_127_3477_n2110), .CI(DP_OP_425J2_127_3477_n2960), .CO(
        DP_OP_425J2_127_3477_n1648), .S(DP_OP_425J2_127_3477_n1649) );
  FADDX1_HVT DP_OP_425J2_127_3477_U981 ( .A(DP_OP_425J2_127_3477_n2506), .B(
        DP_OP_425J2_127_3477_n2117), .CI(DP_OP_425J2_127_3477_n2953), .CO(
        DP_OP_425J2_127_3477_n1646), .S(DP_OP_425J2_127_3477_n1647) );
  FADDX1_HVT DP_OP_425J2_127_3477_U980 ( .A(DP_OP_425J2_127_3477_n2946), .B(
        DP_OP_425J2_127_3477_n2124), .CI(DP_OP_425J2_127_3477_n2154), .CO(
        DP_OP_425J2_127_3477_n1644), .S(DP_OP_425J2_127_3477_n1645) );
  FADDX1_HVT DP_OP_425J2_127_3477_U979 ( .A(DP_OP_425J2_127_3477_n2469), .B(
        DP_OP_425J2_127_3477_n2161), .CI(DP_OP_425J2_127_3477_n2168), .CO(
        DP_OP_425J2_127_3477_n1642), .S(DP_OP_425J2_127_3477_n1643) );
  FADDX1_HVT DP_OP_425J2_127_3477_U978 ( .A(DP_OP_425J2_127_3477_n2550), .B(
        DP_OP_425J2_127_3477_n2198), .CI(DP_OP_425J2_127_3477_n2205), .CO(
        DP_OP_425J2_127_3477_n1640), .S(DP_OP_425J2_127_3477_n1641) );
  FADDX1_HVT DP_OP_425J2_127_3477_U977 ( .A(DP_OP_425J2_127_3477_n2557), .B(
        DP_OP_425J2_127_3477_n2212), .CI(DP_OP_425J2_127_3477_n2242), .CO(
        DP_OP_425J2_127_3477_n1638), .S(DP_OP_425J2_127_3477_n1639) );
  FADDX1_HVT DP_OP_425J2_127_3477_U976 ( .A(DP_OP_425J2_127_3477_n2564), .B(
        DP_OP_425J2_127_3477_n2916), .CI(DP_OP_425J2_127_3477_n2249), .CO(
        DP_OP_425J2_127_3477_n1636), .S(DP_OP_425J2_127_3477_n1637) );
  FADDX1_HVT DP_OP_425J2_127_3477_U975 ( .A(DP_OP_425J2_127_3477_n2594), .B(
        DP_OP_425J2_127_3477_n2256), .CI(DP_OP_425J2_127_3477_n2909), .CO(
        DP_OP_425J2_127_3477_n1634), .S(DP_OP_425J2_127_3477_n1635) );
  FADDX1_HVT DP_OP_425J2_127_3477_U974 ( .A(DP_OP_425J2_127_3477_n2520), .B(
        DP_OP_425J2_127_3477_n2902), .CI(DP_OP_425J2_127_3477_n2872), .CO(
        DP_OP_425J2_127_3477_n1632), .S(DP_OP_425J2_127_3477_n1633) );
  FADDX1_HVT DP_OP_425J2_127_3477_U973 ( .A(DP_OP_425J2_127_3477_n2432), .B(
        DP_OP_425J2_127_3477_n2865), .CI(DP_OP_425J2_127_3477_n2286), .CO(
        DP_OP_425J2_127_3477_n1630), .S(DP_OP_425J2_127_3477_n1631) );
  FADDX1_HVT DP_OP_425J2_127_3477_U972 ( .A(DP_OP_425J2_127_3477_n2858), .B(
        DP_OP_425J2_127_3477_n2293), .CI(DP_OP_425J2_127_3477_n2828), .CO(
        DP_OP_425J2_127_3477_n1628), .S(DP_OP_425J2_127_3477_n1629) );
  FADDX1_HVT DP_OP_425J2_127_3477_U971 ( .A(DP_OP_425J2_127_3477_n2821), .B(
        DP_OP_425J2_127_3477_n2814), .CI(DP_OP_425J2_127_3477_n2300), .CO(
        DP_OP_425J2_127_3477_n1626), .S(DP_OP_425J2_127_3477_n1627) );
  FADDX1_HVT DP_OP_425J2_127_3477_U970 ( .A(DP_OP_425J2_127_3477_n2425), .B(
        DP_OP_425J2_127_3477_n2330), .CI(DP_OP_425J2_127_3477_n2784), .CO(
        DP_OP_425J2_127_3477_n1624), .S(DP_OP_425J2_127_3477_n1625) );
  FADDX1_HVT DP_OP_425J2_127_3477_U969 ( .A(DP_OP_425J2_127_3477_n2418), .B(
        DP_OP_425J2_127_3477_n2777), .CI(DP_OP_425J2_127_3477_n2770), .CO(
        DP_OP_425J2_127_3477_n1622), .S(DP_OP_425J2_127_3477_n1623) );
  FADDX1_HVT DP_OP_425J2_127_3477_U968 ( .A(DP_OP_425J2_127_3477_n2374), .B(
        DP_OP_425J2_127_3477_n2740), .CI(DP_OP_425J2_127_3477_n2733), .CO(
        DP_OP_425J2_127_3477_n1620), .S(DP_OP_425J2_127_3477_n1621) );
  FADDX1_HVT DP_OP_425J2_127_3477_U967 ( .A(DP_OP_425J2_127_3477_n2337), .B(
        DP_OP_425J2_127_3477_n2726), .CI(DP_OP_425J2_127_3477_n2696), .CO(
        DP_OP_425J2_127_3477_n1618), .S(DP_OP_425J2_127_3477_n1619) );
  FADDX1_HVT DP_OP_425J2_127_3477_U966 ( .A(DP_OP_425J2_127_3477_n2608), .B(
        DP_OP_425J2_127_3477_n2689), .CI(DP_OP_425J2_127_3477_n2344), .CO(
        DP_OP_425J2_127_3477_n1616), .S(DP_OP_425J2_127_3477_n1617) );
  FADDX1_HVT DP_OP_425J2_127_3477_U965 ( .A(DP_OP_425J2_127_3477_n2462), .B(
        DP_OP_425J2_127_3477_n2381), .CI(DP_OP_425J2_127_3477_n2682), .CO(
        DP_OP_425J2_127_3477_n1614), .S(DP_OP_425J2_127_3477_n1615) );
  FADDX1_HVT DP_OP_425J2_127_3477_U964 ( .A(DP_OP_425J2_127_3477_n2652), .B(
        DP_OP_425J2_127_3477_n2388), .CI(DP_OP_425J2_127_3477_n2601), .CO(
        DP_OP_425J2_127_3477_n1612), .S(DP_OP_425J2_127_3477_n1613) );
  FADDX1_HVT DP_OP_425J2_127_3477_U963 ( .A(DP_OP_425J2_127_3477_n2645), .B(
        DP_OP_425J2_127_3477_n2638), .CI(DP_OP_425J2_127_3477_n1784), .CO(
        DP_OP_425J2_127_3477_n1610), .S(DP_OP_425J2_127_3477_n1611) );
  FADDX1_HVT DP_OP_425J2_127_3477_U962 ( .A(DP_OP_425J2_127_3477_n1760), .B(
        DP_OP_425J2_127_3477_n1782), .CI(DP_OP_425J2_127_3477_n1736), .CO(
        DP_OP_425J2_127_3477_n1608), .S(DP_OP_425J2_127_3477_n1609) );
  FADDX1_HVT DP_OP_425J2_127_3477_U961 ( .A(DP_OP_425J2_127_3477_n1758), .B(
        DP_OP_425J2_127_3477_n1780), .CI(DP_OP_425J2_127_3477_n1778), .CO(
        DP_OP_425J2_127_3477_n1606), .S(DP_OP_425J2_127_3477_n1607) );
  FADDX1_HVT DP_OP_425J2_127_3477_U960 ( .A(DP_OP_425J2_127_3477_n1752), .B(
        DP_OP_425J2_127_3477_n1776), .CI(DP_OP_425J2_127_3477_n1774), .CO(
        DP_OP_425J2_127_3477_n1604), .S(DP_OP_425J2_127_3477_n1605) );
  FADDX1_HVT DP_OP_425J2_127_3477_U959 ( .A(DP_OP_425J2_127_3477_n1748), .B(
        DP_OP_425J2_127_3477_n1738), .CI(DP_OP_425J2_127_3477_n1740), .CO(
        DP_OP_425J2_127_3477_n1602), .S(DP_OP_425J2_127_3477_n1603) );
  FADDX1_HVT DP_OP_425J2_127_3477_U958 ( .A(DP_OP_425J2_127_3477_n1746), .B(
        DP_OP_425J2_127_3477_n1772), .CI(DP_OP_425J2_127_3477_n1742), .CO(
        DP_OP_425J2_127_3477_n1600), .S(DP_OP_425J2_127_3477_n1601) );
  FADDX1_HVT DP_OP_425J2_127_3477_U957 ( .A(DP_OP_425J2_127_3477_n1744), .B(
        DP_OP_425J2_127_3477_n1770), .CI(DP_OP_425J2_127_3477_n1768), .CO(
        DP_OP_425J2_127_3477_n1598), .S(DP_OP_425J2_127_3477_n1599) );
  FADDX1_HVT DP_OP_425J2_127_3477_U956 ( .A(DP_OP_425J2_127_3477_n1756), .B(
        DP_OP_425J2_127_3477_n1766), .CI(DP_OP_425J2_127_3477_n1750), .CO(
        DP_OP_425J2_127_3477_n1596), .S(DP_OP_425J2_127_3477_n1597) );
  FADDX1_HVT DP_OP_425J2_127_3477_U955 ( .A(DP_OP_425J2_127_3477_n1764), .B(
        DP_OP_425J2_127_3477_n1762), .CI(DP_OP_425J2_127_3477_n1754), .CO(
        DP_OP_425J2_127_3477_n1594), .S(DP_OP_425J2_127_3477_n1595) );
  FADDX1_HVT DP_OP_425J2_127_3477_U954 ( .A(DP_OP_425J2_127_3477_n1673), .B(
        DP_OP_425J2_127_3477_n1675), .CI(DP_OP_425J2_127_3477_n1661), .CO(
        DP_OP_425J2_127_3477_n1592), .S(DP_OP_425J2_127_3477_n1593) );
  FADDX1_HVT DP_OP_425J2_127_3477_U953 ( .A(DP_OP_425J2_127_3477_n1667), .B(
        DP_OP_425J2_127_3477_n1669), .CI(DP_OP_425J2_127_3477_n1734), .CO(
        DP_OP_425J2_127_3477_n1590), .S(DP_OP_425J2_127_3477_n1591) );
  FADDX1_HVT DP_OP_425J2_127_3477_U952 ( .A(DP_OP_425J2_127_3477_n1663), .B(
        DP_OP_425J2_127_3477_n1665), .CI(DP_OP_425J2_127_3477_n1671), .CO(
        DP_OP_425J2_127_3477_n1588), .S(DP_OP_425J2_127_3477_n1589) );
  FADDX1_HVT DP_OP_425J2_127_3477_U951 ( .A(DP_OP_425J2_127_3477_n1677), .B(
        DP_OP_425J2_127_3477_n1627), .CI(DP_OP_425J2_127_3477_n1625), .CO(
        DP_OP_425J2_127_3477_n1586), .S(DP_OP_425J2_127_3477_n1587) );
  FADDX1_HVT DP_OP_425J2_127_3477_U950 ( .A(DP_OP_425J2_127_3477_n1629), .B(
        DP_OP_425J2_127_3477_n1645), .CI(DP_OP_425J2_127_3477_n1653), .CO(
        DP_OP_425J2_127_3477_n1584), .S(DP_OP_425J2_127_3477_n1585) );
  FADDX1_HVT DP_OP_425J2_127_3477_U949 ( .A(DP_OP_425J2_127_3477_n1621), .B(
        DP_OP_425J2_127_3477_n1641), .CI(DP_OP_425J2_127_3477_n1639), .CO(
        DP_OP_425J2_127_3477_n1582), .S(DP_OP_425J2_127_3477_n1583) );
  FADDX1_HVT DP_OP_425J2_127_3477_U948 ( .A(DP_OP_425J2_127_3477_n1619), .B(
        DP_OP_425J2_127_3477_n1655), .CI(DP_OP_425J2_127_3477_n1643), .CO(
        DP_OP_425J2_127_3477_n1580), .S(DP_OP_425J2_127_3477_n1581) );
  FADDX1_HVT DP_OP_425J2_127_3477_U947 ( .A(DP_OP_425J2_127_3477_n1617), .B(
        DP_OP_425J2_127_3477_n1649), .CI(DP_OP_425J2_127_3477_n1651), .CO(
        DP_OP_425J2_127_3477_n1578), .S(DP_OP_425J2_127_3477_n1579) );
  FADDX1_HVT DP_OP_425J2_127_3477_U946 ( .A(DP_OP_425J2_127_3477_n1615), .B(
        DP_OP_425J2_127_3477_n1647), .CI(DP_OP_425J2_127_3477_n1659), .CO(
        DP_OP_425J2_127_3477_n1576), .S(DP_OP_425J2_127_3477_n1577) );
  FADDX1_HVT DP_OP_425J2_127_3477_U945 ( .A(DP_OP_425J2_127_3477_n1637), .B(
        DP_OP_425J2_127_3477_n1657), .CI(DP_OP_425J2_127_3477_n1613), .CO(
        DP_OP_425J2_127_3477_n1574), .S(DP_OP_425J2_127_3477_n1575) );
  FADDX1_HVT DP_OP_425J2_127_3477_U944 ( .A(DP_OP_425J2_127_3477_n1623), .B(
        DP_OP_425J2_127_3477_n1633), .CI(DP_OP_425J2_127_3477_n1635), .CO(
        DP_OP_425J2_127_3477_n1572), .S(DP_OP_425J2_127_3477_n1573) );
  FADDX1_HVT DP_OP_425J2_127_3477_U943 ( .A(DP_OP_425J2_127_3477_n1631), .B(
        DP_OP_425J2_127_3477_n1611), .CI(DP_OP_425J2_127_3477_n1732), .CO(
        DP_OP_425J2_127_3477_n1570), .S(DP_OP_425J2_127_3477_n1571) );
  FADDX1_HVT DP_OP_425J2_127_3477_U942 ( .A(DP_OP_425J2_127_3477_n1730), .B(
        DP_OP_425J2_127_3477_n1728), .CI(DP_OP_425J2_127_3477_n1726), .CO(
        DP_OP_425J2_127_3477_n1568), .S(DP_OP_425J2_127_3477_n1569) );
  FADDX1_HVT DP_OP_425J2_127_3477_U941 ( .A(DP_OP_425J2_127_3477_n1724), .B(
        DP_OP_425J2_127_3477_n1722), .CI(DP_OP_425J2_127_3477_n1710), .CO(
        DP_OP_425J2_127_3477_n1566), .S(DP_OP_425J2_127_3477_n1567) );
  FADDX1_HVT DP_OP_425J2_127_3477_U940 ( .A(DP_OP_425J2_127_3477_n1708), .B(
        DP_OP_425J2_127_3477_n1609), .CI(DP_OP_425J2_127_3477_n1706), .CO(
        DP_OP_425J2_127_3477_n1564), .S(DP_OP_425J2_127_3477_n1565) );
  FADDX1_HVT DP_OP_425J2_127_3477_U939 ( .A(DP_OP_425J2_127_3477_n1720), .B(
        DP_OP_425J2_127_3477_n1599), .CI(DP_OP_425J2_127_3477_n1607), .CO(
        DP_OP_425J2_127_3477_n1562), .S(DP_OP_425J2_127_3477_n1563) );
  FADDX1_HVT DP_OP_425J2_127_3477_U938 ( .A(DP_OP_425J2_127_3477_n1718), .B(
        DP_OP_425J2_127_3477_n1597), .CI(DP_OP_425J2_127_3477_n1601), .CO(
        DP_OP_425J2_127_3477_n1560), .S(DP_OP_425J2_127_3477_n1561) );
  FADDX1_HVT DP_OP_425J2_127_3477_U937 ( .A(DP_OP_425J2_127_3477_n1714), .B(
        DP_OP_425J2_127_3477_n1605), .CI(DP_OP_425J2_127_3477_n1603), .CO(
        DP_OP_425J2_127_3477_n1558), .S(DP_OP_425J2_127_3477_n1559) );
  FADDX1_HVT DP_OP_425J2_127_3477_U936 ( .A(DP_OP_425J2_127_3477_n1712), .B(
        DP_OP_425J2_127_3477_n1716), .CI(DP_OP_425J2_127_3477_n1595), .CO(
        DP_OP_425J2_127_3477_n1556), .S(DP_OP_425J2_127_3477_n1557) );
  FADDX1_HVT DP_OP_425J2_127_3477_U935 ( .A(DP_OP_425J2_127_3477_n1591), .B(
        DP_OP_425J2_127_3477_n1593), .CI(DP_OP_425J2_127_3477_n1587), .CO(
        DP_OP_425J2_127_3477_n1554), .S(DP_OP_425J2_127_3477_n1555) );
  FADDX1_HVT DP_OP_425J2_127_3477_U934 ( .A(DP_OP_425J2_127_3477_n1589), .B(
        DP_OP_425J2_127_3477_n1575), .CI(DP_OP_425J2_127_3477_n1577), .CO(
        DP_OP_425J2_127_3477_n1552), .S(DP_OP_425J2_127_3477_n1553) );
  FADDX1_HVT DP_OP_425J2_127_3477_U933 ( .A(DP_OP_425J2_127_3477_n1583), .B(
        DP_OP_425J2_127_3477_n1581), .CI(DP_OP_425J2_127_3477_n1704), .CO(
        DP_OP_425J2_127_3477_n1550), .S(DP_OP_425J2_127_3477_n1551) );
  FADDX1_HVT DP_OP_425J2_127_3477_U932 ( .A(DP_OP_425J2_127_3477_n1579), .B(
        DP_OP_425J2_127_3477_n1573), .CI(DP_OP_425J2_127_3477_n1585), .CO(
        DP_OP_425J2_127_3477_n1548), .S(DP_OP_425J2_127_3477_n1549) );
  FADDX1_HVT DP_OP_425J2_127_3477_U931 ( .A(DP_OP_425J2_127_3477_n1571), .B(
        DP_OP_425J2_127_3477_n1702), .CI(DP_OP_425J2_127_3477_n1698), .CO(
        DP_OP_425J2_127_3477_n1546), .S(DP_OP_425J2_127_3477_n1547) );
  FADDX1_HVT DP_OP_425J2_127_3477_U930 ( .A(DP_OP_425J2_127_3477_n1700), .B(
        DP_OP_425J2_127_3477_n1569), .CI(DP_OP_425J2_127_3477_n1696), .CO(
        DP_OP_425J2_127_3477_n1544), .S(DP_OP_425J2_127_3477_n1545) );
  FADDX1_HVT DP_OP_425J2_127_3477_U929 ( .A(DP_OP_425J2_127_3477_n1567), .B(
        DP_OP_425J2_127_3477_n1557), .CI(DP_OP_425J2_127_3477_n1559), .CO(
        DP_OP_425J2_127_3477_n1542), .S(DP_OP_425J2_127_3477_n1543) );
  FADDX1_HVT DP_OP_425J2_127_3477_U928 ( .A(DP_OP_425J2_127_3477_n1694), .B(
        DP_OP_425J2_127_3477_n1561), .CI(DP_OP_425J2_127_3477_n1692), .CO(
        DP_OP_425J2_127_3477_n1540), .S(DP_OP_425J2_127_3477_n1541) );
  FADDX1_HVT DP_OP_425J2_127_3477_U927 ( .A(DP_OP_425J2_127_3477_n1565), .B(
        DP_OP_425J2_127_3477_n1563), .CI(DP_OP_425J2_127_3477_n1555), .CO(
        DP_OP_425J2_127_3477_n1538), .S(DP_OP_425J2_127_3477_n1539) );
  FADDX1_HVT DP_OP_425J2_127_3477_U926 ( .A(DP_OP_425J2_127_3477_n1690), .B(
        DP_OP_425J2_127_3477_n1553), .CI(DP_OP_425J2_127_3477_n1549), .CO(
        DP_OP_425J2_127_3477_n1536), .S(DP_OP_425J2_127_3477_n1537) );
  FADDX1_HVT DP_OP_425J2_127_3477_U925 ( .A(DP_OP_425J2_127_3477_n1551), .B(
        DP_OP_425J2_127_3477_n1688), .CI(DP_OP_425J2_127_3477_n1547), .CO(
        DP_OP_425J2_127_3477_n1534), .S(DP_OP_425J2_127_3477_n1535) );
  FADDX1_HVT DP_OP_425J2_127_3477_U924 ( .A(DP_OP_425J2_127_3477_n1686), .B(
        DP_OP_425J2_127_3477_n1545), .CI(DP_OP_425J2_127_3477_n1684), .CO(
        DP_OP_425J2_127_3477_n1532), .S(DP_OP_425J2_127_3477_n1533) );
  FADDX1_HVT DP_OP_425J2_127_3477_U923 ( .A(DP_OP_425J2_127_3477_n1543), .B(
        DP_OP_425J2_127_3477_n1541), .CI(DP_OP_425J2_127_3477_n1539), .CO(
        DP_OP_425J2_127_3477_n1530), .S(DP_OP_425J2_127_3477_n1531) );
  FADDX1_HVT DP_OP_425J2_127_3477_U922 ( .A(DP_OP_425J2_127_3477_n1537), .B(
        DP_OP_425J2_127_3477_n1682), .CI(DP_OP_425J2_127_3477_n1535), .CO(
        DP_OP_425J2_127_3477_n1528), .S(DP_OP_425J2_127_3477_n1529) );
  FADDX1_HVT DP_OP_425J2_127_3477_U921 ( .A(DP_OP_425J2_127_3477_n1680), .B(
        DP_OP_425J2_127_3477_n1533), .CI(DP_OP_425J2_127_3477_n1531), .CO(
        DP_OP_425J2_127_3477_n1526), .S(DP_OP_425J2_127_3477_n1527) );
  FADDX1_HVT DP_OP_425J2_127_3477_U920 ( .A(DP_OP_425J2_127_3477_n1678), .B(
        DP_OP_425J2_127_3477_n1926), .CI(DP_OP_425J2_127_3477_n1882), .CO(
        DP_OP_425J2_127_3477_n1524), .S(DP_OP_425J2_127_3477_n1525) );
  FADDX1_HVT DP_OP_425J2_127_3477_U919 ( .A(DP_OP_425J2_127_3477_n2981), .B(
        DP_OP_425J2_127_3477_n2498), .CI(DP_OP_425J2_127_3477_n2366), .CO(
        DP_OP_425J2_127_3477_n1522), .S(DP_OP_425J2_127_3477_n1523) );
  FADDX1_HVT DP_OP_425J2_127_3477_U918 ( .A(DP_OP_425J2_127_3477_n2894), .B(
        DP_OP_425J2_127_3477_n2630), .CI(DP_OP_425J2_127_3477_n2278), .CO(
        DP_OP_425J2_127_3477_n1520), .S(DP_OP_425J2_127_3477_n1521) );
  FADDX1_HVT DP_OP_425J2_127_3477_U917 ( .A(DP_OP_425J2_127_3477_n2058), .B(
        DP_OP_425J2_127_3477_n2586), .CI(DP_OP_425J2_127_3477_n2806), .CO(
        DP_OP_425J2_127_3477_n1518), .S(DP_OP_425J2_127_3477_n1519) );
  FADDX1_HVT DP_OP_425J2_127_3477_U916 ( .A(DP_OP_425J2_127_3477_n2146), .B(
        DP_OP_425J2_127_3477_n2322), .CI(DP_OP_425J2_127_3477_n2410), .CO(
        DP_OP_425J2_127_3477_n1516), .S(DP_OP_425J2_127_3477_n1517) );
  FADDX1_HVT DP_OP_425J2_127_3477_U915 ( .A(DP_OP_425J2_127_3477_n2762), .B(
        DP_OP_425J2_127_3477_n2234), .CI(DP_OP_425J2_127_3477_n2850), .CO(
        DP_OP_425J2_127_3477_n1514), .S(DP_OP_425J2_127_3477_n1515) );
  FADDX1_HVT DP_OP_425J2_127_3477_U914 ( .A(DP_OP_425J2_127_3477_n2102), .B(
        DP_OP_425J2_127_3477_n2454), .CI(DP_OP_425J2_127_3477_n2542), .CO(
        DP_OP_425J2_127_3477_n1512), .S(DP_OP_425J2_127_3477_n1513) );
  FADDX1_HVT DP_OP_425J2_127_3477_U913 ( .A(DP_OP_425J2_127_3477_n2938), .B(
        DP_OP_425J2_127_3477_n2674), .CI(DP_OP_425J2_127_3477_n2718), .CO(
        DP_OP_425J2_127_3477_n1510), .S(DP_OP_425J2_127_3477_n1511) );
  FADDX1_HVT DP_OP_425J2_127_3477_U912 ( .A(DP_OP_425J2_127_3477_n2014), .B(
        DP_OP_425J2_127_3477_n2190), .CI(DP_OP_425J2_127_3477_n1970), .CO(
        DP_OP_425J2_127_3477_n1508), .S(DP_OP_425J2_127_3477_n1509) );
  FADDX1_HVT DP_OP_425J2_127_3477_U911 ( .A(DP_OP_425J2_127_3477_n2505), .B(
        DP_OP_425J2_127_3477_n1940), .CI(DP_OP_425J2_127_3477_n1933), .CO(
        DP_OP_425J2_127_3477_n1506), .S(DP_OP_425J2_127_3477_n1507) );
  FADDX1_HVT DP_OP_425J2_127_3477_U910 ( .A(DP_OP_425J2_127_3477_n3001), .B(
        DP_OP_425J2_127_3477_n1947), .CI(DP_OP_425J2_127_3477_n1977), .CO(
        DP_OP_425J2_127_3477_n1504), .S(DP_OP_425J2_127_3477_n1505) );
  FADDX1_HVT DP_OP_425J2_127_3477_U909 ( .A(DP_OP_425J2_127_3477_n2387), .B(
        DP_OP_425J2_127_3477_n2994), .CI(DP_OP_425J2_127_3477_n1984), .CO(
        DP_OP_425J2_127_3477_n1502), .S(DP_OP_425J2_127_3477_n1503) );
  FADDX1_HVT DP_OP_425J2_127_3477_U908 ( .A(DP_OP_425J2_127_3477_n2380), .B(
        DP_OP_425J2_127_3477_n2987), .CI(DP_OP_425J2_127_3477_n1991), .CO(
        DP_OP_425J2_127_3477_n1500), .S(DP_OP_425J2_127_3477_n1501) );
  FADDX1_HVT DP_OP_425J2_127_3477_U907 ( .A(DP_OP_425J2_127_3477_n2959), .B(
        DP_OP_425J2_127_3477_n2021), .CI(DP_OP_425J2_127_3477_n2028), .CO(
        DP_OP_425J2_127_3477_n1498), .S(DP_OP_425J2_127_3477_n1499) );
  FADDX1_HVT DP_OP_425J2_127_3477_U906 ( .A(DP_OP_425J2_127_3477_n2417), .B(
        DP_OP_425J2_127_3477_n2952), .CI(DP_OP_425J2_127_3477_n2945), .CO(
        DP_OP_425J2_127_3477_n1496), .S(DP_OP_425J2_127_3477_n1497) );
  FADDX1_HVT DP_OP_425J2_127_3477_U905 ( .A(DP_OP_425J2_127_3477_n2343), .B(
        DP_OP_425J2_127_3477_n2915), .CI(DP_OP_425J2_127_3477_n2908), .CO(
        DP_OP_425J2_127_3477_n1494), .S(DP_OP_425J2_127_3477_n1495) );
  FADDX1_HVT DP_OP_425J2_127_3477_U904 ( .A(DP_OP_425J2_127_3477_n2336), .B(
        DP_OP_425J2_127_3477_n2901), .CI(DP_OP_425J2_127_3477_n2035), .CO(
        DP_OP_425J2_127_3477_n1492), .S(DP_OP_425J2_127_3477_n1493) );
  FADDX1_HVT DP_OP_425J2_127_3477_U903 ( .A(DP_OP_425J2_127_3477_n2329), .B(
        DP_OP_425J2_127_3477_n2871), .CI(DP_OP_425J2_127_3477_n2864), .CO(
        DP_OP_425J2_127_3477_n1490), .S(DP_OP_425J2_127_3477_n1491) );
  FADDX1_HVT DP_OP_425J2_127_3477_U902 ( .A(DP_OP_425J2_127_3477_n2299), .B(
        DP_OP_425J2_127_3477_n2857), .CI(DP_OP_425J2_127_3477_n2065), .CO(
        DP_OP_425J2_127_3477_n1488), .S(DP_OP_425J2_127_3477_n1489) );
  FADDX1_HVT DP_OP_425J2_127_3477_U901 ( .A(DP_OP_425J2_127_3477_n2292), .B(
        DP_OP_425J2_127_3477_n2072), .CI(DP_OP_425J2_127_3477_n2079), .CO(
        DP_OP_425J2_127_3477_n1486), .S(DP_OP_425J2_127_3477_n1487) );
  FADDX1_HVT DP_OP_425J2_127_3477_U900 ( .A(DP_OP_425J2_127_3477_n2373), .B(
        DP_OP_425J2_127_3477_n2109), .CI(DP_OP_425J2_127_3477_n2827), .CO(
        DP_OP_425J2_127_3477_n1484), .S(DP_OP_425J2_127_3477_n1485) );
  FADDX1_HVT DP_OP_425J2_127_3477_U899 ( .A(DP_OP_425J2_127_3477_n2424), .B(
        DP_OP_425J2_127_3477_n2820), .CI(DP_OP_425J2_127_3477_n2813), .CO(
        DP_OP_425J2_127_3477_n1482), .S(DP_OP_425J2_127_3477_n1483) );
  FADDX1_HVT DP_OP_425J2_127_3477_U898 ( .A(DP_OP_425J2_127_3477_n2783), .B(
        DP_OP_425J2_127_3477_n2116), .CI(DP_OP_425J2_127_3477_n2123), .CO(
        DP_OP_425J2_127_3477_n1480), .S(DP_OP_425J2_127_3477_n1481) );
  FADDX1_HVT DP_OP_425J2_127_3477_U897 ( .A(DP_OP_425J2_127_3477_n2556), .B(
        DP_OP_425J2_127_3477_n2153), .CI(DP_OP_425J2_127_3477_n2160), .CO(
        DP_OP_425J2_127_3477_n1478), .S(DP_OP_425J2_127_3477_n1479) );
  FADDX1_HVT DP_OP_425J2_127_3477_U896 ( .A(DP_OP_425J2_127_3477_n2776), .B(
        DP_OP_425J2_127_3477_n2167), .CI(DP_OP_425J2_127_3477_n2197), .CO(
        DP_OP_425J2_127_3477_n1476), .S(DP_OP_425J2_127_3477_n1477) );
  FADDX1_HVT DP_OP_425J2_127_3477_U895 ( .A(DP_OP_425J2_127_3477_n2769), .B(
        DP_OP_425J2_127_3477_n2204), .CI(DP_OP_425J2_127_3477_n2211), .CO(
        DP_OP_425J2_127_3477_n1474), .S(DP_OP_425J2_127_3477_n1475) );
  FADDX1_HVT DP_OP_425J2_127_3477_U894 ( .A(DP_OP_425J2_127_3477_n2739), .B(
        DP_OP_425J2_127_3477_n2241), .CI(DP_OP_425J2_127_3477_n2248), .CO(
        DP_OP_425J2_127_3477_n1472), .S(DP_OP_425J2_127_3477_n1473) );
  FADDX1_HVT DP_OP_425J2_127_3477_U893 ( .A(DP_OP_425J2_127_3477_n2732), .B(
        DP_OP_425J2_127_3477_n2255), .CI(DP_OP_425J2_127_3477_n2285), .CO(
        DP_OP_425J2_127_3477_n1470), .S(DP_OP_425J2_127_3477_n1471) );
  FADDX1_HVT DP_OP_425J2_127_3477_U892 ( .A(DP_OP_425J2_127_3477_n2725), .B(
        DP_OP_425J2_127_3477_n2431), .CI(DP_OP_425J2_127_3477_n2461), .CO(
        DP_OP_425J2_127_3477_n1468), .S(DP_OP_425J2_127_3477_n1469) );
  FADDX1_HVT DP_OP_425J2_127_3477_U891 ( .A(DP_OP_425J2_127_3477_n2695), .B(
        DP_OP_425J2_127_3477_n2468), .CI(DP_OP_425J2_127_3477_n2688), .CO(
        DP_OP_425J2_127_3477_n1466), .S(DP_OP_425J2_127_3477_n1467) );
  FADDX1_HVT DP_OP_425J2_127_3477_U890 ( .A(DP_OP_425J2_127_3477_n2593), .B(
        DP_OP_425J2_127_3477_n2475), .CI(DP_OP_425J2_127_3477_n2512), .CO(
        DP_OP_425J2_127_3477_n1464), .S(DP_OP_425J2_127_3477_n1465) );
  FADDX1_HVT DP_OP_425J2_127_3477_U889 ( .A(DP_OP_425J2_127_3477_n2563), .B(
        DP_OP_425J2_127_3477_n2519), .CI(DP_OP_425J2_127_3477_n2681), .CO(
        DP_OP_425J2_127_3477_n1462), .S(DP_OP_425J2_127_3477_n1463) );
  FADDX1_HVT DP_OP_425J2_127_3477_U888 ( .A(DP_OP_425J2_127_3477_n2637), .B(
        DP_OP_425J2_127_3477_n2549), .CI(DP_OP_425J2_127_3477_n2651), .CO(
        DP_OP_425J2_127_3477_n1460), .S(DP_OP_425J2_127_3477_n1461) );
  FADDX1_HVT DP_OP_425J2_127_3477_U887 ( .A(DP_OP_425J2_127_3477_n2600), .B(
        DP_OP_425J2_127_3477_n2607), .CI(DP_OP_425J2_127_3477_n2644), .CO(
        DP_OP_425J2_127_3477_n1458), .S(DP_OP_425J2_127_3477_n1459) );
  FADDX1_HVT DP_OP_425J2_127_3477_U886 ( .A(DP_OP_425J2_127_3477_n1666), .B(
        DP_OP_425J2_127_3477_n1662), .CI(DP_OP_425J2_127_3477_n1660), .CO(
        DP_OP_425J2_127_3477_n1456), .S(DP_OP_425J2_127_3477_n1457) );
  FADDX1_HVT DP_OP_425J2_127_3477_U885 ( .A(DP_OP_425J2_127_3477_n1664), .B(
        DP_OP_425J2_127_3477_n1668), .CI(DP_OP_425J2_127_3477_n1670), .CO(
        DP_OP_425J2_127_3477_n1454), .S(DP_OP_425J2_127_3477_n1455) );
  FADDX1_HVT DP_OP_425J2_127_3477_U884 ( .A(DP_OP_425J2_127_3477_n1672), .B(
        DP_OP_425J2_127_3477_n1674), .CI(DP_OP_425J2_127_3477_n1676), .CO(
        DP_OP_425J2_127_3477_n1452), .S(DP_OP_425J2_127_3477_n1453) );
  FADDX1_HVT DP_OP_425J2_127_3477_U883 ( .A(DP_OP_425J2_127_3477_n1636), .B(
        DP_OP_425J2_127_3477_n1658), .CI(DP_OP_425J2_127_3477_n1656), .CO(
        DP_OP_425J2_127_3477_n1450), .S(DP_OP_425J2_127_3477_n1451) );
  FADDX1_HVT DP_OP_425J2_127_3477_U882 ( .A(DP_OP_425J2_127_3477_n1632), .B(
        DP_OP_425J2_127_3477_n1654), .CI(DP_OP_425J2_127_3477_n1652), .CO(
        DP_OP_425J2_127_3477_n1448), .S(DP_OP_425J2_127_3477_n1449) );
  FADDX1_HVT DP_OP_425J2_127_3477_U881 ( .A(DP_OP_425J2_127_3477_n1626), .B(
        DP_OP_425J2_127_3477_n1650), .CI(DP_OP_425J2_127_3477_n1648), .CO(
        DP_OP_425J2_127_3477_n1446), .S(DP_OP_425J2_127_3477_n1447) );
  FADDX1_HVT DP_OP_425J2_127_3477_U880 ( .A(DP_OP_425J2_127_3477_n1622), .B(
        DP_OP_425J2_127_3477_n1646), .CI(DP_OP_425J2_127_3477_n1612), .CO(
        DP_OP_425J2_127_3477_n1444), .S(DP_OP_425J2_127_3477_n1445) );
  FADDX1_HVT DP_OP_425J2_127_3477_U879 ( .A(DP_OP_425J2_127_3477_n1618), .B(
        DP_OP_425J2_127_3477_n1644), .CI(DP_OP_425J2_127_3477_n1642), .CO(
        DP_OP_425J2_127_3477_n1442), .S(DP_OP_425J2_127_3477_n1443) );
  FADDX1_HVT DP_OP_425J2_127_3477_U878 ( .A(DP_OP_425J2_127_3477_n1628), .B(
        DP_OP_425J2_127_3477_n1640), .CI(DP_OP_425J2_127_3477_n1638), .CO(
        DP_OP_425J2_127_3477_n1440), .S(DP_OP_425J2_127_3477_n1441) );
  FADDX1_HVT DP_OP_425J2_127_3477_U877 ( .A(DP_OP_425J2_127_3477_n1620), .B(
        DP_OP_425J2_127_3477_n1634), .CI(DP_OP_425J2_127_3477_n1630), .CO(
        DP_OP_425J2_127_3477_n1438), .S(DP_OP_425J2_127_3477_n1439) );
  FADDX1_HVT DP_OP_425J2_127_3477_U876 ( .A(DP_OP_425J2_127_3477_n1616), .B(
        DP_OP_425J2_127_3477_n1624), .CI(DP_OP_425J2_127_3477_n1614), .CO(
        DP_OP_425J2_127_3477_n1436), .S(DP_OP_425J2_127_3477_n1437) );
  FADDX1_HVT DP_OP_425J2_127_3477_U875 ( .A(DP_OP_425J2_127_3477_n1525), .B(
        DP_OP_425J2_127_3477_n1509), .CI(DP_OP_425J2_127_3477_n1610), .CO(
        DP_OP_425J2_127_3477_n1434), .S(DP_OP_425J2_127_3477_n1435) );
  FADDX1_HVT DP_OP_425J2_127_3477_U874 ( .A(DP_OP_425J2_127_3477_n1523), .B(
        DP_OP_425J2_127_3477_n1511), .CI(DP_OP_425J2_127_3477_n1513), .CO(
        DP_OP_425J2_127_3477_n1432), .S(DP_OP_425J2_127_3477_n1433) );
  FADDX1_HVT DP_OP_425J2_127_3477_U873 ( .A(DP_OP_425J2_127_3477_n1519), .B(
        DP_OP_425J2_127_3477_n1517), .CI(DP_OP_425J2_127_3477_n1521), .CO(
        DP_OP_425J2_127_3477_n1430), .S(DP_OP_425J2_127_3477_n1431) );
  FADDX1_HVT DP_OP_425J2_127_3477_U872 ( .A(DP_OP_425J2_127_3477_n1515), .B(
        DP_OP_425J2_127_3477_n1495), .CI(DP_OP_425J2_127_3477_n1499), .CO(
        DP_OP_425J2_127_3477_n1428), .S(DP_OP_425J2_127_3477_n1429) );
  FADDX1_HVT DP_OP_425J2_127_3477_U871 ( .A(DP_OP_425J2_127_3477_n1497), .B(
        DP_OP_425J2_127_3477_n1505), .CI(DP_OP_425J2_127_3477_n1503), .CO(
        DP_OP_425J2_127_3477_n1426), .S(DP_OP_425J2_127_3477_n1427) );
  FADDX1_HVT DP_OP_425J2_127_3477_U870 ( .A(DP_OP_425J2_127_3477_n1507), .B(
        DP_OP_425J2_127_3477_n1485), .CI(DP_OP_425J2_127_3477_n1479), .CO(
        DP_OP_425J2_127_3477_n1424), .S(DP_OP_425J2_127_3477_n1425) );
  FADDX1_HVT DP_OP_425J2_127_3477_U869 ( .A(DP_OP_425J2_127_3477_n1487), .B(
        DP_OP_425J2_127_3477_n1483), .CI(DP_OP_425J2_127_3477_n1477), .CO(
        DP_OP_425J2_127_3477_n1422), .S(DP_OP_425J2_127_3477_n1423) );
  FADDX1_HVT DP_OP_425J2_127_3477_U868 ( .A(DP_OP_425J2_127_3477_n1489), .B(
        DP_OP_425J2_127_3477_n1463), .CI(DP_OP_425J2_127_3477_n1461), .CO(
        DP_OP_425J2_127_3477_n1420), .S(DP_OP_425J2_127_3477_n1421) );
  FADDX1_HVT DP_OP_425J2_127_3477_U867 ( .A(DP_OP_425J2_127_3477_n1475), .B(
        DP_OP_425J2_127_3477_n1471), .CI(DP_OP_425J2_127_3477_n1473), .CO(
        DP_OP_425J2_127_3477_n1418), .S(DP_OP_425J2_127_3477_n1419) );
  FADDX1_HVT DP_OP_425J2_127_3477_U866 ( .A(DP_OP_425J2_127_3477_n1481), .B(
        DP_OP_425J2_127_3477_n1459), .CI(DP_OP_425J2_127_3477_n1467), .CO(
        DP_OP_425J2_127_3477_n1416), .S(DP_OP_425J2_127_3477_n1417) );
  FADDX1_HVT DP_OP_425J2_127_3477_U865 ( .A(DP_OP_425J2_127_3477_n1469), .B(
        DP_OP_425J2_127_3477_n1493), .CI(DP_OP_425J2_127_3477_n1501), .CO(
        DP_OP_425J2_127_3477_n1414), .S(DP_OP_425J2_127_3477_n1415) );
  FADDX1_HVT DP_OP_425J2_127_3477_U864 ( .A(DP_OP_425J2_127_3477_n1465), .B(
        DP_OP_425J2_127_3477_n1491), .CI(DP_OP_425J2_127_3477_n1608), .CO(
        DP_OP_425J2_127_3477_n1412), .S(DP_OP_425J2_127_3477_n1413) );
  FADDX1_HVT DP_OP_425J2_127_3477_U863 ( .A(DP_OP_425J2_127_3477_n1606), .B(
        DP_OP_425J2_127_3477_n1604), .CI(DP_OP_425J2_127_3477_n1602), .CO(
        DP_OP_425J2_127_3477_n1410), .S(DP_OP_425J2_127_3477_n1411) );
  FADDX1_HVT DP_OP_425J2_127_3477_U862 ( .A(DP_OP_425J2_127_3477_n1594), .B(
        DP_OP_425J2_127_3477_n1600), .CI(DP_OP_425J2_127_3477_n1596), .CO(
        DP_OP_425J2_127_3477_n1408), .S(DP_OP_425J2_127_3477_n1409) );
  FADDX1_HVT DP_OP_425J2_127_3477_U861 ( .A(DP_OP_425J2_127_3477_n1598), .B(
        DP_OP_425J2_127_3477_n1592), .CI(DP_OP_425J2_127_3477_n1453), .CO(
        DP_OP_425J2_127_3477_n1406), .S(DP_OP_425J2_127_3477_n1407) );
  FADDX1_HVT DP_OP_425J2_127_3477_U860 ( .A(DP_OP_425J2_127_3477_n1455), .B(
        DP_OP_425J2_127_3477_n1590), .CI(DP_OP_425J2_127_3477_n1586), .CO(
        DP_OP_425J2_127_3477_n1404), .S(DP_OP_425J2_127_3477_n1405) );
  FADDX1_HVT DP_OP_425J2_127_3477_U859 ( .A(DP_OP_425J2_127_3477_n1457), .B(
        DP_OP_425J2_127_3477_n1588), .CI(DP_OP_425J2_127_3477_n1584), .CO(
        DP_OP_425J2_127_3477_n1402), .S(DP_OP_425J2_127_3477_n1403) );
  FADDX1_HVT DP_OP_425J2_127_3477_U858 ( .A(DP_OP_425J2_127_3477_n1574), .B(
        DP_OP_425J2_127_3477_n1437), .CI(DP_OP_425J2_127_3477_n1449), .CO(
        DP_OP_425J2_127_3477_n1400), .S(DP_OP_425J2_127_3477_n1401) );
  FADDX1_HVT DP_OP_425J2_127_3477_U857 ( .A(DP_OP_425J2_127_3477_n1582), .B(
        DP_OP_425J2_127_3477_n1451), .CI(DP_OP_425J2_127_3477_n1447), .CO(
        DP_OP_425J2_127_3477_n1398), .S(DP_OP_425J2_127_3477_n1399) );
  FADDX1_HVT DP_OP_425J2_127_3477_U856 ( .A(DP_OP_425J2_127_3477_n1580), .B(
        DP_OP_425J2_127_3477_n1439), .CI(DP_OP_425J2_127_3477_n1441), .CO(
        DP_OP_425J2_127_3477_n1396), .S(DP_OP_425J2_127_3477_n1397) );
  FADDX1_HVT DP_OP_425J2_127_3477_U855 ( .A(DP_OP_425J2_127_3477_n1578), .B(
        DP_OP_425J2_127_3477_n1445), .CI(DP_OP_425J2_127_3477_n1443), .CO(
        DP_OP_425J2_127_3477_n1394), .S(DP_OP_425J2_127_3477_n1395) );
  FADDX1_HVT DP_OP_425J2_127_3477_U854 ( .A(DP_OP_425J2_127_3477_n1576), .B(
        DP_OP_425J2_127_3477_n1572), .CI(DP_OP_425J2_127_3477_n1433), .CO(
        DP_OP_425J2_127_3477_n1392), .S(DP_OP_425J2_127_3477_n1393) );
  FADDX1_HVT DP_OP_425J2_127_3477_U853 ( .A(DP_OP_425J2_127_3477_n1435), .B(
        DP_OP_425J2_127_3477_n1431), .CI(DP_OP_425J2_127_3477_n1429), .CO(
        DP_OP_425J2_127_3477_n1390), .S(DP_OP_425J2_127_3477_n1391) );
  FADDX1_HVT DP_OP_425J2_127_3477_U852 ( .A(DP_OP_425J2_127_3477_n1570), .B(
        DP_OP_425J2_127_3477_n1421), .CI(DP_OP_425J2_127_3477_n1419), .CO(
        DP_OP_425J2_127_3477_n1388), .S(DP_OP_425J2_127_3477_n1389) );
  FADDX1_HVT DP_OP_425J2_127_3477_U851 ( .A(DP_OP_425J2_127_3477_n1425), .B(
        DP_OP_425J2_127_3477_n1415), .CI(DP_OP_425J2_127_3477_n1417), .CO(
        DP_OP_425J2_127_3477_n1386), .S(DP_OP_425J2_127_3477_n1387) );
  FADDX1_HVT DP_OP_425J2_127_3477_U850 ( .A(DP_OP_425J2_127_3477_n1423), .B(
        DP_OP_425J2_127_3477_n1427), .CI(DP_OP_425J2_127_3477_n1568), .CO(
        DP_OP_425J2_127_3477_n1384), .S(DP_OP_425J2_127_3477_n1385) );
  FADDX1_HVT DP_OP_425J2_127_3477_U849 ( .A(DP_OP_425J2_127_3477_n1566), .B(
        DP_OP_425J2_127_3477_n1413), .CI(DP_OP_425J2_127_3477_n1564), .CO(
        DP_OP_425J2_127_3477_n1382), .S(DP_OP_425J2_127_3477_n1383) );
  FADDX1_HVT DP_OP_425J2_127_3477_U848 ( .A(DP_OP_425J2_127_3477_n1562), .B(
        DP_OP_425J2_127_3477_n1409), .CI(DP_OP_425J2_127_3477_n1411), .CO(
        DP_OP_425J2_127_3477_n1380), .S(DP_OP_425J2_127_3477_n1381) );
  FADDX1_HVT DP_OP_425J2_127_3477_U847 ( .A(DP_OP_425J2_127_3477_n1560), .B(
        DP_OP_425J2_127_3477_n1556), .CI(DP_OP_425J2_127_3477_n1558), .CO(
        DP_OP_425J2_127_3477_n1378), .S(DP_OP_425J2_127_3477_n1379) );
  FADDX1_HVT DP_OP_425J2_127_3477_U846 ( .A(DP_OP_425J2_127_3477_n1407), .B(
        DP_OP_425J2_127_3477_n1554), .CI(DP_OP_425J2_127_3477_n1552), .CO(
        DP_OP_425J2_127_3477_n1376), .S(DP_OP_425J2_127_3477_n1377) );
  FADDX1_HVT DP_OP_425J2_127_3477_U845 ( .A(DP_OP_425J2_127_3477_n1405), .B(
        DP_OP_425J2_127_3477_n1403), .CI(DP_OP_425J2_127_3477_n1399), .CO(
        DP_OP_425J2_127_3477_n1374), .S(DP_OP_425J2_127_3477_n1375) );
  FADDX1_HVT DP_OP_425J2_127_3477_U844 ( .A(DP_OP_425J2_127_3477_n1401), .B(
        DP_OP_425J2_127_3477_n1397), .CI(DP_OP_425J2_127_3477_n1393), .CO(
        DP_OP_425J2_127_3477_n1372), .S(DP_OP_425J2_127_3477_n1373) );
  FADDX1_HVT DP_OP_425J2_127_3477_U843 ( .A(DP_OP_425J2_127_3477_n1550), .B(
        DP_OP_425J2_127_3477_n1395), .CI(DP_OP_425J2_127_3477_n1548), .CO(
        DP_OP_425J2_127_3477_n1370), .S(DP_OP_425J2_127_3477_n1371) );
  FADDX1_HVT DP_OP_425J2_127_3477_U842 ( .A(DP_OP_425J2_127_3477_n1391), .B(
        DP_OP_425J2_127_3477_n1389), .CI(DP_OP_425J2_127_3477_n1387), .CO(
        DP_OP_425J2_127_3477_n1368), .S(DP_OP_425J2_127_3477_n1369) );
  FADDX1_HVT DP_OP_425J2_127_3477_U841 ( .A(DP_OP_425J2_127_3477_n1546), .B(
        DP_OP_425J2_127_3477_n1385), .CI(DP_OP_425J2_127_3477_n1544), .CO(
        DP_OP_425J2_127_3477_n1366), .S(DP_OP_425J2_127_3477_n1367) );
  FADDX1_HVT DP_OP_425J2_127_3477_U840 ( .A(DP_OP_425J2_127_3477_n1383), .B(
        DP_OP_425J2_127_3477_n1542), .CI(DP_OP_425J2_127_3477_n1540), .CO(
        DP_OP_425J2_127_3477_n1364), .S(DP_OP_425J2_127_3477_n1365) );
  FADDX1_HVT DP_OP_425J2_127_3477_U839 ( .A(DP_OP_425J2_127_3477_n1379), .B(
        DP_OP_425J2_127_3477_n1381), .CI(DP_OP_425J2_127_3477_n1538), .CO(
        DP_OP_425J2_127_3477_n1362), .S(DP_OP_425J2_127_3477_n1363) );
  FADDX1_HVT DP_OP_425J2_127_3477_U838 ( .A(DP_OP_425J2_127_3477_n1377), .B(
        DP_OP_425J2_127_3477_n1375), .CI(DP_OP_425J2_127_3477_n1536), .CO(
        DP_OP_425J2_127_3477_n1360), .S(DP_OP_425J2_127_3477_n1361) );
  FADDX1_HVT DP_OP_425J2_127_3477_U837 ( .A(DP_OP_425J2_127_3477_n1371), .B(
        DP_OP_425J2_127_3477_n1373), .CI(DP_OP_425J2_127_3477_n1534), .CO(
        DP_OP_425J2_127_3477_n1358), .S(DP_OP_425J2_127_3477_n1359) );
  FADDX1_HVT DP_OP_425J2_127_3477_U836 ( .A(DP_OP_425J2_127_3477_n1369), .B(
        DP_OP_425J2_127_3477_n1367), .CI(DP_OP_425J2_127_3477_n1532), .CO(
        DP_OP_425J2_127_3477_n1356), .S(DP_OP_425J2_127_3477_n1357) );
  FADDX1_HVT DP_OP_425J2_127_3477_U835 ( .A(DP_OP_425J2_127_3477_n1365), .B(
        DP_OP_425J2_127_3477_n1530), .CI(DP_OP_425J2_127_3477_n1363), .CO(
        DP_OP_425J2_127_3477_n1354), .S(DP_OP_425J2_127_3477_n1355) );
  FADDX1_HVT DP_OP_425J2_127_3477_U834 ( .A(DP_OP_425J2_127_3477_n1361), .B(
        DP_OP_425J2_127_3477_n1528), .CI(DP_OP_425J2_127_3477_n1359), .CO(
        DP_OP_425J2_127_3477_n1352), .S(DP_OP_425J2_127_3477_n1353) );
  FADDX1_HVT DP_OP_425J2_127_3477_U833 ( .A(DP_OP_425J2_127_3477_n1357), .B(
        DP_OP_425J2_127_3477_n1526), .CI(DP_OP_425J2_127_3477_n1355), .CO(
        DP_OP_425J2_127_3477_n1350), .S(DP_OP_425J2_127_3477_n1351) );
  HADDX1_HVT DP_OP_425J2_127_3477_U832 ( .A0(DP_OP_425J2_127_3477_n2980), .B0(
        DP_OP_425J2_127_3477_n1925), .C1(DP_OP_425J2_127_3477_n1348), .SO(
        DP_OP_425J2_127_3477_n1349) );
  FADDX1_HVT DP_OP_425J2_127_3477_U831 ( .A(DP_OP_425J2_127_3477_n2453), .B(
        DP_OP_425J2_127_3477_n2365), .CI(DP_OP_425J2_127_3477_n1881), .CO(
        DP_OP_425J2_127_3477_n1346), .S(DP_OP_425J2_127_3477_n1347) );
  FADDX1_HVT DP_OP_425J2_127_3477_U830 ( .A(DP_OP_425J2_127_3477_n2497), .B(
        DP_OP_425J2_127_3477_n2277), .CI(DP_OP_425J2_127_3477_n2321), .CO(
        DP_OP_425J2_127_3477_n1344), .S(DP_OP_425J2_127_3477_n1345) );
  FADDX1_HVT DP_OP_425J2_127_3477_U829 ( .A(DP_OP_425J2_127_3477_n2805), .B(
        DP_OP_425J2_127_3477_n1969), .CI(DP_OP_425J2_127_3477_n2057), .CO(
        DP_OP_425J2_127_3477_n1342), .S(DP_OP_425J2_127_3477_n1343) );
  FADDX1_HVT DP_OP_425J2_127_3477_U828 ( .A(DP_OP_425J2_127_3477_n2541), .B(
        DP_OP_425J2_127_3477_n2101), .CI(DP_OP_425J2_127_3477_n2629), .CO(
        DP_OP_425J2_127_3477_n1340), .S(DP_OP_425J2_127_3477_n1341) );
  FADDX1_HVT DP_OP_425J2_127_3477_U827 ( .A(DP_OP_425J2_127_3477_n2013), .B(
        DP_OP_425J2_127_3477_n2849), .CI(DP_OP_425J2_127_3477_n2145), .CO(
        DP_OP_425J2_127_3477_n1338), .S(DP_OP_425J2_127_3477_n1339) );
  FADDX1_HVT DP_OP_425J2_127_3477_U826 ( .A(DP_OP_425J2_127_3477_n2409), .B(
        DP_OP_425J2_127_3477_n2893), .CI(DP_OP_425J2_127_3477_n2717), .CO(
        DP_OP_425J2_127_3477_n1336), .S(DP_OP_425J2_127_3477_n1337) );
  FADDX1_HVT DP_OP_425J2_127_3477_U825 ( .A(DP_OP_425J2_127_3477_n2233), .B(
        DP_OP_425J2_127_3477_n2189), .CI(DP_OP_425J2_127_3477_n2673), .CO(
        DP_OP_425J2_127_3477_n1334), .S(DP_OP_425J2_127_3477_n1335) );
  FADDX1_HVT DP_OP_425J2_127_3477_U824 ( .A(DP_OP_425J2_127_3477_n2937), .B(
        DP_OP_425J2_127_3477_n2585), .CI(DP_OP_425J2_127_3477_n2761), .CO(
        DP_OP_425J2_127_3477_n1332), .S(DP_OP_425J2_127_3477_n1333) );
  FADDX1_HVT DP_OP_425J2_127_3477_U823 ( .A(DP_OP_425J2_127_3477_n2379), .B(
        DP_OP_425J2_127_3477_n3000), .CI(DP_OP_425J2_127_3477_n1932), .CO(
        DP_OP_425J2_127_3477_n1330), .S(DP_OP_425J2_127_3477_n1331) );
  FADDX1_HVT DP_OP_425J2_127_3477_U822 ( .A(DP_OP_425J2_127_3477_n2372), .B(
        DP_OP_425J2_127_3477_n1939), .CI(DP_OP_425J2_127_3477_n1946), .CO(
        DP_OP_425J2_127_3477_n1328), .S(DP_OP_425J2_127_3477_n1329) );
  FADDX1_HVT DP_OP_425J2_127_3477_U821 ( .A(DP_OP_425J2_127_3477_n2386), .B(
        DP_OP_425J2_127_3477_n1976), .CI(DP_OP_425J2_127_3477_n2993), .CO(
        DP_OP_425J2_127_3477_n1326), .S(DP_OP_425J2_127_3477_n1327) );
  FADDX1_HVT DP_OP_425J2_127_3477_U820 ( .A(DP_OP_425J2_127_3477_n2342), .B(
        DP_OP_425J2_127_3477_n2986), .CI(DP_OP_425J2_127_3477_n2958), .CO(
        DP_OP_425J2_127_3477_n1324), .S(DP_OP_425J2_127_3477_n1325) );
  FADDX1_HVT DP_OP_425J2_127_3477_U819 ( .A(DP_OP_425J2_127_3477_n2335), .B(
        DP_OP_425J2_127_3477_n2951), .CI(DP_OP_425J2_127_3477_n2944), .CO(
        DP_OP_425J2_127_3477_n1322), .S(DP_OP_425J2_127_3477_n1323) );
  FADDX1_HVT DP_OP_425J2_127_3477_U818 ( .A(DP_OP_425J2_127_3477_n2298), .B(
        DP_OP_425J2_127_3477_n2914), .CI(DP_OP_425J2_127_3477_n2907), .CO(
        DP_OP_425J2_127_3477_n1320), .S(DP_OP_425J2_127_3477_n1321) );
  FADDX1_HVT DP_OP_425J2_127_3477_U817 ( .A(DP_OP_425J2_127_3477_n2291), .B(
        DP_OP_425J2_127_3477_n1983), .CI(DP_OP_425J2_127_3477_n2900), .CO(
        DP_OP_425J2_127_3477_n1318), .S(DP_OP_425J2_127_3477_n1319) );
  FADDX1_HVT DP_OP_425J2_127_3477_U816 ( .A(DP_OP_425J2_127_3477_n2284), .B(
        DP_OP_425J2_127_3477_n2870), .CI(DP_OP_425J2_127_3477_n2863), .CO(
        DP_OP_425J2_127_3477_n1316), .S(DP_OP_425J2_127_3477_n1317) );
  FADDX1_HVT DP_OP_425J2_127_3477_U815 ( .A(DP_OP_425J2_127_3477_n2254), .B(
        DP_OP_425J2_127_3477_n2856), .CI(DP_OP_425J2_127_3477_n1990), .CO(
        DP_OP_425J2_127_3477_n1314), .S(DP_OP_425J2_127_3477_n1315) );
  FADDX1_HVT DP_OP_425J2_127_3477_U814 ( .A(DP_OP_425J2_127_3477_n2247), .B(
        DP_OP_425J2_127_3477_n2020), .CI(DP_OP_425J2_127_3477_n2027), .CO(
        DP_OP_425J2_127_3477_n1312), .S(DP_OP_425J2_127_3477_n1313) );
  FADDX1_HVT DP_OP_425J2_127_3477_U813 ( .A(DP_OP_425J2_127_3477_n2328), .B(
        DP_OP_425J2_127_3477_n2034), .CI(DP_OP_425J2_127_3477_n2826), .CO(
        DP_OP_425J2_127_3477_n1310), .S(DP_OP_425J2_127_3477_n1311) );
  FADDX1_HVT DP_OP_425J2_127_3477_U812 ( .A(DP_OP_425J2_127_3477_n2416), .B(
        DP_OP_425J2_127_3477_n2819), .CI(DP_OP_425J2_127_3477_n2064), .CO(
        DP_OP_425J2_127_3477_n1308), .S(DP_OP_425J2_127_3477_n1309) );
  FADDX1_HVT DP_OP_425J2_127_3477_U811 ( .A(DP_OP_425J2_127_3477_n2812), .B(
        DP_OP_425J2_127_3477_n2071), .CI(DP_OP_425J2_127_3477_n2078), .CO(
        DP_OP_425J2_127_3477_n1306), .S(DP_OP_425J2_127_3477_n1307) );
  FADDX1_HVT DP_OP_425J2_127_3477_U810 ( .A(DP_OP_425J2_127_3477_n2782), .B(
        DP_OP_425J2_127_3477_n2108), .CI(DP_OP_425J2_127_3477_n2115), .CO(
        DP_OP_425J2_127_3477_n1304), .S(DP_OP_425J2_127_3477_n1305) );
  FADDX1_HVT DP_OP_425J2_127_3477_U809 ( .A(DP_OP_425J2_127_3477_n2775), .B(
        DP_OP_425J2_127_3477_n2122), .CI(DP_OP_425J2_127_3477_n2152), .CO(
        DP_OP_425J2_127_3477_n1302), .S(DP_OP_425J2_127_3477_n1303) );
  FADDX1_HVT DP_OP_425J2_127_3477_U808 ( .A(DP_OP_425J2_127_3477_n2768), .B(
        DP_OP_425J2_127_3477_n2159), .CI(DP_OP_425J2_127_3477_n2166), .CO(
        DP_OP_425J2_127_3477_n1300), .S(DP_OP_425J2_127_3477_n1301) );
  FADDX1_HVT DP_OP_425J2_127_3477_U807 ( .A(DP_OP_425J2_127_3477_n2738), .B(
        DP_OP_425J2_127_3477_n2196), .CI(DP_OP_425J2_127_3477_n2203), .CO(
        DP_OP_425J2_127_3477_n1298), .S(DP_OP_425J2_127_3477_n1299) );
  FADDX1_HVT DP_OP_425J2_127_3477_U806 ( .A(DP_OP_425J2_127_3477_n2731), .B(
        DP_OP_425J2_127_3477_n2210), .CI(DP_OP_425J2_127_3477_n2240), .CO(
        DP_OP_425J2_127_3477_n1296), .S(DP_OP_425J2_127_3477_n1297) );
  FADDX1_HVT DP_OP_425J2_127_3477_U805 ( .A(DP_OP_425J2_127_3477_n2724), .B(
        DP_OP_425J2_127_3477_n2423), .CI(DP_OP_425J2_127_3477_n2430), .CO(
        DP_OP_425J2_127_3477_n1294), .S(DP_OP_425J2_127_3477_n1295) );
  FADDX1_HVT DP_OP_425J2_127_3477_U804 ( .A(DP_OP_425J2_127_3477_n2694), .B(
        DP_OP_425J2_127_3477_n2460), .CI(DP_OP_425J2_127_3477_n2467), .CO(
        DP_OP_425J2_127_3477_n1292), .S(DP_OP_425J2_127_3477_n1293) );
  FADDX1_HVT DP_OP_425J2_127_3477_U803 ( .A(DP_OP_425J2_127_3477_n2687), .B(
        DP_OP_425J2_127_3477_n2474), .CI(DP_OP_425J2_127_3477_n2504), .CO(
        DP_OP_425J2_127_3477_n1290), .S(DP_OP_425J2_127_3477_n1291) );
  FADDX1_HVT DP_OP_425J2_127_3477_U802 ( .A(DP_OP_425J2_127_3477_n2680), .B(
        DP_OP_425J2_127_3477_n2511), .CI(DP_OP_425J2_127_3477_n2518), .CO(
        DP_OP_425J2_127_3477_n1288), .S(DP_OP_425J2_127_3477_n1289) );
  FADDX1_HVT DP_OP_425J2_127_3477_U801 ( .A(DP_OP_425J2_127_3477_n2650), .B(
        DP_OP_425J2_127_3477_n2643), .CI(DP_OP_425J2_127_3477_n2636), .CO(
        DP_OP_425J2_127_3477_n1286), .S(DP_OP_425J2_127_3477_n1287) );
  FADDX1_HVT DP_OP_425J2_127_3477_U800 ( .A(DP_OP_425J2_127_3477_n2592), .B(
        DP_OP_425J2_127_3477_n2606), .CI(DP_OP_425J2_127_3477_n2548), .CO(
        DP_OP_425J2_127_3477_n1284), .S(DP_OP_425J2_127_3477_n1285) );
  FADDX1_HVT DP_OP_425J2_127_3477_U799 ( .A(DP_OP_425J2_127_3477_n2555), .B(
        DP_OP_425J2_127_3477_n2562), .CI(DP_OP_425J2_127_3477_n2599), .CO(
        DP_OP_425J2_127_3477_n1282), .S(DP_OP_425J2_127_3477_n1283) );
  FADDX1_HVT DP_OP_425J2_127_3477_U798 ( .A(DP_OP_425J2_127_3477_n1349), .B(
        DP_OP_425J2_127_3477_n1524), .CI(DP_OP_425J2_127_3477_n1514), .CO(
        DP_OP_425J2_127_3477_n1280), .S(DP_OP_425J2_127_3477_n1281) );
  FADDX1_HVT DP_OP_425J2_127_3477_U797 ( .A(DP_OP_425J2_127_3477_n1522), .B(
        DP_OP_425J2_127_3477_n1520), .CI(DP_OP_425J2_127_3477_n1518), .CO(
        DP_OP_425J2_127_3477_n1278), .S(DP_OP_425J2_127_3477_n1279) );
  FADDX1_HVT DP_OP_425J2_127_3477_U796 ( .A(DP_OP_425J2_127_3477_n1516), .B(
        DP_OP_425J2_127_3477_n1512), .CI(DP_OP_425J2_127_3477_n1508), .CO(
        DP_OP_425J2_127_3477_n1276), .S(DP_OP_425J2_127_3477_n1277) );
  FADDX1_HVT DP_OP_425J2_127_3477_U795 ( .A(DP_OP_425J2_127_3477_n1510), .B(
        DP_OP_425J2_127_3477_n1484), .CI(DP_OP_425J2_127_3477_n1482), .CO(
        DP_OP_425J2_127_3477_n1274), .S(DP_OP_425J2_127_3477_n1275) );
  FADDX1_HVT DP_OP_425J2_127_3477_U794 ( .A(DP_OP_425J2_127_3477_n1486), .B(
        DP_OP_425J2_127_3477_n1458), .CI(DP_OP_425J2_127_3477_n1506), .CO(
        DP_OP_425J2_127_3477_n1272), .S(DP_OP_425J2_127_3477_n1273) );
  FADDX1_HVT DP_OP_425J2_127_3477_U793 ( .A(DP_OP_425J2_127_3477_n1478), .B(
        DP_OP_425J2_127_3477_n1504), .CI(DP_OP_425J2_127_3477_n1502), .CO(
        DP_OP_425J2_127_3477_n1270), .S(DP_OP_425J2_127_3477_n1271) );
  FADDX1_HVT DP_OP_425J2_127_3477_U792 ( .A(DP_OP_425J2_127_3477_n1474), .B(
        DP_OP_425J2_127_3477_n1500), .CI(DP_OP_425J2_127_3477_n1498), .CO(
        DP_OP_425J2_127_3477_n1268), .S(DP_OP_425J2_127_3477_n1269) );
  FADDX1_HVT DP_OP_425J2_127_3477_U791 ( .A(DP_OP_425J2_127_3477_n1468), .B(
        DP_OP_425J2_127_3477_n1460), .CI(DP_OP_425J2_127_3477_n1462), .CO(
        DP_OP_425J2_127_3477_n1266), .S(DP_OP_425J2_127_3477_n1267) );
  FADDX1_HVT DP_OP_425J2_127_3477_U790 ( .A(DP_OP_425J2_127_3477_n1466), .B(
        DP_OP_425J2_127_3477_n1496), .CI(DP_OP_425J2_127_3477_n1494), .CO(
        DP_OP_425J2_127_3477_n1264), .S(DP_OP_425J2_127_3477_n1265) );
  FADDX1_HVT DP_OP_425J2_127_3477_U789 ( .A(DP_OP_425J2_127_3477_n1476), .B(
        DP_OP_425J2_127_3477_n1492), .CI(DP_OP_425J2_127_3477_n1464), .CO(
        DP_OP_425J2_127_3477_n1262), .S(DP_OP_425J2_127_3477_n1263) );
  FADDX1_HVT DP_OP_425J2_127_3477_U788 ( .A(DP_OP_425J2_127_3477_n1472), .B(
        DP_OP_425J2_127_3477_n1490), .CI(DP_OP_425J2_127_3477_n1488), .CO(
        DP_OP_425J2_127_3477_n1260), .S(DP_OP_425J2_127_3477_n1261) );
  FADDX1_HVT DP_OP_425J2_127_3477_U787 ( .A(DP_OP_425J2_127_3477_n1470), .B(
        DP_OP_425J2_127_3477_n1480), .CI(DP_OP_425J2_127_3477_n1339), .CO(
        DP_OP_425J2_127_3477_n1258), .S(DP_OP_425J2_127_3477_n1259) );
  FADDX1_HVT DP_OP_425J2_127_3477_U786 ( .A(DP_OP_425J2_127_3477_n1341), .B(
        DP_OP_425J2_127_3477_n1333), .CI(DP_OP_425J2_127_3477_n1335), .CO(
        DP_OP_425J2_127_3477_n1256), .S(DP_OP_425J2_127_3477_n1257) );
  FADDX1_HVT DP_OP_425J2_127_3477_U785 ( .A(DP_OP_425J2_127_3477_n1345), .B(
        DP_OP_425J2_127_3477_n1343), .CI(DP_OP_425J2_127_3477_n1347), .CO(
        DP_OP_425J2_127_3477_n1254), .S(DP_OP_425J2_127_3477_n1255) );
  FADDX1_HVT DP_OP_425J2_127_3477_U784 ( .A(DP_OP_425J2_127_3477_n1337), .B(
        DP_OP_425J2_127_3477_n1289), .CI(DP_OP_425J2_127_3477_n1287), .CO(
        DP_OP_425J2_127_3477_n1252), .S(DP_OP_425J2_127_3477_n1253) );
  FADDX1_HVT DP_OP_425J2_127_3477_U783 ( .A(DP_OP_425J2_127_3477_n1283), .B(
        DP_OP_425J2_127_3477_n1331), .CI(DP_OP_425J2_127_3477_n1329), .CO(
        DP_OP_425J2_127_3477_n1250), .S(DP_OP_425J2_127_3477_n1251) );
  FADDX1_HVT DP_OP_425J2_127_3477_U782 ( .A(DP_OP_425J2_127_3477_n1319), .B(
        DP_OP_425J2_127_3477_n1309), .CI(DP_OP_425J2_127_3477_n1315), .CO(
        DP_OP_425J2_127_3477_n1248), .S(DP_OP_425J2_127_3477_n1249) );
  FADDX1_HVT DP_OP_425J2_127_3477_U781 ( .A(DP_OP_425J2_127_3477_n1313), .B(
        DP_OP_425J2_127_3477_n1311), .CI(DP_OP_425J2_127_3477_n1295), .CO(
        DP_OP_425J2_127_3477_n1246), .S(DP_OP_425J2_127_3477_n1247) );
  FADDX1_HVT DP_OP_425J2_127_3477_U780 ( .A(DP_OP_425J2_127_3477_n1317), .B(
        DP_OP_425J2_127_3477_n1291), .CI(DP_OP_425J2_127_3477_n1285), .CO(
        DP_OP_425J2_127_3477_n1244), .S(DP_OP_425J2_127_3477_n1245) );
  FADDX1_HVT DP_OP_425J2_127_3477_U779 ( .A(DP_OP_425J2_127_3477_n1321), .B(
        DP_OP_425J2_127_3477_n1303), .CI(DP_OP_425J2_127_3477_n1305), .CO(
        DP_OP_425J2_127_3477_n1242), .S(DP_OP_425J2_127_3477_n1243) );
  FADDX1_HVT DP_OP_425J2_127_3477_U778 ( .A(DP_OP_425J2_127_3477_n1301), .B(
        DP_OP_425J2_127_3477_n1299), .CI(DP_OP_425J2_127_3477_n1293), .CO(
        DP_OP_425J2_127_3477_n1240), .S(DP_OP_425J2_127_3477_n1241) );
  FADDX1_HVT DP_OP_425J2_127_3477_U777 ( .A(DP_OP_425J2_127_3477_n1297), .B(
        DP_OP_425J2_127_3477_n1327), .CI(DP_OP_425J2_127_3477_n1323), .CO(
        DP_OP_425J2_127_3477_n1238), .S(DP_OP_425J2_127_3477_n1239) );
  FADDX1_HVT DP_OP_425J2_127_3477_U776 ( .A(DP_OP_425J2_127_3477_n1325), .B(
        DP_OP_425J2_127_3477_n1307), .CI(DP_OP_425J2_127_3477_n1456), .CO(
        DP_OP_425J2_127_3477_n1236), .S(DP_OP_425J2_127_3477_n1237) );
  FADDX1_HVT DP_OP_425J2_127_3477_U775 ( .A(DP_OP_425J2_127_3477_n1454), .B(
        DP_OP_425J2_127_3477_n1452), .CI(DP_OP_425J2_127_3477_n1450), .CO(
        DP_OP_425J2_127_3477_n1234), .S(DP_OP_425J2_127_3477_n1235) );
  FADDX1_HVT DP_OP_425J2_127_3477_U774 ( .A(DP_OP_425J2_127_3477_n1448), .B(
        DP_OP_425J2_127_3477_n1436), .CI(DP_OP_425J2_127_3477_n1438), .CO(
        DP_OP_425J2_127_3477_n1232), .S(DP_OP_425J2_127_3477_n1233) );
  FADDX1_HVT DP_OP_425J2_127_3477_U773 ( .A(DP_OP_425J2_127_3477_n1442), .B(
        DP_OP_425J2_127_3477_n1446), .CI(DP_OP_425J2_127_3477_n1440), .CO(
        DP_OP_425J2_127_3477_n1230), .S(DP_OP_425J2_127_3477_n1231) );
  FADDX1_HVT DP_OP_425J2_127_3477_U772 ( .A(DP_OP_425J2_127_3477_n1444), .B(
        DP_OP_425J2_127_3477_n1281), .CI(DP_OP_425J2_127_3477_n1434), .CO(
        DP_OP_425J2_127_3477_n1228), .S(DP_OP_425J2_127_3477_n1229) );
  FADDX1_HVT DP_OP_425J2_127_3477_U771 ( .A(DP_OP_425J2_127_3477_n1279), .B(
        DP_OP_425J2_127_3477_n1277), .CI(DP_OP_425J2_127_3477_n1275), .CO(
        DP_OP_425J2_127_3477_n1226), .S(DP_OP_425J2_127_3477_n1227) );
  FADDX1_HVT DP_OP_425J2_127_3477_U770 ( .A(DP_OP_425J2_127_3477_n1432), .B(
        DP_OP_425J2_127_3477_n1430), .CI(DP_OP_425J2_127_3477_n1428), .CO(
        DP_OP_425J2_127_3477_n1224), .S(DP_OP_425J2_127_3477_n1225) );
  FADDX1_HVT DP_OP_425J2_127_3477_U769 ( .A(DP_OP_425J2_127_3477_n1416), .B(
        DP_OP_425J2_127_3477_n1261), .CI(DP_OP_425J2_127_3477_n1259), .CO(
        DP_OP_425J2_127_3477_n1222), .S(DP_OP_425J2_127_3477_n1223) );
  FADDX1_HVT DP_OP_425J2_127_3477_U768 ( .A(DP_OP_425J2_127_3477_n1426), .B(
        DP_OP_425J2_127_3477_n1271), .CI(DP_OP_425J2_127_3477_n1273), .CO(
        DP_OP_425J2_127_3477_n1220), .S(DP_OP_425J2_127_3477_n1221) );
  FADDX1_HVT DP_OP_425J2_127_3477_U767 ( .A(DP_OP_425J2_127_3477_n1424), .B(
        DP_OP_425J2_127_3477_n1267), .CI(DP_OP_425J2_127_3477_n1263), .CO(
        DP_OP_425J2_127_3477_n1218), .S(DP_OP_425J2_127_3477_n1219) );
  FADDX1_HVT DP_OP_425J2_127_3477_U766 ( .A(DP_OP_425J2_127_3477_n1422), .B(
        DP_OP_425J2_127_3477_n1269), .CI(DP_OP_425J2_127_3477_n1265), .CO(
        DP_OP_425J2_127_3477_n1216), .S(DP_OP_425J2_127_3477_n1217) );
  FADDX1_HVT DP_OP_425J2_127_3477_U765 ( .A(DP_OP_425J2_127_3477_n1420), .B(
        DP_OP_425J2_127_3477_n1414), .CI(DP_OP_425J2_127_3477_n1418), .CO(
        DP_OP_425J2_127_3477_n1214), .S(DP_OP_425J2_127_3477_n1215) );
  FADDX1_HVT DP_OP_425J2_127_3477_U764 ( .A(DP_OP_425J2_127_3477_n1255), .B(
        DP_OP_425J2_127_3477_n1257), .CI(DP_OP_425J2_127_3477_n1253), .CO(
        DP_OP_425J2_127_3477_n1212), .S(DP_OP_425J2_127_3477_n1213) );
  FADDX1_HVT DP_OP_425J2_127_3477_U763 ( .A(DP_OP_425J2_127_3477_n1245), .B(
        DP_OP_425J2_127_3477_n1247), .CI(DP_OP_425J2_127_3477_n1412), .CO(
        DP_OP_425J2_127_3477_n1210), .S(DP_OP_425J2_127_3477_n1211) );
  FADDX1_HVT DP_OP_425J2_127_3477_U762 ( .A(DP_OP_425J2_127_3477_n1243), .B(
        DP_OP_425J2_127_3477_n1251), .CI(DP_OP_425J2_127_3477_n1249), .CO(
        DP_OP_425J2_127_3477_n1208), .S(DP_OP_425J2_127_3477_n1209) );
  FADDX1_HVT DP_OP_425J2_127_3477_U761 ( .A(DP_OP_425J2_127_3477_n1239), .B(
        DP_OP_425J2_127_3477_n1241), .CI(DP_OP_425J2_127_3477_n1408), .CO(
        DP_OP_425J2_127_3477_n1206), .S(DP_OP_425J2_127_3477_n1207) );
  FADDX1_HVT DP_OP_425J2_127_3477_U760 ( .A(DP_OP_425J2_127_3477_n1410), .B(
        DP_OP_425J2_127_3477_n1237), .CI(DP_OP_425J2_127_3477_n1406), .CO(
        DP_OP_425J2_127_3477_n1204), .S(DP_OP_425J2_127_3477_n1205) );
  FADDX1_HVT DP_OP_425J2_127_3477_U759 ( .A(DP_OP_425J2_127_3477_n1404), .B(
        DP_OP_425J2_127_3477_n1402), .CI(DP_OP_425J2_127_3477_n1235), .CO(
        DP_OP_425J2_127_3477_n1202), .S(DP_OP_425J2_127_3477_n1203) );
  FADDX1_HVT DP_OP_425J2_127_3477_U758 ( .A(DP_OP_425J2_127_3477_n1400), .B(
        DP_OP_425J2_127_3477_n1392), .CI(DP_OP_425J2_127_3477_n1229), .CO(
        DP_OP_425J2_127_3477_n1200), .S(DP_OP_425J2_127_3477_n1201) );
  FADDX1_HVT DP_OP_425J2_127_3477_U757 ( .A(DP_OP_425J2_127_3477_n1398), .B(
        DP_OP_425J2_127_3477_n1231), .CI(DP_OP_425J2_127_3477_n1233), .CO(
        DP_OP_425J2_127_3477_n1198), .S(DP_OP_425J2_127_3477_n1199) );
  FADDX1_HVT DP_OP_425J2_127_3477_U756 ( .A(DP_OP_425J2_127_3477_n1396), .B(
        DP_OP_425J2_127_3477_n1394), .CI(DP_OP_425J2_127_3477_n1390), .CO(
        DP_OP_425J2_127_3477_n1196), .S(DP_OP_425J2_127_3477_n1197) );
  FADDX1_HVT DP_OP_425J2_127_3477_U755 ( .A(DP_OP_425J2_127_3477_n1225), .B(
        DP_OP_425J2_127_3477_n1227), .CI(DP_OP_425J2_127_3477_n1388), .CO(
        DP_OP_425J2_127_3477_n1194), .S(DP_OP_425J2_127_3477_n1195) );
  FADDX1_HVT DP_OP_425J2_127_3477_U754 ( .A(DP_OP_425J2_127_3477_n1386), .B(
        DP_OP_425J2_127_3477_n1219), .CI(DP_OP_425J2_127_3477_n1384), .CO(
        DP_OP_425J2_127_3477_n1192), .S(DP_OP_425J2_127_3477_n1193) );
  FADDX1_HVT DP_OP_425J2_127_3477_U753 ( .A(DP_OP_425J2_127_3477_n1217), .B(
        DP_OP_425J2_127_3477_n1223), .CI(DP_OP_425J2_127_3477_n1221), .CO(
        DP_OP_425J2_127_3477_n1190), .S(DP_OP_425J2_127_3477_n1191) );
  FADDX1_HVT DP_OP_425J2_127_3477_U752 ( .A(DP_OP_425J2_127_3477_n1215), .B(
        DP_OP_425J2_127_3477_n1213), .CI(DP_OP_425J2_127_3477_n1209), .CO(
        DP_OP_425J2_127_3477_n1188), .S(DP_OP_425J2_127_3477_n1189) );
  FADDX1_HVT DP_OP_425J2_127_3477_U751 ( .A(DP_OP_425J2_127_3477_n1211), .B(
        DP_OP_425J2_127_3477_n1382), .CI(DP_OP_425J2_127_3477_n1207), .CO(
        DP_OP_425J2_127_3477_n1186), .S(DP_OP_425J2_127_3477_n1187) );
  FADDX1_HVT DP_OP_425J2_127_3477_U750 ( .A(DP_OP_425J2_127_3477_n1380), .B(
        DP_OP_425J2_127_3477_n1378), .CI(DP_OP_425J2_127_3477_n1205), .CO(
        DP_OP_425J2_127_3477_n1184), .S(DP_OP_425J2_127_3477_n1185) );
  FADDX1_HVT DP_OP_425J2_127_3477_U749 ( .A(DP_OP_425J2_127_3477_n1376), .B(
        DP_OP_425J2_127_3477_n1374), .CI(DP_OP_425J2_127_3477_n1203), .CO(
        DP_OP_425J2_127_3477_n1182), .S(DP_OP_425J2_127_3477_n1183) );
  FADDX1_HVT DP_OP_425J2_127_3477_U748 ( .A(DP_OP_425J2_127_3477_n1372), .B(
        DP_OP_425J2_127_3477_n1199), .CI(DP_OP_425J2_127_3477_n1197), .CO(
        DP_OP_425J2_127_3477_n1180), .S(DP_OP_425J2_127_3477_n1181) );
  FADDX1_HVT DP_OP_425J2_127_3477_U747 ( .A(DP_OP_425J2_127_3477_n1370), .B(
        DP_OP_425J2_127_3477_n1201), .CI(DP_OP_425J2_127_3477_n1195), .CO(
        DP_OP_425J2_127_3477_n1178), .S(DP_OP_425J2_127_3477_n1179) );
  FADDX1_HVT DP_OP_425J2_127_3477_U746 ( .A(DP_OP_425J2_127_3477_n1368), .B(
        DP_OP_425J2_127_3477_n1191), .CI(DP_OP_425J2_127_3477_n1366), .CO(
        DP_OP_425J2_127_3477_n1176), .S(DP_OP_425J2_127_3477_n1177) );
  FADDX1_HVT DP_OP_425J2_127_3477_U745 ( .A(DP_OP_425J2_127_3477_n1193), .B(
        DP_OP_425J2_127_3477_n1189), .CI(DP_OP_425J2_127_3477_n1187), .CO(
        DP_OP_425J2_127_3477_n1174), .S(DP_OP_425J2_127_3477_n1175) );
  FADDX1_HVT DP_OP_425J2_127_3477_U744 ( .A(DP_OP_425J2_127_3477_n1364), .B(
        DP_OP_425J2_127_3477_n1362), .CI(DP_OP_425J2_127_3477_n1185), .CO(
        DP_OP_425J2_127_3477_n1172), .S(DP_OP_425J2_127_3477_n1173) );
  FADDX1_HVT DP_OP_425J2_127_3477_U743 ( .A(DP_OP_425J2_127_3477_n1360), .B(
        DP_OP_425J2_127_3477_n1183), .CI(DP_OP_425J2_127_3477_n1181), .CO(
        DP_OP_425J2_127_3477_n1170), .S(DP_OP_425J2_127_3477_n1171) );
  FADDX1_HVT DP_OP_425J2_127_3477_U742 ( .A(DP_OP_425J2_127_3477_n1179), .B(
        DP_OP_425J2_127_3477_n1358), .CI(DP_OP_425J2_127_3477_n1177), .CO(
        DP_OP_425J2_127_3477_n1168), .S(DP_OP_425J2_127_3477_n1169) );
  FADDX1_HVT DP_OP_425J2_127_3477_U741 ( .A(DP_OP_425J2_127_3477_n1356), .B(
        DP_OP_425J2_127_3477_n1175), .CI(DP_OP_425J2_127_3477_n1354), .CO(
        DP_OP_425J2_127_3477_n1166), .S(DP_OP_425J2_127_3477_n1167) );
  FADDX1_HVT DP_OP_425J2_127_3477_U740 ( .A(DP_OP_425J2_127_3477_n1173), .B(
        DP_OP_425J2_127_3477_n1171), .CI(DP_OP_425J2_127_3477_n1352), .CO(
        DP_OP_425J2_127_3477_n1164), .S(DP_OP_425J2_127_3477_n1165) );
  FADDX1_HVT DP_OP_425J2_127_3477_U739 ( .A(DP_OP_425J2_127_3477_n1169), .B(
        DP_OP_425J2_127_3477_n1350), .CI(DP_OP_425J2_127_3477_n1167), .CO(
        DP_OP_425J2_127_3477_n1162), .S(DP_OP_425J2_127_3477_n1163) );
  OR2X1_HVT DP_OP_425J2_127_3477_U738 ( .A1(DP_OP_425J2_127_3477_n2979), .A2(
        DP_OP_425J2_127_3477_n2452), .Y(DP_OP_425J2_127_3477_n1160) );
  FADDX1_HVT DP_OP_425J2_127_3477_U736 ( .A(DP_OP_425J2_127_3477_n2144), .B(
        DP_OP_425J2_127_3477_n1924), .CI(DP_OP_425J2_127_3477_n1880), .CO(
        DP_OP_425J2_127_3477_n1158), .S(DP_OP_425J2_127_3477_n1159) );
  FADDX1_HVT DP_OP_425J2_127_3477_U735 ( .A(DP_OP_425J2_127_3477_n2584), .B(
        DP_OP_425J2_127_3477_n2012), .CI(DP_OP_425J2_127_3477_n2364), .CO(
        DP_OP_425J2_127_3477_n1156), .S(DP_OP_425J2_127_3477_n1157) );
  FADDX1_HVT DP_OP_425J2_127_3477_U734 ( .A(DP_OP_425J2_127_3477_n2804), .B(
        DP_OP_425J2_127_3477_n2628), .CI(DP_OP_425J2_127_3477_n2188), .CO(
        DP_OP_425J2_127_3477_n1154), .S(DP_OP_425J2_127_3477_n1155) );
  FADDX1_HVT DP_OP_425J2_127_3477_U733 ( .A(DP_OP_425J2_127_3477_n2276), .B(
        DP_OP_425J2_127_3477_n2100), .CI(DP_OP_425J2_127_3477_n2848), .CO(
        DP_OP_425J2_127_3477_n1152), .S(DP_OP_425J2_127_3477_n1153) );
  FADDX1_HVT DP_OP_425J2_127_3477_U732 ( .A(DP_OP_425J2_127_3477_n2408), .B(
        DP_OP_425J2_127_3477_n2892), .CI(DP_OP_425J2_127_3477_n2672), .CO(
        DP_OP_425J2_127_3477_n1150), .S(DP_OP_425J2_127_3477_n1151) );
  FADDX1_HVT DP_OP_425J2_127_3477_U731 ( .A(DP_OP_425J2_127_3477_n2496), .B(
        DP_OP_425J2_127_3477_n2716), .CI(DP_OP_425J2_127_3477_n2540), .CO(
        DP_OP_425J2_127_3477_n1148), .S(DP_OP_425J2_127_3477_n1149) );
  FADDX1_HVT DP_OP_425J2_127_3477_U730 ( .A(DP_OP_425J2_127_3477_n2232), .B(
        DP_OP_425J2_127_3477_n2056), .CI(DP_OP_425J2_127_3477_n2936), .CO(
        DP_OP_425J2_127_3477_n1146), .S(DP_OP_425J2_127_3477_n1147) );
  FADDX1_HVT DP_OP_425J2_127_3477_U729 ( .A(DP_OP_425J2_127_3477_n2760), .B(
        DP_OP_425J2_127_3477_n1968), .CI(DP_OP_425J2_127_3477_n2320), .CO(
        DP_OP_425J2_127_3477_n1144), .S(DP_OP_425J2_127_3477_n1145) );
  FADDX1_HVT DP_OP_425J2_127_3477_U728 ( .A(DP_OP_425J2_127_3477_n2371), .B(
        DP_OP_425J2_127_3477_n2999), .CI(DP_OP_425J2_127_3477_n1931), .CO(
        DP_OP_425J2_127_3477_n1142), .S(DP_OP_425J2_127_3477_n1143) );
  FADDX1_HVT DP_OP_425J2_127_3477_U727 ( .A(DP_OP_425J2_127_3477_n2378), .B(
        DP_OP_425J2_127_3477_n2992), .CI(DP_OP_425J2_127_3477_n2985), .CO(
        DP_OP_425J2_127_3477_n1140), .S(DP_OP_425J2_127_3477_n1141) );
  FADDX1_HVT DP_OP_425J2_127_3477_U726 ( .A(DP_OP_425J2_127_3477_n2334), .B(
        DP_OP_425J2_127_3477_n2957), .CI(DP_OP_425J2_127_3477_n2950), .CO(
        DP_OP_425J2_127_3477_n1138), .S(DP_OP_425J2_127_3477_n1139) );
  FADDX1_HVT DP_OP_425J2_127_3477_U725 ( .A(DP_OP_425J2_127_3477_n2297), .B(
        DP_OP_425J2_127_3477_n2943), .CI(DP_OP_425J2_127_3477_n2913), .CO(
        DP_OP_425J2_127_3477_n1136), .S(DP_OP_425J2_127_3477_n1137) );
  FADDX1_HVT DP_OP_425J2_127_3477_U724 ( .A(DP_OP_425J2_127_3477_n2290), .B(
        DP_OP_425J2_127_3477_n1938), .CI(DP_OP_425J2_127_3477_n2906), .CO(
        DP_OP_425J2_127_3477_n1134), .S(DP_OP_425J2_127_3477_n1135) );
  FADDX1_HVT DP_OP_425J2_127_3477_U723 ( .A(DP_OP_425J2_127_3477_n2327), .B(
        DP_OP_425J2_127_3477_n2899), .CI(DP_OP_425J2_127_3477_n1945), .CO(
        DP_OP_425J2_127_3477_n1132), .S(DP_OP_425J2_127_3477_n1133) );
  FADDX1_HVT DP_OP_425J2_127_3477_U722 ( .A(DP_OP_425J2_127_3477_n2283), .B(
        DP_OP_425J2_127_3477_n2869), .CI(DP_OP_425J2_127_3477_n1975), .CO(
        DP_OP_425J2_127_3477_n1130), .S(DP_OP_425J2_127_3477_n1131) );
  FADDX1_HVT DP_OP_425J2_127_3477_U721 ( .A(DP_OP_425J2_127_3477_n2253), .B(
        DP_OP_425J2_127_3477_n2862), .CI(DP_OP_425J2_127_3477_n2855), .CO(
        DP_OP_425J2_127_3477_n1128), .S(DP_OP_425J2_127_3477_n1129) );
  FADDX1_HVT DP_OP_425J2_127_3477_U720 ( .A(DP_OP_425J2_127_3477_n2246), .B(
        DP_OP_425J2_127_3477_n1982), .CI(DP_OP_425J2_127_3477_n2825), .CO(
        DP_OP_425J2_127_3477_n1126), .S(DP_OP_425J2_127_3477_n1127) );
  FADDX1_HVT DP_OP_425J2_127_3477_U719 ( .A(DP_OP_425J2_127_3477_n2239), .B(
        DP_OP_425J2_127_3477_n1989), .CI(DP_OP_425J2_127_3477_n2818), .CO(
        DP_OP_425J2_127_3477_n1124), .S(DP_OP_425J2_127_3477_n1125) );
  FADDX1_HVT DP_OP_425J2_127_3477_U718 ( .A(DP_OP_425J2_127_3477_n2019), .B(
        DP_OP_425J2_127_3477_n2026), .CI(DP_OP_425J2_127_3477_n2033), .CO(
        DP_OP_425J2_127_3477_n1122), .S(DP_OP_425J2_127_3477_n1123) );
  FADDX1_HVT DP_OP_425J2_127_3477_U717 ( .A(DP_OP_425J2_127_3477_n2811), .B(
        DP_OP_425J2_127_3477_n2063), .CI(DP_OP_425J2_127_3477_n2070), .CO(
        DP_OP_425J2_127_3477_n1120), .S(DP_OP_425J2_127_3477_n1121) );
  FADDX1_HVT DP_OP_425J2_127_3477_U716 ( .A(DP_OP_425J2_127_3477_n2781), .B(
        DP_OP_425J2_127_3477_n2077), .CI(DP_OP_425J2_127_3477_n2107), .CO(
        DP_OP_425J2_127_3477_n1118), .S(DP_OP_425J2_127_3477_n1119) );
  FADDX1_HVT DP_OP_425J2_127_3477_U715 ( .A(DP_OP_425J2_127_3477_n2774), .B(
        DP_OP_425J2_127_3477_n2114), .CI(DP_OP_425J2_127_3477_n2121), .CO(
        DP_OP_425J2_127_3477_n1116), .S(DP_OP_425J2_127_3477_n1117) );
  FADDX1_HVT DP_OP_425J2_127_3477_U714 ( .A(DP_OP_425J2_127_3477_n2767), .B(
        DP_OP_425J2_127_3477_n2151), .CI(DP_OP_425J2_127_3477_n2158), .CO(
        DP_OP_425J2_127_3477_n1114), .S(DP_OP_425J2_127_3477_n1115) );
  FADDX1_HVT DP_OP_425J2_127_3477_U713 ( .A(DP_OP_425J2_127_3477_n2737), .B(
        DP_OP_425J2_127_3477_n2165), .CI(DP_OP_425J2_127_3477_n2195), .CO(
        DP_OP_425J2_127_3477_n1112), .S(DP_OP_425J2_127_3477_n1113) );
  FADDX1_HVT DP_OP_425J2_127_3477_U712 ( .A(DP_OP_425J2_127_3477_n2730), .B(
        DP_OP_425J2_127_3477_n2202), .CI(DP_OP_425J2_127_3477_n2209), .CO(
        DP_OP_425J2_127_3477_n1110), .S(DP_OP_425J2_127_3477_n1111) );
  FADDX1_HVT DP_OP_425J2_127_3477_U711 ( .A(DP_OP_425J2_127_3477_n2723), .B(
        DP_OP_425J2_127_3477_n2341), .CI(DP_OP_425J2_127_3477_n2385), .CO(
        DP_OP_425J2_127_3477_n1108), .S(DP_OP_425J2_127_3477_n1109) );
  FADDX1_HVT DP_OP_425J2_127_3477_U710 ( .A(DP_OP_425J2_127_3477_n2693), .B(
        DP_OP_425J2_127_3477_n2415), .CI(DP_OP_425J2_127_3477_n2422), .CO(
        DP_OP_425J2_127_3477_n1106), .S(DP_OP_425J2_127_3477_n1107) );
  FADDX1_HVT DP_OP_425J2_127_3477_U709 ( .A(DP_OP_425J2_127_3477_n2686), .B(
        DP_OP_425J2_127_3477_n2429), .CI(DP_OP_425J2_127_3477_n2459), .CO(
        DP_OP_425J2_127_3477_n1104), .S(DP_OP_425J2_127_3477_n1105) );
  FADDX1_HVT DP_OP_425J2_127_3477_U708 ( .A(DP_OP_425J2_127_3477_n2679), .B(
        DP_OP_425J2_127_3477_n2466), .CI(DP_OP_425J2_127_3477_n2473), .CO(
        DP_OP_425J2_127_3477_n1102), .S(DP_OP_425J2_127_3477_n1103) );
  FADDX1_HVT DP_OP_425J2_127_3477_U707 ( .A(DP_OP_425J2_127_3477_n2649), .B(
        DP_OP_425J2_127_3477_n2503), .CI(DP_OP_425J2_127_3477_n2510), .CO(
        DP_OP_425J2_127_3477_n1100), .S(DP_OP_425J2_127_3477_n1101) );
  FADDX1_HVT DP_OP_425J2_127_3477_U706 ( .A(DP_OP_425J2_127_3477_n2642), .B(
        DP_OP_425J2_127_3477_n2517), .CI(DP_OP_425J2_127_3477_n2547), .CO(
        DP_OP_425J2_127_3477_n1098), .S(DP_OP_425J2_127_3477_n1099) );
  FADDX1_HVT DP_OP_425J2_127_3477_U705 ( .A(DP_OP_425J2_127_3477_n2635), .B(
        DP_OP_425J2_127_3477_n2554), .CI(DP_OP_425J2_127_3477_n2561), .CO(
        DP_OP_425J2_127_3477_n1096), .S(DP_OP_425J2_127_3477_n1097) );
  FADDX1_HVT DP_OP_425J2_127_3477_U704 ( .A(DP_OP_425J2_127_3477_n2591), .B(
        DP_OP_425J2_127_3477_n2598), .CI(DP_OP_425J2_127_3477_n2605), .CO(
        DP_OP_425J2_127_3477_n1094), .S(DP_OP_425J2_127_3477_n1095) );
  FADDX1_HVT DP_OP_425J2_127_3477_U703 ( .A(DP_OP_425J2_127_3477_n1348), .B(
        DP_OP_425J2_127_3477_n1336), .CI(DP_OP_425J2_127_3477_n1334), .CO(
        DP_OP_425J2_127_3477_n1092), .S(DP_OP_425J2_127_3477_n1093) );
  FADDX1_HVT DP_OP_425J2_127_3477_U702 ( .A(DP_OP_425J2_127_3477_n1332), .B(
        DP_OP_425J2_127_3477_n1338), .CI(DP_OP_425J2_127_3477_n1161), .CO(
        DP_OP_425J2_127_3477_n1090), .S(DP_OP_425J2_127_3477_n1091) );
  FADDX1_HVT DP_OP_425J2_127_3477_U701 ( .A(DP_OP_425J2_127_3477_n1342), .B(
        DP_OP_425J2_127_3477_n1346), .CI(DP_OP_425J2_127_3477_n1340), .CO(
        DP_OP_425J2_127_3477_n1088), .S(DP_OP_425J2_127_3477_n1089) );
  FADDX1_HVT DP_OP_425J2_127_3477_U700 ( .A(DP_OP_425J2_127_3477_n1344), .B(
        DP_OP_425J2_127_3477_n1308), .CI(DP_OP_425J2_127_3477_n1306), .CO(
        DP_OP_425J2_127_3477_n1086), .S(DP_OP_425J2_127_3477_n1087) );
  FADDX1_HVT DP_OP_425J2_127_3477_U699 ( .A(DP_OP_425J2_127_3477_n1310), .B(
        DP_OP_425J2_127_3477_n1282), .CI(DP_OP_425J2_127_3477_n1330), .CO(
        DP_OP_425J2_127_3477_n1084), .S(DP_OP_425J2_127_3477_n1085) );
  FADDX1_HVT DP_OP_425J2_127_3477_U698 ( .A(DP_OP_425J2_127_3477_n1302), .B(
        DP_OP_425J2_127_3477_n1284), .CI(DP_OP_425J2_127_3477_n1328), .CO(
        DP_OP_425J2_127_3477_n1082), .S(DP_OP_425J2_127_3477_n1083) );
  FADDX1_HVT DP_OP_425J2_127_3477_U697 ( .A(DP_OP_425J2_127_3477_n1300), .B(
        DP_OP_425J2_127_3477_n1286), .CI(DP_OP_425J2_127_3477_n1326), .CO(
        DP_OP_425J2_127_3477_n1080), .S(DP_OP_425J2_127_3477_n1081) );
  FADDX1_HVT DP_OP_425J2_127_3477_U696 ( .A(DP_OP_425J2_127_3477_n1296), .B(
        DP_OP_425J2_127_3477_n1324), .CI(DP_OP_425J2_127_3477_n1322), .CO(
        DP_OP_425J2_127_3477_n1078), .S(DP_OP_425J2_127_3477_n1079) );
  FADDX1_HVT DP_OP_425J2_127_3477_U695 ( .A(DP_OP_425J2_127_3477_n1290), .B(
        DP_OP_425J2_127_3477_n1320), .CI(DP_OP_425J2_127_3477_n1318), .CO(
        DP_OP_425J2_127_3477_n1076), .S(DP_OP_425J2_127_3477_n1077) );
  FADDX1_HVT DP_OP_425J2_127_3477_U694 ( .A(DP_OP_425J2_127_3477_n1298), .B(
        DP_OP_425J2_127_3477_n1316), .CI(DP_OP_425J2_127_3477_n1314), .CO(
        DP_OP_425J2_127_3477_n1074), .S(DP_OP_425J2_127_3477_n1075) );
  FADDX1_HVT DP_OP_425J2_127_3477_U693 ( .A(DP_OP_425J2_127_3477_n1292), .B(
        DP_OP_425J2_127_3477_n1312), .CI(DP_OP_425J2_127_3477_n1304), .CO(
        DP_OP_425J2_127_3477_n1072), .S(DP_OP_425J2_127_3477_n1073) );
  FADDX1_HVT DP_OP_425J2_127_3477_U692 ( .A(DP_OP_425J2_127_3477_n1294), .B(
        DP_OP_425J2_127_3477_n1288), .CI(DP_OP_425J2_127_3477_n1151), .CO(
        DP_OP_425J2_127_3477_n1070), .S(DP_OP_425J2_127_3477_n1071) );
  FADDX1_HVT DP_OP_425J2_127_3477_U691 ( .A(DP_OP_425J2_127_3477_n1147), .B(
        DP_OP_425J2_127_3477_n1145), .CI(DP_OP_425J2_127_3477_n1149), .CO(
        DP_OP_425J2_127_3477_n1068), .S(DP_OP_425J2_127_3477_n1069) );
  FADDX1_HVT DP_OP_425J2_127_3477_U690 ( .A(DP_OP_425J2_127_3477_n1157), .B(
        DP_OP_425J2_127_3477_n1155), .CI(DP_OP_425J2_127_3477_n1159), .CO(
        DP_OP_425J2_127_3477_n1066), .S(DP_OP_425J2_127_3477_n1067) );
  FADDX1_HVT DP_OP_425J2_127_3477_U689 ( .A(DP_OP_425J2_127_3477_n1153), .B(
        DP_OP_425J2_127_3477_n1101), .CI(DP_OP_425J2_127_3477_n1103), .CO(
        DP_OP_425J2_127_3477_n1064), .S(DP_OP_425J2_127_3477_n1065) );
  FADDX1_HVT DP_OP_425J2_127_3477_U688 ( .A(DP_OP_425J2_127_3477_n1099), .B(
        DP_OP_425J2_127_3477_n1135), .CI(DP_OP_425J2_127_3477_n1131), .CO(
        DP_OP_425J2_127_3477_n1062), .S(DP_OP_425J2_127_3477_n1063) );
  FADDX1_HVT DP_OP_425J2_127_3477_U687 ( .A(DP_OP_425J2_127_3477_n1137), .B(
        DP_OP_425J2_127_3477_n1121), .CI(DP_OP_425J2_127_3477_n1127), .CO(
        DP_OP_425J2_127_3477_n1060), .S(DP_OP_425J2_127_3477_n1061) );
  FADDX1_HVT DP_OP_425J2_127_3477_U686 ( .A(DP_OP_425J2_127_3477_n1125), .B(
        DP_OP_425J2_127_3477_n1123), .CI(DP_OP_425J2_127_3477_n1107), .CO(
        DP_OP_425J2_127_3477_n1058), .S(DP_OP_425J2_127_3477_n1059) );
  FADDX1_HVT DP_OP_425J2_127_3477_U685 ( .A(DP_OP_425J2_127_3477_n1129), .B(
        DP_OP_425J2_127_3477_n1097), .CI(DP_OP_425J2_127_3477_n1095), .CO(
        DP_OP_425J2_127_3477_n1056), .S(DP_OP_425J2_127_3477_n1057) );
  FADDX1_HVT DP_OP_425J2_127_3477_U684 ( .A(DP_OP_425J2_127_3477_n1133), .B(
        DP_OP_425J2_127_3477_n1115), .CI(DP_OP_425J2_127_3477_n1117), .CO(
        DP_OP_425J2_127_3477_n1054), .S(DP_OP_425J2_127_3477_n1055) );
  FADDX1_HVT DP_OP_425J2_127_3477_U683 ( .A(DP_OP_425J2_127_3477_n1113), .B(
        DP_OP_425J2_127_3477_n1111), .CI(DP_OP_425J2_127_3477_n1105), .CO(
        DP_OP_425J2_127_3477_n1052), .S(DP_OP_425J2_127_3477_n1053) );
  FADDX1_HVT DP_OP_425J2_127_3477_U682 ( .A(DP_OP_425J2_127_3477_n1109), .B(
        DP_OP_425J2_127_3477_n1143), .CI(DP_OP_425J2_127_3477_n1141), .CO(
        DP_OP_425J2_127_3477_n1050), .S(DP_OP_425J2_127_3477_n1051) );
  FADDX1_HVT DP_OP_425J2_127_3477_U681 ( .A(DP_OP_425J2_127_3477_n1139), .B(
        DP_OP_425J2_127_3477_n1119), .CI(DP_OP_425J2_127_3477_n1280), .CO(
        DP_OP_425J2_127_3477_n1048), .S(DP_OP_425J2_127_3477_n1049) );
  FADDX1_HVT DP_OP_425J2_127_3477_U680 ( .A(DP_OP_425J2_127_3477_n1278), .B(
        DP_OP_425J2_127_3477_n1276), .CI(DP_OP_425J2_127_3477_n1274), .CO(
        DP_OP_425J2_127_3477_n1046), .S(DP_OP_425J2_127_3477_n1047) );
  FADDX1_HVT DP_OP_425J2_127_3477_U679 ( .A(DP_OP_425J2_127_3477_n1272), .B(
        DP_OP_425J2_127_3477_n1260), .CI(DP_OP_425J2_127_3477_n1258), .CO(
        DP_OP_425J2_127_3477_n1044), .S(DP_OP_425J2_127_3477_n1045) );
  FADDX1_HVT DP_OP_425J2_127_3477_U678 ( .A(DP_OP_425J2_127_3477_n1264), .B(
        DP_OP_425J2_127_3477_n1262), .CI(DP_OP_425J2_127_3477_n1270), .CO(
        DP_OP_425J2_127_3477_n1042), .S(DP_OP_425J2_127_3477_n1043) );
  FADDX1_HVT DP_OP_425J2_127_3477_U677 ( .A(DP_OP_425J2_127_3477_n1268), .B(
        DP_OP_425J2_127_3477_n1266), .CI(DP_OP_425J2_127_3477_n1093), .CO(
        DP_OP_425J2_127_3477_n1040), .S(DP_OP_425J2_127_3477_n1041) );
  FADDX1_HVT DP_OP_425J2_127_3477_U676 ( .A(DP_OP_425J2_127_3477_n1256), .B(
        DP_OP_425J2_127_3477_n1254), .CI(DP_OP_425J2_127_3477_n1087), .CO(
        DP_OP_425J2_127_3477_n1038), .S(DP_OP_425J2_127_3477_n1039) );
  FADDX1_HVT DP_OP_425J2_127_3477_U675 ( .A(DP_OP_425J2_127_3477_n1091), .B(
        DP_OP_425J2_127_3477_n1089), .CI(DP_OP_425J2_127_3477_n1252), .CO(
        DP_OP_425J2_127_3477_n1036), .S(DP_OP_425J2_127_3477_n1037) );
  FADDX1_HVT DP_OP_425J2_127_3477_U674 ( .A(DP_OP_425J2_127_3477_n1240), .B(
        DP_OP_425J2_127_3477_n1085), .CI(DP_OP_425J2_127_3477_n1071), .CO(
        DP_OP_425J2_127_3477_n1034), .S(DP_OP_425J2_127_3477_n1035) );
  FADDX1_HVT DP_OP_425J2_127_3477_U673 ( .A(DP_OP_425J2_127_3477_n1238), .B(
        DP_OP_425J2_127_3477_n1081), .CI(DP_OP_425J2_127_3477_n1083), .CO(
        DP_OP_425J2_127_3477_n1032), .S(DP_OP_425J2_127_3477_n1033) );
  FADDX1_HVT DP_OP_425J2_127_3477_U672 ( .A(DP_OP_425J2_127_3477_n1242), .B(
        DP_OP_425J2_127_3477_n1079), .CI(DP_OP_425J2_127_3477_n1077), .CO(
        DP_OP_425J2_127_3477_n1030), .S(DP_OP_425J2_127_3477_n1031) );
  FADDX1_HVT DP_OP_425J2_127_3477_U671 ( .A(DP_OP_425J2_127_3477_n1250), .B(
        DP_OP_425J2_127_3477_n1073), .CI(DP_OP_425J2_127_3477_n1075), .CO(
        DP_OP_425J2_127_3477_n1028), .S(DP_OP_425J2_127_3477_n1029) );
  FADDX1_HVT DP_OP_425J2_127_3477_U670 ( .A(DP_OP_425J2_127_3477_n1248), .B(
        DP_OP_425J2_127_3477_n1244), .CI(DP_OP_425J2_127_3477_n1246), .CO(
        DP_OP_425J2_127_3477_n1026), .S(DP_OP_425J2_127_3477_n1027) );
  FADDX1_HVT DP_OP_425J2_127_3477_U669 ( .A(DP_OP_425J2_127_3477_n1067), .B(
        DP_OP_425J2_127_3477_n1236), .CI(DP_OP_425J2_127_3477_n1065), .CO(
        DP_OP_425J2_127_3477_n1024), .S(DP_OP_425J2_127_3477_n1025) );
  FADDX1_HVT DP_OP_425J2_127_3477_U668 ( .A(DP_OP_425J2_127_3477_n1069), .B(
        DP_OP_425J2_127_3477_n1059), .CI(DP_OP_425J2_127_3477_n1061), .CO(
        DP_OP_425J2_127_3477_n1022), .S(DP_OP_425J2_127_3477_n1023) );
  FADDX1_HVT DP_OP_425J2_127_3477_U667 ( .A(DP_OP_425J2_127_3477_n1057), .B(
        DP_OP_425J2_127_3477_n1051), .CI(DP_OP_425J2_127_3477_n1234), .CO(
        DP_OP_425J2_127_3477_n1020), .S(DP_OP_425J2_127_3477_n1021) );
  FADDX1_HVT DP_OP_425J2_127_3477_U666 ( .A(DP_OP_425J2_127_3477_n1053), .B(
        DP_OP_425J2_127_3477_n1063), .CI(DP_OP_425J2_127_3477_n1055), .CO(
        DP_OP_425J2_127_3477_n1018), .S(DP_OP_425J2_127_3477_n1019) );
  FADDX1_HVT DP_OP_425J2_127_3477_U665 ( .A(DP_OP_425J2_127_3477_n1049), .B(
        DP_OP_425J2_127_3477_n1232), .CI(DP_OP_425J2_127_3477_n1228), .CO(
        DP_OP_425J2_127_3477_n1016), .S(DP_OP_425J2_127_3477_n1017) );
  FADDX1_HVT DP_OP_425J2_127_3477_U664 ( .A(DP_OP_425J2_127_3477_n1230), .B(
        DP_OP_425J2_127_3477_n1226), .CI(DP_OP_425J2_127_3477_n1224), .CO(
        DP_OP_425J2_127_3477_n1014), .S(DP_OP_425J2_127_3477_n1015) );
  FADDX1_HVT DP_OP_425J2_127_3477_U663 ( .A(DP_OP_425J2_127_3477_n1047), .B(
        DP_OP_425J2_127_3477_n1222), .CI(DP_OP_425J2_127_3477_n1220), .CO(
        DP_OP_425J2_127_3477_n1012), .S(DP_OP_425J2_127_3477_n1013) );
  FADDX1_HVT DP_OP_425J2_127_3477_U662 ( .A(DP_OP_425J2_127_3477_n1218), .B(
        DP_OP_425J2_127_3477_n1043), .CI(DP_OP_425J2_127_3477_n1041), .CO(
        DP_OP_425J2_127_3477_n1010), .S(DP_OP_425J2_127_3477_n1011) );
  FADDX1_HVT DP_OP_425J2_127_3477_U661 ( .A(DP_OP_425J2_127_3477_n1216), .B(
        DP_OP_425J2_127_3477_n1214), .CI(DP_OP_425J2_127_3477_n1045), .CO(
        DP_OP_425J2_127_3477_n1008), .S(DP_OP_425J2_127_3477_n1009) );
  FADDX1_HVT DP_OP_425J2_127_3477_U660 ( .A(DP_OP_425J2_127_3477_n1037), .B(
        DP_OP_425J2_127_3477_n1212), .CI(DP_OP_425J2_127_3477_n1039), .CO(
        DP_OP_425J2_127_3477_n1006), .S(DP_OP_425J2_127_3477_n1007) );
  FADDX1_HVT DP_OP_425J2_127_3477_U659 ( .A(DP_OP_425J2_127_3477_n1031), .B(
        DP_OP_425J2_127_3477_n1035), .CI(DP_OP_425J2_127_3477_n1206), .CO(
        DP_OP_425J2_127_3477_n1004), .S(DP_OP_425J2_127_3477_n1005) );
  FADDX1_HVT DP_OP_425J2_127_3477_U658 ( .A(DP_OP_425J2_127_3477_n1210), .B(
        DP_OP_425J2_127_3477_n1029), .CI(DP_OP_425J2_127_3477_n1033), .CO(
        DP_OP_425J2_127_3477_n1002), .S(DP_OP_425J2_127_3477_n1003) );
  FADDX1_HVT DP_OP_425J2_127_3477_U657 ( .A(DP_OP_425J2_127_3477_n1208), .B(
        DP_OP_425J2_127_3477_n1027), .CI(DP_OP_425J2_127_3477_n1204), .CO(
        DP_OP_425J2_127_3477_n1000), .S(DP_OP_425J2_127_3477_n1001) );
  FADDX1_HVT DP_OP_425J2_127_3477_U656 ( .A(DP_OP_425J2_127_3477_n1025), .B(
        DP_OP_425J2_127_3477_n1023), .CI(DP_OP_425J2_127_3477_n1021), .CO(
        DP_OP_425J2_127_3477_n998), .S(DP_OP_425J2_127_3477_n999) );
  FADDX1_HVT DP_OP_425J2_127_3477_U655 ( .A(DP_OP_425J2_127_3477_n1019), .B(
        DP_OP_425J2_127_3477_n1202), .CI(DP_OP_425J2_127_3477_n1017), .CO(
        DP_OP_425J2_127_3477_n996), .S(DP_OP_425J2_127_3477_n997) );
  FADDX1_HVT DP_OP_425J2_127_3477_U654 ( .A(DP_OP_425J2_127_3477_n1200), .B(
        DP_OP_425J2_127_3477_n1198), .CI(DP_OP_425J2_127_3477_n1196), .CO(
        DP_OP_425J2_127_3477_n994), .S(DP_OP_425J2_127_3477_n995) );
  FADDX1_HVT DP_OP_425J2_127_3477_U653 ( .A(DP_OP_425J2_127_3477_n1015), .B(
        DP_OP_425J2_127_3477_n1194), .CI(DP_OP_425J2_127_3477_n1013), .CO(
        DP_OP_425J2_127_3477_n992), .S(DP_OP_425J2_127_3477_n993) );
  FADDX1_HVT DP_OP_425J2_127_3477_U652 ( .A(DP_OP_425J2_127_3477_n1192), .B(
        DP_OP_425J2_127_3477_n1009), .CI(DP_OP_425J2_127_3477_n1011), .CO(
        DP_OP_425J2_127_3477_n990), .S(DP_OP_425J2_127_3477_n991) );
  FADDX1_HVT DP_OP_425J2_127_3477_U651 ( .A(DP_OP_425J2_127_3477_n1190), .B(
        DP_OP_425J2_127_3477_n1188), .CI(DP_OP_425J2_127_3477_n1007), .CO(
        DP_OP_425J2_127_3477_n988), .S(DP_OP_425J2_127_3477_n989) );
  FADDX1_HVT DP_OP_425J2_127_3477_U650 ( .A(DP_OP_425J2_127_3477_n1186), .B(
        DP_OP_425J2_127_3477_n1003), .CI(DP_OP_425J2_127_3477_n1001), .CO(
        DP_OP_425J2_127_3477_n986), .S(DP_OP_425J2_127_3477_n987) );
  FADDX1_HVT DP_OP_425J2_127_3477_U649 ( .A(DP_OP_425J2_127_3477_n1005), .B(
        DP_OP_425J2_127_3477_n1184), .CI(DP_OP_425J2_127_3477_n999), .CO(
        DP_OP_425J2_127_3477_n984), .S(DP_OP_425J2_127_3477_n985) );
  FADDX1_HVT DP_OP_425J2_127_3477_U648 ( .A(DP_OP_425J2_127_3477_n1182), .B(
        DP_OP_425J2_127_3477_n997), .CI(DP_OP_425J2_127_3477_n1180), .CO(
        DP_OP_425J2_127_3477_n982), .S(DP_OP_425J2_127_3477_n983) );
  FADDX1_HVT DP_OP_425J2_127_3477_U647 ( .A(DP_OP_425J2_127_3477_n995), .B(
        DP_OP_425J2_127_3477_n1178), .CI(DP_OP_425J2_127_3477_n993), .CO(
        DP_OP_425J2_127_3477_n980), .S(DP_OP_425J2_127_3477_n981) );
  FADDX1_HVT DP_OP_425J2_127_3477_U646 ( .A(DP_OP_425J2_127_3477_n1176), .B(
        DP_OP_425J2_127_3477_n991), .CI(DP_OP_425J2_127_3477_n989), .CO(
        DP_OP_425J2_127_3477_n978), .S(DP_OP_425J2_127_3477_n979) );
  FADDX1_HVT DP_OP_425J2_127_3477_U645 ( .A(DP_OP_425J2_127_3477_n1174), .B(
        DP_OP_425J2_127_3477_n987), .CI(DP_OP_425J2_127_3477_n1172), .CO(
        DP_OP_425J2_127_3477_n976), .S(DP_OP_425J2_127_3477_n977) );
  FADDX1_HVT DP_OP_425J2_127_3477_U644 ( .A(DP_OP_425J2_127_3477_n985), .B(
        DP_OP_425J2_127_3477_n1170), .CI(DP_OP_425J2_127_3477_n983), .CO(
        DP_OP_425J2_127_3477_n974), .S(DP_OP_425J2_127_3477_n975) );
  FADDX1_HVT DP_OP_425J2_127_3477_U643 ( .A(DP_OP_425J2_127_3477_n981), .B(
        DP_OP_425J2_127_3477_n1168), .CI(DP_OP_425J2_127_3477_n979), .CO(
        DP_OP_425J2_127_3477_n972), .S(DP_OP_425J2_127_3477_n973) );
  FADDX1_HVT DP_OP_425J2_127_3477_U642 ( .A(DP_OP_425J2_127_3477_n1166), .B(
        DP_OP_425J2_127_3477_n977), .CI(DP_OP_425J2_127_3477_n975), .CO(
        DP_OP_425J2_127_3477_n970), .S(DP_OP_425J2_127_3477_n971) );
  FADDX1_HVT DP_OP_425J2_127_3477_U641 ( .A(DP_OP_425J2_127_3477_n1164), .B(
        DP_OP_425J2_127_3477_n973), .CI(DP_OP_425J2_127_3477_n1162), .CO(
        DP_OP_425J2_127_3477_n968), .S(DP_OP_425J2_127_3477_n969) );
  FADDX1_HVT DP_OP_425J2_127_3477_U640 ( .A(DP_OP_425J2_127_3477_n2978), .B(
        DP_OP_425J2_127_3477_n1923), .CI(DP_OP_425J2_127_3477_n1879), .CO(
        DP_OP_425J2_127_3477_n966), .S(DP_OP_425J2_127_3477_n967) );
  FADDX1_HVT DP_OP_425J2_127_3477_U639 ( .A(DP_OP_425J2_127_3477_n2803), .B(
        DP_OP_425J2_127_3477_n2120), .CI(DP_OP_425J2_127_3477_n2384), .CO(
        DP_OP_425J2_127_3477_n964), .S(DP_OP_425J2_127_3477_n965) );
  FADDX1_HVT DP_OP_425J2_127_3477_U638 ( .A(DP_OP_425J2_127_3477_n2011), .B(
        DP_OP_425J2_127_3477_n2428), .CI(DP_OP_425J2_127_3477_n1988), .CO(
        DP_OP_425J2_127_3477_n962), .S(DP_OP_425J2_127_3477_n963) );
  FADDX1_HVT DP_OP_425J2_127_3477_U637 ( .A(DP_OP_425J2_127_3477_n2319), .B(
        DP_OP_425J2_127_3477_n1944), .CI(DP_OP_425J2_127_3477_n2912), .CO(
        DP_OP_425J2_127_3477_n960), .S(DP_OP_425J2_127_3477_n961) );
  FADDX1_HVT DP_OP_425J2_127_3477_U636 ( .A(DP_OP_425J2_127_3477_n2275), .B(
        DP_OP_425J2_127_3477_n2252), .CI(DP_OP_425J2_127_3477_n2604), .CO(
        DP_OP_425J2_127_3477_n958), .S(DP_OP_425J2_127_3477_n959) );
  FADDX1_HVT DP_OP_425J2_127_3477_U635 ( .A(DP_OP_425J2_127_3477_n2187), .B(
        DP_OP_425J2_127_3477_n2296), .CI(DP_OP_425J2_127_3477_n2956), .CO(
        DP_OP_425J2_127_3477_n956), .S(DP_OP_425J2_127_3477_n957) );
  FADDX1_HVT DP_OP_425J2_127_3477_U634 ( .A(DP_OP_425J2_127_3477_n1967), .B(
        DP_OP_425J2_127_3477_n2032), .CI(DP_OP_425J2_127_3477_n2472), .CO(
        DP_OP_425J2_127_3477_n954), .S(DP_OP_425J2_127_3477_n955) );
  FADDX1_HVT DP_OP_425J2_127_3477_U633 ( .A(DP_OP_425J2_127_3477_n2055), .B(
        DP_OP_425J2_127_3477_n2736), .CI(DP_OP_425J2_127_3477_n2780), .CO(
        DP_OP_425J2_127_3477_n952), .S(DP_OP_425J2_127_3477_n953) );
  FADDX1_HVT DP_OP_425J2_127_3477_U632 ( .A(DP_OP_425J2_127_3477_n2143), .B(
        DP_OP_425J2_127_3477_n2692), .CI(DP_OP_425J2_127_3477_n2560), .CO(
        DP_OP_425J2_127_3477_n950), .S(DP_OP_425J2_127_3477_n951) );
  FADDX1_HVT DP_OP_425J2_127_3477_U631 ( .A(DP_OP_425J2_127_3477_n2495), .B(
        DP_OP_425J2_127_3477_n2340), .CI(DP_OP_425J2_127_3477_n2824), .CO(
        DP_OP_425J2_127_3477_n948), .S(DP_OP_425J2_127_3477_n949) );
  FADDX1_HVT DP_OP_425J2_127_3477_U630 ( .A(DP_OP_425J2_127_3477_n2891), .B(
        DP_OP_425J2_127_3477_n2164), .CI(DP_OP_425J2_127_3477_n2076), .CO(
        DP_OP_425J2_127_3477_n946), .S(DP_OP_425J2_127_3477_n947) );
  FADDX1_HVT DP_OP_425J2_127_3477_U629 ( .A(DP_OP_425J2_127_3477_n2627), .B(
        DP_OP_425J2_127_3477_n2868), .CI(DP_OP_425J2_127_3477_n2516), .CO(
        DP_OP_425J2_127_3477_n944), .S(DP_OP_425J2_127_3477_n945) );
  FADDX1_HVT DP_OP_425J2_127_3477_U628 ( .A(DP_OP_425J2_127_3477_n2407), .B(
        DP_OP_425J2_127_3477_n2998), .CI(DP_OP_425J2_127_3477_n2208), .CO(
        DP_OP_425J2_127_3477_n942), .S(DP_OP_425J2_127_3477_n943) );
  FADDX1_HVT DP_OP_425J2_127_3477_U627 ( .A(DP_OP_425J2_127_3477_n2099), .B(
        DP_OP_425J2_127_3477_n2363), .CI(DP_OP_425J2_127_3477_n2648), .CO(
        DP_OP_425J2_127_3477_n940), .S(DP_OP_425J2_127_3477_n941) );
  FADDX1_HVT DP_OP_425J2_127_3477_U626 ( .A(DP_OP_425J2_127_3477_n2715), .B(
        DP_OP_425J2_127_3477_n2759), .CI(DP_OP_425J2_127_3477_n2847), .CO(
        DP_OP_425J2_127_3477_n938), .S(DP_OP_425J2_127_3477_n939) );
  FADDX1_HVT DP_OP_425J2_127_3477_U625 ( .A(DP_OP_425J2_127_3477_n2451), .B(
        DP_OP_425J2_127_3477_n2539), .CI(DP_OP_425J2_127_3477_n2935), .CO(
        DP_OP_425J2_127_3477_n936), .S(DP_OP_425J2_127_3477_n937) );
  FADDX1_HVT DP_OP_425J2_127_3477_U624 ( .A(DP_OP_425J2_127_3477_n2583), .B(
        DP_OP_425J2_127_3477_n2231), .CI(DP_OP_425J2_127_3477_n2671), .CO(
        DP_OP_425J2_127_3477_n934), .S(DP_OP_425J2_127_3477_n935) );
  FADDX1_HVT DP_OP_425J2_127_3477_U623 ( .A(DP_OP_425J2_127_3477_n2991), .B(
        DP_OP_425J2_127_3477_n1937), .CI(DP_OP_425J2_127_3477_n1930), .CO(
        DP_OP_425J2_127_3477_n932), .S(DP_OP_425J2_127_3477_n933) );
  FADDX1_HVT DP_OP_425J2_127_3477_U622 ( .A(DP_OP_425J2_127_3477_n2984), .B(
        DP_OP_425J2_127_3477_n2949), .CI(DP_OP_425J2_127_3477_n2942), .CO(
        DP_OP_425J2_127_3477_n930), .S(DP_OP_425J2_127_3477_n931) );
  FADDX1_HVT DP_OP_425J2_127_3477_U621 ( .A(DP_OP_425J2_127_3477_n2465), .B(
        DP_OP_425J2_127_3477_n2905), .CI(DP_OP_425J2_127_3477_n2898), .CO(
        DP_OP_425J2_127_3477_n928), .S(DP_OP_425J2_127_3477_n929) );
  FADDX1_HVT DP_OP_425J2_127_3477_U620 ( .A(DP_OP_425J2_127_3477_n2861), .B(
        DP_OP_425J2_127_3477_n1974), .CI(DP_OP_425J2_127_3477_n1981), .CO(
        DP_OP_425J2_127_3477_n926), .S(DP_OP_425J2_127_3477_n927) );
  FADDX1_HVT DP_OP_425J2_127_3477_U619 ( .A(DP_OP_425J2_127_3477_n2854), .B(
        DP_OP_425J2_127_3477_n2018), .CI(DP_OP_425J2_127_3477_n2025), .CO(
        DP_OP_425J2_127_3477_n924), .S(DP_OP_425J2_127_3477_n925) );
  FADDX1_HVT DP_OP_425J2_127_3477_U618 ( .A(DP_OP_425J2_127_3477_n2817), .B(
        DP_OP_425J2_127_3477_n2062), .CI(DP_OP_425J2_127_3477_n2069), .CO(
        DP_OP_425J2_127_3477_n922), .S(DP_OP_425J2_127_3477_n923) );
  FADDX1_HVT DP_OP_425J2_127_3477_U617 ( .A(DP_OP_425J2_127_3477_n2810), .B(
        DP_OP_425J2_127_3477_n2106), .CI(DP_OP_425J2_127_3477_n2113), .CO(
        DP_OP_425J2_127_3477_n920), .S(DP_OP_425J2_127_3477_n921) );
  FADDX1_HVT DP_OP_425J2_127_3477_U616 ( .A(DP_OP_425J2_127_3477_n2773), .B(
        DP_OP_425J2_127_3477_n2150), .CI(DP_OP_425J2_127_3477_n2157), .CO(
        DP_OP_425J2_127_3477_n918), .S(DP_OP_425J2_127_3477_n919) );
  FADDX1_HVT DP_OP_425J2_127_3477_U615 ( .A(DP_OP_425J2_127_3477_n2766), .B(
        DP_OP_425J2_127_3477_n2194), .CI(DP_OP_425J2_127_3477_n2201), .CO(
        DP_OP_425J2_127_3477_n916), .S(DP_OP_425J2_127_3477_n917) );
  FADDX1_HVT DP_OP_425J2_127_3477_U614 ( .A(DP_OP_425J2_127_3477_n2729), .B(
        DP_OP_425J2_127_3477_n2238), .CI(DP_OP_425J2_127_3477_n2245), .CO(
        DP_OP_425J2_127_3477_n914), .S(DP_OP_425J2_127_3477_n915) );
  FADDX1_HVT DP_OP_425J2_127_3477_U613 ( .A(DP_OP_425J2_127_3477_n2722), .B(
        DP_OP_425J2_127_3477_n2282), .CI(DP_OP_425J2_127_3477_n2289), .CO(
        DP_OP_425J2_127_3477_n912), .S(DP_OP_425J2_127_3477_n913) );
  FADDX1_HVT DP_OP_425J2_127_3477_U612 ( .A(DP_OP_425J2_127_3477_n2685), .B(
        DP_OP_425J2_127_3477_n2326), .CI(DP_OP_425J2_127_3477_n2333), .CO(
        DP_OP_425J2_127_3477_n910), .S(DP_OP_425J2_127_3477_n911) );
  FADDX1_HVT DP_OP_425J2_127_3477_U611 ( .A(DP_OP_425J2_127_3477_n2678), .B(
        DP_OP_425J2_127_3477_n2370), .CI(DP_OP_425J2_127_3477_n2377), .CO(
        DP_OP_425J2_127_3477_n908), .S(DP_OP_425J2_127_3477_n909) );
  FADDX1_HVT DP_OP_425J2_127_3477_U610 ( .A(DP_OP_425J2_127_3477_n2641), .B(
        DP_OP_425J2_127_3477_n2414), .CI(DP_OP_425J2_127_3477_n2421), .CO(
        DP_OP_425J2_127_3477_n906), .S(DP_OP_425J2_127_3477_n907) );
  FADDX1_HVT DP_OP_425J2_127_3477_U609 ( .A(DP_OP_425J2_127_3477_n2634), .B(
        DP_OP_425J2_127_3477_n2458), .CI(DP_OP_425J2_127_3477_n2502), .CO(
        DP_OP_425J2_127_3477_n904), .S(DP_OP_425J2_127_3477_n905) );
  FADDX1_HVT DP_OP_425J2_127_3477_U608 ( .A(DP_OP_425J2_127_3477_n2597), .B(
        DP_OP_425J2_127_3477_n2509), .CI(DP_OP_425J2_127_3477_n2546), .CO(
        DP_OP_425J2_127_3477_n902), .S(DP_OP_425J2_127_3477_n903) );
  FADDX1_HVT DP_OP_425J2_127_3477_U607 ( .A(DP_OP_425J2_127_3477_n2590), .B(
        DP_OP_425J2_127_3477_n2553), .CI(DP_OP_425J2_127_3477_n1160), .CO(
        DP_OP_425J2_127_3477_n900), .S(DP_OP_425J2_127_3477_n901) );
  FADDX1_HVT DP_OP_425J2_127_3477_U606 ( .A(DP_OP_425J2_127_3477_n1148), .B(
        DP_OP_425J2_127_3477_n1144), .CI(DP_OP_425J2_127_3477_n1158), .CO(
        DP_OP_425J2_127_3477_n898), .S(DP_OP_425J2_127_3477_n899) );
  FADDX1_HVT DP_OP_425J2_127_3477_U605 ( .A(DP_OP_425J2_127_3477_n1156), .B(
        DP_OP_425J2_127_3477_n1146), .CI(DP_OP_425J2_127_3477_n1154), .CO(
        DP_OP_425J2_127_3477_n896), .S(DP_OP_425J2_127_3477_n897) );
  FADDX1_HVT DP_OP_425J2_127_3477_U604 ( .A(DP_OP_425J2_127_3477_n1152), .B(
        DP_OP_425J2_127_3477_n1150), .CI(DP_OP_425J2_127_3477_n1120), .CO(
        DP_OP_425J2_127_3477_n894), .S(DP_OP_425J2_127_3477_n895) );
  FADDX1_HVT DP_OP_425J2_127_3477_U603 ( .A(DP_OP_425J2_127_3477_n1118), .B(
        DP_OP_425J2_127_3477_n1094), .CI(DP_OP_425J2_127_3477_n1142), .CO(
        DP_OP_425J2_127_3477_n892), .S(DP_OP_425J2_127_3477_n893) );
  FADDX1_HVT DP_OP_425J2_127_3477_U602 ( .A(DP_OP_425J2_127_3477_n1116), .B(
        DP_OP_425J2_127_3477_n1140), .CI(DP_OP_425J2_127_3477_n1138), .CO(
        DP_OP_425J2_127_3477_n890), .S(DP_OP_425J2_127_3477_n891) );
  FADDX1_HVT DP_OP_425J2_127_3477_U601 ( .A(DP_OP_425J2_127_3477_n1110), .B(
        DP_OP_425J2_127_3477_n1136), .CI(DP_OP_425J2_127_3477_n1134), .CO(
        DP_OP_425J2_127_3477_n888), .S(DP_OP_425J2_127_3477_n889) );
  FADDX1_HVT DP_OP_425J2_127_3477_U600 ( .A(DP_OP_425J2_127_3477_n1132), .B(
        DP_OP_425J2_127_3477_n1130), .CI(DP_OP_425J2_127_3477_n1128), .CO(
        DP_OP_425J2_127_3477_n886), .S(DP_OP_425J2_127_3477_n887) );
  FADDX1_HVT DP_OP_425J2_127_3477_U599 ( .A(DP_OP_425J2_127_3477_n1100), .B(
        DP_OP_425J2_127_3477_n1126), .CI(DP_OP_425J2_127_3477_n1124), .CO(
        DP_OP_425J2_127_3477_n884), .S(DP_OP_425J2_127_3477_n885) );
  FADDX1_HVT DP_OP_425J2_127_3477_U598 ( .A(DP_OP_425J2_127_3477_n1106), .B(
        DP_OP_425J2_127_3477_n1122), .CI(DP_OP_425J2_127_3477_n1114), .CO(
        DP_OP_425J2_127_3477_n882), .S(DP_OP_425J2_127_3477_n883) );
  FADDX1_HVT DP_OP_425J2_127_3477_U597 ( .A(DP_OP_425J2_127_3477_n1098), .B(
        DP_OP_425J2_127_3477_n1112), .CI(DP_OP_425J2_127_3477_n1108), .CO(
        DP_OP_425J2_127_3477_n880), .S(DP_OP_425J2_127_3477_n881) );
  FADDX1_HVT DP_OP_425J2_127_3477_U596 ( .A(DP_OP_425J2_127_3477_n1102), .B(
        DP_OP_425J2_127_3477_n1096), .CI(DP_OP_425J2_127_3477_n1104), .CO(
        DP_OP_425J2_127_3477_n878), .S(DP_OP_425J2_127_3477_n879) );
  FADDX1_HVT DP_OP_425J2_127_3477_U595 ( .A(DP_OP_425J2_127_3477_n967), .B(
        DP_OP_425J2_127_3477_n953), .CI(DP_OP_425J2_127_3477_n955), .CO(
        DP_OP_425J2_127_3477_n876), .S(DP_OP_425J2_127_3477_n877) );
  FADDX1_HVT DP_OP_425J2_127_3477_U594 ( .A(DP_OP_425J2_127_3477_n959), .B(
        DP_OP_425J2_127_3477_n937), .CI(DP_OP_425J2_127_3477_n935), .CO(
        DP_OP_425J2_127_3477_n874), .S(DP_OP_425J2_127_3477_n875) );
  FADDX1_HVT DP_OP_425J2_127_3477_U593 ( .A(DP_OP_425J2_127_3477_n951), .B(
        DP_OP_425J2_127_3477_n949), .CI(DP_OP_425J2_127_3477_n945), .CO(
        DP_OP_425J2_127_3477_n872), .S(DP_OP_425J2_127_3477_n873) );
  FADDX1_HVT DP_OP_425J2_127_3477_U592 ( .A(DP_OP_425J2_127_3477_n957), .B(
        DP_OP_425J2_127_3477_n939), .CI(DP_OP_425J2_127_3477_n943), .CO(
        DP_OP_425J2_127_3477_n870), .S(DP_OP_425J2_127_3477_n871) );
  FADDX1_HVT DP_OP_425J2_127_3477_U591 ( .A(DP_OP_425J2_127_3477_n947), .B(
        DP_OP_425J2_127_3477_n965), .CI(DP_OP_425J2_127_3477_n961), .CO(
        DP_OP_425J2_127_3477_n868), .S(DP_OP_425J2_127_3477_n869) );
  FADDX1_HVT DP_OP_425J2_127_3477_U590 ( .A(DP_OP_425J2_127_3477_n941), .B(
        DP_OP_425J2_127_3477_n963), .CI(DP_OP_425J2_127_3477_n923), .CO(
        DP_OP_425J2_127_3477_n866), .S(DP_OP_425J2_127_3477_n867) );
  FADDX1_HVT DP_OP_425J2_127_3477_U589 ( .A(DP_OP_425J2_127_3477_n925), .B(
        DP_OP_425J2_127_3477_n907), .CI(DP_OP_425J2_127_3477_n901), .CO(
        DP_OP_425J2_127_3477_n864), .S(DP_OP_425J2_127_3477_n865) );
  FADDX1_HVT DP_OP_425J2_127_3477_U588 ( .A(DP_OP_425J2_127_3477_n927), .B(
        DP_OP_425J2_127_3477_n903), .CI(DP_OP_425J2_127_3477_n919), .CO(
        DP_OP_425J2_127_3477_n862), .S(DP_OP_425J2_127_3477_n863) );
  FADDX1_HVT DP_OP_425J2_127_3477_U587 ( .A(DP_OP_425J2_127_3477_n917), .B(
        DP_OP_425J2_127_3477_n915), .CI(DP_OP_425J2_127_3477_n905), .CO(
        DP_OP_425J2_127_3477_n860), .S(DP_OP_425J2_127_3477_n861) );
  FADDX1_HVT DP_OP_425J2_127_3477_U586 ( .A(DP_OP_425J2_127_3477_n921), .B(
        DP_OP_425J2_127_3477_n909), .CI(DP_OP_425J2_127_3477_n911), .CO(
        DP_OP_425J2_127_3477_n858), .S(DP_OP_425J2_127_3477_n859) );
  FADDX1_HVT DP_OP_425J2_127_3477_U585 ( .A(DP_OP_425J2_127_3477_n929), .B(
        DP_OP_425J2_127_3477_n933), .CI(DP_OP_425J2_127_3477_n931), .CO(
        DP_OP_425J2_127_3477_n856), .S(DP_OP_425J2_127_3477_n857) );
  FADDX1_HVT DP_OP_425J2_127_3477_U584 ( .A(DP_OP_425J2_127_3477_n913), .B(
        DP_OP_425J2_127_3477_n1092), .CI(DP_OP_425J2_127_3477_n1090), .CO(
        DP_OP_425J2_127_3477_n854), .S(DP_OP_425J2_127_3477_n855) );
  FADDX1_HVT DP_OP_425J2_127_3477_U583 ( .A(DP_OP_425J2_127_3477_n1088), .B(
        DP_OP_425J2_127_3477_n1086), .CI(DP_OP_425J2_127_3477_n1072), .CO(
        DP_OP_425J2_127_3477_n852), .S(DP_OP_425J2_127_3477_n853) );
  FADDX1_HVT DP_OP_425J2_127_3477_U582 ( .A(DP_OP_425J2_127_3477_n1084), .B(
        DP_OP_425J2_127_3477_n1082), .CI(DP_OP_425J2_127_3477_n1070), .CO(
        DP_OP_425J2_127_3477_n850), .S(DP_OP_425J2_127_3477_n851) );
  FADDX1_HVT DP_OP_425J2_127_3477_U581 ( .A(DP_OP_425J2_127_3477_n1080), .B(
        DP_OP_425J2_127_3477_n1074), .CI(DP_OP_425J2_127_3477_n1076), .CO(
        DP_OP_425J2_127_3477_n848), .S(DP_OP_425J2_127_3477_n849) );
  FADDX1_HVT DP_OP_425J2_127_3477_U580 ( .A(DP_OP_425J2_127_3477_n1078), .B(
        DP_OP_425J2_127_3477_n1068), .CI(DP_OP_425J2_127_3477_n1066), .CO(
        DP_OP_425J2_127_3477_n846), .S(DP_OP_425J2_127_3477_n847) );
  FADDX1_HVT DP_OP_425J2_127_3477_U579 ( .A(DP_OP_425J2_127_3477_n899), .B(
        DP_OP_425J2_127_3477_n895), .CI(DP_OP_425J2_127_3477_n1064), .CO(
        DP_OP_425J2_127_3477_n844), .S(DP_OP_425J2_127_3477_n845) );
  FADDX1_HVT DP_OP_425J2_127_3477_U578 ( .A(DP_OP_425J2_127_3477_n897), .B(
        DP_OP_425J2_127_3477_n1052), .CI(DP_OP_425J2_127_3477_n1050), .CO(
        DP_OP_425J2_127_3477_n842), .S(DP_OP_425J2_127_3477_n843) );
  FADDX1_HVT DP_OP_425J2_127_3477_U577 ( .A(DP_OP_425J2_127_3477_n1058), .B(
        DP_OP_425J2_127_3477_n893), .CI(DP_OP_425J2_127_3477_n1048), .CO(
        DP_OP_425J2_127_3477_n840), .S(DP_OP_425J2_127_3477_n841) );
  FADDX1_HVT DP_OP_425J2_127_3477_U576 ( .A(DP_OP_425J2_127_3477_n1056), .B(
        DP_OP_425J2_127_3477_n889), .CI(DP_OP_425J2_127_3477_n879), .CO(
        DP_OP_425J2_127_3477_n838), .S(DP_OP_425J2_127_3477_n839) );
  FADDX1_HVT DP_OP_425J2_127_3477_U575 ( .A(DP_OP_425J2_127_3477_n1062), .B(
        DP_OP_425J2_127_3477_n885), .CI(DP_OP_425J2_127_3477_n887), .CO(
        DP_OP_425J2_127_3477_n836), .S(DP_OP_425J2_127_3477_n837) );
  FADDX1_HVT DP_OP_425J2_127_3477_U574 ( .A(DP_OP_425J2_127_3477_n1060), .B(
        DP_OP_425J2_127_3477_n881), .CI(DP_OP_425J2_127_3477_n883), .CO(
        DP_OP_425J2_127_3477_n834), .S(DP_OP_425J2_127_3477_n835) );
  FADDX1_HVT DP_OP_425J2_127_3477_U573 ( .A(DP_OP_425J2_127_3477_n1054), .B(
        DP_OP_425J2_127_3477_n891), .CI(DP_OP_425J2_127_3477_n877), .CO(
        DP_OP_425J2_127_3477_n832), .S(DP_OP_425J2_127_3477_n833) );
  FADDX1_HVT DP_OP_425J2_127_3477_U572 ( .A(DP_OP_425J2_127_3477_n871), .B(
        DP_OP_425J2_127_3477_n875), .CI(DP_OP_425J2_127_3477_n867), .CO(
        DP_OP_425J2_127_3477_n830), .S(DP_OP_425J2_127_3477_n831) );
  FADDX1_HVT DP_OP_425J2_127_3477_U571 ( .A(DP_OP_425J2_127_3477_n869), .B(
        DP_OP_425J2_127_3477_n873), .CI(DP_OP_425J2_127_3477_n861), .CO(
        DP_OP_425J2_127_3477_n828), .S(DP_OP_425J2_127_3477_n829) );
  FADDX1_HVT DP_OP_425J2_127_3477_U570 ( .A(DP_OP_425J2_127_3477_n859), .B(
        DP_OP_425J2_127_3477_n865), .CI(DP_OP_425J2_127_3477_n1046), .CO(
        DP_OP_425J2_127_3477_n826), .S(DP_OP_425J2_127_3477_n827) );
  FADDX1_HVT DP_OP_425J2_127_3477_U569 ( .A(DP_OP_425J2_127_3477_n857), .B(
        DP_OP_425J2_127_3477_n863), .CI(DP_OP_425J2_127_3477_n1042), .CO(
        DP_OP_425J2_127_3477_n824), .S(DP_OP_425J2_127_3477_n825) );
  FADDX1_HVT DP_OP_425J2_127_3477_U568 ( .A(DP_OP_425J2_127_3477_n1044), .B(
        DP_OP_425J2_127_3477_n1040), .CI(DP_OP_425J2_127_3477_n855), .CO(
        DP_OP_425J2_127_3477_n822), .S(DP_OP_425J2_127_3477_n823) );
  FADDX1_HVT DP_OP_425J2_127_3477_U567 ( .A(DP_OP_425J2_127_3477_n1038), .B(
        DP_OP_425J2_127_3477_n1036), .CI(DP_OP_425J2_127_3477_n853), .CO(
        DP_OP_425J2_127_3477_n820), .S(DP_OP_425J2_127_3477_n821) );
  FADDX1_HVT DP_OP_425J2_127_3477_U566 ( .A(DP_OP_425J2_127_3477_n1034), .B(
        DP_OP_425J2_127_3477_n851), .CI(DP_OP_425J2_127_3477_n849), .CO(
        DP_OP_425J2_127_3477_n818), .S(DP_OP_425J2_127_3477_n819) );
  FADDX1_HVT DP_OP_425J2_127_3477_U565 ( .A(DP_OP_425J2_127_3477_n1032), .B(
        DP_OP_425J2_127_3477_n1026), .CI(DP_OP_425J2_127_3477_n1028), .CO(
        DP_OP_425J2_127_3477_n816), .S(DP_OP_425J2_127_3477_n817) );
  FADDX1_HVT DP_OP_425J2_127_3477_U564 ( .A(DP_OP_425J2_127_3477_n1030), .B(
        DP_OP_425J2_127_3477_n847), .CI(DP_OP_425J2_127_3477_n1024), .CO(
        DP_OP_425J2_127_3477_n814), .S(DP_OP_425J2_127_3477_n815) );
  FADDX1_HVT DP_OP_425J2_127_3477_U563 ( .A(DP_OP_425J2_127_3477_n845), .B(
        DP_OP_425J2_127_3477_n1022), .CI(DP_OP_425J2_127_3477_n843), .CO(
        DP_OP_425J2_127_3477_n812), .S(DP_OP_425J2_127_3477_n813) );
  FADDX1_HVT DP_OP_425J2_127_3477_U562 ( .A(DP_OP_425J2_127_3477_n1020), .B(
        DP_OP_425J2_127_3477_n837), .CI(DP_OP_425J2_127_3477_n833), .CO(
        DP_OP_425J2_127_3477_n810), .S(DP_OP_425J2_127_3477_n811) );
  FADDX1_HVT DP_OP_425J2_127_3477_U561 ( .A(DP_OP_425J2_127_3477_n1018), .B(
        DP_OP_425J2_127_3477_n841), .CI(DP_OP_425J2_127_3477_n839), .CO(
        DP_OP_425J2_127_3477_n808), .S(DP_OP_425J2_127_3477_n809) );
  FADDX1_HVT DP_OP_425J2_127_3477_U560 ( .A(DP_OP_425J2_127_3477_n835), .B(
        DP_OP_425J2_127_3477_n1016), .CI(DP_OP_425J2_127_3477_n831), .CO(
        DP_OP_425J2_127_3477_n806), .S(DP_OP_425J2_127_3477_n807) );
  FADDX1_HVT DP_OP_425J2_127_3477_U559 ( .A(DP_OP_425J2_127_3477_n829), .B(
        DP_OP_425J2_127_3477_n1014), .CI(DP_OP_425J2_127_3477_n827), .CO(
        DP_OP_425J2_127_3477_n804), .S(DP_OP_425J2_127_3477_n805) );
  FADDX1_HVT DP_OP_425J2_127_3477_U558 ( .A(DP_OP_425J2_127_3477_n825), .B(
        DP_OP_425J2_127_3477_n1012), .CI(DP_OP_425J2_127_3477_n1008), .CO(
        DP_OP_425J2_127_3477_n802), .S(DP_OP_425J2_127_3477_n803) );
  FADDX1_HVT DP_OP_425J2_127_3477_U557 ( .A(DP_OP_425J2_127_3477_n1010), .B(
        DP_OP_425J2_127_3477_n823), .CI(DP_OP_425J2_127_3477_n1006), .CO(
        DP_OP_425J2_127_3477_n800), .S(DP_OP_425J2_127_3477_n801) );
  FADDX1_HVT DP_OP_425J2_127_3477_U556 ( .A(DP_OP_425J2_127_3477_n821), .B(
        DP_OP_425J2_127_3477_n1004), .CI(DP_OP_425J2_127_3477_n1002), .CO(
        DP_OP_425J2_127_3477_n798), .S(DP_OP_425J2_127_3477_n799) );
  FADDX1_HVT DP_OP_425J2_127_3477_U555 ( .A(DP_OP_425J2_127_3477_n819), .B(
        DP_OP_425J2_127_3477_n1000), .CI(DP_OP_425J2_127_3477_n815), .CO(
        DP_OP_425J2_127_3477_n796), .S(DP_OP_425J2_127_3477_n797) );
  FADDX1_HVT DP_OP_425J2_127_3477_U554 ( .A(DP_OP_425J2_127_3477_n817), .B(
        DP_OP_425J2_127_3477_n998), .CI(DP_OP_425J2_127_3477_n813), .CO(
        DP_OP_425J2_127_3477_n794), .S(DP_OP_425J2_127_3477_n795) );
  FADDX1_HVT DP_OP_425J2_127_3477_U553 ( .A(DP_OP_425J2_127_3477_n996), .B(
        DP_OP_425J2_127_3477_n811), .CI(DP_OP_425J2_127_3477_n807), .CO(
        DP_OP_425J2_127_3477_n792), .S(DP_OP_425J2_127_3477_n793) );
  FADDX1_HVT DP_OP_425J2_127_3477_U552 ( .A(DP_OP_425J2_127_3477_n809), .B(
        DP_OP_425J2_127_3477_n994), .CI(DP_OP_425J2_127_3477_n805), .CO(
        DP_OP_425J2_127_3477_n790), .S(DP_OP_425J2_127_3477_n791) );
  FADDX1_HVT DP_OP_425J2_127_3477_U551 ( .A(DP_OP_425J2_127_3477_n992), .B(
        DP_OP_425J2_127_3477_n803), .CI(DP_OP_425J2_127_3477_n990), .CO(
        DP_OP_425J2_127_3477_n788), .S(DP_OP_425J2_127_3477_n789) );
  FADDX1_HVT DP_OP_425J2_127_3477_U550 ( .A(DP_OP_425J2_127_3477_n801), .B(
        DP_OP_425J2_127_3477_n988), .CI(DP_OP_425J2_127_3477_n799), .CO(
        DP_OP_425J2_127_3477_n786), .S(DP_OP_425J2_127_3477_n787) );
  FADDX1_HVT DP_OP_425J2_127_3477_U549 ( .A(DP_OP_425J2_127_3477_n986), .B(
        DP_OP_425J2_127_3477_n797), .CI(DP_OP_425J2_127_3477_n984), .CO(
        DP_OP_425J2_127_3477_n784), .S(DP_OP_425J2_127_3477_n785) );
  FADDX1_HVT DP_OP_425J2_127_3477_U548 ( .A(DP_OP_425J2_127_3477_n795), .B(
        DP_OP_425J2_127_3477_n793), .CI(DP_OP_425J2_127_3477_n982), .CO(
        DP_OP_425J2_127_3477_n782), .S(DP_OP_425J2_127_3477_n783) );
  FADDX1_HVT DP_OP_425J2_127_3477_U547 ( .A(DP_OP_425J2_127_3477_n791), .B(
        DP_OP_425J2_127_3477_n980), .CI(DP_OP_425J2_127_3477_n789), .CO(
        DP_OP_425J2_127_3477_n780), .S(DP_OP_425J2_127_3477_n781) );
  FADDX1_HVT DP_OP_425J2_127_3477_U546 ( .A(DP_OP_425J2_127_3477_n978), .B(
        DP_OP_425J2_127_3477_n787), .CI(DP_OP_425J2_127_3477_n976), .CO(
        DP_OP_425J2_127_3477_n778), .S(DP_OP_425J2_127_3477_n779) );
  FADDX1_HVT DP_OP_425J2_127_3477_U545 ( .A(DP_OP_425J2_127_3477_n785), .B(
        DP_OP_425J2_127_3477_n974), .CI(DP_OP_425J2_127_3477_n783), .CO(
        DP_OP_425J2_127_3477_n776), .S(DP_OP_425J2_127_3477_n777) );
  FADDX1_HVT DP_OP_425J2_127_3477_U544 ( .A(DP_OP_425J2_127_3477_n781), .B(
        DP_OP_425J2_127_3477_n972), .CI(DP_OP_425J2_127_3477_n779), .CO(
        DP_OP_425J2_127_3477_n774), .S(DP_OP_425J2_127_3477_n775) );
  FADDX1_HVT DP_OP_425J2_127_3477_U543 ( .A(DP_OP_425J2_127_3477_n970), .B(
        DP_OP_425J2_127_3477_n777), .CI(DP_OP_425J2_127_3477_n775), .CO(
        DP_OP_425J2_127_3477_n772), .S(DP_OP_425J2_127_3477_n773) );
  FADDX1_HVT DP_OP_425J2_127_3477_U541 ( .A(DP_OP_425J2_127_3477_n2186), .B(
        DP_OP_425J2_127_3477_n1922), .CI(DP_OP_425J2_127_3477_n1878), .CO(
        DP_OP_425J2_127_3477_n768), .S(DP_OP_425J2_127_3477_n769) );
  FADDX1_HVT DP_OP_425J2_127_3477_U540 ( .A(DP_OP_425J2_127_3477_n2758), .B(
        DP_OP_425J2_127_3477_n1980), .CI(DP_OP_425J2_127_3477_n2244), .CO(
        DP_OP_425J2_127_3477_n766), .S(DP_OP_425J2_127_3477_n767) );
  FADDX1_HVT DP_OP_425J2_127_3477_U539 ( .A(DP_OP_425J2_127_3477_n2230), .B(
        DP_OP_425J2_127_3477_n2990), .CI(DP_OP_425J2_127_3477_n2640), .CO(
        DP_OP_425J2_127_3477_n764), .S(DP_OP_425J2_127_3477_n765) );
  FADDX1_HVT DP_OP_425J2_127_3477_U538 ( .A(DP_OP_425J2_127_3477_n2450), .B(
        DP_OP_425J2_127_3477_n2024), .CI(DP_OP_425J2_127_3477_n2068), .CO(
        DP_OP_425J2_127_3477_n762), .S(DP_OP_425J2_127_3477_n763) );
  FADDX1_HVT DP_OP_425J2_127_3477_U537 ( .A(DP_OP_425J2_127_3477_n2010), .B(
        DP_OP_425J2_127_3477_n2112), .CI(DP_OP_425J2_127_3477_n2156), .CO(
        DP_OP_425J2_127_3477_n760), .S(DP_OP_425J2_127_3477_n761) );
  FADDX1_HVT DP_OP_425J2_127_3477_U536 ( .A(DP_OP_425J2_127_3477_n2714), .B(
        DP_OP_425J2_127_3477_n2816), .CI(DP_OP_425J2_127_3477_n2860), .CO(
        DP_OP_425J2_127_3477_n758), .S(DP_OP_425J2_127_3477_n759) );
  FADDX1_HVT DP_OP_425J2_127_3477_U535 ( .A(DP_OP_425J2_127_3477_n2054), .B(
        DP_OP_425J2_127_3477_n2772), .CI(DP_OP_425J2_127_3477_n2596), .CO(
        DP_OP_425J2_127_3477_n756), .S(DP_OP_425J2_127_3477_n757) );
  FADDX1_HVT DP_OP_425J2_127_3477_U534 ( .A(DP_OP_425J2_127_3477_n2142), .B(
        DP_OP_425J2_127_3477_n2420), .CI(DP_OP_425J2_127_3477_n2948), .CO(
        DP_OP_425J2_127_3477_n754), .S(DP_OP_425J2_127_3477_n755) );
  FADDX1_HVT DP_OP_425J2_127_3477_U533 ( .A(DP_OP_425J2_127_3477_n2670), .B(
        DP_OP_425J2_127_3477_n2904), .CI(DP_OP_425J2_127_3477_n2464), .CO(
        DP_OP_425J2_127_3477_n752), .S(DP_OP_425J2_127_3477_n753) );
  FADDX1_HVT DP_OP_425J2_127_3477_U532 ( .A(DP_OP_425J2_127_3477_n2626), .B(
        DP_OP_425J2_127_3477_n2376), .CI(DP_OP_425J2_127_3477_n2728), .CO(
        DP_OP_425J2_127_3477_n750), .S(DP_OP_425J2_127_3477_n751) );
  FADDX1_HVT DP_OP_425J2_127_3477_U531 ( .A(DP_OP_425J2_127_3477_n2846), .B(
        DP_OP_425J2_127_3477_n2508), .CI(DP_OP_425J2_127_3477_n2332), .CO(
        DP_OP_425J2_127_3477_n748), .S(DP_OP_425J2_127_3477_n749) );
  FADDX1_HVT DP_OP_425J2_127_3477_U530 ( .A(DP_OP_425J2_127_3477_n2318), .B(
        DP_OP_425J2_127_3477_n2288), .CI(DP_OP_425J2_127_3477_n1936), .CO(
        DP_OP_425J2_127_3477_n746), .S(DP_OP_425J2_127_3477_n747) );
  FADDX1_HVT DP_OP_425J2_127_3477_U529 ( .A(DP_OP_425J2_127_3477_n2538), .B(
        DP_OP_425J2_127_3477_n2200), .CI(DP_OP_425J2_127_3477_n2552), .CO(
        DP_OP_425J2_127_3477_n744), .S(DP_OP_425J2_127_3477_n745) );
  FADDX1_HVT DP_OP_425J2_127_3477_U528 ( .A(DP_OP_425J2_127_3477_n2494), .B(
        DP_OP_425J2_127_3477_n2362), .CI(DP_OP_425J2_127_3477_n2684), .CO(
        DP_OP_425J2_127_3477_n742), .S(DP_OP_425J2_127_3477_n743) );
  FADDX1_HVT DP_OP_425J2_127_3477_U527 ( .A(DP_OP_425J2_127_3477_n2802), .B(
        DP_OP_425J2_127_3477_n2098), .CI(DP_OP_425J2_127_3477_n2274), .CO(
        DP_OP_425J2_127_3477_n740), .S(DP_OP_425J2_127_3477_n741) );
  FADDX1_HVT DP_OP_425J2_127_3477_U526 ( .A(DP_OP_425J2_127_3477_n1966), .B(
        DP_OP_425J2_127_3477_n2582), .CI(DP_OP_425J2_127_3477_n2934), .CO(
        DP_OP_425J2_127_3477_n738), .S(DP_OP_425J2_127_3477_n739) );
  FADDX1_HVT DP_OP_425J2_127_3477_U525 ( .A(DP_OP_425J2_127_3477_n2890), .B(
        DP_OP_425J2_127_3477_n2406), .CI(DP_OP_425J2_127_3477_n771), .CO(
        DP_OP_425J2_127_3477_n736), .S(DP_OP_425J2_127_3477_n737) );
  FADDX1_HVT DP_OP_425J2_127_3477_U524 ( .A(DP_OP_425J2_127_3477_n2237), .B(
        DP_OP_425J2_127_3477_n1973), .CI(DP_OP_425J2_127_3477_n1929), .CO(
        DP_OP_425J2_127_3477_n734), .S(DP_OP_425J2_127_3477_n735) );
  FADDX1_HVT DP_OP_425J2_127_3477_U523 ( .A(DP_OP_425J2_127_3477_n2983), .B(
        DP_OP_425J2_127_3477_n2017), .CI(DP_OP_425J2_127_3477_n2061), .CO(
        DP_OP_425J2_127_3477_n732), .S(DP_OP_425J2_127_3477_n733) );
  FADDX1_HVT DP_OP_425J2_127_3477_U522 ( .A(DP_OP_425J2_127_3477_n2941), .B(
        DP_OP_425J2_127_3477_n2105), .CI(DP_OP_425J2_127_3477_n2149), .CO(
        DP_OP_425J2_127_3477_n730), .S(DP_OP_425J2_127_3477_n731) );
  FADDX1_HVT DP_OP_425J2_127_3477_U521 ( .A(DP_OP_425J2_127_3477_n2897), .B(
        DP_OP_425J2_127_3477_n2193), .CI(DP_OP_425J2_127_3477_n2281), .CO(
        DP_OP_425J2_127_3477_n728), .S(DP_OP_425J2_127_3477_n729) );
  FADDX1_HVT DP_OP_425J2_127_3477_U520 ( .A(DP_OP_425J2_127_3477_n2853), .B(
        DP_OP_425J2_127_3477_n2325), .CI(DP_OP_425J2_127_3477_n2369), .CO(
        DP_OP_425J2_127_3477_n726), .S(DP_OP_425J2_127_3477_n727) );
  FADDX1_HVT DP_OP_425J2_127_3477_U519 ( .A(DP_OP_425J2_127_3477_n2809), .B(
        DP_OP_425J2_127_3477_n2413), .CI(DP_OP_425J2_127_3477_n2457), .CO(
        DP_OP_425J2_127_3477_n724), .S(DP_OP_425J2_127_3477_n725) );
  FADDX1_HVT DP_OP_425J2_127_3477_U518 ( .A(DP_OP_425J2_127_3477_n2765), .B(
        DP_OP_425J2_127_3477_n2501), .CI(DP_OP_425J2_127_3477_n2545), .CO(
        DP_OP_425J2_127_3477_n722), .S(DP_OP_425J2_127_3477_n723) );
  FADDX1_HVT DP_OP_425J2_127_3477_U517 ( .A(DP_OP_425J2_127_3477_n2721), .B(
        DP_OP_425J2_127_3477_n2589), .CI(DP_OP_425J2_127_3477_n2633), .CO(
        DP_OP_425J2_127_3477_n720), .S(DP_OP_425J2_127_3477_n721) );
  FADDX1_HVT DP_OP_425J2_127_3477_U516 ( .A(DP_OP_425J2_127_3477_n2677), .B(
        DP_OP_425J2_127_3477_n966), .CI(DP_OP_425J2_127_3477_n964), .CO(
        DP_OP_425J2_127_3477_n718), .S(DP_OP_425J2_127_3477_n719) );
  FADDX1_HVT DP_OP_425J2_127_3477_U515 ( .A(DP_OP_425J2_127_3477_n962), .B(
        DP_OP_425J2_127_3477_n934), .CI(DP_OP_425J2_127_3477_n936), .CO(
        DP_OP_425J2_127_3477_n716), .S(DP_OP_425J2_127_3477_n717) );
  FADDX1_HVT DP_OP_425J2_127_3477_U514 ( .A(DP_OP_425J2_127_3477_n960), .B(
        DP_OP_425J2_127_3477_n938), .CI(DP_OP_425J2_127_3477_n940), .CO(
        DP_OP_425J2_127_3477_n714), .S(DP_OP_425J2_127_3477_n715) );
  FADDX1_HVT DP_OP_425J2_127_3477_U513 ( .A(DP_OP_425J2_127_3477_n958), .B(
        DP_OP_425J2_127_3477_n942), .CI(DP_OP_425J2_127_3477_n944), .CO(
        DP_OP_425J2_127_3477_n712), .S(DP_OP_425J2_127_3477_n713) );
  FADDX1_HVT DP_OP_425J2_127_3477_U512 ( .A(DP_OP_425J2_127_3477_n950), .B(
        DP_OP_425J2_127_3477_n956), .CI(DP_OP_425J2_127_3477_n946), .CO(
        DP_OP_425J2_127_3477_n710), .S(DP_OP_425J2_127_3477_n711) );
  FADDX1_HVT DP_OP_425J2_127_3477_U511 ( .A(DP_OP_425J2_127_3477_n948), .B(
        DP_OP_425J2_127_3477_n952), .CI(DP_OP_425J2_127_3477_n954), .CO(
        DP_OP_425J2_127_3477_n708), .S(DP_OP_425J2_127_3477_n709) );
  FADDX1_HVT DP_OP_425J2_127_3477_U510 ( .A(DP_OP_425J2_127_3477_n932), .B(
        DP_OP_425J2_127_3477_n930), .CI(DP_OP_425J2_127_3477_n900), .CO(
        DP_OP_425J2_127_3477_n706), .S(DP_OP_425J2_127_3477_n707) );
  FADDX1_HVT DP_OP_425J2_127_3477_U509 ( .A(DP_OP_425J2_127_3477_n914), .B(
        DP_OP_425J2_127_3477_n902), .CI(DP_OP_425J2_127_3477_n904), .CO(
        DP_OP_425J2_127_3477_n704), .S(DP_OP_425J2_127_3477_n705) );
  FADDX1_HVT DP_OP_425J2_127_3477_U508 ( .A(DP_OP_425J2_127_3477_n912), .B(
        DP_OP_425J2_127_3477_n906), .CI(DP_OP_425J2_127_3477_n908), .CO(
        DP_OP_425J2_127_3477_n702), .S(DP_OP_425J2_127_3477_n703) );
  FADDX1_HVT DP_OP_425J2_127_3477_U507 ( .A(DP_OP_425J2_127_3477_n910), .B(
        DP_OP_425J2_127_3477_n928), .CI(DP_OP_425J2_127_3477_n926), .CO(
        DP_OP_425J2_127_3477_n700), .S(DP_OP_425J2_127_3477_n701) );
  FADDX1_HVT DP_OP_425J2_127_3477_U506 ( .A(DP_OP_425J2_127_3477_n920), .B(
        DP_OP_425J2_127_3477_n916), .CI(DP_OP_425J2_127_3477_n918), .CO(
        DP_OP_425J2_127_3477_n698), .S(DP_OP_425J2_127_3477_n699) );
  FADDX1_HVT DP_OP_425J2_127_3477_U505 ( .A(DP_OP_425J2_127_3477_n924), .B(
        DP_OP_425J2_127_3477_n922), .CI(DP_OP_425J2_127_3477_n763), .CO(
        DP_OP_425J2_127_3477_n696), .S(DP_OP_425J2_127_3477_n697) );
  FADDX1_HVT DP_OP_425J2_127_3477_U504 ( .A(DP_OP_425J2_127_3477_n759), .B(
        DP_OP_425J2_127_3477_n755), .CI(DP_OP_425J2_127_3477_n737), .CO(
        DP_OP_425J2_127_3477_n694), .S(DP_OP_425J2_127_3477_n695) );
  FADDX1_HVT DP_OP_425J2_127_3477_U503 ( .A(DP_OP_425J2_127_3477_n761), .B(
        DP_OP_425J2_127_3477_n743), .CI(DP_OP_425J2_127_3477_n741), .CO(
        DP_OP_425J2_127_3477_n692), .S(DP_OP_425J2_127_3477_n693) );
  FADDX1_HVT DP_OP_425J2_127_3477_U502 ( .A(DP_OP_425J2_127_3477_n753), .B(
        DP_OP_425J2_127_3477_n757), .CI(DP_OP_425J2_127_3477_n749), .CO(
        DP_OP_425J2_127_3477_n690), .S(DP_OP_425J2_127_3477_n691) );
  FADDX1_HVT DP_OP_425J2_127_3477_U501 ( .A(DP_OP_425J2_127_3477_n765), .B(
        DP_OP_425J2_127_3477_n745), .CI(DP_OP_425J2_127_3477_n739), .CO(
        DP_OP_425J2_127_3477_n688), .S(DP_OP_425J2_127_3477_n689) );
  FADDX1_HVT DP_OP_425J2_127_3477_U500 ( .A(DP_OP_425J2_127_3477_n747), .B(
        DP_OP_425J2_127_3477_n769), .CI(DP_OP_425J2_127_3477_n767), .CO(
        DP_OP_425J2_127_3477_n686), .S(DP_OP_425J2_127_3477_n687) );
  FADDX1_HVT DP_OP_425J2_127_3477_U499 ( .A(DP_OP_425J2_127_3477_n751), .B(
        DP_OP_425J2_127_3477_n731), .CI(DP_OP_425J2_127_3477_n727), .CO(
        DP_OP_425J2_127_3477_n684), .S(DP_OP_425J2_127_3477_n685) );
  FADDX1_HVT DP_OP_425J2_127_3477_U498 ( .A(DP_OP_425J2_127_3477_n723), .B(
        DP_OP_425J2_127_3477_n721), .CI(DP_OP_425J2_127_3477_n733), .CO(
        DP_OP_425J2_127_3477_n682), .S(DP_OP_425J2_127_3477_n683) );
  FADDX1_HVT DP_OP_425J2_127_3477_U497 ( .A(DP_OP_425J2_127_3477_n729), .B(
        DP_OP_425J2_127_3477_n725), .CI(DP_OP_425J2_127_3477_n735), .CO(
        DP_OP_425J2_127_3477_n680), .S(DP_OP_425J2_127_3477_n681) );
  FADDX1_HVT DP_OP_425J2_127_3477_U496 ( .A(DP_OP_425J2_127_3477_n898), .B(
        DP_OP_425J2_127_3477_n894), .CI(DP_OP_425J2_127_3477_n896), .CO(
        DP_OP_425J2_127_3477_n678), .S(DP_OP_425J2_127_3477_n679) );
  FADDX1_HVT DP_OP_425J2_127_3477_U495 ( .A(DP_OP_425J2_127_3477_n892), .B(
        DP_OP_425J2_127_3477_n878), .CI(DP_OP_425J2_127_3477_n880), .CO(
        DP_OP_425J2_127_3477_n676), .S(DP_OP_425J2_127_3477_n677) );
  FADDX1_HVT DP_OP_425J2_127_3477_U494 ( .A(DP_OP_425J2_127_3477_n890), .B(
        DP_OP_425J2_127_3477_n882), .CI(DP_OP_425J2_127_3477_n888), .CO(
        DP_OP_425J2_127_3477_n674), .S(DP_OP_425J2_127_3477_n675) );
  FADDX1_HVT DP_OP_425J2_127_3477_U493 ( .A(DP_OP_425J2_127_3477_n886), .B(
        DP_OP_425J2_127_3477_n884), .CI(DP_OP_425J2_127_3477_n719), .CO(
        DP_OP_425J2_127_3477_n672), .S(DP_OP_425J2_127_3477_n673) );
  FADDX1_HVT DP_OP_425J2_127_3477_U492 ( .A(DP_OP_425J2_127_3477_n876), .B(
        DP_OP_425J2_127_3477_n717), .CI(DP_OP_425J2_127_3477_n715), .CO(
        DP_OP_425J2_127_3477_n670), .S(DP_OP_425J2_127_3477_n671) );
  FADDX1_HVT DP_OP_425J2_127_3477_U491 ( .A(DP_OP_425J2_127_3477_n874), .B(
        DP_OP_425J2_127_3477_n711), .CI(DP_OP_425J2_127_3477_n713), .CO(
        DP_OP_425J2_127_3477_n668), .S(DP_OP_425J2_127_3477_n669) );
  FADDX1_HVT DP_OP_425J2_127_3477_U490 ( .A(DP_OP_425J2_127_3477_n872), .B(
        DP_OP_425J2_127_3477_n709), .CI(DP_OP_425J2_127_3477_n866), .CO(
        DP_OP_425J2_127_3477_n666), .S(DP_OP_425J2_127_3477_n667) );
  FADDX1_HVT DP_OP_425J2_127_3477_U489 ( .A(DP_OP_425J2_127_3477_n870), .B(
        DP_OP_425J2_127_3477_n868), .CI(DP_OP_425J2_127_3477_n856), .CO(
        DP_OP_425J2_127_3477_n664), .S(DP_OP_425J2_127_3477_n665) );
  FADDX1_HVT DP_OP_425J2_127_3477_U488 ( .A(DP_OP_425J2_127_3477_n864), .B(
        DP_OP_425J2_127_3477_n707), .CI(DP_OP_425J2_127_3477_n697), .CO(
        DP_OP_425J2_127_3477_n662), .S(DP_OP_425J2_127_3477_n663) );
  FADDX1_HVT DP_OP_425J2_127_3477_U487 ( .A(DP_OP_425J2_127_3477_n862), .B(
        DP_OP_425J2_127_3477_n703), .CI(DP_OP_425J2_127_3477_n699), .CO(
        DP_OP_425J2_127_3477_n660), .S(DP_OP_425J2_127_3477_n661) );
  FADDX1_HVT DP_OP_425J2_127_3477_U486 ( .A(DP_OP_425J2_127_3477_n860), .B(
        DP_OP_425J2_127_3477_n705), .CI(DP_OP_425J2_127_3477_n701), .CO(
        DP_OP_425J2_127_3477_n658), .S(DP_OP_425J2_127_3477_n659) );
  FADDX1_HVT DP_OP_425J2_127_3477_U485 ( .A(DP_OP_425J2_127_3477_n858), .B(
        DP_OP_425J2_127_3477_n693), .CI(DP_OP_425J2_127_3477_n689), .CO(
        DP_OP_425J2_127_3477_n656), .S(DP_OP_425J2_127_3477_n657) );
  FADDX1_HVT DP_OP_425J2_127_3477_U484 ( .A(DP_OP_425J2_127_3477_n691), .B(
        DP_OP_425J2_127_3477_n854), .CI(DP_OP_425J2_127_3477_n685), .CO(
        DP_OP_425J2_127_3477_n654), .S(DP_OP_425J2_127_3477_n655) );
  FADDX1_HVT DP_OP_425J2_127_3477_U483 ( .A(DP_OP_425J2_127_3477_n687), .B(
        DP_OP_425J2_127_3477_n695), .CI(DP_OP_425J2_127_3477_n681), .CO(
        DP_OP_425J2_127_3477_n652), .S(DP_OP_425J2_127_3477_n653) );
  FADDX1_HVT DP_OP_425J2_127_3477_U482 ( .A(DP_OP_425J2_127_3477_n683), .B(
        DP_OP_425J2_127_3477_n852), .CI(DP_OP_425J2_127_3477_n850), .CO(
        DP_OP_425J2_127_3477_n650), .S(DP_OP_425J2_127_3477_n651) );
  FADDX1_HVT DP_OP_425J2_127_3477_U481 ( .A(DP_OP_425J2_127_3477_n848), .B(
        DP_OP_425J2_127_3477_n846), .CI(DP_OP_425J2_127_3477_n679), .CO(
        DP_OP_425J2_127_3477_n648), .S(DP_OP_425J2_127_3477_n649) );
  FADDX1_HVT DP_OP_425J2_127_3477_U480 ( .A(DP_OP_425J2_127_3477_n844), .B(
        DP_OP_425J2_127_3477_n842), .CI(DP_OP_425J2_127_3477_n840), .CO(
        DP_OP_425J2_127_3477_n646), .S(DP_OP_425J2_127_3477_n647) );
  FADDX1_HVT DP_OP_425J2_127_3477_U479 ( .A(DP_OP_425J2_127_3477_n838), .B(
        DP_OP_425J2_127_3477_n673), .CI(DP_OP_425J2_127_3477_n832), .CO(
        DP_OP_425J2_127_3477_n644), .S(DP_OP_425J2_127_3477_n645) );
  FADDX1_HVT DP_OP_425J2_127_3477_U478 ( .A(DP_OP_425J2_127_3477_n836), .B(
        DP_OP_425J2_127_3477_n675), .CI(DP_OP_425J2_127_3477_n677), .CO(
        DP_OP_425J2_127_3477_n642), .S(DP_OP_425J2_127_3477_n643) );
  FADDX1_HVT DP_OP_425J2_127_3477_U477 ( .A(DP_OP_425J2_127_3477_n834), .B(
        DP_OP_425J2_127_3477_n671), .CI(DP_OP_425J2_127_3477_n667), .CO(
        DP_OP_425J2_127_3477_n640), .S(DP_OP_425J2_127_3477_n641) );
  FADDX1_HVT DP_OP_425J2_127_3477_U476 ( .A(DP_OP_425J2_127_3477_n830), .B(
        DP_OP_425J2_127_3477_n669), .CI(DP_OP_425J2_127_3477_n665), .CO(
        DP_OP_425J2_127_3477_n638), .S(DP_OP_425J2_127_3477_n639) );
  FADDX1_HVT DP_OP_425J2_127_3477_U475 ( .A(DP_OP_425J2_127_3477_n828), .B(
        DP_OP_425J2_127_3477_n826), .CI(DP_OP_425J2_127_3477_n661), .CO(
        DP_OP_425J2_127_3477_n636), .S(DP_OP_425J2_127_3477_n637) );
  FADDX1_HVT DP_OP_425J2_127_3477_U474 ( .A(DP_OP_425J2_127_3477_n659), .B(
        DP_OP_425J2_127_3477_n663), .CI(DP_OP_425J2_127_3477_n824), .CO(
        DP_OP_425J2_127_3477_n634), .S(DP_OP_425J2_127_3477_n635) );
  FADDX1_HVT DP_OP_425J2_127_3477_U473 ( .A(DP_OP_425J2_127_3477_n657), .B(
        DP_OP_425J2_127_3477_n822), .CI(DP_OP_425J2_127_3477_n653), .CO(
        DP_OP_425J2_127_3477_n632), .S(DP_OP_425J2_127_3477_n633) );
  FADDX1_HVT DP_OP_425J2_127_3477_U472 ( .A(DP_OP_425J2_127_3477_n655), .B(
        DP_OP_425J2_127_3477_n820), .CI(DP_OP_425J2_127_3477_n651), .CO(
        DP_OP_425J2_127_3477_n630), .S(DP_OP_425J2_127_3477_n631) );
  FADDX1_HVT DP_OP_425J2_127_3477_U471 ( .A(DP_OP_425J2_127_3477_n818), .B(
        DP_OP_425J2_127_3477_n816), .CI(DP_OP_425J2_127_3477_n649), .CO(
        DP_OP_425J2_127_3477_n628), .S(DP_OP_425J2_127_3477_n629) );
  FADDX1_HVT DP_OP_425J2_127_3477_U470 ( .A(DP_OP_425J2_127_3477_n814), .B(
        DP_OP_425J2_127_3477_n812), .CI(DP_OP_425J2_127_3477_n647), .CO(
        DP_OP_425J2_127_3477_n626), .S(DP_OP_425J2_127_3477_n627) );
  FADDX1_HVT DP_OP_425J2_127_3477_U469 ( .A(DP_OP_425J2_127_3477_n810), .B(
        DP_OP_425J2_127_3477_n643), .CI(DP_OP_425J2_127_3477_n806), .CO(
        DP_OP_425J2_127_3477_n624), .S(DP_OP_425J2_127_3477_n625) );
  FADDX1_HVT DP_OP_425J2_127_3477_U468 ( .A(DP_OP_425J2_127_3477_n808), .B(
        DP_OP_425J2_127_3477_n645), .CI(DP_OP_425J2_127_3477_n641), .CO(
        DP_OP_425J2_127_3477_n622), .S(DP_OP_425J2_127_3477_n623) );
  FADDX1_HVT DP_OP_425J2_127_3477_U467 ( .A(DP_OP_425J2_127_3477_n639), .B(
        DP_OP_425J2_127_3477_n804), .CI(DP_OP_425J2_127_3477_n637), .CO(
        DP_OP_425J2_127_3477_n620), .S(DP_OP_425J2_127_3477_n621) );
  FADDX1_HVT DP_OP_425J2_127_3477_U466 ( .A(DP_OP_425J2_127_3477_n635), .B(
        DP_OP_425J2_127_3477_n802), .CI(DP_OP_425J2_127_3477_n633), .CO(
        DP_OP_425J2_127_3477_n618), .S(DP_OP_425J2_127_3477_n619) );
  FADDX1_HVT DP_OP_425J2_127_3477_U465 ( .A(DP_OP_425J2_127_3477_n800), .B(
        DP_OP_425J2_127_3477_n631), .CI(DP_OP_425J2_127_3477_n798), .CO(
        DP_OP_425J2_127_3477_n616), .S(DP_OP_425J2_127_3477_n617) );
  FADDX1_HVT DP_OP_425J2_127_3477_U464 ( .A(DP_OP_425J2_127_3477_n796), .B(
        DP_OP_425J2_127_3477_n629), .CI(DP_OP_425J2_127_3477_n794), .CO(
        DP_OP_425J2_127_3477_n614), .S(DP_OP_425J2_127_3477_n615) );
  FADDX1_HVT DP_OP_425J2_127_3477_U463 ( .A(DP_OP_425J2_127_3477_n627), .B(
        DP_OP_425J2_127_3477_n792), .CI(DP_OP_425J2_127_3477_n625), .CO(
        DP_OP_425J2_127_3477_n612), .S(DP_OP_425J2_127_3477_n613) );
  FADDX1_HVT DP_OP_425J2_127_3477_U462 ( .A(DP_OP_425J2_127_3477_n623), .B(
        DP_OP_425J2_127_3477_n790), .CI(DP_OP_425J2_127_3477_n621), .CO(
        DP_OP_425J2_127_3477_n610), .S(DP_OP_425J2_127_3477_n611) );
  FADDX1_HVT DP_OP_425J2_127_3477_U461 ( .A(DP_OP_425J2_127_3477_n788), .B(
        DP_OP_425J2_127_3477_n619), .CI(DP_OP_425J2_127_3477_n786), .CO(
        DP_OP_425J2_127_3477_n608), .S(DP_OP_425J2_127_3477_n609) );
  FADDX1_HVT DP_OP_425J2_127_3477_U460 ( .A(DP_OP_425J2_127_3477_n617), .B(
        DP_OP_425J2_127_3477_n784), .CI(DP_OP_425J2_127_3477_n615), .CO(
        DP_OP_425J2_127_3477_n606), .S(DP_OP_425J2_127_3477_n607) );
  FADDX1_HVT DP_OP_425J2_127_3477_U459 ( .A(DP_OP_425J2_127_3477_n782), .B(
        DP_OP_425J2_127_3477_n613), .CI(DP_OP_425J2_127_3477_n611), .CO(
        DP_OP_425J2_127_3477_n604), .S(DP_OP_425J2_127_3477_n605) );
  FADDX1_HVT DP_OP_425J2_127_3477_U458 ( .A(DP_OP_425J2_127_3477_n780), .B(
        DP_OP_425J2_127_3477_n609), .CI(DP_OP_425J2_127_3477_n778), .CO(
        DP_OP_425J2_127_3477_n602), .S(DP_OP_425J2_127_3477_n603) );
  FADDX1_HVT DP_OP_425J2_127_3477_U457 ( .A(DP_OP_425J2_127_3477_n607), .B(
        DP_OP_425J2_127_3477_n776), .CI(DP_OP_425J2_127_3477_n605), .CO(
        DP_OP_425J2_127_3477_n600), .S(DP_OP_425J2_127_3477_n601) );
  FADDX1_HVT DP_OP_425J2_127_3477_U456 ( .A(DP_OP_425J2_127_3477_n774), .B(
        DP_OP_425J2_127_3477_n603), .CI(DP_OP_425J2_127_3477_n601), .CO(
        DP_OP_425J2_127_3477_n598), .S(DP_OP_425J2_127_3477_n599) );
  FADDX1_HVT DP_OP_425J2_127_3477_U455 ( .A(DP_OP_425J2_127_3477_n2977), .B(
        DP_OP_425J2_127_3477_n1921), .CI(DP_OP_425J2_127_3477_n1877), .CO(
        DP_OP_425J2_127_3477_n596), .S(DP_OP_425J2_127_3477_n597) );
  FADDX1_HVT DP_OP_425J2_127_3477_U454 ( .A(DP_OP_425J2_127_3477_n770), .B(
        DP_OP_425J2_127_3477_n2236), .CI(DP_OP_425J2_127_3477_n1928), .CO(
        DP_OP_425J2_127_3477_n594), .S(DP_OP_425J2_127_3477_n595) );
  FADDX1_HVT DP_OP_425J2_127_3477_U453 ( .A(DP_OP_425J2_127_3477_n2317), .B(
        DP_OP_425J2_127_3477_n2982), .CI(DP_OP_425J2_127_3477_n2632), .CO(
        DP_OP_425J2_127_3477_n592), .S(DP_OP_425J2_127_3477_n593) );
  FADDX1_HVT DP_OP_425J2_127_3477_U452 ( .A(DP_OP_425J2_127_3477_n2009), .B(
        DP_OP_425J2_127_3477_n2544), .CI(DP_OP_425J2_127_3477_n2764), .CO(
        DP_OP_425J2_127_3477_n590), .S(DP_OP_425J2_127_3477_n591) );
  FADDX1_HVT DP_OP_425J2_127_3477_U451 ( .A(DP_OP_425J2_127_3477_n2229), .B(
        DP_OP_425J2_127_3477_n2324), .CI(DP_OP_425J2_127_3477_n2940), .CO(
        DP_OP_425J2_127_3477_n588), .S(DP_OP_425J2_127_3477_n589) );
  FADDX1_HVT DP_OP_425J2_127_3477_U450 ( .A(DP_OP_425J2_127_3477_n1965), .B(
        DP_OP_425J2_127_3477_n2852), .CI(DP_OP_425J2_127_3477_n2016), .CO(
        DP_OP_425J2_127_3477_n586), .S(DP_OP_425J2_127_3477_n587) );
  FADDX1_HVT DP_OP_425J2_127_3477_U449 ( .A(DP_OP_425J2_127_3477_n2097), .B(
        DP_OP_425J2_127_3477_n1972), .CI(DP_OP_425J2_127_3477_n2808), .CO(
        DP_OP_425J2_127_3477_n584), .S(DP_OP_425J2_127_3477_n585) );
  FADDX1_HVT DP_OP_425J2_127_3477_U448 ( .A(DP_OP_425J2_127_3477_n2933), .B(
        DP_OP_425J2_127_3477_n2368), .CI(DP_OP_425J2_127_3477_n2456), .CO(
        DP_OP_425J2_127_3477_n582), .S(DP_OP_425J2_127_3477_n583) );
  FADDX1_HVT DP_OP_425J2_127_3477_U447 ( .A(DP_OP_425J2_127_3477_n2449), .B(
        DP_OP_425J2_127_3477_n2500), .CI(DP_OP_425J2_127_3477_n2896), .CO(
        DP_OP_425J2_127_3477_n580), .S(DP_OP_425J2_127_3477_n581) );
  FADDX1_HVT DP_OP_425J2_127_3477_U446 ( .A(DP_OP_425J2_127_3477_n2713), .B(
        DP_OP_425J2_127_3477_n2192), .CI(DP_OP_425J2_127_3477_n2720), .CO(
        DP_OP_425J2_127_3477_n578), .S(DP_OP_425J2_127_3477_n579) );
  FADDX1_HVT DP_OP_425J2_127_3477_U445 ( .A(DP_OP_425J2_127_3477_n2889), .B(
        DP_OP_425J2_127_3477_n2412), .CI(DP_OP_425J2_127_3477_n2588), .CO(
        DP_OP_425J2_127_3477_n576), .S(DP_OP_425J2_127_3477_n577) );
  FADDX1_HVT DP_OP_425J2_127_3477_U444 ( .A(DP_OP_425J2_127_3477_n2185), .B(
        DP_OP_425J2_127_3477_n2060), .CI(DP_OP_425J2_127_3477_n2676), .CO(
        DP_OP_425J2_127_3477_n574), .S(DP_OP_425J2_127_3477_n575) );
  FADDX1_HVT DP_OP_425J2_127_3477_U443 ( .A(DP_OP_425J2_127_3477_n2141), .B(
        DP_OP_425J2_127_3477_n2280), .CI(DP_OP_425J2_127_3477_n2148), .CO(
        DP_OP_425J2_127_3477_n572), .S(DP_OP_425J2_127_3477_n573) );
  FADDX1_HVT DP_OP_425J2_127_3477_U442 ( .A(DP_OP_425J2_127_3477_n2537), .B(
        DP_OP_425J2_127_3477_n2361), .CI(DP_OP_425J2_127_3477_n2104), .CO(
        DP_OP_425J2_127_3477_n570), .S(DP_OP_425J2_127_3477_n571) );
  FADDX1_HVT DP_OP_425J2_127_3477_U441 ( .A(DP_OP_425J2_127_3477_n2845), .B(
        DP_OP_425J2_127_3477_n2053), .CI(DP_OP_425J2_127_3477_n2273), .CO(
        DP_OP_425J2_127_3477_n568), .S(DP_OP_425J2_127_3477_n569) );
  FADDX1_HVT DP_OP_425J2_127_3477_U440 ( .A(DP_OP_425J2_127_3477_n2801), .B(
        DP_OP_425J2_127_3477_n2405), .CI(DP_OP_425J2_127_3477_n2493), .CO(
        DP_OP_425J2_127_3477_n566), .S(DP_OP_425J2_127_3477_n567) );
  FADDX1_HVT DP_OP_425J2_127_3477_U439 ( .A(DP_OP_425J2_127_3477_n2757), .B(
        DP_OP_425J2_127_3477_n2581), .CI(DP_OP_425J2_127_3477_n2625), .CO(
        DP_OP_425J2_127_3477_n564), .S(DP_OP_425J2_127_3477_n565) );
  FADDX1_HVT DP_OP_425J2_127_3477_U438 ( .A(DP_OP_425J2_127_3477_n2669), .B(
        DP_OP_425J2_127_3477_n768), .CI(DP_OP_425J2_127_3477_n766), .CO(
        DP_OP_425J2_127_3477_n562), .S(DP_OP_425J2_127_3477_n563) );
  FADDX1_HVT DP_OP_425J2_127_3477_U437 ( .A(DP_OP_425J2_127_3477_n764), .B(
        DP_OP_425J2_127_3477_n736), .CI(DP_OP_425J2_127_3477_n738), .CO(
        DP_OP_425J2_127_3477_n560), .S(DP_OP_425J2_127_3477_n561) );
  FADDX1_HVT DP_OP_425J2_127_3477_U436 ( .A(DP_OP_425J2_127_3477_n762), .B(
        DP_OP_425J2_127_3477_n740), .CI(DP_OP_425J2_127_3477_n742), .CO(
        DP_OP_425J2_127_3477_n558), .S(DP_OP_425J2_127_3477_n559) );
  FADDX1_HVT DP_OP_425J2_127_3477_U435 ( .A(DP_OP_425J2_127_3477_n760), .B(
        DP_OP_425J2_127_3477_n744), .CI(DP_OP_425J2_127_3477_n746), .CO(
        DP_OP_425J2_127_3477_n556), .S(DP_OP_425J2_127_3477_n557) );
  FADDX1_HVT DP_OP_425J2_127_3477_U434 ( .A(DP_OP_425J2_127_3477_n758), .B(
        DP_OP_425J2_127_3477_n748), .CI(DP_OP_425J2_127_3477_n750), .CO(
        DP_OP_425J2_127_3477_n554), .S(DP_OP_425J2_127_3477_n555) );
  FADDX1_HVT DP_OP_425J2_127_3477_U433 ( .A(DP_OP_425J2_127_3477_n756), .B(
        DP_OP_425J2_127_3477_n752), .CI(DP_OP_425J2_127_3477_n754), .CO(
        DP_OP_425J2_127_3477_n552), .S(DP_OP_425J2_127_3477_n553) );
  FADDX1_HVT DP_OP_425J2_127_3477_U432 ( .A(DP_OP_425J2_127_3477_n734), .B(
        DP_OP_425J2_127_3477_n720), .CI(DP_OP_425J2_127_3477_n732), .CO(
        DP_OP_425J2_127_3477_n550), .S(DP_OP_425J2_127_3477_n551) );
  FADDX1_HVT DP_OP_425J2_127_3477_U431 ( .A(DP_OP_425J2_127_3477_n726), .B(
        DP_OP_425J2_127_3477_n722), .CI(DP_OP_425J2_127_3477_n724), .CO(
        DP_OP_425J2_127_3477_n548), .S(DP_OP_425J2_127_3477_n549) );
  FADDX1_HVT DP_OP_425J2_127_3477_U430 ( .A(DP_OP_425J2_127_3477_n730), .B(
        DP_OP_425J2_127_3477_n728), .CI(DP_OP_425J2_127_3477_n595), .CO(
        DP_OP_425J2_127_3477_n546), .S(DP_OP_425J2_127_3477_n547) );
  FADDX1_HVT DP_OP_425J2_127_3477_U429 ( .A(DP_OP_425J2_127_3477_n597), .B(
        DP_OP_425J2_127_3477_n583), .CI(DP_OP_425J2_127_3477_n589), .CO(
        DP_OP_425J2_127_3477_n544), .S(DP_OP_425J2_127_3477_n545) );
  FADDX1_HVT DP_OP_425J2_127_3477_U428 ( .A(DP_OP_425J2_127_3477_n565), .B(
        DP_OP_425J2_127_3477_n587), .CI(DP_OP_425J2_127_3477_n585), .CO(
        DP_OP_425J2_127_3477_n542), .S(DP_OP_425J2_127_3477_n543) );
  FADDX1_HVT DP_OP_425J2_127_3477_U427 ( .A(DP_OP_425J2_127_3477_n591), .B(
        DP_OP_425J2_127_3477_n573), .CI(DP_OP_425J2_127_3477_n575), .CO(
        DP_OP_425J2_127_3477_n540), .S(DP_OP_425J2_127_3477_n541) );
  FADDX1_HVT DP_OP_425J2_127_3477_U426 ( .A(DP_OP_425J2_127_3477_n577), .B(
        DP_OP_425J2_127_3477_n567), .CI(DP_OP_425J2_127_3477_n569), .CO(
        DP_OP_425J2_127_3477_n538), .S(DP_OP_425J2_127_3477_n539) );
  FADDX1_HVT DP_OP_425J2_127_3477_U425 ( .A(DP_OP_425J2_127_3477_n571), .B(
        DP_OP_425J2_127_3477_n593), .CI(DP_OP_425J2_127_3477_n581), .CO(
        DP_OP_425J2_127_3477_n536), .S(DP_OP_425J2_127_3477_n537) );
  FADDX1_HVT DP_OP_425J2_127_3477_U424 ( .A(DP_OP_425J2_127_3477_n579), .B(
        DP_OP_425J2_127_3477_n718), .CI(DP_OP_425J2_127_3477_n716), .CO(
        DP_OP_425J2_127_3477_n534), .S(DP_OP_425J2_127_3477_n535) );
  FADDX1_HVT DP_OP_425J2_127_3477_U423 ( .A(DP_OP_425J2_127_3477_n714), .B(
        DP_OP_425J2_127_3477_n708), .CI(DP_OP_425J2_127_3477_n710), .CO(
        DP_OP_425J2_127_3477_n532), .S(DP_OP_425J2_127_3477_n533) );
  FADDX1_HVT DP_OP_425J2_127_3477_U422 ( .A(DP_OP_425J2_127_3477_n712), .B(
        DP_OP_425J2_127_3477_n706), .CI(DP_OP_425J2_127_3477_n704), .CO(
        DP_OP_425J2_127_3477_n530), .S(DP_OP_425J2_127_3477_n531) );
  FADDX1_HVT DP_OP_425J2_127_3477_U421 ( .A(DP_OP_425J2_127_3477_n702), .B(
        DP_OP_425J2_127_3477_n698), .CI(DP_OP_425J2_127_3477_n696), .CO(
        DP_OP_425J2_127_3477_n528), .S(DP_OP_425J2_127_3477_n529) );
  FADDX1_HVT DP_OP_425J2_127_3477_U420 ( .A(DP_OP_425J2_127_3477_n700), .B(
        DP_OP_425J2_127_3477_n563), .CI(DP_OP_425J2_127_3477_n557), .CO(
        DP_OP_425J2_127_3477_n526), .S(DP_OP_425J2_127_3477_n527) );
  FADDX1_HVT DP_OP_425J2_127_3477_U419 ( .A(DP_OP_425J2_127_3477_n559), .B(
        DP_OP_425J2_127_3477_n553), .CI(DP_OP_425J2_127_3477_n684), .CO(
        DP_OP_425J2_127_3477_n524), .S(DP_OP_425J2_127_3477_n525) );
  FADDX1_HVT DP_OP_425J2_127_3477_U418 ( .A(DP_OP_425J2_127_3477_n694), .B(
        DP_OP_425J2_127_3477_n561), .CI(DP_OP_425J2_127_3477_n555), .CO(
        DP_OP_425J2_127_3477_n522), .S(DP_OP_425J2_127_3477_n523) );
  FADDX1_HVT DP_OP_425J2_127_3477_U417 ( .A(DP_OP_425J2_127_3477_n688), .B(
        DP_OP_425J2_127_3477_n692), .CI(DP_OP_425J2_127_3477_n686), .CO(
        DP_OP_425J2_127_3477_n520), .S(DP_OP_425J2_127_3477_n521) );
  FADDX1_HVT DP_OP_425J2_127_3477_U416 ( .A(DP_OP_425J2_127_3477_n690), .B(
        DP_OP_425J2_127_3477_n682), .CI(DP_OP_425J2_127_3477_n680), .CO(
        DP_OP_425J2_127_3477_n518), .S(DP_OP_425J2_127_3477_n519) );
  FADDX1_HVT DP_OP_425J2_127_3477_U415 ( .A(DP_OP_425J2_127_3477_n549), .B(
        DP_OP_425J2_127_3477_n551), .CI(DP_OP_425J2_127_3477_n547), .CO(
        DP_OP_425J2_127_3477_n516), .S(DP_OP_425J2_127_3477_n517) );
  FADDX1_HVT DP_OP_425J2_127_3477_U414 ( .A(DP_OP_425J2_127_3477_n545), .B(
        DP_OP_425J2_127_3477_n539), .CI(DP_OP_425J2_127_3477_n543), .CO(
        DP_OP_425J2_127_3477_n514), .S(DP_OP_425J2_127_3477_n515) );
  FADDX1_HVT DP_OP_425J2_127_3477_U413 ( .A(DP_OP_425J2_127_3477_n537), .B(
        DP_OP_425J2_127_3477_n541), .CI(DP_OP_425J2_127_3477_n678), .CO(
        DP_OP_425J2_127_3477_n512), .S(DP_OP_425J2_127_3477_n513) );
  FADDX1_HVT DP_OP_425J2_127_3477_U412 ( .A(DP_OP_425J2_127_3477_n676), .B(
        DP_OP_425J2_127_3477_n672), .CI(DP_OP_425J2_127_3477_n535), .CO(
        DP_OP_425J2_127_3477_n510), .S(DP_OP_425J2_127_3477_n511) );
  FADDX1_HVT DP_OP_425J2_127_3477_U411 ( .A(DP_OP_425J2_127_3477_n674), .B(
        DP_OP_425J2_127_3477_n670), .CI(DP_OP_425J2_127_3477_n668), .CO(
        DP_OP_425J2_127_3477_n508), .S(DP_OP_425J2_127_3477_n509) );
  FADDX1_HVT DP_OP_425J2_127_3477_U410 ( .A(DP_OP_425J2_127_3477_n666), .B(
        DP_OP_425J2_127_3477_n533), .CI(DP_OP_425J2_127_3477_n531), .CO(
        DP_OP_425J2_127_3477_n506), .S(DP_OP_425J2_127_3477_n507) );
  FADDX1_HVT DP_OP_425J2_127_3477_U409 ( .A(DP_OP_425J2_127_3477_n664), .B(
        DP_OP_425J2_127_3477_n662), .CI(DP_OP_425J2_127_3477_n660), .CO(
        DP_OP_425J2_127_3477_n504), .S(DP_OP_425J2_127_3477_n505) );
  FADDX1_HVT DP_OP_425J2_127_3477_U408 ( .A(DP_OP_425J2_127_3477_n658), .B(
        DP_OP_425J2_127_3477_n529), .CI(DP_OP_425J2_127_3477_n656), .CO(
        DP_OP_425J2_127_3477_n502), .S(DP_OP_425J2_127_3477_n503) );
  FADDX1_HVT DP_OP_425J2_127_3477_U407 ( .A(DP_OP_425J2_127_3477_n527), .B(
        DP_OP_425J2_127_3477_n654), .CI(DP_OP_425J2_127_3477_n525), .CO(
        DP_OP_425J2_127_3477_n500), .S(DP_OP_425J2_127_3477_n501) );
  FADDX1_HVT DP_OP_425J2_127_3477_U406 ( .A(DP_OP_425J2_127_3477_n652), .B(
        DP_OP_425J2_127_3477_n521), .CI(DP_OP_425J2_127_3477_n519), .CO(
        DP_OP_425J2_127_3477_n498), .S(DP_OP_425J2_127_3477_n499) );
  FADDX1_HVT DP_OP_425J2_127_3477_U405 ( .A(DP_OP_425J2_127_3477_n523), .B(
        DP_OP_425J2_127_3477_n517), .CI(DP_OP_425J2_127_3477_n650), .CO(
        DP_OP_425J2_127_3477_n496), .S(DP_OP_425J2_127_3477_n497) );
  FADDX1_HVT DP_OP_425J2_127_3477_U404 ( .A(DP_OP_425J2_127_3477_n515), .B(
        DP_OP_425J2_127_3477_n648), .CI(DP_OP_425J2_127_3477_n513), .CO(
        DP_OP_425J2_127_3477_n494), .S(DP_OP_425J2_127_3477_n495) );
  FADDX1_HVT DP_OP_425J2_127_3477_U403 ( .A(DP_OP_425J2_127_3477_n646), .B(
        DP_OP_425J2_127_3477_n644), .CI(DP_OP_425J2_127_3477_n642), .CO(
        DP_OP_425J2_127_3477_n492), .S(DP_OP_425J2_127_3477_n493) );
  FADDX1_HVT DP_OP_425J2_127_3477_U402 ( .A(DP_OP_425J2_127_3477_n511), .B(
        DP_OP_425J2_127_3477_n640), .CI(DP_OP_425J2_127_3477_n509), .CO(
        DP_OP_425J2_127_3477_n490), .S(DP_OP_425J2_127_3477_n491) );
  FADDX1_HVT DP_OP_425J2_127_3477_U401 ( .A(DP_OP_425J2_127_3477_n638), .B(
        DP_OP_425J2_127_3477_n507), .CI(DP_OP_425J2_127_3477_n505), .CO(
        DP_OP_425J2_127_3477_n488), .S(DP_OP_425J2_127_3477_n489) );
  FADDX1_HVT DP_OP_425J2_127_3477_U400 ( .A(DP_OP_425J2_127_3477_n636), .B(
        DP_OP_425J2_127_3477_n634), .CI(DP_OP_425J2_127_3477_n503), .CO(
        DP_OP_425J2_127_3477_n486), .S(DP_OP_425J2_127_3477_n487) );
  FADDX1_HVT DP_OP_425J2_127_3477_U399 ( .A(DP_OP_425J2_127_3477_n632), .B(
        DP_OP_425J2_127_3477_n501), .CI(DP_OP_425J2_127_3477_n499), .CO(
        DP_OP_425J2_127_3477_n484), .S(DP_OP_425J2_127_3477_n485) );
  FADDX1_HVT DP_OP_425J2_127_3477_U398 ( .A(DP_OP_425J2_127_3477_n630), .B(
        DP_OP_425J2_127_3477_n497), .CI(DP_OP_425J2_127_3477_n628), .CO(
        DP_OP_425J2_127_3477_n482), .S(DP_OP_425J2_127_3477_n483) );
  FADDX1_HVT DP_OP_425J2_127_3477_U397 ( .A(DP_OP_425J2_127_3477_n495), .B(
        DP_OP_425J2_127_3477_n626), .CI(DP_OP_425J2_127_3477_n493), .CO(
        DP_OP_425J2_127_3477_n480), .S(DP_OP_425J2_127_3477_n481) );
  FADDX1_HVT DP_OP_425J2_127_3477_U396 ( .A(DP_OP_425J2_127_3477_n624), .B(
        DP_OP_425J2_127_3477_n622), .CI(DP_OP_425J2_127_3477_n491), .CO(
        DP_OP_425J2_127_3477_n478), .S(DP_OP_425J2_127_3477_n479) );
  FADDX1_HVT DP_OP_425J2_127_3477_U395 ( .A(DP_OP_425J2_127_3477_n620), .B(
        DP_OP_425J2_127_3477_n489), .CI(DP_OP_425J2_127_3477_n487), .CO(
        DP_OP_425J2_127_3477_n476), .S(DP_OP_425J2_127_3477_n477) );
  FADDX1_HVT DP_OP_425J2_127_3477_U394 ( .A(DP_OP_425J2_127_3477_n618), .B(
        DP_OP_425J2_127_3477_n485), .CI(DP_OP_425J2_127_3477_n616), .CO(
        DP_OP_425J2_127_3477_n474), .S(DP_OP_425J2_127_3477_n475) );
  FADDX1_HVT DP_OP_425J2_127_3477_U393 ( .A(DP_OP_425J2_127_3477_n483), .B(
        DP_OP_425J2_127_3477_n614), .CI(DP_OP_425J2_127_3477_n481), .CO(
        DP_OP_425J2_127_3477_n472), .S(DP_OP_425J2_127_3477_n473) );
  FADDX1_HVT DP_OP_425J2_127_3477_U392 ( .A(DP_OP_425J2_127_3477_n612), .B(
        DP_OP_425J2_127_3477_n479), .CI(DP_OP_425J2_127_3477_n610), .CO(
        DP_OP_425J2_127_3477_n470), .S(DP_OP_425J2_127_3477_n471) );
  FADDX1_HVT DP_OP_425J2_127_3477_U391 ( .A(DP_OP_425J2_127_3477_n477), .B(
        DP_OP_425J2_127_3477_n608), .CI(DP_OP_425J2_127_3477_n475), .CO(
        DP_OP_425J2_127_3477_n468), .S(DP_OP_425J2_127_3477_n469) );
  FADDX1_HVT DP_OP_425J2_127_3477_U390 ( .A(DP_OP_425J2_127_3477_n606), .B(
        DP_OP_425J2_127_3477_n473), .CI(DP_OP_425J2_127_3477_n604), .CO(
        DP_OP_425J2_127_3477_n466), .S(DP_OP_425J2_127_3477_n467) );
  FADDX1_HVT DP_OP_425J2_127_3477_U389 ( .A(DP_OP_425J2_127_3477_n471), .B(
        DP_OP_425J2_127_3477_n469), .CI(DP_OP_425J2_127_3477_n602), .CO(
        DP_OP_425J2_127_3477_n464), .S(DP_OP_425J2_127_3477_n465) );
  FADDX1_HVT DP_OP_425J2_127_3477_U388 ( .A(DP_OP_425J2_127_3477_n600), .B(
        DP_OP_425J2_127_3477_n467), .CI(DP_OP_425J2_127_3477_n465), .CO(
        DP_OP_425J2_127_3477_n462), .S(DP_OP_425J2_127_3477_n463) );
  FADDX1_HVT DP_OP_425J2_127_3477_U386 ( .A(DP_OP_425J2_127_3477_n2976), .B(
        DP_OP_425J2_127_3477_n1920), .CI(DP_OP_425J2_127_3477_n461), .CO(
        DP_OP_425J2_127_3477_n458), .S(DP_OP_425J2_127_3477_n459) );
  FADDX1_HVT DP_OP_425J2_127_3477_U385 ( .A(DP_OP_425J2_127_3477_n2008), .B(
        DP_OP_425J2_127_3477_n2932), .CI(DP_OP_425J2_127_3477_n2360), .CO(
        DP_OP_425J2_127_3477_n456), .S(DP_OP_425J2_127_3477_n457) );
  FADDX1_HVT DP_OP_425J2_127_3477_U384 ( .A(DP_OP_425J2_127_3477_n2492), .B(
        DP_OP_425J2_127_3477_n2888), .CI(DP_OP_425J2_127_3477_n2844), .CO(
        DP_OP_425J2_127_3477_n454), .S(DP_OP_425J2_127_3477_n455) );
  FADDX1_HVT DP_OP_425J2_127_3477_U383 ( .A(DP_OP_425J2_127_3477_n2316), .B(
        DP_OP_425J2_127_3477_n2800), .CI(DP_OP_425J2_127_3477_n2756), .CO(
        DP_OP_425J2_127_3477_n452), .S(DP_OP_425J2_127_3477_n453) );
  FADDX1_HVT DP_OP_425J2_127_3477_U382 ( .A(DP_OP_425J2_127_3477_n2184), .B(
        DP_OP_425J2_127_3477_n1964), .CI(DP_OP_425J2_127_3477_n2712), .CO(
        DP_OP_425J2_127_3477_n450), .S(DP_OP_425J2_127_3477_n451) );
  FADDX1_HVT DP_OP_425J2_127_3477_U381 ( .A(DP_OP_425J2_127_3477_n2668), .B(
        DP_OP_425J2_127_3477_n2624), .CI(DP_OP_425J2_127_3477_n2580), .CO(
        DP_OP_425J2_127_3477_n448), .S(DP_OP_425J2_127_3477_n449) );
  FADDX1_HVT DP_OP_425J2_127_3477_U380 ( .A(DP_OP_425J2_127_3477_n2228), .B(
        DP_OP_425J2_127_3477_n2052), .CI(DP_OP_425J2_127_3477_n2096), .CO(
        DP_OP_425J2_127_3477_n446), .S(DP_OP_425J2_127_3477_n447) );
  FADDX1_HVT DP_OP_425J2_127_3477_U379 ( .A(DP_OP_425J2_127_3477_n2140), .B(
        DP_OP_425J2_127_3477_n2536), .CI(DP_OP_425J2_127_3477_n2448), .CO(
        DP_OP_425J2_127_3477_n444), .S(DP_OP_425J2_127_3477_n445) );
  FADDX1_HVT DP_OP_425J2_127_3477_U378 ( .A(DP_OP_425J2_127_3477_n2272), .B(
        DP_OP_425J2_127_3477_n2404), .CI(DP_OP_425J2_127_3477_n596), .CO(
        DP_OP_425J2_127_3477_n442), .S(DP_OP_425J2_127_3477_n443) );
  FADDX1_HVT DP_OP_425J2_127_3477_U377 ( .A(DP_OP_425J2_127_3477_n594), .B(
        DP_OP_425J2_127_3477_n564), .CI(DP_OP_425J2_127_3477_n592), .CO(
        DP_OP_425J2_127_3477_n440), .S(DP_OP_425J2_127_3477_n441) );
  FADDX1_HVT DP_OP_425J2_127_3477_U376 ( .A(DP_OP_425J2_127_3477_n590), .B(
        DP_OP_425J2_127_3477_n566), .CI(DP_OP_425J2_127_3477_n568), .CO(
        DP_OP_425J2_127_3477_n438), .S(DP_OP_425J2_127_3477_n439) );
  FADDX1_HVT DP_OP_425J2_127_3477_U375 ( .A(DP_OP_425J2_127_3477_n588), .B(
        DP_OP_425J2_127_3477_n570), .CI(DP_OP_425J2_127_3477_n572), .CO(
        DP_OP_425J2_127_3477_n436), .S(DP_OP_425J2_127_3477_n437) );
  FADDX1_HVT DP_OP_425J2_127_3477_U374 ( .A(DP_OP_425J2_127_3477_n586), .B(
        DP_OP_425J2_127_3477_n574), .CI(DP_OP_425J2_127_3477_n576), .CO(
        DP_OP_425J2_127_3477_n434), .S(DP_OP_425J2_127_3477_n435) );
  FADDX1_HVT DP_OP_425J2_127_3477_U373 ( .A(DP_OP_425J2_127_3477_n584), .B(
        DP_OP_425J2_127_3477_n578), .CI(DP_OP_425J2_127_3477_n580), .CO(
        DP_OP_425J2_127_3477_n432), .S(DP_OP_425J2_127_3477_n433) );
  FADDX1_HVT DP_OP_425J2_127_3477_U372 ( .A(DP_OP_425J2_127_3477_n582), .B(
        DP_OP_425J2_127_3477_n459), .CI(DP_OP_425J2_127_3477_n455), .CO(
        DP_OP_425J2_127_3477_n430), .S(DP_OP_425J2_127_3477_n431) );
  FADDX1_HVT DP_OP_425J2_127_3477_U371 ( .A(DP_OP_425J2_127_3477_n451), .B(
        DP_OP_425J2_127_3477_n445), .CI(DP_OP_425J2_127_3477_n447), .CO(
        DP_OP_425J2_127_3477_n428), .S(DP_OP_425J2_127_3477_n429) );
  FADDX1_HVT DP_OP_425J2_127_3477_U370 ( .A(DP_OP_425J2_127_3477_n449), .B(
        DP_OP_425J2_127_3477_n457), .CI(DP_OP_425J2_127_3477_n453), .CO(
        DP_OP_425J2_127_3477_n426), .S(DP_OP_425J2_127_3477_n427) );
  FADDX1_HVT DP_OP_425J2_127_3477_U369 ( .A(DP_OP_425J2_127_3477_n562), .B(
        DP_OP_425J2_127_3477_n560), .CI(DP_OP_425J2_127_3477_n552), .CO(
        DP_OP_425J2_127_3477_n424), .S(DP_OP_425J2_127_3477_n425) );
  FADDX1_HVT DP_OP_425J2_127_3477_U368 ( .A(DP_OP_425J2_127_3477_n558), .B(
        DP_OP_425J2_127_3477_n554), .CI(DP_OP_425J2_127_3477_n556), .CO(
        DP_OP_425J2_127_3477_n422), .S(DP_OP_425J2_127_3477_n423) );
  FADDX1_HVT DP_OP_425J2_127_3477_U367 ( .A(DP_OP_425J2_127_3477_n550), .B(
        DP_OP_425J2_127_3477_n546), .CI(DP_OP_425J2_127_3477_n443), .CO(
        DP_OP_425J2_127_3477_n420), .S(DP_OP_425J2_127_3477_n421) );
  FADDX1_HVT DP_OP_425J2_127_3477_U366 ( .A(DP_OP_425J2_127_3477_n548), .B(
        DP_OP_425J2_127_3477_n544), .CI(DP_OP_425J2_127_3477_n441), .CO(
        DP_OP_425J2_127_3477_n418), .S(DP_OP_425J2_127_3477_n419) );
  FADDX1_HVT DP_OP_425J2_127_3477_U365 ( .A(DP_OP_425J2_127_3477_n542), .B(
        DP_OP_425J2_127_3477_n435), .CI(DP_OP_425J2_127_3477_n437), .CO(
        DP_OP_425J2_127_3477_n416), .S(DP_OP_425J2_127_3477_n417) );
  FADDX1_HVT DP_OP_425J2_127_3477_U364 ( .A(DP_OP_425J2_127_3477_n540), .B(
        DP_OP_425J2_127_3477_n439), .CI(DP_OP_425J2_127_3477_n433), .CO(
        DP_OP_425J2_127_3477_n414), .S(DP_OP_425J2_127_3477_n415) );
  FADDX1_HVT DP_OP_425J2_127_3477_U363 ( .A(DP_OP_425J2_127_3477_n538), .B(
        DP_OP_425J2_127_3477_n536), .CI(DP_OP_425J2_127_3477_n534), .CO(
        DP_OP_425J2_127_3477_n412), .S(DP_OP_425J2_127_3477_n413) );
  FADDX1_HVT DP_OP_425J2_127_3477_U362 ( .A(DP_OP_425J2_127_3477_n431), .B(
        DP_OP_425J2_127_3477_n427), .CI(DP_OP_425J2_127_3477_n532), .CO(
        DP_OP_425J2_127_3477_n410), .S(DP_OP_425J2_127_3477_n411) );
  FADDX1_HVT DP_OP_425J2_127_3477_U361 ( .A(DP_OP_425J2_127_3477_n429), .B(
        DP_OP_425J2_127_3477_n530), .CI(DP_OP_425J2_127_3477_n528), .CO(
        DP_OP_425J2_127_3477_n408), .S(DP_OP_425J2_127_3477_n409) );
  FADDX1_HVT DP_OP_425J2_127_3477_U360 ( .A(DP_OP_425J2_127_3477_n526), .B(
        DP_OP_425J2_127_3477_n425), .CI(DP_OP_425J2_127_3477_n423), .CO(
        DP_OP_425J2_127_3477_n406), .S(DP_OP_425J2_127_3477_n407) );
  FADDX1_HVT DP_OP_425J2_127_3477_U359 ( .A(DP_OP_425J2_127_3477_n524), .B(
        DP_OP_425J2_127_3477_n520), .CI(DP_OP_425J2_127_3477_n518), .CO(
        DP_OP_425J2_127_3477_n404), .S(DP_OP_425J2_127_3477_n405) );
  FADDX1_HVT DP_OP_425J2_127_3477_U358 ( .A(DP_OP_425J2_127_3477_n522), .B(
        DP_OP_425J2_127_3477_n516), .CI(DP_OP_425J2_127_3477_n421), .CO(
        DP_OP_425J2_127_3477_n402), .S(DP_OP_425J2_127_3477_n403) );
  FADDX1_HVT DP_OP_425J2_127_3477_U357 ( .A(DP_OP_425J2_127_3477_n419), .B(
        DP_OP_425J2_127_3477_n514), .CI(DP_OP_425J2_127_3477_n512), .CO(
        DP_OP_425J2_127_3477_n400), .S(DP_OP_425J2_127_3477_n401) );
  FADDX1_HVT DP_OP_425J2_127_3477_U356 ( .A(DP_OP_425J2_127_3477_n417), .B(
        DP_OP_425J2_127_3477_n415), .CI(DP_OP_425J2_127_3477_n413), .CO(
        DP_OP_425J2_127_3477_n398), .S(DP_OP_425J2_127_3477_n399) );
  FADDX1_HVT DP_OP_425J2_127_3477_U355 ( .A(DP_OP_425J2_127_3477_n510), .B(
        DP_OP_425J2_127_3477_n508), .CI(DP_OP_425J2_127_3477_n411), .CO(
        DP_OP_425J2_127_3477_n396), .S(DP_OP_425J2_127_3477_n397) );
  FADDX1_HVT DP_OP_425J2_127_3477_U354 ( .A(DP_OP_425J2_127_3477_n506), .B(
        DP_OP_425J2_127_3477_n409), .CI(DP_OP_425J2_127_3477_n504), .CO(
        DP_OP_425J2_127_3477_n394), .S(DP_OP_425J2_127_3477_n395) );
  FADDX1_HVT DP_OP_425J2_127_3477_U353 ( .A(DP_OP_425J2_127_3477_n502), .B(
        DP_OP_425J2_127_3477_n407), .CI(DP_OP_425J2_127_3477_n500), .CO(
        DP_OP_425J2_127_3477_n392), .S(DP_OP_425J2_127_3477_n393) );
  FADDX1_HVT DP_OP_425J2_127_3477_U352 ( .A(DP_OP_425J2_127_3477_n498), .B(
        DP_OP_425J2_127_3477_n405), .CI(DP_OP_425J2_127_3477_n403), .CO(
        DP_OP_425J2_127_3477_n390), .S(DP_OP_425J2_127_3477_n391) );
  FADDX1_HVT DP_OP_425J2_127_3477_U351 ( .A(DP_OP_425J2_127_3477_n496), .B(
        DP_OP_425J2_127_3477_n401), .CI(DP_OP_425J2_127_3477_n494), .CO(
        DP_OP_425J2_127_3477_n388), .S(DP_OP_425J2_127_3477_n389) );
  FADDX1_HVT DP_OP_425J2_127_3477_U350 ( .A(DP_OP_425J2_127_3477_n399), .B(
        DP_OP_425J2_127_3477_n492), .CI(DP_OP_425J2_127_3477_n490), .CO(
        DP_OP_425J2_127_3477_n386), .S(DP_OP_425J2_127_3477_n387) );
  FADDX1_HVT DP_OP_425J2_127_3477_U349 ( .A(DP_OP_425J2_127_3477_n397), .B(
        DP_OP_425J2_127_3477_n488), .CI(DP_OP_425J2_127_3477_n395), .CO(
        DP_OP_425J2_127_3477_n384), .S(DP_OP_425J2_127_3477_n385) );
  FADDX1_HVT DP_OP_425J2_127_3477_U348 ( .A(DP_OP_425J2_127_3477_n486), .B(
        DP_OP_425J2_127_3477_n393), .CI(DP_OP_425J2_127_3477_n484), .CO(
        DP_OP_425J2_127_3477_n382), .S(DP_OP_425J2_127_3477_n383) );
  FADDX1_HVT DP_OP_425J2_127_3477_U347 ( .A(DP_OP_425J2_127_3477_n391), .B(
        DP_OP_425J2_127_3477_n482), .CI(DP_OP_425J2_127_3477_n389), .CO(
        DP_OP_425J2_127_3477_n380), .S(DP_OP_425J2_127_3477_n381) );
  FADDX1_HVT DP_OP_425J2_127_3477_U346 ( .A(DP_OP_425J2_127_3477_n480), .B(
        DP_OP_425J2_127_3477_n387), .CI(DP_OP_425J2_127_3477_n478), .CO(
        DP_OP_425J2_127_3477_n378), .S(DP_OP_425J2_127_3477_n379) );
  FADDX1_HVT DP_OP_425J2_127_3477_U345 ( .A(DP_OP_425J2_127_3477_n385), .B(
        DP_OP_425J2_127_3477_n476), .CI(DP_OP_425J2_127_3477_n383), .CO(
        DP_OP_425J2_127_3477_n376), .S(DP_OP_425J2_127_3477_n377) );
  FADDX1_HVT DP_OP_425J2_127_3477_U344 ( .A(DP_OP_425J2_127_3477_n474), .B(
        DP_OP_425J2_127_3477_n381), .CI(DP_OP_425J2_127_3477_n472), .CO(
        DP_OP_425J2_127_3477_n374), .S(DP_OP_425J2_127_3477_n375) );
  FADDX1_HVT DP_OP_425J2_127_3477_U343 ( .A(DP_OP_425J2_127_3477_n379), .B(
        DP_OP_425J2_127_3477_n470), .CI(DP_OP_425J2_127_3477_n377), .CO(
        DP_OP_425J2_127_3477_n372), .S(DP_OP_425J2_127_3477_n373) );
  FADDX1_HVT DP_OP_425J2_127_3477_U342 ( .A(DP_OP_425J2_127_3477_n468), .B(
        DP_OP_425J2_127_3477_n375), .CI(DP_OP_425J2_127_3477_n466), .CO(
        DP_OP_425J2_127_3477_n370), .S(DP_OP_425J2_127_3477_n371) );
  FADDX1_HVT DP_OP_425J2_127_3477_U341 ( .A(DP_OP_425J2_127_3477_n373), .B(
        DP_OP_425J2_127_3477_n464), .CI(DP_OP_425J2_127_3477_n371), .CO(
        DP_OP_425J2_127_3477_n368), .S(DP_OP_425J2_127_3477_n369) );
  FADDX1_HVT DP_OP_425J2_127_3477_U340 ( .A(DP_OP_425J2_127_3477_n1876), .B(
        DP_OP_425J2_127_3477_n460), .CI(DP_OP_425J2_127_3477_n458), .CO(
        DP_OP_425J2_127_3477_n366), .S(DP_OP_425J2_127_3477_n367) );
  FADDX1_HVT DP_OP_425J2_127_3477_U339 ( .A(DP_OP_425J2_127_3477_n448), .B(
        DP_OP_425J2_127_3477_n444), .CI(DP_OP_425J2_127_3477_n456), .CO(
        DP_OP_425J2_127_3477_n364), .S(DP_OP_425J2_127_3477_n365) );
  FADDX1_HVT DP_OP_425J2_127_3477_U338 ( .A(DP_OP_425J2_127_3477_n454), .B(
        DP_OP_425J2_127_3477_n452), .CI(DP_OP_425J2_127_3477_n450), .CO(
        DP_OP_425J2_127_3477_n362), .S(DP_OP_425J2_127_3477_n363) );
  FADDX1_HVT DP_OP_425J2_127_3477_U337 ( .A(DP_OP_425J2_127_3477_n446), .B(
        DP_OP_425J2_127_3477_n442), .CI(DP_OP_425J2_127_3477_n440), .CO(
        DP_OP_425J2_127_3477_n360), .S(DP_OP_425J2_127_3477_n361) );
  FADDX1_HVT DP_OP_425J2_127_3477_U336 ( .A(DP_OP_425J2_127_3477_n438), .B(
        DP_OP_425J2_127_3477_n436), .CI(DP_OP_425J2_127_3477_n434), .CO(
        DP_OP_425J2_127_3477_n358), .S(DP_OP_425J2_127_3477_n359) );
  FADDX1_HVT DP_OP_425J2_127_3477_U335 ( .A(DP_OP_425J2_127_3477_n432), .B(
        DP_OP_425J2_127_3477_n367), .CI(DP_OP_425J2_127_3477_n430), .CO(
        DP_OP_425J2_127_3477_n356), .S(DP_OP_425J2_127_3477_n357) );
  FADDX1_HVT DP_OP_425J2_127_3477_U334 ( .A(DP_OP_425J2_127_3477_n428), .B(
        DP_OP_425J2_127_3477_n363), .CI(DP_OP_425J2_127_3477_n365), .CO(
        DP_OP_425J2_127_3477_n354), .S(DP_OP_425J2_127_3477_n355) );
  FADDX1_HVT DP_OP_425J2_127_3477_U333 ( .A(DP_OP_425J2_127_3477_n426), .B(
        DP_OP_425J2_127_3477_n424), .CI(DP_OP_425J2_127_3477_n422), .CO(
        DP_OP_425J2_127_3477_n352), .S(DP_OP_425J2_127_3477_n353) );
  FADDX1_HVT DP_OP_425J2_127_3477_U332 ( .A(DP_OP_425J2_127_3477_n420), .B(
        DP_OP_425J2_127_3477_n361), .CI(DP_OP_425J2_127_3477_n418), .CO(
        DP_OP_425J2_127_3477_n350), .S(DP_OP_425J2_127_3477_n351) );
  FADDX1_HVT DP_OP_425J2_127_3477_U331 ( .A(DP_OP_425J2_127_3477_n416), .B(
        DP_OP_425J2_127_3477_n359), .CI(DP_OP_425J2_127_3477_n414), .CO(
        DP_OP_425J2_127_3477_n348), .S(DP_OP_425J2_127_3477_n349) );
  FADDX1_HVT DP_OP_425J2_127_3477_U330 ( .A(DP_OP_425J2_127_3477_n412), .B(
        DP_OP_425J2_127_3477_n357), .CI(DP_OP_425J2_127_3477_n410), .CO(
        DP_OP_425J2_127_3477_n346), .S(DP_OP_425J2_127_3477_n347) );
  FADDX1_HVT DP_OP_425J2_127_3477_U329 ( .A(DP_OP_425J2_127_3477_n355), .B(
        DP_OP_425J2_127_3477_n408), .CI(DP_OP_425J2_127_3477_n406), .CO(
        DP_OP_425J2_127_3477_n344), .S(DP_OP_425J2_127_3477_n345) );
  FADDX1_HVT DP_OP_425J2_127_3477_U328 ( .A(DP_OP_425J2_127_3477_n353), .B(
        DP_OP_425J2_127_3477_n404), .CI(DP_OP_425J2_127_3477_n402), .CO(
        DP_OP_425J2_127_3477_n342), .S(DP_OP_425J2_127_3477_n343) );
  FADDX1_HVT DP_OP_425J2_127_3477_U327 ( .A(DP_OP_425J2_127_3477_n351), .B(
        DP_OP_425J2_127_3477_n400), .CI(DP_OP_425J2_127_3477_n349), .CO(
        DP_OP_425J2_127_3477_n340), .S(DP_OP_425J2_127_3477_n341) );
  FADDX1_HVT DP_OP_425J2_127_3477_U326 ( .A(DP_OP_425J2_127_3477_n398), .B(
        DP_OP_425J2_127_3477_n347), .CI(DP_OP_425J2_127_3477_n396), .CO(
        DP_OP_425J2_127_3477_n338), .S(DP_OP_425J2_127_3477_n339) );
  FADDX1_HVT DP_OP_425J2_127_3477_U325 ( .A(DP_OP_425J2_127_3477_n394), .B(
        DP_OP_425J2_127_3477_n345), .CI(DP_OP_425J2_127_3477_n392), .CO(
        DP_OP_425J2_127_3477_n336), .S(DP_OP_425J2_127_3477_n337) );
  FADDX1_HVT DP_OP_425J2_127_3477_U324 ( .A(DP_OP_425J2_127_3477_n343), .B(
        DP_OP_425J2_127_3477_n390), .CI(DP_OP_425J2_127_3477_n388), .CO(
        DP_OP_425J2_127_3477_n334), .S(DP_OP_425J2_127_3477_n335) );
  FADDX1_HVT DP_OP_425J2_127_3477_U323 ( .A(DP_OP_425J2_127_3477_n341), .B(
        DP_OP_425J2_127_3477_n386), .CI(DP_OP_425J2_127_3477_n339), .CO(
        DP_OP_425J2_127_3477_n332), .S(DP_OP_425J2_127_3477_n333) );
  FADDX1_HVT DP_OP_425J2_127_3477_U322 ( .A(DP_OP_425J2_127_3477_n384), .B(
        DP_OP_425J2_127_3477_n337), .CI(DP_OP_425J2_127_3477_n382), .CO(
        DP_OP_425J2_127_3477_n330), .S(DP_OP_425J2_127_3477_n331) );
  FADDX1_HVT DP_OP_425J2_127_3477_U321 ( .A(DP_OP_425J2_127_3477_n380), .B(
        DP_OP_425J2_127_3477_n335), .CI(DP_OP_425J2_127_3477_n333), .CO(
        DP_OP_425J2_127_3477_n328), .S(DP_OP_425J2_127_3477_n329) );
  FADDX1_HVT DP_OP_425J2_127_3477_U320 ( .A(DP_OP_425J2_127_3477_n378), .B(
        DP_OP_425J2_127_3477_n331), .CI(DP_OP_425J2_127_3477_n376), .CO(
        DP_OP_425J2_127_3477_n326), .S(DP_OP_425J2_127_3477_n327) );
  FADDX1_HVT DP_OP_425J2_127_3477_U319 ( .A(DP_OP_425J2_127_3477_n374), .B(
        DP_OP_425J2_127_3477_n329), .CI(DP_OP_425J2_127_3477_n372), .CO(
        DP_OP_425J2_127_3477_n324), .S(DP_OP_425J2_127_3477_n325) );
  FADDX1_HVT DP_OP_425J2_127_3477_U318 ( .A(DP_OP_425J2_127_3477_n327), .B(
        DP_OP_425J2_127_3477_n370), .CI(DP_OP_425J2_127_3477_n325), .CO(
        DP_OP_425J2_127_3477_n322), .S(DP_OP_425J2_127_3477_n323) );
  FADDX1_HVT DP_OP_425J2_127_3477_U317 ( .A(DP_OP_425J2_127_3477_n1875), .B(
        DP_OP_425J2_127_3477_n366), .CI(DP_OP_425J2_127_3477_n364), .CO(
        DP_OP_425J2_127_3477_n320), .S(DP_OP_425J2_127_3477_n321) );
  FADDX1_HVT DP_OP_425J2_127_3477_U316 ( .A(DP_OP_425J2_127_3477_n362), .B(
        DP_OP_425J2_127_3477_n360), .CI(DP_OP_425J2_127_3477_n358), .CO(
        DP_OP_425J2_127_3477_n318), .S(DP_OP_425J2_127_3477_n319) );
  FADDX1_HVT DP_OP_425J2_127_3477_U315 ( .A(DP_OP_425J2_127_3477_n356), .B(
        DP_OP_425J2_127_3477_n321), .CI(DP_OP_425J2_127_3477_n354), .CO(
        DP_OP_425J2_127_3477_n316), .S(DP_OP_425J2_127_3477_n317) );
  FADDX1_HVT DP_OP_425J2_127_3477_U314 ( .A(DP_OP_425J2_127_3477_n352), .B(
        DP_OP_425J2_127_3477_n350), .CI(DP_OP_425J2_127_3477_n319), .CO(
        DP_OP_425J2_127_3477_n314), .S(DP_OP_425J2_127_3477_n315) );
  FADDX1_HVT DP_OP_425J2_127_3477_U313 ( .A(DP_OP_425J2_127_3477_n348), .B(
        DP_OP_425J2_127_3477_n346), .CI(DP_OP_425J2_127_3477_n317), .CO(
        DP_OP_425J2_127_3477_n312), .S(DP_OP_425J2_127_3477_n313) );
  FADDX1_HVT DP_OP_425J2_127_3477_U312 ( .A(DP_OP_425J2_127_3477_n344), .B(
        DP_OP_425J2_127_3477_n342), .CI(DP_OP_425J2_127_3477_n315), .CO(
        DP_OP_425J2_127_3477_n310), .S(DP_OP_425J2_127_3477_n311) );
  FADDX1_HVT DP_OP_425J2_127_3477_U311 ( .A(DP_OP_425J2_127_3477_n340), .B(
        DP_OP_425J2_127_3477_n313), .CI(DP_OP_425J2_127_3477_n338), .CO(
        DP_OP_425J2_127_3477_n308), .S(DP_OP_425J2_127_3477_n309) );
  FADDX1_HVT DP_OP_425J2_127_3477_U310 ( .A(DP_OP_425J2_127_3477_n336), .B(
        DP_OP_425J2_127_3477_n311), .CI(DP_OP_425J2_127_3477_n334), .CO(
        DP_OP_425J2_127_3477_n306), .S(DP_OP_425J2_127_3477_n307) );
  FADDX1_HVT DP_OP_425J2_127_3477_U309 ( .A(DP_OP_425J2_127_3477_n332), .B(
        DP_OP_425J2_127_3477_n309), .CI(DP_OP_425J2_127_3477_n330), .CO(
        DP_OP_425J2_127_3477_n304), .S(DP_OP_425J2_127_3477_n305) );
  FADDX1_HVT DP_OP_425J2_127_3477_U308 ( .A(DP_OP_425J2_127_3477_n307), .B(
        DP_OP_425J2_127_3477_n328), .CI(DP_OP_425J2_127_3477_n305), .CO(
        DP_OP_425J2_127_3477_n302), .S(DP_OP_425J2_127_3477_n303) );
  FADDX1_HVT DP_OP_425J2_127_3477_U307 ( .A(DP_OP_425J2_127_3477_n326), .B(
        DP_OP_425J2_127_3477_n324), .CI(DP_OP_425J2_127_3477_n303), .CO(
        DP_OP_425J2_127_3477_n300), .S(DP_OP_425J2_127_3477_n301) );
  FADDX1_HVT DP_OP_425J2_127_3477_U306 ( .A(DP_OP_425J2_127_3477_n1874), .B(
        DP_OP_425J2_127_3477_n320), .CI(DP_OP_425J2_127_3477_n318), .CO(
        DP_OP_425J2_127_3477_n298), .S(DP_OP_425J2_127_3477_n299) );
  FADDX1_HVT DP_OP_425J2_127_3477_U305 ( .A(DP_OP_425J2_127_3477_n316), .B(
        DP_OP_425J2_127_3477_n299), .CI(DP_OP_425J2_127_3477_n314), .CO(
        DP_OP_425J2_127_3477_n296), .S(DP_OP_425J2_127_3477_n297) );
  FADDX1_HVT DP_OP_425J2_127_3477_U304 ( .A(DP_OP_425J2_127_3477_n312), .B(
        DP_OP_425J2_127_3477_n310), .CI(DP_OP_425J2_127_3477_n297), .CO(
        DP_OP_425J2_127_3477_n294), .S(DP_OP_425J2_127_3477_n295) );
  FADDX1_HVT DP_OP_425J2_127_3477_U303 ( .A(DP_OP_425J2_127_3477_n308), .B(
        DP_OP_425J2_127_3477_n295), .CI(DP_OP_425J2_127_3477_n306), .CO(
        DP_OP_425J2_127_3477_n292), .S(DP_OP_425J2_127_3477_n293) );
  FADDX1_HVT DP_OP_425J2_127_3477_U302 ( .A(DP_OP_425J2_127_3477_n304), .B(
        DP_OP_425J2_127_3477_n293), .CI(DP_OP_425J2_127_3477_n302), .CO(
        DP_OP_425J2_127_3477_n290), .S(DP_OP_425J2_127_3477_n291) );
  FADDX1_HVT DP_OP_425J2_127_3477_U300 ( .A(DP_OP_425J2_127_3477_n289), .B(
        DP_OP_425J2_127_3477_n298), .CI(DP_OP_425J2_127_3477_n296), .CO(
        DP_OP_425J2_127_3477_n286), .S(DP_OP_425J2_127_3477_n287) );
  FADDX1_HVT DP_OP_425J2_127_3477_U299 ( .A(DP_OP_425J2_127_3477_n287), .B(
        DP_OP_425J2_127_3477_n294), .CI(DP_OP_425J2_127_3477_n292), .CO(
        DP_OP_425J2_127_3477_n284), .S(DP_OP_425J2_127_3477_n285) );
  FADDX1_HVT DP_OP_425J2_127_3477_U298 ( .A(DP_OP_425J2_127_3477_n1873), .B(
        DP_OP_425J2_127_3477_n288), .CI(DP_OP_425J2_127_3477_n286), .CO(
        DP_OP_425J2_127_3477_n282), .S(DP_OP_425J2_127_3477_n283) );
  FADDX1_HVT DP_OP_425J2_127_3477_U281 ( .A(DP_OP_425J2_127_3477_n1853), .B(
        DP_OP_425J2_127_3477_n1851), .CI(DP_OP_425J2_127_3477_n1849), .CO(
        DP_OP_425J2_127_3477_n219), .S(n_conv2_sum_d[0]) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U280 ( .A1(DP_OP_425J2_127_3477_n1787), 
        .A2(DP_OP_425J2_127_3477_n1789), .Y(DP_OP_425J2_127_3477_n218) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U279 ( .A1(DP_OP_425J2_127_3477_n1789), .A2(
        DP_OP_425J2_127_3477_n1787), .Y(DP_OP_425J2_127_3477_n217) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U273 ( .A1(DP_OP_425J2_127_3477_n1681), 
        .A2(DP_OP_425J2_127_3477_n1683), .Y(DP_OP_425J2_127_3477_n215) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U265 ( .A1(DP_OP_425J2_127_3477_n1527), 
        .A2(DP_OP_425J2_127_3477_n1529), .Y(DP_OP_425J2_127_3477_n210) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U264 ( .A1(DP_OP_425J2_127_3477_n1529), .A2(
        DP_OP_425J2_127_3477_n1527), .Y(DP_OP_425J2_127_3477_n209) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U259 ( .A1(DP_OP_425J2_127_3477_n1351), 
        .A2(DP_OP_425J2_127_3477_n1353), .Y(DP_OP_425J2_127_3477_n207) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U251 ( .A1(DP_OP_425J2_127_3477_n1163), 
        .A2(DP_OP_425J2_127_3477_n1165), .Y(DP_OP_425J2_127_3477_n202) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U250 ( .A1(DP_OP_425J2_127_3477_n1165), .A2(
        DP_OP_425J2_127_3477_n1163), .Y(DP_OP_425J2_127_3477_n201) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U245 ( .A1(DP_OP_425J2_127_3477_n969), .A2(
        DP_OP_425J2_127_3477_n971), .Y(DP_OP_425J2_127_3477_n199) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U237 ( .A1(DP_OP_425J2_127_3477_n773), .A2(
        DP_OP_425J2_127_3477_n968), .Y(DP_OP_425J2_127_3477_n194) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U236 ( .A1(DP_OP_425J2_127_3477_n968), .A2(
        DP_OP_425J2_127_3477_n773), .Y(DP_OP_425J2_127_3477_n193) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U230 ( .A1(DP_OP_425J2_127_3477_n599), .A2(
        DP_OP_425J2_127_3477_n772), .Y(DP_OP_425J2_127_3477_n190) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U229 ( .A1(DP_OP_425J2_127_3477_n772), .A2(
        DP_OP_425J2_127_3477_n599), .Y(DP_OP_425J2_127_3477_n189) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U224 ( .A1(DP_OP_425J2_127_3477_n463), .A2(
        DP_OP_425J2_127_3477_n598), .Y(DP_OP_425J2_127_3477_n187) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U223 ( .A1(DP_OP_425J2_127_3477_n598), .A2(
        DP_OP_425J2_127_3477_n463), .Y(DP_OP_425J2_127_3477_n186) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U219 ( .A1(DP_OP_425J2_127_3477_n189), .A2(
        DP_OP_425J2_127_3477_n186), .Y(DP_OP_425J2_127_3477_n184) );
  AOI21X1_HVT DP_OP_425J2_127_3477_U218 ( .A1(DP_OP_425J2_127_3477_n184), .A2(
        DP_OP_425J2_127_3477_n192), .A3(DP_OP_425J2_127_3477_n185), .Y(
        DP_OP_425J2_127_3477_n183) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U215 ( .A1(DP_OP_425J2_127_3477_n369), .A2(
        DP_OP_425J2_127_3477_n462), .Y(DP_OP_425J2_127_3477_n181) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U214 ( .A1(DP_OP_425J2_127_3477_n462), .A2(
        DP_OP_425J2_127_3477_n369), .Y(DP_OP_425J2_127_3477_n180) );
  AOI21X1_HVT DP_OP_425J2_127_3477_U209 ( .A1(DP_OP_425J2_127_3477_n182), .A2(
        DP_OP_425J2_127_3477_n241), .A3(DP_OP_425J2_127_3477_n179), .Y(
        DP_OP_425J2_127_3477_n177) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U207 ( .A1(DP_OP_425J2_127_3477_n323), .A2(
        DP_OP_425J2_127_3477_n368), .Y(DP_OP_425J2_127_3477_n176) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U206 ( .A1(DP_OP_425J2_127_3477_n368), .A2(
        DP_OP_425J2_127_3477_n323), .Y(DP_OP_425J2_127_3477_n175) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U204 ( .A1(DP_OP_425J2_127_3477_n240), .A2(
        DP_OP_425J2_127_3477_n176), .Y(DP_OP_425J2_127_3477_n25) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U202 ( .A1(DP_OP_425J2_127_3477_n175), .A2(
        DP_OP_425J2_127_3477_n180), .Y(DP_OP_425J2_127_3477_n173) );
  AOI21X1_HVT DP_OP_425J2_127_3477_U201 ( .A1(DP_OP_425J2_127_3477_n182), .A2(
        DP_OP_425J2_127_3477_n173), .A3(DP_OP_425J2_127_3477_n174), .Y(
        DP_OP_425J2_127_3477_n172) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U199 ( .A1(DP_OP_425J2_127_3477_n301), .A2(
        DP_OP_425J2_127_3477_n322), .Y(DP_OP_425J2_127_3477_n171) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U198 ( .A1(DP_OP_425J2_127_3477_n322), .A2(
        DP_OP_425J2_127_3477_n301), .Y(DP_OP_425J2_127_3477_n170) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U193 ( .A1(DP_OP_425J2_127_3477_n300), .A2(
        DP_OP_425J2_127_3477_n291), .Y(DP_OP_425J2_127_3477_n168) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U192 ( .A1(DP_OP_425J2_127_3477_n291), .A2(
        DP_OP_425J2_127_3477_n300), .Y(DP_OP_425J2_127_3477_n167) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U188 ( .A1(DP_OP_425J2_127_3477_n167), .A2(
        DP_OP_425J2_127_3477_n170), .Y(DP_OP_425J2_127_3477_n165) );
  AOI21X1_HVT DP_OP_425J2_127_3477_U187 ( .A1(DP_OP_425J2_127_3477_n174), .A2(
        DP_OP_425J2_127_3477_n165), .A3(DP_OP_425J2_127_3477_n166), .Y(
        DP_OP_425J2_127_3477_n164) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U186 ( .A1(DP_OP_425J2_127_3477_n173), .A2(
        DP_OP_425J2_127_3477_n165), .Y(DP_OP_425J2_127_3477_n163) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U182 ( .A1(DP_OP_425J2_127_3477_n290), .A2(
        DP_OP_425J2_127_3477_n285), .Y(DP_OP_425J2_127_3477_n152) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U181 ( .A1(DP_OP_425J2_127_3477_n285), .A2(
        DP_OP_425J2_127_3477_n290), .Y(DP_OP_425J2_127_3477_n151) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U168 ( .A1(DP_OP_425J2_127_3477_n284), .A2(
        DP_OP_425J2_127_3477_n283), .Y(DP_OP_425J2_127_3477_n149) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U167 ( .A1(DP_OP_425J2_127_3477_n283), .A2(
        DP_OP_425J2_127_3477_n284), .Y(DP_OP_425J2_127_3477_n148) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U161 ( .A1(DP_OP_425J2_127_3477_n237), .A2(
        DP_OP_425J2_127_3477_n236), .Y(DP_OP_425J2_127_3477_n144) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U156 ( .A1(DP_OP_425J2_127_3477_n282), .A2(
        DP_OP_425J2_127_3477_n281), .Y(DP_OP_425J2_127_3477_n140) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U153 ( .A1(DP_OP_425J2_127_3477_n235), .A2(
        DP_OP_425J2_127_3477_n140), .Y(DP_OP_425J2_127_3477_n20) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U146 ( .A1(DP_OP_425J2_127_3477_n279), .A2(
        DP_OP_425J2_127_3477_n280), .Y(DP_OP_425J2_127_3477_n133) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U145 ( .A1(DP_OP_425J2_127_3477_n280), .A2(
        DP_OP_425J2_127_3477_n279), .Y(DP_OP_425J2_127_3477_n132) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U143 ( .A1(DP_OP_425J2_127_3477_n234), .A2(
        DP_OP_425J2_127_3477_n133), .Y(DP_OP_425J2_127_3477_n19) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U140 ( .A1(DP_OP_425J2_127_3477_n277), .A2(
        DP_OP_425J2_127_3477_n278), .Y(DP_OP_425J2_127_3477_n130) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U139 ( .A1(DP_OP_425J2_127_3477_n278), .A2(
        DP_OP_425J2_127_3477_n277), .Y(DP_OP_425J2_127_3477_n129) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U137 ( .A1(DP_OP_425J2_127_3477_n233), .A2(
        DP_OP_425J2_127_3477_n130), .Y(DP_OP_425J2_127_3477_n18) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U135 ( .A1(DP_OP_425J2_127_3477_n129), .A2(
        DP_OP_425J2_127_3477_n132), .Y(DP_OP_425J2_127_3477_n127) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U130 ( .A1(DP_OP_425J2_127_3477_n275), .A2(
        DP_OP_425J2_127_3477_n276), .Y(DP_OP_425J2_127_3477_n123) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U127 ( .A1(n462), .A2(
        DP_OP_425J2_127_3477_n123), .Y(DP_OP_425J2_127_3477_n17) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U123 ( .A1(DP_OP_425J2_127_3477_n127), .A2(
        n462), .Y(DP_OP_425J2_127_3477_n118) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U120 ( .A1(DP_OP_425J2_127_3477_n273), .A2(
        DP_OP_425J2_127_3477_n274), .Y(DP_OP_425J2_127_3477_n116) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U119 ( .A1(DP_OP_425J2_127_3477_n274), .A2(
        DP_OP_425J2_127_3477_n273), .Y(DP_OP_425J2_127_3477_n115) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U110 ( .A1(DP_OP_425J2_127_3477_n271), .A2(
        DP_OP_425J2_127_3477_n272), .Y(DP_OP_425J2_127_3477_n109) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U103 ( .A1(DP_OP_425J2_127_3477_n113), .A2(
        n461), .Y(DP_OP_425J2_127_3477_n104) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U100 ( .A1(DP_OP_425J2_127_3477_n269), .A2(
        DP_OP_425J2_127_3477_n270), .Y(DP_OP_425J2_127_3477_n102) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U99 ( .A1(DP_OP_425J2_127_3477_n270), .A2(
        DP_OP_425J2_127_3477_n269), .Y(DP_OP_425J2_127_3477_n101) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U90 ( .A1(DP_OP_425J2_127_3477_n267), .A2(
        DP_OP_425J2_127_3477_n268), .Y(DP_OP_425J2_127_3477_n95) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U83 ( .A1(DP_OP_425J2_127_3477_n99), .A2(
        n457), .Y(DP_OP_425J2_127_3477_n90) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U80 ( .A1(DP_OP_425J2_127_3477_n265), .A2(
        DP_OP_425J2_127_3477_n266), .Y(DP_OP_425J2_127_3477_n88) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U79 ( .A1(DP_OP_425J2_127_3477_n266), .A2(
        DP_OP_425J2_127_3477_n265), .Y(DP_OP_425J2_127_3477_n87) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U70 ( .A1(DP_OP_425J2_127_3477_n263), .A2(
        DP_OP_425J2_127_3477_n264), .Y(DP_OP_425J2_127_3477_n81) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U63 ( .A1(DP_OP_425J2_127_3477_n85), .A2(
        n456), .Y(DP_OP_425J2_127_3477_n76) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U61 ( .A1(DP_OP_425J2_127_3477_n76), .A2(
        DP_OP_425J2_127_3477_n137), .Y(DP_OP_425J2_127_3477_n74) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U56 ( .A1(DP_OP_425J2_127_3477_n261), .A2(
        DP_OP_425J2_127_3477_n262), .Y(DP_OP_425J2_127_3477_n70) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U49 ( .A1(DP_OP_425J2_127_3477_n74), .A2(
        n455), .Y(DP_OP_425J2_127_3477_n65) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U45 ( .A1(DP_OP_425J2_127_3477_n237), .A2(
        DP_OP_425J2_127_3477_n63), .Y(DP_OP_425J2_127_3477_n61) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U42 ( .A1(DP_OP_425J2_127_3477_n259), .A2(
        DP_OP_425J2_127_3477_n260), .Y(DP_OP_425J2_127_3477_n59) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U41 ( .A1(DP_OP_425J2_127_3477_n260), .A2(
        DP_OP_425J2_127_3477_n259), .Y(DP_OP_425J2_127_3477_n58) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U32 ( .A1(DP_OP_425J2_127_3477_n257), .A2(
        DP_OP_425J2_127_3477_n258), .Y(DP_OP_425J2_127_3477_n52) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U25 ( .A1(DP_OP_425J2_127_3477_n56), .A2(
        n454), .Y(DP_OP_425J2_127_3477_n47) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U22 ( .A1(DP_OP_425J2_127_3477_n255), .A2(
        DP_OP_425J2_127_3477_n256), .Y(DP_OP_425J2_127_3477_n45) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U21 ( .A1(DP_OP_425J2_127_3477_n256), .A2(
        DP_OP_425J2_127_3477_n255), .Y(DP_OP_425J2_127_3477_n44) );
  AOI21X1_HVT DP_OP_425J2_127_3477_U16 ( .A1(DP_OP_425J2_127_3477_n162), .A2(
        DP_OP_425J2_127_3477_n42), .A3(DP_OP_425J2_127_3477_n43), .Y(
        DP_OP_425J2_127_3477_n41) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U14 ( .A1(DP_OP_425J2_127_3477_n253), .A2(
        DP_OP_425J2_127_3477_n254), .Y(DP_OP_425J2_127_3477_n40) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U13 ( .A1(DP_OP_425J2_127_3477_n254), .A2(
        DP_OP_425J2_127_3477_n253), .Y(DP_OP_425J2_127_3477_n39) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U8 ( .A1(n463), .A2(
        DP_OP_425J2_127_3477_n252), .Y(DP_OP_425J2_127_3477_n37) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U96 ( .A1(DP_OP_424J2_126_3477_n101), .A2(
        DP_OP_424J2_126_3477_n105), .A3(DP_OP_424J2_126_3477_n102), .Y(
        DP_OP_424J2_126_3477_n100) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U261 ( .A1(DP_OP_424J2_126_3477_n211), .A2(
        DP_OP_424J2_126_3477_n209), .A3(DP_OP_424J2_126_3477_n210), .Y(
        DP_OP_424J2_126_3477_n208) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U76 ( .A1(DP_OP_424J2_126_3477_n87), .A2(
        DP_OP_424J2_126_3477_n91), .A3(DP_OP_424J2_126_3477_n88), .Y(
        DP_OP_424J2_126_3477_n86) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U116 ( .A1(DP_OP_424J2_126_3477_n115), .A2(
        DP_OP_424J2_126_3477_n119), .A3(DP_OP_424J2_126_3477_n116), .Y(
        DP_OP_424J2_126_3477_n114) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U136 ( .A1(DP_OP_424J2_126_3477_n133), .A2(
        DP_OP_424J2_126_3477_n129), .A3(DP_OP_424J2_126_3477_n130), .Y(
        DP_OP_424J2_126_3477_n128) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U275 ( .A1(DP_OP_424J2_126_3477_n4), .A2(
        DP_OP_424J2_126_3477_n217), .A3(DP_OP_424J2_126_3477_n218), .Y(
        DP_OP_424J2_126_3477_n216) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1111 ( .A1(n501), .A2(n385), .Y(
        DP_OP_424J2_126_3477_n288) );
  XNOR2X1_HVT DP_OP_424J2_126_3477_U737 ( .A1(DP_OP_424J2_126_3477_n2452), 
        .A2(DP_OP_424J2_126_3477_n2979), .Y(DP_OP_424J2_126_3477_n1161) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1109 ( .A1(n338), .A2(
        DP_OP_425J2_127_3477_n2), .Y(DP_OP_424J2_126_3477_n280) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2239 ( .A1(DP_OP_424J2_126_3477_n3006), .A2(
        DP_OP_425J2_127_3477_n3017), .Y(DP_OP_424J2_126_3477_n2998) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2231 ( .A1(DP_OP_424J2_126_3477_n3006), .A2(
        DP_OP_424J2_126_3477_n3016), .Y(DP_OP_424J2_126_3477_n2990) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2223 ( .A1(DP_OP_424J2_126_3477_n3006), .A2(
        DP_OP_424J2_126_3477_n3015), .Y(DP_OP_424J2_126_3477_n2982) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2222 ( .A1(DP_OP_424J2_126_3477_n3013), .A2(
        DP_OP_423J2_125_3477_n3014), .Y(DP_OP_424J2_126_3477_n1678) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2221 ( .A1(DP_OP_424J2_126_3477_n3012), .A2(
        DP_OP_425J2_127_3477_n3014), .Y(DP_OP_424J2_126_3477_n2981) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2220 ( .A1(DP_OP_424J2_126_3477_n3011), .A2(
        DP_OP_422J2_124_3477_n3014), .Y(DP_OP_424J2_126_3477_n2980) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2219 ( .A1(DP_OP_424J2_126_3477_n3010), .A2(
        DP_OP_422J2_124_3477_n3014), .Y(DP_OP_424J2_126_3477_n2979) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2218 ( .A1(DP_OP_424J2_126_3477_n3009), .A2(
        DP_OP_425J2_127_3477_n3014), .Y(DP_OP_424J2_126_3477_n2978) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2217 ( .A1(DP_OP_424J2_126_3477_n3008), .A2(
        DP_OP_423J2_125_3477_n3014), .Y(DP_OP_424J2_126_3477_n770) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2216 ( .A1(DP_OP_424J2_126_3477_n3007), .A2(
        DP_OP_422J2_124_3477_n3014), .Y(DP_OP_424J2_126_3477_n2977) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2215 ( .A1(DP_OP_424J2_126_3477_n3006), 
        .A2(DP_OP_423J2_125_3477_n3014), .Y(DP_OP_424J2_126_3477_n2976) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2195 ( .A1(DP_OP_424J2_126_3477_n2964), .A2(
        DP_OP_424J2_126_3477_n2975), .Y(DP_OP_424J2_126_3477_n2956) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2187 ( .A1(DP_OP_424J2_126_3477_n2964), .A2(
        DP_OP_425J2_127_3477_n2974), .Y(DP_OP_424J2_126_3477_n2948) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2179 ( .A1(DP_OP_424J2_126_3477_n2964), .A2(
        DP_OP_425J2_127_3477_n2973), .Y(DP_OP_424J2_126_3477_n2940) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2178 ( .A1(DP_OP_425J2_127_3477_n2003), .A2(
        DP_OP_423J2_125_3477_n2972), .Y(DP_OP_424J2_126_3477_n2939) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2177 ( .A1(DP_OP_424J2_126_3477_n2970), .A2(
        DP_OP_422J2_124_3477_n2972), .Y(DP_OP_424J2_126_3477_n2938) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2176 ( .A1(DP_OP_424J2_126_3477_n2969), .A2(
        DP_OP_425J2_127_3477_n2972), .Y(DP_OP_424J2_126_3477_n2937) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2175 ( .A1(DP_OP_425J2_127_3477_n2000), .A2(
        DP_OP_425J2_127_3477_n2972), .Y(DP_OP_424J2_126_3477_n2936) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2174 ( .A1(DP_OP_424J2_126_3477_n2967), .A2(
        DP_OP_423J2_125_3477_n2972), .Y(DP_OP_424J2_126_3477_n2935) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2173 ( .A1(DP_OP_425J2_127_3477_n1998), .A2(
        DP_OP_422J2_124_3477_n2972), .Y(DP_OP_424J2_126_3477_n2934) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2172 ( .A1(DP_OP_425J2_127_3477_n1997), .A2(
        DP_OP_422J2_124_3477_n2972), .Y(DP_OP_424J2_126_3477_n2933) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2171 ( .A1(DP_OP_424J2_126_3477_n2964), 
        .A2(DP_OP_423J2_125_3477_n2972), .Y(DP_OP_424J2_126_3477_n2932) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2151 ( .A1(DP_OP_424J2_126_3477_n2920), .A2(
        DP_OP_425J2_127_3477_n2931), .Y(DP_OP_424J2_126_3477_n2912) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2143 ( .A1(DP_OP_424J2_126_3477_n2920), .A2(
        DP_OP_422J2_124_3477_n2930), .Y(DP_OP_424J2_126_3477_n2904) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2135 ( .A1(DP_OP_424J2_126_3477_n2920), .A2(
        DP_OP_424J2_126_3477_n2929), .Y(DP_OP_424J2_126_3477_n2896) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2134 ( .A1(DP_OP_424J2_126_3477_n2927), .A2(
        DP_OP_422J2_124_3477_n2928), .Y(DP_OP_424J2_126_3477_n2895) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2133 ( .A1(DP_OP_424J2_126_3477_n2926), .A2(
        DP_OP_425J2_127_3477_n2928), .Y(DP_OP_424J2_126_3477_n2894) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2132 ( .A1(DP_OP_424J2_126_3477_n2925), .A2(
        DP_OP_422J2_124_3477_n2928), .Y(DP_OP_424J2_126_3477_n2893) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2131 ( .A1(DP_OP_424J2_126_3477_n2924), .A2(
        DP_OP_423J2_125_3477_n2928), .Y(DP_OP_424J2_126_3477_n2892) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2130 ( .A1(DP_OP_424J2_126_3477_n2923), .A2(
        DP_OP_423J2_125_3477_n2928), .Y(DP_OP_424J2_126_3477_n2891) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2129 ( .A1(DP_OP_424J2_126_3477_n2922), .A2(
        DP_OP_425J2_127_3477_n2928), .Y(DP_OP_424J2_126_3477_n2890) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2128 ( .A1(DP_OP_424J2_126_3477_n2921), .A2(
        DP_OP_422J2_124_3477_n2928), .Y(DP_OP_424J2_126_3477_n2889) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2127 ( .A1(DP_OP_424J2_126_3477_n2920), 
        .A2(DP_OP_423J2_125_3477_n2928), .Y(DP_OP_424J2_126_3477_n2888) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2107 ( .A1(DP_OP_425J2_127_3477_n2084), .A2(
        DP_OP_424J2_126_3477_n2887), .Y(DP_OP_424J2_126_3477_n2868) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2099 ( .A1(DP_OP_425J2_127_3477_n2084), .A2(
        DP_OP_424J2_126_3477_n2886), .Y(DP_OP_424J2_126_3477_n2860) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2092 ( .A1(DP_OP_424J2_126_3477_n2877), 
        .A2(DP_OP_424J2_126_3477_n2885), .Y(DP_OP_424J2_126_3477_n2853) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2091 ( .A1(DP_OP_423J2_125_3477_n2964), .A2(
        DP_OP_424J2_126_3477_n2885), .Y(DP_OP_424J2_126_3477_n2852) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2090 ( .A1(DP_OP_424J2_126_3477_n2883), .A2(
        DP_OP_422J2_124_3477_n2884), .Y(DP_OP_424J2_126_3477_n2851) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2089 ( .A1(DP_OP_423J2_125_3477_n2970), .A2(
        DP_OP_422J2_124_3477_n2884), .Y(DP_OP_424J2_126_3477_n2850) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2088 ( .A1(DP_OP_423J2_125_3477_n2969), .A2(
        DP_OP_423J2_125_3477_n2884), .Y(DP_OP_424J2_126_3477_n2849) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2087 ( .A1(DP_OP_424J2_126_3477_n2880), .A2(
        DP_OP_425J2_127_3477_n2884), .Y(DP_OP_424J2_126_3477_n2848) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2086 ( .A1(DP_OP_425J2_127_3477_n2087), .A2(
        DP_OP_425J2_127_3477_n2884), .Y(DP_OP_424J2_126_3477_n2847) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2085 ( .A1(DP_OP_424J2_126_3477_n2878), .A2(
        DP_OP_423J2_125_3477_n2884), .Y(DP_OP_424J2_126_3477_n2846) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2084 ( .A1(DP_OP_424J2_126_3477_n2877), .A2(
        DP_OP_423J2_125_3477_n2884), .Y(DP_OP_424J2_126_3477_n2845) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2083 ( .A1(DP_OP_423J2_125_3477_n2964), 
        .A2(DP_OP_422J2_124_3477_n2884), .Y(DP_OP_424J2_126_3477_n2844) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2063 ( .A1(DP_OP_423J2_125_3477_n2920), .A2(
        DP_OP_422J2_124_3477_n2843), .Y(DP_OP_424J2_126_3477_n2824) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2055 ( .A1(DP_OP_423J2_125_3477_n2920), .A2(
        DP_OP_425J2_127_3477_n2842), .Y(DP_OP_424J2_126_3477_n2816) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2048 ( .A1(DP_OP_424J2_126_3477_n2833), 
        .A2(DP_OP_423J2_125_3477_n2841), .Y(DP_OP_424J2_126_3477_n2809) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2047 ( .A1(DP_OP_425J2_127_3477_n2128), .A2(
        DP_OP_423J2_125_3477_n2841), .Y(DP_OP_424J2_126_3477_n2808) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2046 ( .A1(DP_OP_425J2_127_3477_n2135), .A2(
        DP_OP_423J2_125_3477_n2840), .Y(DP_OP_424J2_126_3477_n2807) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2045 ( .A1(DP_OP_425J2_127_3477_n2134), .A2(
        DP_OP_423J2_125_3477_n2840), .Y(DP_OP_424J2_126_3477_n2806) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2044 ( .A1(DP_OP_424J2_126_3477_n2837), .A2(
        DP_OP_425J2_127_3477_n2840), .Y(DP_OP_424J2_126_3477_n2805) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2043 ( .A1(DP_OP_422J2_124_3477_n2000), .A2(
        DP_OP_425J2_127_3477_n2840), .Y(DP_OP_424J2_126_3477_n2804) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2042 ( .A1(DP_OP_424J2_126_3477_n2835), .A2(
        DP_OP_422J2_124_3477_n2840), .Y(DP_OP_424J2_126_3477_n2803) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2041 ( .A1(DP_OP_424J2_126_3477_n2834), .A2(
        DP_OP_422J2_124_3477_n2840), .Y(DP_OP_424J2_126_3477_n2802) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2040 ( .A1(DP_OP_424J2_126_3477_n2833), .A2(
        DP_OP_423J2_125_3477_n2840), .Y(DP_OP_424J2_126_3477_n2801) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2039 ( .A1(DP_OP_425J2_127_3477_n2128), 
        .A2(DP_OP_422J2_124_3477_n2840), .Y(DP_OP_424J2_126_3477_n2800) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2019 ( .A1(DP_OP_422J2_124_3477_n2040), .A2(
        DP_OP_424J2_126_3477_n2799), .Y(DP_OP_424J2_126_3477_n2780) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2011 ( .A1(DP_OP_422J2_124_3477_n2040), .A2(
        DP_OP_425J2_127_3477_n2798), .Y(DP_OP_424J2_126_3477_n2772) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2004 ( .A1(DP_OP_424J2_126_3477_n2789), 
        .A2(DP_OP_424J2_126_3477_n2797), .Y(DP_OP_424J2_126_3477_n2765) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2003 ( .A1(DP_OP_422J2_124_3477_n2040), .A2(
        DP_OP_424J2_126_3477_n2797), .Y(DP_OP_424J2_126_3477_n2764) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2002 ( .A1(DP_OP_424J2_126_3477_n2795), .A2(
        DP_OP_422J2_124_3477_n2796), .Y(DP_OP_424J2_126_3477_n2763) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2001 ( .A1(DP_OP_424J2_126_3477_n2794), .A2(
        DP_OP_425J2_127_3477_n2796), .Y(DP_OP_424J2_126_3477_n2762) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2000 ( .A1(DP_OP_424J2_126_3477_n2793), .A2(
        DP_OP_423J2_125_3477_n2796), .Y(DP_OP_424J2_126_3477_n2761) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1999 ( .A1(DP_OP_423J2_125_3477_n2880), .A2(
        DP_OP_422J2_124_3477_n2796), .Y(DP_OP_424J2_126_3477_n2760) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1998 ( .A1(DP_OP_424J2_126_3477_n2791), .A2(
        DP_OP_423J2_125_3477_n2796), .Y(DP_OP_424J2_126_3477_n2759) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1997 ( .A1(DP_OP_424J2_126_3477_n2790), .A2(
        DP_OP_425J2_127_3477_n2796), .Y(DP_OP_424J2_126_3477_n2758) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1996 ( .A1(DP_OP_424J2_126_3477_n2789), .A2(
        DP_OP_422J2_124_3477_n2796), .Y(DP_OP_424J2_126_3477_n2757) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1995 ( .A1(DP_OP_422J2_124_3477_n2040), 
        .A2(DP_OP_425J2_127_3477_n2796), .Y(DP_OP_424J2_126_3477_n2756) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1982 ( .A1(DP_OP_424J2_126_3477_n2751), 
        .A2(DP_OP_424J2_126_3477_n2755), .Y(DP_OP_424J2_126_3477_n2743) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1981 ( .A1(DP_OP_424J2_126_3477_n2750), 
        .A2(DP_OP_424J2_126_3477_n2755), .Y(DP_OP_424J2_126_3477_n2742) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1980 ( .A1(DP_OP_424J2_126_3477_n2749), 
        .A2(DP_OP_424J2_126_3477_n2755), .Y(DP_OP_424J2_126_3477_n2741) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1979 ( .A1(DP_OP_425J2_127_3477_n2220), 
        .A2(DP_OP_424J2_126_3477_n2755), .Y(DP_OP_424J2_126_3477_n2740) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1978 ( .A1(DP_OP_424J2_126_3477_n2747), 
        .A2(DP_OP_424J2_126_3477_n2755), .Y(DP_OP_424J2_126_3477_n2739) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1977 ( .A1(DP_OP_423J2_125_3477_n2834), 
        .A2(DP_OP_424J2_126_3477_n2755), .Y(DP_OP_424J2_126_3477_n2738) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1976 ( .A1(DP_OP_424J2_126_3477_n2745), 
        .A2(DP_OP_424J2_126_3477_n2755), .Y(DP_OP_424J2_126_3477_n2737) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1975 ( .A1(DP_OP_425J2_127_3477_n2216), .A2(
        DP_OP_424J2_126_3477_n2755), .Y(DP_OP_424J2_126_3477_n2736) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1968 ( .A1(DP_OP_424J2_126_3477_n2745), 
        .A2(DP_OP_425J2_127_3477_n2754), .Y(DP_OP_424J2_126_3477_n2729) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1967 ( .A1(DP_OP_422J2_124_3477_n2084), .A2(
        DP_OP_423J2_125_3477_n2754), .Y(DP_OP_424J2_126_3477_n2728) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1959 ( .A1(DP_OP_425J2_127_3477_n2216), .A2(
        DP_OP_424J2_126_3477_n2753), .Y(DP_OP_424J2_126_3477_n2720) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1958 ( .A1(DP_OP_424J2_126_3477_n2751), .A2(
        DP_OP_425J2_127_3477_n2752), .Y(DP_OP_424J2_126_3477_n2719) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1957 ( .A1(DP_OP_424J2_126_3477_n2750), .A2(
        DP_OP_423J2_125_3477_n2752), .Y(DP_OP_424J2_126_3477_n2718) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1956 ( .A1(DP_OP_424J2_126_3477_n2749), .A2(
        DP_OP_423J2_125_3477_n2752), .Y(DP_OP_424J2_126_3477_n2717) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1955 ( .A1(DP_OP_422J2_124_3477_n2088), .A2(
        DP_OP_422J2_124_3477_n2752), .Y(DP_OP_424J2_126_3477_n2716) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1954 ( .A1(DP_OP_424J2_126_3477_n2747), .A2(
        DP_OP_422J2_124_3477_n2752), .Y(DP_OP_424J2_126_3477_n2715) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1953 ( .A1(DP_OP_423J2_125_3477_n2834), .A2(
        DP_OP_425J2_127_3477_n2752), .Y(DP_OP_424J2_126_3477_n2714) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1952 ( .A1(DP_OP_424J2_126_3477_n2745), .A2(
        DP_OP_425J2_127_3477_n2752), .Y(DP_OP_424J2_126_3477_n2713) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1951 ( .A1(DP_OP_425J2_127_3477_n2216), 
        .A2(DP_OP_422J2_124_3477_n2752), .Y(DP_OP_424J2_126_3477_n2712) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1931 ( .A1(DP_OP_424J2_126_3477_n2700), .A2(
        DP_OP_424J2_126_3477_n2711), .Y(DP_OP_424J2_126_3477_n2692) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1923 ( .A1(DP_OP_424J2_126_3477_n2700), .A2(
        DP_OP_423J2_125_3477_n2710), .Y(DP_OP_424J2_126_3477_n2684) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1915 ( .A1(DP_OP_424J2_126_3477_n2700), .A2(
        DP_OP_425J2_127_3477_n2709), .Y(DP_OP_424J2_126_3477_n2676) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1914 ( .A1(DP_OP_422J2_124_3477_n2135), .A2(
        DP_OP_422J2_124_3477_n2708), .Y(DP_OP_424J2_126_3477_n2675) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1913 ( .A1(DP_OP_422J2_124_3477_n2134), .A2(
        DP_OP_423J2_125_3477_n2708), .Y(DP_OP_424J2_126_3477_n2674) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1912 ( .A1(DP_OP_424J2_126_3477_n2705), .A2(
        DP_OP_422J2_124_3477_n2708), .Y(DP_OP_424J2_126_3477_n2673) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1911 ( .A1(DP_OP_422J2_124_3477_n2132), .A2(
        DP_OP_425J2_127_3477_n2708), .Y(DP_OP_424J2_126_3477_n2672) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1910 ( .A1(DP_OP_424J2_126_3477_n2703), .A2(
        DP_OP_422J2_124_3477_n2708), .Y(DP_OP_424J2_126_3477_n2671) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1909 ( .A1(DP_OP_422J2_124_3477_n2130), .A2(
        DP_OP_425J2_127_3477_n2708), .Y(DP_OP_424J2_126_3477_n2670) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1908 ( .A1(DP_OP_422J2_124_3477_n2129), .A2(
        DP_OP_425J2_127_3477_n2708), .Y(DP_OP_424J2_126_3477_n2669) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1907 ( .A1(DP_OP_424J2_126_3477_n2700), 
        .A2(DP_OP_423J2_125_3477_n2708), .Y(DP_OP_424J2_126_3477_n2668) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1887 ( .A1(DP_OP_425J2_127_3477_n2304), .A2(
        DP_OP_422J2_124_3477_n2667), .Y(DP_OP_424J2_126_3477_n2648) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1879 ( .A1(DP_OP_422J2_124_3477_n2172), .A2(
        DP_OP_424J2_126_3477_n2666), .Y(DP_OP_424J2_126_3477_n2640) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1871 ( .A1(DP_OP_422J2_124_3477_n2172), .A2(
        DP_OP_424J2_126_3477_n2665), .Y(DP_OP_424J2_126_3477_n2632) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1870 ( .A1(DP_OP_424J2_126_3477_n2663), .A2(
        DP_OP_422J2_124_3477_n2664), .Y(DP_OP_424J2_126_3477_n2631) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1869 ( .A1(DP_OP_423J2_125_3477_n2750), .A2(
        DP_OP_423J2_125_3477_n2664), .Y(DP_OP_424J2_126_3477_n2630) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1868 ( .A1(DP_OP_423J2_125_3477_n2749), .A2(
        DP_OP_422J2_124_3477_n2664), .Y(DP_OP_424J2_126_3477_n2629) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1867 ( .A1(DP_OP_423J2_125_3477_n2748), .A2(
        DP_OP_425J2_127_3477_n2664), .Y(DP_OP_424J2_126_3477_n2628) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1866 ( .A1(DP_OP_425J2_127_3477_n2307), .A2(
        DP_OP_425J2_127_3477_n2664), .Y(DP_OP_424J2_126_3477_n2627) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1865 ( .A1(DP_OP_424J2_126_3477_n2658), .A2(
        DP_OP_422J2_124_3477_n2664), .Y(DP_OP_424J2_126_3477_n2626) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1864 ( .A1(DP_OP_425J2_127_3477_n2305), .A2(
        DP_OP_425J2_127_3477_n2664), .Y(DP_OP_424J2_126_3477_n2625) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1863 ( .A1(DP_OP_422J2_124_3477_n2172), 
        .A2(DP_OP_423J2_125_3477_n2664), .Y(DP_OP_424J2_126_3477_n2624) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1843 ( .A1(DP_OP_424J2_126_3477_n2612), .A2(
        DP_OP_424J2_126_3477_n2623), .Y(DP_OP_424J2_126_3477_n2604) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1842 ( .A1(DP_OP_423J2_125_3477_n2707), 
        .A2(DP_OP_424J2_126_3477_n2622), .Y(DP_OP_424J2_126_3477_n2603) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1841 ( .A1(DP_OP_424J2_126_3477_n2618), 
        .A2(DP_OP_424J2_126_3477_n2622), .Y(DP_OP_424J2_126_3477_n2602) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1840 ( .A1(DP_OP_425J2_127_3477_n2353), 
        .A2(DP_OP_424J2_126_3477_n2622), .Y(DP_OP_424J2_126_3477_n2601) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1839 ( .A1(DP_OP_424J2_126_3477_n2616), 
        .A2(DP_OP_424J2_126_3477_n2622), .Y(DP_OP_424J2_126_3477_n2600) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1838 ( .A1(DP_OP_425J2_127_3477_n2351), 
        .A2(DP_OP_424J2_126_3477_n2622), .Y(DP_OP_424J2_126_3477_n2599) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1837 ( .A1(DP_OP_423J2_125_3477_n2702), 
        .A2(DP_OP_424J2_126_3477_n2622), .Y(DP_OP_424J2_126_3477_n2598) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1836 ( .A1(DP_OP_424J2_126_3477_n2613), 
        .A2(DP_OP_424J2_126_3477_n2622), .Y(DP_OP_424J2_126_3477_n2597) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1835 ( .A1(DP_OP_424J2_126_3477_n2612), .A2(
        DP_OP_424J2_126_3477_n2622), .Y(DP_OP_424J2_126_3477_n2596) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1827 ( .A1(DP_OP_424J2_126_3477_n2612), .A2(
        DP_OP_425J2_127_3477_n2621), .Y(DP_OP_424J2_126_3477_n2588) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1825 ( .A1(DP_OP_424J2_126_3477_n2618), .A2(
        DP_OP_424J2_126_3477_n2620), .Y(DP_OP_424J2_126_3477_n2586) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1824 ( .A1(DP_OP_423J2_125_3477_n2705), .A2(
        DP_OP_424J2_126_3477_n2620), .Y(DP_OP_424J2_126_3477_n2585) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1823 ( .A1(DP_OP_424J2_126_3477_n2616), .A2(
        DP_OP_424J2_126_3477_n2620), .Y(DP_OP_424J2_126_3477_n2584) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1822 ( .A1(DP_OP_425J2_127_3477_n2351), .A2(
        DP_OP_424J2_126_3477_n2620), .Y(DP_OP_424J2_126_3477_n2583) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1821 ( .A1(DP_OP_422J2_124_3477_n2218), .A2(
        DP_OP_424J2_126_3477_n2620), .Y(DP_OP_424J2_126_3477_n2582) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1820 ( .A1(DP_OP_424J2_126_3477_n2613), .A2(
        DP_OP_424J2_126_3477_n2620), .Y(DP_OP_424J2_126_3477_n2581) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1819 ( .A1(DP_OP_424J2_126_3477_n2612), 
        .A2(DP_OP_424J2_126_3477_n2620), .Y(DP_OP_424J2_126_3477_n2580) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1800 ( .A1(DP_OP_424J2_126_3477_n2569), 
        .A2(DP_OP_425J2_127_3477_n2579), .Y(DP_OP_424J2_126_3477_n2561) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1799 ( .A1(DP_OP_423J2_125_3477_n2656), .A2(
        DP_OP_425J2_127_3477_n2579), .Y(DP_OP_424J2_126_3477_n2560) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1791 ( .A1(DP_OP_422J2_124_3477_n2260), .A2(
        DP_OP_424J2_126_3477_n2578), .Y(DP_OP_424J2_126_3477_n2552) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1783 ( .A1(DP_OP_422J2_124_3477_n2260), .A2(
        DP_OP_423J2_125_3477_n2577), .Y(DP_OP_424J2_126_3477_n2544) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1782 ( .A1(DP_OP_422J2_124_3477_n2267), .A2(
        DP_OP_422J2_124_3477_n2576), .Y(DP_OP_424J2_126_3477_n2543) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1781 ( .A1(DP_OP_425J2_127_3477_n2398), .A2(
        DP_OP_422J2_124_3477_n2576), .Y(DP_OP_424J2_126_3477_n2542) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1780 ( .A1(DP_OP_422J2_124_3477_n2265), .A2(
        DP_OP_425J2_127_3477_n2576), .Y(DP_OP_424J2_126_3477_n2541) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1779 ( .A1(DP_OP_424J2_126_3477_n2572), .A2(
        DP_OP_423J2_125_3477_n2576), .Y(DP_OP_424J2_126_3477_n2540) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1778 ( .A1(DP_OP_422J2_124_3477_n2263), .A2(
        DP_OP_425J2_127_3477_n2576), .Y(DP_OP_424J2_126_3477_n2539) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1777 ( .A1(DP_OP_423J2_125_3477_n2658), .A2(
        DP_OP_423J2_125_3477_n2576), .Y(DP_OP_424J2_126_3477_n2538) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1776 ( .A1(DP_OP_424J2_126_3477_n2569), .A2(
        DP_OP_422J2_124_3477_n2576), .Y(DP_OP_424J2_126_3477_n2537) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1775 ( .A1(DP_OP_423J2_125_3477_n2656), 
        .A2(DP_OP_423J2_125_3477_n2576), .Y(DP_OP_424J2_126_3477_n2536) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1755 ( .A1(DP_OP_423J2_125_3477_n2612), .A2(
        DP_OP_425J2_127_3477_n2535), .Y(DP_OP_424J2_126_3477_n2516) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1747 ( .A1(DP_OP_423J2_125_3477_n2612), .A2(
        DP_OP_425J2_127_3477_n2534), .Y(DP_OP_424J2_126_3477_n2508) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1740 ( .A1(DP_OP_422J2_124_3477_n2305), 
        .A2(DP_OP_424J2_126_3477_n2533), .Y(DP_OP_424J2_126_3477_n2501) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1739 ( .A1(DP_OP_422J2_124_3477_n2304), .A2(
        DP_OP_424J2_126_3477_n2533), .Y(DP_OP_424J2_126_3477_n2500) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1738 ( .A1(DP_OP_423J2_125_3477_n2619), .A2(
        DP_OP_424J2_126_3477_n2532), .Y(DP_OP_424J2_126_3477_n2499) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1737 ( .A1(DP_OP_424J2_126_3477_n2530), .A2(
        DP_OP_424J2_126_3477_n2532), .Y(DP_OP_424J2_126_3477_n2498) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1736 ( .A1(DP_OP_423J2_125_3477_n2617), .A2(
        DP_OP_424J2_126_3477_n2532), .Y(DP_OP_424J2_126_3477_n2497) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1735 ( .A1(DP_OP_424J2_126_3477_n2528), .A2(
        DP_OP_424J2_126_3477_n2532), .Y(DP_OP_424J2_126_3477_n2496) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1734 ( .A1(DP_OP_422J2_124_3477_n2307), .A2(
        DP_OP_424J2_126_3477_n2532), .Y(DP_OP_424J2_126_3477_n2495) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1733 ( .A1(DP_OP_424J2_126_3477_n2526), .A2(
        DP_OP_424J2_126_3477_n2532), .Y(DP_OP_424J2_126_3477_n2494) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1732 ( .A1(DP_OP_423J2_125_3477_n2613), .A2(
        DP_OP_424J2_126_3477_n2532), .Y(DP_OP_424J2_126_3477_n2493) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1731 ( .A1(DP_OP_423J2_125_3477_n2612), 
        .A2(DP_OP_424J2_126_3477_n2532), .Y(DP_OP_424J2_126_3477_n2492) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1711 ( .A1(DP_OP_422J2_124_3477_n2348), .A2(
        DP_OP_422J2_124_3477_n2491), .Y(DP_OP_424J2_126_3477_n2472) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1703 ( .A1(DP_OP_422J2_124_3477_n2348), .A2(
        DP_OP_422J2_124_3477_n2490), .Y(DP_OP_424J2_126_3477_n2464) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1695 ( .A1(DP_OP_422J2_124_3477_n2348), .A2(
        DP_OP_424J2_126_3477_n2489), .Y(DP_OP_424J2_126_3477_n2456) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1694 ( .A1(DP_OP_422J2_124_3477_n2355), .A2(
        DP_OP_424J2_126_3477_n2488), .Y(DP_OP_424J2_126_3477_n2455) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1693 ( .A1(DP_OP_422J2_124_3477_n2354), .A2(
        DP_OP_424J2_126_3477_n2488), .Y(DP_OP_424J2_126_3477_n2454) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1692 ( .A1(DP_OP_422J2_124_3477_n2353), .A2(
        DP_OP_424J2_126_3477_n2488), .Y(DP_OP_424J2_126_3477_n2453) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1691 ( .A1(DP_OP_424J2_126_3477_n2484), .A2(
        DP_OP_424J2_126_3477_n2488), .Y(DP_OP_424J2_126_3477_n2452) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1690 ( .A1(DP_OP_422J2_124_3477_n2351), .A2(
        DP_OP_424J2_126_3477_n2488), .Y(DP_OP_424J2_126_3477_n2451) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1689 ( .A1(DP_OP_424J2_126_3477_n2482), .A2(
        DP_OP_424J2_126_3477_n2488), .Y(DP_OP_424J2_126_3477_n2450) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1688 ( .A1(DP_OP_424J2_126_3477_n2481), .A2(
        DP_OP_424J2_126_3477_n2488), .Y(DP_OP_424J2_126_3477_n2449) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1687 ( .A1(DP_OP_422J2_124_3477_n2348), 
        .A2(DP_OP_424J2_126_3477_n2488), .Y(DP_OP_424J2_126_3477_n2448) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1667 ( .A1(DP_OP_422J2_124_3477_n2612), .A2(
        DP_OP_424J2_126_3477_n2447), .Y(DP_OP_424J2_126_3477_n2428) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1659 ( .A1(DP_OP_423J2_125_3477_n2348), .A2(
        DP_OP_424J2_126_3477_n2446), .Y(DP_OP_424J2_126_3477_n2420) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1651 ( .A1(DP_OP_423J2_125_3477_n2348), .A2(
        DP_OP_424J2_126_3477_n2445), .Y(DP_OP_424J2_126_3477_n2412) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1650 ( .A1(DP_OP_423J2_125_3477_n2355), .A2(
        DP_OP_424J2_126_3477_n2444), .Y(DP_OP_424J2_126_3477_n2411) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1649 ( .A1(DP_OP_424J2_126_3477_n2442), .A2(
        DP_OP_424J2_126_3477_n2444), .Y(DP_OP_424J2_126_3477_n2410) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1648 ( .A1(DP_OP_423J2_125_3477_n2353), .A2(
        DP_OP_424J2_126_3477_n2444), .Y(DP_OP_424J2_126_3477_n2409) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1647 ( .A1(DP_OP_425J2_127_3477_n2484), .A2(
        DP_OP_424J2_126_3477_n2444), .Y(DP_OP_424J2_126_3477_n2408) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1646 ( .A1(DP_OP_424J2_126_3477_n2439), .A2(
        DP_OP_424J2_126_3477_n2444), .Y(DP_OP_424J2_126_3477_n2407) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1645 ( .A1(DP_OP_425J2_127_3477_n2482), .A2(
        DP_OP_424J2_126_3477_n2444), .Y(DP_OP_424J2_126_3477_n2406) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1644 ( .A1(DP_OP_425J2_127_3477_n2481), .A2(
        DP_OP_424J2_126_3477_n2444), .Y(DP_OP_424J2_126_3477_n2405) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1643 ( .A1(DP_OP_422J2_124_3477_n2612), 
        .A2(DP_OP_424J2_126_3477_n2444), .Y(DP_OP_424J2_126_3477_n2404) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1623 ( .A1(DP_OP_422J2_124_3477_n2656), .A2(
        DP_OP_423J2_125_3477_n2403), .Y(DP_OP_424J2_126_3477_n2384) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1615 ( .A1(DP_OP_422J2_124_3477_n2656), .A2(
        DP_OP_424J2_126_3477_n2402), .Y(DP_OP_424J2_126_3477_n2376) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1607 ( .A1(DP_OP_423J2_125_3477_n2304), .A2(
        DP_OP_424J2_126_3477_n2401), .Y(DP_OP_424J2_126_3477_n2368) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1606 ( .A1(DP_OP_423J2_125_3477_n2311), .A2(
        DP_OP_423J2_125_3477_n2400), .Y(DP_OP_424J2_126_3477_n2367) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1605 ( .A1(DP_OP_425J2_127_3477_n2530), .A2(
        DP_OP_422J2_124_3477_n2400), .Y(DP_OP_424J2_126_3477_n2366) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1604 ( .A1(DP_OP_424J2_126_3477_n2397), .A2(
        DP_OP_423J2_125_3477_n2400), .Y(DP_OP_424J2_126_3477_n2365) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1603 ( .A1(DP_OP_425J2_127_3477_n2528), .A2(
        DP_OP_425J2_127_3477_n2400), .Y(DP_OP_424J2_126_3477_n2364) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1602 ( .A1(DP_OP_422J2_124_3477_n2659), .A2(
        DP_OP_422J2_124_3477_n2400), .Y(DP_OP_424J2_126_3477_n2363) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1601 ( .A1(DP_OP_422J2_124_3477_n2658), .A2(
        DP_OP_425J2_127_3477_n2400), .Y(DP_OP_424J2_126_3477_n2362) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1600 ( .A1(DP_OP_423J2_125_3477_n2305), .A2(
        DP_OP_422J2_124_3477_n2400), .Y(DP_OP_424J2_126_3477_n2361) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1599 ( .A1(DP_OP_423J2_125_3477_n2304), 
        .A2(DP_OP_423J2_125_3477_n2400), .Y(DP_OP_424J2_126_3477_n2360) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1579 ( .A1(DP_OP_422J2_124_3477_n2700), .A2(
        DP_OP_423J2_125_3477_n2359), .Y(DP_OP_424J2_126_3477_n2340) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1571 ( .A1(DP_OP_422J2_124_3477_n2700), .A2(
        DP_OP_424J2_126_3477_n2358), .Y(DP_OP_424J2_126_3477_n2332) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1563 ( .A1(DP_OP_422J2_124_3477_n2700), .A2(
        DP_OP_424J2_126_3477_n2357), .Y(DP_OP_424J2_126_3477_n2324) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1562 ( .A1(DP_OP_422J2_124_3477_n2707), .A2(
        DP_OP_422J2_124_3477_n2356), .Y(DP_OP_424J2_126_3477_n2323) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1561 ( .A1(DP_OP_424J2_126_3477_n2354), .A2(
        DP_OP_425J2_127_3477_n2356), .Y(DP_OP_424J2_126_3477_n2322) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1560 ( .A1(DP_OP_424J2_126_3477_n2353), .A2(
        DP_OP_425J2_127_3477_n2356), .Y(DP_OP_424J2_126_3477_n2321) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1559 ( .A1(DP_OP_422J2_124_3477_n2704), .A2(
        DP_OP_423J2_125_3477_n2356), .Y(DP_OP_424J2_126_3477_n2320) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1558 ( .A1(DP_OP_424J2_126_3477_n2351), .A2(
        DP_OP_423J2_125_3477_n2356), .Y(DP_OP_424J2_126_3477_n2319) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1557 ( .A1(DP_OP_422J2_124_3477_n2702), .A2(
        DP_OP_422J2_124_3477_n2356), .Y(DP_OP_424J2_126_3477_n2318) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1556 ( .A1(DP_OP_422J2_124_3477_n2701), .A2(
        DP_OP_423J2_125_3477_n2356), .Y(DP_OP_424J2_126_3477_n2317) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1555 ( .A1(DP_OP_422J2_124_3477_n2700), 
        .A2(DP_OP_422J2_124_3477_n2356), .Y(DP_OP_424J2_126_3477_n2316) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1535 ( .A1(DP_OP_424J2_126_3477_n2304), .A2(
        DP_OP_424J2_126_3477_n2315), .Y(DP_OP_424J2_126_3477_n2296) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1527 ( .A1(DP_OP_424J2_126_3477_n2304), .A2(
        DP_OP_424J2_126_3477_n2314), .Y(DP_OP_424J2_126_3477_n2288) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1519 ( .A1(DP_OP_424J2_126_3477_n2304), .A2(
        DP_OP_423J2_125_3477_n2313), .Y(DP_OP_424J2_126_3477_n2280) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1518 ( .A1(DP_OP_425J2_127_3477_n2619), .A2(
        DP_OP_422J2_124_3477_n2312), .Y(DP_OP_424J2_126_3477_n2279) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1517 ( .A1(DP_OP_424J2_126_3477_n2310), .A2(
        DP_OP_423J2_125_3477_n2312), .Y(DP_OP_424J2_126_3477_n2278) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1516 ( .A1(DP_OP_425J2_127_3477_n2617), .A2(
        DP_OP_423J2_125_3477_n2312), .Y(DP_OP_424J2_126_3477_n2277) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1515 ( .A1(DP_OP_424J2_126_3477_n2308), .A2(
        DP_OP_422J2_124_3477_n2312), .Y(DP_OP_424J2_126_3477_n2276) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1514 ( .A1(DP_OP_422J2_124_3477_n2747), .A2(
        DP_OP_425J2_127_3477_n2312), .Y(DP_OP_424J2_126_3477_n2275) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1513 ( .A1(DP_OP_422J2_124_3477_n2746), .A2(
        DP_OP_425J2_127_3477_n2312), .Y(DP_OP_424J2_126_3477_n2274) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1512 ( .A1(DP_OP_423J2_125_3477_n2217), .A2(
        DP_OP_422J2_124_3477_n2312), .Y(DP_OP_424J2_126_3477_n2273) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1511 ( .A1(DP_OP_424J2_126_3477_n2304), 
        .A2(DP_OP_425J2_127_3477_n2312), .Y(DP_OP_424J2_126_3477_n2272) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1492 ( .A1(DP_OP_424J2_126_3477_n2261), 
        .A2(DP_OP_424J2_126_3477_n2271), .Y(DP_OP_424J2_126_3477_n2253) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1491 ( .A1(DP_OP_424J2_126_3477_n2260), .A2(
        DP_OP_424J2_126_3477_n2271), .Y(DP_OP_424J2_126_3477_n2252) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1483 ( .A1(DP_OP_424J2_126_3477_n2260), .A2(
        DP_OP_424J2_126_3477_n2270), .Y(DP_OP_424J2_126_3477_n2244) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1475 ( .A1(DP_OP_424J2_126_3477_n2260), .A2(
        DP_OP_424J2_126_3477_n2269), .Y(DP_OP_424J2_126_3477_n2236) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1474 ( .A1(DP_OP_425J2_127_3477_n2663), .A2(
        DP_OP_422J2_124_3477_n2268), .Y(DP_OP_424J2_126_3477_n2235) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1473 ( .A1(DP_OP_425J2_127_3477_n2662), .A2(
        DP_OP_422J2_124_3477_n2268), .Y(DP_OP_424J2_126_3477_n2234) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1472 ( .A1(DP_OP_424J2_126_3477_n2265), .A2(
        DP_OP_423J2_125_3477_n2268), .Y(DP_OP_424J2_126_3477_n2233) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1471 ( .A1(DP_OP_424J2_126_3477_n2264), .A2(
        DP_OP_423J2_125_3477_n2268), .Y(DP_OP_424J2_126_3477_n2232) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1470 ( .A1(DP_OP_422J2_124_3477_n2791), .A2(
        DP_OP_425J2_127_3477_n2268), .Y(DP_OP_424J2_126_3477_n2231) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1469 ( .A1(DP_OP_425J2_127_3477_n2658), .A2(
        DP_OP_425J2_127_3477_n2268), .Y(DP_OP_424J2_126_3477_n2230) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1468 ( .A1(DP_OP_424J2_126_3477_n2261), .A2(
        DP_OP_422J2_124_3477_n2268), .Y(DP_OP_424J2_126_3477_n2229) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1467 ( .A1(DP_OP_424J2_126_3477_n2260), 
        .A2(DP_OP_425J2_127_3477_n2268), .Y(DP_OP_424J2_126_3477_n2228) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1447 ( .A1(DP_OP_423J2_125_3477_n2128), .A2(
        DP_OP_424J2_126_3477_n2227), .Y(DP_OP_424J2_126_3477_n2208) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1439 ( .A1(DP_OP_425J2_127_3477_n2700), .A2(
        DP_OP_424J2_126_3477_n2226), .Y(DP_OP_424J2_126_3477_n2200) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1432 ( .A1(DP_OP_424J2_126_3477_n2217), 
        .A2(DP_OP_424J2_126_3477_n2225), .Y(DP_OP_424J2_126_3477_n2193) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1431 ( .A1(DP_OP_425J2_127_3477_n2700), .A2(
        DP_OP_424J2_126_3477_n2225), .Y(DP_OP_424J2_126_3477_n2192) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1430 ( .A1(DP_OP_425J2_127_3477_n2707), .A2(
        DP_OP_422J2_124_3477_n2224), .Y(DP_OP_424J2_126_3477_n2191) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1429 ( .A1(DP_OP_423J2_125_3477_n2134), .A2(
        DP_OP_423J2_125_3477_n2224), .Y(DP_OP_424J2_126_3477_n2190) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1428 ( .A1(DP_OP_422J2_124_3477_n2837), .A2(
        DP_OP_425J2_127_3477_n2224), .Y(DP_OP_424J2_126_3477_n2189) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1427 ( .A1(DP_OP_424J2_126_3477_n2220), .A2(
        DP_OP_422J2_124_3477_n2224), .Y(DP_OP_424J2_126_3477_n2188) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1426 ( .A1(DP_OP_424J2_126_3477_n2219), .A2(
        DP_OP_422J2_124_3477_n2224), .Y(DP_OP_424J2_126_3477_n2187) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1425 ( .A1(DP_OP_424J2_126_3477_n2218), .A2(
        DP_OP_425J2_127_3477_n2224), .Y(DP_OP_424J2_126_3477_n2186) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1424 ( .A1(DP_OP_424J2_126_3477_n2217), .A2(
        DP_OP_425J2_127_3477_n2224), .Y(DP_OP_424J2_126_3477_n2185) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1423 ( .A1(DP_OP_425J2_127_3477_n2700), 
        .A2(DP_OP_423J2_125_3477_n2224), .Y(DP_OP_424J2_126_3477_n2184) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1403 ( .A1(DP_OP_424J2_126_3477_n2172), .A2(
        DP_OP_424J2_126_3477_n2183), .Y(DP_OP_424J2_126_3477_n2164) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1395 ( .A1(DP_OP_424J2_126_3477_n2172), .A2(
        DP_OP_424J2_126_3477_n2182), .Y(DP_OP_424J2_126_3477_n2156) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1387 ( .A1(DP_OP_424J2_126_3477_n2172), .A2(
        DP_OP_425J2_127_3477_n2181), .Y(DP_OP_424J2_126_3477_n2148) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1386 ( .A1(DP_OP_424J2_126_3477_n2179), .A2(
        DP_OP_422J2_124_3477_n2180), .Y(DP_OP_424J2_126_3477_n2147) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1385 ( .A1(DP_OP_424J2_126_3477_n2178), .A2(
        DP_OP_425J2_127_3477_n2180), .Y(DP_OP_424J2_126_3477_n2146) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1384 ( .A1(DP_OP_424J2_126_3477_n2177), .A2(
        DP_OP_423J2_125_3477_n2180), .Y(DP_OP_424J2_126_3477_n2145) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1383 ( .A1(DP_OP_423J2_125_3477_n2088), .A2(
        DP_OP_423J2_125_3477_n2180), .Y(DP_OP_424J2_126_3477_n2144) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1382 ( .A1(DP_OP_423J2_125_3477_n2087), .A2(
        DP_OP_422J2_124_3477_n2180), .Y(DP_OP_424J2_126_3477_n2143) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1381 ( .A1(DP_OP_422J2_124_3477_n2878), .A2(
        DP_OP_425J2_127_3477_n2180), .Y(DP_OP_424J2_126_3477_n2142) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1380 ( .A1(DP_OP_425J2_127_3477_n2745), .A2(
        DP_OP_425J2_127_3477_n2180), .Y(DP_OP_424J2_126_3477_n2141) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1379 ( .A1(DP_OP_424J2_126_3477_n2172), 
        .A2(DP_OP_422J2_124_3477_n2180), .Y(DP_OP_424J2_126_3477_n2140) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1359 ( .A1(DP_OP_424J2_126_3477_n2128), .A2(
        DP_OP_423J2_125_3477_n2139), .Y(DP_OP_424J2_126_3477_n2120) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1351 ( .A1(DP_OP_424J2_126_3477_n2128), .A2(
        DP_OP_422J2_124_3477_n2138), .Y(DP_OP_424J2_126_3477_n2112) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1344 ( .A1(DP_OP_422J2_124_3477_n2921), 
        .A2(DP_OP_424J2_126_3477_n2137), .Y(DP_OP_424J2_126_3477_n2105) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1343 ( .A1(DP_OP_424J2_126_3477_n2128), .A2(
        DP_OP_424J2_126_3477_n2137), .Y(DP_OP_424J2_126_3477_n2104) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1342 ( .A1(DP_OP_422J2_124_3477_n2927), .A2(
        DP_OP_422J2_124_3477_n2136), .Y(DP_OP_424J2_126_3477_n2103) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1341 ( .A1(DP_OP_422J2_124_3477_n2926), .A2(
        DP_OP_423J2_125_3477_n2136), .Y(DP_OP_424J2_126_3477_n2102) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1340 ( .A1(DP_OP_424J2_126_3477_n2133), .A2(
        DP_OP_425J2_127_3477_n2136), .Y(DP_OP_424J2_126_3477_n2101) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1339 ( .A1(DP_OP_422J2_124_3477_n2924), .A2(
        DP_OP_423J2_125_3477_n2136), .Y(DP_OP_424J2_126_3477_n2100) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1338 ( .A1(DP_OP_422J2_124_3477_n2923), .A2(
        DP_OP_425J2_127_3477_n2136), .Y(DP_OP_424J2_126_3477_n2099) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1337 ( .A1(DP_OP_422J2_124_3477_n2922), .A2(
        DP_OP_422J2_124_3477_n2136), .Y(DP_OP_424J2_126_3477_n2098) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1336 ( .A1(DP_OP_422J2_124_3477_n2921), .A2(
        DP_OP_422J2_124_3477_n2136), .Y(DP_OP_424J2_126_3477_n2097) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1335 ( .A1(DP_OP_424J2_126_3477_n2128), 
        .A2(DP_OP_423J2_125_3477_n2136), .Y(DP_OP_424J2_126_3477_n2096) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1322 ( .A1(DP_OP_423J2_125_3477_n2003), 
        .A2(DP_OP_424J2_126_3477_n2095), .Y(DP_OP_424J2_126_3477_n2083) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1321 ( .A1(DP_OP_424J2_126_3477_n2090), 
        .A2(DP_OP_424J2_126_3477_n2095), .Y(DP_OP_424J2_126_3477_n2082) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1320 ( .A1(DP_OP_422J2_124_3477_n2969), 
        .A2(DP_OP_424J2_126_3477_n2095), .Y(DP_OP_424J2_126_3477_n2081) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1319 ( .A1(DP_OP_424J2_126_3477_n2088), 
        .A2(DP_OP_424J2_126_3477_n2095), .Y(DP_OP_424J2_126_3477_n2080) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1318 ( .A1(DP_OP_424J2_126_3477_n2087), 
        .A2(DP_OP_424J2_126_3477_n2095), .Y(DP_OP_424J2_126_3477_n2079) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1317 ( .A1(DP_OP_423J2_125_3477_n1998), 
        .A2(DP_OP_424J2_126_3477_n2095), .Y(DP_OP_424J2_126_3477_n2078) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1316 ( .A1(DP_OP_423J2_125_3477_n1997), 
        .A2(DP_OP_424J2_126_3477_n2095), .Y(DP_OP_424J2_126_3477_n2077) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1315 ( .A1(DP_OP_424J2_126_3477_n2084), .A2(
        DP_OP_424J2_126_3477_n2095), .Y(DP_OP_424J2_126_3477_n2076) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1314 ( .A1(DP_OP_422J2_124_3477_n2971), 
        .A2(DP_OP_424J2_126_3477_n2094), .Y(DP_OP_424J2_126_3477_n2075) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1313 ( .A1(DP_OP_424J2_126_3477_n2090), 
        .A2(DP_OP_424J2_126_3477_n2094), .Y(DP_OP_424J2_126_3477_n2074) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1312 ( .A1(DP_OP_422J2_124_3477_n2969), 
        .A2(DP_OP_424J2_126_3477_n2094), .Y(DP_OP_424J2_126_3477_n2073) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1311 ( .A1(DP_OP_424J2_126_3477_n2088), 
        .A2(DP_OP_424J2_126_3477_n2094), .Y(DP_OP_424J2_126_3477_n2072) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1310 ( .A1(DP_OP_424J2_126_3477_n2087), 
        .A2(DP_OP_424J2_126_3477_n2094), .Y(DP_OP_424J2_126_3477_n2071) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1309 ( .A1(DP_OP_425J2_127_3477_n2834), 
        .A2(DP_OP_424J2_126_3477_n2094), .Y(DP_OP_424J2_126_3477_n2070) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1308 ( .A1(DP_OP_423J2_125_3477_n1997), 
        .A2(DP_OP_424J2_126_3477_n2094), .Y(DP_OP_424J2_126_3477_n2069) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1307 ( .A1(DP_OP_424J2_126_3477_n2084), .A2(
        DP_OP_424J2_126_3477_n2094), .Y(DP_OP_424J2_126_3477_n2068) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1299 ( .A1(DP_OP_424J2_126_3477_n2084), .A2(
        DP_OP_425J2_127_3477_n2093), .Y(DP_OP_424J2_126_3477_n2060) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1298 ( .A1(DP_OP_423J2_125_3477_n2003), .A2(
        DP_OP_425J2_127_3477_n2092), .Y(DP_OP_424J2_126_3477_n2059) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1297 ( .A1(DP_OP_424J2_126_3477_n2090), .A2(
        DP_OP_422J2_124_3477_n2092), .Y(DP_OP_424J2_126_3477_n2058) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1296 ( .A1(DP_OP_425J2_127_3477_n2837), .A2(
        DP_OP_423J2_125_3477_n2092), .Y(DP_OP_424J2_126_3477_n2057) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1295 ( .A1(DP_OP_424J2_126_3477_n2088), .A2(
        DP_OP_423J2_125_3477_n2092), .Y(DP_OP_424J2_126_3477_n2056) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1294 ( .A1(DP_OP_424J2_126_3477_n2087), .A2(
        DP_OP_422J2_124_3477_n2092), .Y(DP_OP_424J2_126_3477_n2055) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1293 ( .A1(DP_OP_425J2_127_3477_n2834), .A2(
        DP_OP_425J2_127_3477_n2092), .Y(DP_OP_424J2_126_3477_n2054) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1292 ( .A1(DP_OP_425J2_127_3477_n2833), .A2(
        DP_OP_422J2_124_3477_n2092), .Y(DP_OP_424J2_126_3477_n2053) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1291 ( .A1(DP_OP_424J2_126_3477_n2084), 
        .A2(DP_OP_425J2_127_3477_n2092), .Y(DP_OP_424J2_126_3477_n2052) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1275 ( .A1(DP_OP_424J2_126_3477_n2044), 
        .A2(DP_OP_424J2_126_3477_n2051), .Y(DP_OP_424J2_126_3477_n2036) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1263 ( .A1(DP_OP_423J2_125_3477_n1952), .A2(
        DP_OP_423J2_125_3477_n2050), .Y(DP_OP_424J2_126_3477_n2024) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1255 ( .A1(DP_OP_422J2_124_3477_n3006), .A2(
        DP_OP_424J2_126_3477_n2049), .Y(DP_OP_424J2_126_3477_n2016) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1254 ( .A1(DP_OP_424J2_126_3477_n2047), .A2(
        DP_OP_422J2_124_3477_n2048), .Y(DP_OP_424J2_126_3477_n2015) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1253 ( .A1(DP_OP_423J2_125_3477_n1958), .A2(
        DP_OP_422J2_124_3477_n2048), .Y(DP_OP_424J2_126_3477_n2014) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1252 ( .A1(DP_OP_423J2_125_3477_n1957), .A2(
        DP_OP_423J2_125_3477_n2048), .Y(DP_OP_424J2_126_3477_n2013) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1251 ( .A1(DP_OP_424J2_126_3477_n2044), .A2(
        DP_OP_423J2_125_3477_n2048), .Y(DP_OP_424J2_126_3477_n2012) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1250 ( .A1(DP_OP_422J2_124_3477_n3009), .A2(
        DP_OP_425J2_127_3477_n2048), .Y(DP_OP_424J2_126_3477_n2011) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1249 ( .A1(DP_OP_425J2_127_3477_n2878), .A2(
        DP_OP_425J2_127_3477_n2048), .Y(DP_OP_424J2_126_3477_n2010) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1248 ( .A1(DP_OP_422J2_124_3477_n3007), .A2(
        DP_OP_425J2_127_3477_n2048), .Y(DP_OP_424J2_126_3477_n2009) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1247 ( .A1(DP_OP_423J2_125_3477_n1952), 
        .A2(DP_OP_422J2_124_3477_n2048), .Y(DP_OP_424J2_126_3477_n2008) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1227 ( .A1(DP_OP_425J2_127_3477_n2920), .A2(
        DP_OP_423J2_125_3477_n2007), .Y(DP_OP_424J2_126_3477_n1988) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1219 ( .A1(DP_OP_425J2_127_3477_n2920), .A2(
        DP_OP_422J2_124_3477_n2006), .Y(DP_OP_424J2_126_3477_n1980) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1212 ( .A1(DP_OP_425J2_127_3477_n2921), 
        .A2(DP_OP_423J2_125_3477_n2005), .Y(DP_OP_424J2_126_3477_n1973) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1211 ( .A1(DP_OP_425J2_127_3477_n2920), .A2(
        DP_OP_425J2_127_3477_n2005), .Y(DP_OP_424J2_126_3477_n1972) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1210 ( .A1(DP_OP_425J2_127_3477_n2927), .A2(
        DP_OP_422J2_124_3477_n2004), .Y(DP_OP_424J2_126_3477_n1971) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1209 ( .A1(DP_OP_425J2_127_3477_n2926), .A2(
        DP_OP_425J2_127_3477_n2004), .Y(DP_OP_424J2_126_3477_n1970) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1208 ( .A1(DP_OP_424J2_126_3477_n2001), .A2(
        DP_OP_425J2_127_3477_n2004), .Y(DP_OP_424J2_126_3477_n1969) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1207 ( .A1(DP_OP_425J2_127_3477_n2924), .A2(
        DP_OP_422J2_124_3477_n2004), .Y(DP_OP_424J2_126_3477_n1968) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1206 ( .A1(DP_OP_425J2_127_3477_n2923), .A2(
        DP_OP_423J2_125_3477_n2004), .Y(DP_OP_424J2_126_3477_n1967) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1205 ( .A1(DP_OP_425J2_127_3477_n2922), .A2(
        DP_OP_423J2_125_3477_n2004), .Y(DP_OP_424J2_126_3477_n1966) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1204 ( .A1(DP_OP_425J2_127_3477_n2921), .A2(
        DP_OP_425J2_127_3477_n2004), .Y(DP_OP_424J2_126_3477_n1965) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1203 ( .A1(DP_OP_425J2_127_3477_n2920), 
        .A2(DP_OP_422J2_124_3477_n2004), .Y(DP_OP_424J2_126_3477_n1964) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1184 ( .A1(DP_OP_425J2_127_3477_n2965), 
        .A2(DP_OP_425J2_127_3477_n1963), .Y(DP_OP_424J2_126_3477_n1945) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1183 ( .A1(DP_OP_425J2_127_3477_n2964), .A2(
        DP_OP_422J2_124_3477_n1963), .Y(DP_OP_424J2_126_3477_n1944) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1175 ( .A1(DP_OP_425J2_127_3477_n2964), .A2(
        DP_OP_424J2_126_3477_n1962), .Y(DP_OP_424J2_126_3477_n1936) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1167 ( .A1(DP_OP_425J2_127_3477_n2964), .A2(
        DP_OP_424J2_126_3477_n1961), .Y(DP_OP_424J2_126_3477_n1928) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1166 ( .A1(DP_OP_425J2_127_3477_n2971), .A2(
        DP_OP_423J2_125_3477_n1960), .Y(DP_OP_424J2_126_3477_n1927) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1165 ( .A1(DP_OP_424J2_126_3477_n1958), .A2(
        DP_OP_425J2_127_3477_n1960), .Y(DP_OP_424J2_126_3477_n1926) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1164 ( .A1(DP_OP_424J2_126_3477_n1957), .A2(
        DP_OP_422J2_124_3477_n1960), .Y(DP_OP_424J2_126_3477_n1925) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1163 ( .A1(DP_OP_424J2_126_3477_n1956), .A2(
        DP_OP_423J2_125_3477_n1960), .Y(DP_OP_424J2_126_3477_n1924) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1162 ( .A1(DP_OP_425J2_127_3477_n2967), .A2(
        DP_OP_422J2_124_3477_n1960), .Y(DP_OP_424J2_126_3477_n1923) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1161 ( .A1(DP_OP_424J2_126_3477_n1954), .A2(
        DP_OP_425J2_127_3477_n1960), .Y(DP_OP_424J2_126_3477_n1922) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1160 ( .A1(DP_OP_425J2_127_3477_n2965), .A2(
        DP_OP_422J2_124_3477_n1960), .Y(DP_OP_424J2_126_3477_n1921) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1159 ( .A1(DP_OP_425J2_127_3477_n2964), 
        .A2(DP_OP_425J2_127_3477_n1960), .Y(DP_OP_424J2_126_3477_n1920) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1110 ( .A1(n513), .A2(n391), .Y(
        DP_OP_424J2_126_3477_n1873) );
  HADDX1_HVT DP_OP_424J2_126_3477_U1093 ( .A0(DP_OP_424J2_126_3477_n1886), 
        .B0(DP_OP_424J2_126_3477_n1995), .C1(DP_OP_424J2_126_3477_n1870), .SO(
        DP_OP_424J2_126_3477_n1871) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1092 ( .A(DP_OP_424J2_126_3477_n2039), .B(
        DP_OP_424J2_126_3477_n1951), .CI(DP_OP_424J2_126_3477_n2083), .CO(
        DP_OP_424J2_126_3477_n1868), .S(DP_OP_424J2_126_3477_n1869) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1091 ( .A(DP_OP_424J2_126_3477_n2171), .B(
        DP_OP_424J2_126_3477_n2127), .CI(DP_OP_424J2_126_3477_n2215), .CO(
        DP_OP_424J2_126_3477_n1866), .S(DP_OP_424J2_126_3477_n1867) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1090 ( .A(DP_OP_424J2_126_3477_n2303), .B(
        DP_OP_424J2_126_3477_n2259), .CI(DP_OP_424J2_126_3477_n2347), .CO(
        DP_OP_424J2_126_3477_n1864), .S(DP_OP_424J2_126_3477_n1865) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1089 ( .A(DP_OP_424J2_126_3477_n2435), .B(
        DP_OP_424J2_126_3477_n2391), .CI(DP_OP_424J2_126_3477_n2479), .CO(
        DP_OP_424J2_126_3477_n1862), .S(DP_OP_424J2_126_3477_n1863) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1088 ( .A(DP_OP_424J2_126_3477_n2567), .B(
        DP_OP_424J2_126_3477_n2523), .CI(DP_OP_424J2_126_3477_n2611), .CO(
        DP_OP_424J2_126_3477_n1860), .S(DP_OP_424J2_126_3477_n1861) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1087 ( .A(DP_OP_424J2_126_3477_n2699), .B(
        DP_OP_424J2_126_3477_n2655), .CI(DP_OP_424J2_126_3477_n2743), .CO(
        DP_OP_424J2_126_3477_n1858), .S(DP_OP_424J2_126_3477_n1859) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1086 ( .A(DP_OP_424J2_126_3477_n3005), .B(
        DP_OP_424J2_126_3477_n2787), .CI(DP_OP_424J2_126_3477_n2831), .CO(
        DP_OP_424J2_126_3477_n1856), .S(DP_OP_424J2_126_3477_n1857) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1085 ( .A(DP_OP_424J2_126_3477_n2963), .B(
        DP_OP_424J2_126_3477_n2875), .CI(DP_OP_424J2_126_3477_n2919), .CO(
        DP_OP_424J2_126_3477_n1854), .S(DP_OP_424J2_126_3477_n1855) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1084 ( .A(DP_OP_424J2_126_3477_n1871), .B(
        DP_OP_424J2_126_3477_n1857), .CI(DP_OP_424J2_126_3477_n1859), .CO(
        DP_OP_424J2_126_3477_n1852), .S(DP_OP_424J2_126_3477_n1853) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1083 ( .A(DP_OP_424J2_126_3477_n1861), .B(
        DP_OP_424J2_126_3477_n1855), .CI(DP_OP_424J2_126_3477_n1863), .CO(
        DP_OP_424J2_126_3477_n1850), .S(DP_OP_424J2_126_3477_n1851) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1082 ( .A(DP_OP_424J2_126_3477_n1869), .B(
        DP_OP_424J2_126_3477_n1865), .CI(DP_OP_424J2_126_3477_n1867), .CO(
        DP_OP_424J2_126_3477_n1848), .S(DP_OP_424J2_126_3477_n1849) );
  HADDX1_HVT DP_OP_424J2_126_3477_U1081 ( .A0(DP_OP_424J2_126_3477_n1885), 
        .B0(DP_OP_424J2_126_3477_n1950), .C1(DP_OP_424J2_126_3477_n1846), .SO(
        DP_OP_424J2_126_3477_n1847) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1080 ( .A(DP_OP_424J2_126_3477_n1987), .B(
        DP_OP_424J2_126_3477_n1943), .CI(DP_OP_424J2_126_3477_n1994), .CO(
        DP_OP_424J2_126_3477_n1844), .S(DP_OP_424J2_126_3477_n1845) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1079 ( .A(DP_OP_424J2_126_3477_n2038), .B(
        DP_OP_424J2_126_3477_n2031), .CI(DP_OP_424J2_126_3477_n2075), .CO(
        DP_OP_424J2_126_3477_n1842), .S(DP_OP_424J2_126_3477_n1843) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1078 ( .A(DP_OP_424J2_126_3477_n2119), .B(
        DP_OP_424J2_126_3477_n2082), .CI(DP_OP_424J2_126_3477_n2126), .CO(
        DP_OP_424J2_126_3477_n1840), .S(DP_OP_424J2_126_3477_n1841) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1077 ( .A(DP_OP_424J2_126_3477_n2170), .B(
        DP_OP_424J2_126_3477_n2163), .CI(DP_OP_424J2_126_3477_n2207), .CO(
        DP_OP_424J2_126_3477_n1838), .S(DP_OP_424J2_126_3477_n1839) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1076 ( .A(DP_OP_424J2_126_3477_n2251), .B(
        DP_OP_424J2_126_3477_n2214), .CI(DP_OP_424J2_126_3477_n2258), .CO(
        DP_OP_424J2_126_3477_n1836), .S(DP_OP_424J2_126_3477_n1837) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1075 ( .A(DP_OP_424J2_126_3477_n2302), .B(
        DP_OP_424J2_126_3477_n2295), .CI(DP_OP_424J2_126_3477_n2339), .CO(
        DP_OP_424J2_126_3477_n1834), .S(DP_OP_424J2_126_3477_n1835) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1074 ( .A(DP_OP_424J2_126_3477_n2383), .B(
        DP_OP_424J2_126_3477_n2346), .CI(DP_OP_424J2_126_3477_n2390), .CO(
        DP_OP_424J2_126_3477_n1832), .S(DP_OP_424J2_126_3477_n1833) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1073 ( .A(DP_OP_424J2_126_3477_n2434), .B(
        DP_OP_424J2_126_3477_n2427), .CI(DP_OP_424J2_126_3477_n2471), .CO(
        DP_OP_424J2_126_3477_n1830), .S(DP_OP_424J2_126_3477_n1831) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1072 ( .A(DP_OP_424J2_126_3477_n2515), .B(
        DP_OP_424J2_126_3477_n2478), .CI(DP_OP_424J2_126_3477_n2522), .CO(
        DP_OP_424J2_126_3477_n1828), .S(DP_OP_424J2_126_3477_n1829) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1071 ( .A(DP_OP_424J2_126_3477_n3004), .B(
        DP_OP_424J2_126_3477_n2559), .CI(DP_OP_424J2_126_3477_n2997), .CO(
        DP_OP_424J2_126_3477_n1826), .S(DP_OP_424J2_126_3477_n1827) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1070 ( .A(DP_OP_424J2_126_3477_n2742), .B(
        DP_OP_424J2_126_3477_n2566), .CI(DP_OP_424J2_126_3477_n2603), .CO(
        DP_OP_424J2_126_3477_n1824), .S(DP_OP_424J2_126_3477_n1825) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1069 ( .A(DP_OP_424J2_126_3477_n2779), .B(
        DP_OP_424J2_126_3477_n2962), .CI(DP_OP_424J2_126_3477_n2955), .CO(
        DP_OP_424J2_126_3477_n1822), .S(DP_OP_424J2_126_3477_n1823) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1068 ( .A(DP_OP_424J2_126_3477_n2698), .B(
        DP_OP_424J2_126_3477_n2918), .CI(DP_OP_424J2_126_3477_n2911), .CO(
        DP_OP_424J2_126_3477_n1820), .S(DP_OP_424J2_126_3477_n1821) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1067 ( .A(DP_OP_424J2_126_3477_n2691), .B(
        DP_OP_424J2_126_3477_n2874), .CI(DP_OP_424J2_126_3477_n2610), .CO(
        DP_OP_424J2_126_3477_n1818), .S(DP_OP_424J2_126_3477_n1819) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1066 ( .A(DP_OP_424J2_126_3477_n2867), .B(
        DP_OP_424J2_126_3477_n2647), .CI(DP_OP_424J2_126_3477_n2654), .CO(
        DP_OP_424J2_126_3477_n1816), .S(DP_OP_424J2_126_3477_n1817) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1065 ( .A(DP_OP_424J2_126_3477_n2823), .B(
        DP_OP_424J2_126_3477_n2735), .CI(DP_OP_424J2_126_3477_n2786), .CO(
        DP_OP_424J2_126_3477_n1814), .S(DP_OP_424J2_126_3477_n1815) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1064 ( .A(DP_OP_424J2_126_3477_n2830), .B(
        DP_OP_424J2_126_3477_n1870), .CI(DP_OP_424J2_126_3477_n1847), .CO(
        DP_OP_424J2_126_3477_n1812), .S(DP_OP_424J2_126_3477_n1813) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1063 ( .A(DP_OP_424J2_126_3477_n1854), .B(
        DP_OP_424J2_126_3477_n1868), .CI(DP_OP_424J2_126_3477_n1866), .CO(
        DP_OP_424J2_126_3477_n1810), .S(DP_OP_424J2_126_3477_n1811) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1062 ( .A(DP_OP_424J2_126_3477_n1860), .B(
        DP_OP_424J2_126_3477_n1856), .CI(DP_OP_424J2_126_3477_n1864), .CO(
        DP_OP_424J2_126_3477_n1808), .S(DP_OP_424J2_126_3477_n1809) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1061 ( .A(DP_OP_424J2_126_3477_n1862), .B(
        DP_OP_424J2_126_3477_n1858), .CI(DP_OP_424J2_126_3477_n1815), .CO(
        DP_OP_424J2_126_3477_n1806), .S(DP_OP_424J2_126_3477_n1807) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1060 ( .A(DP_OP_424J2_126_3477_n1837), .B(
        DP_OP_424J2_126_3477_n1823), .CI(DP_OP_424J2_126_3477_n1821), .CO(
        DP_OP_424J2_126_3477_n1804), .S(DP_OP_424J2_126_3477_n1805) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1059 ( .A(DP_OP_424J2_126_3477_n1841), .B(
        DP_OP_424J2_126_3477_n1825), .CI(DP_OP_424J2_126_3477_n1829), .CO(
        DP_OP_424J2_126_3477_n1802), .S(DP_OP_424J2_126_3477_n1803) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1058 ( .A(DP_OP_424J2_126_3477_n1843), .B(
        DP_OP_424J2_126_3477_n1831), .CI(DP_OP_424J2_126_3477_n1827), .CO(
        DP_OP_424J2_126_3477_n1800), .S(DP_OP_424J2_126_3477_n1801) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1057 ( .A(DP_OP_424J2_126_3477_n1845), .B(
        DP_OP_424J2_126_3477_n1835), .CI(DP_OP_424J2_126_3477_n1819), .CO(
        DP_OP_424J2_126_3477_n1798), .S(DP_OP_424J2_126_3477_n1799) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1056 ( .A(DP_OP_424J2_126_3477_n1839), .B(
        DP_OP_424J2_126_3477_n1833), .CI(DP_OP_424J2_126_3477_n1817), .CO(
        DP_OP_424J2_126_3477_n1796), .S(DP_OP_424J2_126_3477_n1797) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1055 ( .A(DP_OP_424J2_126_3477_n1813), .B(
        DP_OP_424J2_126_3477_n1852), .CI(DP_OP_424J2_126_3477_n1850), .CO(
        DP_OP_424J2_126_3477_n1794), .S(DP_OP_424J2_126_3477_n1795) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1054 ( .A(DP_OP_424J2_126_3477_n1848), .B(
        DP_OP_424J2_126_3477_n1809), .CI(DP_OP_424J2_126_3477_n1811), .CO(
        DP_OP_424J2_126_3477_n1792), .S(DP_OP_424J2_126_3477_n1793) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1053 ( .A(DP_OP_424J2_126_3477_n1807), .B(
        DP_OP_424J2_126_3477_n1799), .CI(DP_OP_424J2_126_3477_n1801), .CO(
        DP_OP_424J2_126_3477_n1790), .S(DP_OP_424J2_126_3477_n1791) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1052 ( .A(DP_OP_424J2_126_3477_n1805), .B(
        DP_OP_424J2_126_3477_n1797), .CI(DP_OP_424J2_126_3477_n1803), .CO(
        DP_OP_424J2_126_3477_n1788), .S(DP_OP_424J2_126_3477_n1789) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1051 ( .A(DP_OP_424J2_126_3477_n1795), .B(
        DP_OP_424J2_126_3477_n1793), .CI(DP_OP_424J2_126_3477_n1791), .CO(
        DP_OP_424J2_126_3477_n1786), .S(DP_OP_424J2_126_3477_n1787) );
  HADDX1_HVT DP_OP_424J2_126_3477_U1050 ( .A0(DP_OP_424J2_126_3477_n1884), 
        .B0(DP_OP_424J2_126_3477_n1949), .C1(DP_OP_424J2_126_3477_n1784), .SO(
        DP_OP_424J2_126_3477_n1785) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1049 ( .A(DP_OP_424J2_126_3477_n1979), .B(
        DP_OP_424J2_126_3477_n1942), .CI(DP_OP_424J2_126_3477_n1935), .CO(
        DP_OP_424J2_126_3477_n1782), .S(DP_OP_424J2_126_3477_n1783) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1048 ( .A(DP_OP_424J2_126_3477_n1993), .B(
        DP_OP_424J2_126_3477_n1986), .CI(DP_OP_424J2_126_3477_n2023), .CO(
        DP_OP_424J2_126_3477_n1780), .S(DP_OP_424J2_126_3477_n1781) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1047 ( .A(DP_OP_424J2_126_3477_n2037), .B(
        DP_OP_424J2_126_3477_n2030), .CI(DP_OP_424J2_126_3477_n2067), .CO(
        DP_OP_424J2_126_3477_n1778), .S(DP_OP_424J2_126_3477_n1779) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1046 ( .A(DP_OP_424J2_126_3477_n2081), .B(
        DP_OP_424J2_126_3477_n2074), .CI(DP_OP_424J2_126_3477_n2111), .CO(
        DP_OP_424J2_126_3477_n1776), .S(DP_OP_424J2_126_3477_n1777) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1045 ( .A(DP_OP_424J2_126_3477_n2125), .B(
        DP_OP_424J2_126_3477_n2118), .CI(DP_OP_424J2_126_3477_n2155), .CO(
        DP_OP_424J2_126_3477_n1774), .S(DP_OP_424J2_126_3477_n1775) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1044 ( .A(DP_OP_424J2_126_3477_n2169), .B(
        DP_OP_424J2_126_3477_n2162), .CI(DP_OP_424J2_126_3477_n2199), .CO(
        DP_OP_424J2_126_3477_n1772), .S(DP_OP_424J2_126_3477_n1773) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1043 ( .A(DP_OP_424J2_126_3477_n2213), .B(
        DP_OP_424J2_126_3477_n2206), .CI(DP_OP_424J2_126_3477_n2243), .CO(
        DP_OP_424J2_126_3477_n1770), .S(DP_OP_424J2_126_3477_n1771) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1042 ( .A(DP_OP_424J2_126_3477_n2257), .B(
        DP_OP_424J2_126_3477_n2250), .CI(DP_OP_424J2_126_3477_n2287), .CO(
        DP_OP_424J2_126_3477_n1768), .S(DP_OP_424J2_126_3477_n1769) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1041 ( .A(DP_OP_424J2_126_3477_n2301), .B(
        DP_OP_424J2_126_3477_n2294), .CI(DP_OP_424J2_126_3477_n2331), .CO(
        DP_OP_424J2_126_3477_n1766), .S(DP_OP_424J2_126_3477_n1767) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1040 ( .A(DP_OP_424J2_126_3477_n2345), .B(
        DP_OP_424J2_126_3477_n2338), .CI(DP_OP_424J2_126_3477_n2375), .CO(
        DP_OP_424J2_126_3477_n1764), .S(DP_OP_424J2_126_3477_n1765) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1039 ( .A(DP_OP_424J2_126_3477_n2389), .B(
        DP_OP_424J2_126_3477_n2382), .CI(DP_OP_424J2_126_3477_n2419), .CO(
        DP_OP_424J2_126_3477_n1762), .S(DP_OP_424J2_126_3477_n1763) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1038 ( .A(DP_OP_424J2_126_3477_n2690), .B(
        DP_OP_424J2_126_3477_n3003), .CI(DP_OP_424J2_126_3477_n2996), .CO(
        DP_OP_424J2_126_3477_n1760), .S(DP_OP_424J2_126_3477_n1761) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1037 ( .A(DP_OP_424J2_126_3477_n2653), .B(
        DP_OP_424J2_126_3477_n2426), .CI(DP_OP_424J2_126_3477_n2989), .CO(
        DP_OP_424J2_126_3477_n1758), .S(DP_OP_424J2_126_3477_n1759) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1036 ( .A(DP_OP_424J2_126_3477_n2646), .B(
        DP_OP_424J2_126_3477_n2961), .CI(DP_OP_424J2_126_3477_n2433), .CO(
        DP_OP_424J2_126_3477_n1756), .S(DP_OP_424J2_126_3477_n1757) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1035 ( .A(DP_OP_424J2_126_3477_n2683), .B(
        DP_OP_424J2_126_3477_n2463), .CI(DP_OP_424J2_126_3477_n2470), .CO(
        DP_OP_424J2_126_3477_n1754), .S(DP_OP_424J2_126_3477_n1755) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1034 ( .A(DP_OP_424J2_126_3477_n2697), .B(
        DP_OP_424J2_126_3477_n2477), .CI(DP_OP_424J2_126_3477_n2954), .CO(
        DP_OP_424J2_126_3477_n1752), .S(DP_OP_424J2_126_3477_n1753) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1033 ( .A(DP_OP_424J2_126_3477_n2727), .B(
        DP_OP_424J2_126_3477_n2507), .CI(DP_OP_424J2_126_3477_n2947), .CO(
        DP_OP_424J2_126_3477_n1750), .S(DP_OP_424J2_126_3477_n1751) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1032 ( .A(DP_OP_424J2_126_3477_n2639), .B(
        DP_OP_424J2_126_3477_n2514), .CI(DP_OP_424J2_126_3477_n2917), .CO(
        DP_OP_424J2_126_3477_n1748), .S(DP_OP_424J2_126_3477_n1749) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1031 ( .A(DP_OP_424J2_126_3477_n2609), .B(
        DP_OP_424J2_126_3477_n2521), .CI(DP_OP_424J2_126_3477_n2910), .CO(
        DP_OP_424J2_126_3477_n1746), .S(DP_OP_424J2_126_3477_n1747) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1030 ( .A(DP_OP_424J2_126_3477_n2903), .B(
        DP_OP_424J2_126_3477_n2551), .CI(DP_OP_424J2_126_3477_n2558), .CO(
        DP_OP_424J2_126_3477_n1744), .S(DP_OP_424J2_126_3477_n1745) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1029 ( .A(DP_OP_424J2_126_3477_n2873), .B(
        DP_OP_424J2_126_3477_n2565), .CI(DP_OP_424J2_126_3477_n2595), .CO(
        DP_OP_424J2_126_3477_n1742), .S(DP_OP_424J2_126_3477_n1743) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1028 ( .A(DP_OP_424J2_126_3477_n2866), .B(
        DP_OP_424J2_126_3477_n2602), .CI(DP_OP_424J2_126_3477_n2734), .CO(
        DP_OP_424J2_126_3477_n1740), .S(DP_OP_424J2_126_3477_n1741) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1027 ( .A(DP_OP_424J2_126_3477_n2859), .B(
        DP_OP_424J2_126_3477_n2741), .CI(DP_OP_424J2_126_3477_n2771), .CO(
        DP_OP_424J2_126_3477_n1738), .S(DP_OP_424J2_126_3477_n1739) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1026 ( .A(DP_OP_424J2_126_3477_n2829), .B(
        DP_OP_424J2_126_3477_n2778), .CI(DP_OP_424J2_126_3477_n2785), .CO(
        DP_OP_424J2_126_3477_n1736), .S(DP_OP_424J2_126_3477_n1737) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1025 ( .A(DP_OP_424J2_126_3477_n2822), .B(
        DP_OP_424J2_126_3477_n2815), .CI(DP_OP_424J2_126_3477_n1846), .CO(
        DP_OP_424J2_126_3477_n1734), .S(DP_OP_424J2_126_3477_n1735) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1024 ( .A(DP_OP_424J2_126_3477_n1785), .B(
        DP_OP_424J2_126_3477_n1814), .CI(DP_OP_424J2_126_3477_n1816), .CO(
        DP_OP_424J2_126_3477_n1732), .S(DP_OP_424J2_126_3477_n1733) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1023 ( .A(DP_OP_424J2_126_3477_n1832), .B(
        DP_OP_424J2_126_3477_n1844), .CI(DP_OP_424J2_126_3477_n1818), .CO(
        DP_OP_424J2_126_3477_n1730), .S(DP_OP_424J2_126_3477_n1731) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1022 ( .A(DP_OP_424J2_126_3477_n1830), .B(
        DP_OP_424J2_126_3477_n1842), .CI(DP_OP_424J2_126_3477_n1820), .CO(
        DP_OP_424J2_126_3477_n1728), .S(DP_OP_424J2_126_3477_n1729) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1021 ( .A(DP_OP_424J2_126_3477_n1826), .B(
        DP_OP_424J2_126_3477_n1840), .CI(DP_OP_424J2_126_3477_n1822), .CO(
        DP_OP_424J2_126_3477_n1726), .S(DP_OP_424J2_126_3477_n1727) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1020 ( .A(DP_OP_424J2_126_3477_n1838), .B(
        DP_OP_424J2_126_3477_n1836), .CI(DP_OP_424J2_126_3477_n1834), .CO(
        DP_OP_424J2_126_3477_n1724), .S(DP_OP_424J2_126_3477_n1725) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1019 ( .A(DP_OP_424J2_126_3477_n1828), .B(
        DP_OP_424J2_126_3477_n1824), .CI(DP_OP_424J2_126_3477_n1757), .CO(
        DP_OP_424J2_126_3477_n1722), .S(DP_OP_424J2_126_3477_n1723) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1018 ( .A(DP_OP_424J2_126_3477_n1751), .B(
        DP_OP_424J2_126_3477_n1765), .CI(DP_OP_424J2_126_3477_n1769), .CO(
        DP_OP_424J2_126_3477_n1720), .S(DP_OP_424J2_126_3477_n1721) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1017 ( .A(DP_OP_424J2_126_3477_n1747), .B(
        DP_OP_424J2_126_3477_n1775), .CI(DP_OP_424J2_126_3477_n1777), .CO(
        DP_OP_424J2_126_3477_n1718), .S(DP_OP_424J2_126_3477_n1719) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1016 ( .A(DP_OP_424J2_126_3477_n1745), .B(
        DP_OP_424J2_126_3477_n1767), .CI(DP_OP_424J2_126_3477_n1781), .CO(
        DP_OP_424J2_126_3477_n1716), .S(DP_OP_424J2_126_3477_n1717) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1015 ( .A(DP_OP_424J2_126_3477_n1743), .B(
        DP_OP_424J2_126_3477_n1761), .CI(DP_OP_424J2_126_3477_n1779), .CO(
        DP_OP_424J2_126_3477_n1714), .S(DP_OP_424J2_126_3477_n1715) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1014 ( .A(DP_OP_424J2_126_3477_n1741), .B(
        DP_OP_424J2_126_3477_n1771), .CI(DP_OP_424J2_126_3477_n1759), .CO(
        DP_OP_424J2_126_3477_n1712), .S(DP_OP_424J2_126_3477_n1713) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1013 ( .A(DP_OP_424J2_126_3477_n1739), .B(
        DP_OP_424J2_126_3477_n1773), .CI(DP_OP_424J2_126_3477_n1783), .CO(
        DP_OP_424J2_126_3477_n1710), .S(DP_OP_424J2_126_3477_n1711) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1012 ( .A(DP_OP_424J2_126_3477_n1737), .B(
        DP_OP_424J2_126_3477_n1763), .CI(DP_OP_424J2_126_3477_n1749), .CO(
        DP_OP_424J2_126_3477_n1708), .S(DP_OP_424J2_126_3477_n1709) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1011 ( .A(DP_OP_424J2_126_3477_n1755), .B(
        DP_OP_424J2_126_3477_n1753), .CI(DP_OP_424J2_126_3477_n1812), .CO(
        DP_OP_424J2_126_3477_n1706), .S(DP_OP_424J2_126_3477_n1707) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1010 ( .A(DP_OP_424J2_126_3477_n1735), .B(
        DP_OP_424J2_126_3477_n1810), .CI(DP_OP_424J2_126_3477_n1808), .CO(
        DP_OP_424J2_126_3477_n1704), .S(DP_OP_424J2_126_3477_n1705) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1009 ( .A(DP_OP_424J2_126_3477_n1806), .B(
        DP_OP_424J2_126_3477_n1733), .CI(DP_OP_424J2_126_3477_n1800), .CO(
        DP_OP_424J2_126_3477_n1702), .S(DP_OP_424J2_126_3477_n1703) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1008 ( .A(DP_OP_424J2_126_3477_n1804), .B(
        DP_OP_424J2_126_3477_n1725), .CI(DP_OP_424J2_126_3477_n1731), .CO(
        DP_OP_424J2_126_3477_n1700), .S(DP_OP_424J2_126_3477_n1701) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1007 ( .A(DP_OP_424J2_126_3477_n1802), .B(
        DP_OP_424J2_126_3477_n1729), .CI(DP_OP_424J2_126_3477_n1727), .CO(
        DP_OP_424J2_126_3477_n1698), .S(DP_OP_424J2_126_3477_n1699) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1006 ( .A(DP_OP_424J2_126_3477_n1798), .B(
        DP_OP_424J2_126_3477_n1796), .CI(DP_OP_424J2_126_3477_n1723), .CO(
        DP_OP_424J2_126_3477_n1696), .S(DP_OP_424J2_126_3477_n1697) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1005 ( .A(DP_OP_424J2_126_3477_n1721), .B(
        DP_OP_424J2_126_3477_n1709), .CI(DP_OP_424J2_126_3477_n1707), .CO(
        DP_OP_424J2_126_3477_n1694), .S(DP_OP_424J2_126_3477_n1695) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1004 ( .A(DP_OP_424J2_126_3477_n1711), .B(
        DP_OP_424J2_126_3477_n1719), .CI(DP_OP_424J2_126_3477_n1717), .CO(
        DP_OP_424J2_126_3477_n1692), .S(DP_OP_424J2_126_3477_n1693) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1003 ( .A(DP_OP_424J2_126_3477_n1713), .B(
        DP_OP_424J2_126_3477_n1715), .CI(DP_OP_424J2_126_3477_n1794), .CO(
        DP_OP_424J2_126_3477_n1690), .S(DP_OP_424J2_126_3477_n1691) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1002 ( .A(DP_OP_424J2_126_3477_n1705), .B(
        DP_OP_424J2_126_3477_n1792), .CI(DP_OP_424J2_126_3477_n1703), .CO(
        DP_OP_424J2_126_3477_n1688), .S(DP_OP_424J2_126_3477_n1689) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1001 ( .A(DP_OP_424J2_126_3477_n1790), .B(
        DP_OP_424J2_126_3477_n1788), .CI(DP_OP_424J2_126_3477_n1699), .CO(
        DP_OP_424J2_126_3477_n1686), .S(DP_OP_424J2_126_3477_n1687) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1000 ( .A(DP_OP_424J2_126_3477_n1701), .B(
        DP_OP_424J2_126_3477_n1697), .CI(DP_OP_424J2_126_3477_n1695), .CO(
        DP_OP_424J2_126_3477_n1684), .S(DP_OP_424J2_126_3477_n1685) );
  FADDX1_HVT DP_OP_424J2_126_3477_U999 ( .A(DP_OP_424J2_126_3477_n1693), .B(
        DP_OP_424J2_126_3477_n1691), .CI(DP_OP_424J2_126_3477_n1689), .CO(
        DP_OP_424J2_126_3477_n1682), .S(DP_OP_424J2_126_3477_n1683) );
  FADDX1_HVT DP_OP_424J2_126_3477_U998 ( .A(DP_OP_424J2_126_3477_n1786), .B(
        DP_OP_424J2_126_3477_n1687), .CI(DP_OP_424J2_126_3477_n1685), .CO(
        DP_OP_424J2_126_3477_n1680), .S(DP_OP_424J2_126_3477_n1681) );
  FADDX1_HVT DP_OP_424J2_126_3477_U996 ( .A(DP_OP_424J2_126_3477_n2455), .B(
        DP_OP_424J2_126_3477_n1927), .CI(DP_OP_424J2_126_3477_n1883), .CO(
        DP_OP_424J2_126_3477_n1676), .S(DP_OP_424J2_126_3477_n1677) );
  FADDX1_HVT DP_OP_424J2_126_3477_U995 ( .A(DP_OP_424J2_126_3477_n2147), .B(
        DP_OP_424J2_126_3477_n2587), .CI(DP_OP_424J2_126_3477_n2367), .CO(
        DP_OP_424J2_126_3477_n1674), .S(DP_OP_424J2_126_3477_n1675) );
  FADDX1_HVT DP_OP_424J2_126_3477_U994 ( .A(DP_OP_424J2_126_3477_n2895), .B(
        DP_OP_424J2_126_3477_n2103), .CI(DP_OP_424J2_126_3477_n2323), .CO(
        DP_OP_424J2_126_3477_n1672), .S(DP_OP_424J2_126_3477_n1673) );
  FADDX1_HVT DP_OP_424J2_126_3477_U993 ( .A(DP_OP_424J2_126_3477_n2499), .B(
        DP_OP_424J2_126_3477_n2807), .CI(DP_OP_424J2_126_3477_n2411), .CO(
        DP_OP_424J2_126_3477_n1670), .S(DP_OP_424J2_126_3477_n1671) );
  FADDX1_HVT DP_OP_424J2_126_3477_U992 ( .A(DP_OP_424J2_126_3477_n2235), .B(
        DP_OP_424J2_126_3477_n2279), .CI(DP_OP_424J2_126_3477_n2059), .CO(
        DP_OP_424J2_126_3477_n1668), .S(DP_OP_424J2_126_3477_n1669) );
  FADDX1_HVT DP_OP_424J2_126_3477_U991 ( .A(DP_OP_424J2_126_3477_n2763), .B(
        DP_OP_424J2_126_3477_n2631), .CI(DP_OP_424J2_126_3477_n2675), .CO(
        DP_OP_424J2_126_3477_n1666), .S(DP_OP_424J2_126_3477_n1667) );
  FADDX1_HVT DP_OP_424J2_126_3477_U990 ( .A(DP_OP_424J2_126_3477_n2015), .B(
        DP_OP_424J2_126_3477_n2851), .CI(DP_OP_424J2_126_3477_n2719), .CO(
        DP_OP_424J2_126_3477_n1664), .S(DP_OP_424J2_126_3477_n1665) );
  FADDX1_HVT DP_OP_424J2_126_3477_U989 ( .A(DP_OP_424J2_126_3477_n2543), .B(
        DP_OP_424J2_126_3477_n2939), .CI(DP_OP_424J2_126_3477_n2191), .CO(
        DP_OP_424J2_126_3477_n1662), .S(DP_OP_424J2_126_3477_n1663) );
  FADDX1_HVT DP_OP_424J2_126_3477_U988 ( .A(DP_OP_424J2_126_3477_n1971), .B(
        DP_OP_424J2_126_3477_n1679), .CI(DP_OP_424J2_126_3477_n1948), .CO(
        DP_OP_424J2_126_3477_n1660), .S(DP_OP_424J2_126_3477_n1661) );
  FADDX1_HVT DP_OP_424J2_126_3477_U987 ( .A(DP_OP_424J2_126_3477_n1978), .B(
        DP_OP_424J2_126_3477_n1941), .CI(DP_OP_424J2_126_3477_n1934), .CO(
        DP_OP_424J2_126_3477_n1658), .S(DP_OP_424J2_126_3477_n1659) );
  FADDX1_HVT DP_OP_424J2_126_3477_U986 ( .A(DP_OP_424J2_126_3477_n1992), .B(
        DP_OP_424J2_126_3477_n1985), .CI(DP_OP_424J2_126_3477_n2022), .CO(
        DP_OP_424J2_126_3477_n1656), .S(DP_OP_424J2_126_3477_n1657) );
  FADDX1_HVT DP_OP_424J2_126_3477_U985 ( .A(DP_OP_424J2_126_3477_n2036), .B(
        DP_OP_424J2_126_3477_n2029), .CI(DP_OP_424J2_126_3477_n2066), .CO(
        DP_OP_424J2_126_3477_n1654), .S(DP_OP_424J2_126_3477_n1655) );
  FADDX1_HVT DP_OP_424J2_126_3477_U984 ( .A(DP_OP_424J2_126_3477_n3002), .B(
        DP_OP_424J2_126_3477_n2073), .CI(DP_OP_424J2_126_3477_n2080), .CO(
        DP_OP_424J2_126_3477_n1652), .S(DP_OP_424J2_126_3477_n1653) );
  FADDX1_HVT DP_OP_424J2_126_3477_U983 ( .A(DP_OP_424J2_126_3477_n2513), .B(
        DP_OP_424J2_126_3477_n2995), .CI(DP_OP_424J2_126_3477_n2988), .CO(
        DP_OP_424J2_126_3477_n1650), .S(DP_OP_424J2_126_3477_n1651) );
  FADDX1_HVT DP_OP_424J2_126_3477_U982 ( .A(DP_OP_424J2_126_3477_n2476), .B(
        DP_OP_424J2_126_3477_n2110), .CI(DP_OP_424J2_126_3477_n2960), .CO(
        DP_OP_424J2_126_3477_n1648), .S(DP_OP_424J2_126_3477_n1649) );
  FADDX1_HVT DP_OP_424J2_126_3477_U981 ( .A(DP_OP_424J2_126_3477_n2506), .B(
        DP_OP_424J2_126_3477_n2117), .CI(DP_OP_424J2_126_3477_n2953), .CO(
        DP_OP_424J2_126_3477_n1646), .S(DP_OP_424J2_126_3477_n1647) );
  FADDX1_HVT DP_OP_424J2_126_3477_U980 ( .A(DP_OP_424J2_126_3477_n2946), .B(
        DP_OP_424J2_126_3477_n2124), .CI(DP_OP_424J2_126_3477_n2154), .CO(
        DP_OP_424J2_126_3477_n1644), .S(DP_OP_424J2_126_3477_n1645) );
  FADDX1_HVT DP_OP_424J2_126_3477_U979 ( .A(DP_OP_424J2_126_3477_n2469), .B(
        DP_OP_424J2_126_3477_n2161), .CI(DP_OP_424J2_126_3477_n2168), .CO(
        DP_OP_424J2_126_3477_n1642), .S(DP_OP_424J2_126_3477_n1643) );
  FADDX1_HVT DP_OP_424J2_126_3477_U978 ( .A(DP_OP_424J2_126_3477_n2550), .B(
        DP_OP_424J2_126_3477_n2198), .CI(DP_OP_424J2_126_3477_n2205), .CO(
        DP_OP_424J2_126_3477_n1640), .S(DP_OP_424J2_126_3477_n1641) );
  FADDX1_HVT DP_OP_424J2_126_3477_U977 ( .A(DP_OP_424J2_126_3477_n2557), .B(
        DP_OP_424J2_126_3477_n2212), .CI(DP_OP_424J2_126_3477_n2242), .CO(
        DP_OP_424J2_126_3477_n1638), .S(DP_OP_424J2_126_3477_n1639) );
  FADDX1_HVT DP_OP_424J2_126_3477_U976 ( .A(DP_OP_424J2_126_3477_n2564), .B(
        DP_OP_424J2_126_3477_n2916), .CI(DP_OP_424J2_126_3477_n2249), .CO(
        DP_OP_424J2_126_3477_n1636), .S(DP_OP_424J2_126_3477_n1637) );
  FADDX1_HVT DP_OP_424J2_126_3477_U975 ( .A(DP_OP_424J2_126_3477_n2594), .B(
        DP_OP_424J2_126_3477_n2256), .CI(DP_OP_424J2_126_3477_n2909), .CO(
        DP_OP_424J2_126_3477_n1634), .S(DP_OP_424J2_126_3477_n1635) );
  FADDX1_HVT DP_OP_424J2_126_3477_U974 ( .A(DP_OP_424J2_126_3477_n2520), .B(
        DP_OP_424J2_126_3477_n2902), .CI(DP_OP_424J2_126_3477_n2872), .CO(
        DP_OP_424J2_126_3477_n1632), .S(DP_OP_424J2_126_3477_n1633) );
  FADDX1_HVT DP_OP_424J2_126_3477_U973 ( .A(DP_OP_424J2_126_3477_n2432), .B(
        DP_OP_424J2_126_3477_n2865), .CI(DP_OP_424J2_126_3477_n2286), .CO(
        DP_OP_424J2_126_3477_n1630), .S(DP_OP_424J2_126_3477_n1631) );
  FADDX1_HVT DP_OP_424J2_126_3477_U972 ( .A(DP_OP_424J2_126_3477_n2858), .B(
        DP_OP_424J2_126_3477_n2293), .CI(DP_OP_424J2_126_3477_n2828), .CO(
        DP_OP_424J2_126_3477_n1628), .S(DP_OP_424J2_126_3477_n1629) );
  FADDX1_HVT DP_OP_424J2_126_3477_U971 ( .A(DP_OP_424J2_126_3477_n2821), .B(
        DP_OP_424J2_126_3477_n2814), .CI(DP_OP_424J2_126_3477_n2300), .CO(
        DP_OP_424J2_126_3477_n1626), .S(DP_OP_424J2_126_3477_n1627) );
  FADDX1_HVT DP_OP_424J2_126_3477_U970 ( .A(DP_OP_424J2_126_3477_n2425), .B(
        DP_OP_424J2_126_3477_n2330), .CI(DP_OP_424J2_126_3477_n2784), .CO(
        DP_OP_424J2_126_3477_n1624), .S(DP_OP_424J2_126_3477_n1625) );
  FADDX1_HVT DP_OP_424J2_126_3477_U969 ( .A(DP_OP_424J2_126_3477_n2418), .B(
        DP_OP_424J2_126_3477_n2777), .CI(DP_OP_424J2_126_3477_n2770), .CO(
        DP_OP_424J2_126_3477_n1622), .S(DP_OP_424J2_126_3477_n1623) );
  FADDX1_HVT DP_OP_424J2_126_3477_U968 ( .A(DP_OP_424J2_126_3477_n2374), .B(
        DP_OP_424J2_126_3477_n2740), .CI(DP_OP_424J2_126_3477_n2733), .CO(
        DP_OP_424J2_126_3477_n1620), .S(DP_OP_424J2_126_3477_n1621) );
  FADDX1_HVT DP_OP_424J2_126_3477_U967 ( .A(DP_OP_424J2_126_3477_n2337), .B(
        DP_OP_424J2_126_3477_n2726), .CI(DP_OP_424J2_126_3477_n2696), .CO(
        DP_OP_424J2_126_3477_n1618), .S(DP_OP_424J2_126_3477_n1619) );
  FADDX1_HVT DP_OP_424J2_126_3477_U966 ( .A(DP_OP_424J2_126_3477_n2608), .B(
        DP_OP_424J2_126_3477_n2689), .CI(DP_OP_424J2_126_3477_n2344), .CO(
        DP_OP_424J2_126_3477_n1616), .S(DP_OP_424J2_126_3477_n1617) );
  FADDX1_HVT DP_OP_424J2_126_3477_U965 ( .A(DP_OP_424J2_126_3477_n2462), .B(
        DP_OP_424J2_126_3477_n2381), .CI(DP_OP_424J2_126_3477_n2682), .CO(
        DP_OP_424J2_126_3477_n1614), .S(DP_OP_424J2_126_3477_n1615) );
  FADDX1_HVT DP_OP_424J2_126_3477_U964 ( .A(DP_OP_424J2_126_3477_n2652), .B(
        DP_OP_424J2_126_3477_n2388), .CI(DP_OP_424J2_126_3477_n2601), .CO(
        DP_OP_424J2_126_3477_n1612), .S(DP_OP_424J2_126_3477_n1613) );
  FADDX1_HVT DP_OP_424J2_126_3477_U963 ( .A(DP_OP_424J2_126_3477_n2645), .B(
        DP_OP_424J2_126_3477_n2638), .CI(DP_OP_424J2_126_3477_n1784), .CO(
        DP_OP_424J2_126_3477_n1610), .S(DP_OP_424J2_126_3477_n1611) );
  FADDX1_HVT DP_OP_424J2_126_3477_U962 ( .A(DP_OP_424J2_126_3477_n1760), .B(
        DP_OP_424J2_126_3477_n1782), .CI(DP_OP_424J2_126_3477_n1736), .CO(
        DP_OP_424J2_126_3477_n1608), .S(DP_OP_424J2_126_3477_n1609) );
  FADDX1_HVT DP_OP_424J2_126_3477_U961 ( .A(DP_OP_424J2_126_3477_n1758), .B(
        DP_OP_424J2_126_3477_n1780), .CI(DP_OP_424J2_126_3477_n1778), .CO(
        DP_OP_424J2_126_3477_n1606), .S(DP_OP_424J2_126_3477_n1607) );
  FADDX1_HVT DP_OP_424J2_126_3477_U960 ( .A(DP_OP_424J2_126_3477_n1752), .B(
        DP_OP_424J2_126_3477_n1776), .CI(DP_OP_424J2_126_3477_n1774), .CO(
        DP_OP_424J2_126_3477_n1604), .S(DP_OP_424J2_126_3477_n1605) );
  FADDX1_HVT DP_OP_424J2_126_3477_U959 ( .A(DP_OP_424J2_126_3477_n1748), .B(
        DP_OP_424J2_126_3477_n1738), .CI(DP_OP_424J2_126_3477_n1740), .CO(
        DP_OP_424J2_126_3477_n1602), .S(DP_OP_424J2_126_3477_n1603) );
  FADDX1_HVT DP_OP_424J2_126_3477_U958 ( .A(DP_OP_424J2_126_3477_n1746), .B(
        DP_OP_424J2_126_3477_n1772), .CI(DP_OP_424J2_126_3477_n1742), .CO(
        DP_OP_424J2_126_3477_n1600), .S(DP_OP_424J2_126_3477_n1601) );
  FADDX1_HVT DP_OP_424J2_126_3477_U957 ( .A(DP_OP_424J2_126_3477_n1744), .B(
        DP_OP_424J2_126_3477_n1770), .CI(DP_OP_424J2_126_3477_n1768), .CO(
        DP_OP_424J2_126_3477_n1598), .S(DP_OP_424J2_126_3477_n1599) );
  FADDX1_HVT DP_OP_424J2_126_3477_U956 ( .A(DP_OP_424J2_126_3477_n1756), .B(
        DP_OP_424J2_126_3477_n1766), .CI(DP_OP_424J2_126_3477_n1750), .CO(
        DP_OP_424J2_126_3477_n1596), .S(DP_OP_424J2_126_3477_n1597) );
  FADDX1_HVT DP_OP_424J2_126_3477_U955 ( .A(DP_OP_424J2_126_3477_n1764), .B(
        DP_OP_424J2_126_3477_n1762), .CI(DP_OP_424J2_126_3477_n1754), .CO(
        DP_OP_424J2_126_3477_n1594), .S(DP_OP_424J2_126_3477_n1595) );
  FADDX1_HVT DP_OP_424J2_126_3477_U954 ( .A(DP_OP_424J2_126_3477_n1673), .B(
        DP_OP_424J2_126_3477_n1675), .CI(DP_OP_424J2_126_3477_n1661), .CO(
        DP_OP_424J2_126_3477_n1592), .S(DP_OP_424J2_126_3477_n1593) );
  FADDX1_HVT DP_OP_424J2_126_3477_U953 ( .A(DP_OP_424J2_126_3477_n1667), .B(
        DP_OP_424J2_126_3477_n1669), .CI(DP_OP_424J2_126_3477_n1734), .CO(
        DP_OP_424J2_126_3477_n1590), .S(DP_OP_424J2_126_3477_n1591) );
  FADDX1_HVT DP_OP_424J2_126_3477_U952 ( .A(DP_OP_424J2_126_3477_n1663), .B(
        DP_OP_424J2_126_3477_n1665), .CI(DP_OP_424J2_126_3477_n1671), .CO(
        DP_OP_424J2_126_3477_n1588), .S(DP_OP_424J2_126_3477_n1589) );
  FADDX1_HVT DP_OP_424J2_126_3477_U951 ( .A(DP_OP_424J2_126_3477_n1677), .B(
        DP_OP_424J2_126_3477_n1627), .CI(DP_OP_424J2_126_3477_n1625), .CO(
        DP_OP_424J2_126_3477_n1586), .S(DP_OP_424J2_126_3477_n1587) );
  FADDX1_HVT DP_OP_424J2_126_3477_U950 ( .A(DP_OP_424J2_126_3477_n1629), .B(
        DP_OP_424J2_126_3477_n1645), .CI(DP_OP_424J2_126_3477_n1653), .CO(
        DP_OP_424J2_126_3477_n1584), .S(DP_OP_424J2_126_3477_n1585) );
  FADDX1_HVT DP_OP_424J2_126_3477_U949 ( .A(DP_OP_424J2_126_3477_n1621), .B(
        DP_OP_424J2_126_3477_n1641), .CI(DP_OP_424J2_126_3477_n1639), .CO(
        DP_OP_424J2_126_3477_n1582), .S(DP_OP_424J2_126_3477_n1583) );
  FADDX1_HVT DP_OP_424J2_126_3477_U948 ( .A(DP_OP_424J2_126_3477_n1619), .B(
        DP_OP_424J2_126_3477_n1655), .CI(DP_OP_424J2_126_3477_n1643), .CO(
        DP_OP_424J2_126_3477_n1580), .S(DP_OP_424J2_126_3477_n1581) );
  FADDX1_HVT DP_OP_424J2_126_3477_U947 ( .A(DP_OP_424J2_126_3477_n1617), .B(
        DP_OP_424J2_126_3477_n1649), .CI(DP_OP_424J2_126_3477_n1651), .CO(
        DP_OP_424J2_126_3477_n1578), .S(DP_OP_424J2_126_3477_n1579) );
  FADDX1_HVT DP_OP_424J2_126_3477_U946 ( .A(DP_OP_424J2_126_3477_n1615), .B(
        DP_OP_424J2_126_3477_n1647), .CI(DP_OP_424J2_126_3477_n1659), .CO(
        DP_OP_424J2_126_3477_n1576), .S(DP_OP_424J2_126_3477_n1577) );
  FADDX1_HVT DP_OP_424J2_126_3477_U945 ( .A(DP_OP_424J2_126_3477_n1637), .B(
        DP_OP_424J2_126_3477_n1657), .CI(DP_OP_424J2_126_3477_n1613), .CO(
        DP_OP_424J2_126_3477_n1574), .S(DP_OP_424J2_126_3477_n1575) );
  FADDX1_HVT DP_OP_424J2_126_3477_U944 ( .A(DP_OP_424J2_126_3477_n1623), .B(
        DP_OP_424J2_126_3477_n1633), .CI(DP_OP_424J2_126_3477_n1635), .CO(
        DP_OP_424J2_126_3477_n1572), .S(DP_OP_424J2_126_3477_n1573) );
  FADDX1_HVT DP_OP_424J2_126_3477_U943 ( .A(DP_OP_424J2_126_3477_n1631), .B(
        DP_OP_424J2_126_3477_n1611), .CI(DP_OP_424J2_126_3477_n1732), .CO(
        DP_OP_424J2_126_3477_n1570), .S(DP_OP_424J2_126_3477_n1571) );
  FADDX1_HVT DP_OP_424J2_126_3477_U942 ( .A(DP_OP_424J2_126_3477_n1730), .B(
        DP_OP_424J2_126_3477_n1728), .CI(DP_OP_424J2_126_3477_n1726), .CO(
        DP_OP_424J2_126_3477_n1568), .S(DP_OP_424J2_126_3477_n1569) );
  FADDX1_HVT DP_OP_424J2_126_3477_U941 ( .A(DP_OP_424J2_126_3477_n1724), .B(
        DP_OP_424J2_126_3477_n1722), .CI(DP_OP_424J2_126_3477_n1710), .CO(
        DP_OP_424J2_126_3477_n1566), .S(DP_OP_424J2_126_3477_n1567) );
  FADDX1_HVT DP_OP_424J2_126_3477_U940 ( .A(DP_OP_424J2_126_3477_n1708), .B(
        DP_OP_424J2_126_3477_n1609), .CI(DP_OP_424J2_126_3477_n1706), .CO(
        DP_OP_424J2_126_3477_n1564), .S(DP_OP_424J2_126_3477_n1565) );
  FADDX1_HVT DP_OP_424J2_126_3477_U939 ( .A(DP_OP_424J2_126_3477_n1720), .B(
        DP_OP_424J2_126_3477_n1599), .CI(DP_OP_424J2_126_3477_n1607), .CO(
        DP_OP_424J2_126_3477_n1562), .S(DP_OP_424J2_126_3477_n1563) );
  FADDX1_HVT DP_OP_424J2_126_3477_U938 ( .A(DP_OP_424J2_126_3477_n1718), .B(
        DP_OP_424J2_126_3477_n1597), .CI(DP_OP_424J2_126_3477_n1601), .CO(
        DP_OP_424J2_126_3477_n1560), .S(DP_OP_424J2_126_3477_n1561) );
  FADDX1_HVT DP_OP_424J2_126_3477_U937 ( .A(DP_OP_424J2_126_3477_n1714), .B(
        DP_OP_424J2_126_3477_n1605), .CI(DP_OP_424J2_126_3477_n1603), .CO(
        DP_OP_424J2_126_3477_n1558), .S(DP_OP_424J2_126_3477_n1559) );
  FADDX1_HVT DP_OP_424J2_126_3477_U936 ( .A(DP_OP_424J2_126_3477_n1712), .B(
        DP_OP_424J2_126_3477_n1716), .CI(DP_OP_424J2_126_3477_n1595), .CO(
        DP_OP_424J2_126_3477_n1556), .S(DP_OP_424J2_126_3477_n1557) );
  FADDX1_HVT DP_OP_424J2_126_3477_U935 ( .A(DP_OP_424J2_126_3477_n1591), .B(
        DP_OP_424J2_126_3477_n1593), .CI(DP_OP_424J2_126_3477_n1587), .CO(
        DP_OP_424J2_126_3477_n1554), .S(DP_OP_424J2_126_3477_n1555) );
  FADDX1_HVT DP_OP_424J2_126_3477_U934 ( .A(DP_OP_424J2_126_3477_n1589), .B(
        DP_OP_424J2_126_3477_n1575), .CI(DP_OP_424J2_126_3477_n1577), .CO(
        DP_OP_424J2_126_3477_n1552), .S(DP_OP_424J2_126_3477_n1553) );
  FADDX1_HVT DP_OP_424J2_126_3477_U933 ( .A(DP_OP_424J2_126_3477_n1583), .B(
        DP_OP_424J2_126_3477_n1581), .CI(DP_OP_424J2_126_3477_n1704), .CO(
        DP_OP_424J2_126_3477_n1550), .S(DP_OP_424J2_126_3477_n1551) );
  FADDX1_HVT DP_OP_424J2_126_3477_U932 ( .A(DP_OP_424J2_126_3477_n1579), .B(
        DP_OP_424J2_126_3477_n1573), .CI(DP_OP_424J2_126_3477_n1585), .CO(
        DP_OP_424J2_126_3477_n1548), .S(DP_OP_424J2_126_3477_n1549) );
  FADDX1_HVT DP_OP_424J2_126_3477_U931 ( .A(DP_OP_424J2_126_3477_n1571), .B(
        DP_OP_424J2_126_3477_n1702), .CI(DP_OP_424J2_126_3477_n1698), .CO(
        DP_OP_424J2_126_3477_n1546), .S(DP_OP_424J2_126_3477_n1547) );
  FADDX1_HVT DP_OP_424J2_126_3477_U930 ( .A(DP_OP_424J2_126_3477_n1700), .B(
        DP_OP_424J2_126_3477_n1569), .CI(DP_OP_424J2_126_3477_n1696), .CO(
        DP_OP_424J2_126_3477_n1544), .S(DP_OP_424J2_126_3477_n1545) );
  FADDX1_HVT DP_OP_424J2_126_3477_U929 ( .A(DP_OP_424J2_126_3477_n1567), .B(
        DP_OP_424J2_126_3477_n1557), .CI(DP_OP_424J2_126_3477_n1559), .CO(
        DP_OP_424J2_126_3477_n1542), .S(DP_OP_424J2_126_3477_n1543) );
  FADDX1_HVT DP_OP_424J2_126_3477_U928 ( .A(DP_OP_424J2_126_3477_n1694), .B(
        DP_OP_424J2_126_3477_n1561), .CI(DP_OP_424J2_126_3477_n1692), .CO(
        DP_OP_424J2_126_3477_n1540), .S(DP_OP_424J2_126_3477_n1541) );
  FADDX1_HVT DP_OP_424J2_126_3477_U927 ( .A(DP_OP_424J2_126_3477_n1565), .B(
        DP_OP_424J2_126_3477_n1563), .CI(DP_OP_424J2_126_3477_n1555), .CO(
        DP_OP_424J2_126_3477_n1538), .S(DP_OP_424J2_126_3477_n1539) );
  FADDX1_HVT DP_OP_424J2_126_3477_U926 ( .A(DP_OP_424J2_126_3477_n1690), .B(
        DP_OP_424J2_126_3477_n1553), .CI(DP_OP_424J2_126_3477_n1549), .CO(
        DP_OP_424J2_126_3477_n1536), .S(DP_OP_424J2_126_3477_n1537) );
  FADDX1_HVT DP_OP_424J2_126_3477_U925 ( .A(DP_OP_424J2_126_3477_n1551), .B(
        DP_OP_424J2_126_3477_n1688), .CI(DP_OP_424J2_126_3477_n1547), .CO(
        DP_OP_424J2_126_3477_n1534), .S(DP_OP_424J2_126_3477_n1535) );
  FADDX1_HVT DP_OP_424J2_126_3477_U924 ( .A(DP_OP_424J2_126_3477_n1686), .B(
        DP_OP_424J2_126_3477_n1545), .CI(DP_OP_424J2_126_3477_n1684), .CO(
        DP_OP_424J2_126_3477_n1532), .S(DP_OP_424J2_126_3477_n1533) );
  FADDX1_HVT DP_OP_424J2_126_3477_U923 ( .A(DP_OP_424J2_126_3477_n1543), .B(
        DP_OP_424J2_126_3477_n1541), .CI(DP_OP_424J2_126_3477_n1539), .CO(
        DP_OP_424J2_126_3477_n1530), .S(DP_OP_424J2_126_3477_n1531) );
  FADDX1_HVT DP_OP_424J2_126_3477_U922 ( .A(DP_OP_424J2_126_3477_n1537), .B(
        DP_OP_424J2_126_3477_n1682), .CI(DP_OP_424J2_126_3477_n1535), .CO(
        DP_OP_424J2_126_3477_n1528), .S(DP_OP_424J2_126_3477_n1529) );
  FADDX1_HVT DP_OP_424J2_126_3477_U921 ( .A(DP_OP_424J2_126_3477_n1680), .B(
        DP_OP_424J2_126_3477_n1533), .CI(DP_OP_424J2_126_3477_n1531), .CO(
        DP_OP_424J2_126_3477_n1526), .S(DP_OP_424J2_126_3477_n1527) );
  FADDX1_HVT DP_OP_424J2_126_3477_U920 ( .A(DP_OP_424J2_126_3477_n1678), .B(
        DP_OP_424J2_126_3477_n1926), .CI(DP_OP_424J2_126_3477_n1882), .CO(
        DP_OP_424J2_126_3477_n1524), .S(DP_OP_424J2_126_3477_n1525) );
  FADDX1_HVT DP_OP_424J2_126_3477_U919 ( .A(DP_OP_424J2_126_3477_n2981), .B(
        DP_OP_424J2_126_3477_n2498), .CI(DP_OP_424J2_126_3477_n2366), .CO(
        DP_OP_424J2_126_3477_n1522), .S(DP_OP_424J2_126_3477_n1523) );
  FADDX1_HVT DP_OP_424J2_126_3477_U918 ( .A(DP_OP_424J2_126_3477_n2894), .B(
        DP_OP_424J2_126_3477_n2630), .CI(DP_OP_424J2_126_3477_n2278), .CO(
        DP_OP_424J2_126_3477_n1520), .S(DP_OP_424J2_126_3477_n1521) );
  FADDX1_HVT DP_OP_424J2_126_3477_U917 ( .A(DP_OP_424J2_126_3477_n2058), .B(
        DP_OP_424J2_126_3477_n2586), .CI(DP_OP_424J2_126_3477_n2806), .CO(
        DP_OP_424J2_126_3477_n1518), .S(DP_OP_424J2_126_3477_n1519) );
  FADDX1_HVT DP_OP_424J2_126_3477_U916 ( .A(DP_OP_424J2_126_3477_n2146), .B(
        DP_OP_424J2_126_3477_n2322), .CI(DP_OP_424J2_126_3477_n2410), .CO(
        DP_OP_424J2_126_3477_n1516), .S(DP_OP_424J2_126_3477_n1517) );
  FADDX1_HVT DP_OP_424J2_126_3477_U915 ( .A(DP_OP_424J2_126_3477_n2762), .B(
        DP_OP_424J2_126_3477_n2234), .CI(DP_OP_424J2_126_3477_n2850), .CO(
        DP_OP_424J2_126_3477_n1514), .S(DP_OP_424J2_126_3477_n1515) );
  FADDX1_HVT DP_OP_424J2_126_3477_U914 ( .A(DP_OP_424J2_126_3477_n2102), .B(
        DP_OP_424J2_126_3477_n2454), .CI(DP_OP_424J2_126_3477_n2542), .CO(
        DP_OP_424J2_126_3477_n1512), .S(DP_OP_424J2_126_3477_n1513) );
  FADDX1_HVT DP_OP_424J2_126_3477_U913 ( .A(DP_OP_424J2_126_3477_n2938), .B(
        DP_OP_424J2_126_3477_n2674), .CI(DP_OP_424J2_126_3477_n2718), .CO(
        DP_OP_424J2_126_3477_n1510), .S(DP_OP_424J2_126_3477_n1511) );
  FADDX1_HVT DP_OP_424J2_126_3477_U912 ( .A(DP_OP_424J2_126_3477_n2014), .B(
        DP_OP_424J2_126_3477_n2190), .CI(DP_OP_424J2_126_3477_n1970), .CO(
        DP_OP_424J2_126_3477_n1508), .S(DP_OP_424J2_126_3477_n1509) );
  FADDX1_HVT DP_OP_424J2_126_3477_U911 ( .A(DP_OP_424J2_126_3477_n2505), .B(
        DP_OP_424J2_126_3477_n1940), .CI(DP_OP_424J2_126_3477_n1933), .CO(
        DP_OP_424J2_126_3477_n1506), .S(DP_OP_424J2_126_3477_n1507) );
  FADDX1_HVT DP_OP_424J2_126_3477_U910 ( .A(DP_OP_424J2_126_3477_n3001), .B(
        DP_OP_424J2_126_3477_n1947), .CI(DP_OP_424J2_126_3477_n1977), .CO(
        DP_OP_424J2_126_3477_n1504), .S(DP_OP_424J2_126_3477_n1505) );
  FADDX1_HVT DP_OP_424J2_126_3477_U909 ( .A(DP_OP_424J2_126_3477_n2387), .B(
        DP_OP_424J2_126_3477_n2994), .CI(DP_OP_424J2_126_3477_n1984), .CO(
        DP_OP_424J2_126_3477_n1502), .S(DP_OP_424J2_126_3477_n1503) );
  FADDX1_HVT DP_OP_424J2_126_3477_U908 ( .A(DP_OP_424J2_126_3477_n2380), .B(
        DP_OP_424J2_126_3477_n2987), .CI(DP_OP_424J2_126_3477_n1991), .CO(
        DP_OP_424J2_126_3477_n1500), .S(DP_OP_424J2_126_3477_n1501) );
  FADDX1_HVT DP_OP_424J2_126_3477_U907 ( .A(DP_OP_424J2_126_3477_n2959), .B(
        DP_OP_424J2_126_3477_n2021), .CI(DP_OP_424J2_126_3477_n2028), .CO(
        DP_OP_424J2_126_3477_n1498), .S(DP_OP_424J2_126_3477_n1499) );
  FADDX1_HVT DP_OP_424J2_126_3477_U906 ( .A(DP_OP_424J2_126_3477_n2417), .B(
        DP_OP_424J2_126_3477_n2952), .CI(DP_OP_424J2_126_3477_n2945), .CO(
        DP_OP_424J2_126_3477_n1496), .S(DP_OP_424J2_126_3477_n1497) );
  FADDX1_HVT DP_OP_424J2_126_3477_U905 ( .A(DP_OP_424J2_126_3477_n2343), .B(
        DP_OP_424J2_126_3477_n2915), .CI(DP_OP_424J2_126_3477_n2908), .CO(
        DP_OP_424J2_126_3477_n1494), .S(DP_OP_424J2_126_3477_n1495) );
  FADDX1_HVT DP_OP_424J2_126_3477_U904 ( .A(DP_OP_424J2_126_3477_n2336), .B(
        DP_OP_424J2_126_3477_n2901), .CI(DP_OP_424J2_126_3477_n2035), .CO(
        DP_OP_424J2_126_3477_n1492), .S(DP_OP_424J2_126_3477_n1493) );
  FADDX1_HVT DP_OP_424J2_126_3477_U903 ( .A(DP_OP_424J2_126_3477_n2329), .B(
        DP_OP_424J2_126_3477_n2871), .CI(DP_OP_424J2_126_3477_n2864), .CO(
        DP_OP_424J2_126_3477_n1490), .S(DP_OP_424J2_126_3477_n1491) );
  FADDX1_HVT DP_OP_424J2_126_3477_U902 ( .A(DP_OP_424J2_126_3477_n2299), .B(
        DP_OP_424J2_126_3477_n2857), .CI(DP_OP_424J2_126_3477_n2065), .CO(
        DP_OP_424J2_126_3477_n1488), .S(DP_OP_424J2_126_3477_n1489) );
  FADDX1_HVT DP_OP_424J2_126_3477_U901 ( .A(DP_OP_424J2_126_3477_n2292), .B(
        DP_OP_424J2_126_3477_n2072), .CI(DP_OP_424J2_126_3477_n2079), .CO(
        DP_OP_424J2_126_3477_n1486), .S(DP_OP_424J2_126_3477_n1487) );
  FADDX1_HVT DP_OP_424J2_126_3477_U900 ( .A(DP_OP_424J2_126_3477_n2373), .B(
        DP_OP_424J2_126_3477_n2109), .CI(DP_OP_424J2_126_3477_n2827), .CO(
        DP_OP_424J2_126_3477_n1484), .S(DP_OP_424J2_126_3477_n1485) );
  FADDX1_HVT DP_OP_424J2_126_3477_U899 ( .A(DP_OP_424J2_126_3477_n2424), .B(
        DP_OP_424J2_126_3477_n2820), .CI(DP_OP_424J2_126_3477_n2813), .CO(
        DP_OP_424J2_126_3477_n1482), .S(DP_OP_424J2_126_3477_n1483) );
  FADDX1_HVT DP_OP_424J2_126_3477_U898 ( .A(DP_OP_424J2_126_3477_n2783), .B(
        DP_OP_424J2_126_3477_n2116), .CI(DP_OP_424J2_126_3477_n2123), .CO(
        DP_OP_424J2_126_3477_n1480), .S(DP_OP_424J2_126_3477_n1481) );
  FADDX1_HVT DP_OP_424J2_126_3477_U897 ( .A(DP_OP_424J2_126_3477_n2556), .B(
        DP_OP_424J2_126_3477_n2153), .CI(DP_OP_424J2_126_3477_n2160), .CO(
        DP_OP_424J2_126_3477_n1478), .S(DP_OP_424J2_126_3477_n1479) );
  FADDX1_HVT DP_OP_424J2_126_3477_U896 ( .A(DP_OP_424J2_126_3477_n2776), .B(
        DP_OP_424J2_126_3477_n2167), .CI(DP_OP_424J2_126_3477_n2197), .CO(
        DP_OP_424J2_126_3477_n1476), .S(DP_OP_424J2_126_3477_n1477) );
  FADDX1_HVT DP_OP_424J2_126_3477_U895 ( .A(DP_OP_424J2_126_3477_n2769), .B(
        DP_OP_424J2_126_3477_n2204), .CI(DP_OP_424J2_126_3477_n2211), .CO(
        DP_OP_424J2_126_3477_n1474), .S(DP_OP_424J2_126_3477_n1475) );
  FADDX1_HVT DP_OP_424J2_126_3477_U894 ( .A(DP_OP_424J2_126_3477_n2739), .B(
        DP_OP_424J2_126_3477_n2241), .CI(DP_OP_424J2_126_3477_n2248), .CO(
        DP_OP_424J2_126_3477_n1472), .S(DP_OP_424J2_126_3477_n1473) );
  FADDX1_HVT DP_OP_424J2_126_3477_U893 ( .A(DP_OP_424J2_126_3477_n2732), .B(
        DP_OP_424J2_126_3477_n2255), .CI(DP_OP_424J2_126_3477_n2285), .CO(
        DP_OP_424J2_126_3477_n1470), .S(DP_OP_424J2_126_3477_n1471) );
  FADDX1_HVT DP_OP_424J2_126_3477_U892 ( .A(DP_OP_424J2_126_3477_n2725), .B(
        DP_OP_424J2_126_3477_n2431), .CI(DP_OP_424J2_126_3477_n2461), .CO(
        DP_OP_424J2_126_3477_n1468), .S(DP_OP_424J2_126_3477_n1469) );
  FADDX1_HVT DP_OP_424J2_126_3477_U891 ( .A(DP_OP_424J2_126_3477_n2695), .B(
        DP_OP_424J2_126_3477_n2468), .CI(DP_OP_424J2_126_3477_n2688), .CO(
        DP_OP_424J2_126_3477_n1466), .S(DP_OP_424J2_126_3477_n1467) );
  FADDX1_HVT DP_OP_424J2_126_3477_U890 ( .A(DP_OP_424J2_126_3477_n2593), .B(
        DP_OP_424J2_126_3477_n2475), .CI(DP_OP_424J2_126_3477_n2512), .CO(
        DP_OP_424J2_126_3477_n1464), .S(DP_OP_424J2_126_3477_n1465) );
  FADDX1_HVT DP_OP_424J2_126_3477_U889 ( .A(DP_OP_424J2_126_3477_n2563), .B(
        DP_OP_424J2_126_3477_n2519), .CI(DP_OP_424J2_126_3477_n2681), .CO(
        DP_OP_424J2_126_3477_n1462), .S(DP_OP_424J2_126_3477_n1463) );
  FADDX1_HVT DP_OP_424J2_126_3477_U888 ( .A(DP_OP_424J2_126_3477_n2637), .B(
        DP_OP_424J2_126_3477_n2549), .CI(DP_OP_424J2_126_3477_n2651), .CO(
        DP_OP_424J2_126_3477_n1460), .S(DP_OP_424J2_126_3477_n1461) );
  FADDX1_HVT DP_OP_424J2_126_3477_U887 ( .A(DP_OP_424J2_126_3477_n2600), .B(
        DP_OP_424J2_126_3477_n2607), .CI(DP_OP_424J2_126_3477_n2644), .CO(
        DP_OP_424J2_126_3477_n1458), .S(DP_OP_424J2_126_3477_n1459) );
  FADDX1_HVT DP_OP_424J2_126_3477_U886 ( .A(DP_OP_424J2_126_3477_n1666), .B(
        DP_OP_424J2_126_3477_n1662), .CI(DP_OP_424J2_126_3477_n1660), .CO(
        DP_OP_424J2_126_3477_n1456), .S(DP_OP_424J2_126_3477_n1457) );
  FADDX1_HVT DP_OP_424J2_126_3477_U885 ( .A(DP_OP_424J2_126_3477_n1664), .B(
        DP_OP_424J2_126_3477_n1668), .CI(DP_OP_424J2_126_3477_n1670), .CO(
        DP_OP_424J2_126_3477_n1454), .S(DP_OP_424J2_126_3477_n1455) );
  FADDX1_HVT DP_OP_424J2_126_3477_U884 ( .A(DP_OP_424J2_126_3477_n1672), .B(
        DP_OP_424J2_126_3477_n1674), .CI(DP_OP_424J2_126_3477_n1676), .CO(
        DP_OP_424J2_126_3477_n1452), .S(DP_OP_424J2_126_3477_n1453) );
  FADDX1_HVT DP_OP_424J2_126_3477_U883 ( .A(DP_OP_424J2_126_3477_n1636), .B(
        DP_OP_424J2_126_3477_n1658), .CI(DP_OP_424J2_126_3477_n1656), .CO(
        DP_OP_424J2_126_3477_n1450), .S(DP_OP_424J2_126_3477_n1451) );
  FADDX1_HVT DP_OP_424J2_126_3477_U882 ( .A(DP_OP_424J2_126_3477_n1632), .B(
        DP_OP_424J2_126_3477_n1654), .CI(DP_OP_424J2_126_3477_n1652), .CO(
        DP_OP_424J2_126_3477_n1448), .S(DP_OP_424J2_126_3477_n1449) );
  FADDX1_HVT DP_OP_424J2_126_3477_U881 ( .A(DP_OP_424J2_126_3477_n1626), .B(
        DP_OP_424J2_126_3477_n1650), .CI(DP_OP_424J2_126_3477_n1648), .CO(
        DP_OP_424J2_126_3477_n1446), .S(DP_OP_424J2_126_3477_n1447) );
  FADDX1_HVT DP_OP_424J2_126_3477_U880 ( .A(DP_OP_424J2_126_3477_n1622), .B(
        DP_OP_424J2_126_3477_n1646), .CI(DP_OP_424J2_126_3477_n1612), .CO(
        DP_OP_424J2_126_3477_n1444), .S(DP_OP_424J2_126_3477_n1445) );
  FADDX1_HVT DP_OP_424J2_126_3477_U879 ( .A(DP_OP_424J2_126_3477_n1618), .B(
        DP_OP_424J2_126_3477_n1644), .CI(DP_OP_424J2_126_3477_n1642), .CO(
        DP_OP_424J2_126_3477_n1442), .S(DP_OP_424J2_126_3477_n1443) );
  FADDX1_HVT DP_OP_424J2_126_3477_U878 ( .A(DP_OP_424J2_126_3477_n1628), .B(
        DP_OP_424J2_126_3477_n1640), .CI(DP_OP_424J2_126_3477_n1638), .CO(
        DP_OP_424J2_126_3477_n1440), .S(DP_OP_424J2_126_3477_n1441) );
  FADDX1_HVT DP_OP_424J2_126_3477_U877 ( .A(DP_OP_424J2_126_3477_n1620), .B(
        DP_OP_424J2_126_3477_n1634), .CI(DP_OP_424J2_126_3477_n1630), .CO(
        DP_OP_424J2_126_3477_n1438), .S(DP_OP_424J2_126_3477_n1439) );
  FADDX1_HVT DP_OP_424J2_126_3477_U876 ( .A(DP_OP_424J2_126_3477_n1616), .B(
        DP_OP_424J2_126_3477_n1624), .CI(DP_OP_424J2_126_3477_n1614), .CO(
        DP_OP_424J2_126_3477_n1436), .S(DP_OP_424J2_126_3477_n1437) );
  FADDX1_HVT DP_OP_424J2_126_3477_U875 ( .A(DP_OP_424J2_126_3477_n1525), .B(
        DP_OP_424J2_126_3477_n1509), .CI(DP_OP_424J2_126_3477_n1610), .CO(
        DP_OP_424J2_126_3477_n1434), .S(DP_OP_424J2_126_3477_n1435) );
  FADDX1_HVT DP_OP_424J2_126_3477_U874 ( .A(DP_OP_424J2_126_3477_n1523), .B(
        DP_OP_424J2_126_3477_n1511), .CI(DP_OP_424J2_126_3477_n1513), .CO(
        DP_OP_424J2_126_3477_n1432), .S(DP_OP_424J2_126_3477_n1433) );
  FADDX1_HVT DP_OP_424J2_126_3477_U873 ( .A(DP_OP_424J2_126_3477_n1519), .B(
        DP_OP_424J2_126_3477_n1517), .CI(DP_OP_424J2_126_3477_n1521), .CO(
        DP_OP_424J2_126_3477_n1430), .S(DP_OP_424J2_126_3477_n1431) );
  FADDX1_HVT DP_OP_424J2_126_3477_U872 ( .A(DP_OP_424J2_126_3477_n1515), .B(
        DP_OP_424J2_126_3477_n1495), .CI(DP_OP_424J2_126_3477_n1499), .CO(
        DP_OP_424J2_126_3477_n1428), .S(DP_OP_424J2_126_3477_n1429) );
  FADDX1_HVT DP_OP_424J2_126_3477_U871 ( .A(DP_OP_424J2_126_3477_n1497), .B(
        DP_OP_424J2_126_3477_n1505), .CI(DP_OP_424J2_126_3477_n1503), .CO(
        DP_OP_424J2_126_3477_n1426), .S(DP_OP_424J2_126_3477_n1427) );
  FADDX1_HVT DP_OP_424J2_126_3477_U870 ( .A(DP_OP_424J2_126_3477_n1507), .B(
        DP_OP_424J2_126_3477_n1485), .CI(DP_OP_424J2_126_3477_n1479), .CO(
        DP_OP_424J2_126_3477_n1424), .S(DP_OP_424J2_126_3477_n1425) );
  FADDX1_HVT DP_OP_424J2_126_3477_U869 ( .A(DP_OP_424J2_126_3477_n1487), .B(
        DP_OP_424J2_126_3477_n1483), .CI(DP_OP_424J2_126_3477_n1477), .CO(
        DP_OP_424J2_126_3477_n1422), .S(DP_OP_424J2_126_3477_n1423) );
  FADDX1_HVT DP_OP_424J2_126_3477_U868 ( .A(DP_OP_424J2_126_3477_n1489), .B(
        DP_OP_424J2_126_3477_n1463), .CI(DP_OP_424J2_126_3477_n1461), .CO(
        DP_OP_424J2_126_3477_n1420), .S(DP_OP_424J2_126_3477_n1421) );
  FADDX1_HVT DP_OP_424J2_126_3477_U867 ( .A(DP_OP_424J2_126_3477_n1475), .B(
        DP_OP_424J2_126_3477_n1471), .CI(DP_OP_424J2_126_3477_n1473), .CO(
        DP_OP_424J2_126_3477_n1418), .S(DP_OP_424J2_126_3477_n1419) );
  FADDX1_HVT DP_OP_424J2_126_3477_U866 ( .A(DP_OP_424J2_126_3477_n1481), .B(
        DP_OP_424J2_126_3477_n1459), .CI(DP_OP_424J2_126_3477_n1467), .CO(
        DP_OP_424J2_126_3477_n1416), .S(DP_OP_424J2_126_3477_n1417) );
  FADDX1_HVT DP_OP_424J2_126_3477_U865 ( .A(DP_OP_424J2_126_3477_n1469), .B(
        DP_OP_424J2_126_3477_n1493), .CI(DP_OP_424J2_126_3477_n1501), .CO(
        DP_OP_424J2_126_3477_n1414), .S(DP_OP_424J2_126_3477_n1415) );
  FADDX1_HVT DP_OP_424J2_126_3477_U864 ( .A(DP_OP_424J2_126_3477_n1465), .B(
        DP_OP_424J2_126_3477_n1491), .CI(DP_OP_424J2_126_3477_n1608), .CO(
        DP_OP_424J2_126_3477_n1412), .S(DP_OP_424J2_126_3477_n1413) );
  FADDX1_HVT DP_OP_424J2_126_3477_U863 ( .A(DP_OP_424J2_126_3477_n1606), .B(
        DP_OP_424J2_126_3477_n1604), .CI(DP_OP_424J2_126_3477_n1602), .CO(
        DP_OP_424J2_126_3477_n1410), .S(DP_OP_424J2_126_3477_n1411) );
  FADDX1_HVT DP_OP_424J2_126_3477_U862 ( .A(DP_OP_424J2_126_3477_n1594), .B(
        DP_OP_424J2_126_3477_n1600), .CI(DP_OP_424J2_126_3477_n1596), .CO(
        DP_OP_424J2_126_3477_n1408), .S(DP_OP_424J2_126_3477_n1409) );
  FADDX1_HVT DP_OP_424J2_126_3477_U861 ( .A(DP_OP_424J2_126_3477_n1598), .B(
        DP_OP_424J2_126_3477_n1592), .CI(DP_OP_424J2_126_3477_n1453), .CO(
        DP_OP_424J2_126_3477_n1406), .S(DP_OP_424J2_126_3477_n1407) );
  FADDX1_HVT DP_OP_424J2_126_3477_U860 ( .A(DP_OP_424J2_126_3477_n1455), .B(
        DP_OP_424J2_126_3477_n1590), .CI(DP_OP_424J2_126_3477_n1586), .CO(
        DP_OP_424J2_126_3477_n1404), .S(DP_OP_424J2_126_3477_n1405) );
  FADDX1_HVT DP_OP_424J2_126_3477_U859 ( .A(DP_OP_424J2_126_3477_n1457), .B(
        DP_OP_424J2_126_3477_n1588), .CI(DP_OP_424J2_126_3477_n1584), .CO(
        DP_OP_424J2_126_3477_n1402), .S(DP_OP_424J2_126_3477_n1403) );
  FADDX1_HVT DP_OP_424J2_126_3477_U858 ( .A(DP_OP_424J2_126_3477_n1574), .B(
        DP_OP_424J2_126_3477_n1437), .CI(DP_OP_424J2_126_3477_n1449), .CO(
        DP_OP_424J2_126_3477_n1400), .S(DP_OP_424J2_126_3477_n1401) );
  FADDX1_HVT DP_OP_424J2_126_3477_U857 ( .A(DP_OP_424J2_126_3477_n1582), .B(
        DP_OP_424J2_126_3477_n1451), .CI(DP_OP_424J2_126_3477_n1447), .CO(
        DP_OP_424J2_126_3477_n1398), .S(DP_OP_424J2_126_3477_n1399) );
  FADDX1_HVT DP_OP_424J2_126_3477_U856 ( .A(DP_OP_424J2_126_3477_n1580), .B(
        DP_OP_424J2_126_3477_n1439), .CI(DP_OP_424J2_126_3477_n1441), .CO(
        DP_OP_424J2_126_3477_n1396), .S(DP_OP_424J2_126_3477_n1397) );
  FADDX1_HVT DP_OP_424J2_126_3477_U855 ( .A(DP_OP_424J2_126_3477_n1578), .B(
        DP_OP_424J2_126_3477_n1445), .CI(DP_OP_424J2_126_3477_n1443), .CO(
        DP_OP_424J2_126_3477_n1394), .S(DP_OP_424J2_126_3477_n1395) );
  FADDX1_HVT DP_OP_424J2_126_3477_U854 ( .A(DP_OP_424J2_126_3477_n1576), .B(
        DP_OP_424J2_126_3477_n1572), .CI(DP_OP_424J2_126_3477_n1433), .CO(
        DP_OP_424J2_126_3477_n1392), .S(DP_OP_424J2_126_3477_n1393) );
  FADDX1_HVT DP_OP_424J2_126_3477_U853 ( .A(DP_OP_424J2_126_3477_n1435), .B(
        DP_OP_424J2_126_3477_n1431), .CI(DP_OP_424J2_126_3477_n1429), .CO(
        DP_OP_424J2_126_3477_n1390), .S(DP_OP_424J2_126_3477_n1391) );
  FADDX1_HVT DP_OP_424J2_126_3477_U852 ( .A(DP_OP_424J2_126_3477_n1570), .B(
        DP_OP_424J2_126_3477_n1421), .CI(DP_OP_424J2_126_3477_n1419), .CO(
        DP_OP_424J2_126_3477_n1388), .S(DP_OP_424J2_126_3477_n1389) );
  FADDX1_HVT DP_OP_424J2_126_3477_U851 ( .A(DP_OP_424J2_126_3477_n1425), .B(
        DP_OP_424J2_126_3477_n1415), .CI(DP_OP_424J2_126_3477_n1417), .CO(
        DP_OP_424J2_126_3477_n1386), .S(DP_OP_424J2_126_3477_n1387) );
  FADDX1_HVT DP_OP_424J2_126_3477_U850 ( .A(DP_OP_424J2_126_3477_n1423), .B(
        DP_OP_424J2_126_3477_n1427), .CI(DP_OP_424J2_126_3477_n1568), .CO(
        DP_OP_424J2_126_3477_n1384), .S(DP_OP_424J2_126_3477_n1385) );
  FADDX1_HVT DP_OP_424J2_126_3477_U849 ( .A(DP_OP_424J2_126_3477_n1566), .B(
        DP_OP_424J2_126_3477_n1413), .CI(DP_OP_424J2_126_3477_n1564), .CO(
        DP_OP_424J2_126_3477_n1382), .S(DP_OP_424J2_126_3477_n1383) );
  FADDX1_HVT DP_OP_424J2_126_3477_U848 ( .A(DP_OP_424J2_126_3477_n1562), .B(
        DP_OP_424J2_126_3477_n1409), .CI(DP_OP_424J2_126_3477_n1411), .CO(
        DP_OP_424J2_126_3477_n1380), .S(DP_OP_424J2_126_3477_n1381) );
  FADDX1_HVT DP_OP_424J2_126_3477_U847 ( .A(DP_OP_424J2_126_3477_n1560), .B(
        DP_OP_424J2_126_3477_n1556), .CI(DP_OP_424J2_126_3477_n1558), .CO(
        DP_OP_424J2_126_3477_n1378), .S(DP_OP_424J2_126_3477_n1379) );
  FADDX1_HVT DP_OP_424J2_126_3477_U846 ( .A(DP_OP_424J2_126_3477_n1407), .B(
        DP_OP_424J2_126_3477_n1554), .CI(DP_OP_424J2_126_3477_n1552), .CO(
        DP_OP_424J2_126_3477_n1376), .S(DP_OP_424J2_126_3477_n1377) );
  FADDX1_HVT DP_OP_424J2_126_3477_U845 ( .A(DP_OP_424J2_126_3477_n1405), .B(
        DP_OP_424J2_126_3477_n1403), .CI(DP_OP_424J2_126_3477_n1399), .CO(
        DP_OP_424J2_126_3477_n1374), .S(DP_OP_424J2_126_3477_n1375) );
  FADDX1_HVT DP_OP_424J2_126_3477_U844 ( .A(DP_OP_424J2_126_3477_n1401), .B(
        DP_OP_424J2_126_3477_n1397), .CI(DP_OP_424J2_126_3477_n1393), .CO(
        DP_OP_424J2_126_3477_n1372), .S(DP_OP_424J2_126_3477_n1373) );
  FADDX1_HVT DP_OP_424J2_126_3477_U843 ( .A(DP_OP_424J2_126_3477_n1550), .B(
        DP_OP_424J2_126_3477_n1395), .CI(DP_OP_424J2_126_3477_n1548), .CO(
        DP_OP_424J2_126_3477_n1370), .S(DP_OP_424J2_126_3477_n1371) );
  FADDX1_HVT DP_OP_424J2_126_3477_U842 ( .A(DP_OP_424J2_126_3477_n1391), .B(
        DP_OP_424J2_126_3477_n1389), .CI(DP_OP_424J2_126_3477_n1387), .CO(
        DP_OP_424J2_126_3477_n1368), .S(DP_OP_424J2_126_3477_n1369) );
  FADDX1_HVT DP_OP_424J2_126_3477_U841 ( .A(DP_OP_424J2_126_3477_n1546), .B(
        DP_OP_424J2_126_3477_n1385), .CI(DP_OP_424J2_126_3477_n1544), .CO(
        DP_OP_424J2_126_3477_n1366), .S(DP_OP_424J2_126_3477_n1367) );
  FADDX1_HVT DP_OP_424J2_126_3477_U840 ( .A(DP_OP_424J2_126_3477_n1383), .B(
        DP_OP_424J2_126_3477_n1542), .CI(DP_OP_424J2_126_3477_n1540), .CO(
        DP_OP_424J2_126_3477_n1364), .S(DP_OP_424J2_126_3477_n1365) );
  FADDX1_HVT DP_OP_424J2_126_3477_U839 ( .A(DP_OP_424J2_126_3477_n1379), .B(
        DP_OP_424J2_126_3477_n1381), .CI(DP_OP_424J2_126_3477_n1538), .CO(
        DP_OP_424J2_126_3477_n1362), .S(DP_OP_424J2_126_3477_n1363) );
  FADDX1_HVT DP_OP_424J2_126_3477_U838 ( .A(DP_OP_424J2_126_3477_n1377), .B(
        DP_OP_424J2_126_3477_n1375), .CI(DP_OP_424J2_126_3477_n1536), .CO(
        DP_OP_424J2_126_3477_n1360), .S(DP_OP_424J2_126_3477_n1361) );
  FADDX1_HVT DP_OP_424J2_126_3477_U837 ( .A(DP_OP_424J2_126_3477_n1371), .B(
        DP_OP_424J2_126_3477_n1373), .CI(DP_OP_424J2_126_3477_n1534), .CO(
        DP_OP_424J2_126_3477_n1358), .S(DP_OP_424J2_126_3477_n1359) );
  FADDX1_HVT DP_OP_424J2_126_3477_U836 ( .A(DP_OP_424J2_126_3477_n1369), .B(
        DP_OP_424J2_126_3477_n1367), .CI(DP_OP_424J2_126_3477_n1532), .CO(
        DP_OP_424J2_126_3477_n1356), .S(DP_OP_424J2_126_3477_n1357) );
  FADDX1_HVT DP_OP_424J2_126_3477_U835 ( .A(DP_OP_424J2_126_3477_n1365), .B(
        DP_OP_424J2_126_3477_n1530), .CI(DP_OP_424J2_126_3477_n1363), .CO(
        DP_OP_424J2_126_3477_n1354), .S(DP_OP_424J2_126_3477_n1355) );
  FADDX1_HVT DP_OP_424J2_126_3477_U834 ( .A(DP_OP_424J2_126_3477_n1361), .B(
        DP_OP_424J2_126_3477_n1528), .CI(DP_OP_424J2_126_3477_n1359), .CO(
        DP_OP_424J2_126_3477_n1352), .S(DP_OP_424J2_126_3477_n1353) );
  FADDX1_HVT DP_OP_424J2_126_3477_U833 ( .A(DP_OP_424J2_126_3477_n1357), .B(
        DP_OP_424J2_126_3477_n1526), .CI(DP_OP_424J2_126_3477_n1355), .CO(
        DP_OP_424J2_126_3477_n1350), .S(DP_OP_424J2_126_3477_n1351) );
  HADDX1_HVT DP_OP_424J2_126_3477_U832 ( .A0(DP_OP_424J2_126_3477_n2980), .B0(
        DP_OP_424J2_126_3477_n1925), .C1(DP_OP_424J2_126_3477_n1348), .SO(
        DP_OP_424J2_126_3477_n1349) );
  FADDX1_HVT DP_OP_424J2_126_3477_U831 ( .A(DP_OP_424J2_126_3477_n2453), .B(
        DP_OP_424J2_126_3477_n2365), .CI(DP_OP_424J2_126_3477_n1881), .CO(
        DP_OP_424J2_126_3477_n1346), .S(DP_OP_424J2_126_3477_n1347) );
  FADDX1_HVT DP_OP_424J2_126_3477_U830 ( .A(DP_OP_424J2_126_3477_n2497), .B(
        DP_OP_424J2_126_3477_n2277), .CI(DP_OP_424J2_126_3477_n2321), .CO(
        DP_OP_424J2_126_3477_n1344), .S(DP_OP_424J2_126_3477_n1345) );
  FADDX1_HVT DP_OP_424J2_126_3477_U829 ( .A(DP_OP_424J2_126_3477_n2805), .B(
        DP_OP_424J2_126_3477_n1969), .CI(DP_OP_424J2_126_3477_n2057), .CO(
        DP_OP_424J2_126_3477_n1342), .S(DP_OP_424J2_126_3477_n1343) );
  FADDX1_HVT DP_OP_424J2_126_3477_U828 ( .A(DP_OP_424J2_126_3477_n2541), .B(
        DP_OP_424J2_126_3477_n2101), .CI(DP_OP_424J2_126_3477_n2629), .CO(
        DP_OP_424J2_126_3477_n1340), .S(DP_OP_424J2_126_3477_n1341) );
  FADDX1_HVT DP_OP_424J2_126_3477_U827 ( .A(DP_OP_424J2_126_3477_n2013), .B(
        DP_OP_424J2_126_3477_n2849), .CI(DP_OP_424J2_126_3477_n2145), .CO(
        DP_OP_424J2_126_3477_n1338), .S(DP_OP_424J2_126_3477_n1339) );
  FADDX1_HVT DP_OP_424J2_126_3477_U826 ( .A(DP_OP_424J2_126_3477_n2409), .B(
        DP_OP_424J2_126_3477_n2893), .CI(DP_OP_424J2_126_3477_n2717), .CO(
        DP_OP_424J2_126_3477_n1336), .S(DP_OP_424J2_126_3477_n1337) );
  FADDX1_HVT DP_OP_424J2_126_3477_U825 ( .A(DP_OP_424J2_126_3477_n2233), .B(
        DP_OP_424J2_126_3477_n2189), .CI(DP_OP_424J2_126_3477_n2673), .CO(
        DP_OP_424J2_126_3477_n1334), .S(DP_OP_424J2_126_3477_n1335) );
  FADDX1_HVT DP_OP_424J2_126_3477_U824 ( .A(DP_OP_424J2_126_3477_n2937), .B(
        DP_OP_424J2_126_3477_n2585), .CI(DP_OP_424J2_126_3477_n2761), .CO(
        DP_OP_424J2_126_3477_n1332), .S(DP_OP_424J2_126_3477_n1333) );
  FADDX1_HVT DP_OP_424J2_126_3477_U823 ( .A(DP_OP_424J2_126_3477_n2379), .B(
        DP_OP_424J2_126_3477_n3000), .CI(DP_OP_424J2_126_3477_n1932), .CO(
        DP_OP_424J2_126_3477_n1330), .S(DP_OP_424J2_126_3477_n1331) );
  FADDX1_HVT DP_OP_424J2_126_3477_U822 ( .A(DP_OP_424J2_126_3477_n2372), .B(
        DP_OP_424J2_126_3477_n1939), .CI(DP_OP_424J2_126_3477_n1946), .CO(
        DP_OP_424J2_126_3477_n1328), .S(DP_OP_424J2_126_3477_n1329) );
  FADDX1_HVT DP_OP_424J2_126_3477_U821 ( .A(DP_OP_424J2_126_3477_n2386), .B(
        DP_OP_424J2_126_3477_n1976), .CI(DP_OP_424J2_126_3477_n2993), .CO(
        DP_OP_424J2_126_3477_n1326), .S(DP_OP_424J2_126_3477_n1327) );
  FADDX1_HVT DP_OP_424J2_126_3477_U820 ( .A(DP_OP_424J2_126_3477_n2342), .B(
        DP_OP_424J2_126_3477_n2986), .CI(DP_OP_424J2_126_3477_n2958), .CO(
        DP_OP_424J2_126_3477_n1324), .S(DP_OP_424J2_126_3477_n1325) );
  FADDX1_HVT DP_OP_424J2_126_3477_U819 ( .A(DP_OP_424J2_126_3477_n2335), .B(
        DP_OP_424J2_126_3477_n2951), .CI(DP_OP_424J2_126_3477_n2944), .CO(
        DP_OP_424J2_126_3477_n1322), .S(DP_OP_424J2_126_3477_n1323) );
  FADDX1_HVT DP_OP_424J2_126_3477_U818 ( .A(DP_OP_424J2_126_3477_n2298), .B(
        DP_OP_424J2_126_3477_n2914), .CI(DP_OP_424J2_126_3477_n2907), .CO(
        DP_OP_424J2_126_3477_n1320), .S(DP_OP_424J2_126_3477_n1321) );
  FADDX1_HVT DP_OP_424J2_126_3477_U817 ( .A(DP_OP_424J2_126_3477_n2291), .B(
        DP_OP_424J2_126_3477_n1983), .CI(DP_OP_424J2_126_3477_n2900), .CO(
        DP_OP_424J2_126_3477_n1318), .S(DP_OP_424J2_126_3477_n1319) );
  FADDX1_HVT DP_OP_424J2_126_3477_U816 ( .A(DP_OP_424J2_126_3477_n2284), .B(
        DP_OP_424J2_126_3477_n2870), .CI(DP_OP_424J2_126_3477_n2863), .CO(
        DP_OP_424J2_126_3477_n1316), .S(DP_OP_424J2_126_3477_n1317) );
  FADDX1_HVT DP_OP_424J2_126_3477_U815 ( .A(DP_OP_424J2_126_3477_n2254), .B(
        DP_OP_424J2_126_3477_n2856), .CI(DP_OP_424J2_126_3477_n1990), .CO(
        DP_OP_424J2_126_3477_n1314), .S(DP_OP_424J2_126_3477_n1315) );
  FADDX1_HVT DP_OP_424J2_126_3477_U814 ( .A(DP_OP_424J2_126_3477_n2247), .B(
        DP_OP_424J2_126_3477_n2020), .CI(DP_OP_424J2_126_3477_n2027), .CO(
        DP_OP_424J2_126_3477_n1312), .S(DP_OP_424J2_126_3477_n1313) );
  FADDX1_HVT DP_OP_424J2_126_3477_U813 ( .A(DP_OP_424J2_126_3477_n2328), .B(
        DP_OP_424J2_126_3477_n2034), .CI(DP_OP_424J2_126_3477_n2826), .CO(
        DP_OP_424J2_126_3477_n1310), .S(DP_OP_424J2_126_3477_n1311) );
  FADDX1_HVT DP_OP_424J2_126_3477_U812 ( .A(DP_OP_424J2_126_3477_n2416), .B(
        DP_OP_424J2_126_3477_n2819), .CI(DP_OP_424J2_126_3477_n2064), .CO(
        DP_OP_424J2_126_3477_n1308), .S(DP_OP_424J2_126_3477_n1309) );
  FADDX1_HVT DP_OP_424J2_126_3477_U811 ( .A(DP_OP_424J2_126_3477_n2812), .B(
        DP_OP_424J2_126_3477_n2071), .CI(DP_OP_424J2_126_3477_n2078), .CO(
        DP_OP_424J2_126_3477_n1306), .S(DP_OP_424J2_126_3477_n1307) );
  FADDX1_HVT DP_OP_424J2_126_3477_U810 ( .A(DP_OP_424J2_126_3477_n2782), .B(
        DP_OP_424J2_126_3477_n2108), .CI(DP_OP_424J2_126_3477_n2115), .CO(
        DP_OP_424J2_126_3477_n1304), .S(DP_OP_424J2_126_3477_n1305) );
  FADDX1_HVT DP_OP_424J2_126_3477_U809 ( .A(DP_OP_424J2_126_3477_n2775), .B(
        DP_OP_424J2_126_3477_n2122), .CI(DP_OP_424J2_126_3477_n2152), .CO(
        DP_OP_424J2_126_3477_n1302), .S(DP_OP_424J2_126_3477_n1303) );
  FADDX1_HVT DP_OP_424J2_126_3477_U808 ( .A(DP_OP_424J2_126_3477_n2768), .B(
        DP_OP_424J2_126_3477_n2159), .CI(DP_OP_424J2_126_3477_n2166), .CO(
        DP_OP_424J2_126_3477_n1300), .S(DP_OP_424J2_126_3477_n1301) );
  FADDX1_HVT DP_OP_424J2_126_3477_U807 ( .A(DP_OP_424J2_126_3477_n2738), .B(
        DP_OP_424J2_126_3477_n2196), .CI(DP_OP_424J2_126_3477_n2203), .CO(
        DP_OP_424J2_126_3477_n1298), .S(DP_OP_424J2_126_3477_n1299) );
  FADDX1_HVT DP_OP_424J2_126_3477_U806 ( .A(DP_OP_424J2_126_3477_n2731), .B(
        DP_OP_424J2_126_3477_n2210), .CI(DP_OP_424J2_126_3477_n2240), .CO(
        DP_OP_424J2_126_3477_n1296), .S(DP_OP_424J2_126_3477_n1297) );
  FADDX1_HVT DP_OP_424J2_126_3477_U805 ( .A(DP_OP_424J2_126_3477_n2724), .B(
        DP_OP_424J2_126_3477_n2423), .CI(DP_OP_424J2_126_3477_n2430), .CO(
        DP_OP_424J2_126_3477_n1294), .S(DP_OP_424J2_126_3477_n1295) );
  FADDX1_HVT DP_OP_424J2_126_3477_U804 ( .A(DP_OP_424J2_126_3477_n2694), .B(
        DP_OP_424J2_126_3477_n2460), .CI(DP_OP_424J2_126_3477_n2467), .CO(
        DP_OP_424J2_126_3477_n1292), .S(DP_OP_424J2_126_3477_n1293) );
  FADDX1_HVT DP_OP_424J2_126_3477_U803 ( .A(DP_OP_424J2_126_3477_n2687), .B(
        DP_OP_424J2_126_3477_n2474), .CI(DP_OP_424J2_126_3477_n2504), .CO(
        DP_OP_424J2_126_3477_n1290), .S(DP_OP_424J2_126_3477_n1291) );
  FADDX1_HVT DP_OP_424J2_126_3477_U802 ( .A(DP_OP_424J2_126_3477_n2680), .B(
        DP_OP_424J2_126_3477_n2511), .CI(DP_OP_424J2_126_3477_n2518), .CO(
        DP_OP_424J2_126_3477_n1288), .S(DP_OP_424J2_126_3477_n1289) );
  FADDX1_HVT DP_OP_424J2_126_3477_U801 ( .A(DP_OP_424J2_126_3477_n2650), .B(
        DP_OP_424J2_126_3477_n2643), .CI(DP_OP_424J2_126_3477_n2636), .CO(
        DP_OP_424J2_126_3477_n1286), .S(DP_OP_424J2_126_3477_n1287) );
  FADDX1_HVT DP_OP_424J2_126_3477_U800 ( .A(DP_OP_424J2_126_3477_n2592), .B(
        DP_OP_424J2_126_3477_n2606), .CI(DP_OP_424J2_126_3477_n2548), .CO(
        DP_OP_424J2_126_3477_n1284), .S(DP_OP_424J2_126_3477_n1285) );
  FADDX1_HVT DP_OP_424J2_126_3477_U799 ( .A(DP_OP_424J2_126_3477_n2555), .B(
        DP_OP_424J2_126_3477_n2562), .CI(DP_OP_424J2_126_3477_n2599), .CO(
        DP_OP_424J2_126_3477_n1282), .S(DP_OP_424J2_126_3477_n1283) );
  FADDX1_HVT DP_OP_424J2_126_3477_U798 ( .A(DP_OP_424J2_126_3477_n1349), .B(
        DP_OP_424J2_126_3477_n1524), .CI(DP_OP_424J2_126_3477_n1514), .CO(
        DP_OP_424J2_126_3477_n1280), .S(DP_OP_424J2_126_3477_n1281) );
  FADDX1_HVT DP_OP_424J2_126_3477_U797 ( .A(DP_OP_424J2_126_3477_n1522), .B(
        DP_OP_424J2_126_3477_n1520), .CI(DP_OP_424J2_126_3477_n1518), .CO(
        DP_OP_424J2_126_3477_n1278), .S(DP_OP_424J2_126_3477_n1279) );
  FADDX1_HVT DP_OP_424J2_126_3477_U796 ( .A(DP_OP_424J2_126_3477_n1516), .B(
        DP_OP_424J2_126_3477_n1512), .CI(DP_OP_424J2_126_3477_n1508), .CO(
        DP_OP_424J2_126_3477_n1276), .S(DP_OP_424J2_126_3477_n1277) );
  FADDX1_HVT DP_OP_424J2_126_3477_U795 ( .A(DP_OP_424J2_126_3477_n1510), .B(
        DP_OP_424J2_126_3477_n1484), .CI(DP_OP_424J2_126_3477_n1482), .CO(
        DP_OP_424J2_126_3477_n1274), .S(DP_OP_424J2_126_3477_n1275) );
  FADDX1_HVT DP_OP_424J2_126_3477_U794 ( .A(DP_OP_424J2_126_3477_n1486), .B(
        DP_OP_424J2_126_3477_n1458), .CI(DP_OP_424J2_126_3477_n1506), .CO(
        DP_OP_424J2_126_3477_n1272), .S(DP_OP_424J2_126_3477_n1273) );
  FADDX1_HVT DP_OP_424J2_126_3477_U793 ( .A(DP_OP_424J2_126_3477_n1478), .B(
        DP_OP_424J2_126_3477_n1504), .CI(DP_OP_424J2_126_3477_n1502), .CO(
        DP_OP_424J2_126_3477_n1270), .S(DP_OP_424J2_126_3477_n1271) );
  FADDX1_HVT DP_OP_424J2_126_3477_U792 ( .A(DP_OP_424J2_126_3477_n1474), .B(
        DP_OP_424J2_126_3477_n1500), .CI(DP_OP_424J2_126_3477_n1498), .CO(
        DP_OP_424J2_126_3477_n1268), .S(DP_OP_424J2_126_3477_n1269) );
  FADDX1_HVT DP_OP_424J2_126_3477_U791 ( .A(DP_OP_424J2_126_3477_n1468), .B(
        DP_OP_424J2_126_3477_n1460), .CI(DP_OP_424J2_126_3477_n1462), .CO(
        DP_OP_424J2_126_3477_n1266), .S(DP_OP_424J2_126_3477_n1267) );
  FADDX1_HVT DP_OP_424J2_126_3477_U790 ( .A(DP_OP_424J2_126_3477_n1466), .B(
        DP_OP_424J2_126_3477_n1496), .CI(DP_OP_424J2_126_3477_n1494), .CO(
        DP_OP_424J2_126_3477_n1264), .S(DP_OP_424J2_126_3477_n1265) );
  FADDX1_HVT DP_OP_424J2_126_3477_U789 ( .A(DP_OP_424J2_126_3477_n1476), .B(
        DP_OP_424J2_126_3477_n1492), .CI(DP_OP_424J2_126_3477_n1464), .CO(
        DP_OP_424J2_126_3477_n1262), .S(DP_OP_424J2_126_3477_n1263) );
  FADDX1_HVT DP_OP_424J2_126_3477_U788 ( .A(DP_OP_424J2_126_3477_n1472), .B(
        DP_OP_424J2_126_3477_n1490), .CI(DP_OP_424J2_126_3477_n1488), .CO(
        DP_OP_424J2_126_3477_n1260), .S(DP_OP_424J2_126_3477_n1261) );
  FADDX1_HVT DP_OP_424J2_126_3477_U787 ( .A(DP_OP_424J2_126_3477_n1470), .B(
        DP_OP_424J2_126_3477_n1480), .CI(DP_OP_424J2_126_3477_n1339), .CO(
        DP_OP_424J2_126_3477_n1258), .S(DP_OP_424J2_126_3477_n1259) );
  FADDX1_HVT DP_OP_424J2_126_3477_U786 ( .A(DP_OP_424J2_126_3477_n1341), .B(
        DP_OP_424J2_126_3477_n1333), .CI(DP_OP_424J2_126_3477_n1335), .CO(
        DP_OP_424J2_126_3477_n1256), .S(DP_OP_424J2_126_3477_n1257) );
  FADDX1_HVT DP_OP_424J2_126_3477_U785 ( .A(DP_OP_424J2_126_3477_n1345), .B(
        DP_OP_424J2_126_3477_n1343), .CI(DP_OP_424J2_126_3477_n1347), .CO(
        DP_OP_424J2_126_3477_n1254), .S(DP_OP_424J2_126_3477_n1255) );
  FADDX1_HVT DP_OP_424J2_126_3477_U784 ( .A(DP_OP_424J2_126_3477_n1337), .B(
        DP_OP_424J2_126_3477_n1289), .CI(DP_OP_424J2_126_3477_n1287), .CO(
        DP_OP_424J2_126_3477_n1252), .S(DP_OP_424J2_126_3477_n1253) );
  FADDX1_HVT DP_OP_424J2_126_3477_U783 ( .A(DP_OP_424J2_126_3477_n1283), .B(
        DP_OP_424J2_126_3477_n1331), .CI(DP_OP_424J2_126_3477_n1329), .CO(
        DP_OP_424J2_126_3477_n1250), .S(DP_OP_424J2_126_3477_n1251) );
  FADDX1_HVT DP_OP_424J2_126_3477_U782 ( .A(DP_OP_424J2_126_3477_n1319), .B(
        DP_OP_424J2_126_3477_n1309), .CI(DP_OP_424J2_126_3477_n1315), .CO(
        DP_OP_424J2_126_3477_n1248), .S(DP_OP_424J2_126_3477_n1249) );
  FADDX1_HVT DP_OP_424J2_126_3477_U781 ( .A(DP_OP_424J2_126_3477_n1313), .B(
        DP_OP_424J2_126_3477_n1311), .CI(DP_OP_424J2_126_3477_n1295), .CO(
        DP_OP_424J2_126_3477_n1246), .S(DP_OP_424J2_126_3477_n1247) );
  FADDX1_HVT DP_OP_424J2_126_3477_U780 ( .A(DP_OP_424J2_126_3477_n1317), .B(
        DP_OP_424J2_126_3477_n1291), .CI(DP_OP_424J2_126_3477_n1285), .CO(
        DP_OP_424J2_126_3477_n1244), .S(DP_OP_424J2_126_3477_n1245) );
  FADDX1_HVT DP_OP_424J2_126_3477_U779 ( .A(DP_OP_424J2_126_3477_n1321), .B(
        DP_OP_424J2_126_3477_n1303), .CI(DP_OP_424J2_126_3477_n1305), .CO(
        DP_OP_424J2_126_3477_n1242), .S(DP_OP_424J2_126_3477_n1243) );
  FADDX1_HVT DP_OP_424J2_126_3477_U778 ( .A(DP_OP_424J2_126_3477_n1301), .B(
        DP_OP_424J2_126_3477_n1299), .CI(DP_OP_424J2_126_3477_n1293), .CO(
        DP_OP_424J2_126_3477_n1240), .S(DP_OP_424J2_126_3477_n1241) );
  FADDX1_HVT DP_OP_424J2_126_3477_U777 ( .A(DP_OP_424J2_126_3477_n1297), .B(
        DP_OP_424J2_126_3477_n1327), .CI(DP_OP_424J2_126_3477_n1323), .CO(
        DP_OP_424J2_126_3477_n1238), .S(DP_OP_424J2_126_3477_n1239) );
  FADDX1_HVT DP_OP_424J2_126_3477_U776 ( .A(DP_OP_424J2_126_3477_n1325), .B(
        DP_OP_424J2_126_3477_n1307), .CI(DP_OP_424J2_126_3477_n1456), .CO(
        DP_OP_424J2_126_3477_n1236), .S(DP_OP_424J2_126_3477_n1237) );
  FADDX1_HVT DP_OP_424J2_126_3477_U775 ( .A(DP_OP_424J2_126_3477_n1454), .B(
        DP_OP_424J2_126_3477_n1452), .CI(DP_OP_424J2_126_3477_n1450), .CO(
        DP_OP_424J2_126_3477_n1234), .S(DP_OP_424J2_126_3477_n1235) );
  FADDX1_HVT DP_OP_424J2_126_3477_U774 ( .A(DP_OP_424J2_126_3477_n1448), .B(
        DP_OP_424J2_126_3477_n1436), .CI(DP_OP_424J2_126_3477_n1438), .CO(
        DP_OP_424J2_126_3477_n1232), .S(DP_OP_424J2_126_3477_n1233) );
  FADDX1_HVT DP_OP_424J2_126_3477_U773 ( .A(DP_OP_424J2_126_3477_n1442), .B(
        DP_OP_424J2_126_3477_n1446), .CI(DP_OP_424J2_126_3477_n1440), .CO(
        DP_OP_424J2_126_3477_n1230), .S(DP_OP_424J2_126_3477_n1231) );
  FADDX1_HVT DP_OP_424J2_126_3477_U772 ( .A(DP_OP_424J2_126_3477_n1444), .B(
        DP_OP_424J2_126_3477_n1281), .CI(DP_OP_424J2_126_3477_n1434), .CO(
        DP_OP_424J2_126_3477_n1228), .S(DP_OP_424J2_126_3477_n1229) );
  FADDX1_HVT DP_OP_424J2_126_3477_U771 ( .A(DP_OP_424J2_126_3477_n1279), .B(
        DP_OP_424J2_126_3477_n1277), .CI(DP_OP_424J2_126_3477_n1275), .CO(
        DP_OP_424J2_126_3477_n1226), .S(DP_OP_424J2_126_3477_n1227) );
  FADDX1_HVT DP_OP_424J2_126_3477_U770 ( .A(DP_OP_424J2_126_3477_n1432), .B(
        DP_OP_424J2_126_3477_n1430), .CI(DP_OP_424J2_126_3477_n1428), .CO(
        DP_OP_424J2_126_3477_n1224), .S(DP_OP_424J2_126_3477_n1225) );
  FADDX1_HVT DP_OP_424J2_126_3477_U769 ( .A(DP_OP_424J2_126_3477_n1416), .B(
        DP_OP_424J2_126_3477_n1261), .CI(DP_OP_424J2_126_3477_n1259), .CO(
        DP_OP_424J2_126_3477_n1222), .S(DP_OP_424J2_126_3477_n1223) );
  FADDX1_HVT DP_OP_424J2_126_3477_U768 ( .A(DP_OP_424J2_126_3477_n1426), .B(
        DP_OP_424J2_126_3477_n1271), .CI(DP_OP_424J2_126_3477_n1273), .CO(
        DP_OP_424J2_126_3477_n1220), .S(DP_OP_424J2_126_3477_n1221) );
  FADDX1_HVT DP_OP_424J2_126_3477_U767 ( .A(DP_OP_424J2_126_3477_n1424), .B(
        DP_OP_424J2_126_3477_n1267), .CI(DP_OP_424J2_126_3477_n1263), .CO(
        DP_OP_424J2_126_3477_n1218), .S(DP_OP_424J2_126_3477_n1219) );
  FADDX1_HVT DP_OP_424J2_126_3477_U766 ( .A(DP_OP_424J2_126_3477_n1422), .B(
        DP_OP_424J2_126_3477_n1269), .CI(DP_OP_424J2_126_3477_n1265), .CO(
        DP_OP_424J2_126_3477_n1216), .S(DP_OP_424J2_126_3477_n1217) );
  FADDX1_HVT DP_OP_424J2_126_3477_U765 ( .A(DP_OP_424J2_126_3477_n1420), .B(
        DP_OP_424J2_126_3477_n1414), .CI(DP_OP_424J2_126_3477_n1418), .CO(
        DP_OP_424J2_126_3477_n1214), .S(DP_OP_424J2_126_3477_n1215) );
  FADDX1_HVT DP_OP_424J2_126_3477_U764 ( .A(DP_OP_424J2_126_3477_n1255), .B(
        DP_OP_424J2_126_3477_n1257), .CI(DP_OP_424J2_126_3477_n1253), .CO(
        DP_OP_424J2_126_3477_n1212), .S(DP_OP_424J2_126_3477_n1213) );
  FADDX1_HVT DP_OP_424J2_126_3477_U763 ( .A(DP_OP_424J2_126_3477_n1245), .B(
        DP_OP_424J2_126_3477_n1247), .CI(DP_OP_424J2_126_3477_n1412), .CO(
        DP_OP_424J2_126_3477_n1210), .S(DP_OP_424J2_126_3477_n1211) );
  FADDX1_HVT DP_OP_424J2_126_3477_U762 ( .A(DP_OP_424J2_126_3477_n1243), .B(
        DP_OP_424J2_126_3477_n1251), .CI(DP_OP_424J2_126_3477_n1249), .CO(
        DP_OP_424J2_126_3477_n1208), .S(DP_OP_424J2_126_3477_n1209) );
  FADDX1_HVT DP_OP_424J2_126_3477_U761 ( .A(DP_OP_424J2_126_3477_n1239), .B(
        DP_OP_424J2_126_3477_n1241), .CI(DP_OP_424J2_126_3477_n1408), .CO(
        DP_OP_424J2_126_3477_n1206), .S(DP_OP_424J2_126_3477_n1207) );
  FADDX1_HVT DP_OP_424J2_126_3477_U760 ( .A(DP_OP_424J2_126_3477_n1410), .B(
        DP_OP_424J2_126_3477_n1237), .CI(DP_OP_424J2_126_3477_n1406), .CO(
        DP_OP_424J2_126_3477_n1204), .S(DP_OP_424J2_126_3477_n1205) );
  FADDX1_HVT DP_OP_424J2_126_3477_U759 ( .A(DP_OP_424J2_126_3477_n1404), .B(
        DP_OP_424J2_126_3477_n1402), .CI(DP_OP_424J2_126_3477_n1235), .CO(
        DP_OP_424J2_126_3477_n1202), .S(DP_OP_424J2_126_3477_n1203) );
  FADDX1_HVT DP_OP_424J2_126_3477_U758 ( .A(DP_OP_424J2_126_3477_n1400), .B(
        DP_OP_424J2_126_3477_n1392), .CI(DP_OP_424J2_126_3477_n1229), .CO(
        DP_OP_424J2_126_3477_n1200), .S(DP_OP_424J2_126_3477_n1201) );
  FADDX1_HVT DP_OP_424J2_126_3477_U757 ( .A(DP_OP_424J2_126_3477_n1398), .B(
        DP_OP_424J2_126_3477_n1231), .CI(DP_OP_424J2_126_3477_n1233), .CO(
        DP_OP_424J2_126_3477_n1198), .S(DP_OP_424J2_126_3477_n1199) );
  FADDX1_HVT DP_OP_424J2_126_3477_U756 ( .A(DP_OP_424J2_126_3477_n1396), .B(
        DP_OP_424J2_126_3477_n1394), .CI(DP_OP_424J2_126_3477_n1390), .CO(
        DP_OP_424J2_126_3477_n1196), .S(DP_OP_424J2_126_3477_n1197) );
  FADDX1_HVT DP_OP_424J2_126_3477_U755 ( .A(DP_OP_424J2_126_3477_n1225), .B(
        DP_OP_424J2_126_3477_n1227), .CI(DP_OP_424J2_126_3477_n1388), .CO(
        DP_OP_424J2_126_3477_n1194), .S(DP_OP_424J2_126_3477_n1195) );
  FADDX1_HVT DP_OP_424J2_126_3477_U754 ( .A(DP_OP_424J2_126_3477_n1386), .B(
        DP_OP_424J2_126_3477_n1219), .CI(DP_OP_424J2_126_3477_n1384), .CO(
        DP_OP_424J2_126_3477_n1192), .S(DP_OP_424J2_126_3477_n1193) );
  FADDX1_HVT DP_OP_424J2_126_3477_U753 ( .A(DP_OP_424J2_126_3477_n1217), .B(
        DP_OP_424J2_126_3477_n1223), .CI(DP_OP_424J2_126_3477_n1221), .CO(
        DP_OP_424J2_126_3477_n1190), .S(DP_OP_424J2_126_3477_n1191) );
  FADDX1_HVT DP_OP_424J2_126_3477_U752 ( .A(DP_OP_424J2_126_3477_n1215), .B(
        DP_OP_424J2_126_3477_n1213), .CI(DP_OP_424J2_126_3477_n1209), .CO(
        DP_OP_424J2_126_3477_n1188), .S(DP_OP_424J2_126_3477_n1189) );
  FADDX1_HVT DP_OP_424J2_126_3477_U751 ( .A(DP_OP_424J2_126_3477_n1211), .B(
        DP_OP_424J2_126_3477_n1382), .CI(DP_OP_424J2_126_3477_n1207), .CO(
        DP_OP_424J2_126_3477_n1186), .S(DP_OP_424J2_126_3477_n1187) );
  FADDX1_HVT DP_OP_424J2_126_3477_U750 ( .A(DP_OP_424J2_126_3477_n1380), .B(
        DP_OP_424J2_126_3477_n1378), .CI(DP_OP_424J2_126_3477_n1205), .CO(
        DP_OP_424J2_126_3477_n1184), .S(DP_OP_424J2_126_3477_n1185) );
  FADDX1_HVT DP_OP_424J2_126_3477_U749 ( .A(DP_OP_424J2_126_3477_n1376), .B(
        DP_OP_424J2_126_3477_n1374), .CI(DP_OP_424J2_126_3477_n1203), .CO(
        DP_OP_424J2_126_3477_n1182), .S(DP_OP_424J2_126_3477_n1183) );
  FADDX1_HVT DP_OP_424J2_126_3477_U748 ( .A(DP_OP_424J2_126_3477_n1372), .B(
        DP_OP_424J2_126_3477_n1199), .CI(DP_OP_424J2_126_3477_n1197), .CO(
        DP_OP_424J2_126_3477_n1180), .S(DP_OP_424J2_126_3477_n1181) );
  FADDX1_HVT DP_OP_424J2_126_3477_U747 ( .A(DP_OP_424J2_126_3477_n1370), .B(
        DP_OP_424J2_126_3477_n1201), .CI(DP_OP_424J2_126_3477_n1195), .CO(
        DP_OP_424J2_126_3477_n1178), .S(DP_OP_424J2_126_3477_n1179) );
  FADDX1_HVT DP_OP_424J2_126_3477_U746 ( .A(DP_OP_424J2_126_3477_n1368), .B(
        DP_OP_424J2_126_3477_n1191), .CI(DP_OP_424J2_126_3477_n1366), .CO(
        DP_OP_424J2_126_3477_n1176), .S(DP_OP_424J2_126_3477_n1177) );
  FADDX1_HVT DP_OP_424J2_126_3477_U745 ( .A(DP_OP_424J2_126_3477_n1193), .B(
        DP_OP_424J2_126_3477_n1189), .CI(DP_OP_424J2_126_3477_n1187), .CO(
        DP_OP_424J2_126_3477_n1174), .S(DP_OP_424J2_126_3477_n1175) );
  FADDX1_HVT DP_OP_424J2_126_3477_U744 ( .A(DP_OP_424J2_126_3477_n1364), .B(
        DP_OP_424J2_126_3477_n1362), .CI(DP_OP_424J2_126_3477_n1185), .CO(
        DP_OP_424J2_126_3477_n1172), .S(DP_OP_424J2_126_3477_n1173) );
  FADDX1_HVT DP_OP_424J2_126_3477_U743 ( .A(DP_OP_424J2_126_3477_n1360), .B(
        DP_OP_424J2_126_3477_n1183), .CI(DP_OP_424J2_126_3477_n1181), .CO(
        DP_OP_424J2_126_3477_n1170), .S(DP_OP_424J2_126_3477_n1171) );
  FADDX1_HVT DP_OP_424J2_126_3477_U742 ( .A(DP_OP_424J2_126_3477_n1179), .B(
        DP_OP_424J2_126_3477_n1358), .CI(DP_OP_424J2_126_3477_n1177), .CO(
        DP_OP_424J2_126_3477_n1168), .S(DP_OP_424J2_126_3477_n1169) );
  FADDX1_HVT DP_OP_424J2_126_3477_U741 ( .A(DP_OP_424J2_126_3477_n1356), .B(
        DP_OP_424J2_126_3477_n1175), .CI(DP_OP_424J2_126_3477_n1354), .CO(
        DP_OP_424J2_126_3477_n1166), .S(DP_OP_424J2_126_3477_n1167) );
  FADDX1_HVT DP_OP_424J2_126_3477_U740 ( .A(DP_OP_424J2_126_3477_n1173), .B(
        DP_OP_424J2_126_3477_n1171), .CI(DP_OP_424J2_126_3477_n1352), .CO(
        DP_OP_424J2_126_3477_n1164), .S(DP_OP_424J2_126_3477_n1165) );
  FADDX1_HVT DP_OP_424J2_126_3477_U739 ( .A(DP_OP_424J2_126_3477_n1169), .B(
        DP_OP_424J2_126_3477_n1350), .CI(DP_OP_424J2_126_3477_n1167), .CO(
        DP_OP_424J2_126_3477_n1162), .S(DP_OP_424J2_126_3477_n1163) );
  OR2X1_HVT DP_OP_424J2_126_3477_U738 ( .A1(DP_OP_424J2_126_3477_n2979), .A2(
        DP_OP_424J2_126_3477_n2452), .Y(DP_OP_424J2_126_3477_n1160) );
  FADDX1_HVT DP_OP_424J2_126_3477_U736 ( .A(DP_OP_424J2_126_3477_n2144), .B(
        DP_OP_424J2_126_3477_n1924), .CI(DP_OP_424J2_126_3477_n1880), .CO(
        DP_OP_424J2_126_3477_n1158), .S(DP_OP_424J2_126_3477_n1159) );
  FADDX1_HVT DP_OP_424J2_126_3477_U735 ( .A(DP_OP_424J2_126_3477_n2584), .B(
        DP_OP_424J2_126_3477_n2012), .CI(DP_OP_424J2_126_3477_n2364), .CO(
        DP_OP_424J2_126_3477_n1156), .S(DP_OP_424J2_126_3477_n1157) );
  FADDX1_HVT DP_OP_424J2_126_3477_U734 ( .A(DP_OP_424J2_126_3477_n2804), .B(
        DP_OP_424J2_126_3477_n2628), .CI(DP_OP_424J2_126_3477_n2188), .CO(
        DP_OP_424J2_126_3477_n1154), .S(DP_OP_424J2_126_3477_n1155) );
  FADDX1_HVT DP_OP_424J2_126_3477_U733 ( .A(DP_OP_424J2_126_3477_n2276), .B(
        DP_OP_424J2_126_3477_n2100), .CI(DP_OP_424J2_126_3477_n2848), .CO(
        DP_OP_424J2_126_3477_n1152), .S(DP_OP_424J2_126_3477_n1153) );
  FADDX1_HVT DP_OP_424J2_126_3477_U732 ( .A(DP_OP_424J2_126_3477_n2408), .B(
        DP_OP_424J2_126_3477_n2892), .CI(DP_OP_424J2_126_3477_n2672), .CO(
        DP_OP_424J2_126_3477_n1150), .S(DP_OP_424J2_126_3477_n1151) );
  FADDX1_HVT DP_OP_424J2_126_3477_U731 ( .A(DP_OP_424J2_126_3477_n2496), .B(
        DP_OP_424J2_126_3477_n2716), .CI(DP_OP_424J2_126_3477_n2540), .CO(
        DP_OP_424J2_126_3477_n1148), .S(DP_OP_424J2_126_3477_n1149) );
  FADDX1_HVT DP_OP_424J2_126_3477_U730 ( .A(DP_OP_424J2_126_3477_n2232), .B(
        DP_OP_424J2_126_3477_n2056), .CI(DP_OP_424J2_126_3477_n2936), .CO(
        DP_OP_424J2_126_3477_n1146), .S(DP_OP_424J2_126_3477_n1147) );
  FADDX1_HVT DP_OP_424J2_126_3477_U729 ( .A(DP_OP_424J2_126_3477_n2760), .B(
        DP_OP_424J2_126_3477_n1968), .CI(DP_OP_424J2_126_3477_n2320), .CO(
        DP_OP_424J2_126_3477_n1144), .S(DP_OP_424J2_126_3477_n1145) );
  FADDX1_HVT DP_OP_424J2_126_3477_U728 ( .A(DP_OP_424J2_126_3477_n2371), .B(
        DP_OP_424J2_126_3477_n2999), .CI(DP_OP_424J2_126_3477_n1931), .CO(
        DP_OP_424J2_126_3477_n1142), .S(DP_OP_424J2_126_3477_n1143) );
  FADDX1_HVT DP_OP_424J2_126_3477_U727 ( .A(DP_OP_424J2_126_3477_n2378), .B(
        DP_OP_424J2_126_3477_n2992), .CI(DP_OP_424J2_126_3477_n2985), .CO(
        DP_OP_424J2_126_3477_n1140), .S(DP_OP_424J2_126_3477_n1141) );
  FADDX1_HVT DP_OP_424J2_126_3477_U726 ( .A(DP_OP_424J2_126_3477_n2334), .B(
        DP_OP_424J2_126_3477_n2957), .CI(DP_OP_424J2_126_3477_n2950), .CO(
        DP_OP_424J2_126_3477_n1138), .S(DP_OP_424J2_126_3477_n1139) );
  FADDX1_HVT DP_OP_424J2_126_3477_U725 ( .A(DP_OP_424J2_126_3477_n2297), .B(
        DP_OP_424J2_126_3477_n2943), .CI(DP_OP_424J2_126_3477_n2913), .CO(
        DP_OP_424J2_126_3477_n1136), .S(DP_OP_424J2_126_3477_n1137) );
  FADDX1_HVT DP_OP_424J2_126_3477_U724 ( .A(DP_OP_424J2_126_3477_n2290), .B(
        DP_OP_424J2_126_3477_n1938), .CI(DP_OP_424J2_126_3477_n2906), .CO(
        DP_OP_424J2_126_3477_n1134), .S(DP_OP_424J2_126_3477_n1135) );
  FADDX1_HVT DP_OP_424J2_126_3477_U723 ( .A(DP_OP_424J2_126_3477_n2327), .B(
        DP_OP_424J2_126_3477_n2899), .CI(DP_OP_424J2_126_3477_n1945), .CO(
        DP_OP_424J2_126_3477_n1132), .S(DP_OP_424J2_126_3477_n1133) );
  FADDX1_HVT DP_OP_424J2_126_3477_U722 ( .A(DP_OP_424J2_126_3477_n2283), .B(
        DP_OP_424J2_126_3477_n2869), .CI(DP_OP_424J2_126_3477_n1975), .CO(
        DP_OP_424J2_126_3477_n1130), .S(DP_OP_424J2_126_3477_n1131) );
  FADDX1_HVT DP_OP_424J2_126_3477_U721 ( .A(DP_OP_424J2_126_3477_n2253), .B(
        DP_OP_424J2_126_3477_n2862), .CI(DP_OP_424J2_126_3477_n2855), .CO(
        DP_OP_424J2_126_3477_n1128), .S(DP_OP_424J2_126_3477_n1129) );
  FADDX1_HVT DP_OP_424J2_126_3477_U720 ( .A(DP_OP_424J2_126_3477_n2246), .B(
        DP_OP_424J2_126_3477_n1982), .CI(DP_OP_424J2_126_3477_n2825), .CO(
        DP_OP_424J2_126_3477_n1126), .S(DP_OP_424J2_126_3477_n1127) );
  FADDX1_HVT DP_OP_424J2_126_3477_U719 ( .A(DP_OP_424J2_126_3477_n2239), .B(
        DP_OP_424J2_126_3477_n1989), .CI(DP_OP_424J2_126_3477_n2818), .CO(
        DP_OP_424J2_126_3477_n1124), .S(DP_OP_424J2_126_3477_n1125) );
  FADDX1_HVT DP_OP_424J2_126_3477_U718 ( .A(DP_OP_424J2_126_3477_n2019), .B(
        DP_OP_424J2_126_3477_n2026), .CI(DP_OP_424J2_126_3477_n2033), .CO(
        DP_OP_424J2_126_3477_n1122), .S(DP_OP_424J2_126_3477_n1123) );
  FADDX1_HVT DP_OP_424J2_126_3477_U717 ( .A(DP_OP_424J2_126_3477_n2811), .B(
        DP_OP_424J2_126_3477_n2063), .CI(DP_OP_424J2_126_3477_n2070), .CO(
        DP_OP_424J2_126_3477_n1120), .S(DP_OP_424J2_126_3477_n1121) );
  FADDX1_HVT DP_OP_424J2_126_3477_U716 ( .A(DP_OP_424J2_126_3477_n2781), .B(
        DP_OP_424J2_126_3477_n2077), .CI(DP_OP_424J2_126_3477_n2107), .CO(
        DP_OP_424J2_126_3477_n1118), .S(DP_OP_424J2_126_3477_n1119) );
  FADDX1_HVT DP_OP_424J2_126_3477_U715 ( .A(DP_OP_424J2_126_3477_n2774), .B(
        DP_OP_424J2_126_3477_n2114), .CI(DP_OP_424J2_126_3477_n2121), .CO(
        DP_OP_424J2_126_3477_n1116), .S(DP_OP_424J2_126_3477_n1117) );
  FADDX1_HVT DP_OP_424J2_126_3477_U714 ( .A(DP_OP_424J2_126_3477_n2767), .B(
        DP_OP_424J2_126_3477_n2151), .CI(DP_OP_424J2_126_3477_n2158), .CO(
        DP_OP_424J2_126_3477_n1114), .S(DP_OP_424J2_126_3477_n1115) );
  FADDX1_HVT DP_OP_424J2_126_3477_U713 ( .A(DP_OP_424J2_126_3477_n2737), .B(
        DP_OP_424J2_126_3477_n2165), .CI(DP_OP_424J2_126_3477_n2195), .CO(
        DP_OP_424J2_126_3477_n1112), .S(DP_OP_424J2_126_3477_n1113) );
  FADDX1_HVT DP_OP_424J2_126_3477_U712 ( .A(DP_OP_424J2_126_3477_n2730), .B(
        DP_OP_424J2_126_3477_n2202), .CI(DP_OP_424J2_126_3477_n2209), .CO(
        DP_OP_424J2_126_3477_n1110), .S(DP_OP_424J2_126_3477_n1111) );
  FADDX1_HVT DP_OP_424J2_126_3477_U711 ( .A(DP_OP_424J2_126_3477_n2723), .B(
        DP_OP_424J2_126_3477_n2341), .CI(DP_OP_424J2_126_3477_n2385), .CO(
        DP_OP_424J2_126_3477_n1108), .S(DP_OP_424J2_126_3477_n1109) );
  FADDX1_HVT DP_OP_424J2_126_3477_U710 ( .A(DP_OP_424J2_126_3477_n2693), .B(
        DP_OP_424J2_126_3477_n2415), .CI(DP_OP_424J2_126_3477_n2422), .CO(
        DP_OP_424J2_126_3477_n1106), .S(DP_OP_424J2_126_3477_n1107) );
  FADDX1_HVT DP_OP_424J2_126_3477_U709 ( .A(DP_OP_424J2_126_3477_n2686), .B(
        DP_OP_424J2_126_3477_n2429), .CI(DP_OP_424J2_126_3477_n2459), .CO(
        DP_OP_424J2_126_3477_n1104), .S(DP_OP_424J2_126_3477_n1105) );
  FADDX1_HVT DP_OP_424J2_126_3477_U708 ( .A(DP_OP_424J2_126_3477_n2679), .B(
        DP_OP_424J2_126_3477_n2466), .CI(DP_OP_424J2_126_3477_n2473), .CO(
        DP_OP_424J2_126_3477_n1102), .S(DP_OP_424J2_126_3477_n1103) );
  FADDX1_HVT DP_OP_424J2_126_3477_U707 ( .A(DP_OP_424J2_126_3477_n2649), .B(
        DP_OP_424J2_126_3477_n2503), .CI(DP_OP_424J2_126_3477_n2510), .CO(
        DP_OP_424J2_126_3477_n1100), .S(DP_OP_424J2_126_3477_n1101) );
  FADDX1_HVT DP_OP_424J2_126_3477_U706 ( .A(DP_OP_424J2_126_3477_n2642), .B(
        DP_OP_424J2_126_3477_n2517), .CI(DP_OP_424J2_126_3477_n2547), .CO(
        DP_OP_424J2_126_3477_n1098), .S(DP_OP_424J2_126_3477_n1099) );
  FADDX1_HVT DP_OP_424J2_126_3477_U705 ( .A(DP_OP_424J2_126_3477_n2635), .B(
        DP_OP_424J2_126_3477_n2554), .CI(DP_OP_424J2_126_3477_n2561), .CO(
        DP_OP_424J2_126_3477_n1096), .S(DP_OP_424J2_126_3477_n1097) );
  FADDX1_HVT DP_OP_424J2_126_3477_U704 ( .A(DP_OP_424J2_126_3477_n2591), .B(
        DP_OP_424J2_126_3477_n2598), .CI(DP_OP_424J2_126_3477_n2605), .CO(
        DP_OP_424J2_126_3477_n1094), .S(DP_OP_424J2_126_3477_n1095) );
  FADDX1_HVT DP_OP_424J2_126_3477_U703 ( .A(DP_OP_424J2_126_3477_n1348), .B(
        DP_OP_424J2_126_3477_n1336), .CI(DP_OP_424J2_126_3477_n1334), .CO(
        DP_OP_424J2_126_3477_n1092), .S(DP_OP_424J2_126_3477_n1093) );
  FADDX1_HVT DP_OP_424J2_126_3477_U702 ( .A(DP_OP_424J2_126_3477_n1332), .B(
        DP_OP_424J2_126_3477_n1338), .CI(DP_OP_424J2_126_3477_n1161), .CO(
        DP_OP_424J2_126_3477_n1090), .S(DP_OP_424J2_126_3477_n1091) );
  FADDX1_HVT DP_OP_424J2_126_3477_U701 ( .A(DP_OP_424J2_126_3477_n1342), .B(
        DP_OP_424J2_126_3477_n1346), .CI(DP_OP_424J2_126_3477_n1340), .CO(
        DP_OP_424J2_126_3477_n1088), .S(DP_OP_424J2_126_3477_n1089) );
  FADDX1_HVT DP_OP_424J2_126_3477_U700 ( .A(DP_OP_424J2_126_3477_n1344), .B(
        DP_OP_424J2_126_3477_n1308), .CI(DP_OP_424J2_126_3477_n1306), .CO(
        DP_OP_424J2_126_3477_n1086), .S(DP_OP_424J2_126_3477_n1087) );
  FADDX1_HVT DP_OP_424J2_126_3477_U699 ( .A(DP_OP_424J2_126_3477_n1310), .B(
        DP_OP_424J2_126_3477_n1282), .CI(DP_OP_424J2_126_3477_n1330), .CO(
        DP_OP_424J2_126_3477_n1084), .S(DP_OP_424J2_126_3477_n1085) );
  FADDX1_HVT DP_OP_424J2_126_3477_U698 ( .A(DP_OP_424J2_126_3477_n1302), .B(
        DP_OP_424J2_126_3477_n1284), .CI(DP_OP_424J2_126_3477_n1328), .CO(
        DP_OP_424J2_126_3477_n1082), .S(DP_OP_424J2_126_3477_n1083) );
  FADDX1_HVT DP_OP_424J2_126_3477_U697 ( .A(DP_OP_424J2_126_3477_n1300), .B(
        DP_OP_424J2_126_3477_n1286), .CI(DP_OP_424J2_126_3477_n1326), .CO(
        DP_OP_424J2_126_3477_n1080), .S(DP_OP_424J2_126_3477_n1081) );
  FADDX1_HVT DP_OP_424J2_126_3477_U696 ( .A(DP_OP_424J2_126_3477_n1296), .B(
        DP_OP_424J2_126_3477_n1324), .CI(DP_OP_424J2_126_3477_n1322), .CO(
        DP_OP_424J2_126_3477_n1078), .S(DP_OP_424J2_126_3477_n1079) );
  FADDX1_HVT DP_OP_424J2_126_3477_U695 ( .A(DP_OP_424J2_126_3477_n1290), .B(
        DP_OP_424J2_126_3477_n1320), .CI(DP_OP_424J2_126_3477_n1318), .CO(
        DP_OP_424J2_126_3477_n1076), .S(DP_OP_424J2_126_3477_n1077) );
  FADDX1_HVT DP_OP_424J2_126_3477_U694 ( .A(DP_OP_424J2_126_3477_n1298), .B(
        DP_OP_424J2_126_3477_n1316), .CI(DP_OP_424J2_126_3477_n1314), .CO(
        DP_OP_424J2_126_3477_n1074), .S(DP_OP_424J2_126_3477_n1075) );
  FADDX1_HVT DP_OP_424J2_126_3477_U693 ( .A(DP_OP_424J2_126_3477_n1292), .B(
        DP_OP_424J2_126_3477_n1312), .CI(DP_OP_424J2_126_3477_n1304), .CO(
        DP_OP_424J2_126_3477_n1072), .S(DP_OP_424J2_126_3477_n1073) );
  FADDX1_HVT DP_OP_424J2_126_3477_U692 ( .A(DP_OP_424J2_126_3477_n1294), .B(
        DP_OP_424J2_126_3477_n1288), .CI(DP_OP_424J2_126_3477_n1151), .CO(
        DP_OP_424J2_126_3477_n1070), .S(DP_OP_424J2_126_3477_n1071) );
  FADDX1_HVT DP_OP_424J2_126_3477_U691 ( .A(DP_OP_424J2_126_3477_n1147), .B(
        DP_OP_424J2_126_3477_n1145), .CI(DP_OP_424J2_126_3477_n1149), .CO(
        DP_OP_424J2_126_3477_n1068), .S(DP_OP_424J2_126_3477_n1069) );
  FADDX1_HVT DP_OP_424J2_126_3477_U690 ( .A(DP_OP_424J2_126_3477_n1157), .B(
        DP_OP_424J2_126_3477_n1155), .CI(DP_OP_424J2_126_3477_n1159), .CO(
        DP_OP_424J2_126_3477_n1066), .S(DP_OP_424J2_126_3477_n1067) );
  FADDX1_HVT DP_OP_424J2_126_3477_U689 ( .A(DP_OP_424J2_126_3477_n1153), .B(
        DP_OP_424J2_126_3477_n1101), .CI(DP_OP_424J2_126_3477_n1103), .CO(
        DP_OP_424J2_126_3477_n1064), .S(DP_OP_424J2_126_3477_n1065) );
  FADDX1_HVT DP_OP_424J2_126_3477_U688 ( .A(DP_OP_424J2_126_3477_n1099), .B(
        DP_OP_424J2_126_3477_n1135), .CI(DP_OP_424J2_126_3477_n1131), .CO(
        DP_OP_424J2_126_3477_n1062), .S(DP_OP_424J2_126_3477_n1063) );
  FADDX1_HVT DP_OP_424J2_126_3477_U687 ( .A(DP_OP_424J2_126_3477_n1137), .B(
        DP_OP_424J2_126_3477_n1121), .CI(DP_OP_424J2_126_3477_n1127), .CO(
        DP_OP_424J2_126_3477_n1060), .S(DP_OP_424J2_126_3477_n1061) );
  FADDX1_HVT DP_OP_424J2_126_3477_U686 ( .A(DP_OP_424J2_126_3477_n1125), .B(
        DP_OP_424J2_126_3477_n1123), .CI(DP_OP_424J2_126_3477_n1107), .CO(
        DP_OP_424J2_126_3477_n1058), .S(DP_OP_424J2_126_3477_n1059) );
  FADDX1_HVT DP_OP_424J2_126_3477_U685 ( .A(DP_OP_424J2_126_3477_n1129), .B(
        DP_OP_424J2_126_3477_n1097), .CI(DP_OP_424J2_126_3477_n1095), .CO(
        DP_OP_424J2_126_3477_n1056), .S(DP_OP_424J2_126_3477_n1057) );
  FADDX1_HVT DP_OP_424J2_126_3477_U684 ( .A(DP_OP_424J2_126_3477_n1133), .B(
        DP_OP_424J2_126_3477_n1115), .CI(DP_OP_424J2_126_3477_n1117), .CO(
        DP_OP_424J2_126_3477_n1054), .S(DP_OP_424J2_126_3477_n1055) );
  FADDX1_HVT DP_OP_424J2_126_3477_U683 ( .A(DP_OP_424J2_126_3477_n1113), .B(
        DP_OP_424J2_126_3477_n1111), .CI(DP_OP_424J2_126_3477_n1105), .CO(
        DP_OP_424J2_126_3477_n1052), .S(DP_OP_424J2_126_3477_n1053) );
  FADDX1_HVT DP_OP_424J2_126_3477_U682 ( .A(DP_OP_424J2_126_3477_n1109), .B(
        DP_OP_424J2_126_3477_n1143), .CI(DP_OP_424J2_126_3477_n1141), .CO(
        DP_OP_424J2_126_3477_n1050), .S(DP_OP_424J2_126_3477_n1051) );
  FADDX1_HVT DP_OP_424J2_126_3477_U681 ( .A(DP_OP_424J2_126_3477_n1139), .B(
        DP_OP_424J2_126_3477_n1119), .CI(DP_OP_424J2_126_3477_n1280), .CO(
        DP_OP_424J2_126_3477_n1048), .S(DP_OP_424J2_126_3477_n1049) );
  FADDX1_HVT DP_OP_424J2_126_3477_U680 ( .A(DP_OP_424J2_126_3477_n1278), .B(
        DP_OP_424J2_126_3477_n1276), .CI(DP_OP_424J2_126_3477_n1274), .CO(
        DP_OP_424J2_126_3477_n1046), .S(DP_OP_424J2_126_3477_n1047) );
  FADDX1_HVT DP_OP_424J2_126_3477_U679 ( .A(DP_OP_424J2_126_3477_n1272), .B(
        DP_OP_424J2_126_3477_n1260), .CI(DP_OP_424J2_126_3477_n1258), .CO(
        DP_OP_424J2_126_3477_n1044), .S(DP_OP_424J2_126_3477_n1045) );
  FADDX1_HVT DP_OP_424J2_126_3477_U678 ( .A(DP_OP_424J2_126_3477_n1264), .B(
        DP_OP_424J2_126_3477_n1262), .CI(DP_OP_424J2_126_3477_n1270), .CO(
        DP_OP_424J2_126_3477_n1042), .S(DP_OP_424J2_126_3477_n1043) );
  FADDX1_HVT DP_OP_424J2_126_3477_U677 ( .A(DP_OP_424J2_126_3477_n1268), .B(
        DP_OP_424J2_126_3477_n1266), .CI(DP_OP_424J2_126_3477_n1093), .CO(
        DP_OP_424J2_126_3477_n1040), .S(DP_OP_424J2_126_3477_n1041) );
  FADDX1_HVT DP_OP_424J2_126_3477_U676 ( .A(DP_OP_424J2_126_3477_n1256), .B(
        DP_OP_424J2_126_3477_n1254), .CI(DP_OP_424J2_126_3477_n1087), .CO(
        DP_OP_424J2_126_3477_n1038), .S(DP_OP_424J2_126_3477_n1039) );
  FADDX1_HVT DP_OP_424J2_126_3477_U675 ( .A(DP_OP_424J2_126_3477_n1091), .B(
        DP_OP_424J2_126_3477_n1089), .CI(DP_OP_424J2_126_3477_n1252), .CO(
        DP_OP_424J2_126_3477_n1036), .S(DP_OP_424J2_126_3477_n1037) );
  FADDX1_HVT DP_OP_424J2_126_3477_U674 ( .A(DP_OP_424J2_126_3477_n1240), .B(
        DP_OP_424J2_126_3477_n1085), .CI(DP_OP_424J2_126_3477_n1071), .CO(
        DP_OP_424J2_126_3477_n1034), .S(DP_OP_424J2_126_3477_n1035) );
  FADDX1_HVT DP_OP_424J2_126_3477_U673 ( .A(DP_OP_424J2_126_3477_n1238), .B(
        DP_OP_424J2_126_3477_n1081), .CI(DP_OP_424J2_126_3477_n1083), .CO(
        DP_OP_424J2_126_3477_n1032), .S(DP_OP_424J2_126_3477_n1033) );
  FADDX1_HVT DP_OP_424J2_126_3477_U672 ( .A(DP_OP_424J2_126_3477_n1242), .B(
        DP_OP_424J2_126_3477_n1079), .CI(DP_OP_424J2_126_3477_n1077), .CO(
        DP_OP_424J2_126_3477_n1030), .S(DP_OP_424J2_126_3477_n1031) );
  FADDX1_HVT DP_OP_424J2_126_3477_U671 ( .A(DP_OP_424J2_126_3477_n1250), .B(
        DP_OP_424J2_126_3477_n1073), .CI(DP_OP_424J2_126_3477_n1075), .CO(
        DP_OP_424J2_126_3477_n1028), .S(DP_OP_424J2_126_3477_n1029) );
  FADDX1_HVT DP_OP_424J2_126_3477_U670 ( .A(DP_OP_424J2_126_3477_n1248), .B(
        DP_OP_424J2_126_3477_n1244), .CI(DP_OP_424J2_126_3477_n1246), .CO(
        DP_OP_424J2_126_3477_n1026), .S(DP_OP_424J2_126_3477_n1027) );
  FADDX1_HVT DP_OP_424J2_126_3477_U669 ( .A(DP_OP_424J2_126_3477_n1067), .B(
        DP_OP_424J2_126_3477_n1236), .CI(DP_OP_424J2_126_3477_n1065), .CO(
        DP_OP_424J2_126_3477_n1024), .S(DP_OP_424J2_126_3477_n1025) );
  FADDX1_HVT DP_OP_424J2_126_3477_U668 ( .A(DP_OP_424J2_126_3477_n1069), .B(
        DP_OP_424J2_126_3477_n1059), .CI(DP_OP_424J2_126_3477_n1061), .CO(
        DP_OP_424J2_126_3477_n1022), .S(DP_OP_424J2_126_3477_n1023) );
  FADDX1_HVT DP_OP_424J2_126_3477_U667 ( .A(DP_OP_424J2_126_3477_n1057), .B(
        DP_OP_424J2_126_3477_n1051), .CI(DP_OP_424J2_126_3477_n1234), .CO(
        DP_OP_424J2_126_3477_n1020), .S(DP_OP_424J2_126_3477_n1021) );
  FADDX1_HVT DP_OP_424J2_126_3477_U666 ( .A(DP_OP_424J2_126_3477_n1053), .B(
        DP_OP_424J2_126_3477_n1063), .CI(DP_OP_424J2_126_3477_n1055), .CO(
        DP_OP_424J2_126_3477_n1018), .S(DP_OP_424J2_126_3477_n1019) );
  FADDX1_HVT DP_OP_424J2_126_3477_U665 ( .A(DP_OP_424J2_126_3477_n1049), .B(
        DP_OP_424J2_126_3477_n1232), .CI(DP_OP_424J2_126_3477_n1228), .CO(
        DP_OP_424J2_126_3477_n1016), .S(DP_OP_424J2_126_3477_n1017) );
  FADDX1_HVT DP_OP_424J2_126_3477_U664 ( .A(DP_OP_424J2_126_3477_n1230), .B(
        DP_OP_424J2_126_3477_n1226), .CI(DP_OP_424J2_126_3477_n1224), .CO(
        DP_OP_424J2_126_3477_n1014), .S(DP_OP_424J2_126_3477_n1015) );
  FADDX1_HVT DP_OP_424J2_126_3477_U663 ( .A(DP_OP_424J2_126_3477_n1047), .B(
        DP_OP_424J2_126_3477_n1222), .CI(DP_OP_424J2_126_3477_n1220), .CO(
        DP_OP_424J2_126_3477_n1012), .S(DP_OP_424J2_126_3477_n1013) );
  FADDX1_HVT DP_OP_424J2_126_3477_U662 ( .A(DP_OP_424J2_126_3477_n1218), .B(
        DP_OP_424J2_126_3477_n1043), .CI(DP_OP_424J2_126_3477_n1041), .CO(
        DP_OP_424J2_126_3477_n1010), .S(DP_OP_424J2_126_3477_n1011) );
  FADDX1_HVT DP_OP_424J2_126_3477_U661 ( .A(DP_OP_424J2_126_3477_n1216), .B(
        DP_OP_424J2_126_3477_n1214), .CI(DP_OP_424J2_126_3477_n1045), .CO(
        DP_OP_424J2_126_3477_n1008), .S(DP_OP_424J2_126_3477_n1009) );
  FADDX1_HVT DP_OP_424J2_126_3477_U660 ( .A(DP_OP_424J2_126_3477_n1037), .B(
        DP_OP_424J2_126_3477_n1212), .CI(DP_OP_424J2_126_3477_n1039), .CO(
        DP_OP_424J2_126_3477_n1006), .S(DP_OP_424J2_126_3477_n1007) );
  FADDX1_HVT DP_OP_424J2_126_3477_U659 ( .A(DP_OP_424J2_126_3477_n1031), .B(
        DP_OP_424J2_126_3477_n1035), .CI(DP_OP_424J2_126_3477_n1206), .CO(
        DP_OP_424J2_126_3477_n1004), .S(DP_OP_424J2_126_3477_n1005) );
  FADDX1_HVT DP_OP_424J2_126_3477_U658 ( .A(DP_OP_424J2_126_3477_n1210), .B(
        DP_OP_424J2_126_3477_n1029), .CI(DP_OP_424J2_126_3477_n1033), .CO(
        DP_OP_424J2_126_3477_n1002), .S(DP_OP_424J2_126_3477_n1003) );
  FADDX1_HVT DP_OP_424J2_126_3477_U657 ( .A(DP_OP_424J2_126_3477_n1208), .B(
        DP_OP_424J2_126_3477_n1027), .CI(DP_OP_424J2_126_3477_n1204), .CO(
        DP_OP_424J2_126_3477_n1000), .S(DP_OP_424J2_126_3477_n1001) );
  FADDX1_HVT DP_OP_424J2_126_3477_U656 ( .A(DP_OP_424J2_126_3477_n1025), .B(
        DP_OP_424J2_126_3477_n1023), .CI(DP_OP_424J2_126_3477_n1021), .CO(
        DP_OP_424J2_126_3477_n998), .S(DP_OP_424J2_126_3477_n999) );
  FADDX1_HVT DP_OP_424J2_126_3477_U655 ( .A(DP_OP_424J2_126_3477_n1019), .B(
        DP_OP_424J2_126_3477_n1202), .CI(DP_OP_424J2_126_3477_n1017), .CO(
        DP_OP_424J2_126_3477_n996), .S(DP_OP_424J2_126_3477_n997) );
  FADDX1_HVT DP_OP_424J2_126_3477_U654 ( .A(DP_OP_424J2_126_3477_n1200), .B(
        DP_OP_424J2_126_3477_n1198), .CI(DP_OP_424J2_126_3477_n1196), .CO(
        DP_OP_424J2_126_3477_n994), .S(DP_OP_424J2_126_3477_n995) );
  FADDX1_HVT DP_OP_424J2_126_3477_U653 ( .A(DP_OP_424J2_126_3477_n1015), .B(
        DP_OP_424J2_126_3477_n1194), .CI(DP_OP_424J2_126_3477_n1013), .CO(
        DP_OP_424J2_126_3477_n992), .S(DP_OP_424J2_126_3477_n993) );
  FADDX1_HVT DP_OP_424J2_126_3477_U652 ( .A(DP_OP_424J2_126_3477_n1192), .B(
        DP_OP_424J2_126_3477_n1009), .CI(DP_OP_424J2_126_3477_n1011), .CO(
        DP_OP_424J2_126_3477_n990), .S(DP_OP_424J2_126_3477_n991) );
  FADDX1_HVT DP_OP_424J2_126_3477_U651 ( .A(DP_OP_424J2_126_3477_n1190), .B(
        DP_OP_424J2_126_3477_n1188), .CI(DP_OP_424J2_126_3477_n1007), .CO(
        DP_OP_424J2_126_3477_n988), .S(DP_OP_424J2_126_3477_n989) );
  FADDX1_HVT DP_OP_424J2_126_3477_U650 ( .A(DP_OP_424J2_126_3477_n1186), .B(
        DP_OP_424J2_126_3477_n1003), .CI(DP_OP_424J2_126_3477_n1001), .CO(
        DP_OP_424J2_126_3477_n986), .S(DP_OP_424J2_126_3477_n987) );
  FADDX1_HVT DP_OP_424J2_126_3477_U649 ( .A(DP_OP_424J2_126_3477_n1005), .B(
        DP_OP_424J2_126_3477_n1184), .CI(DP_OP_424J2_126_3477_n999), .CO(
        DP_OP_424J2_126_3477_n984), .S(DP_OP_424J2_126_3477_n985) );
  FADDX1_HVT DP_OP_424J2_126_3477_U648 ( .A(DP_OP_424J2_126_3477_n1182), .B(
        DP_OP_424J2_126_3477_n997), .CI(DP_OP_424J2_126_3477_n1180), .CO(
        DP_OP_424J2_126_3477_n982), .S(DP_OP_424J2_126_3477_n983) );
  FADDX1_HVT DP_OP_424J2_126_3477_U647 ( .A(DP_OP_424J2_126_3477_n995), .B(
        DP_OP_424J2_126_3477_n1178), .CI(DP_OP_424J2_126_3477_n993), .CO(
        DP_OP_424J2_126_3477_n980), .S(DP_OP_424J2_126_3477_n981) );
  FADDX1_HVT DP_OP_424J2_126_3477_U646 ( .A(DP_OP_424J2_126_3477_n1176), .B(
        DP_OP_424J2_126_3477_n991), .CI(DP_OP_424J2_126_3477_n989), .CO(
        DP_OP_424J2_126_3477_n978), .S(DP_OP_424J2_126_3477_n979) );
  FADDX1_HVT DP_OP_424J2_126_3477_U645 ( .A(DP_OP_424J2_126_3477_n1174), .B(
        DP_OP_424J2_126_3477_n987), .CI(DP_OP_424J2_126_3477_n1172), .CO(
        DP_OP_424J2_126_3477_n976), .S(DP_OP_424J2_126_3477_n977) );
  FADDX1_HVT DP_OP_424J2_126_3477_U644 ( .A(DP_OP_424J2_126_3477_n985), .B(
        DP_OP_424J2_126_3477_n1170), .CI(DP_OP_424J2_126_3477_n983), .CO(
        DP_OP_424J2_126_3477_n974), .S(DP_OP_424J2_126_3477_n975) );
  FADDX1_HVT DP_OP_424J2_126_3477_U643 ( .A(DP_OP_424J2_126_3477_n981), .B(
        DP_OP_424J2_126_3477_n1168), .CI(DP_OP_424J2_126_3477_n979), .CO(
        DP_OP_424J2_126_3477_n972), .S(DP_OP_424J2_126_3477_n973) );
  FADDX1_HVT DP_OP_424J2_126_3477_U642 ( .A(DP_OP_424J2_126_3477_n1166), .B(
        DP_OP_424J2_126_3477_n977), .CI(DP_OP_424J2_126_3477_n975), .CO(
        DP_OP_424J2_126_3477_n970), .S(DP_OP_424J2_126_3477_n971) );
  FADDX1_HVT DP_OP_424J2_126_3477_U641 ( .A(DP_OP_424J2_126_3477_n1164), .B(
        DP_OP_424J2_126_3477_n973), .CI(DP_OP_424J2_126_3477_n1162), .CO(
        DP_OP_424J2_126_3477_n968), .S(DP_OP_424J2_126_3477_n969) );
  FADDX1_HVT DP_OP_424J2_126_3477_U640 ( .A(DP_OP_424J2_126_3477_n2978), .B(
        DP_OP_424J2_126_3477_n1923), .CI(DP_OP_424J2_126_3477_n1879), .CO(
        DP_OP_424J2_126_3477_n966), .S(DP_OP_424J2_126_3477_n967) );
  FADDX1_HVT DP_OP_424J2_126_3477_U639 ( .A(DP_OP_424J2_126_3477_n2803), .B(
        DP_OP_424J2_126_3477_n2120), .CI(DP_OP_424J2_126_3477_n2384), .CO(
        DP_OP_424J2_126_3477_n964), .S(DP_OP_424J2_126_3477_n965) );
  FADDX1_HVT DP_OP_424J2_126_3477_U638 ( .A(DP_OP_424J2_126_3477_n2011), .B(
        DP_OP_424J2_126_3477_n2428), .CI(DP_OP_424J2_126_3477_n1988), .CO(
        DP_OP_424J2_126_3477_n962), .S(DP_OP_424J2_126_3477_n963) );
  FADDX1_HVT DP_OP_424J2_126_3477_U637 ( .A(DP_OP_424J2_126_3477_n2319), .B(
        DP_OP_424J2_126_3477_n1944), .CI(DP_OP_424J2_126_3477_n2912), .CO(
        DP_OP_424J2_126_3477_n960), .S(DP_OP_424J2_126_3477_n961) );
  FADDX1_HVT DP_OP_424J2_126_3477_U636 ( .A(DP_OP_424J2_126_3477_n2275), .B(
        DP_OP_424J2_126_3477_n2252), .CI(DP_OP_424J2_126_3477_n2604), .CO(
        DP_OP_424J2_126_3477_n958), .S(DP_OP_424J2_126_3477_n959) );
  FADDX1_HVT DP_OP_424J2_126_3477_U635 ( .A(DP_OP_424J2_126_3477_n2187), .B(
        DP_OP_424J2_126_3477_n2296), .CI(DP_OP_424J2_126_3477_n2956), .CO(
        DP_OP_424J2_126_3477_n956), .S(DP_OP_424J2_126_3477_n957) );
  FADDX1_HVT DP_OP_424J2_126_3477_U634 ( .A(DP_OP_424J2_126_3477_n1967), .B(
        DP_OP_424J2_126_3477_n2032), .CI(DP_OP_424J2_126_3477_n2472), .CO(
        DP_OP_424J2_126_3477_n954), .S(DP_OP_424J2_126_3477_n955) );
  FADDX1_HVT DP_OP_424J2_126_3477_U633 ( .A(DP_OP_424J2_126_3477_n2055), .B(
        DP_OP_424J2_126_3477_n2736), .CI(DP_OP_424J2_126_3477_n2780), .CO(
        DP_OP_424J2_126_3477_n952), .S(DP_OP_424J2_126_3477_n953) );
  FADDX1_HVT DP_OP_424J2_126_3477_U632 ( .A(DP_OP_424J2_126_3477_n2143), .B(
        DP_OP_424J2_126_3477_n2692), .CI(DP_OP_424J2_126_3477_n2560), .CO(
        DP_OP_424J2_126_3477_n950), .S(DP_OP_424J2_126_3477_n951) );
  FADDX1_HVT DP_OP_424J2_126_3477_U631 ( .A(DP_OP_424J2_126_3477_n2495), .B(
        DP_OP_424J2_126_3477_n2340), .CI(DP_OP_424J2_126_3477_n2824), .CO(
        DP_OP_424J2_126_3477_n948), .S(DP_OP_424J2_126_3477_n949) );
  FADDX1_HVT DP_OP_424J2_126_3477_U630 ( .A(DP_OP_424J2_126_3477_n2891), .B(
        DP_OP_424J2_126_3477_n2164), .CI(DP_OP_424J2_126_3477_n2076), .CO(
        DP_OP_424J2_126_3477_n946), .S(DP_OP_424J2_126_3477_n947) );
  FADDX1_HVT DP_OP_424J2_126_3477_U629 ( .A(DP_OP_424J2_126_3477_n2627), .B(
        DP_OP_424J2_126_3477_n2868), .CI(DP_OP_424J2_126_3477_n2516), .CO(
        DP_OP_424J2_126_3477_n944), .S(DP_OP_424J2_126_3477_n945) );
  FADDX1_HVT DP_OP_424J2_126_3477_U628 ( .A(DP_OP_424J2_126_3477_n2407), .B(
        DP_OP_424J2_126_3477_n2998), .CI(DP_OP_424J2_126_3477_n2208), .CO(
        DP_OP_424J2_126_3477_n942), .S(DP_OP_424J2_126_3477_n943) );
  FADDX1_HVT DP_OP_424J2_126_3477_U627 ( .A(DP_OP_424J2_126_3477_n2099), .B(
        DP_OP_424J2_126_3477_n2363), .CI(DP_OP_424J2_126_3477_n2648), .CO(
        DP_OP_424J2_126_3477_n940), .S(DP_OP_424J2_126_3477_n941) );
  FADDX1_HVT DP_OP_424J2_126_3477_U626 ( .A(DP_OP_424J2_126_3477_n2715), .B(
        DP_OP_424J2_126_3477_n2759), .CI(DP_OP_424J2_126_3477_n2847), .CO(
        DP_OP_424J2_126_3477_n938), .S(DP_OP_424J2_126_3477_n939) );
  FADDX1_HVT DP_OP_424J2_126_3477_U625 ( .A(DP_OP_424J2_126_3477_n2451), .B(
        DP_OP_424J2_126_3477_n2539), .CI(DP_OP_424J2_126_3477_n2935), .CO(
        DP_OP_424J2_126_3477_n936), .S(DP_OP_424J2_126_3477_n937) );
  FADDX1_HVT DP_OP_424J2_126_3477_U624 ( .A(DP_OP_424J2_126_3477_n2583), .B(
        DP_OP_424J2_126_3477_n2231), .CI(DP_OP_424J2_126_3477_n2671), .CO(
        DP_OP_424J2_126_3477_n934), .S(DP_OP_424J2_126_3477_n935) );
  FADDX1_HVT DP_OP_424J2_126_3477_U623 ( .A(DP_OP_424J2_126_3477_n2991), .B(
        DP_OP_424J2_126_3477_n1937), .CI(DP_OP_424J2_126_3477_n1930), .CO(
        DP_OP_424J2_126_3477_n932), .S(DP_OP_424J2_126_3477_n933) );
  FADDX1_HVT DP_OP_424J2_126_3477_U622 ( .A(DP_OP_424J2_126_3477_n2984), .B(
        DP_OP_424J2_126_3477_n2949), .CI(DP_OP_424J2_126_3477_n2942), .CO(
        DP_OP_424J2_126_3477_n930), .S(DP_OP_424J2_126_3477_n931) );
  FADDX1_HVT DP_OP_424J2_126_3477_U621 ( .A(DP_OP_424J2_126_3477_n2465), .B(
        DP_OP_424J2_126_3477_n2905), .CI(DP_OP_424J2_126_3477_n2898), .CO(
        DP_OP_424J2_126_3477_n928), .S(DP_OP_424J2_126_3477_n929) );
  FADDX1_HVT DP_OP_424J2_126_3477_U620 ( .A(DP_OP_424J2_126_3477_n2861), .B(
        DP_OP_424J2_126_3477_n1974), .CI(DP_OP_424J2_126_3477_n1981), .CO(
        DP_OP_424J2_126_3477_n926), .S(DP_OP_424J2_126_3477_n927) );
  FADDX1_HVT DP_OP_424J2_126_3477_U619 ( .A(DP_OP_424J2_126_3477_n2854), .B(
        DP_OP_424J2_126_3477_n2018), .CI(DP_OP_424J2_126_3477_n2025), .CO(
        DP_OP_424J2_126_3477_n924), .S(DP_OP_424J2_126_3477_n925) );
  FADDX1_HVT DP_OP_424J2_126_3477_U618 ( .A(DP_OP_424J2_126_3477_n2817), .B(
        DP_OP_424J2_126_3477_n2062), .CI(DP_OP_424J2_126_3477_n2069), .CO(
        DP_OP_424J2_126_3477_n922), .S(DP_OP_424J2_126_3477_n923) );
  FADDX1_HVT DP_OP_424J2_126_3477_U617 ( .A(DP_OP_424J2_126_3477_n2810), .B(
        DP_OP_424J2_126_3477_n2106), .CI(DP_OP_424J2_126_3477_n2113), .CO(
        DP_OP_424J2_126_3477_n920), .S(DP_OP_424J2_126_3477_n921) );
  FADDX1_HVT DP_OP_424J2_126_3477_U616 ( .A(DP_OP_424J2_126_3477_n2773), .B(
        DP_OP_424J2_126_3477_n2150), .CI(DP_OP_424J2_126_3477_n2157), .CO(
        DP_OP_424J2_126_3477_n918), .S(DP_OP_424J2_126_3477_n919) );
  FADDX1_HVT DP_OP_424J2_126_3477_U615 ( .A(DP_OP_424J2_126_3477_n2766), .B(
        DP_OP_424J2_126_3477_n2194), .CI(DP_OP_424J2_126_3477_n2201), .CO(
        DP_OP_424J2_126_3477_n916), .S(DP_OP_424J2_126_3477_n917) );
  FADDX1_HVT DP_OP_424J2_126_3477_U614 ( .A(DP_OP_424J2_126_3477_n2729), .B(
        DP_OP_424J2_126_3477_n2238), .CI(DP_OP_424J2_126_3477_n2245), .CO(
        DP_OP_424J2_126_3477_n914), .S(DP_OP_424J2_126_3477_n915) );
  FADDX1_HVT DP_OP_424J2_126_3477_U613 ( .A(DP_OP_424J2_126_3477_n2722), .B(
        DP_OP_424J2_126_3477_n2282), .CI(DP_OP_424J2_126_3477_n2289), .CO(
        DP_OP_424J2_126_3477_n912), .S(DP_OP_424J2_126_3477_n913) );
  FADDX1_HVT DP_OP_424J2_126_3477_U612 ( .A(DP_OP_424J2_126_3477_n2685), .B(
        DP_OP_424J2_126_3477_n2326), .CI(DP_OP_424J2_126_3477_n2333), .CO(
        DP_OP_424J2_126_3477_n910), .S(DP_OP_424J2_126_3477_n911) );
  FADDX1_HVT DP_OP_424J2_126_3477_U611 ( .A(DP_OP_424J2_126_3477_n2678), .B(
        DP_OP_424J2_126_3477_n2370), .CI(DP_OP_424J2_126_3477_n2377), .CO(
        DP_OP_424J2_126_3477_n908), .S(DP_OP_424J2_126_3477_n909) );
  FADDX1_HVT DP_OP_424J2_126_3477_U610 ( .A(DP_OP_424J2_126_3477_n2641), .B(
        DP_OP_424J2_126_3477_n2414), .CI(DP_OP_424J2_126_3477_n2421), .CO(
        DP_OP_424J2_126_3477_n906), .S(DP_OP_424J2_126_3477_n907) );
  FADDX1_HVT DP_OP_424J2_126_3477_U609 ( .A(DP_OP_424J2_126_3477_n2634), .B(
        DP_OP_424J2_126_3477_n2458), .CI(DP_OP_424J2_126_3477_n2502), .CO(
        DP_OP_424J2_126_3477_n904), .S(DP_OP_424J2_126_3477_n905) );
  FADDX1_HVT DP_OP_424J2_126_3477_U608 ( .A(DP_OP_424J2_126_3477_n2597), .B(
        DP_OP_424J2_126_3477_n2509), .CI(DP_OP_424J2_126_3477_n2546), .CO(
        DP_OP_424J2_126_3477_n902), .S(DP_OP_424J2_126_3477_n903) );
  FADDX1_HVT DP_OP_424J2_126_3477_U607 ( .A(DP_OP_424J2_126_3477_n2590), .B(
        DP_OP_424J2_126_3477_n2553), .CI(DP_OP_424J2_126_3477_n1160), .CO(
        DP_OP_424J2_126_3477_n900), .S(DP_OP_424J2_126_3477_n901) );
  FADDX1_HVT DP_OP_424J2_126_3477_U606 ( .A(DP_OP_424J2_126_3477_n1148), .B(
        DP_OP_424J2_126_3477_n1144), .CI(DP_OP_424J2_126_3477_n1158), .CO(
        DP_OP_424J2_126_3477_n898), .S(DP_OP_424J2_126_3477_n899) );
  FADDX1_HVT DP_OP_424J2_126_3477_U605 ( .A(DP_OP_424J2_126_3477_n1156), .B(
        DP_OP_424J2_126_3477_n1146), .CI(DP_OP_424J2_126_3477_n1154), .CO(
        DP_OP_424J2_126_3477_n896), .S(DP_OP_424J2_126_3477_n897) );
  FADDX1_HVT DP_OP_424J2_126_3477_U604 ( .A(DP_OP_424J2_126_3477_n1152), .B(
        DP_OP_424J2_126_3477_n1150), .CI(DP_OP_424J2_126_3477_n1120), .CO(
        DP_OP_424J2_126_3477_n894), .S(DP_OP_424J2_126_3477_n895) );
  FADDX1_HVT DP_OP_424J2_126_3477_U603 ( .A(DP_OP_424J2_126_3477_n1118), .B(
        DP_OP_424J2_126_3477_n1094), .CI(DP_OP_424J2_126_3477_n1142), .CO(
        DP_OP_424J2_126_3477_n892), .S(DP_OP_424J2_126_3477_n893) );
  FADDX1_HVT DP_OP_424J2_126_3477_U602 ( .A(DP_OP_424J2_126_3477_n1116), .B(
        DP_OP_424J2_126_3477_n1140), .CI(DP_OP_424J2_126_3477_n1138), .CO(
        DP_OP_424J2_126_3477_n890), .S(DP_OP_424J2_126_3477_n891) );
  FADDX1_HVT DP_OP_424J2_126_3477_U601 ( .A(DP_OP_424J2_126_3477_n1110), .B(
        DP_OP_424J2_126_3477_n1136), .CI(DP_OP_424J2_126_3477_n1134), .CO(
        DP_OP_424J2_126_3477_n888), .S(DP_OP_424J2_126_3477_n889) );
  FADDX1_HVT DP_OP_424J2_126_3477_U600 ( .A(DP_OP_424J2_126_3477_n1132), .B(
        DP_OP_424J2_126_3477_n1130), .CI(DP_OP_424J2_126_3477_n1128), .CO(
        DP_OP_424J2_126_3477_n886), .S(DP_OP_424J2_126_3477_n887) );
  FADDX1_HVT DP_OP_424J2_126_3477_U599 ( .A(DP_OP_424J2_126_3477_n1100), .B(
        DP_OP_424J2_126_3477_n1126), .CI(DP_OP_424J2_126_3477_n1124), .CO(
        DP_OP_424J2_126_3477_n884), .S(DP_OP_424J2_126_3477_n885) );
  FADDX1_HVT DP_OP_424J2_126_3477_U598 ( .A(DP_OP_424J2_126_3477_n1106), .B(
        DP_OP_424J2_126_3477_n1122), .CI(DP_OP_424J2_126_3477_n1114), .CO(
        DP_OP_424J2_126_3477_n882), .S(DP_OP_424J2_126_3477_n883) );
  FADDX1_HVT DP_OP_424J2_126_3477_U597 ( .A(DP_OP_424J2_126_3477_n1098), .B(
        DP_OP_424J2_126_3477_n1112), .CI(DP_OP_424J2_126_3477_n1108), .CO(
        DP_OP_424J2_126_3477_n880), .S(DP_OP_424J2_126_3477_n881) );
  FADDX1_HVT DP_OP_424J2_126_3477_U596 ( .A(DP_OP_424J2_126_3477_n1102), .B(
        DP_OP_424J2_126_3477_n1096), .CI(DP_OP_424J2_126_3477_n1104), .CO(
        DP_OP_424J2_126_3477_n878), .S(DP_OP_424J2_126_3477_n879) );
  FADDX1_HVT DP_OP_424J2_126_3477_U595 ( .A(DP_OP_424J2_126_3477_n967), .B(
        DP_OP_424J2_126_3477_n953), .CI(DP_OP_424J2_126_3477_n955), .CO(
        DP_OP_424J2_126_3477_n876), .S(DP_OP_424J2_126_3477_n877) );
  FADDX1_HVT DP_OP_424J2_126_3477_U594 ( .A(DP_OP_424J2_126_3477_n959), .B(
        DP_OP_424J2_126_3477_n937), .CI(DP_OP_424J2_126_3477_n935), .CO(
        DP_OP_424J2_126_3477_n874), .S(DP_OP_424J2_126_3477_n875) );
  FADDX1_HVT DP_OP_424J2_126_3477_U593 ( .A(DP_OP_424J2_126_3477_n951), .B(
        DP_OP_424J2_126_3477_n949), .CI(DP_OP_424J2_126_3477_n945), .CO(
        DP_OP_424J2_126_3477_n872), .S(DP_OP_424J2_126_3477_n873) );
  FADDX1_HVT DP_OP_424J2_126_3477_U592 ( .A(DP_OP_424J2_126_3477_n957), .B(
        DP_OP_424J2_126_3477_n939), .CI(DP_OP_424J2_126_3477_n943), .CO(
        DP_OP_424J2_126_3477_n870), .S(DP_OP_424J2_126_3477_n871) );
  FADDX1_HVT DP_OP_424J2_126_3477_U591 ( .A(DP_OP_424J2_126_3477_n947), .B(
        DP_OP_424J2_126_3477_n965), .CI(DP_OP_424J2_126_3477_n961), .CO(
        DP_OP_424J2_126_3477_n868), .S(DP_OP_424J2_126_3477_n869) );
  FADDX1_HVT DP_OP_424J2_126_3477_U590 ( .A(DP_OP_424J2_126_3477_n941), .B(
        DP_OP_424J2_126_3477_n963), .CI(DP_OP_424J2_126_3477_n923), .CO(
        DP_OP_424J2_126_3477_n866), .S(DP_OP_424J2_126_3477_n867) );
  FADDX1_HVT DP_OP_424J2_126_3477_U589 ( .A(DP_OP_424J2_126_3477_n925), .B(
        DP_OP_424J2_126_3477_n907), .CI(DP_OP_424J2_126_3477_n901), .CO(
        DP_OP_424J2_126_3477_n864), .S(DP_OP_424J2_126_3477_n865) );
  FADDX1_HVT DP_OP_424J2_126_3477_U588 ( .A(DP_OP_424J2_126_3477_n927), .B(
        DP_OP_424J2_126_3477_n903), .CI(DP_OP_424J2_126_3477_n919), .CO(
        DP_OP_424J2_126_3477_n862), .S(DP_OP_424J2_126_3477_n863) );
  FADDX1_HVT DP_OP_424J2_126_3477_U587 ( .A(DP_OP_424J2_126_3477_n917), .B(
        DP_OP_424J2_126_3477_n915), .CI(DP_OP_424J2_126_3477_n905), .CO(
        DP_OP_424J2_126_3477_n860), .S(DP_OP_424J2_126_3477_n861) );
  FADDX1_HVT DP_OP_424J2_126_3477_U586 ( .A(DP_OP_424J2_126_3477_n921), .B(
        DP_OP_424J2_126_3477_n909), .CI(DP_OP_424J2_126_3477_n911), .CO(
        DP_OP_424J2_126_3477_n858), .S(DP_OP_424J2_126_3477_n859) );
  FADDX1_HVT DP_OP_424J2_126_3477_U585 ( .A(DP_OP_424J2_126_3477_n929), .B(
        DP_OP_424J2_126_3477_n933), .CI(DP_OP_424J2_126_3477_n931), .CO(
        DP_OP_424J2_126_3477_n856), .S(DP_OP_424J2_126_3477_n857) );
  FADDX1_HVT DP_OP_424J2_126_3477_U584 ( .A(DP_OP_424J2_126_3477_n913), .B(
        DP_OP_424J2_126_3477_n1092), .CI(DP_OP_424J2_126_3477_n1090), .CO(
        DP_OP_424J2_126_3477_n854), .S(DP_OP_424J2_126_3477_n855) );
  FADDX1_HVT DP_OP_424J2_126_3477_U583 ( .A(DP_OP_424J2_126_3477_n1088), .B(
        DP_OP_424J2_126_3477_n1086), .CI(DP_OP_424J2_126_3477_n1072), .CO(
        DP_OP_424J2_126_3477_n852), .S(DP_OP_424J2_126_3477_n853) );
  FADDX1_HVT DP_OP_424J2_126_3477_U582 ( .A(DP_OP_424J2_126_3477_n1084), .B(
        DP_OP_424J2_126_3477_n1082), .CI(DP_OP_424J2_126_3477_n1070), .CO(
        DP_OP_424J2_126_3477_n850), .S(DP_OP_424J2_126_3477_n851) );
  FADDX1_HVT DP_OP_424J2_126_3477_U581 ( .A(DP_OP_424J2_126_3477_n1080), .B(
        DP_OP_424J2_126_3477_n1074), .CI(DP_OP_424J2_126_3477_n1076), .CO(
        DP_OP_424J2_126_3477_n848), .S(DP_OP_424J2_126_3477_n849) );
  FADDX1_HVT DP_OP_424J2_126_3477_U580 ( .A(DP_OP_424J2_126_3477_n1078), .B(
        DP_OP_424J2_126_3477_n1068), .CI(DP_OP_424J2_126_3477_n1066), .CO(
        DP_OP_424J2_126_3477_n846), .S(DP_OP_424J2_126_3477_n847) );
  FADDX1_HVT DP_OP_424J2_126_3477_U579 ( .A(DP_OP_424J2_126_3477_n899), .B(
        DP_OP_424J2_126_3477_n895), .CI(DP_OP_424J2_126_3477_n1064), .CO(
        DP_OP_424J2_126_3477_n844), .S(DP_OP_424J2_126_3477_n845) );
  FADDX1_HVT DP_OP_424J2_126_3477_U578 ( .A(DP_OP_424J2_126_3477_n897), .B(
        DP_OP_424J2_126_3477_n1052), .CI(DP_OP_424J2_126_3477_n1050), .CO(
        DP_OP_424J2_126_3477_n842), .S(DP_OP_424J2_126_3477_n843) );
  FADDX1_HVT DP_OP_424J2_126_3477_U577 ( .A(DP_OP_424J2_126_3477_n1058), .B(
        DP_OP_424J2_126_3477_n893), .CI(DP_OP_424J2_126_3477_n1048), .CO(
        DP_OP_424J2_126_3477_n840), .S(DP_OP_424J2_126_3477_n841) );
  FADDX1_HVT DP_OP_424J2_126_3477_U576 ( .A(DP_OP_424J2_126_3477_n1056), .B(
        DP_OP_424J2_126_3477_n889), .CI(DP_OP_424J2_126_3477_n879), .CO(
        DP_OP_424J2_126_3477_n838), .S(DP_OP_424J2_126_3477_n839) );
  FADDX1_HVT DP_OP_424J2_126_3477_U575 ( .A(DP_OP_424J2_126_3477_n1062), .B(
        DP_OP_424J2_126_3477_n885), .CI(DP_OP_424J2_126_3477_n887), .CO(
        DP_OP_424J2_126_3477_n836), .S(DP_OP_424J2_126_3477_n837) );
  FADDX1_HVT DP_OP_424J2_126_3477_U574 ( .A(DP_OP_424J2_126_3477_n1060), .B(
        DP_OP_424J2_126_3477_n881), .CI(DP_OP_424J2_126_3477_n883), .CO(
        DP_OP_424J2_126_3477_n834), .S(DP_OP_424J2_126_3477_n835) );
  FADDX1_HVT DP_OP_424J2_126_3477_U573 ( .A(DP_OP_424J2_126_3477_n1054), .B(
        DP_OP_424J2_126_3477_n891), .CI(DP_OP_424J2_126_3477_n877), .CO(
        DP_OP_424J2_126_3477_n832), .S(DP_OP_424J2_126_3477_n833) );
  FADDX1_HVT DP_OP_424J2_126_3477_U572 ( .A(DP_OP_424J2_126_3477_n871), .B(
        DP_OP_424J2_126_3477_n875), .CI(DP_OP_424J2_126_3477_n867), .CO(
        DP_OP_424J2_126_3477_n830), .S(DP_OP_424J2_126_3477_n831) );
  FADDX1_HVT DP_OP_424J2_126_3477_U571 ( .A(DP_OP_424J2_126_3477_n869), .B(
        DP_OP_424J2_126_3477_n873), .CI(DP_OP_424J2_126_3477_n861), .CO(
        DP_OP_424J2_126_3477_n828), .S(DP_OP_424J2_126_3477_n829) );
  FADDX1_HVT DP_OP_424J2_126_3477_U570 ( .A(DP_OP_424J2_126_3477_n859), .B(
        DP_OP_424J2_126_3477_n865), .CI(DP_OP_424J2_126_3477_n1046), .CO(
        DP_OP_424J2_126_3477_n826), .S(DP_OP_424J2_126_3477_n827) );
  FADDX1_HVT DP_OP_424J2_126_3477_U569 ( .A(DP_OP_424J2_126_3477_n857), .B(
        DP_OP_424J2_126_3477_n863), .CI(DP_OP_424J2_126_3477_n1042), .CO(
        DP_OP_424J2_126_3477_n824), .S(DP_OP_424J2_126_3477_n825) );
  FADDX1_HVT DP_OP_424J2_126_3477_U568 ( .A(DP_OP_424J2_126_3477_n1044), .B(
        DP_OP_424J2_126_3477_n1040), .CI(DP_OP_424J2_126_3477_n855), .CO(
        DP_OP_424J2_126_3477_n822), .S(DP_OP_424J2_126_3477_n823) );
  FADDX1_HVT DP_OP_424J2_126_3477_U567 ( .A(DP_OP_424J2_126_3477_n1038), .B(
        DP_OP_424J2_126_3477_n1036), .CI(DP_OP_424J2_126_3477_n853), .CO(
        DP_OP_424J2_126_3477_n820), .S(DP_OP_424J2_126_3477_n821) );
  FADDX1_HVT DP_OP_424J2_126_3477_U566 ( .A(DP_OP_424J2_126_3477_n1034), .B(
        DP_OP_424J2_126_3477_n851), .CI(DP_OP_424J2_126_3477_n849), .CO(
        DP_OP_424J2_126_3477_n818), .S(DP_OP_424J2_126_3477_n819) );
  FADDX1_HVT DP_OP_424J2_126_3477_U565 ( .A(DP_OP_424J2_126_3477_n1032), .B(
        DP_OP_424J2_126_3477_n1026), .CI(DP_OP_424J2_126_3477_n1028), .CO(
        DP_OP_424J2_126_3477_n816), .S(DP_OP_424J2_126_3477_n817) );
  FADDX1_HVT DP_OP_424J2_126_3477_U564 ( .A(DP_OP_424J2_126_3477_n1030), .B(
        DP_OP_424J2_126_3477_n847), .CI(DP_OP_424J2_126_3477_n1024), .CO(
        DP_OP_424J2_126_3477_n814), .S(DP_OP_424J2_126_3477_n815) );
  FADDX1_HVT DP_OP_424J2_126_3477_U563 ( .A(DP_OP_424J2_126_3477_n845), .B(
        DP_OP_424J2_126_3477_n1022), .CI(DP_OP_424J2_126_3477_n843), .CO(
        DP_OP_424J2_126_3477_n812), .S(DP_OP_424J2_126_3477_n813) );
  FADDX1_HVT DP_OP_424J2_126_3477_U562 ( .A(DP_OP_424J2_126_3477_n1020), .B(
        DP_OP_424J2_126_3477_n837), .CI(DP_OP_424J2_126_3477_n833), .CO(
        DP_OP_424J2_126_3477_n810), .S(DP_OP_424J2_126_3477_n811) );
  FADDX1_HVT DP_OP_424J2_126_3477_U561 ( .A(DP_OP_424J2_126_3477_n1018), .B(
        DP_OP_424J2_126_3477_n841), .CI(DP_OP_424J2_126_3477_n839), .CO(
        DP_OP_424J2_126_3477_n808), .S(DP_OP_424J2_126_3477_n809) );
  FADDX1_HVT DP_OP_424J2_126_3477_U560 ( .A(DP_OP_424J2_126_3477_n835), .B(
        DP_OP_424J2_126_3477_n1016), .CI(DP_OP_424J2_126_3477_n831), .CO(
        DP_OP_424J2_126_3477_n806), .S(DP_OP_424J2_126_3477_n807) );
  FADDX1_HVT DP_OP_424J2_126_3477_U559 ( .A(DP_OP_424J2_126_3477_n829), .B(
        DP_OP_424J2_126_3477_n1014), .CI(DP_OP_424J2_126_3477_n827), .CO(
        DP_OP_424J2_126_3477_n804), .S(DP_OP_424J2_126_3477_n805) );
  FADDX1_HVT DP_OP_424J2_126_3477_U558 ( .A(DP_OP_424J2_126_3477_n825), .B(
        DP_OP_424J2_126_3477_n1012), .CI(DP_OP_424J2_126_3477_n1008), .CO(
        DP_OP_424J2_126_3477_n802), .S(DP_OP_424J2_126_3477_n803) );
  FADDX1_HVT DP_OP_424J2_126_3477_U557 ( .A(DP_OP_424J2_126_3477_n1010), .B(
        DP_OP_424J2_126_3477_n823), .CI(DP_OP_424J2_126_3477_n1006), .CO(
        DP_OP_424J2_126_3477_n800), .S(DP_OP_424J2_126_3477_n801) );
  FADDX1_HVT DP_OP_424J2_126_3477_U556 ( .A(DP_OP_424J2_126_3477_n821), .B(
        DP_OP_424J2_126_3477_n1004), .CI(DP_OP_424J2_126_3477_n1002), .CO(
        DP_OP_424J2_126_3477_n798), .S(DP_OP_424J2_126_3477_n799) );
  FADDX1_HVT DP_OP_424J2_126_3477_U555 ( .A(DP_OP_424J2_126_3477_n819), .B(
        DP_OP_424J2_126_3477_n1000), .CI(DP_OP_424J2_126_3477_n815), .CO(
        DP_OP_424J2_126_3477_n796), .S(DP_OP_424J2_126_3477_n797) );
  FADDX1_HVT DP_OP_424J2_126_3477_U554 ( .A(DP_OP_424J2_126_3477_n817), .B(
        DP_OP_424J2_126_3477_n998), .CI(DP_OP_424J2_126_3477_n813), .CO(
        DP_OP_424J2_126_3477_n794), .S(DP_OP_424J2_126_3477_n795) );
  FADDX1_HVT DP_OP_424J2_126_3477_U553 ( .A(DP_OP_424J2_126_3477_n996), .B(
        DP_OP_424J2_126_3477_n811), .CI(DP_OP_424J2_126_3477_n807), .CO(
        DP_OP_424J2_126_3477_n792), .S(DP_OP_424J2_126_3477_n793) );
  FADDX1_HVT DP_OP_424J2_126_3477_U552 ( .A(DP_OP_424J2_126_3477_n809), .B(
        DP_OP_424J2_126_3477_n994), .CI(DP_OP_424J2_126_3477_n805), .CO(
        DP_OP_424J2_126_3477_n790), .S(DP_OP_424J2_126_3477_n791) );
  FADDX1_HVT DP_OP_424J2_126_3477_U551 ( .A(DP_OP_424J2_126_3477_n992), .B(
        DP_OP_424J2_126_3477_n803), .CI(DP_OP_424J2_126_3477_n990), .CO(
        DP_OP_424J2_126_3477_n788), .S(DP_OP_424J2_126_3477_n789) );
  FADDX1_HVT DP_OP_424J2_126_3477_U550 ( .A(DP_OP_424J2_126_3477_n801), .B(
        DP_OP_424J2_126_3477_n988), .CI(DP_OP_424J2_126_3477_n799), .CO(
        DP_OP_424J2_126_3477_n786), .S(DP_OP_424J2_126_3477_n787) );
  FADDX1_HVT DP_OP_424J2_126_3477_U549 ( .A(DP_OP_424J2_126_3477_n986), .B(
        DP_OP_424J2_126_3477_n797), .CI(DP_OP_424J2_126_3477_n984), .CO(
        DP_OP_424J2_126_3477_n784), .S(DP_OP_424J2_126_3477_n785) );
  FADDX1_HVT DP_OP_424J2_126_3477_U548 ( .A(DP_OP_424J2_126_3477_n795), .B(
        DP_OP_424J2_126_3477_n793), .CI(DP_OP_424J2_126_3477_n982), .CO(
        DP_OP_424J2_126_3477_n782), .S(DP_OP_424J2_126_3477_n783) );
  FADDX1_HVT DP_OP_424J2_126_3477_U547 ( .A(DP_OP_424J2_126_3477_n791), .B(
        DP_OP_424J2_126_3477_n980), .CI(DP_OP_424J2_126_3477_n789), .CO(
        DP_OP_424J2_126_3477_n780), .S(DP_OP_424J2_126_3477_n781) );
  FADDX1_HVT DP_OP_424J2_126_3477_U546 ( .A(DP_OP_424J2_126_3477_n978), .B(
        DP_OP_424J2_126_3477_n787), .CI(DP_OP_424J2_126_3477_n976), .CO(
        DP_OP_424J2_126_3477_n778), .S(DP_OP_424J2_126_3477_n779) );
  FADDX1_HVT DP_OP_424J2_126_3477_U545 ( .A(DP_OP_424J2_126_3477_n785), .B(
        DP_OP_424J2_126_3477_n974), .CI(DP_OP_424J2_126_3477_n783), .CO(
        DP_OP_424J2_126_3477_n776), .S(DP_OP_424J2_126_3477_n777) );
  FADDX1_HVT DP_OP_424J2_126_3477_U544 ( .A(DP_OP_424J2_126_3477_n781), .B(
        DP_OP_424J2_126_3477_n972), .CI(DP_OP_424J2_126_3477_n779), .CO(
        DP_OP_424J2_126_3477_n774), .S(DP_OP_424J2_126_3477_n775) );
  FADDX1_HVT DP_OP_424J2_126_3477_U543 ( .A(DP_OP_424J2_126_3477_n970), .B(
        DP_OP_424J2_126_3477_n777), .CI(DP_OP_424J2_126_3477_n775), .CO(
        DP_OP_424J2_126_3477_n772), .S(DP_OP_424J2_126_3477_n773) );
  FADDX1_HVT DP_OP_424J2_126_3477_U541 ( .A(DP_OP_424J2_126_3477_n2186), .B(
        DP_OP_424J2_126_3477_n1922), .CI(DP_OP_424J2_126_3477_n1878), .CO(
        DP_OP_424J2_126_3477_n768), .S(DP_OP_424J2_126_3477_n769) );
  FADDX1_HVT DP_OP_424J2_126_3477_U540 ( .A(DP_OP_424J2_126_3477_n2758), .B(
        DP_OP_424J2_126_3477_n1980), .CI(DP_OP_424J2_126_3477_n2244), .CO(
        DP_OP_424J2_126_3477_n766), .S(DP_OP_424J2_126_3477_n767) );
  FADDX1_HVT DP_OP_424J2_126_3477_U539 ( .A(DP_OP_424J2_126_3477_n2230), .B(
        DP_OP_424J2_126_3477_n2990), .CI(DP_OP_424J2_126_3477_n2640), .CO(
        DP_OP_424J2_126_3477_n764), .S(DP_OP_424J2_126_3477_n765) );
  FADDX1_HVT DP_OP_424J2_126_3477_U538 ( .A(DP_OP_424J2_126_3477_n2450), .B(
        DP_OP_424J2_126_3477_n2024), .CI(DP_OP_424J2_126_3477_n2068), .CO(
        DP_OP_424J2_126_3477_n762), .S(DP_OP_424J2_126_3477_n763) );
  FADDX1_HVT DP_OP_424J2_126_3477_U537 ( .A(DP_OP_424J2_126_3477_n2010), .B(
        DP_OP_424J2_126_3477_n2112), .CI(DP_OP_424J2_126_3477_n2156), .CO(
        DP_OP_424J2_126_3477_n760), .S(DP_OP_424J2_126_3477_n761) );
  FADDX1_HVT DP_OP_424J2_126_3477_U536 ( .A(DP_OP_424J2_126_3477_n2714), .B(
        DP_OP_424J2_126_3477_n2816), .CI(DP_OP_424J2_126_3477_n2860), .CO(
        DP_OP_424J2_126_3477_n758), .S(DP_OP_424J2_126_3477_n759) );
  FADDX1_HVT DP_OP_424J2_126_3477_U535 ( .A(DP_OP_424J2_126_3477_n2054), .B(
        DP_OP_424J2_126_3477_n2772), .CI(DP_OP_424J2_126_3477_n2596), .CO(
        DP_OP_424J2_126_3477_n756), .S(DP_OP_424J2_126_3477_n757) );
  FADDX1_HVT DP_OP_424J2_126_3477_U534 ( .A(DP_OP_424J2_126_3477_n2142), .B(
        DP_OP_424J2_126_3477_n2420), .CI(DP_OP_424J2_126_3477_n2948), .CO(
        DP_OP_424J2_126_3477_n754), .S(DP_OP_424J2_126_3477_n755) );
  FADDX1_HVT DP_OP_424J2_126_3477_U533 ( .A(DP_OP_424J2_126_3477_n2670), .B(
        DP_OP_424J2_126_3477_n2904), .CI(DP_OP_424J2_126_3477_n2464), .CO(
        DP_OP_424J2_126_3477_n752), .S(DP_OP_424J2_126_3477_n753) );
  FADDX1_HVT DP_OP_424J2_126_3477_U532 ( .A(DP_OP_424J2_126_3477_n2626), .B(
        DP_OP_424J2_126_3477_n2376), .CI(DP_OP_424J2_126_3477_n2728), .CO(
        DP_OP_424J2_126_3477_n750), .S(DP_OP_424J2_126_3477_n751) );
  FADDX1_HVT DP_OP_424J2_126_3477_U531 ( .A(DP_OP_424J2_126_3477_n2846), .B(
        DP_OP_424J2_126_3477_n2508), .CI(DP_OP_424J2_126_3477_n2332), .CO(
        DP_OP_424J2_126_3477_n748), .S(DP_OP_424J2_126_3477_n749) );
  FADDX1_HVT DP_OP_424J2_126_3477_U530 ( .A(DP_OP_424J2_126_3477_n2318), .B(
        DP_OP_424J2_126_3477_n2288), .CI(DP_OP_424J2_126_3477_n1936), .CO(
        DP_OP_424J2_126_3477_n746), .S(DP_OP_424J2_126_3477_n747) );
  FADDX1_HVT DP_OP_424J2_126_3477_U529 ( .A(DP_OP_424J2_126_3477_n2538), .B(
        DP_OP_424J2_126_3477_n2200), .CI(DP_OP_424J2_126_3477_n2552), .CO(
        DP_OP_424J2_126_3477_n744), .S(DP_OP_424J2_126_3477_n745) );
  FADDX1_HVT DP_OP_424J2_126_3477_U528 ( .A(DP_OP_424J2_126_3477_n2494), .B(
        DP_OP_424J2_126_3477_n2362), .CI(DP_OP_424J2_126_3477_n2684), .CO(
        DP_OP_424J2_126_3477_n742), .S(DP_OP_424J2_126_3477_n743) );
  FADDX1_HVT DP_OP_424J2_126_3477_U527 ( .A(DP_OP_424J2_126_3477_n2802), .B(
        DP_OP_424J2_126_3477_n2098), .CI(DP_OP_424J2_126_3477_n2274), .CO(
        DP_OP_424J2_126_3477_n740), .S(DP_OP_424J2_126_3477_n741) );
  FADDX1_HVT DP_OP_424J2_126_3477_U526 ( .A(DP_OP_424J2_126_3477_n1966), .B(
        DP_OP_424J2_126_3477_n2582), .CI(DP_OP_424J2_126_3477_n2934), .CO(
        DP_OP_424J2_126_3477_n738), .S(DP_OP_424J2_126_3477_n739) );
  FADDX1_HVT DP_OP_424J2_126_3477_U525 ( .A(DP_OP_424J2_126_3477_n2890), .B(
        DP_OP_424J2_126_3477_n2406), .CI(DP_OP_424J2_126_3477_n771), .CO(
        DP_OP_424J2_126_3477_n736), .S(DP_OP_424J2_126_3477_n737) );
  FADDX1_HVT DP_OP_424J2_126_3477_U524 ( .A(DP_OP_424J2_126_3477_n2237), .B(
        DP_OP_424J2_126_3477_n1973), .CI(DP_OP_424J2_126_3477_n1929), .CO(
        DP_OP_424J2_126_3477_n734), .S(DP_OP_424J2_126_3477_n735) );
  FADDX1_HVT DP_OP_424J2_126_3477_U523 ( .A(DP_OP_424J2_126_3477_n2983), .B(
        DP_OP_424J2_126_3477_n2017), .CI(DP_OP_424J2_126_3477_n2061), .CO(
        DP_OP_424J2_126_3477_n732), .S(DP_OP_424J2_126_3477_n733) );
  FADDX1_HVT DP_OP_424J2_126_3477_U522 ( .A(DP_OP_424J2_126_3477_n2941), .B(
        DP_OP_424J2_126_3477_n2105), .CI(DP_OP_424J2_126_3477_n2149), .CO(
        DP_OP_424J2_126_3477_n730), .S(DP_OP_424J2_126_3477_n731) );
  FADDX1_HVT DP_OP_424J2_126_3477_U521 ( .A(DP_OP_424J2_126_3477_n2897), .B(
        DP_OP_424J2_126_3477_n2193), .CI(DP_OP_424J2_126_3477_n2281), .CO(
        DP_OP_424J2_126_3477_n728), .S(DP_OP_424J2_126_3477_n729) );
  FADDX1_HVT DP_OP_424J2_126_3477_U520 ( .A(DP_OP_424J2_126_3477_n2853), .B(
        DP_OP_424J2_126_3477_n2325), .CI(DP_OP_424J2_126_3477_n2369), .CO(
        DP_OP_424J2_126_3477_n726), .S(DP_OP_424J2_126_3477_n727) );
  FADDX1_HVT DP_OP_424J2_126_3477_U519 ( .A(DP_OP_424J2_126_3477_n2809), .B(
        DP_OP_424J2_126_3477_n2413), .CI(DP_OP_424J2_126_3477_n2457), .CO(
        DP_OP_424J2_126_3477_n724), .S(DP_OP_424J2_126_3477_n725) );
  FADDX1_HVT DP_OP_424J2_126_3477_U518 ( .A(DP_OP_424J2_126_3477_n2765), .B(
        DP_OP_424J2_126_3477_n2501), .CI(DP_OP_424J2_126_3477_n2545), .CO(
        DP_OP_424J2_126_3477_n722), .S(DP_OP_424J2_126_3477_n723) );
  FADDX1_HVT DP_OP_424J2_126_3477_U517 ( .A(DP_OP_424J2_126_3477_n2721), .B(
        DP_OP_424J2_126_3477_n2589), .CI(DP_OP_424J2_126_3477_n2633), .CO(
        DP_OP_424J2_126_3477_n720), .S(DP_OP_424J2_126_3477_n721) );
  FADDX1_HVT DP_OP_424J2_126_3477_U516 ( .A(DP_OP_424J2_126_3477_n2677), .B(
        DP_OP_424J2_126_3477_n966), .CI(DP_OP_424J2_126_3477_n964), .CO(
        DP_OP_424J2_126_3477_n718), .S(DP_OP_424J2_126_3477_n719) );
  FADDX1_HVT DP_OP_424J2_126_3477_U515 ( .A(DP_OP_424J2_126_3477_n962), .B(
        DP_OP_424J2_126_3477_n934), .CI(DP_OP_424J2_126_3477_n936), .CO(
        DP_OP_424J2_126_3477_n716), .S(DP_OP_424J2_126_3477_n717) );
  FADDX1_HVT DP_OP_424J2_126_3477_U514 ( .A(DP_OP_424J2_126_3477_n960), .B(
        DP_OP_424J2_126_3477_n938), .CI(DP_OP_424J2_126_3477_n940), .CO(
        DP_OP_424J2_126_3477_n714), .S(DP_OP_424J2_126_3477_n715) );
  FADDX1_HVT DP_OP_424J2_126_3477_U513 ( .A(DP_OP_424J2_126_3477_n958), .B(
        DP_OP_424J2_126_3477_n942), .CI(DP_OP_424J2_126_3477_n944), .CO(
        DP_OP_424J2_126_3477_n712), .S(DP_OP_424J2_126_3477_n713) );
  FADDX1_HVT DP_OP_424J2_126_3477_U512 ( .A(DP_OP_424J2_126_3477_n950), .B(
        DP_OP_424J2_126_3477_n956), .CI(DP_OP_424J2_126_3477_n946), .CO(
        DP_OP_424J2_126_3477_n710), .S(DP_OP_424J2_126_3477_n711) );
  FADDX1_HVT DP_OP_424J2_126_3477_U511 ( .A(DP_OP_424J2_126_3477_n948), .B(
        DP_OP_424J2_126_3477_n952), .CI(DP_OP_424J2_126_3477_n954), .CO(
        DP_OP_424J2_126_3477_n708), .S(DP_OP_424J2_126_3477_n709) );
  FADDX1_HVT DP_OP_424J2_126_3477_U510 ( .A(DP_OP_424J2_126_3477_n932), .B(
        DP_OP_424J2_126_3477_n930), .CI(DP_OP_424J2_126_3477_n900), .CO(
        DP_OP_424J2_126_3477_n706), .S(DP_OP_424J2_126_3477_n707) );
  FADDX1_HVT DP_OP_424J2_126_3477_U509 ( .A(DP_OP_424J2_126_3477_n914), .B(
        DP_OP_424J2_126_3477_n902), .CI(DP_OP_424J2_126_3477_n904), .CO(
        DP_OP_424J2_126_3477_n704), .S(DP_OP_424J2_126_3477_n705) );
  FADDX1_HVT DP_OP_424J2_126_3477_U508 ( .A(DP_OP_424J2_126_3477_n912), .B(
        DP_OP_424J2_126_3477_n906), .CI(DP_OP_424J2_126_3477_n908), .CO(
        DP_OP_424J2_126_3477_n702), .S(DP_OP_424J2_126_3477_n703) );
  FADDX1_HVT DP_OP_424J2_126_3477_U507 ( .A(DP_OP_424J2_126_3477_n910), .B(
        DP_OP_424J2_126_3477_n928), .CI(DP_OP_424J2_126_3477_n926), .CO(
        DP_OP_424J2_126_3477_n700), .S(DP_OP_424J2_126_3477_n701) );
  FADDX1_HVT DP_OP_424J2_126_3477_U506 ( .A(DP_OP_424J2_126_3477_n920), .B(
        DP_OP_424J2_126_3477_n916), .CI(DP_OP_424J2_126_3477_n918), .CO(
        DP_OP_424J2_126_3477_n698), .S(DP_OP_424J2_126_3477_n699) );
  FADDX1_HVT DP_OP_424J2_126_3477_U505 ( .A(DP_OP_424J2_126_3477_n924), .B(
        DP_OP_424J2_126_3477_n922), .CI(DP_OP_424J2_126_3477_n763), .CO(
        DP_OP_424J2_126_3477_n696), .S(DP_OP_424J2_126_3477_n697) );
  FADDX1_HVT DP_OP_424J2_126_3477_U504 ( .A(DP_OP_424J2_126_3477_n759), .B(
        DP_OP_424J2_126_3477_n755), .CI(DP_OP_424J2_126_3477_n737), .CO(
        DP_OP_424J2_126_3477_n694), .S(DP_OP_424J2_126_3477_n695) );
  FADDX1_HVT DP_OP_424J2_126_3477_U503 ( .A(DP_OP_424J2_126_3477_n761), .B(
        DP_OP_424J2_126_3477_n743), .CI(DP_OP_424J2_126_3477_n741), .CO(
        DP_OP_424J2_126_3477_n692), .S(DP_OP_424J2_126_3477_n693) );
  FADDX1_HVT DP_OP_424J2_126_3477_U502 ( .A(DP_OP_424J2_126_3477_n753), .B(
        DP_OP_424J2_126_3477_n757), .CI(DP_OP_424J2_126_3477_n749), .CO(
        DP_OP_424J2_126_3477_n690), .S(DP_OP_424J2_126_3477_n691) );
  FADDX1_HVT DP_OP_424J2_126_3477_U501 ( .A(DP_OP_424J2_126_3477_n765), .B(
        DP_OP_424J2_126_3477_n745), .CI(DP_OP_424J2_126_3477_n739), .CO(
        DP_OP_424J2_126_3477_n688), .S(DP_OP_424J2_126_3477_n689) );
  FADDX1_HVT DP_OP_424J2_126_3477_U500 ( .A(DP_OP_424J2_126_3477_n747), .B(
        DP_OP_424J2_126_3477_n769), .CI(DP_OP_424J2_126_3477_n767), .CO(
        DP_OP_424J2_126_3477_n686), .S(DP_OP_424J2_126_3477_n687) );
  FADDX1_HVT DP_OP_424J2_126_3477_U499 ( .A(DP_OP_424J2_126_3477_n751), .B(
        DP_OP_424J2_126_3477_n731), .CI(DP_OP_424J2_126_3477_n727), .CO(
        DP_OP_424J2_126_3477_n684), .S(DP_OP_424J2_126_3477_n685) );
  FADDX1_HVT DP_OP_424J2_126_3477_U498 ( .A(DP_OP_424J2_126_3477_n723), .B(
        DP_OP_424J2_126_3477_n721), .CI(DP_OP_424J2_126_3477_n733), .CO(
        DP_OP_424J2_126_3477_n682), .S(DP_OP_424J2_126_3477_n683) );
  FADDX1_HVT DP_OP_424J2_126_3477_U497 ( .A(DP_OP_424J2_126_3477_n729), .B(
        DP_OP_424J2_126_3477_n725), .CI(DP_OP_424J2_126_3477_n735), .CO(
        DP_OP_424J2_126_3477_n680), .S(DP_OP_424J2_126_3477_n681) );
  FADDX1_HVT DP_OP_424J2_126_3477_U496 ( .A(DP_OP_424J2_126_3477_n898), .B(
        DP_OP_424J2_126_3477_n894), .CI(DP_OP_424J2_126_3477_n896), .CO(
        DP_OP_424J2_126_3477_n678), .S(DP_OP_424J2_126_3477_n679) );
  FADDX1_HVT DP_OP_424J2_126_3477_U495 ( .A(DP_OP_424J2_126_3477_n892), .B(
        DP_OP_424J2_126_3477_n878), .CI(DP_OP_424J2_126_3477_n880), .CO(
        DP_OP_424J2_126_3477_n676), .S(DP_OP_424J2_126_3477_n677) );
  FADDX1_HVT DP_OP_424J2_126_3477_U494 ( .A(DP_OP_424J2_126_3477_n890), .B(
        DP_OP_424J2_126_3477_n882), .CI(DP_OP_424J2_126_3477_n888), .CO(
        DP_OP_424J2_126_3477_n674), .S(DP_OP_424J2_126_3477_n675) );
  FADDX1_HVT DP_OP_424J2_126_3477_U493 ( .A(DP_OP_424J2_126_3477_n886), .B(
        DP_OP_424J2_126_3477_n884), .CI(DP_OP_424J2_126_3477_n719), .CO(
        DP_OP_424J2_126_3477_n672), .S(DP_OP_424J2_126_3477_n673) );
  FADDX1_HVT DP_OP_424J2_126_3477_U492 ( .A(DP_OP_424J2_126_3477_n876), .B(
        DP_OP_424J2_126_3477_n717), .CI(DP_OP_424J2_126_3477_n715), .CO(
        DP_OP_424J2_126_3477_n670), .S(DP_OP_424J2_126_3477_n671) );
  FADDX1_HVT DP_OP_424J2_126_3477_U491 ( .A(DP_OP_424J2_126_3477_n874), .B(
        DP_OP_424J2_126_3477_n711), .CI(DP_OP_424J2_126_3477_n713), .CO(
        DP_OP_424J2_126_3477_n668), .S(DP_OP_424J2_126_3477_n669) );
  FADDX1_HVT DP_OP_424J2_126_3477_U490 ( .A(DP_OP_424J2_126_3477_n872), .B(
        DP_OP_424J2_126_3477_n709), .CI(DP_OP_424J2_126_3477_n866), .CO(
        DP_OP_424J2_126_3477_n666), .S(DP_OP_424J2_126_3477_n667) );
  FADDX1_HVT DP_OP_424J2_126_3477_U489 ( .A(DP_OP_424J2_126_3477_n870), .B(
        DP_OP_424J2_126_3477_n868), .CI(DP_OP_424J2_126_3477_n856), .CO(
        DP_OP_424J2_126_3477_n664), .S(DP_OP_424J2_126_3477_n665) );
  FADDX1_HVT DP_OP_424J2_126_3477_U488 ( .A(DP_OP_424J2_126_3477_n864), .B(
        DP_OP_424J2_126_3477_n707), .CI(DP_OP_424J2_126_3477_n697), .CO(
        DP_OP_424J2_126_3477_n662), .S(DP_OP_424J2_126_3477_n663) );
  FADDX1_HVT DP_OP_424J2_126_3477_U487 ( .A(DP_OP_424J2_126_3477_n862), .B(
        DP_OP_424J2_126_3477_n703), .CI(DP_OP_424J2_126_3477_n699), .CO(
        DP_OP_424J2_126_3477_n660), .S(DP_OP_424J2_126_3477_n661) );
  FADDX1_HVT DP_OP_424J2_126_3477_U486 ( .A(DP_OP_424J2_126_3477_n860), .B(
        DP_OP_424J2_126_3477_n705), .CI(DP_OP_424J2_126_3477_n701), .CO(
        DP_OP_424J2_126_3477_n658), .S(DP_OP_424J2_126_3477_n659) );
  FADDX1_HVT DP_OP_424J2_126_3477_U485 ( .A(DP_OP_424J2_126_3477_n858), .B(
        DP_OP_424J2_126_3477_n693), .CI(DP_OP_424J2_126_3477_n689), .CO(
        DP_OP_424J2_126_3477_n656), .S(DP_OP_424J2_126_3477_n657) );
  FADDX1_HVT DP_OP_424J2_126_3477_U484 ( .A(DP_OP_424J2_126_3477_n691), .B(
        DP_OP_424J2_126_3477_n854), .CI(DP_OP_424J2_126_3477_n685), .CO(
        DP_OP_424J2_126_3477_n654), .S(DP_OP_424J2_126_3477_n655) );
  FADDX1_HVT DP_OP_424J2_126_3477_U483 ( .A(DP_OP_424J2_126_3477_n687), .B(
        DP_OP_424J2_126_3477_n695), .CI(DP_OP_424J2_126_3477_n681), .CO(
        DP_OP_424J2_126_3477_n652), .S(DP_OP_424J2_126_3477_n653) );
  FADDX1_HVT DP_OP_424J2_126_3477_U482 ( .A(DP_OP_424J2_126_3477_n683), .B(
        DP_OP_424J2_126_3477_n852), .CI(DP_OP_424J2_126_3477_n850), .CO(
        DP_OP_424J2_126_3477_n650), .S(DP_OP_424J2_126_3477_n651) );
  FADDX1_HVT DP_OP_424J2_126_3477_U481 ( .A(DP_OP_424J2_126_3477_n848), .B(
        DP_OP_424J2_126_3477_n846), .CI(DP_OP_424J2_126_3477_n679), .CO(
        DP_OP_424J2_126_3477_n648), .S(DP_OP_424J2_126_3477_n649) );
  FADDX1_HVT DP_OP_424J2_126_3477_U480 ( .A(DP_OP_424J2_126_3477_n844), .B(
        DP_OP_424J2_126_3477_n842), .CI(DP_OP_424J2_126_3477_n840), .CO(
        DP_OP_424J2_126_3477_n646), .S(DP_OP_424J2_126_3477_n647) );
  FADDX1_HVT DP_OP_424J2_126_3477_U479 ( .A(DP_OP_424J2_126_3477_n838), .B(
        DP_OP_424J2_126_3477_n673), .CI(DP_OP_424J2_126_3477_n832), .CO(
        DP_OP_424J2_126_3477_n644), .S(DP_OP_424J2_126_3477_n645) );
  FADDX1_HVT DP_OP_424J2_126_3477_U478 ( .A(DP_OP_424J2_126_3477_n836), .B(
        DP_OP_424J2_126_3477_n675), .CI(DP_OP_424J2_126_3477_n677), .CO(
        DP_OP_424J2_126_3477_n642), .S(DP_OP_424J2_126_3477_n643) );
  FADDX1_HVT DP_OP_424J2_126_3477_U477 ( .A(DP_OP_424J2_126_3477_n834), .B(
        DP_OP_424J2_126_3477_n671), .CI(DP_OP_424J2_126_3477_n667), .CO(
        DP_OP_424J2_126_3477_n640), .S(DP_OP_424J2_126_3477_n641) );
  FADDX1_HVT DP_OP_424J2_126_3477_U476 ( .A(DP_OP_424J2_126_3477_n830), .B(
        DP_OP_424J2_126_3477_n669), .CI(DP_OP_424J2_126_3477_n665), .CO(
        DP_OP_424J2_126_3477_n638), .S(DP_OP_424J2_126_3477_n639) );
  FADDX1_HVT DP_OP_424J2_126_3477_U475 ( .A(DP_OP_424J2_126_3477_n828), .B(
        DP_OP_424J2_126_3477_n826), .CI(DP_OP_424J2_126_3477_n661), .CO(
        DP_OP_424J2_126_3477_n636), .S(DP_OP_424J2_126_3477_n637) );
  FADDX1_HVT DP_OP_424J2_126_3477_U474 ( .A(DP_OP_424J2_126_3477_n659), .B(
        DP_OP_424J2_126_3477_n663), .CI(DP_OP_424J2_126_3477_n824), .CO(
        DP_OP_424J2_126_3477_n634), .S(DP_OP_424J2_126_3477_n635) );
  FADDX1_HVT DP_OP_424J2_126_3477_U473 ( .A(DP_OP_424J2_126_3477_n657), .B(
        DP_OP_424J2_126_3477_n822), .CI(DP_OP_424J2_126_3477_n653), .CO(
        DP_OP_424J2_126_3477_n632), .S(DP_OP_424J2_126_3477_n633) );
  FADDX1_HVT DP_OP_424J2_126_3477_U472 ( .A(DP_OP_424J2_126_3477_n655), .B(
        DP_OP_424J2_126_3477_n820), .CI(DP_OP_424J2_126_3477_n651), .CO(
        DP_OP_424J2_126_3477_n630), .S(DP_OP_424J2_126_3477_n631) );
  FADDX1_HVT DP_OP_424J2_126_3477_U471 ( .A(DP_OP_424J2_126_3477_n818), .B(
        DP_OP_424J2_126_3477_n816), .CI(DP_OP_424J2_126_3477_n649), .CO(
        DP_OP_424J2_126_3477_n628), .S(DP_OP_424J2_126_3477_n629) );
  FADDX1_HVT DP_OP_424J2_126_3477_U470 ( .A(DP_OP_424J2_126_3477_n814), .B(
        DP_OP_424J2_126_3477_n812), .CI(DP_OP_424J2_126_3477_n647), .CO(
        DP_OP_424J2_126_3477_n626), .S(DP_OP_424J2_126_3477_n627) );
  FADDX1_HVT DP_OP_424J2_126_3477_U469 ( .A(DP_OP_424J2_126_3477_n810), .B(
        DP_OP_424J2_126_3477_n643), .CI(DP_OP_424J2_126_3477_n806), .CO(
        DP_OP_424J2_126_3477_n624), .S(DP_OP_424J2_126_3477_n625) );
  FADDX1_HVT DP_OP_424J2_126_3477_U468 ( .A(DP_OP_424J2_126_3477_n808), .B(
        DP_OP_424J2_126_3477_n645), .CI(DP_OP_424J2_126_3477_n641), .CO(
        DP_OP_424J2_126_3477_n622), .S(DP_OP_424J2_126_3477_n623) );
  FADDX1_HVT DP_OP_424J2_126_3477_U467 ( .A(DP_OP_424J2_126_3477_n639), .B(
        DP_OP_424J2_126_3477_n804), .CI(DP_OP_424J2_126_3477_n637), .CO(
        DP_OP_424J2_126_3477_n620), .S(DP_OP_424J2_126_3477_n621) );
  FADDX1_HVT DP_OP_424J2_126_3477_U466 ( .A(DP_OP_424J2_126_3477_n635), .B(
        DP_OP_424J2_126_3477_n802), .CI(DP_OP_424J2_126_3477_n633), .CO(
        DP_OP_424J2_126_3477_n618), .S(DP_OP_424J2_126_3477_n619) );
  FADDX1_HVT DP_OP_424J2_126_3477_U465 ( .A(DP_OP_424J2_126_3477_n800), .B(
        DP_OP_424J2_126_3477_n631), .CI(DP_OP_424J2_126_3477_n798), .CO(
        DP_OP_424J2_126_3477_n616), .S(DP_OP_424J2_126_3477_n617) );
  FADDX1_HVT DP_OP_424J2_126_3477_U464 ( .A(DP_OP_424J2_126_3477_n796), .B(
        DP_OP_424J2_126_3477_n629), .CI(DP_OP_424J2_126_3477_n794), .CO(
        DP_OP_424J2_126_3477_n614), .S(DP_OP_424J2_126_3477_n615) );
  FADDX1_HVT DP_OP_424J2_126_3477_U463 ( .A(DP_OP_424J2_126_3477_n627), .B(
        DP_OP_424J2_126_3477_n792), .CI(DP_OP_424J2_126_3477_n625), .CO(
        DP_OP_424J2_126_3477_n612), .S(DP_OP_424J2_126_3477_n613) );
  FADDX1_HVT DP_OP_424J2_126_3477_U462 ( .A(DP_OP_424J2_126_3477_n623), .B(
        DP_OP_424J2_126_3477_n790), .CI(DP_OP_424J2_126_3477_n621), .CO(
        DP_OP_424J2_126_3477_n610), .S(DP_OP_424J2_126_3477_n611) );
  FADDX1_HVT DP_OP_424J2_126_3477_U461 ( .A(DP_OP_424J2_126_3477_n788), .B(
        DP_OP_424J2_126_3477_n619), .CI(DP_OP_424J2_126_3477_n786), .CO(
        DP_OP_424J2_126_3477_n608), .S(DP_OP_424J2_126_3477_n609) );
  FADDX1_HVT DP_OP_424J2_126_3477_U460 ( .A(DP_OP_424J2_126_3477_n617), .B(
        DP_OP_424J2_126_3477_n784), .CI(DP_OP_424J2_126_3477_n615), .CO(
        DP_OP_424J2_126_3477_n606), .S(DP_OP_424J2_126_3477_n607) );
  FADDX1_HVT DP_OP_424J2_126_3477_U459 ( .A(DP_OP_424J2_126_3477_n782), .B(
        DP_OP_424J2_126_3477_n613), .CI(DP_OP_424J2_126_3477_n611), .CO(
        DP_OP_424J2_126_3477_n604), .S(DP_OP_424J2_126_3477_n605) );
  FADDX1_HVT DP_OP_424J2_126_3477_U458 ( .A(DP_OP_424J2_126_3477_n780), .B(
        DP_OP_424J2_126_3477_n609), .CI(DP_OP_424J2_126_3477_n778), .CO(
        DP_OP_424J2_126_3477_n602), .S(DP_OP_424J2_126_3477_n603) );
  FADDX1_HVT DP_OP_424J2_126_3477_U457 ( .A(DP_OP_424J2_126_3477_n607), .B(
        DP_OP_424J2_126_3477_n776), .CI(DP_OP_424J2_126_3477_n605), .CO(
        DP_OP_424J2_126_3477_n600), .S(DP_OP_424J2_126_3477_n601) );
  FADDX1_HVT DP_OP_424J2_126_3477_U456 ( .A(DP_OP_424J2_126_3477_n774), .B(
        DP_OP_424J2_126_3477_n603), .CI(DP_OP_424J2_126_3477_n601), .CO(
        DP_OP_424J2_126_3477_n598), .S(DP_OP_424J2_126_3477_n599) );
  FADDX1_HVT DP_OP_424J2_126_3477_U455 ( .A(DP_OP_424J2_126_3477_n2977), .B(
        DP_OP_424J2_126_3477_n1921), .CI(DP_OP_424J2_126_3477_n1877), .CO(
        DP_OP_424J2_126_3477_n596), .S(DP_OP_424J2_126_3477_n597) );
  FADDX1_HVT DP_OP_424J2_126_3477_U454 ( .A(DP_OP_424J2_126_3477_n770), .B(
        DP_OP_424J2_126_3477_n2236), .CI(DP_OP_424J2_126_3477_n1928), .CO(
        DP_OP_424J2_126_3477_n594), .S(DP_OP_424J2_126_3477_n595) );
  FADDX1_HVT DP_OP_424J2_126_3477_U453 ( .A(DP_OP_424J2_126_3477_n2317), .B(
        DP_OP_424J2_126_3477_n2982), .CI(DP_OP_424J2_126_3477_n2632), .CO(
        DP_OP_424J2_126_3477_n592), .S(DP_OP_424J2_126_3477_n593) );
  FADDX1_HVT DP_OP_424J2_126_3477_U452 ( .A(DP_OP_424J2_126_3477_n2009), .B(
        DP_OP_424J2_126_3477_n2544), .CI(DP_OP_424J2_126_3477_n2764), .CO(
        DP_OP_424J2_126_3477_n590), .S(DP_OP_424J2_126_3477_n591) );
  FADDX1_HVT DP_OP_424J2_126_3477_U451 ( .A(DP_OP_424J2_126_3477_n2229), .B(
        DP_OP_424J2_126_3477_n2324), .CI(DP_OP_424J2_126_3477_n2940), .CO(
        DP_OP_424J2_126_3477_n588), .S(DP_OP_424J2_126_3477_n589) );
  FADDX1_HVT DP_OP_424J2_126_3477_U450 ( .A(DP_OP_424J2_126_3477_n1965), .B(
        DP_OP_424J2_126_3477_n2852), .CI(DP_OP_424J2_126_3477_n2016), .CO(
        DP_OP_424J2_126_3477_n586), .S(DP_OP_424J2_126_3477_n587) );
  FADDX1_HVT DP_OP_424J2_126_3477_U449 ( .A(DP_OP_424J2_126_3477_n2097), .B(
        DP_OP_424J2_126_3477_n1972), .CI(DP_OP_424J2_126_3477_n2808), .CO(
        DP_OP_424J2_126_3477_n584), .S(DP_OP_424J2_126_3477_n585) );
  FADDX1_HVT DP_OP_424J2_126_3477_U448 ( .A(DP_OP_424J2_126_3477_n2933), .B(
        DP_OP_424J2_126_3477_n2368), .CI(DP_OP_424J2_126_3477_n2456), .CO(
        DP_OP_424J2_126_3477_n582), .S(DP_OP_424J2_126_3477_n583) );
  FADDX1_HVT DP_OP_424J2_126_3477_U447 ( .A(DP_OP_424J2_126_3477_n2449), .B(
        DP_OP_424J2_126_3477_n2500), .CI(DP_OP_424J2_126_3477_n2896), .CO(
        DP_OP_424J2_126_3477_n580), .S(DP_OP_424J2_126_3477_n581) );
  FADDX1_HVT DP_OP_424J2_126_3477_U446 ( .A(DP_OP_424J2_126_3477_n2713), .B(
        DP_OP_424J2_126_3477_n2192), .CI(DP_OP_424J2_126_3477_n2720), .CO(
        DP_OP_424J2_126_3477_n578), .S(DP_OP_424J2_126_3477_n579) );
  FADDX1_HVT DP_OP_424J2_126_3477_U445 ( .A(DP_OP_424J2_126_3477_n2889), .B(
        DP_OP_424J2_126_3477_n2412), .CI(DP_OP_424J2_126_3477_n2588), .CO(
        DP_OP_424J2_126_3477_n576), .S(DP_OP_424J2_126_3477_n577) );
  FADDX1_HVT DP_OP_424J2_126_3477_U444 ( .A(DP_OP_424J2_126_3477_n2185), .B(
        DP_OP_424J2_126_3477_n2060), .CI(DP_OP_424J2_126_3477_n2676), .CO(
        DP_OP_424J2_126_3477_n574), .S(DP_OP_424J2_126_3477_n575) );
  FADDX1_HVT DP_OP_424J2_126_3477_U443 ( .A(DP_OP_424J2_126_3477_n2141), .B(
        DP_OP_424J2_126_3477_n2280), .CI(DP_OP_424J2_126_3477_n2148), .CO(
        DP_OP_424J2_126_3477_n572), .S(DP_OP_424J2_126_3477_n573) );
  FADDX1_HVT DP_OP_424J2_126_3477_U442 ( .A(DP_OP_424J2_126_3477_n2537), .B(
        DP_OP_424J2_126_3477_n2361), .CI(DP_OP_424J2_126_3477_n2104), .CO(
        DP_OP_424J2_126_3477_n570), .S(DP_OP_424J2_126_3477_n571) );
  FADDX1_HVT DP_OP_424J2_126_3477_U441 ( .A(DP_OP_424J2_126_3477_n2845), .B(
        DP_OP_424J2_126_3477_n2053), .CI(DP_OP_424J2_126_3477_n2273), .CO(
        DP_OP_424J2_126_3477_n568), .S(DP_OP_424J2_126_3477_n569) );
  FADDX1_HVT DP_OP_424J2_126_3477_U440 ( .A(DP_OP_424J2_126_3477_n2801), .B(
        DP_OP_424J2_126_3477_n2405), .CI(DP_OP_424J2_126_3477_n2493), .CO(
        DP_OP_424J2_126_3477_n566), .S(DP_OP_424J2_126_3477_n567) );
  FADDX1_HVT DP_OP_424J2_126_3477_U439 ( .A(DP_OP_424J2_126_3477_n2757), .B(
        DP_OP_424J2_126_3477_n2581), .CI(DP_OP_424J2_126_3477_n2625), .CO(
        DP_OP_424J2_126_3477_n564), .S(DP_OP_424J2_126_3477_n565) );
  FADDX1_HVT DP_OP_424J2_126_3477_U438 ( .A(DP_OP_424J2_126_3477_n2669), .B(
        DP_OP_424J2_126_3477_n768), .CI(DP_OP_424J2_126_3477_n766), .CO(
        DP_OP_424J2_126_3477_n562), .S(DP_OP_424J2_126_3477_n563) );
  FADDX1_HVT DP_OP_424J2_126_3477_U437 ( .A(DP_OP_424J2_126_3477_n764), .B(
        DP_OP_424J2_126_3477_n736), .CI(DP_OP_424J2_126_3477_n738), .CO(
        DP_OP_424J2_126_3477_n560), .S(DP_OP_424J2_126_3477_n561) );
  FADDX1_HVT DP_OP_424J2_126_3477_U436 ( .A(DP_OP_424J2_126_3477_n762), .B(
        DP_OP_424J2_126_3477_n740), .CI(DP_OP_424J2_126_3477_n742), .CO(
        DP_OP_424J2_126_3477_n558), .S(DP_OP_424J2_126_3477_n559) );
  FADDX1_HVT DP_OP_424J2_126_3477_U435 ( .A(DP_OP_424J2_126_3477_n760), .B(
        DP_OP_424J2_126_3477_n744), .CI(DP_OP_424J2_126_3477_n746), .CO(
        DP_OP_424J2_126_3477_n556), .S(DP_OP_424J2_126_3477_n557) );
  FADDX1_HVT DP_OP_424J2_126_3477_U434 ( .A(DP_OP_424J2_126_3477_n758), .B(
        DP_OP_424J2_126_3477_n748), .CI(DP_OP_424J2_126_3477_n750), .CO(
        DP_OP_424J2_126_3477_n554), .S(DP_OP_424J2_126_3477_n555) );
  FADDX1_HVT DP_OP_424J2_126_3477_U433 ( .A(DP_OP_424J2_126_3477_n756), .B(
        DP_OP_424J2_126_3477_n752), .CI(DP_OP_424J2_126_3477_n754), .CO(
        DP_OP_424J2_126_3477_n552), .S(DP_OP_424J2_126_3477_n553) );
  FADDX1_HVT DP_OP_424J2_126_3477_U432 ( .A(DP_OP_424J2_126_3477_n734), .B(
        DP_OP_424J2_126_3477_n720), .CI(DP_OP_424J2_126_3477_n732), .CO(
        DP_OP_424J2_126_3477_n550), .S(DP_OP_424J2_126_3477_n551) );
  FADDX1_HVT DP_OP_424J2_126_3477_U431 ( .A(DP_OP_424J2_126_3477_n726), .B(
        DP_OP_424J2_126_3477_n722), .CI(DP_OP_424J2_126_3477_n724), .CO(
        DP_OP_424J2_126_3477_n548), .S(DP_OP_424J2_126_3477_n549) );
  FADDX1_HVT DP_OP_424J2_126_3477_U430 ( .A(DP_OP_424J2_126_3477_n730), .B(
        DP_OP_424J2_126_3477_n728), .CI(DP_OP_424J2_126_3477_n595), .CO(
        DP_OP_424J2_126_3477_n546), .S(DP_OP_424J2_126_3477_n547) );
  FADDX1_HVT DP_OP_424J2_126_3477_U429 ( .A(DP_OP_424J2_126_3477_n597), .B(
        DP_OP_424J2_126_3477_n583), .CI(DP_OP_424J2_126_3477_n589), .CO(
        DP_OP_424J2_126_3477_n544), .S(DP_OP_424J2_126_3477_n545) );
  FADDX1_HVT DP_OP_424J2_126_3477_U428 ( .A(DP_OP_424J2_126_3477_n565), .B(
        DP_OP_424J2_126_3477_n587), .CI(DP_OP_424J2_126_3477_n585), .CO(
        DP_OP_424J2_126_3477_n542), .S(DP_OP_424J2_126_3477_n543) );
  FADDX1_HVT DP_OP_424J2_126_3477_U427 ( .A(DP_OP_424J2_126_3477_n591), .B(
        DP_OP_424J2_126_3477_n573), .CI(DP_OP_424J2_126_3477_n575), .CO(
        DP_OP_424J2_126_3477_n540), .S(DP_OP_424J2_126_3477_n541) );
  FADDX1_HVT DP_OP_424J2_126_3477_U426 ( .A(DP_OP_424J2_126_3477_n577), .B(
        DP_OP_424J2_126_3477_n567), .CI(DP_OP_424J2_126_3477_n569), .CO(
        DP_OP_424J2_126_3477_n538), .S(DP_OP_424J2_126_3477_n539) );
  FADDX1_HVT DP_OP_424J2_126_3477_U425 ( .A(DP_OP_424J2_126_3477_n571), .B(
        DP_OP_424J2_126_3477_n593), .CI(DP_OP_424J2_126_3477_n581), .CO(
        DP_OP_424J2_126_3477_n536), .S(DP_OP_424J2_126_3477_n537) );
  FADDX1_HVT DP_OP_424J2_126_3477_U424 ( .A(DP_OP_424J2_126_3477_n579), .B(
        DP_OP_424J2_126_3477_n718), .CI(DP_OP_424J2_126_3477_n716), .CO(
        DP_OP_424J2_126_3477_n534), .S(DP_OP_424J2_126_3477_n535) );
  FADDX1_HVT DP_OP_424J2_126_3477_U423 ( .A(DP_OP_424J2_126_3477_n714), .B(
        DP_OP_424J2_126_3477_n708), .CI(DP_OP_424J2_126_3477_n710), .CO(
        DP_OP_424J2_126_3477_n532), .S(DP_OP_424J2_126_3477_n533) );
  FADDX1_HVT DP_OP_424J2_126_3477_U422 ( .A(DP_OP_424J2_126_3477_n712), .B(
        DP_OP_424J2_126_3477_n706), .CI(DP_OP_424J2_126_3477_n704), .CO(
        DP_OP_424J2_126_3477_n530), .S(DP_OP_424J2_126_3477_n531) );
  FADDX1_HVT DP_OP_424J2_126_3477_U421 ( .A(DP_OP_424J2_126_3477_n702), .B(
        DP_OP_424J2_126_3477_n698), .CI(DP_OP_424J2_126_3477_n696), .CO(
        DP_OP_424J2_126_3477_n528), .S(DP_OP_424J2_126_3477_n529) );
  FADDX1_HVT DP_OP_424J2_126_3477_U420 ( .A(DP_OP_424J2_126_3477_n700), .B(
        DP_OP_424J2_126_3477_n563), .CI(DP_OP_424J2_126_3477_n557), .CO(
        DP_OP_424J2_126_3477_n526), .S(DP_OP_424J2_126_3477_n527) );
  FADDX1_HVT DP_OP_424J2_126_3477_U419 ( .A(DP_OP_424J2_126_3477_n559), .B(
        DP_OP_424J2_126_3477_n553), .CI(DP_OP_424J2_126_3477_n684), .CO(
        DP_OP_424J2_126_3477_n524), .S(DP_OP_424J2_126_3477_n525) );
  FADDX1_HVT DP_OP_424J2_126_3477_U418 ( .A(DP_OP_424J2_126_3477_n694), .B(
        DP_OP_424J2_126_3477_n561), .CI(DP_OP_424J2_126_3477_n555), .CO(
        DP_OP_424J2_126_3477_n522), .S(DP_OP_424J2_126_3477_n523) );
  FADDX1_HVT DP_OP_424J2_126_3477_U417 ( .A(DP_OP_424J2_126_3477_n688), .B(
        DP_OP_424J2_126_3477_n692), .CI(DP_OP_424J2_126_3477_n686), .CO(
        DP_OP_424J2_126_3477_n520), .S(DP_OP_424J2_126_3477_n521) );
  FADDX1_HVT DP_OP_424J2_126_3477_U416 ( .A(DP_OP_424J2_126_3477_n690), .B(
        DP_OP_424J2_126_3477_n682), .CI(DP_OP_424J2_126_3477_n680), .CO(
        DP_OP_424J2_126_3477_n518), .S(DP_OP_424J2_126_3477_n519) );
  FADDX1_HVT DP_OP_424J2_126_3477_U415 ( .A(DP_OP_424J2_126_3477_n549), .B(
        DP_OP_424J2_126_3477_n551), .CI(DP_OP_424J2_126_3477_n547), .CO(
        DP_OP_424J2_126_3477_n516), .S(DP_OP_424J2_126_3477_n517) );
  FADDX1_HVT DP_OP_424J2_126_3477_U414 ( .A(DP_OP_424J2_126_3477_n545), .B(
        DP_OP_424J2_126_3477_n539), .CI(DP_OP_424J2_126_3477_n543), .CO(
        DP_OP_424J2_126_3477_n514), .S(DP_OP_424J2_126_3477_n515) );
  FADDX1_HVT DP_OP_424J2_126_3477_U413 ( .A(DP_OP_424J2_126_3477_n537), .B(
        DP_OP_424J2_126_3477_n541), .CI(DP_OP_424J2_126_3477_n678), .CO(
        DP_OP_424J2_126_3477_n512), .S(DP_OP_424J2_126_3477_n513) );
  FADDX1_HVT DP_OP_424J2_126_3477_U412 ( .A(DP_OP_424J2_126_3477_n676), .B(
        DP_OP_424J2_126_3477_n672), .CI(DP_OP_424J2_126_3477_n535), .CO(
        DP_OP_424J2_126_3477_n510), .S(DP_OP_424J2_126_3477_n511) );
  FADDX1_HVT DP_OP_424J2_126_3477_U411 ( .A(DP_OP_424J2_126_3477_n674), .B(
        DP_OP_424J2_126_3477_n670), .CI(DP_OP_424J2_126_3477_n668), .CO(
        DP_OP_424J2_126_3477_n508), .S(DP_OP_424J2_126_3477_n509) );
  FADDX1_HVT DP_OP_424J2_126_3477_U410 ( .A(DP_OP_424J2_126_3477_n666), .B(
        DP_OP_424J2_126_3477_n533), .CI(DP_OP_424J2_126_3477_n531), .CO(
        DP_OP_424J2_126_3477_n506), .S(DP_OP_424J2_126_3477_n507) );
  FADDX1_HVT DP_OP_424J2_126_3477_U409 ( .A(DP_OP_424J2_126_3477_n664), .B(
        DP_OP_424J2_126_3477_n662), .CI(DP_OP_424J2_126_3477_n660), .CO(
        DP_OP_424J2_126_3477_n504), .S(DP_OP_424J2_126_3477_n505) );
  FADDX1_HVT DP_OP_424J2_126_3477_U408 ( .A(DP_OP_424J2_126_3477_n658), .B(
        DP_OP_424J2_126_3477_n529), .CI(DP_OP_424J2_126_3477_n656), .CO(
        DP_OP_424J2_126_3477_n502), .S(DP_OP_424J2_126_3477_n503) );
  FADDX1_HVT DP_OP_424J2_126_3477_U407 ( .A(DP_OP_424J2_126_3477_n527), .B(
        DP_OP_424J2_126_3477_n654), .CI(DP_OP_424J2_126_3477_n525), .CO(
        DP_OP_424J2_126_3477_n500), .S(DP_OP_424J2_126_3477_n501) );
  FADDX1_HVT DP_OP_424J2_126_3477_U406 ( .A(DP_OP_424J2_126_3477_n652), .B(
        DP_OP_424J2_126_3477_n521), .CI(DP_OP_424J2_126_3477_n519), .CO(
        DP_OP_424J2_126_3477_n498), .S(DP_OP_424J2_126_3477_n499) );
  FADDX1_HVT DP_OP_424J2_126_3477_U405 ( .A(DP_OP_424J2_126_3477_n523), .B(
        DP_OP_424J2_126_3477_n517), .CI(DP_OP_424J2_126_3477_n650), .CO(
        DP_OP_424J2_126_3477_n496), .S(DP_OP_424J2_126_3477_n497) );
  FADDX1_HVT DP_OP_424J2_126_3477_U404 ( .A(DP_OP_424J2_126_3477_n515), .B(
        DP_OP_424J2_126_3477_n648), .CI(DP_OP_424J2_126_3477_n513), .CO(
        DP_OP_424J2_126_3477_n494), .S(DP_OP_424J2_126_3477_n495) );
  FADDX1_HVT DP_OP_424J2_126_3477_U403 ( .A(DP_OP_424J2_126_3477_n646), .B(
        DP_OP_424J2_126_3477_n644), .CI(DP_OP_424J2_126_3477_n642), .CO(
        DP_OP_424J2_126_3477_n492), .S(DP_OP_424J2_126_3477_n493) );
  FADDX1_HVT DP_OP_424J2_126_3477_U402 ( .A(DP_OP_424J2_126_3477_n511), .B(
        DP_OP_424J2_126_3477_n640), .CI(DP_OP_424J2_126_3477_n509), .CO(
        DP_OP_424J2_126_3477_n490), .S(DP_OP_424J2_126_3477_n491) );
  FADDX1_HVT DP_OP_424J2_126_3477_U401 ( .A(DP_OP_424J2_126_3477_n638), .B(
        DP_OP_424J2_126_3477_n507), .CI(DP_OP_424J2_126_3477_n505), .CO(
        DP_OP_424J2_126_3477_n488), .S(DP_OP_424J2_126_3477_n489) );
  FADDX1_HVT DP_OP_424J2_126_3477_U400 ( .A(DP_OP_424J2_126_3477_n636), .B(
        DP_OP_424J2_126_3477_n634), .CI(DP_OP_424J2_126_3477_n503), .CO(
        DP_OP_424J2_126_3477_n486), .S(DP_OP_424J2_126_3477_n487) );
  FADDX1_HVT DP_OP_424J2_126_3477_U399 ( .A(DP_OP_424J2_126_3477_n632), .B(
        DP_OP_424J2_126_3477_n501), .CI(DP_OP_424J2_126_3477_n499), .CO(
        DP_OP_424J2_126_3477_n484), .S(DP_OP_424J2_126_3477_n485) );
  FADDX1_HVT DP_OP_424J2_126_3477_U398 ( .A(DP_OP_424J2_126_3477_n630), .B(
        DP_OP_424J2_126_3477_n497), .CI(DP_OP_424J2_126_3477_n628), .CO(
        DP_OP_424J2_126_3477_n482), .S(DP_OP_424J2_126_3477_n483) );
  FADDX1_HVT DP_OP_424J2_126_3477_U397 ( .A(DP_OP_424J2_126_3477_n495), .B(
        DP_OP_424J2_126_3477_n626), .CI(DP_OP_424J2_126_3477_n493), .CO(
        DP_OP_424J2_126_3477_n480), .S(DP_OP_424J2_126_3477_n481) );
  FADDX1_HVT DP_OP_424J2_126_3477_U396 ( .A(DP_OP_424J2_126_3477_n624), .B(
        DP_OP_424J2_126_3477_n622), .CI(DP_OP_424J2_126_3477_n491), .CO(
        DP_OP_424J2_126_3477_n478), .S(DP_OP_424J2_126_3477_n479) );
  FADDX1_HVT DP_OP_424J2_126_3477_U395 ( .A(DP_OP_424J2_126_3477_n620), .B(
        DP_OP_424J2_126_3477_n489), .CI(DP_OP_424J2_126_3477_n487), .CO(
        DP_OP_424J2_126_3477_n476), .S(DP_OP_424J2_126_3477_n477) );
  FADDX1_HVT DP_OP_424J2_126_3477_U394 ( .A(DP_OP_424J2_126_3477_n618), .B(
        DP_OP_424J2_126_3477_n485), .CI(DP_OP_424J2_126_3477_n616), .CO(
        DP_OP_424J2_126_3477_n474), .S(DP_OP_424J2_126_3477_n475) );
  FADDX1_HVT DP_OP_424J2_126_3477_U393 ( .A(DP_OP_424J2_126_3477_n483), .B(
        DP_OP_424J2_126_3477_n614), .CI(DP_OP_424J2_126_3477_n481), .CO(
        DP_OP_424J2_126_3477_n472), .S(DP_OP_424J2_126_3477_n473) );
  FADDX1_HVT DP_OP_424J2_126_3477_U392 ( .A(DP_OP_424J2_126_3477_n612), .B(
        DP_OP_424J2_126_3477_n479), .CI(DP_OP_424J2_126_3477_n610), .CO(
        DP_OP_424J2_126_3477_n470), .S(DP_OP_424J2_126_3477_n471) );
  FADDX1_HVT DP_OP_424J2_126_3477_U391 ( .A(DP_OP_424J2_126_3477_n477), .B(
        DP_OP_424J2_126_3477_n608), .CI(DP_OP_424J2_126_3477_n475), .CO(
        DP_OP_424J2_126_3477_n468), .S(DP_OP_424J2_126_3477_n469) );
  FADDX1_HVT DP_OP_424J2_126_3477_U390 ( .A(DP_OP_424J2_126_3477_n606), .B(
        DP_OP_424J2_126_3477_n473), .CI(DP_OP_424J2_126_3477_n604), .CO(
        DP_OP_424J2_126_3477_n466), .S(DP_OP_424J2_126_3477_n467) );
  FADDX1_HVT DP_OP_424J2_126_3477_U389 ( .A(DP_OP_424J2_126_3477_n471), .B(
        DP_OP_424J2_126_3477_n469), .CI(DP_OP_424J2_126_3477_n602), .CO(
        DP_OP_424J2_126_3477_n464), .S(DP_OP_424J2_126_3477_n465) );
  FADDX1_HVT DP_OP_424J2_126_3477_U388 ( .A(DP_OP_424J2_126_3477_n600), .B(
        DP_OP_424J2_126_3477_n467), .CI(DP_OP_424J2_126_3477_n465), .CO(
        DP_OP_424J2_126_3477_n462), .S(DP_OP_424J2_126_3477_n463) );
  FADDX1_HVT DP_OP_424J2_126_3477_U386 ( .A(DP_OP_424J2_126_3477_n2976), .B(
        DP_OP_424J2_126_3477_n1920), .CI(DP_OP_424J2_126_3477_n461), .CO(
        DP_OP_424J2_126_3477_n458), .S(DP_OP_424J2_126_3477_n459) );
  FADDX1_HVT DP_OP_424J2_126_3477_U385 ( .A(DP_OP_424J2_126_3477_n2008), .B(
        DP_OP_424J2_126_3477_n2932), .CI(DP_OP_424J2_126_3477_n2360), .CO(
        DP_OP_424J2_126_3477_n456), .S(DP_OP_424J2_126_3477_n457) );
  FADDX1_HVT DP_OP_424J2_126_3477_U384 ( .A(DP_OP_424J2_126_3477_n2492), .B(
        DP_OP_424J2_126_3477_n2888), .CI(DP_OP_424J2_126_3477_n2844), .CO(
        DP_OP_424J2_126_3477_n454), .S(DP_OP_424J2_126_3477_n455) );
  FADDX1_HVT DP_OP_424J2_126_3477_U383 ( .A(DP_OP_424J2_126_3477_n2316), .B(
        DP_OP_424J2_126_3477_n2800), .CI(DP_OP_424J2_126_3477_n2756), .CO(
        DP_OP_424J2_126_3477_n452), .S(DP_OP_424J2_126_3477_n453) );
  FADDX1_HVT DP_OP_424J2_126_3477_U382 ( .A(DP_OP_424J2_126_3477_n2184), .B(
        DP_OP_424J2_126_3477_n1964), .CI(DP_OP_424J2_126_3477_n2712), .CO(
        DP_OP_424J2_126_3477_n450), .S(DP_OP_424J2_126_3477_n451) );
  FADDX1_HVT DP_OP_424J2_126_3477_U381 ( .A(DP_OP_424J2_126_3477_n2668), .B(
        DP_OP_424J2_126_3477_n2624), .CI(DP_OP_424J2_126_3477_n2580), .CO(
        DP_OP_424J2_126_3477_n448), .S(DP_OP_424J2_126_3477_n449) );
  FADDX1_HVT DP_OP_424J2_126_3477_U380 ( .A(DP_OP_424J2_126_3477_n2228), .B(
        DP_OP_424J2_126_3477_n2052), .CI(DP_OP_424J2_126_3477_n2096), .CO(
        DP_OP_424J2_126_3477_n446), .S(DP_OP_424J2_126_3477_n447) );
  FADDX1_HVT DP_OP_424J2_126_3477_U379 ( .A(DP_OP_424J2_126_3477_n2140), .B(
        DP_OP_424J2_126_3477_n2536), .CI(DP_OP_424J2_126_3477_n2448), .CO(
        DP_OP_424J2_126_3477_n444), .S(DP_OP_424J2_126_3477_n445) );
  FADDX1_HVT DP_OP_424J2_126_3477_U378 ( .A(DP_OP_424J2_126_3477_n2272), .B(
        DP_OP_424J2_126_3477_n2404), .CI(DP_OP_424J2_126_3477_n596), .CO(
        DP_OP_424J2_126_3477_n442), .S(DP_OP_424J2_126_3477_n443) );
  FADDX1_HVT DP_OP_424J2_126_3477_U377 ( .A(DP_OP_424J2_126_3477_n594), .B(
        DP_OP_424J2_126_3477_n564), .CI(DP_OP_424J2_126_3477_n592), .CO(
        DP_OP_424J2_126_3477_n440), .S(DP_OP_424J2_126_3477_n441) );
  FADDX1_HVT DP_OP_424J2_126_3477_U376 ( .A(DP_OP_424J2_126_3477_n590), .B(
        DP_OP_424J2_126_3477_n566), .CI(DP_OP_424J2_126_3477_n568), .CO(
        DP_OP_424J2_126_3477_n438), .S(DP_OP_424J2_126_3477_n439) );
  FADDX1_HVT DP_OP_424J2_126_3477_U375 ( .A(DP_OP_424J2_126_3477_n588), .B(
        DP_OP_424J2_126_3477_n570), .CI(DP_OP_424J2_126_3477_n572), .CO(
        DP_OP_424J2_126_3477_n436), .S(DP_OP_424J2_126_3477_n437) );
  FADDX1_HVT DP_OP_424J2_126_3477_U374 ( .A(DP_OP_424J2_126_3477_n586), .B(
        DP_OP_424J2_126_3477_n574), .CI(DP_OP_424J2_126_3477_n576), .CO(
        DP_OP_424J2_126_3477_n434), .S(DP_OP_424J2_126_3477_n435) );
  FADDX1_HVT DP_OP_424J2_126_3477_U373 ( .A(DP_OP_424J2_126_3477_n584), .B(
        DP_OP_424J2_126_3477_n578), .CI(DP_OP_424J2_126_3477_n580), .CO(
        DP_OP_424J2_126_3477_n432), .S(DP_OP_424J2_126_3477_n433) );
  FADDX1_HVT DP_OP_424J2_126_3477_U372 ( .A(DP_OP_424J2_126_3477_n582), .B(
        DP_OP_424J2_126_3477_n459), .CI(DP_OP_424J2_126_3477_n455), .CO(
        DP_OP_424J2_126_3477_n430), .S(DP_OP_424J2_126_3477_n431) );
  FADDX1_HVT DP_OP_424J2_126_3477_U371 ( .A(DP_OP_424J2_126_3477_n451), .B(
        DP_OP_424J2_126_3477_n445), .CI(DP_OP_424J2_126_3477_n447), .CO(
        DP_OP_424J2_126_3477_n428), .S(DP_OP_424J2_126_3477_n429) );
  FADDX1_HVT DP_OP_424J2_126_3477_U370 ( .A(DP_OP_424J2_126_3477_n449), .B(
        DP_OP_424J2_126_3477_n457), .CI(DP_OP_424J2_126_3477_n453), .CO(
        DP_OP_424J2_126_3477_n426), .S(DP_OP_424J2_126_3477_n427) );
  FADDX1_HVT DP_OP_424J2_126_3477_U369 ( .A(DP_OP_424J2_126_3477_n562), .B(
        DP_OP_424J2_126_3477_n560), .CI(DP_OP_424J2_126_3477_n552), .CO(
        DP_OP_424J2_126_3477_n424), .S(DP_OP_424J2_126_3477_n425) );
  FADDX1_HVT DP_OP_424J2_126_3477_U368 ( .A(DP_OP_424J2_126_3477_n558), .B(
        DP_OP_424J2_126_3477_n554), .CI(DP_OP_424J2_126_3477_n556), .CO(
        DP_OP_424J2_126_3477_n422), .S(DP_OP_424J2_126_3477_n423) );
  FADDX1_HVT DP_OP_424J2_126_3477_U367 ( .A(DP_OP_424J2_126_3477_n550), .B(
        DP_OP_424J2_126_3477_n546), .CI(DP_OP_424J2_126_3477_n443), .CO(
        DP_OP_424J2_126_3477_n420), .S(DP_OP_424J2_126_3477_n421) );
  FADDX1_HVT DP_OP_424J2_126_3477_U366 ( .A(DP_OP_424J2_126_3477_n548), .B(
        DP_OP_424J2_126_3477_n544), .CI(DP_OP_424J2_126_3477_n441), .CO(
        DP_OP_424J2_126_3477_n418), .S(DP_OP_424J2_126_3477_n419) );
  FADDX1_HVT DP_OP_424J2_126_3477_U365 ( .A(DP_OP_424J2_126_3477_n542), .B(
        DP_OP_424J2_126_3477_n435), .CI(DP_OP_424J2_126_3477_n437), .CO(
        DP_OP_424J2_126_3477_n416), .S(DP_OP_424J2_126_3477_n417) );
  FADDX1_HVT DP_OP_424J2_126_3477_U364 ( .A(DP_OP_424J2_126_3477_n540), .B(
        DP_OP_424J2_126_3477_n439), .CI(DP_OP_424J2_126_3477_n433), .CO(
        DP_OP_424J2_126_3477_n414), .S(DP_OP_424J2_126_3477_n415) );
  FADDX1_HVT DP_OP_424J2_126_3477_U363 ( .A(DP_OP_424J2_126_3477_n538), .B(
        DP_OP_424J2_126_3477_n536), .CI(DP_OP_424J2_126_3477_n534), .CO(
        DP_OP_424J2_126_3477_n412), .S(DP_OP_424J2_126_3477_n413) );
  FADDX1_HVT DP_OP_424J2_126_3477_U362 ( .A(DP_OP_424J2_126_3477_n431), .B(
        DP_OP_424J2_126_3477_n427), .CI(DP_OP_424J2_126_3477_n532), .CO(
        DP_OP_424J2_126_3477_n410), .S(DP_OP_424J2_126_3477_n411) );
  FADDX1_HVT DP_OP_424J2_126_3477_U361 ( .A(DP_OP_424J2_126_3477_n429), .B(
        DP_OP_424J2_126_3477_n530), .CI(DP_OP_424J2_126_3477_n528), .CO(
        DP_OP_424J2_126_3477_n408), .S(DP_OP_424J2_126_3477_n409) );
  FADDX1_HVT DP_OP_424J2_126_3477_U360 ( .A(DP_OP_424J2_126_3477_n526), .B(
        DP_OP_424J2_126_3477_n425), .CI(DP_OP_424J2_126_3477_n423), .CO(
        DP_OP_424J2_126_3477_n406), .S(DP_OP_424J2_126_3477_n407) );
  FADDX1_HVT DP_OP_424J2_126_3477_U359 ( .A(DP_OP_424J2_126_3477_n524), .B(
        DP_OP_424J2_126_3477_n520), .CI(DP_OP_424J2_126_3477_n518), .CO(
        DP_OP_424J2_126_3477_n404), .S(DP_OP_424J2_126_3477_n405) );
  FADDX1_HVT DP_OP_424J2_126_3477_U358 ( .A(DP_OP_424J2_126_3477_n522), .B(
        DP_OP_424J2_126_3477_n516), .CI(DP_OP_424J2_126_3477_n421), .CO(
        DP_OP_424J2_126_3477_n402), .S(DP_OP_424J2_126_3477_n403) );
  FADDX1_HVT DP_OP_424J2_126_3477_U357 ( .A(DP_OP_424J2_126_3477_n419), .B(
        DP_OP_424J2_126_3477_n514), .CI(DP_OP_424J2_126_3477_n512), .CO(
        DP_OP_424J2_126_3477_n400), .S(DP_OP_424J2_126_3477_n401) );
  FADDX1_HVT DP_OP_424J2_126_3477_U356 ( .A(DP_OP_424J2_126_3477_n417), .B(
        DP_OP_424J2_126_3477_n415), .CI(DP_OP_424J2_126_3477_n413), .CO(
        DP_OP_424J2_126_3477_n398), .S(DP_OP_424J2_126_3477_n399) );
  FADDX1_HVT DP_OP_424J2_126_3477_U355 ( .A(DP_OP_424J2_126_3477_n510), .B(
        DP_OP_424J2_126_3477_n508), .CI(DP_OP_424J2_126_3477_n411), .CO(
        DP_OP_424J2_126_3477_n396), .S(DP_OP_424J2_126_3477_n397) );
  FADDX1_HVT DP_OP_424J2_126_3477_U354 ( .A(DP_OP_424J2_126_3477_n506), .B(
        DP_OP_424J2_126_3477_n409), .CI(DP_OP_424J2_126_3477_n504), .CO(
        DP_OP_424J2_126_3477_n394), .S(DP_OP_424J2_126_3477_n395) );
  FADDX1_HVT DP_OP_424J2_126_3477_U353 ( .A(DP_OP_424J2_126_3477_n502), .B(
        DP_OP_424J2_126_3477_n407), .CI(DP_OP_424J2_126_3477_n500), .CO(
        DP_OP_424J2_126_3477_n392), .S(DP_OP_424J2_126_3477_n393) );
  FADDX1_HVT DP_OP_424J2_126_3477_U352 ( .A(DP_OP_424J2_126_3477_n498), .B(
        DP_OP_424J2_126_3477_n405), .CI(DP_OP_424J2_126_3477_n403), .CO(
        DP_OP_424J2_126_3477_n390), .S(DP_OP_424J2_126_3477_n391) );
  FADDX1_HVT DP_OP_424J2_126_3477_U351 ( .A(DP_OP_424J2_126_3477_n496), .B(
        DP_OP_424J2_126_3477_n401), .CI(DP_OP_424J2_126_3477_n494), .CO(
        DP_OP_424J2_126_3477_n388), .S(DP_OP_424J2_126_3477_n389) );
  FADDX1_HVT DP_OP_424J2_126_3477_U350 ( .A(DP_OP_424J2_126_3477_n399), .B(
        DP_OP_424J2_126_3477_n492), .CI(DP_OP_424J2_126_3477_n490), .CO(
        DP_OP_424J2_126_3477_n386), .S(DP_OP_424J2_126_3477_n387) );
  FADDX1_HVT DP_OP_424J2_126_3477_U349 ( .A(DP_OP_424J2_126_3477_n397), .B(
        DP_OP_424J2_126_3477_n488), .CI(DP_OP_424J2_126_3477_n395), .CO(
        DP_OP_424J2_126_3477_n384), .S(DP_OP_424J2_126_3477_n385) );
  FADDX1_HVT DP_OP_424J2_126_3477_U348 ( .A(DP_OP_424J2_126_3477_n486), .B(
        DP_OP_424J2_126_3477_n393), .CI(DP_OP_424J2_126_3477_n484), .CO(
        DP_OP_424J2_126_3477_n382), .S(DP_OP_424J2_126_3477_n383) );
  FADDX1_HVT DP_OP_424J2_126_3477_U347 ( .A(DP_OP_424J2_126_3477_n391), .B(
        DP_OP_424J2_126_3477_n482), .CI(DP_OP_424J2_126_3477_n389), .CO(
        DP_OP_424J2_126_3477_n380), .S(DP_OP_424J2_126_3477_n381) );
  FADDX1_HVT DP_OP_424J2_126_3477_U346 ( .A(DP_OP_424J2_126_3477_n480), .B(
        DP_OP_424J2_126_3477_n387), .CI(DP_OP_424J2_126_3477_n478), .CO(
        DP_OP_424J2_126_3477_n378), .S(DP_OP_424J2_126_3477_n379) );
  FADDX1_HVT DP_OP_424J2_126_3477_U345 ( .A(DP_OP_424J2_126_3477_n385), .B(
        DP_OP_424J2_126_3477_n476), .CI(DP_OP_424J2_126_3477_n383), .CO(
        DP_OP_424J2_126_3477_n376), .S(DP_OP_424J2_126_3477_n377) );
  FADDX1_HVT DP_OP_424J2_126_3477_U344 ( .A(DP_OP_424J2_126_3477_n474), .B(
        DP_OP_424J2_126_3477_n381), .CI(DP_OP_424J2_126_3477_n472), .CO(
        DP_OP_424J2_126_3477_n374), .S(DP_OP_424J2_126_3477_n375) );
  FADDX1_HVT DP_OP_424J2_126_3477_U343 ( .A(DP_OP_424J2_126_3477_n379), .B(
        DP_OP_424J2_126_3477_n470), .CI(DP_OP_424J2_126_3477_n377), .CO(
        DP_OP_424J2_126_3477_n372), .S(DP_OP_424J2_126_3477_n373) );
  FADDX1_HVT DP_OP_424J2_126_3477_U342 ( .A(DP_OP_424J2_126_3477_n468), .B(
        DP_OP_424J2_126_3477_n375), .CI(DP_OP_424J2_126_3477_n466), .CO(
        DP_OP_424J2_126_3477_n370), .S(DP_OP_424J2_126_3477_n371) );
  FADDX1_HVT DP_OP_424J2_126_3477_U341 ( .A(DP_OP_424J2_126_3477_n373), .B(
        DP_OP_424J2_126_3477_n464), .CI(DP_OP_424J2_126_3477_n371), .CO(
        DP_OP_424J2_126_3477_n368), .S(DP_OP_424J2_126_3477_n369) );
  FADDX1_HVT DP_OP_424J2_126_3477_U340 ( .A(DP_OP_424J2_126_3477_n1876), .B(
        DP_OP_424J2_126_3477_n460), .CI(DP_OP_424J2_126_3477_n458), .CO(
        DP_OP_424J2_126_3477_n366), .S(DP_OP_424J2_126_3477_n367) );
  FADDX1_HVT DP_OP_424J2_126_3477_U339 ( .A(DP_OP_424J2_126_3477_n448), .B(
        DP_OP_424J2_126_3477_n444), .CI(DP_OP_424J2_126_3477_n456), .CO(
        DP_OP_424J2_126_3477_n364), .S(DP_OP_424J2_126_3477_n365) );
  FADDX1_HVT DP_OP_424J2_126_3477_U338 ( .A(DP_OP_424J2_126_3477_n454), .B(
        DP_OP_424J2_126_3477_n452), .CI(DP_OP_424J2_126_3477_n450), .CO(
        DP_OP_424J2_126_3477_n362), .S(DP_OP_424J2_126_3477_n363) );
  FADDX1_HVT DP_OP_424J2_126_3477_U337 ( .A(DP_OP_424J2_126_3477_n446), .B(
        DP_OP_424J2_126_3477_n442), .CI(DP_OP_424J2_126_3477_n440), .CO(
        DP_OP_424J2_126_3477_n360), .S(DP_OP_424J2_126_3477_n361) );
  FADDX1_HVT DP_OP_424J2_126_3477_U336 ( .A(DP_OP_424J2_126_3477_n438), .B(
        DP_OP_424J2_126_3477_n436), .CI(DP_OP_424J2_126_3477_n434), .CO(
        DP_OP_424J2_126_3477_n358), .S(DP_OP_424J2_126_3477_n359) );
  FADDX1_HVT DP_OP_424J2_126_3477_U335 ( .A(DP_OP_424J2_126_3477_n432), .B(
        DP_OP_424J2_126_3477_n367), .CI(DP_OP_424J2_126_3477_n430), .CO(
        DP_OP_424J2_126_3477_n356), .S(DP_OP_424J2_126_3477_n357) );
  FADDX1_HVT DP_OP_424J2_126_3477_U334 ( .A(DP_OP_424J2_126_3477_n428), .B(
        DP_OP_424J2_126_3477_n363), .CI(DP_OP_424J2_126_3477_n365), .CO(
        DP_OP_424J2_126_3477_n354), .S(DP_OP_424J2_126_3477_n355) );
  FADDX1_HVT DP_OP_424J2_126_3477_U333 ( .A(DP_OP_424J2_126_3477_n426), .B(
        DP_OP_424J2_126_3477_n424), .CI(DP_OP_424J2_126_3477_n422), .CO(
        DP_OP_424J2_126_3477_n352), .S(DP_OP_424J2_126_3477_n353) );
  FADDX1_HVT DP_OP_424J2_126_3477_U332 ( .A(DP_OP_424J2_126_3477_n420), .B(
        DP_OP_424J2_126_3477_n361), .CI(DP_OP_424J2_126_3477_n418), .CO(
        DP_OP_424J2_126_3477_n350), .S(DP_OP_424J2_126_3477_n351) );
  FADDX1_HVT DP_OP_424J2_126_3477_U331 ( .A(DP_OP_424J2_126_3477_n416), .B(
        DP_OP_424J2_126_3477_n359), .CI(DP_OP_424J2_126_3477_n414), .CO(
        DP_OP_424J2_126_3477_n348), .S(DP_OP_424J2_126_3477_n349) );
  FADDX1_HVT DP_OP_424J2_126_3477_U330 ( .A(DP_OP_424J2_126_3477_n412), .B(
        DP_OP_424J2_126_3477_n357), .CI(DP_OP_424J2_126_3477_n410), .CO(
        DP_OP_424J2_126_3477_n346), .S(DP_OP_424J2_126_3477_n347) );
  FADDX1_HVT DP_OP_424J2_126_3477_U329 ( .A(DP_OP_424J2_126_3477_n355), .B(
        DP_OP_424J2_126_3477_n408), .CI(DP_OP_424J2_126_3477_n406), .CO(
        DP_OP_424J2_126_3477_n344), .S(DP_OP_424J2_126_3477_n345) );
  FADDX1_HVT DP_OP_424J2_126_3477_U328 ( .A(DP_OP_424J2_126_3477_n353), .B(
        DP_OP_424J2_126_3477_n404), .CI(DP_OP_424J2_126_3477_n402), .CO(
        DP_OP_424J2_126_3477_n342), .S(DP_OP_424J2_126_3477_n343) );
  FADDX1_HVT DP_OP_424J2_126_3477_U327 ( .A(DP_OP_424J2_126_3477_n351), .B(
        DP_OP_424J2_126_3477_n400), .CI(DP_OP_424J2_126_3477_n349), .CO(
        DP_OP_424J2_126_3477_n340), .S(DP_OP_424J2_126_3477_n341) );
  FADDX1_HVT DP_OP_424J2_126_3477_U326 ( .A(DP_OP_424J2_126_3477_n398), .B(
        DP_OP_424J2_126_3477_n347), .CI(DP_OP_424J2_126_3477_n396), .CO(
        DP_OP_424J2_126_3477_n338), .S(DP_OP_424J2_126_3477_n339) );
  FADDX1_HVT DP_OP_424J2_126_3477_U325 ( .A(DP_OP_424J2_126_3477_n394), .B(
        DP_OP_424J2_126_3477_n345), .CI(DP_OP_424J2_126_3477_n392), .CO(
        DP_OP_424J2_126_3477_n336), .S(DP_OP_424J2_126_3477_n337) );
  FADDX1_HVT DP_OP_424J2_126_3477_U324 ( .A(DP_OP_424J2_126_3477_n343), .B(
        DP_OP_424J2_126_3477_n390), .CI(DP_OP_424J2_126_3477_n388), .CO(
        DP_OP_424J2_126_3477_n334), .S(DP_OP_424J2_126_3477_n335) );
  FADDX1_HVT DP_OP_424J2_126_3477_U323 ( .A(DP_OP_424J2_126_3477_n341), .B(
        DP_OP_424J2_126_3477_n386), .CI(DP_OP_424J2_126_3477_n339), .CO(
        DP_OP_424J2_126_3477_n332), .S(DP_OP_424J2_126_3477_n333) );
  FADDX1_HVT DP_OP_424J2_126_3477_U322 ( .A(DP_OP_424J2_126_3477_n384), .B(
        DP_OP_424J2_126_3477_n337), .CI(DP_OP_424J2_126_3477_n382), .CO(
        DP_OP_424J2_126_3477_n330), .S(DP_OP_424J2_126_3477_n331) );
  FADDX1_HVT DP_OP_424J2_126_3477_U321 ( .A(DP_OP_424J2_126_3477_n380), .B(
        DP_OP_424J2_126_3477_n335), .CI(DP_OP_424J2_126_3477_n333), .CO(
        DP_OP_424J2_126_3477_n328), .S(DP_OP_424J2_126_3477_n329) );
  FADDX1_HVT DP_OP_424J2_126_3477_U320 ( .A(DP_OP_424J2_126_3477_n378), .B(
        DP_OP_424J2_126_3477_n331), .CI(DP_OP_424J2_126_3477_n376), .CO(
        DP_OP_424J2_126_3477_n326), .S(DP_OP_424J2_126_3477_n327) );
  FADDX1_HVT DP_OP_424J2_126_3477_U319 ( .A(DP_OP_424J2_126_3477_n374), .B(
        DP_OP_424J2_126_3477_n329), .CI(DP_OP_424J2_126_3477_n372), .CO(
        DP_OP_424J2_126_3477_n324), .S(DP_OP_424J2_126_3477_n325) );
  FADDX1_HVT DP_OP_424J2_126_3477_U318 ( .A(DP_OP_424J2_126_3477_n327), .B(
        DP_OP_424J2_126_3477_n370), .CI(DP_OP_424J2_126_3477_n325), .CO(
        DP_OP_424J2_126_3477_n322), .S(DP_OP_424J2_126_3477_n323) );
  FADDX1_HVT DP_OP_424J2_126_3477_U317 ( .A(DP_OP_424J2_126_3477_n1875), .B(
        DP_OP_424J2_126_3477_n366), .CI(DP_OP_424J2_126_3477_n364), .CO(
        DP_OP_424J2_126_3477_n320), .S(DP_OP_424J2_126_3477_n321) );
  FADDX1_HVT DP_OP_424J2_126_3477_U316 ( .A(DP_OP_424J2_126_3477_n362), .B(
        DP_OP_424J2_126_3477_n360), .CI(DP_OP_424J2_126_3477_n358), .CO(
        DP_OP_424J2_126_3477_n318), .S(DP_OP_424J2_126_3477_n319) );
  FADDX1_HVT DP_OP_424J2_126_3477_U315 ( .A(DP_OP_424J2_126_3477_n356), .B(
        DP_OP_424J2_126_3477_n321), .CI(DP_OP_424J2_126_3477_n354), .CO(
        DP_OP_424J2_126_3477_n316), .S(DP_OP_424J2_126_3477_n317) );
  FADDX1_HVT DP_OP_424J2_126_3477_U314 ( .A(DP_OP_424J2_126_3477_n352), .B(
        DP_OP_424J2_126_3477_n350), .CI(DP_OP_424J2_126_3477_n319), .CO(
        DP_OP_424J2_126_3477_n314), .S(DP_OP_424J2_126_3477_n315) );
  FADDX1_HVT DP_OP_424J2_126_3477_U313 ( .A(DP_OP_424J2_126_3477_n348), .B(
        DP_OP_424J2_126_3477_n346), .CI(DP_OP_424J2_126_3477_n317), .CO(
        DP_OP_424J2_126_3477_n312), .S(DP_OP_424J2_126_3477_n313) );
  FADDX1_HVT DP_OP_424J2_126_3477_U312 ( .A(DP_OP_424J2_126_3477_n344), .B(
        DP_OP_424J2_126_3477_n342), .CI(DP_OP_424J2_126_3477_n315), .CO(
        DP_OP_424J2_126_3477_n310), .S(DP_OP_424J2_126_3477_n311) );
  FADDX1_HVT DP_OP_424J2_126_3477_U311 ( .A(DP_OP_424J2_126_3477_n340), .B(
        DP_OP_424J2_126_3477_n313), .CI(DP_OP_424J2_126_3477_n338), .CO(
        DP_OP_424J2_126_3477_n308), .S(DP_OP_424J2_126_3477_n309) );
  FADDX1_HVT DP_OP_424J2_126_3477_U310 ( .A(DP_OP_424J2_126_3477_n336), .B(
        DP_OP_424J2_126_3477_n311), .CI(DP_OP_424J2_126_3477_n334), .CO(
        DP_OP_424J2_126_3477_n306), .S(DP_OP_424J2_126_3477_n307) );
  FADDX1_HVT DP_OP_424J2_126_3477_U309 ( .A(DP_OP_424J2_126_3477_n332), .B(
        DP_OP_424J2_126_3477_n309), .CI(DP_OP_424J2_126_3477_n330), .CO(
        DP_OP_424J2_126_3477_n304), .S(DP_OP_424J2_126_3477_n305) );
  FADDX1_HVT DP_OP_424J2_126_3477_U308 ( .A(DP_OP_424J2_126_3477_n307), .B(
        DP_OP_424J2_126_3477_n328), .CI(DP_OP_424J2_126_3477_n305), .CO(
        DP_OP_424J2_126_3477_n302), .S(DP_OP_424J2_126_3477_n303) );
  FADDX1_HVT DP_OP_424J2_126_3477_U307 ( .A(DP_OP_424J2_126_3477_n326), .B(
        DP_OP_424J2_126_3477_n324), .CI(DP_OP_424J2_126_3477_n303), .CO(
        DP_OP_424J2_126_3477_n300), .S(DP_OP_424J2_126_3477_n301) );
  FADDX1_HVT DP_OP_424J2_126_3477_U306 ( .A(DP_OP_424J2_126_3477_n1874), .B(
        DP_OP_424J2_126_3477_n320), .CI(DP_OP_424J2_126_3477_n318), .CO(
        DP_OP_424J2_126_3477_n298), .S(DP_OP_424J2_126_3477_n299) );
  FADDX1_HVT DP_OP_424J2_126_3477_U305 ( .A(DP_OP_424J2_126_3477_n316), .B(
        DP_OP_424J2_126_3477_n299), .CI(DP_OP_424J2_126_3477_n314), .CO(
        DP_OP_424J2_126_3477_n296), .S(DP_OP_424J2_126_3477_n297) );
  FADDX1_HVT DP_OP_424J2_126_3477_U304 ( .A(DP_OP_424J2_126_3477_n312), .B(
        DP_OP_424J2_126_3477_n310), .CI(DP_OP_424J2_126_3477_n297), .CO(
        DP_OP_424J2_126_3477_n294), .S(DP_OP_424J2_126_3477_n295) );
  FADDX1_HVT DP_OP_424J2_126_3477_U303 ( .A(DP_OP_424J2_126_3477_n308), .B(
        DP_OP_424J2_126_3477_n295), .CI(DP_OP_424J2_126_3477_n306), .CO(
        DP_OP_424J2_126_3477_n292), .S(DP_OP_424J2_126_3477_n293) );
  FADDX1_HVT DP_OP_424J2_126_3477_U302 ( .A(DP_OP_424J2_126_3477_n304), .B(
        DP_OP_424J2_126_3477_n293), .CI(DP_OP_424J2_126_3477_n302), .CO(
        DP_OP_424J2_126_3477_n290), .S(DP_OP_424J2_126_3477_n291) );
  FADDX1_HVT DP_OP_424J2_126_3477_U300 ( .A(DP_OP_424J2_126_3477_n289), .B(
        DP_OP_424J2_126_3477_n298), .CI(DP_OP_424J2_126_3477_n296), .CO(
        DP_OP_424J2_126_3477_n286), .S(DP_OP_424J2_126_3477_n287) );
  FADDX1_HVT DP_OP_424J2_126_3477_U299 ( .A(DP_OP_424J2_126_3477_n287), .B(
        DP_OP_424J2_126_3477_n294), .CI(DP_OP_424J2_126_3477_n292), .CO(
        DP_OP_424J2_126_3477_n284), .S(DP_OP_424J2_126_3477_n285) );
  FADDX1_HVT DP_OP_424J2_126_3477_U298 ( .A(DP_OP_424J2_126_3477_n1873), .B(
        DP_OP_424J2_126_3477_n288), .CI(DP_OP_424J2_126_3477_n286), .CO(
        DP_OP_424J2_126_3477_n282), .S(DP_OP_424J2_126_3477_n283) );
  FADDX1_HVT DP_OP_424J2_126_3477_U281 ( .A(DP_OP_424J2_126_3477_n1853), .B(
        DP_OP_424J2_126_3477_n1851), .CI(DP_OP_424J2_126_3477_n1849), .CO(
        DP_OP_424J2_126_3477_n219), .S(n_conv2_sum_c[0]) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U280 ( .A1(DP_OP_424J2_126_3477_n1787), 
        .A2(DP_OP_424J2_126_3477_n1789), .Y(DP_OP_424J2_126_3477_n218) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U279 ( .A1(DP_OP_424J2_126_3477_n1789), .A2(
        DP_OP_424J2_126_3477_n1787), .Y(DP_OP_424J2_126_3477_n217) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U273 ( .A1(DP_OP_424J2_126_3477_n1681), 
        .A2(DP_OP_424J2_126_3477_n1683), .Y(DP_OP_424J2_126_3477_n215) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U265 ( .A1(DP_OP_424J2_126_3477_n1527), 
        .A2(DP_OP_424J2_126_3477_n1529), .Y(DP_OP_424J2_126_3477_n210) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U264 ( .A1(DP_OP_424J2_126_3477_n1529), .A2(
        DP_OP_424J2_126_3477_n1527), .Y(DP_OP_424J2_126_3477_n209) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U259 ( .A1(DP_OP_424J2_126_3477_n1351), 
        .A2(DP_OP_424J2_126_3477_n1353), .Y(DP_OP_424J2_126_3477_n207) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U251 ( .A1(DP_OP_424J2_126_3477_n1163), 
        .A2(DP_OP_424J2_126_3477_n1165), .Y(DP_OP_424J2_126_3477_n202) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U250 ( .A1(DP_OP_424J2_126_3477_n1165), .A2(
        DP_OP_424J2_126_3477_n1163), .Y(DP_OP_424J2_126_3477_n201) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U245 ( .A1(DP_OP_424J2_126_3477_n969), .A2(
        DP_OP_424J2_126_3477_n971), .Y(DP_OP_424J2_126_3477_n199) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U237 ( .A1(DP_OP_424J2_126_3477_n773), .A2(
        DP_OP_424J2_126_3477_n968), .Y(DP_OP_424J2_126_3477_n194) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U236 ( .A1(DP_OP_424J2_126_3477_n968), .A2(
        DP_OP_424J2_126_3477_n773), .Y(DP_OP_424J2_126_3477_n193) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U230 ( .A1(DP_OP_424J2_126_3477_n599), .A2(
        DP_OP_424J2_126_3477_n772), .Y(DP_OP_424J2_126_3477_n190) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U229 ( .A1(DP_OP_424J2_126_3477_n772), .A2(
        DP_OP_424J2_126_3477_n599), .Y(DP_OP_424J2_126_3477_n189) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U224 ( .A1(DP_OP_424J2_126_3477_n463), .A2(
        DP_OP_424J2_126_3477_n598), .Y(DP_OP_424J2_126_3477_n187) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U223 ( .A1(DP_OP_424J2_126_3477_n598), .A2(
        DP_OP_424J2_126_3477_n463), .Y(DP_OP_424J2_126_3477_n186) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U219 ( .A1(DP_OP_424J2_126_3477_n189), .A2(
        DP_OP_424J2_126_3477_n186), .Y(DP_OP_424J2_126_3477_n184) );
  AOI21X1_HVT DP_OP_424J2_126_3477_U218 ( .A1(DP_OP_424J2_126_3477_n184), .A2(
        DP_OP_424J2_126_3477_n192), .A3(DP_OP_424J2_126_3477_n185), .Y(
        DP_OP_424J2_126_3477_n183) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U215 ( .A1(DP_OP_424J2_126_3477_n369), .A2(
        DP_OP_424J2_126_3477_n462), .Y(DP_OP_424J2_126_3477_n181) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U214 ( .A1(DP_OP_424J2_126_3477_n462), .A2(
        DP_OP_424J2_126_3477_n369), .Y(DP_OP_424J2_126_3477_n180) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U212 ( .A1(DP_OP_424J2_126_3477_n241), .A2(
        DP_OP_424J2_126_3477_n181), .Y(DP_OP_424J2_126_3477_n26) );
  AOI21X1_HVT DP_OP_424J2_126_3477_U209 ( .A1(DP_OP_424J2_126_3477_n182), .A2(
        DP_OP_424J2_126_3477_n241), .A3(DP_OP_424J2_126_3477_n179), .Y(
        DP_OP_424J2_126_3477_n177) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U207 ( .A1(DP_OP_424J2_126_3477_n323), .A2(
        DP_OP_424J2_126_3477_n368), .Y(DP_OP_424J2_126_3477_n176) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U206 ( .A1(DP_OP_424J2_126_3477_n368), .A2(
        DP_OP_424J2_126_3477_n323), .Y(DP_OP_424J2_126_3477_n175) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U204 ( .A1(DP_OP_424J2_126_3477_n240), .A2(
        DP_OP_424J2_126_3477_n176), .Y(DP_OP_424J2_126_3477_n25) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U202 ( .A1(DP_OP_424J2_126_3477_n175), .A2(
        DP_OP_424J2_126_3477_n180), .Y(DP_OP_424J2_126_3477_n173) );
  AOI21X1_HVT DP_OP_424J2_126_3477_U201 ( .A1(DP_OP_424J2_126_3477_n182), .A2(
        DP_OP_424J2_126_3477_n173), .A3(DP_OP_424J2_126_3477_n174), .Y(
        DP_OP_424J2_126_3477_n172) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U199 ( .A1(DP_OP_424J2_126_3477_n301), .A2(
        DP_OP_424J2_126_3477_n322), .Y(DP_OP_424J2_126_3477_n171) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U198 ( .A1(DP_OP_424J2_126_3477_n322), .A2(
        DP_OP_424J2_126_3477_n301), .Y(DP_OP_424J2_126_3477_n170) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U193 ( .A1(DP_OP_424J2_126_3477_n300), .A2(
        DP_OP_424J2_126_3477_n291), .Y(DP_OP_424J2_126_3477_n168) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U192 ( .A1(DP_OP_424J2_126_3477_n291), .A2(
        DP_OP_424J2_126_3477_n300), .Y(DP_OP_424J2_126_3477_n167) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U188 ( .A1(DP_OP_424J2_126_3477_n167), .A2(
        DP_OP_424J2_126_3477_n170), .Y(DP_OP_424J2_126_3477_n165) );
  AOI21X1_HVT DP_OP_424J2_126_3477_U187 ( .A1(DP_OP_424J2_126_3477_n174), .A2(
        DP_OP_424J2_126_3477_n165), .A3(DP_OP_424J2_126_3477_n166), .Y(
        DP_OP_424J2_126_3477_n164) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U186 ( .A1(DP_OP_424J2_126_3477_n173), .A2(
        DP_OP_424J2_126_3477_n165), .Y(DP_OP_424J2_126_3477_n163) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U182 ( .A1(DP_OP_424J2_126_3477_n290), .A2(
        DP_OP_424J2_126_3477_n285), .Y(DP_OP_424J2_126_3477_n152) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U181 ( .A1(DP_OP_424J2_126_3477_n285), .A2(
        DP_OP_424J2_126_3477_n290), .Y(DP_OP_424J2_126_3477_n151) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U179 ( .A1(DP_OP_424J2_126_3477_n237), .A2(
        DP_OP_424J2_126_3477_n152), .Y(DP_OP_424J2_126_3477_n22) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U168 ( .A1(DP_OP_424J2_126_3477_n284), .A2(
        DP_OP_424J2_126_3477_n283), .Y(DP_OP_424J2_126_3477_n149) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U167 ( .A1(DP_OP_424J2_126_3477_n283), .A2(
        DP_OP_424J2_126_3477_n284), .Y(DP_OP_424J2_126_3477_n148) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U165 ( .A1(DP_OP_424J2_126_3477_n236), .A2(
        DP_OP_424J2_126_3477_n149), .Y(DP_OP_424J2_126_3477_n21) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U161 ( .A1(DP_OP_424J2_126_3477_n237), .A2(
        DP_OP_424J2_126_3477_n236), .Y(DP_OP_424J2_126_3477_n144) );
  AOI21X1_HVT DP_OP_424J2_126_3477_U158 ( .A1(DP_OP_424J2_126_3477_n162), .A2(
        DP_OP_424J2_126_3477_n142), .A3(DP_OP_424J2_126_3477_n143), .Y(
        DP_OP_424J2_126_3477_n141) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U156 ( .A1(DP_OP_424J2_126_3477_n282), .A2(
        DP_OP_424J2_126_3477_n281), .Y(DP_OP_424J2_126_3477_n140) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U155 ( .A1(DP_OP_424J2_126_3477_n281), .A2(
        DP_OP_424J2_126_3477_n282), .Y(DP_OP_424J2_126_3477_n137) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U146 ( .A1(DP_OP_424J2_126_3477_n279), .A2(
        DP_OP_424J2_126_3477_n280), .Y(DP_OP_424J2_126_3477_n133) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U145 ( .A1(DP_OP_424J2_126_3477_n280), .A2(
        DP_OP_424J2_126_3477_n279), .Y(DP_OP_424J2_126_3477_n132) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U140 ( .A1(DP_OP_424J2_126_3477_n277), .A2(
        DP_OP_424J2_126_3477_n278), .Y(DP_OP_424J2_126_3477_n130) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U139 ( .A1(DP_OP_424J2_126_3477_n278), .A2(
        DP_OP_424J2_126_3477_n277), .Y(DP_OP_424J2_126_3477_n129) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U135 ( .A1(DP_OP_424J2_126_3477_n129), .A2(
        DP_OP_424J2_126_3477_n132), .Y(DP_OP_424J2_126_3477_n127) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U130 ( .A1(DP_OP_424J2_126_3477_n275), .A2(
        DP_OP_424J2_126_3477_n276), .Y(DP_OP_424J2_126_3477_n123) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U123 ( .A1(DP_OP_424J2_126_3477_n127), .A2(
        n452), .Y(DP_OP_424J2_126_3477_n118) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U120 ( .A1(DP_OP_424J2_126_3477_n273), .A2(
        DP_OP_424J2_126_3477_n274), .Y(DP_OP_424J2_126_3477_n116) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U119 ( .A1(DP_OP_424J2_126_3477_n274), .A2(
        DP_OP_424J2_126_3477_n273), .Y(DP_OP_424J2_126_3477_n115) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U110 ( .A1(DP_OP_424J2_126_3477_n271), .A2(
        DP_OP_424J2_126_3477_n272), .Y(DP_OP_424J2_126_3477_n109) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U103 ( .A1(DP_OP_424J2_126_3477_n113), .A2(
        n451), .Y(DP_OP_424J2_126_3477_n104) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U100 ( .A1(DP_OP_424J2_126_3477_n269), .A2(
        DP_OP_424J2_126_3477_n270), .Y(DP_OP_424J2_126_3477_n102) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U99 ( .A1(DP_OP_424J2_126_3477_n270), .A2(
        DP_OP_424J2_126_3477_n269), .Y(DP_OP_424J2_126_3477_n101) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U90 ( .A1(DP_OP_424J2_126_3477_n267), .A2(
        DP_OP_424J2_126_3477_n268), .Y(DP_OP_424J2_126_3477_n95) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U83 ( .A1(DP_OP_424J2_126_3477_n99), .A2(
        n447), .Y(DP_OP_424J2_126_3477_n90) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U80 ( .A1(DP_OP_424J2_126_3477_n265), .A2(
        DP_OP_424J2_126_3477_n266), .Y(DP_OP_424J2_126_3477_n88) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U79 ( .A1(DP_OP_424J2_126_3477_n266), .A2(
        DP_OP_424J2_126_3477_n265), .Y(DP_OP_424J2_126_3477_n87) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U70 ( .A1(DP_OP_424J2_126_3477_n263), .A2(
        DP_OP_424J2_126_3477_n264), .Y(DP_OP_424J2_126_3477_n81) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U63 ( .A1(DP_OP_424J2_126_3477_n85), .A2(
        n446), .Y(DP_OP_424J2_126_3477_n76) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U61 ( .A1(DP_OP_424J2_126_3477_n76), .A2(
        DP_OP_424J2_126_3477_n137), .Y(DP_OP_424J2_126_3477_n74) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U56 ( .A1(DP_OP_424J2_126_3477_n261), .A2(
        DP_OP_424J2_126_3477_n262), .Y(DP_OP_424J2_126_3477_n70) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U49 ( .A1(DP_OP_424J2_126_3477_n74), .A2(
        n445), .Y(DP_OP_424J2_126_3477_n65) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U45 ( .A1(DP_OP_424J2_126_3477_n237), .A2(
        DP_OP_424J2_126_3477_n63), .Y(DP_OP_424J2_126_3477_n61) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U42 ( .A1(DP_OP_424J2_126_3477_n259), .A2(
        DP_OP_424J2_126_3477_n260), .Y(DP_OP_424J2_126_3477_n59) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U41 ( .A1(DP_OP_424J2_126_3477_n260), .A2(
        DP_OP_424J2_126_3477_n259), .Y(DP_OP_424J2_126_3477_n58) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U32 ( .A1(DP_OP_424J2_126_3477_n257), .A2(
        DP_OP_424J2_126_3477_n258), .Y(DP_OP_424J2_126_3477_n52) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U25 ( .A1(DP_OP_424J2_126_3477_n56), .A2(
        n444), .Y(DP_OP_424J2_126_3477_n47) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U22 ( .A1(DP_OP_424J2_126_3477_n255), .A2(
        DP_OP_424J2_126_3477_n256), .Y(DP_OP_424J2_126_3477_n45) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U21 ( .A1(DP_OP_424J2_126_3477_n256), .A2(
        DP_OP_424J2_126_3477_n255), .Y(DP_OP_424J2_126_3477_n44) );
  AOI21X1_HVT DP_OP_424J2_126_3477_U16 ( .A1(DP_OP_424J2_126_3477_n162), .A2(
        DP_OP_424J2_126_3477_n42), .A3(DP_OP_424J2_126_3477_n43), .Y(
        DP_OP_424J2_126_3477_n41) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U14 ( .A1(DP_OP_424J2_126_3477_n253), .A2(
        DP_OP_424J2_126_3477_n254), .Y(DP_OP_424J2_126_3477_n40) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U13 ( .A1(DP_OP_424J2_126_3477_n254), .A2(
        DP_OP_424J2_126_3477_n253), .Y(DP_OP_424J2_126_3477_n39) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U8 ( .A1(n443), .A2(
        DP_OP_424J2_126_3477_n252), .Y(DP_OP_424J2_126_3477_n37) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U96 ( .A1(DP_OP_423J2_125_3477_n101), .A2(
        DP_OP_423J2_125_3477_n105), .A3(DP_OP_423J2_125_3477_n102), .Y(
        DP_OP_423J2_125_3477_n100) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U261 ( .A1(DP_OP_423J2_125_3477_n211), .A2(
        DP_OP_423J2_125_3477_n209), .A3(DP_OP_423J2_125_3477_n210), .Y(
        DP_OP_423J2_125_3477_n208) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U76 ( .A1(DP_OP_423J2_125_3477_n87), .A2(
        DP_OP_423J2_125_3477_n91), .A3(DP_OP_423J2_125_3477_n88), .Y(
        DP_OP_423J2_125_3477_n86) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U116 ( .A1(DP_OP_423J2_125_3477_n115), .A2(
        DP_OP_423J2_125_3477_n119), .A3(DP_OP_423J2_125_3477_n116), .Y(
        DP_OP_423J2_125_3477_n114) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U136 ( .A1(DP_OP_423J2_125_3477_n133), .A2(
        DP_OP_423J2_125_3477_n129), .A3(DP_OP_423J2_125_3477_n130), .Y(
        DP_OP_423J2_125_3477_n128) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U275 ( .A1(DP_OP_423J2_125_3477_n4), .A2(
        DP_OP_423J2_125_3477_n217), .A3(DP_OP_423J2_125_3477_n218), .Y(
        DP_OP_423J2_125_3477_n216) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1111 ( .A1(n363), .A2(n387), .Y(
        DP_OP_423J2_125_3477_n288) );
  XNOR2X1_HVT DP_OP_423J2_125_3477_U737 ( .A1(DP_OP_423J2_125_3477_n2452), 
        .A2(DP_OP_423J2_125_3477_n2979), .Y(DP_OP_423J2_125_3477_n1161) );
  XNOR2X2_HVT DP_OP_423J2_125_3477_U131 ( .A1(DP_OP_423J2_125_3477_n131), .A2(
        DP_OP_423J2_125_3477_n18), .Y(n_conv2_sum_b[18]) );
  OAI21X2_HVT DP_OP_423J2_125_3477_U142 ( .A1(DP_OP_423J2_125_3477_n132), .A2(
        DP_OP_423J2_125_3477_n3), .A3(DP_OP_423J2_125_3477_n133), .Y(
        DP_OP_423J2_125_3477_n131) );
  XNOR2X2_HVT DP_OP_423J2_125_3477_U121 ( .A1(DP_OP_423J2_125_3477_n124), .A2(
        DP_OP_423J2_125_3477_n17), .Y(n_conv2_sum_b[19]) );
  OAI21X2_HVT DP_OP_423J2_125_3477_U132 ( .A1(DP_OP_423J2_125_3477_n125), .A2(
        DP_OP_423J2_125_3477_n3), .A3(DP_OP_423J2_125_3477_n126), .Y(
        DP_OP_423J2_125_3477_n124) );
  OAI21X2_HVT DP_OP_423J2_125_3477_U185 ( .A1(DP_OP_423J2_125_3477_n163), .A2(
        DP_OP_423J2_125_3477_n183), .A3(DP_OP_423J2_125_3477_n164), .Y(
        DP_OP_423J2_125_3477_n162) );
  OAI21X2_HVT DP_OP_423J2_125_3477_U203 ( .A1(DP_OP_423J2_125_3477_n181), .A2(
        DP_OP_423J2_125_3477_n175), .A3(DP_OP_423J2_125_3477_n176), .Y(
        DP_OP_423J2_125_3477_n174) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2240 ( .A1(DP_OP_423J2_125_3477_n3007), 
        .A2(DP_OP_423J2_125_3477_n3017), .Y(DP_OP_423J2_125_3477_n2999) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2239 ( .A1(DP_OP_423J2_125_3477_n3006), .A2(
        DP_OP_423J2_125_3477_n3017), .Y(DP_OP_423J2_125_3477_n2998) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2232 ( .A1(DP_OP_423J2_125_3477_n3007), 
        .A2(DP_OP_423J2_125_3477_n3016), .Y(DP_OP_423J2_125_3477_n2991) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2231 ( .A1(DP_OP_423J2_125_3477_n3006), .A2(
        DP_OP_423J2_125_3477_n3016), .Y(DP_OP_423J2_125_3477_n2990) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2223 ( .A1(DP_OP_423J2_125_3477_n3006), .A2(
        DP_OP_425J2_127_3477_n3015), .Y(DP_OP_423J2_125_3477_n2982) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2222 ( .A1(DP_OP_425J2_127_3477_n2047), .A2(
        DP_OP_423J2_125_3477_n3014), .Y(DP_OP_423J2_125_3477_n1678) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2221 ( .A1(DP_OP_423J2_125_3477_n3012), .A2(
        DP_OP_423J2_125_3477_n3014), .Y(DP_OP_423J2_125_3477_n2981) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2220 ( .A1(DP_OP_423J2_125_3477_n3011), .A2(
        DP_OP_423J2_125_3477_n3014), .Y(DP_OP_423J2_125_3477_n2980) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2219 ( .A1(DP_OP_423J2_125_3477_n3010), .A2(
        DP_OP_423J2_125_3477_n3014), .Y(DP_OP_423J2_125_3477_n2979) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2218 ( .A1(DP_OP_423J2_125_3477_n3009), .A2(
        DP_OP_423J2_125_3477_n3014), .Y(DP_OP_423J2_125_3477_n2978) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2217 ( .A1(DP_OP_423J2_125_3477_n3008), .A2(
        DP_OP_423J2_125_3477_n3014), .Y(DP_OP_423J2_125_3477_n770) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2216 ( .A1(DP_OP_423J2_125_3477_n3007), .A2(
        DP_OP_423J2_125_3477_n3014), .Y(DP_OP_423J2_125_3477_n2977) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2215 ( .A1(DP_OP_423J2_125_3477_n3006), 
        .A2(DP_OP_423J2_125_3477_n3014), .Y(DP_OP_423J2_125_3477_n2976) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2195 ( .A1(DP_OP_423J2_125_3477_n2964), .A2(
        DP_OP_425J2_127_3477_n2975), .Y(DP_OP_423J2_125_3477_n2956) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2187 ( .A1(DP_OP_423J2_125_3477_n2964), .A2(
        DP_OP_423J2_125_3477_n2974), .Y(DP_OP_423J2_125_3477_n2948) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2179 ( .A1(DP_OP_423J2_125_3477_n2964), .A2(
        DP_OP_423J2_125_3477_n2973), .Y(DP_OP_423J2_125_3477_n2940) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2178 ( .A1(DP_OP_423J2_125_3477_n2971), .A2(
        DP_OP_423J2_125_3477_n2972), .Y(DP_OP_423J2_125_3477_n2939) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2177 ( .A1(DP_OP_423J2_125_3477_n2970), .A2(
        DP_OP_423J2_125_3477_n2972), .Y(DP_OP_423J2_125_3477_n2938) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2176 ( .A1(DP_OP_423J2_125_3477_n2969), .A2(
        DP_OP_423J2_125_3477_n2972), .Y(DP_OP_423J2_125_3477_n2937) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2175 ( .A1(DP_OP_424J2_126_3477_n2880), .A2(
        DP_OP_423J2_125_3477_n2972), .Y(DP_OP_423J2_125_3477_n2936) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2174 ( .A1(DP_OP_423J2_125_3477_n2967), .A2(
        DP_OP_423J2_125_3477_n2972), .Y(DP_OP_423J2_125_3477_n2935) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2173 ( .A1(DP_OP_424J2_126_3477_n2878), .A2(
        DP_OP_423J2_125_3477_n2972), .Y(DP_OP_423J2_125_3477_n2934) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2172 ( .A1(DP_OP_425J2_127_3477_n2085), .A2(
        DP_OP_423J2_125_3477_n2972), .Y(DP_OP_423J2_125_3477_n2933) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2171 ( .A1(DP_OP_423J2_125_3477_n2964), 
        .A2(DP_OP_423J2_125_3477_n2972), .Y(DP_OP_423J2_125_3477_n2932) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2151 ( .A1(DP_OP_423J2_125_3477_n2920), .A2(
        DP_OP_423J2_125_3477_n2931), .Y(DP_OP_423J2_125_3477_n2912) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2143 ( .A1(DP_OP_423J2_125_3477_n2920), .A2(
        DP_OP_423J2_125_3477_n2930), .Y(DP_OP_423J2_125_3477_n2904) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2135 ( .A1(DP_OP_423J2_125_3477_n2920), .A2(
        DP_OP_423J2_125_3477_n2929), .Y(DP_OP_423J2_125_3477_n2896) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2134 ( .A1(DP_OP_423J2_125_3477_n2927), .A2(
        DP_OP_423J2_125_3477_n2928), .Y(DP_OP_423J2_125_3477_n2895) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2133 ( .A1(DP_OP_423J2_125_3477_n2926), .A2(
        DP_OP_423J2_125_3477_n2928), .Y(DP_OP_423J2_125_3477_n2894) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2132 ( .A1(DP_OP_425J2_127_3477_n2133), .A2(
        DP_OP_423J2_125_3477_n2928), .Y(DP_OP_423J2_125_3477_n2893) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2131 ( .A1(DP_OP_423J2_125_3477_n2924), .A2(
        DP_OP_423J2_125_3477_n2928), .Y(DP_OP_423J2_125_3477_n2892) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2130 ( .A1(DP_OP_423J2_125_3477_n2923), .A2(
        DP_OP_423J2_125_3477_n2928), .Y(DP_OP_423J2_125_3477_n2891) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2129 ( .A1(DP_OP_423J2_125_3477_n2922), .A2(
        DP_OP_423J2_125_3477_n2928), .Y(DP_OP_423J2_125_3477_n2890) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2128 ( .A1(DP_OP_423J2_125_3477_n2921), .A2(
        DP_OP_423J2_125_3477_n2928), .Y(DP_OP_423J2_125_3477_n2889) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2127 ( .A1(DP_OP_423J2_125_3477_n2920), 
        .A2(DP_OP_423J2_125_3477_n2928), .Y(DP_OP_423J2_125_3477_n2888) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2107 ( .A1(DP_OP_422J2_124_3477_n2040), .A2(
        DP_OP_424J2_126_3477_n2887), .Y(DP_OP_423J2_125_3477_n2868) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2099 ( .A1(DP_OP_422J2_124_3477_n2040), .A2(
        DP_OP_423J2_125_3477_n2886), .Y(DP_OP_423J2_125_3477_n2860) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2092 ( .A1(DP_OP_423J2_125_3477_n2877), 
        .A2(DP_OP_423J2_125_3477_n2885), .Y(DP_OP_423J2_125_3477_n2853) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2091 ( .A1(DP_OP_425J2_127_3477_n2172), .A2(
        DP_OP_423J2_125_3477_n2885), .Y(DP_OP_423J2_125_3477_n2852) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2090 ( .A1(DP_OP_424J2_126_3477_n2795), .A2(
        DP_OP_423J2_125_3477_n2884), .Y(DP_OP_423J2_125_3477_n2851) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2089 ( .A1(DP_OP_425J2_127_3477_n2178), .A2(
        DP_OP_423J2_125_3477_n2884), .Y(DP_OP_423J2_125_3477_n2850) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2088 ( .A1(DP_OP_422J2_124_3477_n2045), .A2(
        DP_OP_423J2_125_3477_n2884), .Y(DP_OP_423J2_125_3477_n2849) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2087 ( .A1(DP_OP_423J2_125_3477_n2880), .A2(
        DP_OP_423J2_125_3477_n2884), .Y(DP_OP_423J2_125_3477_n2848) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2086 ( .A1(DP_OP_424J2_126_3477_n2791), .A2(
        DP_OP_423J2_125_3477_n2884), .Y(DP_OP_423J2_125_3477_n2847) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2085 ( .A1(DP_OP_423J2_125_3477_n2878), .A2(
        DP_OP_423J2_125_3477_n2884), .Y(DP_OP_423J2_125_3477_n2846) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2084 ( .A1(DP_OP_423J2_125_3477_n2877), .A2(
        DP_OP_423J2_125_3477_n2884), .Y(DP_OP_423J2_125_3477_n2845) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2083 ( .A1(DP_OP_422J2_124_3477_n2040), 
        .A2(DP_OP_423J2_125_3477_n2884), .Y(DP_OP_423J2_125_3477_n2844) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2063 ( .A1(DP_OP_425J2_127_3477_n2216), .A2(
        DP_OP_423J2_125_3477_n2843), .Y(DP_OP_423J2_125_3477_n2824) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2055 ( .A1(DP_OP_425J2_127_3477_n2216), .A2(
        DP_OP_423J2_125_3477_n2842), .Y(DP_OP_423J2_125_3477_n2816) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2048 ( .A1(DP_OP_424J2_126_3477_n2745), 
        .A2(DP_OP_425J2_127_3477_n2841), .Y(DP_OP_423J2_125_3477_n2809) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2047 ( .A1(DP_OP_422J2_124_3477_n2084), .A2(
        DP_OP_422J2_124_3477_n2841), .Y(DP_OP_423J2_125_3477_n2808) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2046 ( .A1(DP_OP_422J2_124_3477_n2091), .A2(
        DP_OP_423J2_125_3477_n2840), .Y(DP_OP_423J2_125_3477_n2807) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2045 ( .A1(DP_OP_422J2_124_3477_n2090), .A2(
        DP_OP_423J2_125_3477_n2840), .Y(DP_OP_423J2_125_3477_n2806) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2044 ( .A1(DP_OP_423J2_125_3477_n2837), .A2(
        DP_OP_423J2_125_3477_n2840), .Y(DP_OP_423J2_125_3477_n2805) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2043 ( .A1(DP_OP_425J2_127_3477_n2220), .A2(
        DP_OP_423J2_125_3477_n2840), .Y(DP_OP_423J2_125_3477_n2804) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2042 ( .A1(DP_OP_425J2_127_3477_n2219), .A2(
        DP_OP_423J2_125_3477_n2840), .Y(DP_OP_423J2_125_3477_n2803) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2041 ( .A1(DP_OP_423J2_125_3477_n2834), .A2(
        DP_OP_423J2_125_3477_n2840), .Y(DP_OP_423J2_125_3477_n2802) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2040 ( .A1(DP_OP_425J2_127_3477_n2217), .A2(
        DP_OP_423J2_125_3477_n2840), .Y(DP_OP_423J2_125_3477_n2801) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2039 ( .A1(DP_OP_422J2_124_3477_n2084), 
        .A2(DP_OP_423J2_125_3477_n2840), .Y(DP_OP_423J2_125_3477_n2800) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2020 ( .A1(DP_OP_425J2_127_3477_n2261), 
        .A2(DP_OP_422J2_124_3477_n2799), .Y(DP_OP_423J2_125_3477_n2781) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2019 ( .A1(DP_OP_425J2_127_3477_n2260), .A2(
        DP_OP_425J2_127_3477_n2799), .Y(DP_OP_423J2_125_3477_n2780) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2011 ( .A1(DP_OP_425J2_127_3477_n2260), .A2(
        DP_OP_423J2_125_3477_n2798), .Y(DP_OP_423J2_125_3477_n2772) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2004 ( .A1(DP_OP_425J2_127_3477_n2261), 
        .A2(DP_OP_424J2_126_3477_n2797), .Y(DP_OP_423J2_125_3477_n2765) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2003 ( .A1(DP_OP_425J2_127_3477_n2260), .A2(
        DP_OP_425J2_127_3477_n2797), .Y(DP_OP_423J2_125_3477_n2764) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2002 ( .A1(DP_OP_423J2_125_3477_n2795), .A2(
        DP_OP_423J2_125_3477_n2796), .Y(DP_OP_423J2_125_3477_n2763) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2001 ( .A1(DP_OP_423J2_125_3477_n2794), .A2(
        DP_OP_423J2_125_3477_n2796), .Y(DP_OP_423J2_125_3477_n2762) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2000 ( .A1(DP_OP_423J2_125_3477_n2793), .A2(
        DP_OP_423J2_125_3477_n2796), .Y(DP_OP_423J2_125_3477_n2761) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1999 ( .A1(DP_OP_425J2_127_3477_n2264), .A2(
        DP_OP_423J2_125_3477_n2796), .Y(DP_OP_423J2_125_3477_n2760) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1998 ( .A1(DP_OP_423J2_125_3477_n2791), .A2(
        DP_OP_423J2_125_3477_n2796), .Y(DP_OP_423J2_125_3477_n2759) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1997 ( .A1(DP_OP_423J2_125_3477_n2790), .A2(
        DP_OP_423J2_125_3477_n2796), .Y(DP_OP_423J2_125_3477_n2758) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1996 ( .A1(DP_OP_425J2_127_3477_n2261), .A2(
        DP_OP_423J2_125_3477_n2796), .Y(DP_OP_423J2_125_3477_n2757) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1995 ( .A1(DP_OP_425J2_127_3477_n2260), 
        .A2(DP_OP_423J2_125_3477_n2796), .Y(DP_OP_423J2_125_3477_n2756) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1982 ( .A1(DP_OP_424J2_126_3477_n2663), 
        .A2(DP_OP_423J2_125_3477_n2755), .Y(DP_OP_423J2_125_3477_n2743) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1981 ( .A1(DP_OP_423J2_125_3477_n2750), 
        .A2(DP_OP_423J2_125_3477_n2755), .Y(DP_OP_423J2_125_3477_n2742) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1980 ( .A1(DP_OP_423J2_125_3477_n2749), 
        .A2(DP_OP_423J2_125_3477_n2755), .Y(DP_OP_423J2_125_3477_n2741) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1979 ( .A1(DP_OP_423J2_125_3477_n2748), 
        .A2(DP_OP_423J2_125_3477_n2755), .Y(DP_OP_423J2_125_3477_n2740) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1978 ( .A1(DP_OP_423J2_125_3477_n2747), 
        .A2(DP_OP_423J2_125_3477_n2755), .Y(DP_OP_423J2_125_3477_n2739) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1977 ( .A1(DP_OP_423J2_125_3477_n2746), 
        .A2(DP_OP_423J2_125_3477_n2755), .Y(DP_OP_423J2_125_3477_n2738) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1976 ( .A1(DP_OP_423J2_125_3477_n2745), 
        .A2(DP_OP_423J2_125_3477_n2755), .Y(DP_OP_423J2_125_3477_n2737) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1975 ( .A1(DP_OP_422J2_124_3477_n2172), .A2(
        DP_OP_423J2_125_3477_n2755), .Y(DP_OP_423J2_125_3477_n2736) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1967 ( .A1(DP_OP_425J2_127_3477_n2304), .A2(
        DP_OP_423J2_125_3477_n2754), .Y(DP_OP_423J2_125_3477_n2728) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1959 ( .A1(DP_OP_422J2_124_3477_n2172), .A2(
        DP_OP_423J2_125_3477_n2753), .Y(DP_OP_423J2_125_3477_n2720) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1958 ( .A1(DP_OP_422J2_124_3477_n2179), .A2(
        DP_OP_423J2_125_3477_n2752), .Y(DP_OP_423J2_125_3477_n2719) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1957 ( .A1(DP_OP_423J2_125_3477_n2750), .A2(
        DP_OP_423J2_125_3477_n2752), .Y(DP_OP_423J2_125_3477_n2718) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1956 ( .A1(DP_OP_423J2_125_3477_n2749), .A2(
        DP_OP_423J2_125_3477_n2752), .Y(DP_OP_423J2_125_3477_n2717) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1955 ( .A1(DP_OP_423J2_125_3477_n2748), .A2(
        DP_OP_423J2_125_3477_n2752), .Y(DP_OP_423J2_125_3477_n2716) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1954 ( .A1(DP_OP_423J2_125_3477_n2747), .A2(
        DP_OP_423J2_125_3477_n2752), .Y(DP_OP_423J2_125_3477_n2715) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1953 ( .A1(DP_OP_423J2_125_3477_n2746), .A2(
        DP_OP_423J2_125_3477_n2752), .Y(DP_OP_423J2_125_3477_n2714) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1952 ( .A1(DP_OP_423J2_125_3477_n2745), .A2(
        DP_OP_423J2_125_3477_n2752), .Y(DP_OP_423J2_125_3477_n2713) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1951 ( .A1(DP_OP_425J2_127_3477_n2304), 
        .A2(DP_OP_423J2_125_3477_n2752), .Y(DP_OP_423J2_125_3477_n2712) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1932 ( .A1(DP_OP_424J2_126_3477_n2613), 
        .A2(DP_OP_424J2_126_3477_n2711), .Y(DP_OP_423J2_125_3477_n2693) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1931 ( .A1(DP_OP_423J2_125_3477_n2700), .A2(
        DP_OP_425J2_127_3477_n2711), .Y(DP_OP_423J2_125_3477_n2692) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1923 ( .A1(DP_OP_423J2_125_3477_n2700), .A2(
        DP_OP_423J2_125_3477_n2710), .Y(DP_OP_423J2_125_3477_n2684) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1916 ( .A1(DP_OP_424J2_126_3477_n2613), 
        .A2(DP_OP_423J2_125_3477_n2709), .Y(DP_OP_423J2_125_3477_n2677) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1915 ( .A1(DP_OP_423J2_125_3477_n2700), .A2(
        DP_OP_423J2_125_3477_n2709), .Y(DP_OP_423J2_125_3477_n2676) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1914 ( .A1(DP_OP_423J2_125_3477_n2707), .A2(
        DP_OP_423J2_125_3477_n2708), .Y(DP_OP_423J2_125_3477_n2675) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1913 ( .A1(DP_OP_424J2_126_3477_n2618), .A2(
        DP_OP_423J2_125_3477_n2708), .Y(DP_OP_423J2_125_3477_n2674) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1912 ( .A1(DP_OP_423J2_125_3477_n2705), .A2(
        DP_OP_423J2_125_3477_n2708), .Y(DP_OP_423J2_125_3477_n2673) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1911 ( .A1(DP_OP_422J2_124_3477_n2220), .A2(
        DP_OP_423J2_125_3477_n2708), .Y(DP_OP_423J2_125_3477_n2672) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1910 ( .A1(DP_OP_425J2_127_3477_n2351), .A2(
        DP_OP_423J2_125_3477_n2708), .Y(DP_OP_423J2_125_3477_n2671) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1909 ( .A1(DP_OP_423J2_125_3477_n2702), .A2(
        DP_OP_423J2_125_3477_n2708), .Y(DP_OP_423J2_125_3477_n2670) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1908 ( .A1(DP_OP_422J2_124_3477_n2217), .A2(
        DP_OP_423J2_125_3477_n2708), .Y(DP_OP_423J2_125_3477_n2669) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1907 ( .A1(DP_OP_423J2_125_3477_n2700), 
        .A2(DP_OP_423J2_125_3477_n2708), .Y(DP_OP_423J2_125_3477_n2668) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1888 ( .A1(DP_OP_424J2_126_3477_n2569), 
        .A2(DP_OP_423J2_125_3477_n2667), .Y(DP_OP_423J2_125_3477_n2649) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1887 ( .A1(DP_OP_423J2_125_3477_n2656), .A2(
        DP_OP_423J2_125_3477_n2667), .Y(DP_OP_423J2_125_3477_n2648) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1879 ( .A1(DP_OP_423J2_125_3477_n2656), .A2(
        DP_OP_422J2_124_3477_n2666), .Y(DP_OP_423J2_125_3477_n2640) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1871 ( .A1(DP_OP_423J2_125_3477_n2656), .A2(
        DP_OP_423J2_125_3477_n2665), .Y(DP_OP_423J2_125_3477_n2632) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1870 ( .A1(DP_OP_423J2_125_3477_n2663), .A2(
        DP_OP_423J2_125_3477_n2664), .Y(DP_OP_423J2_125_3477_n2631) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1869 ( .A1(DP_OP_423J2_125_3477_n2662), .A2(
        DP_OP_423J2_125_3477_n2664), .Y(DP_OP_423J2_125_3477_n2630) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1868 ( .A1(DP_OP_422J2_124_3477_n2265), .A2(
        DP_OP_423J2_125_3477_n2664), .Y(DP_OP_423J2_125_3477_n2629) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1867 ( .A1(DP_OP_424J2_126_3477_n2572), .A2(
        DP_OP_423J2_125_3477_n2664), .Y(DP_OP_423J2_125_3477_n2628) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1866 ( .A1(DP_OP_423J2_125_3477_n2659), .A2(
        DP_OP_423J2_125_3477_n2664), .Y(DP_OP_423J2_125_3477_n2627) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1865 ( .A1(DP_OP_423J2_125_3477_n2658), .A2(
        DP_OP_423J2_125_3477_n2664), .Y(DP_OP_423J2_125_3477_n2626) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1864 ( .A1(DP_OP_424J2_126_3477_n2569), .A2(
        DP_OP_423J2_125_3477_n2664), .Y(DP_OP_423J2_125_3477_n2625) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1863 ( .A1(DP_OP_423J2_125_3477_n2656), 
        .A2(DP_OP_423J2_125_3477_n2664), .Y(DP_OP_423J2_125_3477_n2624) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1843 ( .A1(DP_OP_423J2_125_3477_n2612), .A2(
        DP_OP_423J2_125_3477_n2623), .Y(DP_OP_423J2_125_3477_n2604) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1842 ( .A1(DP_OP_423J2_125_3477_n2619), 
        .A2(DP_OP_424J2_126_3477_n2622), .Y(DP_OP_423J2_125_3477_n2603) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1841 ( .A1(DP_OP_425J2_127_3477_n2442), 
        .A2(DP_OP_425J2_127_3477_n2622), .Y(DP_OP_423J2_125_3477_n2602) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1840 ( .A1(DP_OP_423J2_125_3477_n2617), 
        .A2(DP_OP_422J2_124_3477_n2622), .Y(DP_OP_423J2_125_3477_n2601) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1839 ( .A1(DP_OP_424J2_126_3477_n2528), 
        .A2(DP_OP_425J2_127_3477_n2622), .Y(DP_OP_423J2_125_3477_n2600) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1838 ( .A1(DP_OP_422J2_124_3477_n2307), 
        .A2(DP_OP_422J2_124_3477_n2622), .Y(DP_OP_423J2_125_3477_n2599) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1837 ( .A1(DP_OP_425J2_127_3477_n2438), 
        .A2(DP_OP_424J2_126_3477_n2622), .Y(DP_OP_423J2_125_3477_n2598) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1836 ( .A1(DP_OP_423J2_125_3477_n2613), 
        .A2(DP_OP_422J2_124_3477_n2622), .Y(DP_OP_423J2_125_3477_n2597) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1835 ( .A1(DP_OP_423J2_125_3477_n2612), .A2(
        DP_OP_424J2_126_3477_n2622), .Y(DP_OP_423J2_125_3477_n2596) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1827 ( .A1(DP_OP_423J2_125_3477_n2612), .A2(
        DP_OP_423J2_125_3477_n2621), .Y(DP_OP_423J2_125_3477_n2588) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1826 ( .A1(DP_OP_423J2_125_3477_n2619), .A2(
        DP_OP_422J2_124_3477_n2620), .Y(DP_OP_423J2_125_3477_n2587) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1825 ( .A1(DP_OP_425J2_127_3477_n2442), .A2(
        DP_OP_424J2_126_3477_n2620), .Y(DP_OP_423J2_125_3477_n2586) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1824 ( .A1(DP_OP_423J2_125_3477_n2617), .A2(
        DP_OP_424J2_126_3477_n2620), .Y(DP_OP_423J2_125_3477_n2585) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1823 ( .A1(DP_OP_424J2_126_3477_n2528), .A2(
        DP_OP_425J2_127_3477_n2620), .Y(DP_OP_423J2_125_3477_n2584) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1822 ( .A1(DP_OP_422J2_124_3477_n2307), .A2(
        DP_OP_424J2_126_3477_n2620), .Y(DP_OP_423J2_125_3477_n2583) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1821 ( .A1(DP_OP_425J2_127_3477_n2438), .A2(
        DP_OP_422J2_124_3477_n2620), .Y(DP_OP_423J2_125_3477_n2582) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1820 ( .A1(DP_OP_423J2_125_3477_n2613), .A2(
        DP_OP_424J2_126_3477_n2620), .Y(DP_OP_423J2_125_3477_n2581) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1819 ( .A1(DP_OP_423J2_125_3477_n2612), 
        .A2(DP_OP_425J2_127_3477_n2620), .Y(DP_OP_423J2_125_3477_n2580) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1800 ( .A1(DP_OP_423J2_125_3477_n2569), 
        .A2(DP_OP_423J2_125_3477_n2579), .Y(DP_OP_423J2_125_3477_n2561) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1799 ( .A1(DP_OP_423J2_125_3477_n2568), .A2(
        DP_OP_423J2_125_3477_n2579), .Y(DP_OP_423J2_125_3477_n2560) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1791 ( .A1(DP_OP_423J2_125_3477_n2568), .A2(
        DP_OP_425J2_127_3477_n2578), .Y(DP_OP_423J2_125_3477_n2552) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1784 ( .A1(DP_OP_423J2_125_3477_n2569), 
        .A2(DP_OP_423J2_125_3477_n2577), .Y(DP_OP_423J2_125_3477_n2545) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1783 ( .A1(DP_OP_423J2_125_3477_n2568), .A2(
        DP_OP_423J2_125_3477_n2577), .Y(DP_OP_423J2_125_3477_n2544) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1782 ( .A1(DP_OP_423J2_125_3477_n2575), .A2(
        DP_OP_423J2_125_3477_n2576), .Y(DP_OP_423J2_125_3477_n2543) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1781 ( .A1(DP_OP_423J2_125_3477_n2574), .A2(
        DP_OP_423J2_125_3477_n2576), .Y(DP_OP_423J2_125_3477_n2542) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1780 ( .A1(DP_OP_423J2_125_3477_n2573), .A2(
        DP_OP_423J2_125_3477_n2576), .Y(DP_OP_423J2_125_3477_n2541) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1779 ( .A1(DP_OP_423J2_125_3477_n2572), .A2(
        DP_OP_423J2_125_3477_n2576), .Y(DP_OP_423J2_125_3477_n2540) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1778 ( .A1(DP_OP_423J2_125_3477_n2571), .A2(
        DP_OP_423J2_125_3477_n2576), .Y(DP_OP_423J2_125_3477_n2539) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1777 ( .A1(DP_OP_423J2_125_3477_n2570), .A2(
        DP_OP_423J2_125_3477_n2576), .Y(DP_OP_423J2_125_3477_n2538) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1776 ( .A1(DP_OP_423J2_125_3477_n2569), .A2(
        DP_OP_423J2_125_3477_n2576), .Y(DP_OP_423J2_125_3477_n2537) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1775 ( .A1(DP_OP_423J2_125_3477_n2568), 
        .A2(DP_OP_423J2_125_3477_n2576), .Y(DP_OP_423J2_125_3477_n2536) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1755 ( .A1(DP_OP_422J2_124_3477_n2392), .A2(
        DP_OP_423J2_125_3477_n2535), .Y(DP_OP_423J2_125_3477_n2516) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1747 ( .A1(DP_OP_422J2_124_3477_n2392), .A2(
        DP_OP_423J2_125_3477_n2534), .Y(DP_OP_423J2_125_3477_n2508) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1740 ( .A1(DP_OP_423J2_125_3477_n2525), 
        .A2(DP_OP_423J2_125_3477_n2533), .Y(DP_OP_423J2_125_3477_n2501) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1739 ( .A1(DP_OP_422J2_124_3477_n2392), .A2(
        DP_OP_423J2_125_3477_n2533), .Y(DP_OP_423J2_125_3477_n2500) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1738 ( .A1(DP_OP_423J2_125_3477_n2531), .A2(
        DP_OP_423J2_125_3477_n2532), .Y(DP_OP_423J2_125_3477_n2499) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1737 ( .A1(DP_OP_423J2_125_3477_n2530), .A2(
        DP_OP_423J2_125_3477_n2532), .Y(DP_OP_423J2_125_3477_n2498) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1736 ( .A1(DP_OP_423J2_125_3477_n2529), .A2(
        DP_OP_423J2_125_3477_n2532), .Y(DP_OP_423J2_125_3477_n2497) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1735 ( .A1(DP_OP_423J2_125_3477_n2528), .A2(
        DP_OP_423J2_125_3477_n2532), .Y(DP_OP_423J2_125_3477_n2496) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1734 ( .A1(DP_OP_423J2_125_3477_n2527), .A2(
        DP_OP_423J2_125_3477_n2532), .Y(DP_OP_423J2_125_3477_n2495) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1733 ( .A1(DP_OP_423J2_125_3477_n2526), .A2(
        DP_OP_423J2_125_3477_n2532), .Y(DP_OP_423J2_125_3477_n2494) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1732 ( .A1(DP_OP_423J2_125_3477_n2525), .A2(
        DP_OP_423J2_125_3477_n2532), .Y(DP_OP_423J2_125_3477_n2493) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1731 ( .A1(DP_OP_422J2_124_3477_n2392), 
        .A2(DP_OP_423J2_125_3477_n2532), .Y(DP_OP_423J2_125_3477_n2492) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1711 ( .A1(DP_OP_422J2_124_3477_n2436), .A2(
        DP_OP_423J2_125_3477_n2491), .Y(DP_OP_423J2_125_3477_n2472) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1703 ( .A1(DP_OP_422J2_124_3477_n2436), .A2(
        DP_OP_423J2_125_3477_n2490), .Y(DP_OP_423J2_125_3477_n2464) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1695 ( .A1(DP_OP_422J2_124_3477_n2436), .A2(
        DP_OP_423J2_125_3477_n2489), .Y(DP_OP_423J2_125_3477_n2456) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1694 ( .A1(DP_OP_423J2_125_3477_n2487), .A2(
        DP_OP_423J2_125_3477_n2488), .Y(DP_OP_423J2_125_3477_n2455) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1693 ( .A1(DP_OP_422J2_124_3477_n2442), .A2(
        DP_OP_423J2_125_3477_n2488), .Y(DP_OP_423J2_125_3477_n2454) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1692 ( .A1(DP_OP_422J2_124_3477_n2441), .A2(
        DP_OP_423J2_125_3477_n2488), .Y(DP_OP_423J2_125_3477_n2453) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1691 ( .A1(DP_OP_423J2_125_3477_n2484), .A2(
        DP_OP_423J2_125_3477_n2488), .Y(DP_OP_423J2_125_3477_n2452) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1690 ( .A1(DP_OP_422J2_124_3477_n2439), .A2(
        DP_OP_423J2_125_3477_n2488), .Y(DP_OP_423J2_125_3477_n2451) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1689 ( .A1(DP_OP_423J2_125_3477_n2482), .A2(
        DP_OP_423J2_125_3477_n2488), .Y(DP_OP_423J2_125_3477_n2450) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1688 ( .A1(DP_OP_423J2_125_3477_n2481), .A2(
        DP_OP_423J2_125_3477_n2488), .Y(DP_OP_423J2_125_3477_n2449) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1687 ( .A1(DP_OP_422J2_124_3477_n2436), 
        .A2(DP_OP_423J2_125_3477_n2488), .Y(DP_OP_423J2_125_3477_n2448) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1668 ( .A1(DP_OP_423J2_125_3477_n2437), 
        .A2(DP_OP_424J2_126_3477_n2447), .Y(DP_OP_423J2_125_3477_n2429) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1667 ( .A1(DP_OP_423J2_125_3477_n2436), .A2(
        DP_OP_425J2_127_3477_n2447), .Y(DP_OP_423J2_125_3477_n2428) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1659 ( .A1(DP_OP_423J2_125_3477_n2436), .A2(
        DP_OP_423J2_125_3477_n2446), .Y(DP_OP_423J2_125_3477_n2420) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1651 ( .A1(DP_OP_423J2_125_3477_n2436), .A2(
        DP_OP_423J2_125_3477_n2445), .Y(DP_OP_423J2_125_3477_n2412) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1650 ( .A1(DP_OP_422J2_124_3477_n2531), .A2(
        DP_OP_423J2_125_3477_n2444), .Y(DP_OP_423J2_125_3477_n2411) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1649 ( .A1(DP_OP_423J2_125_3477_n2442), .A2(
        DP_OP_423J2_125_3477_n2444), .Y(DP_OP_423J2_125_3477_n2410) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1648 ( .A1(DP_OP_423J2_125_3477_n2441), .A2(
        DP_OP_423J2_125_3477_n2444), .Y(DP_OP_423J2_125_3477_n2409) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1647 ( .A1(DP_OP_422J2_124_3477_n2528), .A2(
        DP_OP_423J2_125_3477_n2444), .Y(DP_OP_423J2_125_3477_n2408) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1646 ( .A1(DP_OP_423J2_125_3477_n2439), .A2(
        DP_OP_423J2_125_3477_n2444), .Y(DP_OP_423J2_125_3477_n2407) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1645 ( .A1(DP_OP_422J2_124_3477_n2526), .A2(
        DP_OP_423J2_125_3477_n2444), .Y(DP_OP_423J2_125_3477_n2406) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1644 ( .A1(DP_OP_423J2_125_3477_n2437), .A2(
        DP_OP_423J2_125_3477_n2444), .Y(DP_OP_423J2_125_3477_n2405) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1643 ( .A1(DP_OP_423J2_125_3477_n2436), 
        .A2(DP_OP_423J2_125_3477_n2444), .Y(DP_OP_423J2_125_3477_n2404) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1623 ( .A1(DP_OP_422J2_124_3477_n2568), .A2(
        DP_OP_423J2_125_3477_n2403), .Y(DP_OP_423J2_125_3477_n2384) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1615 ( .A1(DP_OP_422J2_124_3477_n2568), .A2(
        DP_OP_423J2_125_3477_n2402), .Y(DP_OP_423J2_125_3477_n2376) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1607 ( .A1(DP_OP_422J2_124_3477_n2568), .A2(
        DP_OP_423J2_125_3477_n2401), .Y(DP_OP_423J2_125_3477_n2368) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1606 ( .A1(DP_OP_422J2_124_3477_n2575), .A2(
        DP_OP_423J2_125_3477_n2400), .Y(DP_OP_423J2_125_3477_n2367) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1605 ( .A1(DP_OP_423J2_125_3477_n2398), .A2(
        DP_OP_423J2_125_3477_n2400), .Y(DP_OP_423J2_125_3477_n2366) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1604 ( .A1(DP_OP_423J2_125_3477_n2397), .A2(
        DP_OP_423J2_125_3477_n2400), .Y(DP_OP_423J2_125_3477_n2365) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1603 ( .A1(DP_OP_423J2_125_3477_n2396), .A2(
        DP_OP_423J2_125_3477_n2400), .Y(DP_OP_423J2_125_3477_n2364) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1602 ( .A1(DP_OP_422J2_124_3477_n2571), .A2(
        DP_OP_423J2_125_3477_n2400), .Y(DP_OP_423J2_125_3477_n2363) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1601 ( .A1(DP_OP_422J2_124_3477_n2570), .A2(
        DP_OP_423J2_125_3477_n2400), .Y(DP_OP_423J2_125_3477_n2362) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1600 ( .A1(DP_OP_422J2_124_3477_n2569), .A2(
        DP_OP_423J2_125_3477_n2400), .Y(DP_OP_423J2_125_3477_n2361) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1599 ( .A1(DP_OP_422J2_124_3477_n2568), 
        .A2(DP_OP_423J2_125_3477_n2400), .Y(DP_OP_423J2_125_3477_n2360) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1579 ( .A1(DP_OP_423J2_125_3477_n2348), .A2(
        DP_OP_423J2_125_3477_n2359), .Y(DP_OP_423J2_125_3477_n2340) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1571 ( .A1(DP_OP_423J2_125_3477_n2348), .A2(
        DP_OP_423J2_125_3477_n2358), .Y(DP_OP_423J2_125_3477_n2332) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1563 ( .A1(DP_OP_423J2_125_3477_n2348), .A2(
        DP_OP_423J2_125_3477_n2357), .Y(DP_OP_423J2_125_3477_n2324) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1562 ( .A1(DP_OP_423J2_125_3477_n2355), .A2(
        DP_OP_423J2_125_3477_n2356), .Y(DP_OP_423J2_125_3477_n2323) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1561 ( .A1(DP_OP_423J2_125_3477_n2354), .A2(
        DP_OP_423J2_125_3477_n2356), .Y(DP_OP_423J2_125_3477_n2322) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1560 ( .A1(DP_OP_423J2_125_3477_n2353), .A2(
        DP_OP_423J2_125_3477_n2356), .Y(DP_OP_423J2_125_3477_n2321) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1559 ( .A1(DP_OP_422J2_124_3477_n2616), .A2(
        DP_OP_423J2_125_3477_n2356), .Y(DP_OP_423J2_125_3477_n2320) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1558 ( .A1(DP_OP_423J2_125_3477_n2351), .A2(
        DP_OP_423J2_125_3477_n2356), .Y(DP_OP_423J2_125_3477_n2319) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1557 ( .A1(DP_OP_423J2_125_3477_n2350), .A2(
        DP_OP_423J2_125_3477_n2356), .Y(DP_OP_423J2_125_3477_n2318) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1556 ( .A1(DP_OP_422J2_124_3477_n2613), .A2(
        DP_OP_423J2_125_3477_n2356), .Y(DP_OP_423J2_125_3477_n2317) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1555 ( .A1(DP_OP_423J2_125_3477_n2348), 
        .A2(DP_OP_423J2_125_3477_n2356), .Y(DP_OP_423J2_125_3477_n2316) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1535 ( .A1(DP_OP_423J2_125_3477_n2304), .A2(
        DP_OP_423J2_125_3477_n2315), .Y(DP_OP_423J2_125_3477_n2296) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1527 ( .A1(DP_OP_423J2_125_3477_n2304), .A2(
        DP_OP_423J2_125_3477_n2314), .Y(DP_OP_423J2_125_3477_n2288) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1519 ( .A1(DP_OP_423J2_125_3477_n2304), .A2(
        DP_OP_423J2_125_3477_n2313), .Y(DP_OP_423J2_125_3477_n2280) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1518 ( .A1(DP_OP_423J2_125_3477_n2311), .A2(
        DP_OP_423J2_125_3477_n2312), .Y(DP_OP_423J2_125_3477_n2279) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1517 ( .A1(DP_OP_422J2_124_3477_n2662), .A2(
        DP_OP_423J2_125_3477_n2312), .Y(DP_OP_423J2_125_3477_n2278) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1516 ( .A1(DP_OP_424J2_126_3477_n2397), .A2(
        DP_OP_423J2_125_3477_n2312), .Y(DP_OP_423J2_125_3477_n2277) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1515 ( .A1(DP_OP_423J2_125_3477_n2308), .A2(
        DP_OP_423J2_125_3477_n2312), .Y(DP_OP_423J2_125_3477_n2276) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1514 ( .A1(DP_OP_423J2_125_3477_n2307), .A2(
        DP_OP_423J2_125_3477_n2312), .Y(DP_OP_423J2_125_3477_n2275) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1513 ( .A1(DP_OP_422J2_124_3477_n2658), .A2(
        DP_OP_423J2_125_3477_n2312), .Y(DP_OP_423J2_125_3477_n2274) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1512 ( .A1(DP_OP_423J2_125_3477_n2305), .A2(
        DP_OP_423J2_125_3477_n2312), .Y(DP_OP_423J2_125_3477_n2273) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1511 ( .A1(DP_OP_423J2_125_3477_n2304), 
        .A2(DP_OP_423J2_125_3477_n2312), .Y(DP_OP_423J2_125_3477_n2272) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1492 ( .A1(DP_OP_423J2_125_3477_n2261), 
        .A2(DP_OP_422J2_124_3477_n2271), .Y(DP_OP_423J2_125_3477_n2253) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1491 ( .A1(DP_OP_423J2_125_3477_n2260), .A2(
        DP_OP_424J2_126_3477_n2271), .Y(DP_OP_423J2_125_3477_n2252) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1483 ( .A1(DP_OP_423J2_125_3477_n2260), .A2(
        DP_OP_423J2_125_3477_n2270), .Y(DP_OP_423J2_125_3477_n2244) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1475 ( .A1(DP_OP_423J2_125_3477_n2260), .A2(
        DP_OP_425J2_127_3477_n2269), .Y(DP_OP_423J2_125_3477_n2236) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1474 ( .A1(DP_OP_423J2_125_3477_n2267), .A2(
        DP_OP_423J2_125_3477_n2268), .Y(DP_OP_423J2_125_3477_n2235) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1473 ( .A1(DP_OP_423J2_125_3477_n2266), .A2(
        DP_OP_423J2_125_3477_n2268), .Y(DP_OP_423J2_125_3477_n2234) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1472 ( .A1(DP_OP_423J2_125_3477_n2265), .A2(
        DP_OP_423J2_125_3477_n2268), .Y(DP_OP_423J2_125_3477_n2233) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1471 ( .A1(DP_OP_425J2_127_3477_n2572), .A2(
        DP_OP_423J2_125_3477_n2268), .Y(DP_OP_423J2_125_3477_n2232) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1470 ( .A1(DP_OP_423J2_125_3477_n2263), .A2(
        DP_OP_423J2_125_3477_n2268), .Y(DP_OP_423J2_125_3477_n2231) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1469 ( .A1(DP_OP_423J2_125_3477_n2262), .A2(
        DP_OP_423J2_125_3477_n2268), .Y(DP_OP_423J2_125_3477_n2230) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1468 ( .A1(DP_OP_423J2_125_3477_n2261), .A2(
        DP_OP_423J2_125_3477_n2268), .Y(DP_OP_423J2_125_3477_n2229) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1467 ( .A1(DP_OP_423J2_125_3477_n2260), 
        .A2(DP_OP_423J2_125_3477_n2268), .Y(DP_OP_423J2_125_3477_n2228) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1448 ( .A1(DP_OP_423J2_125_3477_n2217), 
        .A2(DP_OP_424J2_126_3477_n2227), .Y(DP_OP_423J2_125_3477_n2209) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1447 ( .A1(DP_OP_425J2_127_3477_n2612), .A2(
        DP_OP_422J2_124_3477_n2227), .Y(DP_OP_423J2_125_3477_n2208) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1440 ( .A1(DP_OP_423J2_125_3477_n2217), 
        .A2(DP_OP_423J2_125_3477_n2226), .Y(DP_OP_423J2_125_3477_n2201) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1439 ( .A1(DP_OP_425J2_127_3477_n2612), .A2(
        DP_OP_423J2_125_3477_n2226), .Y(DP_OP_423J2_125_3477_n2200) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1431 ( .A1(DP_OP_425J2_127_3477_n2612), .A2(
        DP_OP_423J2_125_3477_n2225), .Y(DP_OP_423J2_125_3477_n2192) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1430 ( .A1(DP_OP_422J2_124_3477_n2751), .A2(
        DP_OP_423J2_125_3477_n2224), .Y(DP_OP_423J2_125_3477_n2191) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1429 ( .A1(DP_OP_424J2_126_3477_n2310), .A2(
        DP_OP_423J2_125_3477_n2224), .Y(DP_OP_423J2_125_3477_n2190) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1428 ( .A1(DP_OP_425J2_127_3477_n2617), .A2(
        DP_OP_423J2_125_3477_n2224), .Y(DP_OP_423J2_125_3477_n2189) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1427 ( .A1(DP_OP_425J2_127_3477_n2616), .A2(
        DP_OP_423J2_125_3477_n2224), .Y(DP_OP_423J2_125_3477_n2188) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1426 ( .A1(DP_OP_423J2_125_3477_n2219), .A2(
        DP_OP_423J2_125_3477_n2224), .Y(DP_OP_423J2_125_3477_n2187) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1425 ( .A1(DP_OP_423J2_125_3477_n2218), .A2(
        DP_OP_423J2_125_3477_n2224), .Y(DP_OP_423J2_125_3477_n2186) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1424 ( .A1(DP_OP_423J2_125_3477_n2217), .A2(
        DP_OP_423J2_125_3477_n2224), .Y(DP_OP_423J2_125_3477_n2185) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1423 ( .A1(DP_OP_425J2_127_3477_n2612), 
        .A2(DP_OP_423J2_125_3477_n2224), .Y(DP_OP_423J2_125_3477_n2184) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1403 ( .A1(DP_OP_423J2_125_3477_n2172), .A2(
        DP_OP_423J2_125_3477_n2183), .Y(DP_OP_423J2_125_3477_n2164) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1395 ( .A1(DP_OP_423J2_125_3477_n2172), .A2(
        DP_OP_425J2_127_3477_n2182), .Y(DP_OP_423J2_125_3477_n2156) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1387 ( .A1(DP_OP_423J2_125_3477_n2172), .A2(
        DP_OP_423J2_125_3477_n2181), .Y(DP_OP_423J2_125_3477_n2148) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1386 ( .A1(DP_OP_422J2_124_3477_n2795), .A2(
        DP_OP_423J2_125_3477_n2180), .Y(DP_OP_423J2_125_3477_n2147) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1385 ( .A1(DP_OP_423J2_125_3477_n2178), .A2(
        DP_OP_423J2_125_3477_n2180), .Y(DP_OP_423J2_125_3477_n2146) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1384 ( .A1(DP_OP_422J2_124_3477_n2793), .A2(
        DP_OP_423J2_125_3477_n2180), .Y(DP_OP_423J2_125_3477_n2145) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1383 ( .A1(DP_OP_424J2_126_3477_n2264), .A2(
        DP_OP_423J2_125_3477_n2180), .Y(DP_OP_423J2_125_3477_n2144) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1382 ( .A1(DP_OP_423J2_125_3477_n2175), .A2(
        DP_OP_423J2_125_3477_n2180), .Y(DP_OP_423J2_125_3477_n2143) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1381 ( .A1(DP_OP_425J2_127_3477_n2658), .A2(
        DP_OP_423J2_125_3477_n2180), .Y(DP_OP_423J2_125_3477_n2142) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1380 ( .A1(DP_OP_424J2_126_3477_n2261), .A2(
        DP_OP_423J2_125_3477_n2180), .Y(DP_OP_423J2_125_3477_n2141) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1379 ( .A1(DP_OP_423J2_125_3477_n2172), 
        .A2(DP_OP_423J2_125_3477_n2180), .Y(DP_OP_423J2_125_3477_n2140) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1359 ( .A1(DP_OP_423J2_125_3477_n2128), .A2(
        DP_OP_423J2_125_3477_n2139), .Y(DP_OP_423J2_125_3477_n2120) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1351 ( .A1(DP_OP_423J2_125_3477_n2128), .A2(
        DP_OP_423J2_125_3477_n2138), .Y(DP_OP_423J2_125_3477_n2112) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1343 ( .A1(DP_OP_423J2_125_3477_n2128), .A2(
        DP_OP_425J2_127_3477_n2137), .Y(DP_OP_423J2_125_3477_n2104) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1342 ( .A1(DP_OP_423J2_125_3477_n2135), .A2(
        DP_OP_423J2_125_3477_n2136), .Y(DP_OP_423J2_125_3477_n2103) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1341 ( .A1(DP_OP_423J2_125_3477_n2134), .A2(
        DP_OP_423J2_125_3477_n2136), .Y(DP_OP_423J2_125_3477_n2102) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1340 ( .A1(DP_OP_425J2_127_3477_n2705), .A2(
        DP_OP_423J2_125_3477_n2136), .Y(DP_OP_423J2_125_3477_n2101) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1339 ( .A1(DP_OP_425J2_127_3477_n2704), .A2(
        DP_OP_423J2_125_3477_n2136), .Y(DP_OP_423J2_125_3477_n2100) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1338 ( .A1(DP_OP_422J2_124_3477_n2835), .A2(
        DP_OP_423J2_125_3477_n2136), .Y(DP_OP_423J2_125_3477_n2099) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1337 ( .A1(DP_OP_424J2_126_3477_n2218), .A2(
        DP_OP_423J2_125_3477_n2136), .Y(DP_OP_423J2_125_3477_n2098) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1336 ( .A1(DP_OP_424J2_126_3477_n2217), .A2(
        DP_OP_423J2_125_3477_n2136), .Y(DP_OP_423J2_125_3477_n2097) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1335 ( .A1(DP_OP_423J2_125_3477_n2128), 
        .A2(DP_OP_423J2_125_3477_n2136), .Y(DP_OP_423J2_125_3477_n2096) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1322 ( .A1(DP_OP_422J2_124_3477_n2883), 
        .A2(DP_OP_425J2_127_3477_n2095), .Y(DP_OP_423J2_125_3477_n2083) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1321 ( .A1(DP_OP_424J2_126_3477_n2178), 
        .A2(DP_OP_424J2_126_3477_n2095), .Y(DP_OP_423J2_125_3477_n2082) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1320 ( .A1(DP_OP_424J2_126_3477_n2177), 
        .A2(DP_OP_422J2_124_3477_n2095), .Y(DP_OP_423J2_125_3477_n2081) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1319 ( .A1(DP_OP_423J2_125_3477_n2088), 
        .A2(DP_OP_424J2_126_3477_n2095), .Y(DP_OP_423J2_125_3477_n2080) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1318 ( .A1(DP_OP_423J2_125_3477_n2087), 
        .A2(DP_OP_425J2_127_3477_n2095), .Y(DP_OP_423J2_125_3477_n2079) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1317 ( .A1(DP_OP_423J2_125_3477_n2086), 
        .A2(DP_OP_422J2_124_3477_n2095), .Y(DP_OP_423J2_125_3477_n2078) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1316 ( .A1(DP_OP_425J2_127_3477_n2745), 
        .A2(DP_OP_425J2_127_3477_n2095), .Y(DP_OP_423J2_125_3477_n2077) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1315 ( .A1(DP_OP_423J2_125_3477_n2084), .A2(
        DP_OP_422J2_124_3477_n2095), .Y(DP_OP_423J2_125_3477_n2076) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1314 ( .A1(DP_OP_424J2_126_3477_n2179), 
        .A2(DP_OP_425J2_127_3477_n2094), .Y(DP_OP_423J2_125_3477_n2075) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1313 ( .A1(DP_OP_425J2_127_3477_n2750), 
        .A2(DP_OP_425J2_127_3477_n2094), .Y(DP_OP_423J2_125_3477_n2074) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1312 ( .A1(DP_OP_424J2_126_3477_n2177), 
        .A2(DP_OP_422J2_124_3477_n2094), .Y(DP_OP_423J2_125_3477_n2073) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1311 ( .A1(DP_OP_423J2_125_3477_n2088), 
        .A2(DP_OP_425J2_127_3477_n2094), .Y(DP_OP_423J2_125_3477_n2072) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1310 ( .A1(DP_OP_423J2_125_3477_n2087), 
        .A2(DP_OP_422J2_124_3477_n2094), .Y(DP_OP_423J2_125_3477_n2071) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1309 ( .A1(DP_OP_423J2_125_3477_n2086), 
        .A2(DP_OP_424J2_126_3477_n2094), .Y(DP_OP_423J2_125_3477_n2070) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1308 ( .A1(DP_OP_422J2_124_3477_n2877), 
        .A2(DP_OP_424J2_126_3477_n2094), .Y(DP_OP_423J2_125_3477_n2069) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1307 ( .A1(DP_OP_423J2_125_3477_n2084), .A2(
        DP_OP_422J2_124_3477_n2094), .Y(DP_OP_423J2_125_3477_n2068) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1299 ( .A1(DP_OP_423J2_125_3477_n2084), .A2(
        DP_OP_423J2_125_3477_n2093), .Y(DP_OP_423J2_125_3477_n2060) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1298 ( .A1(DP_OP_424J2_126_3477_n2179), .A2(
        DP_OP_423J2_125_3477_n2092), .Y(DP_OP_423J2_125_3477_n2059) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1297 ( .A1(DP_OP_424J2_126_3477_n2178), .A2(
        DP_OP_423J2_125_3477_n2092), .Y(DP_OP_423J2_125_3477_n2058) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1296 ( .A1(DP_OP_424J2_126_3477_n2177), .A2(
        DP_OP_423J2_125_3477_n2092), .Y(DP_OP_423J2_125_3477_n2057) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1295 ( .A1(DP_OP_423J2_125_3477_n2088), .A2(
        DP_OP_423J2_125_3477_n2092), .Y(DP_OP_423J2_125_3477_n2056) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1294 ( .A1(DP_OP_423J2_125_3477_n2087), .A2(
        DP_OP_423J2_125_3477_n2092), .Y(DP_OP_423J2_125_3477_n2055) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1293 ( .A1(DP_OP_423J2_125_3477_n2086), .A2(
        DP_OP_423J2_125_3477_n2092), .Y(DP_OP_423J2_125_3477_n2054) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1292 ( .A1(DP_OP_422J2_124_3477_n2877), .A2(
        DP_OP_423J2_125_3477_n2092), .Y(DP_OP_423J2_125_3477_n2053) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1291 ( .A1(DP_OP_423J2_125_3477_n2084), 
        .A2(DP_OP_423J2_125_3477_n2092), .Y(DP_OP_423J2_125_3477_n2052) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1277 ( .A1(DP_OP_425J2_127_3477_n2794), 
        .A2(DP_OP_422J2_124_3477_n2051), .Y(DP_OP_423J2_125_3477_n2038) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1275 ( .A1(DP_OP_423J2_125_3477_n2044), 
        .A2(DP_OP_422J2_124_3477_n2051), .Y(DP_OP_423J2_125_3477_n2036) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1272 ( .A1(DP_OP_425J2_127_3477_n2789), 
        .A2(DP_OP_425J2_127_3477_n2051), .Y(DP_OP_423J2_125_3477_n2033) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1271 ( .A1(DP_OP_423J2_125_3477_n2040), .A2(
        DP_OP_425J2_127_3477_n2051), .Y(DP_OP_423J2_125_3477_n2032) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1263 ( .A1(DP_OP_423J2_125_3477_n2040), .A2(
        DP_OP_423J2_125_3477_n2050), .Y(DP_OP_423J2_125_3477_n2024) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1255 ( .A1(DP_OP_423J2_125_3477_n2040), .A2(
        DP_OP_425J2_127_3477_n2049), .Y(DP_OP_423J2_125_3477_n2016) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1254 ( .A1(DP_OP_425J2_127_3477_n2795), .A2(
        DP_OP_423J2_125_3477_n2048), .Y(DP_OP_423J2_125_3477_n2015) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1253 ( .A1(DP_OP_425J2_127_3477_n2794), .A2(
        DP_OP_423J2_125_3477_n2048), .Y(DP_OP_423J2_125_3477_n2014) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1252 ( .A1(DP_OP_425J2_127_3477_n2793), .A2(
        DP_OP_423J2_125_3477_n2048), .Y(DP_OP_423J2_125_3477_n2013) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1251 ( .A1(DP_OP_423J2_125_3477_n2044), .A2(
        DP_OP_423J2_125_3477_n2048), .Y(DP_OP_423J2_125_3477_n2012) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1250 ( .A1(DP_OP_425J2_127_3477_n2791), .A2(
        DP_OP_423J2_125_3477_n2048), .Y(DP_OP_423J2_125_3477_n2011) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1249 ( .A1(DP_OP_425J2_127_3477_n2790), .A2(
        DP_OP_423J2_125_3477_n2048), .Y(DP_OP_423J2_125_3477_n2010) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1248 ( .A1(DP_OP_425J2_127_3477_n2789), .A2(
        DP_OP_423J2_125_3477_n2048), .Y(DP_OP_423J2_125_3477_n2009) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1247 ( .A1(DP_OP_423J2_125_3477_n2040), 
        .A2(DP_OP_423J2_125_3477_n2048), .Y(DP_OP_423J2_125_3477_n2008) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1227 ( .A1(DP_OP_424J2_126_3477_n2084), .A2(
        DP_OP_423J2_125_3477_n2007), .Y(DP_OP_423J2_125_3477_n1988) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1219 ( .A1(DP_OP_422J2_124_3477_n2964), .A2(
        DP_OP_423J2_125_3477_n2006), .Y(DP_OP_423J2_125_3477_n1980) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1212 ( .A1(DP_OP_423J2_125_3477_n1997), 
        .A2(DP_OP_423J2_125_3477_n2005), .Y(DP_OP_423J2_125_3477_n1973) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1211 ( .A1(DP_OP_424J2_126_3477_n2084), .A2(
        DP_OP_423J2_125_3477_n2005), .Y(DP_OP_423J2_125_3477_n1972) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1210 ( .A1(DP_OP_423J2_125_3477_n2003), .A2(
        DP_OP_423J2_125_3477_n2004), .Y(DP_OP_423J2_125_3477_n1971) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1209 ( .A1(DP_OP_424J2_126_3477_n2090), .A2(
        DP_OP_423J2_125_3477_n2004), .Y(DP_OP_423J2_125_3477_n1970) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1208 ( .A1(DP_OP_422J2_124_3477_n2969), .A2(
        DP_OP_423J2_125_3477_n2004), .Y(DP_OP_423J2_125_3477_n1969) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1207 ( .A1(DP_OP_423J2_125_3477_n2000), .A2(
        DP_OP_423J2_125_3477_n2004), .Y(DP_OP_423J2_125_3477_n1968) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1206 ( .A1(DP_OP_424J2_126_3477_n2087), .A2(
        DP_OP_423J2_125_3477_n2004), .Y(DP_OP_423J2_125_3477_n1967) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1205 ( .A1(DP_OP_423J2_125_3477_n1998), .A2(
        DP_OP_423J2_125_3477_n2004), .Y(DP_OP_423J2_125_3477_n1966) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1204 ( .A1(DP_OP_423J2_125_3477_n1997), .A2(
        DP_OP_423J2_125_3477_n2004), .Y(DP_OP_423J2_125_3477_n1965) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1203 ( .A1(DP_OP_422J2_124_3477_n2964), 
        .A2(DP_OP_423J2_125_3477_n2004), .Y(DP_OP_423J2_125_3477_n1964) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1184 ( .A1(DP_OP_422J2_124_3477_n3007), 
        .A2(DP_OP_423J2_125_3477_n1963), .Y(DP_OP_423J2_125_3477_n1945) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1183 ( .A1(DP_OP_423J2_125_3477_n1952), .A2(
        DP_OP_423J2_125_3477_n1963), .Y(DP_OP_423J2_125_3477_n1944) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1176 ( .A1(DP_OP_422J2_124_3477_n3007), 
        .A2(DP_OP_423J2_125_3477_n1962), .Y(DP_OP_423J2_125_3477_n1937) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1175 ( .A1(DP_OP_423J2_125_3477_n1952), .A2(
        DP_OP_423J2_125_3477_n1962), .Y(DP_OP_423J2_125_3477_n1936) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1167 ( .A1(DP_OP_423J2_125_3477_n1952), .A2(
        DP_OP_425J2_127_3477_n1961), .Y(DP_OP_423J2_125_3477_n1928) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1166 ( .A1(DP_OP_424J2_126_3477_n2047), .A2(
        DP_OP_423J2_125_3477_n1960), .Y(DP_OP_423J2_125_3477_n1927) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1165 ( .A1(DP_OP_423J2_125_3477_n1958), .A2(
        DP_OP_423J2_125_3477_n1960), .Y(DP_OP_423J2_125_3477_n1926) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1164 ( .A1(DP_OP_423J2_125_3477_n1957), .A2(
        DP_OP_423J2_125_3477_n1960), .Y(DP_OP_423J2_125_3477_n1925) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1163 ( .A1(DP_OP_424J2_126_3477_n2044), .A2(
        DP_OP_423J2_125_3477_n1960), .Y(DP_OP_423J2_125_3477_n1924) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1162 ( .A1(DP_OP_422J2_124_3477_n3009), .A2(
        DP_OP_423J2_125_3477_n1960), .Y(DP_OP_423J2_125_3477_n1923) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1161 ( .A1(DP_OP_425J2_127_3477_n2878), .A2(
        DP_OP_423J2_125_3477_n1960), .Y(DP_OP_423J2_125_3477_n1922) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1160 ( .A1(DP_OP_425J2_127_3477_n2877), .A2(
        DP_OP_423J2_125_3477_n1960), .Y(DP_OP_423J2_125_3477_n1921) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1159 ( .A1(DP_OP_423J2_125_3477_n1952), 
        .A2(DP_OP_423J2_125_3477_n1960), .Y(DP_OP_423J2_125_3477_n1920) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1115 ( .A1(n336), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_423J2_125_3477_n460) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1114 ( .A1(n322), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_423J2_125_3477_n1876) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1112 ( .A1(n367), .A2(n391), .Y(
        DP_OP_423J2_125_3477_n1874) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1110 ( .A1(n351), .A2(n388), .Y(
        DP_OP_423J2_125_3477_n1873) );
  HADDX1_HVT DP_OP_423J2_125_3477_U1093 ( .A0(DP_OP_423J2_125_3477_n1886), 
        .B0(DP_OP_423J2_125_3477_n1995), .C1(DP_OP_423J2_125_3477_n1870), .SO(
        DP_OP_423J2_125_3477_n1871) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1092 ( .A(DP_OP_423J2_125_3477_n2039), .B(
        DP_OP_423J2_125_3477_n1951), .CI(DP_OP_423J2_125_3477_n2083), .CO(
        DP_OP_423J2_125_3477_n1868), .S(DP_OP_423J2_125_3477_n1869) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1091 ( .A(DP_OP_423J2_125_3477_n2171), .B(
        DP_OP_423J2_125_3477_n2127), .CI(DP_OP_423J2_125_3477_n2215), .CO(
        DP_OP_423J2_125_3477_n1866), .S(DP_OP_423J2_125_3477_n1867) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1090 ( .A(DP_OP_423J2_125_3477_n2303), .B(
        DP_OP_423J2_125_3477_n2259), .CI(DP_OP_423J2_125_3477_n2347), .CO(
        DP_OP_423J2_125_3477_n1864), .S(DP_OP_423J2_125_3477_n1865) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1089 ( .A(DP_OP_423J2_125_3477_n2435), .B(
        DP_OP_423J2_125_3477_n2391), .CI(DP_OP_423J2_125_3477_n2479), .CO(
        DP_OP_423J2_125_3477_n1862), .S(DP_OP_423J2_125_3477_n1863) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1088 ( .A(DP_OP_423J2_125_3477_n2567), .B(
        DP_OP_423J2_125_3477_n2523), .CI(DP_OP_423J2_125_3477_n2611), .CO(
        DP_OP_423J2_125_3477_n1860), .S(DP_OP_423J2_125_3477_n1861) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1087 ( .A(DP_OP_423J2_125_3477_n2699), .B(
        DP_OP_423J2_125_3477_n2655), .CI(DP_OP_423J2_125_3477_n2743), .CO(
        DP_OP_423J2_125_3477_n1858), .S(DP_OP_423J2_125_3477_n1859) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1086 ( .A(DP_OP_423J2_125_3477_n3005), .B(
        DP_OP_423J2_125_3477_n2787), .CI(DP_OP_423J2_125_3477_n2831), .CO(
        DP_OP_423J2_125_3477_n1856), .S(DP_OP_423J2_125_3477_n1857) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1085 ( .A(DP_OP_423J2_125_3477_n2963), .B(
        DP_OP_423J2_125_3477_n2875), .CI(DP_OP_423J2_125_3477_n2919), .CO(
        DP_OP_423J2_125_3477_n1854), .S(DP_OP_423J2_125_3477_n1855) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1084 ( .A(DP_OP_423J2_125_3477_n1871), .B(
        DP_OP_423J2_125_3477_n1857), .CI(DP_OP_423J2_125_3477_n1859), .CO(
        DP_OP_423J2_125_3477_n1852), .S(DP_OP_423J2_125_3477_n1853) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1083 ( .A(DP_OP_423J2_125_3477_n1861), .B(
        DP_OP_423J2_125_3477_n1855), .CI(DP_OP_423J2_125_3477_n1863), .CO(
        DP_OP_423J2_125_3477_n1850), .S(DP_OP_423J2_125_3477_n1851) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1082 ( .A(DP_OP_423J2_125_3477_n1869), .B(
        DP_OP_423J2_125_3477_n1865), .CI(DP_OP_423J2_125_3477_n1867), .CO(
        DP_OP_423J2_125_3477_n1848), .S(DP_OP_423J2_125_3477_n1849) );
  HADDX1_HVT DP_OP_423J2_125_3477_U1081 ( .A0(DP_OP_423J2_125_3477_n1885), 
        .B0(DP_OP_423J2_125_3477_n1950), .C1(DP_OP_423J2_125_3477_n1846), .SO(
        DP_OP_423J2_125_3477_n1847) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1080 ( .A(DP_OP_423J2_125_3477_n1987), .B(
        DP_OP_423J2_125_3477_n1943), .CI(DP_OP_423J2_125_3477_n1994), .CO(
        DP_OP_423J2_125_3477_n1844), .S(DP_OP_423J2_125_3477_n1845) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1079 ( .A(DP_OP_423J2_125_3477_n2038), .B(
        DP_OP_423J2_125_3477_n2031), .CI(DP_OP_423J2_125_3477_n2075), .CO(
        DP_OP_423J2_125_3477_n1842), .S(DP_OP_423J2_125_3477_n1843) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1078 ( .A(DP_OP_423J2_125_3477_n2119), .B(
        DP_OP_423J2_125_3477_n2082), .CI(DP_OP_423J2_125_3477_n2126), .CO(
        DP_OP_423J2_125_3477_n1840), .S(DP_OP_423J2_125_3477_n1841) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1077 ( .A(DP_OP_423J2_125_3477_n2170), .B(
        DP_OP_423J2_125_3477_n2163), .CI(DP_OP_423J2_125_3477_n2207), .CO(
        DP_OP_423J2_125_3477_n1838), .S(DP_OP_423J2_125_3477_n1839) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1076 ( .A(DP_OP_423J2_125_3477_n2251), .B(
        DP_OP_423J2_125_3477_n2214), .CI(DP_OP_423J2_125_3477_n2258), .CO(
        DP_OP_423J2_125_3477_n1836), .S(DP_OP_423J2_125_3477_n1837) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1075 ( .A(DP_OP_423J2_125_3477_n2302), .B(
        DP_OP_423J2_125_3477_n2295), .CI(DP_OP_423J2_125_3477_n2339), .CO(
        DP_OP_423J2_125_3477_n1834), .S(DP_OP_423J2_125_3477_n1835) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1074 ( .A(DP_OP_423J2_125_3477_n2383), .B(
        DP_OP_423J2_125_3477_n2346), .CI(DP_OP_423J2_125_3477_n2390), .CO(
        DP_OP_423J2_125_3477_n1832), .S(DP_OP_423J2_125_3477_n1833) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1073 ( .A(DP_OP_423J2_125_3477_n2434), .B(
        DP_OP_423J2_125_3477_n2427), .CI(DP_OP_423J2_125_3477_n2471), .CO(
        DP_OP_423J2_125_3477_n1830), .S(DP_OP_423J2_125_3477_n1831) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1072 ( .A(DP_OP_423J2_125_3477_n2515), .B(
        DP_OP_423J2_125_3477_n2478), .CI(DP_OP_423J2_125_3477_n2522), .CO(
        DP_OP_423J2_125_3477_n1828), .S(DP_OP_423J2_125_3477_n1829) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1071 ( .A(DP_OP_423J2_125_3477_n3004), .B(
        DP_OP_423J2_125_3477_n2559), .CI(DP_OP_423J2_125_3477_n2997), .CO(
        DP_OP_423J2_125_3477_n1826), .S(DP_OP_423J2_125_3477_n1827) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1070 ( .A(DP_OP_423J2_125_3477_n2742), .B(
        DP_OP_423J2_125_3477_n2566), .CI(DP_OP_423J2_125_3477_n2603), .CO(
        DP_OP_423J2_125_3477_n1824), .S(DP_OP_423J2_125_3477_n1825) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1069 ( .A(DP_OP_423J2_125_3477_n2779), .B(
        DP_OP_423J2_125_3477_n2962), .CI(DP_OP_423J2_125_3477_n2955), .CO(
        DP_OP_423J2_125_3477_n1822), .S(DP_OP_423J2_125_3477_n1823) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1068 ( .A(DP_OP_423J2_125_3477_n2698), .B(
        DP_OP_423J2_125_3477_n2918), .CI(DP_OP_423J2_125_3477_n2911), .CO(
        DP_OP_423J2_125_3477_n1820), .S(DP_OP_423J2_125_3477_n1821) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1067 ( .A(DP_OP_423J2_125_3477_n2691), .B(
        DP_OP_423J2_125_3477_n2874), .CI(DP_OP_423J2_125_3477_n2610), .CO(
        DP_OP_423J2_125_3477_n1818), .S(DP_OP_423J2_125_3477_n1819) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1066 ( .A(DP_OP_423J2_125_3477_n2867), .B(
        DP_OP_423J2_125_3477_n2647), .CI(DP_OP_423J2_125_3477_n2654), .CO(
        DP_OP_423J2_125_3477_n1816), .S(DP_OP_423J2_125_3477_n1817) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1065 ( .A(DP_OP_423J2_125_3477_n2823), .B(
        DP_OP_423J2_125_3477_n2735), .CI(DP_OP_423J2_125_3477_n2786), .CO(
        DP_OP_423J2_125_3477_n1814), .S(DP_OP_423J2_125_3477_n1815) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1064 ( .A(DP_OP_423J2_125_3477_n2830), .B(
        DP_OP_423J2_125_3477_n1870), .CI(DP_OP_423J2_125_3477_n1847), .CO(
        DP_OP_423J2_125_3477_n1812), .S(DP_OP_423J2_125_3477_n1813) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1063 ( .A(DP_OP_423J2_125_3477_n1854), .B(
        DP_OP_423J2_125_3477_n1868), .CI(DP_OP_423J2_125_3477_n1866), .CO(
        DP_OP_423J2_125_3477_n1810), .S(DP_OP_423J2_125_3477_n1811) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1062 ( .A(DP_OP_423J2_125_3477_n1860), .B(
        DP_OP_423J2_125_3477_n1856), .CI(DP_OP_423J2_125_3477_n1864), .CO(
        DP_OP_423J2_125_3477_n1808), .S(DP_OP_423J2_125_3477_n1809) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1061 ( .A(DP_OP_423J2_125_3477_n1862), .B(
        DP_OP_423J2_125_3477_n1858), .CI(DP_OP_423J2_125_3477_n1815), .CO(
        DP_OP_423J2_125_3477_n1806), .S(DP_OP_423J2_125_3477_n1807) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1060 ( .A(DP_OP_423J2_125_3477_n1837), .B(
        DP_OP_423J2_125_3477_n1823), .CI(DP_OP_423J2_125_3477_n1821), .CO(
        DP_OP_423J2_125_3477_n1804), .S(DP_OP_423J2_125_3477_n1805) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1059 ( .A(DP_OP_423J2_125_3477_n1841), .B(
        DP_OP_423J2_125_3477_n1825), .CI(DP_OP_423J2_125_3477_n1829), .CO(
        DP_OP_423J2_125_3477_n1802), .S(DP_OP_423J2_125_3477_n1803) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1058 ( .A(DP_OP_423J2_125_3477_n1843), .B(
        DP_OP_423J2_125_3477_n1831), .CI(DP_OP_423J2_125_3477_n1827), .CO(
        DP_OP_423J2_125_3477_n1800), .S(DP_OP_423J2_125_3477_n1801) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1057 ( .A(DP_OP_423J2_125_3477_n1845), .B(
        DP_OP_423J2_125_3477_n1835), .CI(DP_OP_423J2_125_3477_n1819), .CO(
        DP_OP_423J2_125_3477_n1798), .S(DP_OP_423J2_125_3477_n1799) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1056 ( .A(DP_OP_423J2_125_3477_n1839), .B(
        DP_OP_423J2_125_3477_n1833), .CI(DP_OP_423J2_125_3477_n1817), .CO(
        DP_OP_423J2_125_3477_n1796), .S(DP_OP_423J2_125_3477_n1797) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1055 ( .A(DP_OP_423J2_125_3477_n1813), .B(
        DP_OP_423J2_125_3477_n1852), .CI(DP_OP_423J2_125_3477_n1850), .CO(
        DP_OP_423J2_125_3477_n1794), .S(DP_OP_423J2_125_3477_n1795) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1054 ( .A(DP_OP_423J2_125_3477_n1848), .B(
        DP_OP_423J2_125_3477_n1809), .CI(DP_OP_423J2_125_3477_n1811), .CO(
        DP_OP_423J2_125_3477_n1792), .S(DP_OP_423J2_125_3477_n1793) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1053 ( .A(DP_OP_423J2_125_3477_n1807), .B(
        DP_OP_423J2_125_3477_n1799), .CI(DP_OP_423J2_125_3477_n1801), .CO(
        DP_OP_423J2_125_3477_n1790), .S(DP_OP_423J2_125_3477_n1791) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1052 ( .A(DP_OP_423J2_125_3477_n1805), .B(
        DP_OP_423J2_125_3477_n1797), .CI(DP_OP_423J2_125_3477_n1803), .CO(
        DP_OP_423J2_125_3477_n1788), .S(DP_OP_423J2_125_3477_n1789) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1051 ( .A(DP_OP_423J2_125_3477_n1795), .B(
        DP_OP_423J2_125_3477_n1793), .CI(DP_OP_423J2_125_3477_n1791), .CO(
        DP_OP_423J2_125_3477_n1786), .S(DP_OP_423J2_125_3477_n1787) );
  HADDX1_HVT DP_OP_423J2_125_3477_U1050 ( .A0(DP_OP_423J2_125_3477_n1884), 
        .B0(DP_OP_423J2_125_3477_n1949), .C1(DP_OP_423J2_125_3477_n1784), .SO(
        DP_OP_423J2_125_3477_n1785) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1049 ( .A(DP_OP_423J2_125_3477_n1979), .B(
        DP_OP_423J2_125_3477_n1942), .CI(DP_OP_423J2_125_3477_n1935), .CO(
        DP_OP_423J2_125_3477_n1782), .S(DP_OP_423J2_125_3477_n1783) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1048 ( .A(DP_OP_423J2_125_3477_n1993), .B(
        DP_OP_423J2_125_3477_n1986), .CI(DP_OP_423J2_125_3477_n2023), .CO(
        DP_OP_423J2_125_3477_n1780), .S(DP_OP_423J2_125_3477_n1781) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1047 ( .A(DP_OP_423J2_125_3477_n2037), .B(
        DP_OP_423J2_125_3477_n2030), .CI(DP_OP_423J2_125_3477_n2067), .CO(
        DP_OP_423J2_125_3477_n1778), .S(DP_OP_423J2_125_3477_n1779) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1046 ( .A(DP_OP_423J2_125_3477_n2081), .B(
        DP_OP_423J2_125_3477_n2074), .CI(DP_OP_423J2_125_3477_n2111), .CO(
        DP_OP_423J2_125_3477_n1776), .S(DP_OP_423J2_125_3477_n1777) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1045 ( .A(DP_OP_423J2_125_3477_n2125), .B(
        DP_OP_423J2_125_3477_n2118), .CI(DP_OP_423J2_125_3477_n2155), .CO(
        DP_OP_423J2_125_3477_n1774), .S(DP_OP_423J2_125_3477_n1775) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1044 ( .A(DP_OP_423J2_125_3477_n2169), .B(
        DP_OP_423J2_125_3477_n2162), .CI(DP_OP_423J2_125_3477_n2199), .CO(
        DP_OP_423J2_125_3477_n1772), .S(DP_OP_423J2_125_3477_n1773) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1043 ( .A(DP_OP_423J2_125_3477_n2213), .B(
        DP_OP_423J2_125_3477_n2206), .CI(DP_OP_423J2_125_3477_n2243), .CO(
        DP_OP_423J2_125_3477_n1770), .S(DP_OP_423J2_125_3477_n1771) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1042 ( .A(DP_OP_423J2_125_3477_n2257), .B(
        DP_OP_423J2_125_3477_n2250), .CI(DP_OP_423J2_125_3477_n2287), .CO(
        DP_OP_423J2_125_3477_n1768), .S(DP_OP_423J2_125_3477_n1769) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1041 ( .A(DP_OP_423J2_125_3477_n2301), .B(
        DP_OP_423J2_125_3477_n2294), .CI(DP_OP_423J2_125_3477_n2331), .CO(
        DP_OP_423J2_125_3477_n1766), .S(DP_OP_423J2_125_3477_n1767) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1040 ( .A(DP_OP_423J2_125_3477_n2345), .B(
        DP_OP_423J2_125_3477_n2338), .CI(DP_OP_423J2_125_3477_n2375), .CO(
        DP_OP_423J2_125_3477_n1764), .S(DP_OP_423J2_125_3477_n1765) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1039 ( .A(DP_OP_423J2_125_3477_n2389), .B(
        DP_OP_423J2_125_3477_n2382), .CI(DP_OP_423J2_125_3477_n2419), .CO(
        DP_OP_423J2_125_3477_n1762), .S(DP_OP_423J2_125_3477_n1763) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1038 ( .A(DP_OP_423J2_125_3477_n2690), .B(
        DP_OP_423J2_125_3477_n3003), .CI(DP_OP_423J2_125_3477_n2996), .CO(
        DP_OP_423J2_125_3477_n1760), .S(DP_OP_423J2_125_3477_n1761) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1037 ( .A(DP_OP_423J2_125_3477_n2653), .B(
        DP_OP_423J2_125_3477_n2426), .CI(DP_OP_423J2_125_3477_n2989), .CO(
        DP_OP_423J2_125_3477_n1758), .S(DP_OP_423J2_125_3477_n1759) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1036 ( .A(DP_OP_423J2_125_3477_n2646), .B(
        DP_OP_423J2_125_3477_n2961), .CI(DP_OP_423J2_125_3477_n2433), .CO(
        DP_OP_423J2_125_3477_n1756), .S(DP_OP_423J2_125_3477_n1757) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1035 ( .A(DP_OP_423J2_125_3477_n2683), .B(
        DP_OP_423J2_125_3477_n2463), .CI(DP_OP_423J2_125_3477_n2470), .CO(
        DP_OP_423J2_125_3477_n1754), .S(DP_OP_423J2_125_3477_n1755) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1034 ( .A(DP_OP_423J2_125_3477_n2697), .B(
        DP_OP_423J2_125_3477_n2477), .CI(DP_OP_423J2_125_3477_n2954), .CO(
        DP_OP_423J2_125_3477_n1752), .S(DP_OP_423J2_125_3477_n1753) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1033 ( .A(DP_OP_423J2_125_3477_n2727), .B(
        DP_OP_423J2_125_3477_n2507), .CI(DP_OP_423J2_125_3477_n2947), .CO(
        DP_OP_423J2_125_3477_n1750), .S(DP_OP_423J2_125_3477_n1751) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1032 ( .A(DP_OP_423J2_125_3477_n2639), .B(
        DP_OP_423J2_125_3477_n2514), .CI(DP_OP_423J2_125_3477_n2917), .CO(
        DP_OP_423J2_125_3477_n1748), .S(DP_OP_423J2_125_3477_n1749) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1031 ( .A(DP_OP_423J2_125_3477_n2609), .B(
        DP_OP_423J2_125_3477_n2521), .CI(DP_OP_423J2_125_3477_n2910), .CO(
        DP_OP_423J2_125_3477_n1746), .S(DP_OP_423J2_125_3477_n1747) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1030 ( .A(DP_OP_423J2_125_3477_n2903), .B(
        DP_OP_423J2_125_3477_n2551), .CI(DP_OP_423J2_125_3477_n2558), .CO(
        DP_OP_423J2_125_3477_n1744), .S(DP_OP_423J2_125_3477_n1745) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1029 ( .A(DP_OP_423J2_125_3477_n2873), .B(
        DP_OP_423J2_125_3477_n2565), .CI(DP_OP_423J2_125_3477_n2595), .CO(
        DP_OP_423J2_125_3477_n1742), .S(DP_OP_423J2_125_3477_n1743) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1028 ( .A(DP_OP_423J2_125_3477_n2866), .B(
        DP_OP_423J2_125_3477_n2602), .CI(DP_OP_423J2_125_3477_n2734), .CO(
        DP_OP_423J2_125_3477_n1740), .S(DP_OP_423J2_125_3477_n1741) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1027 ( .A(DP_OP_423J2_125_3477_n2859), .B(
        DP_OP_423J2_125_3477_n2741), .CI(DP_OP_423J2_125_3477_n2771), .CO(
        DP_OP_423J2_125_3477_n1738), .S(DP_OP_423J2_125_3477_n1739) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1026 ( .A(DP_OP_423J2_125_3477_n2829), .B(
        DP_OP_423J2_125_3477_n2778), .CI(DP_OP_423J2_125_3477_n2785), .CO(
        DP_OP_423J2_125_3477_n1736), .S(DP_OP_423J2_125_3477_n1737) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1025 ( .A(DP_OP_423J2_125_3477_n2822), .B(
        DP_OP_423J2_125_3477_n2815), .CI(DP_OP_423J2_125_3477_n1846), .CO(
        DP_OP_423J2_125_3477_n1734), .S(DP_OP_423J2_125_3477_n1735) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1024 ( .A(DP_OP_423J2_125_3477_n1785), .B(
        DP_OP_423J2_125_3477_n1814), .CI(DP_OP_423J2_125_3477_n1816), .CO(
        DP_OP_423J2_125_3477_n1732), .S(DP_OP_423J2_125_3477_n1733) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1023 ( .A(DP_OP_423J2_125_3477_n1832), .B(
        DP_OP_423J2_125_3477_n1844), .CI(DP_OP_423J2_125_3477_n1818), .CO(
        DP_OP_423J2_125_3477_n1730), .S(DP_OP_423J2_125_3477_n1731) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1022 ( .A(DP_OP_423J2_125_3477_n1830), .B(
        DP_OP_423J2_125_3477_n1842), .CI(DP_OP_423J2_125_3477_n1820), .CO(
        DP_OP_423J2_125_3477_n1728), .S(DP_OP_423J2_125_3477_n1729) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1021 ( .A(DP_OP_423J2_125_3477_n1826), .B(
        DP_OP_423J2_125_3477_n1840), .CI(DP_OP_423J2_125_3477_n1822), .CO(
        DP_OP_423J2_125_3477_n1726), .S(DP_OP_423J2_125_3477_n1727) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1020 ( .A(DP_OP_423J2_125_3477_n1838), .B(
        DP_OP_423J2_125_3477_n1836), .CI(DP_OP_423J2_125_3477_n1834), .CO(
        DP_OP_423J2_125_3477_n1724), .S(DP_OP_423J2_125_3477_n1725) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1019 ( .A(DP_OP_423J2_125_3477_n1828), .B(
        DP_OP_423J2_125_3477_n1824), .CI(DP_OP_423J2_125_3477_n1757), .CO(
        DP_OP_423J2_125_3477_n1722), .S(DP_OP_423J2_125_3477_n1723) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1018 ( .A(DP_OP_423J2_125_3477_n1751), .B(
        DP_OP_423J2_125_3477_n1765), .CI(DP_OP_423J2_125_3477_n1769), .CO(
        DP_OP_423J2_125_3477_n1720), .S(DP_OP_423J2_125_3477_n1721) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1017 ( .A(DP_OP_423J2_125_3477_n1747), .B(
        DP_OP_423J2_125_3477_n1775), .CI(DP_OP_423J2_125_3477_n1777), .CO(
        DP_OP_423J2_125_3477_n1718), .S(DP_OP_423J2_125_3477_n1719) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1016 ( .A(DP_OP_423J2_125_3477_n1745), .B(
        DP_OP_423J2_125_3477_n1767), .CI(DP_OP_423J2_125_3477_n1781), .CO(
        DP_OP_423J2_125_3477_n1716), .S(DP_OP_423J2_125_3477_n1717) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1015 ( .A(DP_OP_423J2_125_3477_n1743), .B(
        DP_OP_423J2_125_3477_n1761), .CI(DP_OP_423J2_125_3477_n1779), .CO(
        DP_OP_423J2_125_3477_n1714), .S(DP_OP_423J2_125_3477_n1715) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1014 ( .A(DP_OP_423J2_125_3477_n1741), .B(
        DP_OP_423J2_125_3477_n1771), .CI(DP_OP_423J2_125_3477_n1759), .CO(
        DP_OP_423J2_125_3477_n1712), .S(DP_OP_423J2_125_3477_n1713) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1013 ( .A(DP_OP_423J2_125_3477_n1739), .B(
        DP_OP_423J2_125_3477_n1773), .CI(DP_OP_423J2_125_3477_n1783), .CO(
        DP_OP_423J2_125_3477_n1710), .S(DP_OP_423J2_125_3477_n1711) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1012 ( .A(DP_OP_423J2_125_3477_n1737), .B(
        DP_OP_423J2_125_3477_n1763), .CI(DP_OP_423J2_125_3477_n1749), .CO(
        DP_OP_423J2_125_3477_n1708), .S(DP_OP_423J2_125_3477_n1709) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1011 ( .A(DP_OP_423J2_125_3477_n1755), .B(
        DP_OP_423J2_125_3477_n1753), .CI(DP_OP_423J2_125_3477_n1812), .CO(
        DP_OP_423J2_125_3477_n1706), .S(DP_OP_423J2_125_3477_n1707) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1010 ( .A(DP_OP_423J2_125_3477_n1735), .B(
        DP_OP_423J2_125_3477_n1810), .CI(DP_OP_423J2_125_3477_n1808), .CO(
        DP_OP_423J2_125_3477_n1704), .S(DP_OP_423J2_125_3477_n1705) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1009 ( .A(DP_OP_423J2_125_3477_n1806), .B(
        DP_OP_423J2_125_3477_n1733), .CI(DP_OP_423J2_125_3477_n1800), .CO(
        DP_OP_423J2_125_3477_n1702), .S(DP_OP_423J2_125_3477_n1703) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1008 ( .A(DP_OP_423J2_125_3477_n1804), .B(
        DP_OP_423J2_125_3477_n1725), .CI(DP_OP_423J2_125_3477_n1731), .CO(
        DP_OP_423J2_125_3477_n1700), .S(DP_OP_423J2_125_3477_n1701) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1007 ( .A(DP_OP_423J2_125_3477_n1802), .B(
        DP_OP_423J2_125_3477_n1729), .CI(DP_OP_423J2_125_3477_n1727), .CO(
        DP_OP_423J2_125_3477_n1698), .S(DP_OP_423J2_125_3477_n1699) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1006 ( .A(DP_OP_423J2_125_3477_n1798), .B(
        DP_OP_423J2_125_3477_n1796), .CI(DP_OP_423J2_125_3477_n1723), .CO(
        DP_OP_423J2_125_3477_n1696), .S(DP_OP_423J2_125_3477_n1697) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1005 ( .A(DP_OP_423J2_125_3477_n1721), .B(
        DP_OP_423J2_125_3477_n1709), .CI(DP_OP_423J2_125_3477_n1707), .CO(
        DP_OP_423J2_125_3477_n1694), .S(DP_OP_423J2_125_3477_n1695) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1004 ( .A(DP_OP_423J2_125_3477_n1711), .B(
        DP_OP_423J2_125_3477_n1719), .CI(DP_OP_423J2_125_3477_n1717), .CO(
        DP_OP_423J2_125_3477_n1692), .S(DP_OP_423J2_125_3477_n1693) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1003 ( .A(DP_OP_423J2_125_3477_n1713), .B(
        DP_OP_423J2_125_3477_n1715), .CI(DP_OP_423J2_125_3477_n1794), .CO(
        DP_OP_423J2_125_3477_n1690), .S(DP_OP_423J2_125_3477_n1691) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1002 ( .A(DP_OP_423J2_125_3477_n1705), .B(
        DP_OP_423J2_125_3477_n1792), .CI(DP_OP_423J2_125_3477_n1703), .CO(
        DP_OP_423J2_125_3477_n1688), .S(DP_OP_423J2_125_3477_n1689) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1001 ( .A(DP_OP_423J2_125_3477_n1790), .B(
        DP_OP_423J2_125_3477_n1788), .CI(DP_OP_423J2_125_3477_n1699), .CO(
        DP_OP_423J2_125_3477_n1686), .S(DP_OP_423J2_125_3477_n1687) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1000 ( .A(DP_OP_423J2_125_3477_n1701), .B(
        DP_OP_423J2_125_3477_n1697), .CI(DP_OP_423J2_125_3477_n1695), .CO(
        DP_OP_423J2_125_3477_n1684), .S(DP_OP_423J2_125_3477_n1685) );
  FADDX1_HVT DP_OP_423J2_125_3477_U999 ( .A(DP_OP_423J2_125_3477_n1693), .B(
        DP_OP_423J2_125_3477_n1691), .CI(DP_OP_423J2_125_3477_n1689), .CO(
        DP_OP_423J2_125_3477_n1682), .S(DP_OP_423J2_125_3477_n1683) );
  FADDX1_HVT DP_OP_423J2_125_3477_U998 ( .A(DP_OP_423J2_125_3477_n1786), .B(
        DP_OP_423J2_125_3477_n1687), .CI(DP_OP_423J2_125_3477_n1685), .CO(
        DP_OP_423J2_125_3477_n1680), .S(DP_OP_423J2_125_3477_n1681) );
  FADDX1_HVT DP_OP_423J2_125_3477_U996 ( .A(DP_OP_423J2_125_3477_n2455), .B(
        DP_OP_423J2_125_3477_n1927), .CI(DP_OP_423J2_125_3477_n1883), .CO(
        DP_OP_423J2_125_3477_n1676), .S(DP_OP_423J2_125_3477_n1677) );
  FADDX1_HVT DP_OP_423J2_125_3477_U995 ( .A(DP_OP_423J2_125_3477_n2147), .B(
        DP_OP_423J2_125_3477_n2587), .CI(DP_OP_423J2_125_3477_n2367), .CO(
        DP_OP_423J2_125_3477_n1674), .S(DP_OP_423J2_125_3477_n1675) );
  FADDX1_HVT DP_OP_423J2_125_3477_U994 ( .A(DP_OP_423J2_125_3477_n2895), .B(
        DP_OP_423J2_125_3477_n2103), .CI(DP_OP_423J2_125_3477_n2323), .CO(
        DP_OP_423J2_125_3477_n1672), .S(DP_OP_423J2_125_3477_n1673) );
  FADDX1_HVT DP_OP_423J2_125_3477_U993 ( .A(DP_OP_423J2_125_3477_n2499), .B(
        DP_OP_423J2_125_3477_n2807), .CI(DP_OP_423J2_125_3477_n2411), .CO(
        DP_OP_423J2_125_3477_n1670), .S(DP_OP_423J2_125_3477_n1671) );
  FADDX1_HVT DP_OP_423J2_125_3477_U992 ( .A(DP_OP_423J2_125_3477_n2235), .B(
        DP_OP_423J2_125_3477_n2279), .CI(DP_OP_423J2_125_3477_n2059), .CO(
        DP_OP_423J2_125_3477_n1668), .S(DP_OP_423J2_125_3477_n1669) );
  FADDX1_HVT DP_OP_423J2_125_3477_U991 ( .A(DP_OP_423J2_125_3477_n2763), .B(
        DP_OP_423J2_125_3477_n2631), .CI(DP_OP_423J2_125_3477_n2675), .CO(
        DP_OP_423J2_125_3477_n1666), .S(DP_OP_423J2_125_3477_n1667) );
  FADDX1_HVT DP_OP_423J2_125_3477_U990 ( .A(DP_OP_423J2_125_3477_n2015), .B(
        DP_OP_423J2_125_3477_n2851), .CI(DP_OP_423J2_125_3477_n2719), .CO(
        DP_OP_423J2_125_3477_n1664), .S(DP_OP_423J2_125_3477_n1665) );
  FADDX1_HVT DP_OP_423J2_125_3477_U989 ( .A(DP_OP_423J2_125_3477_n2543), .B(
        DP_OP_423J2_125_3477_n2939), .CI(DP_OP_423J2_125_3477_n2191), .CO(
        DP_OP_423J2_125_3477_n1662), .S(DP_OP_423J2_125_3477_n1663) );
  FADDX1_HVT DP_OP_423J2_125_3477_U988 ( .A(DP_OP_423J2_125_3477_n1971), .B(
        DP_OP_423J2_125_3477_n1679), .CI(DP_OP_423J2_125_3477_n1948), .CO(
        DP_OP_423J2_125_3477_n1660), .S(DP_OP_423J2_125_3477_n1661) );
  FADDX1_HVT DP_OP_423J2_125_3477_U987 ( .A(DP_OP_423J2_125_3477_n1978), .B(
        DP_OP_423J2_125_3477_n1941), .CI(DP_OP_423J2_125_3477_n1934), .CO(
        DP_OP_423J2_125_3477_n1658), .S(DP_OP_423J2_125_3477_n1659) );
  FADDX1_HVT DP_OP_423J2_125_3477_U986 ( .A(DP_OP_423J2_125_3477_n1992), .B(
        DP_OP_423J2_125_3477_n1985), .CI(DP_OP_423J2_125_3477_n2022), .CO(
        DP_OP_423J2_125_3477_n1656), .S(DP_OP_423J2_125_3477_n1657) );
  FADDX1_HVT DP_OP_423J2_125_3477_U985 ( .A(DP_OP_423J2_125_3477_n2036), .B(
        DP_OP_423J2_125_3477_n2029), .CI(DP_OP_423J2_125_3477_n2066), .CO(
        DP_OP_423J2_125_3477_n1654), .S(DP_OP_423J2_125_3477_n1655) );
  FADDX1_HVT DP_OP_423J2_125_3477_U984 ( .A(DP_OP_423J2_125_3477_n3002), .B(
        DP_OP_423J2_125_3477_n2073), .CI(DP_OP_423J2_125_3477_n2080), .CO(
        DP_OP_423J2_125_3477_n1652), .S(DP_OP_423J2_125_3477_n1653) );
  FADDX1_HVT DP_OP_423J2_125_3477_U983 ( .A(DP_OP_423J2_125_3477_n2513), .B(
        DP_OP_423J2_125_3477_n2995), .CI(DP_OP_423J2_125_3477_n2988), .CO(
        DP_OP_423J2_125_3477_n1650), .S(DP_OP_423J2_125_3477_n1651) );
  FADDX1_HVT DP_OP_423J2_125_3477_U982 ( .A(DP_OP_423J2_125_3477_n2476), .B(
        DP_OP_423J2_125_3477_n2110), .CI(DP_OP_423J2_125_3477_n2960), .CO(
        DP_OP_423J2_125_3477_n1648), .S(DP_OP_423J2_125_3477_n1649) );
  FADDX1_HVT DP_OP_423J2_125_3477_U981 ( .A(DP_OP_423J2_125_3477_n2506), .B(
        DP_OP_423J2_125_3477_n2117), .CI(DP_OP_423J2_125_3477_n2953), .CO(
        DP_OP_423J2_125_3477_n1646), .S(DP_OP_423J2_125_3477_n1647) );
  FADDX1_HVT DP_OP_423J2_125_3477_U980 ( .A(DP_OP_423J2_125_3477_n2946), .B(
        DP_OP_423J2_125_3477_n2124), .CI(DP_OP_423J2_125_3477_n2154), .CO(
        DP_OP_423J2_125_3477_n1644), .S(DP_OP_423J2_125_3477_n1645) );
  FADDX1_HVT DP_OP_423J2_125_3477_U979 ( .A(DP_OP_423J2_125_3477_n2469), .B(
        DP_OP_423J2_125_3477_n2161), .CI(DP_OP_423J2_125_3477_n2168), .CO(
        DP_OP_423J2_125_3477_n1642), .S(DP_OP_423J2_125_3477_n1643) );
  FADDX1_HVT DP_OP_423J2_125_3477_U978 ( .A(DP_OP_423J2_125_3477_n2550), .B(
        DP_OP_423J2_125_3477_n2198), .CI(DP_OP_423J2_125_3477_n2205), .CO(
        DP_OP_423J2_125_3477_n1640), .S(DP_OP_423J2_125_3477_n1641) );
  FADDX1_HVT DP_OP_423J2_125_3477_U977 ( .A(DP_OP_423J2_125_3477_n2557), .B(
        DP_OP_423J2_125_3477_n2212), .CI(DP_OP_423J2_125_3477_n2242), .CO(
        DP_OP_423J2_125_3477_n1638), .S(DP_OP_423J2_125_3477_n1639) );
  FADDX1_HVT DP_OP_423J2_125_3477_U976 ( .A(DP_OP_423J2_125_3477_n2564), .B(
        DP_OP_423J2_125_3477_n2916), .CI(DP_OP_423J2_125_3477_n2249), .CO(
        DP_OP_423J2_125_3477_n1636), .S(DP_OP_423J2_125_3477_n1637) );
  FADDX1_HVT DP_OP_423J2_125_3477_U975 ( .A(DP_OP_423J2_125_3477_n2594), .B(
        DP_OP_423J2_125_3477_n2256), .CI(DP_OP_423J2_125_3477_n2909), .CO(
        DP_OP_423J2_125_3477_n1634), .S(DP_OP_423J2_125_3477_n1635) );
  FADDX1_HVT DP_OP_423J2_125_3477_U974 ( .A(DP_OP_423J2_125_3477_n2520), .B(
        DP_OP_423J2_125_3477_n2902), .CI(DP_OP_423J2_125_3477_n2872), .CO(
        DP_OP_423J2_125_3477_n1632), .S(DP_OP_423J2_125_3477_n1633) );
  FADDX1_HVT DP_OP_423J2_125_3477_U973 ( .A(DP_OP_423J2_125_3477_n2432), .B(
        DP_OP_423J2_125_3477_n2865), .CI(DP_OP_423J2_125_3477_n2286), .CO(
        DP_OP_423J2_125_3477_n1630), .S(DP_OP_423J2_125_3477_n1631) );
  FADDX1_HVT DP_OP_423J2_125_3477_U972 ( .A(DP_OP_423J2_125_3477_n2858), .B(
        DP_OP_423J2_125_3477_n2293), .CI(DP_OP_423J2_125_3477_n2828), .CO(
        DP_OP_423J2_125_3477_n1628), .S(DP_OP_423J2_125_3477_n1629) );
  FADDX1_HVT DP_OP_423J2_125_3477_U971 ( .A(DP_OP_423J2_125_3477_n2821), .B(
        DP_OP_423J2_125_3477_n2814), .CI(DP_OP_423J2_125_3477_n2300), .CO(
        DP_OP_423J2_125_3477_n1626), .S(DP_OP_423J2_125_3477_n1627) );
  FADDX1_HVT DP_OP_423J2_125_3477_U970 ( .A(DP_OP_423J2_125_3477_n2425), .B(
        DP_OP_423J2_125_3477_n2330), .CI(DP_OP_423J2_125_3477_n2784), .CO(
        DP_OP_423J2_125_3477_n1624), .S(DP_OP_423J2_125_3477_n1625) );
  FADDX1_HVT DP_OP_423J2_125_3477_U969 ( .A(DP_OP_423J2_125_3477_n2418), .B(
        DP_OP_423J2_125_3477_n2777), .CI(DP_OP_423J2_125_3477_n2770), .CO(
        DP_OP_423J2_125_3477_n1622), .S(DP_OP_423J2_125_3477_n1623) );
  FADDX1_HVT DP_OP_423J2_125_3477_U968 ( .A(DP_OP_423J2_125_3477_n2374), .B(
        DP_OP_423J2_125_3477_n2740), .CI(DP_OP_423J2_125_3477_n2733), .CO(
        DP_OP_423J2_125_3477_n1620), .S(DP_OP_423J2_125_3477_n1621) );
  FADDX1_HVT DP_OP_423J2_125_3477_U967 ( .A(DP_OP_423J2_125_3477_n2337), .B(
        DP_OP_423J2_125_3477_n2726), .CI(DP_OP_423J2_125_3477_n2696), .CO(
        DP_OP_423J2_125_3477_n1618), .S(DP_OP_423J2_125_3477_n1619) );
  FADDX1_HVT DP_OP_423J2_125_3477_U966 ( .A(DP_OP_423J2_125_3477_n2608), .B(
        DP_OP_423J2_125_3477_n2689), .CI(DP_OP_423J2_125_3477_n2344), .CO(
        DP_OP_423J2_125_3477_n1616), .S(DP_OP_423J2_125_3477_n1617) );
  FADDX1_HVT DP_OP_423J2_125_3477_U965 ( .A(DP_OP_423J2_125_3477_n2462), .B(
        DP_OP_423J2_125_3477_n2381), .CI(DP_OP_423J2_125_3477_n2682), .CO(
        DP_OP_423J2_125_3477_n1614), .S(DP_OP_423J2_125_3477_n1615) );
  FADDX1_HVT DP_OP_423J2_125_3477_U964 ( .A(DP_OP_423J2_125_3477_n2652), .B(
        DP_OP_423J2_125_3477_n2388), .CI(DP_OP_423J2_125_3477_n2601), .CO(
        DP_OP_423J2_125_3477_n1612), .S(DP_OP_423J2_125_3477_n1613) );
  FADDX1_HVT DP_OP_423J2_125_3477_U963 ( .A(DP_OP_423J2_125_3477_n2645), .B(
        DP_OP_423J2_125_3477_n2638), .CI(DP_OP_423J2_125_3477_n1784), .CO(
        DP_OP_423J2_125_3477_n1610), .S(DP_OP_423J2_125_3477_n1611) );
  FADDX1_HVT DP_OP_423J2_125_3477_U962 ( .A(DP_OP_423J2_125_3477_n1760), .B(
        DP_OP_423J2_125_3477_n1782), .CI(DP_OP_423J2_125_3477_n1736), .CO(
        DP_OP_423J2_125_3477_n1608), .S(DP_OP_423J2_125_3477_n1609) );
  FADDX1_HVT DP_OP_423J2_125_3477_U961 ( .A(DP_OP_423J2_125_3477_n1758), .B(
        DP_OP_423J2_125_3477_n1780), .CI(DP_OP_423J2_125_3477_n1778), .CO(
        DP_OP_423J2_125_3477_n1606), .S(DP_OP_423J2_125_3477_n1607) );
  FADDX1_HVT DP_OP_423J2_125_3477_U960 ( .A(DP_OP_423J2_125_3477_n1752), .B(
        DP_OP_423J2_125_3477_n1776), .CI(DP_OP_423J2_125_3477_n1774), .CO(
        DP_OP_423J2_125_3477_n1604), .S(DP_OP_423J2_125_3477_n1605) );
  FADDX1_HVT DP_OP_423J2_125_3477_U959 ( .A(DP_OP_423J2_125_3477_n1748), .B(
        DP_OP_423J2_125_3477_n1738), .CI(DP_OP_423J2_125_3477_n1740), .CO(
        DP_OP_423J2_125_3477_n1602), .S(DP_OP_423J2_125_3477_n1603) );
  FADDX1_HVT DP_OP_423J2_125_3477_U958 ( .A(DP_OP_423J2_125_3477_n1746), .B(
        DP_OP_423J2_125_3477_n1772), .CI(DP_OP_423J2_125_3477_n1742), .CO(
        DP_OP_423J2_125_3477_n1600), .S(DP_OP_423J2_125_3477_n1601) );
  FADDX1_HVT DP_OP_423J2_125_3477_U957 ( .A(DP_OP_423J2_125_3477_n1744), .B(
        DP_OP_423J2_125_3477_n1770), .CI(DP_OP_423J2_125_3477_n1768), .CO(
        DP_OP_423J2_125_3477_n1598), .S(DP_OP_423J2_125_3477_n1599) );
  FADDX1_HVT DP_OP_423J2_125_3477_U956 ( .A(DP_OP_423J2_125_3477_n1756), .B(
        DP_OP_423J2_125_3477_n1766), .CI(DP_OP_423J2_125_3477_n1750), .CO(
        DP_OP_423J2_125_3477_n1596), .S(DP_OP_423J2_125_3477_n1597) );
  FADDX1_HVT DP_OP_423J2_125_3477_U955 ( .A(DP_OP_423J2_125_3477_n1764), .B(
        DP_OP_423J2_125_3477_n1762), .CI(DP_OP_423J2_125_3477_n1754), .CO(
        DP_OP_423J2_125_3477_n1594), .S(DP_OP_423J2_125_3477_n1595) );
  FADDX1_HVT DP_OP_423J2_125_3477_U954 ( .A(DP_OP_423J2_125_3477_n1673), .B(
        DP_OP_423J2_125_3477_n1675), .CI(DP_OP_423J2_125_3477_n1661), .CO(
        DP_OP_423J2_125_3477_n1592), .S(DP_OP_423J2_125_3477_n1593) );
  FADDX1_HVT DP_OP_423J2_125_3477_U953 ( .A(DP_OP_423J2_125_3477_n1667), .B(
        DP_OP_423J2_125_3477_n1669), .CI(DP_OP_423J2_125_3477_n1734), .CO(
        DP_OP_423J2_125_3477_n1590), .S(DP_OP_423J2_125_3477_n1591) );
  FADDX1_HVT DP_OP_423J2_125_3477_U952 ( .A(DP_OP_423J2_125_3477_n1663), .B(
        DP_OP_423J2_125_3477_n1665), .CI(DP_OP_423J2_125_3477_n1671), .CO(
        DP_OP_423J2_125_3477_n1588), .S(DP_OP_423J2_125_3477_n1589) );
  FADDX1_HVT DP_OP_423J2_125_3477_U951 ( .A(DP_OP_423J2_125_3477_n1677), .B(
        DP_OP_423J2_125_3477_n1627), .CI(DP_OP_423J2_125_3477_n1625), .CO(
        DP_OP_423J2_125_3477_n1586), .S(DP_OP_423J2_125_3477_n1587) );
  FADDX1_HVT DP_OP_423J2_125_3477_U950 ( .A(DP_OP_423J2_125_3477_n1629), .B(
        DP_OP_423J2_125_3477_n1645), .CI(DP_OP_423J2_125_3477_n1653), .CO(
        DP_OP_423J2_125_3477_n1584), .S(DP_OP_423J2_125_3477_n1585) );
  FADDX1_HVT DP_OP_423J2_125_3477_U949 ( .A(DP_OP_423J2_125_3477_n1621), .B(
        DP_OP_423J2_125_3477_n1641), .CI(DP_OP_423J2_125_3477_n1639), .CO(
        DP_OP_423J2_125_3477_n1582), .S(DP_OP_423J2_125_3477_n1583) );
  FADDX1_HVT DP_OP_423J2_125_3477_U948 ( .A(DP_OP_423J2_125_3477_n1619), .B(
        DP_OP_423J2_125_3477_n1655), .CI(DP_OP_423J2_125_3477_n1643), .CO(
        DP_OP_423J2_125_3477_n1580), .S(DP_OP_423J2_125_3477_n1581) );
  FADDX1_HVT DP_OP_423J2_125_3477_U947 ( .A(DP_OP_423J2_125_3477_n1617), .B(
        DP_OP_423J2_125_3477_n1649), .CI(DP_OP_423J2_125_3477_n1651), .CO(
        DP_OP_423J2_125_3477_n1578), .S(DP_OP_423J2_125_3477_n1579) );
  FADDX1_HVT DP_OP_423J2_125_3477_U946 ( .A(DP_OP_423J2_125_3477_n1615), .B(
        DP_OP_423J2_125_3477_n1647), .CI(DP_OP_423J2_125_3477_n1659), .CO(
        DP_OP_423J2_125_3477_n1576), .S(DP_OP_423J2_125_3477_n1577) );
  FADDX1_HVT DP_OP_423J2_125_3477_U945 ( .A(DP_OP_423J2_125_3477_n1637), .B(
        DP_OP_423J2_125_3477_n1657), .CI(DP_OP_423J2_125_3477_n1613), .CO(
        DP_OP_423J2_125_3477_n1574), .S(DP_OP_423J2_125_3477_n1575) );
  FADDX1_HVT DP_OP_423J2_125_3477_U944 ( .A(DP_OP_423J2_125_3477_n1623), .B(
        DP_OP_423J2_125_3477_n1633), .CI(DP_OP_423J2_125_3477_n1635), .CO(
        DP_OP_423J2_125_3477_n1572), .S(DP_OP_423J2_125_3477_n1573) );
  FADDX1_HVT DP_OP_423J2_125_3477_U943 ( .A(DP_OP_423J2_125_3477_n1631), .B(
        DP_OP_423J2_125_3477_n1611), .CI(DP_OP_423J2_125_3477_n1732), .CO(
        DP_OP_423J2_125_3477_n1570), .S(DP_OP_423J2_125_3477_n1571) );
  FADDX1_HVT DP_OP_423J2_125_3477_U942 ( .A(DP_OP_423J2_125_3477_n1730), .B(
        DP_OP_423J2_125_3477_n1728), .CI(DP_OP_423J2_125_3477_n1726), .CO(
        DP_OP_423J2_125_3477_n1568), .S(DP_OP_423J2_125_3477_n1569) );
  FADDX1_HVT DP_OP_423J2_125_3477_U941 ( .A(DP_OP_423J2_125_3477_n1724), .B(
        DP_OP_423J2_125_3477_n1722), .CI(DP_OP_423J2_125_3477_n1710), .CO(
        DP_OP_423J2_125_3477_n1566), .S(DP_OP_423J2_125_3477_n1567) );
  FADDX1_HVT DP_OP_423J2_125_3477_U940 ( .A(DP_OP_423J2_125_3477_n1708), .B(
        DP_OP_423J2_125_3477_n1609), .CI(DP_OP_423J2_125_3477_n1706), .CO(
        DP_OP_423J2_125_3477_n1564), .S(DP_OP_423J2_125_3477_n1565) );
  FADDX1_HVT DP_OP_423J2_125_3477_U939 ( .A(DP_OP_423J2_125_3477_n1720), .B(
        DP_OP_423J2_125_3477_n1599), .CI(DP_OP_423J2_125_3477_n1607), .CO(
        DP_OP_423J2_125_3477_n1562), .S(DP_OP_423J2_125_3477_n1563) );
  FADDX1_HVT DP_OP_423J2_125_3477_U938 ( .A(DP_OP_423J2_125_3477_n1718), .B(
        DP_OP_423J2_125_3477_n1597), .CI(DP_OP_423J2_125_3477_n1601), .CO(
        DP_OP_423J2_125_3477_n1560), .S(DP_OP_423J2_125_3477_n1561) );
  FADDX1_HVT DP_OP_423J2_125_3477_U937 ( .A(DP_OP_423J2_125_3477_n1714), .B(
        DP_OP_423J2_125_3477_n1605), .CI(DP_OP_423J2_125_3477_n1603), .CO(
        DP_OP_423J2_125_3477_n1558), .S(DP_OP_423J2_125_3477_n1559) );
  FADDX1_HVT DP_OP_423J2_125_3477_U936 ( .A(DP_OP_423J2_125_3477_n1712), .B(
        DP_OP_423J2_125_3477_n1716), .CI(DP_OP_423J2_125_3477_n1595), .CO(
        DP_OP_423J2_125_3477_n1556), .S(DP_OP_423J2_125_3477_n1557) );
  FADDX1_HVT DP_OP_423J2_125_3477_U935 ( .A(DP_OP_423J2_125_3477_n1591), .B(
        DP_OP_423J2_125_3477_n1593), .CI(DP_OP_423J2_125_3477_n1587), .CO(
        DP_OP_423J2_125_3477_n1554), .S(DP_OP_423J2_125_3477_n1555) );
  FADDX1_HVT DP_OP_423J2_125_3477_U934 ( .A(DP_OP_423J2_125_3477_n1589), .B(
        DP_OP_423J2_125_3477_n1575), .CI(DP_OP_423J2_125_3477_n1577), .CO(
        DP_OP_423J2_125_3477_n1552), .S(DP_OP_423J2_125_3477_n1553) );
  FADDX1_HVT DP_OP_423J2_125_3477_U933 ( .A(DP_OP_423J2_125_3477_n1583), .B(
        DP_OP_423J2_125_3477_n1581), .CI(DP_OP_423J2_125_3477_n1704), .CO(
        DP_OP_423J2_125_3477_n1550), .S(DP_OP_423J2_125_3477_n1551) );
  FADDX1_HVT DP_OP_423J2_125_3477_U932 ( .A(DP_OP_423J2_125_3477_n1579), .B(
        DP_OP_423J2_125_3477_n1573), .CI(DP_OP_423J2_125_3477_n1585), .CO(
        DP_OP_423J2_125_3477_n1548), .S(DP_OP_423J2_125_3477_n1549) );
  FADDX1_HVT DP_OP_423J2_125_3477_U931 ( .A(DP_OP_423J2_125_3477_n1571), .B(
        DP_OP_423J2_125_3477_n1702), .CI(DP_OP_423J2_125_3477_n1698), .CO(
        DP_OP_423J2_125_3477_n1546), .S(DP_OP_423J2_125_3477_n1547) );
  FADDX1_HVT DP_OP_423J2_125_3477_U930 ( .A(DP_OP_423J2_125_3477_n1700), .B(
        DP_OP_423J2_125_3477_n1569), .CI(DP_OP_423J2_125_3477_n1696), .CO(
        DP_OP_423J2_125_3477_n1544), .S(DP_OP_423J2_125_3477_n1545) );
  FADDX1_HVT DP_OP_423J2_125_3477_U929 ( .A(DP_OP_423J2_125_3477_n1567), .B(
        DP_OP_423J2_125_3477_n1557), .CI(DP_OP_423J2_125_3477_n1559), .CO(
        DP_OP_423J2_125_3477_n1542), .S(DP_OP_423J2_125_3477_n1543) );
  FADDX1_HVT DP_OP_423J2_125_3477_U928 ( .A(DP_OP_423J2_125_3477_n1694), .B(
        DP_OP_423J2_125_3477_n1561), .CI(DP_OP_423J2_125_3477_n1692), .CO(
        DP_OP_423J2_125_3477_n1540), .S(DP_OP_423J2_125_3477_n1541) );
  FADDX1_HVT DP_OP_423J2_125_3477_U927 ( .A(DP_OP_423J2_125_3477_n1565), .B(
        DP_OP_423J2_125_3477_n1563), .CI(DP_OP_423J2_125_3477_n1555), .CO(
        DP_OP_423J2_125_3477_n1538), .S(DP_OP_423J2_125_3477_n1539) );
  FADDX1_HVT DP_OP_423J2_125_3477_U926 ( .A(DP_OP_423J2_125_3477_n1690), .B(
        DP_OP_423J2_125_3477_n1553), .CI(DP_OP_423J2_125_3477_n1549), .CO(
        DP_OP_423J2_125_3477_n1536), .S(DP_OP_423J2_125_3477_n1537) );
  FADDX1_HVT DP_OP_423J2_125_3477_U925 ( .A(DP_OP_423J2_125_3477_n1551), .B(
        DP_OP_423J2_125_3477_n1688), .CI(DP_OP_423J2_125_3477_n1547), .CO(
        DP_OP_423J2_125_3477_n1534), .S(DP_OP_423J2_125_3477_n1535) );
  FADDX1_HVT DP_OP_423J2_125_3477_U924 ( .A(DP_OP_423J2_125_3477_n1686), .B(
        DP_OP_423J2_125_3477_n1545), .CI(DP_OP_423J2_125_3477_n1684), .CO(
        DP_OP_423J2_125_3477_n1532), .S(DP_OP_423J2_125_3477_n1533) );
  FADDX1_HVT DP_OP_423J2_125_3477_U923 ( .A(DP_OP_423J2_125_3477_n1543), .B(
        DP_OP_423J2_125_3477_n1541), .CI(DP_OP_423J2_125_3477_n1539), .CO(
        DP_OP_423J2_125_3477_n1530), .S(DP_OP_423J2_125_3477_n1531) );
  FADDX1_HVT DP_OP_423J2_125_3477_U922 ( .A(DP_OP_423J2_125_3477_n1537), .B(
        DP_OP_423J2_125_3477_n1682), .CI(DP_OP_423J2_125_3477_n1535), .CO(
        DP_OP_423J2_125_3477_n1528), .S(DP_OP_423J2_125_3477_n1529) );
  FADDX1_HVT DP_OP_423J2_125_3477_U921 ( .A(DP_OP_423J2_125_3477_n1680), .B(
        DP_OP_423J2_125_3477_n1533), .CI(DP_OP_423J2_125_3477_n1531), .CO(
        DP_OP_423J2_125_3477_n1526), .S(DP_OP_423J2_125_3477_n1527) );
  FADDX1_HVT DP_OP_423J2_125_3477_U920 ( .A(DP_OP_423J2_125_3477_n1678), .B(
        DP_OP_423J2_125_3477_n1926), .CI(DP_OP_423J2_125_3477_n1882), .CO(
        DP_OP_423J2_125_3477_n1524), .S(DP_OP_423J2_125_3477_n1525) );
  FADDX1_HVT DP_OP_423J2_125_3477_U919 ( .A(DP_OP_423J2_125_3477_n2981), .B(
        DP_OP_423J2_125_3477_n2498), .CI(DP_OP_423J2_125_3477_n2366), .CO(
        DP_OP_423J2_125_3477_n1522), .S(DP_OP_423J2_125_3477_n1523) );
  FADDX1_HVT DP_OP_423J2_125_3477_U918 ( .A(DP_OP_423J2_125_3477_n2894), .B(
        DP_OP_423J2_125_3477_n2630), .CI(DP_OP_423J2_125_3477_n2278), .CO(
        DP_OP_423J2_125_3477_n1520), .S(DP_OP_423J2_125_3477_n1521) );
  FADDX1_HVT DP_OP_423J2_125_3477_U917 ( .A(DP_OP_423J2_125_3477_n2058), .B(
        DP_OP_423J2_125_3477_n2586), .CI(DP_OP_423J2_125_3477_n2806), .CO(
        DP_OP_423J2_125_3477_n1518), .S(DP_OP_423J2_125_3477_n1519) );
  FADDX1_HVT DP_OP_423J2_125_3477_U916 ( .A(DP_OP_423J2_125_3477_n2146), .B(
        DP_OP_423J2_125_3477_n2322), .CI(DP_OP_423J2_125_3477_n2410), .CO(
        DP_OP_423J2_125_3477_n1516), .S(DP_OP_423J2_125_3477_n1517) );
  FADDX1_HVT DP_OP_423J2_125_3477_U915 ( .A(DP_OP_423J2_125_3477_n2762), .B(
        DP_OP_423J2_125_3477_n2234), .CI(DP_OP_423J2_125_3477_n2850), .CO(
        DP_OP_423J2_125_3477_n1514), .S(DP_OP_423J2_125_3477_n1515) );
  FADDX1_HVT DP_OP_423J2_125_3477_U914 ( .A(DP_OP_423J2_125_3477_n2102), .B(
        DP_OP_423J2_125_3477_n2454), .CI(DP_OP_423J2_125_3477_n2542), .CO(
        DP_OP_423J2_125_3477_n1512), .S(DP_OP_423J2_125_3477_n1513) );
  FADDX1_HVT DP_OP_423J2_125_3477_U913 ( .A(DP_OP_423J2_125_3477_n2938), .B(
        DP_OP_423J2_125_3477_n2674), .CI(DP_OP_423J2_125_3477_n2718), .CO(
        DP_OP_423J2_125_3477_n1510), .S(DP_OP_423J2_125_3477_n1511) );
  FADDX1_HVT DP_OP_423J2_125_3477_U912 ( .A(DP_OP_423J2_125_3477_n2014), .B(
        DP_OP_423J2_125_3477_n2190), .CI(DP_OP_423J2_125_3477_n1970), .CO(
        DP_OP_423J2_125_3477_n1508), .S(DP_OP_423J2_125_3477_n1509) );
  FADDX1_HVT DP_OP_423J2_125_3477_U911 ( .A(DP_OP_423J2_125_3477_n2505), .B(
        DP_OP_423J2_125_3477_n1940), .CI(DP_OP_423J2_125_3477_n1933), .CO(
        DP_OP_423J2_125_3477_n1506), .S(DP_OP_423J2_125_3477_n1507) );
  FADDX1_HVT DP_OP_423J2_125_3477_U910 ( .A(DP_OP_423J2_125_3477_n3001), .B(
        DP_OP_423J2_125_3477_n1947), .CI(DP_OP_423J2_125_3477_n1977), .CO(
        DP_OP_423J2_125_3477_n1504), .S(DP_OP_423J2_125_3477_n1505) );
  FADDX1_HVT DP_OP_423J2_125_3477_U909 ( .A(DP_OP_423J2_125_3477_n2387), .B(
        DP_OP_423J2_125_3477_n2994), .CI(DP_OP_423J2_125_3477_n1984), .CO(
        DP_OP_423J2_125_3477_n1502), .S(DP_OP_423J2_125_3477_n1503) );
  FADDX1_HVT DP_OP_423J2_125_3477_U908 ( .A(DP_OP_423J2_125_3477_n2380), .B(
        DP_OP_423J2_125_3477_n2987), .CI(DP_OP_423J2_125_3477_n1991), .CO(
        DP_OP_423J2_125_3477_n1500), .S(DP_OP_423J2_125_3477_n1501) );
  FADDX1_HVT DP_OP_423J2_125_3477_U907 ( .A(DP_OP_423J2_125_3477_n2959), .B(
        DP_OP_423J2_125_3477_n2021), .CI(DP_OP_423J2_125_3477_n2028), .CO(
        DP_OP_423J2_125_3477_n1498), .S(DP_OP_423J2_125_3477_n1499) );
  FADDX1_HVT DP_OP_423J2_125_3477_U906 ( .A(DP_OP_423J2_125_3477_n2417), .B(
        DP_OP_423J2_125_3477_n2952), .CI(DP_OP_423J2_125_3477_n2945), .CO(
        DP_OP_423J2_125_3477_n1496), .S(DP_OP_423J2_125_3477_n1497) );
  FADDX1_HVT DP_OP_423J2_125_3477_U905 ( .A(DP_OP_423J2_125_3477_n2343), .B(
        DP_OP_423J2_125_3477_n2915), .CI(DP_OP_423J2_125_3477_n2908), .CO(
        DP_OP_423J2_125_3477_n1494), .S(DP_OP_423J2_125_3477_n1495) );
  FADDX1_HVT DP_OP_423J2_125_3477_U904 ( .A(DP_OP_423J2_125_3477_n2336), .B(
        DP_OP_423J2_125_3477_n2901), .CI(DP_OP_423J2_125_3477_n2035), .CO(
        DP_OP_423J2_125_3477_n1492), .S(DP_OP_423J2_125_3477_n1493) );
  FADDX1_HVT DP_OP_423J2_125_3477_U903 ( .A(DP_OP_423J2_125_3477_n2329), .B(
        DP_OP_423J2_125_3477_n2871), .CI(DP_OP_423J2_125_3477_n2864), .CO(
        DP_OP_423J2_125_3477_n1490), .S(DP_OP_423J2_125_3477_n1491) );
  FADDX1_HVT DP_OP_423J2_125_3477_U902 ( .A(DP_OP_423J2_125_3477_n2299), .B(
        DP_OP_423J2_125_3477_n2857), .CI(DP_OP_423J2_125_3477_n2065), .CO(
        DP_OP_423J2_125_3477_n1488), .S(DP_OP_423J2_125_3477_n1489) );
  FADDX1_HVT DP_OP_423J2_125_3477_U901 ( .A(DP_OP_423J2_125_3477_n2292), .B(
        DP_OP_423J2_125_3477_n2072), .CI(DP_OP_423J2_125_3477_n2079), .CO(
        DP_OP_423J2_125_3477_n1486), .S(DP_OP_423J2_125_3477_n1487) );
  FADDX1_HVT DP_OP_423J2_125_3477_U900 ( .A(DP_OP_423J2_125_3477_n2373), .B(
        DP_OP_423J2_125_3477_n2109), .CI(DP_OP_423J2_125_3477_n2827), .CO(
        DP_OP_423J2_125_3477_n1484), .S(DP_OP_423J2_125_3477_n1485) );
  FADDX1_HVT DP_OP_423J2_125_3477_U899 ( .A(DP_OP_423J2_125_3477_n2424), .B(
        DP_OP_423J2_125_3477_n2820), .CI(DP_OP_423J2_125_3477_n2813), .CO(
        DP_OP_423J2_125_3477_n1482), .S(DP_OP_423J2_125_3477_n1483) );
  FADDX1_HVT DP_OP_423J2_125_3477_U898 ( .A(DP_OP_423J2_125_3477_n2783), .B(
        DP_OP_423J2_125_3477_n2116), .CI(DP_OP_423J2_125_3477_n2123), .CO(
        DP_OP_423J2_125_3477_n1480), .S(DP_OP_423J2_125_3477_n1481) );
  FADDX1_HVT DP_OP_423J2_125_3477_U897 ( .A(DP_OP_423J2_125_3477_n2556), .B(
        DP_OP_423J2_125_3477_n2153), .CI(DP_OP_423J2_125_3477_n2160), .CO(
        DP_OP_423J2_125_3477_n1478), .S(DP_OP_423J2_125_3477_n1479) );
  FADDX1_HVT DP_OP_423J2_125_3477_U896 ( .A(DP_OP_423J2_125_3477_n2776), .B(
        DP_OP_423J2_125_3477_n2167), .CI(DP_OP_423J2_125_3477_n2197), .CO(
        DP_OP_423J2_125_3477_n1476), .S(DP_OP_423J2_125_3477_n1477) );
  FADDX1_HVT DP_OP_423J2_125_3477_U895 ( .A(DP_OP_423J2_125_3477_n2769), .B(
        DP_OP_423J2_125_3477_n2204), .CI(DP_OP_423J2_125_3477_n2211), .CO(
        DP_OP_423J2_125_3477_n1474), .S(DP_OP_423J2_125_3477_n1475) );
  FADDX1_HVT DP_OP_423J2_125_3477_U894 ( .A(DP_OP_423J2_125_3477_n2739), .B(
        DP_OP_423J2_125_3477_n2241), .CI(DP_OP_423J2_125_3477_n2248), .CO(
        DP_OP_423J2_125_3477_n1472), .S(DP_OP_423J2_125_3477_n1473) );
  FADDX1_HVT DP_OP_423J2_125_3477_U893 ( .A(DP_OP_423J2_125_3477_n2732), .B(
        DP_OP_423J2_125_3477_n2255), .CI(DP_OP_423J2_125_3477_n2285), .CO(
        DP_OP_423J2_125_3477_n1470), .S(DP_OP_423J2_125_3477_n1471) );
  FADDX1_HVT DP_OP_423J2_125_3477_U892 ( .A(DP_OP_423J2_125_3477_n2725), .B(
        DP_OP_423J2_125_3477_n2431), .CI(DP_OP_423J2_125_3477_n2461), .CO(
        DP_OP_423J2_125_3477_n1468), .S(DP_OP_423J2_125_3477_n1469) );
  FADDX1_HVT DP_OP_423J2_125_3477_U891 ( .A(DP_OP_423J2_125_3477_n2695), .B(
        DP_OP_423J2_125_3477_n2468), .CI(DP_OP_423J2_125_3477_n2688), .CO(
        DP_OP_423J2_125_3477_n1466), .S(DP_OP_423J2_125_3477_n1467) );
  FADDX1_HVT DP_OP_423J2_125_3477_U890 ( .A(DP_OP_423J2_125_3477_n2593), .B(
        DP_OP_423J2_125_3477_n2475), .CI(DP_OP_423J2_125_3477_n2512), .CO(
        DP_OP_423J2_125_3477_n1464), .S(DP_OP_423J2_125_3477_n1465) );
  FADDX1_HVT DP_OP_423J2_125_3477_U889 ( .A(DP_OP_423J2_125_3477_n2563), .B(
        DP_OP_423J2_125_3477_n2519), .CI(DP_OP_423J2_125_3477_n2681), .CO(
        DP_OP_423J2_125_3477_n1462), .S(DP_OP_423J2_125_3477_n1463) );
  FADDX1_HVT DP_OP_423J2_125_3477_U888 ( .A(DP_OP_423J2_125_3477_n2637), .B(
        DP_OP_423J2_125_3477_n2549), .CI(DP_OP_423J2_125_3477_n2651), .CO(
        DP_OP_423J2_125_3477_n1460), .S(DP_OP_423J2_125_3477_n1461) );
  FADDX1_HVT DP_OP_423J2_125_3477_U887 ( .A(DP_OP_423J2_125_3477_n2600), .B(
        DP_OP_423J2_125_3477_n2607), .CI(DP_OP_423J2_125_3477_n2644), .CO(
        DP_OP_423J2_125_3477_n1458), .S(DP_OP_423J2_125_3477_n1459) );
  FADDX1_HVT DP_OP_423J2_125_3477_U886 ( .A(DP_OP_423J2_125_3477_n1666), .B(
        DP_OP_423J2_125_3477_n1662), .CI(DP_OP_423J2_125_3477_n1660), .CO(
        DP_OP_423J2_125_3477_n1456), .S(DP_OP_423J2_125_3477_n1457) );
  FADDX1_HVT DP_OP_423J2_125_3477_U885 ( .A(DP_OP_423J2_125_3477_n1664), .B(
        DP_OP_423J2_125_3477_n1668), .CI(DP_OP_423J2_125_3477_n1670), .CO(
        DP_OP_423J2_125_3477_n1454), .S(DP_OP_423J2_125_3477_n1455) );
  FADDX1_HVT DP_OP_423J2_125_3477_U884 ( .A(DP_OP_423J2_125_3477_n1672), .B(
        DP_OP_423J2_125_3477_n1674), .CI(DP_OP_423J2_125_3477_n1676), .CO(
        DP_OP_423J2_125_3477_n1452), .S(DP_OP_423J2_125_3477_n1453) );
  FADDX1_HVT DP_OP_423J2_125_3477_U883 ( .A(DP_OP_423J2_125_3477_n1636), .B(
        DP_OP_423J2_125_3477_n1658), .CI(DP_OP_423J2_125_3477_n1656), .CO(
        DP_OP_423J2_125_3477_n1450), .S(DP_OP_423J2_125_3477_n1451) );
  FADDX1_HVT DP_OP_423J2_125_3477_U882 ( .A(DP_OP_423J2_125_3477_n1632), .B(
        DP_OP_423J2_125_3477_n1654), .CI(DP_OP_423J2_125_3477_n1652), .CO(
        DP_OP_423J2_125_3477_n1448), .S(DP_OP_423J2_125_3477_n1449) );
  FADDX1_HVT DP_OP_423J2_125_3477_U881 ( .A(DP_OP_423J2_125_3477_n1626), .B(
        DP_OP_423J2_125_3477_n1650), .CI(DP_OP_423J2_125_3477_n1648), .CO(
        DP_OP_423J2_125_3477_n1446), .S(DP_OP_423J2_125_3477_n1447) );
  FADDX1_HVT DP_OP_423J2_125_3477_U880 ( .A(DP_OP_423J2_125_3477_n1622), .B(
        DP_OP_423J2_125_3477_n1646), .CI(DP_OP_423J2_125_3477_n1612), .CO(
        DP_OP_423J2_125_3477_n1444), .S(DP_OP_423J2_125_3477_n1445) );
  FADDX1_HVT DP_OP_423J2_125_3477_U879 ( .A(DP_OP_423J2_125_3477_n1618), .B(
        DP_OP_423J2_125_3477_n1644), .CI(DP_OP_423J2_125_3477_n1642), .CO(
        DP_OP_423J2_125_3477_n1442), .S(DP_OP_423J2_125_3477_n1443) );
  FADDX1_HVT DP_OP_423J2_125_3477_U878 ( .A(DP_OP_423J2_125_3477_n1628), .B(
        DP_OP_423J2_125_3477_n1640), .CI(DP_OP_423J2_125_3477_n1638), .CO(
        DP_OP_423J2_125_3477_n1440), .S(DP_OP_423J2_125_3477_n1441) );
  FADDX1_HVT DP_OP_423J2_125_3477_U877 ( .A(DP_OP_423J2_125_3477_n1620), .B(
        DP_OP_423J2_125_3477_n1634), .CI(DP_OP_423J2_125_3477_n1630), .CO(
        DP_OP_423J2_125_3477_n1438), .S(DP_OP_423J2_125_3477_n1439) );
  FADDX1_HVT DP_OP_423J2_125_3477_U876 ( .A(DP_OP_423J2_125_3477_n1616), .B(
        DP_OP_423J2_125_3477_n1624), .CI(DP_OP_423J2_125_3477_n1614), .CO(
        DP_OP_423J2_125_3477_n1436), .S(DP_OP_423J2_125_3477_n1437) );
  FADDX1_HVT DP_OP_423J2_125_3477_U875 ( .A(DP_OP_423J2_125_3477_n1525), .B(
        DP_OP_423J2_125_3477_n1509), .CI(DP_OP_423J2_125_3477_n1610), .CO(
        DP_OP_423J2_125_3477_n1434), .S(DP_OP_423J2_125_3477_n1435) );
  FADDX1_HVT DP_OP_423J2_125_3477_U874 ( .A(DP_OP_423J2_125_3477_n1523), .B(
        DP_OP_423J2_125_3477_n1511), .CI(DP_OP_423J2_125_3477_n1513), .CO(
        DP_OP_423J2_125_3477_n1432), .S(DP_OP_423J2_125_3477_n1433) );
  FADDX1_HVT DP_OP_423J2_125_3477_U873 ( .A(DP_OP_423J2_125_3477_n1519), .B(
        DP_OP_423J2_125_3477_n1517), .CI(DP_OP_423J2_125_3477_n1521), .CO(
        DP_OP_423J2_125_3477_n1430), .S(DP_OP_423J2_125_3477_n1431) );
  FADDX1_HVT DP_OP_423J2_125_3477_U872 ( .A(DP_OP_423J2_125_3477_n1515), .B(
        DP_OP_423J2_125_3477_n1495), .CI(DP_OP_423J2_125_3477_n1499), .CO(
        DP_OP_423J2_125_3477_n1428), .S(DP_OP_423J2_125_3477_n1429) );
  FADDX1_HVT DP_OP_423J2_125_3477_U871 ( .A(DP_OP_423J2_125_3477_n1497), .B(
        DP_OP_423J2_125_3477_n1505), .CI(DP_OP_423J2_125_3477_n1503), .CO(
        DP_OP_423J2_125_3477_n1426), .S(DP_OP_423J2_125_3477_n1427) );
  FADDX1_HVT DP_OP_423J2_125_3477_U870 ( .A(DP_OP_423J2_125_3477_n1507), .B(
        DP_OP_423J2_125_3477_n1485), .CI(DP_OP_423J2_125_3477_n1479), .CO(
        DP_OP_423J2_125_3477_n1424), .S(DP_OP_423J2_125_3477_n1425) );
  FADDX1_HVT DP_OP_423J2_125_3477_U869 ( .A(DP_OP_423J2_125_3477_n1487), .B(
        DP_OP_423J2_125_3477_n1483), .CI(DP_OP_423J2_125_3477_n1477), .CO(
        DP_OP_423J2_125_3477_n1422), .S(DP_OP_423J2_125_3477_n1423) );
  FADDX1_HVT DP_OP_423J2_125_3477_U868 ( .A(DP_OP_423J2_125_3477_n1489), .B(
        DP_OP_423J2_125_3477_n1463), .CI(DP_OP_423J2_125_3477_n1461), .CO(
        DP_OP_423J2_125_3477_n1420), .S(DP_OP_423J2_125_3477_n1421) );
  FADDX1_HVT DP_OP_423J2_125_3477_U867 ( .A(DP_OP_423J2_125_3477_n1475), .B(
        DP_OP_423J2_125_3477_n1471), .CI(DP_OP_423J2_125_3477_n1473), .CO(
        DP_OP_423J2_125_3477_n1418), .S(DP_OP_423J2_125_3477_n1419) );
  FADDX1_HVT DP_OP_423J2_125_3477_U866 ( .A(DP_OP_423J2_125_3477_n1481), .B(
        DP_OP_423J2_125_3477_n1459), .CI(DP_OP_423J2_125_3477_n1467), .CO(
        DP_OP_423J2_125_3477_n1416), .S(DP_OP_423J2_125_3477_n1417) );
  FADDX1_HVT DP_OP_423J2_125_3477_U865 ( .A(DP_OP_423J2_125_3477_n1469), .B(
        DP_OP_423J2_125_3477_n1493), .CI(DP_OP_423J2_125_3477_n1501), .CO(
        DP_OP_423J2_125_3477_n1414), .S(DP_OP_423J2_125_3477_n1415) );
  FADDX1_HVT DP_OP_423J2_125_3477_U864 ( .A(DP_OP_423J2_125_3477_n1465), .B(
        DP_OP_423J2_125_3477_n1491), .CI(DP_OP_423J2_125_3477_n1608), .CO(
        DP_OP_423J2_125_3477_n1412), .S(DP_OP_423J2_125_3477_n1413) );
  FADDX1_HVT DP_OP_423J2_125_3477_U863 ( .A(DP_OP_423J2_125_3477_n1606), .B(
        DP_OP_423J2_125_3477_n1604), .CI(DP_OP_423J2_125_3477_n1602), .CO(
        DP_OP_423J2_125_3477_n1410), .S(DP_OP_423J2_125_3477_n1411) );
  FADDX1_HVT DP_OP_423J2_125_3477_U862 ( .A(DP_OP_423J2_125_3477_n1594), .B(
        DP_OP_423J2_125_3477_n1600), .CI(DP_OP_423J2_125_3477_n1596), .CO(
        DP_OP_423J2_125_3477_n1408), .S(DP_OP_423J2_125_3477_n1409) );
  FADDX1_HVT DP_OP_423J2_125_3477_U861 ( .A(DP_OP_423J2_125_3477_n1598), .B(
        DP_OP_423J2_125_3477_n1592), .CI(DP_OP_423J2_125_3477_n1453), .CO(
        DP_OP_423J2_125_3477_n1406), .S(DP_OP_423J2_125_3477_n1407) );
  FADDX1_HVT DP_OP_423J2_125_3477_U860 ( .A(DP_OP_423J2_125_3477_n1455), .B(
        DP_OP_423J2_125_3477_n1590), .CI(DP_OP_423J2_125_3477_n1586), .CO(
        DP_OP_423J2_125_3477_n1404), .S(DP_OP_423J2_125_3477_n1405) );
  FADDX1_HVT DP_OP_423J2_125_3477_U859 ( .A(DP_OP_423J2_125_3477_n1457), .B(
        DP_OP_423J2_125_3477_n1588), .CI(DP_OP_423J2_125_3477_n1584), .CO(
        DP_OP_423J2_125_3477_n1402), .S(DP_OP_423J2_125_3477_n1403) );
  FADDX1_HVT DP_OP_423J2_125_3477_U858 ( .A(DP_OP_423J2_125_3477_n1574), .B(
        DP_OP_423J2_125_3477_n1437), .CI(DP_OP_423J2_125_3477_n1449), .CO(
        DP_OP_423J2_125_3477_n1400), .S(DP_OP_423J2_125_3477_n1401) );
  FADDX1_HVT DP_OP_423J2_125_3477_U857 ( .A(DP_OP_423J2_125_3477_n1582), .B(
        DP_OP_423J2_125_3477_n1451), .CI(DP_OP_423J2_125_3477_n1447), .CO(
        DP_OP_423J2_125_3477_n1398), .S(DP_OP_423J2_125_3477_n1399) );
  FADDX1_HVT DP_OP_423J2_125_3477_U856 ( .A(DP_OP_423J2_125_3477_n1580), .B(
        DP_OP_423J2_125_3477_n1439), .CI(DP_OP_423J2_125_3477_n1441), .CO(
        DP_OP_423J2_125_3477_n1396), .S(DP_OP_423J2_125_3477_n1397) );
  FADDX1_HVT DP_OP_423J2_125_3477_U855 ( .A(DP_OP_423J2_125_3477_n1578), .B(
        DP_OP_423J2_125_3477_n1445), .CI(DP_OP_423J2_125_3477_n1443), .CO(
        DP_OP_423J2_125_3477_n1394), .S(DP_OP_423J2_125_3477_n1395) );
  FADDX1_HVT DP_OP_423J2_125_3477_U854 ( .A(DP_OP_423J2_125_3477_n1576), .B(
        DP_OP_423J2_125_3477_n1572), .CI(DP_OP_423J2_125_3477_n1433), .CO(
        DP_OP_423J2_125_3477_n1392), .S(DP_OP_423J2_125_3477_n1393) );
  FADDX1_HVT DP_OP_423J2_125_3477_U853 ( .A(DP_OP_423J2_125_3477_n1435), .B(
        DP_OP_423J2_125_3477_n1431), .CI(DP_OP_423J2_125_3477_n1429), .CO(
        DP_OP_423J2_125_3477_n1390), .S(DP_OP_423J2_125_3477_n1391) );
  FADDX1_HVT DP_OP_423J2_125_3477_U852 ( .A(DP_OP_423J2_125_3477_n1570), .B(
        DP_OP_423J2_125_3477_n1421), .CI(DP_OP_423J2_125_3477_n1419), .CO(
        DP_OP_423J2_125_3477_n1388), .S(DP_OP_423J2_125_3477_n1389) );
  FADDX1_HVT DP_OP_423J2_125_3477_U851 ( .A(DP_OP_423J2_125_3477_n1425), .B(
        DP_OP_423J2_125_3477_n1415), .CI(DP_OP_423J2_125_3477_n1417), .CO(
        DP_OP_423J2_125_3477_n1386), .S(DP_OP_423J2_125_3477_n1387) );
  FADDX1_HVT DP_OP_423J2_125_3477_U850 ( .A(DP_OP_423J2_125_3477_n1423), .B(
        DP_OP_423J2_125_3477_n1427), .CI(DP_OP_423J2_125_3477_n1568), .CO(
        DP_OP_423J2_125_3477_n1384), .S(DP_OP_423J2_125_3477_n1385) );
  FADDX1_HVT DP_OP_423J2_125_3477_U849 ( .A(DP_OP_423J2_125_3477_n1566), .B(
        DP_OP_423J2_125_3477_n1413), .CI(DP_OP_423J2_125_3477_n1564), .CO(
        DP_OP_423J2_125_3477_n1382), .S(DP_OP_423J2_125_3477_n1383) );
  FADDX1_HVT DP_OP_423J2_125_3477_U848 ( .A(DP_OP_423J2_125_3477_n1562), .B(
        DP_OP_423J2_125_3477_n1409), .CI(DP_OP_423J2_125_3477_n1411), .CO(
        DP_OP_423J2_125_3477_n1380), .S(DP_OP_423J2_125_3477_n1381) );
  FADDX1_HVT DP_OP_423J2_125_3477_U847 ( .A(DP_OP_423J2_125_3477_n1560), .B(
        DP_OP_423J2_125_3477_n1556), .CI(DP_OP_423J2_125_3477_n1558), .CO(
        DP_OP_423J2_125_3477_n1378), .S(DP_OP_423J2_125_3477_n1379) );
  FADDX1_HVT DP_OP_423J2_125_3477_U846 ( .A(DP_OP_423J2_125_3477_n1407), .B(
        DP_OP_423J2_125_3477_n1554), .CI(DP_OP_423J2_125_3477_n1552), .CO(
        DP_OP_423J2_125_3477_n1376), .S(DP_OP_423J2_125_3477_n1377) );
  FADDX1_HVT DP_OP_423J2_125_3477_U845 ( .A(DP_OP_423J2_125_3477_n1405), .B(
        DP_OP_423J2_125_3477_n1403), .CI(DP_OP_423J2_125_3477_n1399), .CO(
        DP_OP_423J2_125_3477_n1374), .S(DP_OP_423J2_125_3477_n1375) );
  FADDX1_HVT DP_OP_423J2_125_3477_U844 ( .A(DP_OP_423J2_125_3477_n1401), .B(
        DP_OP_423J2_125_3477_n1397), .CI(DP_OP_423J2_125_3477_n1393), .CO(
        DP_OP_423J2_125_3477_n1372), .S(DP_OP_423J2_125_3477_n1373) );
  FADDX1_HVT DP_OP_423J2_125_3477_U843 ( .A(DP_OP_423J2_125_3477_n1550), .B(
        DP_OP_423J2_125_3477_n1395), .CI(DP_OP_423J2_125_3477_n1548), .CO(
        DP_OP_423J2_125_3477_n1370), .S(DP_OP_423J2_125_3477_n1371) );
  FADDX1_HVT DP_OP_423J2_125_3477_U842 ( .A(DP_OP_423J2_125_3477_n1391), .B(
        DP_OP_423J2_125_3477_n1389), .CI(DP_OP_423J2_125_3477_n1387), .CO(
        DP_OP_423J2_125_3477_n1368), .S(DP_OP_423J2_125_3477_n1369) );
  FADDX1_HVT DP_OP_423J2_125_3477_U841 ( .A(DP_OP_423J2_125_3477_n1546), .B(
        DP_OP_423J2_125_3477_n1385), .CI(DP_OP_423J2_125_3477_n1544), .CO(
        DP_OP_423J2_125_3477_n1366), .S(DP_OP_423J2_125_3477_n1367) );
  FADDX1_HVT DP_OP_423J2_125_3477_U840 ( .A(DP_OP_423J2_125_3477_n1383), .B(
        DP_OP_423J2_125_3477_n1542), .CI(DP_OP_423J2_125_3477_n1540), .CO(
        DP_OP_423J2_125_3477_n1364), .S(DP_OP_423J2_125_3477_n1365) );
  FADDX1_HVT DP_OP_423J2_125_3477_U839 ( .A(DP_OP_423J2_125_3477_n1379), .B(
        DP_OP_423J2_125_3477_n1381), .CI(DP_OP_423J2_125_3477_n1538), .CO(
        DP_OP_423J2_125_3477_n1362), .S(DP_OP_423J2_125_3477_n1363) );
  FADDX1_HVT DP_OP_423J2_125_3477_U838 ( .A(DP_OP_423J2_125_3477_n1377), .B(
        DP_OP_423J2_125_3477_n1375), .CI(DP_OP_423J2_125_3477_n1536), .CO(
        DP_OP_423J2_125_3477_n1360), .S(DP_OP_423J2_125_3477_n1361) );
  FADDX1_HVT DP_OP_423J2_125_3477_U837 ( .A(DP_OP_423J2_125_3477_n1371), .B(
        DP_OP_423J2_125_3477_n1373), .CI(DP_OP_423J2_125_3477_n1534), .CO(
        DP_OP_423J2_125_3477_n1358), .S(DP_OP_423J2_125_3477_n1359) );
  FADDX1_HVT DP_OP_423J2_125_3477_U836 ( .A(DP_OP_423J2_125_3477_n1369), .B(
        DP_OP_423J2_125_3477_n1367), .CI(DP_OP_423J2_125_3477_n1532), .CO(
        DP_OP_423J2_125_3477_n1356), .S(DP_OP_423J2_125_3477_n1357) );
  FADDX1_HVT DP_OP_423J2_125_3477_U835 ( .A(DP_OP_423J2_125_3477_n1365), .B(
        DP_OP_423J2_125_3477_n1530), .CI(DP_OP_423J2_125_3477_n1363), .CO(
        DP_OP_423J2_125_3477_n1354), .S(DP_OP_423J2_125_3477_n1355) );
  FADDX1_HVT DP_OP_423J2_125_3477_U834 ( .A(DP_OP_423J2_125_3477_n1361), .B(
        DP_OP_423J2_125_3477_n1528), .CI(DP_OP_423J2_125_3477_n1359), .CO(
        DP_OP_423J2_125_3477_n1352), .S(DP_OP_423J2_125_3477_n1353) );
  FADDX1_HVT DP_OP_423J2_125_3477_U833 ( .A(DP_OP_423J2_125_3477_n1357), .B(
        DP_OP_423J2_125_3477_n1526), .CI(DP_OP_423J2_125_3477_n1355), .CO(
        DP_OP_423J2_125_3477_n1350), .S(DP_OP_423J2_125_3477_n1351) );
  HADDX1_HVT DP_OP_423J2_125_3477_U832 ( .A0(DP_OP_423J2_125_3477_n2980), .B0(
        DP_OP_423J2_125_3477_n1925), .C1(DP_OP_423J2_125_3477_n1348), .SO(
        DP_OP_423J2_125_3477_n1349) );
  FADDX1_HVT DP_OP_423J2_125_3477_U831 ( .A(DP_OP_423J2_125_3477_n2453), .B(
        DP_OP_423J2_125_3477_n2365), .CI(DP_OP_423J2_125_3477_n1881), .CO(
        DP_OP_423J2_125_3477_n1346), .S(DP_OP_423J2_125_3477_n1347) );
  FADDX1_HVT DP_OP_423J2_125_3477_U830 ( .A(DP_OP_423J2_125_3477_n2497), .B(
        DP_OP_423J2_125_3477_n2277), .CI(DP_OP_423J2_125_3477_n2321), .CO(
        DP_OP_423J2_125_3477_n1344), .S(DP_OP_423J2_125_3477_n1345) );
  FADDX1_HVT DP_OP_423J2_125_3477_U829 ( .A(DP_OP_423J2_125_3477_n2805), .B(
        DP_OP_423J2_125_3477_n1969), .CI(DP_OP_423J2_125_3477_n2057), .CO(
        DP_OP_423J2_125_3477_n1342), .S(DP_OP_423J2_125_3477_n1343) );
  FADDX1_HVT DP_OP_423J2_125_3477_U828 ( .A(DP_OP_423J2_125_3477_n2541), .B(
        DP_OP_423J2_125_3477_n2101), .CI(DP_OP_423J2_125_3477_n2629), .CO(
        DP_OP_423J2_125_3477_n1340), .S(DP_OP_423J2_125_3477_n1341) );
  FADDX1_HVT DP_OP_423J2_125_3477_U827 ( .A(DP_OP_423J2_125_3477_n2013), .B(
        DP_OP_423J2_125_3477_n2849), .CI(DP_OP_423J2_125_3477_n2145), .CO(
        DP_OP_423J2_125_3477_n1338), .S(DP_OP_423J2_125_3477_n1339) );
  FADDX1_HVT DP_OP_423J2_125_3477_U826 ( .A(DP_OP_423J2_125_3477_n2409), .B(
        DP_OP_423J2_125_3477_n2893), .CI(DP_OP_423J2_125_3477_n2717), .CO(
        DP_OP_423J2_125_3477_n1336), .S(DP_OP_423J2_125_3477_n1337) );
  FADDX1_HVT DP_OP_423J2_125_3477_U825 ( .A(DP_OP_423J2_125_3477_n2233), .B(
        DP_OP_423J2_125_3477_n2189), .CI(DP_OP_423J2_125_3477_n2673), .CO(
        DP_OP_423J2_125_3477_n1334), .S(DP_OP_423J2_125_3477_n1335) );
  FADDX1_HVT DP_OP_423J2_125_3477_U824 ( .A(DP_OP_423J2_125_3477_n2937), .B(
        DP_OP_423J2_125_3477_n2585), .CI(DP_OP_423J2_125_3477_n2761), .CO(
        DP_OP_423J2_125_3477_n1332), .S(DP_OP_423J2_125_3477_n1333) );
  FADDX1_HVT DP_OP_423J2_125_3477_U823 ( .A(DP_OP_423J2_125_3477_n2379), .B(
        DP_OP_423J2_125_3477_n3000), .CI(DP_OP_423J2_125_3477_n1932), .CO(
        DP_OP_423J2_125_3477_n1330), .S(DP_OP_423J2_125_3477_n1331) );
  FADDX1_HVT DP_OP_423J2_125_3477_U822 ( .A(DP_OP_423J2_125_3477_n2372), .B(
        DP_OP_423J2_125_3477_n1939), .CI(DP_OP_423J2_125_3477_n1946), .CO(
        DP_OP_423J2_125_3477_n1328), .S(DP_OP_423J2_125_3477_n1329) );
  FADDX1_HVT DP_OP_423J2_125_3477_U821 ( .A(DP_OP_423J2_125_3477_n2386), .B(
        DP_OP_423J2_125_3477_n1976), .CI(DP_OP_423J2_125_3477_n2993), .CO(
        DP_OP_423J2_125_3477_n1326), .S(DP_OP_423J2_125_3477_n1327) );
  FADDX1_HVT DP_OP_423J2_125_3477_U820 ( .A(DP_OP_423J2_125_3477_n2342), .B(
        DP_OP_423J2_125_3477_n2986), .CI(DP_OP_423J2_125_3477_n2958), .CO(
        DP_OP_423J2_125_3477_n1324), .S(DP_OP_423J2_125_3477_n1325) );
  FADDX1_HVT DP_OP_423J2_125_3477_U819 ( .A(DP_OP_423J2_125_3477_n2335), .B(
        DP_OP_423J2_125_3477_n2951), .CI(DP_OP_423J2_125_3477_n2944), .CO(
        DP_OP_423J2_125_3477_n1322), .S(DP_OP_423J2_125_3477_n1323) );
  FADDX1_HVT DP_OP_423J2_125_3477_U818 ( .A(DP_OP_423J2_125_3477_n2298), .B(
        DP_OP_423J2_125_3477_n2914), .CI(DP_OP_423J2_125_3477_n2907), .CO(
        DP_OP_423J2_125_3477_n1320), .S(DP_OP_423J2_125_3477_n1321) );
  FADDX1_HVT DP_OP_423J2_125_3477_U817 ( .A(DP_OP_423J2_125_3477_n2291), .B(
        DP_OP_423J2_125_3477_n1983), .CI(DP_OP_423J2_125_3477_n2900), .CO(
        DP_OP_423J2_125_3477_n1318), .S(DP_OP_423J2_125_3477_n1319) );
  FADDX1_HVT DP_OP_423J2_125_3477_U816 ( .A(DP_OP_423J2_125_3477_n2284), .B(
        DP_OP_423J2_125_3477_n2870), .CI(DP_OP_423J2_125_3477_n2863), .CO(
        DP_OP_423J2_125_3477_n1316), .S(DP_OP_423J2_125_3477_n1317) );
  FADDX1_HVT DP_OP_423J2_125_3477_U815 ( .A(DP_OP_423J2_125_3477_n2254), .B(
        DP_OP_423J2_125_3477_n2856), .CI(DP_OP_423J2_125_3477_n1990), .CO(
        DP_OP_423J2_125_3477_n1314), .S(DP_OP_423J2_125_3477_n1315) );
  FADDX1_HVT DP_OP_423J2_125_3477_U814 ( .A(DP_OP_423J2_125_3477_n2247), .B(
        DP_OP_423J2_125_3477_n2020), .CI(DP_OP_423J2_125_3477_n2027), .CO(
        DP_OP_423J2_125_3477_n1312), .S(DP_OP_423J2_125_3477_n1313) );
  FADDX1_HVT DP_OP_423J2_125_3477_U813 ( .A(DP_OP_423J2_125_3477_n2328), .B(
        DP_OP_423J2_125_3477_n2034), .CI(DP_OP_423J2_125_3477_n2826), .CO(
        DP_OP_423J2_125_3477_n1310), .S(DP_OP_423J2_125_3477_n1311) );
  FADDX1_HVT DP_OP_423J2_125_3477_U812 ( .A(DP_OP_423J2_125_3477_n2416), .B(
        DP_OP_423J2_125_3477_n2819), .CI(DP_OP_423J2_125_3477_n2064), .CO(
        DP_OP_423J2_125_3477_n1308), .S(DP_OP_423J2_125_3477_n1309) );
  FADDX1_HVT DP_OP_423J2_125_3477_U811 ( .A(DP_OP_423J2_125_3477_n2812), .B(
        DP_OP_423J2_125_3477_n2071), .CI(DP_OP_423J2_125_3477_n2078), .CO(
        DP_OP_423J2_125_3477_n1306), .S(DP_OP_423J2_125_3477_n1307) );
  FADDX1_HVT DP_OP_423J2_125_3477_U810 ( .A(DP_OP_423J2_125_3477_n2782), .B(
        DP_OP_423J2_125_3477_n2108), .CI(DP_OP_423J2_125_3477_n2115), .CO(
        DP_OP_423J2_125_3477_n1304), .S(DP_OP_423J2_125_3477_n1305) );
  FADDX1_HVT DP_OP_423J2_125_3477_U809 ( .A(DP_OP_423J2_125_3477_n2775), .B(
        DP_OP_423J2_125_3477_n2122), .CI(DP_OP_423J2_125_3477_n2152), .CO(
        DP_OP_423J2_125_3477_n1302), .S(DP_OP_423J2_125_3477_n1303) );
  FADDX1_HVT DP_OP_423J2_125_3477_U808 ( .A(DP_OP_423J2_125_3477_n2768), .B(
        DP_OP_423J2_125_3477_n2159), .CI(DP_OP_423J2_125_3477_n2166), .CO(
        DP_OP_423J2_125_3477_n1300), .S(DP_OP_423J2_125_3477_n1301) );
  FADDX1_HVT DP_OP_423J2_125_3477_U807 ( .A(DP_OP_423J2_125_3477_n2738), .B(
        DP_OP_423J2_125_3477_n2196), .CI(DP_OP_423J2_125_3477_n2203), .CO(
        DP_OP_423J2_125_3477_n1298), .S(DP_OP_423J2_125_3477_n1299) );
  FADDX1_HVT DP_OP_423J2_125_3477_U806 ( .A(DP_OP_423J2_125_3477_n2731), .B(
        DP_OP_423J2_125_3477_n2210), .CI(DP_OP_423J2_125_3477_n2240), .CO(
        DP_OP_423J2_125_3477_n1296), .S(DP_OP_423J2_125_3477_n1297) );
  FADDX1_HVT DP_OP_423J2_125_3477_U805 ( .A(DP_OP_423J2_125_3477_n2724), .B(
        DP_OP_423J2_125_3477_n2423), .CI(DP_OP_423J2_125_3477_n2430), .CO(
        DP_OP_423J2_125_3477_n1294), .S(DP_OP_423J2_125_3477_n1295) );
  FADDX1_HVT DP_OP_423J2_125_3477_U804 ( .A(DP_OP_423J2_125_3477_n2694), .B(
        DP_OP_423J2_125_3477_n2460), .CI(DP_OP_423J2_125_3477_n2467), .CO(
        DP_OP_423J2_125_3477_n1292), .S(DP_OP_423J2_125_3477_n1293) );
  FADDX1_HVT DP_OP_423J2_125_3477_U803 ( .A(DP_OP_423J2_125_3477_n2687), .B(
        DP_OP_423J2_125_3477_n2474), .CI(DP_OP_423J2_125_3477_n2504), .CO(
        DP_OP_423J2_125_3477_n1290), .S(DP_OP_423J2_125_3477_n1291) );
  FADDX1_HVT DP_OP_423J2_125_3477_U802 ( .A(DP_OP_423J2_125_3477_n2680), .B(
        DP_OP_423J2_125_3477_n2511), .CI(DP_OP_423J2_125_3477_n2518), .CO(
        DP_OP_423J2_125_3477_n1288), .S(DP_OP_423J2_125_3477_n1289) );
  FADDX1_HVT DP_OP_423J2_125_3477_U801 ( .A(DP_OP_423J2_125_3477_n2650), .B(
        DP_OP_423J2_125_3477_n2643), .CI(DP_OP_423J2_125_3477_n2636), .CO(
        DP_OP_423J2_125_3477_n1286), .S(DP_OP_423J2_125_3477_n1287) );
  FADDX1_HVT DP_OP_423J2_125_3477_U800 ( .A(DP_OP_423J2_125_3477_n2592), .B(
        DP_OP_423J2_125_3477_n2606), .CI(DP_OP_423J2_125_3477_n2548), .CO(
        DP_OP_423J2_125_3477_n1284), .S(DP_OP_423J2_125_3477_n1285) );
  FADDX1_HVT DP_OP_423J2_125_3477_U799 ( .A(DP_OP_423J2_125_3477_n2555), .B(
        DP_OP_423J2_125_3477_n2562), .CI(DP_OP_423J2_125_3477_n2599), .CO(
        DP_OP_423J2_125_3477_n1282), .S(DP_OP_423J2_125_3477_n1283) );
  FADDX1_HVT DP_OP_423J2_125_3477_U798 ( .A(DP_OP_423J2_125_3477_n1349), .B(
        DP_OP_423J2_125_3477_n1524), .CI(DP_OP_423J2_125_3477_n1514), .CO(
        DP_OP_423J2_125_3477_n1280), .S(DP_OP_423J2_125_3477_n1281) );
  FADDX1_HVT DP_OP_423J2_125_3477_U797 ( .A(DP_OP_423J2_125_3477_n1522), .B(
        DP_OP_423J2_125_3477_n1520), .CI(DP_OP_423J2_125_3477_n1518), .CO(
        DP_OP_423J2_125_3477_n1278), .S(DP_OP_423J2_125_3477_n1279) );
  FADDX1_HVT DP_OP_423J2_125_3477_U796 ( .A(DP_OP_423J2_125_3477_n1516), .B(
        DP_OP_423J2_125_3477_n1512), .CI(DP_OP_423J2_125_3477_n1508), .CO(
        DP_OP_423J2_125_3477_n1276), .S(DP_OP_423J2_125_3477_n1277) );
  FADDX1_HVT DP_OP_423J2_125_3477_U795 ( .A(DP_OP_423J2_125_3477_n1510), .B(
        DP_OP_423J2_125_3477_n1484), .CI(DP_OP_423J2_125_3477_n1482), .CO(
        DP_OP_423J2_125_3477_n1274), .S(DP_OP_423J2_125_3477_n1275) );
  FADDX1_HVT DP_OP_423J2_125_3477_U794 ( .A(DP_OP_423J2_125_3477_n1486), .B(
        DP_OP_423J2_125_3477_n1458), .CI(DP_OP_423J2_125_3477_n1506), .CO(
        DP_OP_423J2_125_3477_n1272), .S(DP_OP_423J2_125_3477_n1273) );
  FADDX1_HVT DP_OP_423J2_125_3477_U793 ( .A(DP_OP_423J2_125_3477_n1478), .B(
        DP_OP_423J2_125_3477_n1504), .CI(DP_OP_423J2_125_3477_n1502), .CO(
        DP_OP_423J2_125_3477_n1270), .S(DP_OP_423J2_125_3477_n1271) );
  FADDX1_HVT DP_OP_423J2_125_3477_U792 ( .A(DP_OP_423J2_125_3477_n1474), .B(
        DP_OP_423J2_125_3477_n1500), .CI(DP_OP_423J2_125_3477_n1498), .CO(
        DP_OP_423J2_125_3477_n1268), .S(DP_OP_423J2_125_3477_n1269) );
  FADDX1_HVT DP_OP_423J2_125_3477_U791 ( .A(DP_OP_423J2_125_3477_n1468), .B(
        DP_OP_423J2_125_3477_n1460), .CI(DP_OP_423J2_125_3477_n1462), .CO(
        DP_OP_423J2_125_3477_n1266), .S(DP_OP_423J2_125_3477_n1267) );
  FADDX1_HVT DP_OP_423J2_125_3477_U790 ( .A(DP_OP_423J2_125_3477_n1466), .B(
        DP_OP_423J2_125_3477_n1496), .CI(DP_OP_423J2_125_3477_n1494), .CO(
        DP_OP_423J2_125_3477_n1264), .S(DP_OP_423J2_125_3477_n1265) );
  FADDX1_HVT DP_OP_423J2_125_3477_U789 ( .A(DP_OP_423J2_125_3477_n1476), .B(
        DP_OP_423J2_125_3477_n1492), .CI(DP_OP_423J2_125_3477_n1464), .CO(
        DP_OP_423J2_125_3477_n1262), .S(DP_OP_423J2_125_3477_n1263) );
  FADDX1_HVT DP_OP_423J2_125_3477_U788 ( .A(DP_OP_423J2_125_3477_n1472), .B(
        DP_OP_423J2_125_3477_n1490), .CI(DP_OP_423J2_125_3477_n1488), .CO(
        DP_OP_423J2_125_3477_n1260), .S(DP_OP_423J2_125_3477_n1261) );
  FADDX1_HVT DP_OP_423J2_125_3477_U787 ( .A(DP_OP_423J2_125_3477_n1470), .B(
        DP_OP_423J2_125_3477_n1480), .CI(DP_OP_423J2_125_3477_n1339), .CO(
        DP_OP_423J2_125_3477_n1258), .S(DP_OP_423J2_125_3477_n1259) );
  FADDX1_HVT DP_OP_423J2_125_3477_U786 ( .A(DP_OP_423J2_125_3477_n1341), .B(
        DP_OP_423J2_125_3477_n1333), .CI(DP_OP_423J2_125_3477_n1335), .CO(
        DP_OP_423J2_125_3477_n1256), .S(DP_OP_423J2_125_3477_n1257) );
  FADDX1_HVT DP_OP_423J2_125_3477_U785 ( .A(DP_OP_423J2_125_3477_n1345), .B(
        DP_OP_423J2_125_3477_n1343), .CI(DP_OP_423J2_125_3477_n1347), .CO(
        DP_OP_423J2_125_3477_n1254), .S(DP_OP_423J2_125_3477_n1255) );
  FADDX1_HVT DP_OP_423J2_125_3477_U784 ( .A(DP_OP_423J2_125_3477_n1337), .B(
        DP_OP_423J2_125_3477_n1289), .CI(DP_OP_423J2_125_3477_n1287), .CO(
        DP_OP_423J2_125_3477_n1252), .S(DP_OP_423J2_125_3477_n1253) );
  FADDX1_HVT DP_OP_423J2_125_3477_U783 ( .A(DP_OP_423J2_125_3477_n1283), .B(
        DP_OP_423J2_125_3477_n1331), .CI(DP_OP_423J2_125_3477_n1329), .CO(
        DP_OP_423J2_125_3477_n1250), .S(DP_OP_423J2_125_3477_n1251) );
  FADDX1_HVT DP_OP_423J2_125_3477_U782 ( .A(DP_OP_423J2_125_3477_n1319), .B(
        DP_OP_423J2_125_3477_n1309), .CI(DP_OP_423J2_125_3477_n1315), .CO(
        DP_OP_423J2_125_3477_n1248), .S(DP_OP_423J2_125_3477_n1249) );
  FADDX1_HVT DP_OP_423J2_125_3477_U781 ( .A(DP_OP_423J2_125_3477_n1313), .B(
        DP_OP_423J2_125_3477_n1311), .CI(DP_OP_423J2_125_3477_n1295), .CO(
        DP_OP_423J2_125_3477_n1246), .S(DP_OP_423J2_125_3477_n1247) );
  FADDX1_HVT DP_OP_423J2_125_3477_U780 ( .A(DP_OP_423J2_125_3477_n1317), .B(
        DP_OP_423J2_125_3477_n1291), .CI(DP_OP_423J2_125_3477_n1285), .CO(
        DP_OP_423J2_125_3477_n1244), .S(DP_OP_423J2_125_3477_n1245) );
  FADDX1_HVT DP_OP_423J2_125_3477_U779 ( .A(DP_OP_423J2_125_3477_n1321), .B(
        DP_OP_423J2_125_3477_n1303), .CI(DP_OP_423J2_125_3477_n1305), .CO(
        DP_OP_423J2_125_3477_n1242), .S(DP_OP_423J2_125_3477_n1243) );
  FADDX1_HVT DP_OP_423J2_125_3477_U778 ( .A(DP_OP_423J2_125_3477_n1301), .B(
        DP_OP_423J2_125_3477_n1299), .CI(DP_OP_423J2_125_3477_n1293), .CO(
        DP_OP_423J2_125_3477_n1240), .S(DP_OP_423J2_125_3477_n1241) );
  FADDX1_HVT DP_OP_423J2_125_3477_U777 ( .A(DP_OP_423J2_125_3477_n1297), .B(
        DP_OP_423J2_125_3477_n1327), .CI(DP_OP_423J2_125_3477_n1323), .CO(
        DP_OP_423J2_125_3477_n1238), .S(DP_OP_423J2_125_3477_n1239) );
  FADDX1_HVT DP_OP_423J2_125_3477_U776 ( .A(DP_OP_423J2_125_3477_n1325), .B(
        DP_OP_423J2_125_3477_n1307), .CI(DP_OP_423J2_125_3477_n1456), .CO(
        DP_OP_423J2_125_3477_n1236), .S(DP_OP_423J2_125_3477_n1237) );
  FADDX1_HVT DP_OP_423J2_125_3477_U775 ( .A(DP_OP_423J2_125_3477_n1454), .B(
        DP_OP_423J2_125_3477_n1452), .CI(DP_OP_423J2_125_3477_n1450), .CO(
        DP_OP_423J2_125_3477_n1234), .S(DP_OP_423J2_125_3477_n1235) );
  FADDX1_HVT DP_OP_423J2_125_3477_U774 ( .A(DP_OP_423J2_125_3477_n1448), .B(
        DP_OP_423J2_125_3477_n1436), .CI(DP_OP_423J2_125_3477_n1438), .CO(
        DP_OP_423J2_125_3477_n1232), .S(DP_OP_423J2_125_3477_n1233) );
  FADDX1_HVT DP_OP_423J2_125_3477_U773 ( .A(DP_OP_423J2_125_3477_n1442), .B(
        DP_OP_423J2_125_3477_n1446), .CI(DP_OP_423J2_125_3477_n1440), .CO(
        DP_OP_423J2_125_3477_n1230), .S(DP_OP_423J2_125_3477_n1231) );
  FADDX1_HVT DP_OP_423J2_125_3477_U772 ( .A(DP_OP_423J2_125_3477_n1444), .B(
        DP_OP_423J2_125_3477_n1281), .CI(DP_OP_423J2_125_3477_n1434), .CO(
        DP_OP_423J2_125_3477_n1228), .S(DP_OP_423J2_125_3477_n1229) );
  FADDX1_HVT DP_OP_423J2_125_3477_U771 ( .A(DP_OP_423J2_125_3477_n1279), .B(
        DP_OP_423J2_125_3477_n1277), .CI(DP_OP_423J2_125_3477_n1275), .CO(
        DP_OP_423J2_125_3477_n1226), .S(DP_OP_423J2_125_3477_n1227) );
  FADDX1_HVT DP_OP_423J2_125_3477_U770 ( .A(DP_OP_423J2_125_3477_n1432), .B(
        DP_OP_423J2_125_3477_n1430), .CI(DP_OP_423J2_125_3477_n1428), .CO(
        DP_OP_423J2_125_3477_n1224), .S(DP_OP_423J2_125_3477_n1225) );
  FADDX1_HVT DP_OP_423J2_125_3477_U769 ( .A(DP_OP_423J2_125_3477_n1416), .B(
        DP_OP_423J2_125_3477_n1261), .CI(DP_OP_423J2_125_3477_n1259), .CO(
        DP_OP_423J2_125_3477_n1222), .S(DP_OP_423J2_125_3477_n1223) );
  FADDX1_HVT DP_OP_423J2_125_3477_U768 ( .A(DP_OP_423J2_125_3477_n1426), .B(
        DP_OP_423J2_125_3477_n1271), .CI(DP_OP_423J2_125_3477_n1273), .CO(
        DP_OP_423J2_125_3477_n1220), .S(DP_OP_423J2_125_3477_n1221) );
  FADDX1_HVT DP_OP_423J2_125_3477_U767 ( .A(DP_OP_423J2_125_3477_n1424), .B(
        DP_OP_423J2_125_3477_n1267), .CI(DP_OP_423J2_125_3477_n1263), .CO(
        DP_OP_423J2_125_3477_n1218), .S(DP_OP_423J2_125_3477_n1219) );
  FADDX1_HVT DP_OP_423J2_125_3477_U766 ( .A(DP_OP_423J2_125_3477_n1422), .B(
        DP_OP_423J2_125_3477_n1269), .CI(DP_OP_423J2_125_3477_n1265), .CO(
        DP_OP_423J2_125_3477_n1216), .S(DP_OP_423J2_125_3477_n1217) );
  FADDX1_HVT DP_OP_423J2_125_3477_U765 ( .A(DP_OP_423J2_125_3477_n1420), .B(
        DP_OP_423J2_125_3477_n1414), .CI(DP_OP_423J2_125_3477_n1418), .CO(
        DP_OP_423J2_125_3477_n1214), .S(DP_OP_423J2_125_3477_n1215) );
  FADDX1_HVT DP_OP_423J2_125_3477_U764 ( .A(DP_OP_423J2_125_3477_n1255), .B(
        DP_OP_423J2_125_3477_n1257), .CI(DP_OP_423J2_125_3477_n1253), .CO(
        DP_OP_423J2_125_3477_n1212), .S(DP_OP_423J2_125_3477_n1213) );
  FADDX1_HVT DP_OP_423J2_125_3477_U763 ( .A(DP_OP_423J2_125_3477_n1245), .B(
        DP_OP_423J2_125_3477_n1247), .CI(DP_OP_423J2_125_3477_n1412), .CO(
        DP_OP_423J2_125_3477_n1210), .S(DP_OP_423J2_125_3477_n1211) );
  FADDX1_HVT DP_OP_423J2_125_3477_U762 ( .A(DP_OP_423J2_125_3477_n1243), .B(
        DP_OP_423J2_125_3477_n1251), .CI(DP_OP_423J2_125_3477_n1249), .CO(
        DP_OP_423J2_125_3477_n1208), .S(DP_OP_423J2_125_3477_n1209) );
  FADDX1_HVT DP_OP_423J2_125_3477_U761 ( .A(DP_OP_423J2_125_3477_n1239), .B(
        DP_OP_423J2_125_3477_n1241), .CI(DP_OP_423J2_125_3477_n1408), .CO(
        DP_OP_423J2_125_3477_n1206), .S(DP_OP_423J2_125_3477_n1207) );
  FADDX1_HVT DP_OP_423J2_125_3477_U760 ( .A(DP_OP_423J2_125_3477_n1410), .B(
        DP_OP_423J2_125_3477_n1237), .CI(DP_OP_423J2_125_3477_n1406), .CO(
        DP_OP_423J2_125_3477_n1204), .S(DP_OP_423J2_125_3477_n1205) );
  FADDX1_HVT DP_OP_423J2_125_3477_U759 ( .A(DP_OP_423J2_125_3477_n1404), .B(
        DP_OP_423J2_125_3477_n1402), .CI(DP_OP_423J2_125_3477_n1235), .CO(
        DP_OP_423J2_125_3477_n1202), .S(DP_OP_423J2_125_3477_n1203) );
  FADDX1_HVT DP_OP_423J2_125_3477_U758 ( .A(DP_OP_423J2_125_3477_n1400), .B(
        DP_OP_423J2_125_3477_n1392), .CI(DP_OP_423J2_125_3477_n1229), .CO(
        DP_OP_423J2_125_3477_n1200), .S(DP_OP_423J2_125_3477_n1201) );
  FADDX1_HVT DP_OP_423J2_125_3477_U757 ( .A(DP_OP_423J2_125_3477_n1398), .B(
        DP_OP_423J2_125_3477_n1231), .CI(DP_OP_423J2_125_3477_n1233), .CO(
        DP_OP_423J2_125_3477_n1198), .S(DP_OP_423J2_125_3477_n1199) );
  FADDX1_HVT DP_OP_423J2_125_3477_U756 ( .A(DP_OP_423J2_125_3477_n1396), .B(
        DP_OP_423J2_125_3477_n1394), .CI(DP_OP_423J2_125_3477_n1390), .CO(
        DP_OP_423J2_125_3477_n1196), .S(DP_OP_423J2_125_3477_n1197) );
  FADDX1_HVT DP_OP_423J2_125_3477_U755 ( .A(DP_OP_423J2_125_3477_n1225), .B(
        DP_OP_423J2_125_3477_n1227), .CI(DP_OP_423J2_125_3477_n1388), .CO(
        DP_OP_423J2_125_3477_n1194), .S(DP_OP_423J2_125_3477_n1195) );
  FADDX1_HVT DP_OP_423J2_125_3477_U754 ( .A(DP_OP_423J2_125_3477_n1386), .B(
        DP_OP_423J2_125_3477_n1219), .CI(DP_OP_423J2_125_3477_n1384), .CO(
        DP_OP_423J2_125_3477_n1192), .S(DP_OP_423J2_125_3477_n1193) );
  FADDX1_HVT DP_OP_423J2_125_3477_U753 ( .A(DP_OP_423J2_125_3477_n1217), .B(
        DP_OP_423J2_125_3477_n1223), .CI(DP_OP_423J2_125_3477_n1221), .CO(
        DP_OP_423J2_125_3477_n1190), .S(DP_OP_423J2_125_3477_n1191) );
  FADDX1_HVT DP_OP_423J2_125_3477_U752 ( .A(DP_OP_423J2_125_3477_n1215), .B(
        DP_OP_423J2_125_3477_n1213), .CI(DP_OP_423J2_125_3477_n1209), .CO(
        DP_OP_423J2_125_3477_n1188), .S(DP_OP_423J2_125_3477_n1189) );
  FADDX1_HVT DP_OP_423J2_125_3477_U751 ( .A(DP_OP_423J2_125_3477_n1211), .B(
        DP_OP_423J2_125_3477_n1382), .CI(DP_OP_423J2_125_3477_n1207), .CO(
        DP_OP_423J2_125_3477_n1186), .S(DP_OP_423J2_125_3477_n1187) );
  FADDX1_HVT DP_OP_423J2_125_3477_U750 ( .A(DP_OP_423J2_125_3477_n1380), .B(
        DP_OP_423J2_125_3477_n1378), .CI(DP_OP_423J2_125_3477_n1205), .CO(
        DP_OP_423J2_125_3477_n1184), .S(DP_OP_423J2_125_3477_n1185) );
  FADDX1_HVT DP_OP_423J2_125_3477_U749 ( .A(DP_OP_423J2_125_3477_n1376), .B(
        DP_OP_423J2_125_3477_n1374), .CI(DP_OP_423J2_125_3477_n1203), .CO(
        DP_OP_423J2_125_3477_n1182), .S(DP_OP_423J2_125_3477_n1183) );
  FADDX1_HVT DP_OP_423J2_125_3477_U748 ( .A(DP_OP_423J2_125_3477_n1372), .B(
        DP_OP_423J2_125_3477_n1199), .CI(DP_OP_423J2_125_3477_n1197), .CO(
        DP_OP_423J2_125_3477_n1180), .S(DP_OP_423J2_125_3477_n1181) );
  FADDX1_HVT DP_OP_423J2_125_3477_U747 ( .A(DP_OP_423J2_125_3477_n1370), .B(
        DP_OP_423J2_125_3477_n1201), .CI(DP_OP_423J2_125_3477_n1195), .CO(
        DP_OP_423J2_125_3477_n1178), .S(DP_OP_423J2_125_3477_n1179) );
  FADDX1_HVT DP_OP_423J2_125_3477_U746 ( .A(DP_OP_423J2_125_3477_n1368), .B(
        DP_OP_423J2_125_3477_n1191), .CI(DP_OP_423J2_125_3477_n1366), .CO(
        DP_OP_423J2_125_3477_n1176), .S(DP_OP_423J2_125_3477_n1177) );
  FADDX1_HVT DP_OP_423J2_125_3477_U745 ( .A(DP_OP_423J2_125_3477_n1193), .B(
        DP_OP_423J2_125_3477_n1189), .CI(DP_OP_423J2_125_3477_n1187), .CO(
        DP_OP_423J2_125_3477_n1174), .S(DP_OP_423J2_125_3477_n1175) );
  FADDX1_HVT DP_OP_423J2_125_3477_U744 ( .A(DP_OP_423J2_125_3477_n1364), .B(
        DP_OP_423J2_125_3477_n1362), .CI(DP_OP_423J2_125_3477_n1185), .CO(
        DP_OP_423J2_125_3477_n1172), .S(DP_OP_423J2_125_3477_n1173) );
  FADDX1_HVT DP_OP_423J2_125_3477_U743 ( .A(DP_OP_423J2_125_3477_n1360), .B(
        DP_OP_423J2_125_3477_n1183), .CI(DP_OP_423J2_125_3477_n1181), .CO(
        DP_OP_423J2_125_3477_n1170), .S(DP_OP_423J2_125_3477_n1171) );
  FADDX1_HVT DP_OP_423J2_125_3477_U742 ( .A(DP_OP_423J2_125_3477_n1179), .B(
        DP_OP_423J2_125_3477_n1358), .CI(DP_OP_423J2_125_3477_n1177), .CO(
        DP_OP_423J2_125_3477_n1168), .S(DP_OP_423J2_125_3477_n1169) );
  FADDX1_HVT DP_OP_423J2_125_3477_U741 ( .A(DP_OP_423J2_125_3477_n1356), .B(
        DP_OP_423J2_125_3477_n1175), .CI(DP_OP_423J2_125_3477_n1354), .CO(
        DP_OP_423J2_125_3477_n1166), .S(DP_OP_423J2_125_3477_n1167) );
  FADDX1_HVT DP_OP_423J2_125_3477_U740 ( .A(DP_OP_423J2_125_3477_n1173), .B(
        DP_OP_423J2_125_3477_n1171), .CI(DP_OP_423J2_125_3477_n1352), .CO(
        DP_OP_423J2_125_3477_n1164), .S(DP_OP_423J2_125_3477_n1165) );
  FADDX1_HVT DP_OP_423J2_125_3477_U739 ( .A(DP_OP_423J2_125_3477_n1169), .B(
        DP_OP_423J2_125_3477_n1350), .CI(DP_OP_423J2_125_3477_n1167), .CO(
        DP_OP_423J2_125_3477_n1162), .S(DP_OP_423J2_125_3477_n1163) );
  OR2X1_HVT DP_OP_423J2_125_3477_U738 ( .A1(DP_OP_423J2_125_3477_n2979), .A2(
        DP_OP_423J2_125_3477_n2452), .Y(DP_OP_423J2_125_3477_n1160) );
  FADDX1_HVT DP_OP_423J2_125_3477_U736 ( .A(DP_OP_423J2_125_3477_n2144), .B(
        DP_OP_423J2_125_3477_n1924), .CI(DP_OP_423J2_125_3477_n1880), .CO(
        DP_OP_423J2_125_3477_n1158), .S(DP_OP_423J2_125_3477_n1159) );
  FADDX1_HVT DP_OP_423J2_125_3477_U735 ( .A(DP_OP_423J2_125_3477_n2584), .B(
        DP_OP_423J2_125_3477_n2012), .CI(DP_OP_423J2_125_3477_n2364), .CO(
        DP_OP_423J2_125_3477_n1156), .S(DP_OP_423J2_125_3477_n1157) );
  FADDX1_HVT DP_OP_423J2_125_3477_U734 ( .A(DP_OP_423J2_125_3477_n2804), .B(
        DP_OP_423J2_125_3477_n2628), .CI(DP_OP_423J2_125_3477_n2188), .CO(
        DP_OP_423J2_125_3477_n1154), .S(DP_OP_423J2_125_3477_n1155) );
  FADDX1_HVT DP_OP_423J2_125_3477_U733 ( .A(DP_OP_423J2_125_3477_n2276), .B(
        DP_OP_423J2_125_3477_n2100), .CI(DP_OP_423J2_125_3477_n2848), .CO(
        DP_OP_423J2_125_3477_n1152), .S(DP_OP_423J2_125_3477_n1153) );
  FADDX1_HVT DP_OP_423J2_125_3477_U732 ( .A(DP_OP_423J2_125_3477_n2408), .B(
        DP_OP_423J2_125_3477_n2892), .CI(DP_OP_423J2_125_3477_n2672), .CO(
        DP_OP_423J2_125_3477_n1150), .S(DP_OP_423J2_125_3477_n1151) );
  FADDX1_HVT DP_OP_423J2_125_3477_U731 ( .A(DP_OP_423J2_125_3477_n2496), .B(
        DP_OP_423J2_125_3477_n2716), .CI(DP_OP_423J2_125_3477_n2540), .CO(
        DP_OP_423J2_125_3477_n1148), .S(DP_OP_423J2_125_3477_n1149) );
  FADDX1_HVT DP_OP_423J2_125_3477_U730 ( .A(DP_OP_423J2_125_3477_n2232), .B(
        DP_OP_423J2_125_3477_n2056), .CI(DP_OP_423J2_125_3477_n2936), .CO(
        DP_OP_423J2_125_3477_n1146), .S(DP_OP_423J2_125_3477_n1147) );
  FADDX1_HVT DP_OP_423J2_125_3477_U729 ( .A(DP_OP_423J2_125_3477_n2760), .B(
        DP_OP_423J2_125_3477_n1968), .CI(DP_OP_423J2_125_3477_n2320), .CO(
        DP_OP_423J2_125_3477_n1144), .S(DP_OP_423J2_125_3477_n1145) );
  FADDX1_HVT DP_OP_423J2_125_3477_U728 ( .A(DP_OP_423J2_125_3477_n2371), .B(
        DP_OP_423J2_125_3477_n2999), .CI(DP_OP_423J2_125_3477_n1931), .CO(
        DP_OP_423J2_125_3477_n1142), .S(DP_OP_423J2_125_3477_n1143) );
  FADDX1_HVT DP_OP_423J2_125_3477_U727 ( .A(DP_OP_423J2_125_3477_n2378), .B(
        DP_OP_423J2_125_3477_n2992), .CI(DP_OP_423J2_125_3477_n2985), .CO(
        DP_OP_423J2_125_3477_n1140), .S(DP_OP_423J2_125_3477_n1141) );
  FADDX1_HVT DP_OP_423J2_125_3477_U726 ( .A(DP_OP_423J2_125_3477_n2334), .B(
        DP_OP_423J2_125_3477_n2957), .CI(DP_OP_423J2_125_3477_n2950), .CO(
        DP_OP_423J2_125_3477_n1138), .S(DP_OP_423J2_125_3477_n1139) );
  FADDX1_HVT DP_OP_423J2_125_3477_U725 ( .A(DP_OP_423J2_125_3477_n2297), .B(
        DP_OP_423J2_125_3477_n2943), .CI(DP_OP_423J2_125_3477_n2913), .CO(
        DP_OP_423J2_125_3477_n1136), .S(DP_OP_423J2_125_3477_n1137) );
  FADDX1_HVT DP_OP_423J2_125_3477_U724 ( .A(DP_OP_423J2_125_3477_n2290), .B(
        DP_OP_423J2_125_3477_n1938), .CI(DP_OP_423J2_125_3477_n2906), .CO(
        DP_OP_423J2_125_3477_n1134), .S(DP_OP_423J2_125_3477_n1135) );
  FADDX1_HVT DP_OP_423J2_125_3477_U723 ( .A(DP_OP_423J2_125_3477_n2327), .B(
        DP_OP_423J2_125_3477_n2899), .CI(DP_OP_423J2_125_3477_n1945), .CO(
        DP_OP_423J2_125_3477_n1132), .S(DP_OP_423J2_125_3477_n1133) );
  FADDX1_HVT DP_OP_423J2_125_3477_U722 ( .A(DP_OP_423J2_125_3477_n2283), .B(
        DP_OP_423J2_125_3477_n2869), .CI(DP_OP_423J2_125_3477_n1975), .CO(
        DP_OP_423J2_125_3477_n1130), .S(DP_OP_423J2_125_3477_n1131) );
  FADDX1_HVT DP_OP_423J2_125_3477_U721 ( .A(DP_OP_423J2_125_3477_n2253), .B(
        DP_OP_423J2_125_3477_n2862), .CI(DP_OP_423J2_125_3477_n2855), .CO(
        DP_OP_423J2_125_3477_n1128), .S(DP_OP_423J2_125_3477_n1129) );
  FADDX1_HVT DP_OP_423J2_125_3477_U720 ( .A(DP_OP_423J2_125_3477_n2246), .B(
        DP_OP_423J2_125_3477_n1982), .CI(DP_OP_423J2_125_3477_n2825), .CO(
        DP_OP_423J2_125_3477_n1126), .S(DP_OP_423J2_125_3477_n1127) );
  FADDX1_HVT DP_OP_423J2_125_3477_U719 ( .A(DP_OP_423J2_125_3477_n2239), .B(
        DP_OP_423J2_125_3477_n1989), .CI(DP_OP_423J2_125_3477_n2818), .CO(
        DP_OP_423J2_125_3477_n1124), .S(DP_OP_423J2_125_3477_n1125) );
  FADDX1_HVT DP_OP_423J2_125_3477_U718 ( .A(DP_OP_423J2_125_3477_n2019), .B(
        DP_OP_423J2_125_3477_n2026), .CI(DP_OP_423J2_125_3477_n2033), .CO(
        DP_OP_423J2_125_3477_n1122), .S(DP_OP_423J2_125_3477_n1123) );
  FADDX1_HVT DP_OP_423J2_125_3477_U717 ( .A(DP_OP_423J2_125_3477_n2811), .B(
        DP_OP_423J2_125_3477_n2063), .CI(DP_OP_423J2_125_3477_n2070), .CO(
        DP_OP_423J2_125_3477_n1120), .S(DP_OP_423J2_125_3477_n1121) );
  FADDX1_HVT DP_OP_423J2_125_3477_U716 ( .A(DP_OP_423J2_125_3477_n2781), .B(
        DP_OP_423J2_125_3477_n2077), .CI(DP_OP_423J2_125_3477_n2107), .CO(
        DP_OP_423J2_125_3477_n1118), .S(DP_OP_423J2_125_3477_n1119) );
  FADDX1_HVT DP_OP_423J2_125_3477_U715 ( .A(DP_OP_423J2_125_3477_n2774), .B(
        DP_OP_423J2_125_3477_n2114), .CI(DP_OP_423J2_125_3477_n2121), .CO(
        DP_OP_423J2_125_3477_n1116), .S(DP_OP_423J2_125_3477_n1117) );
  FADDX1_HVT DP_OP_423J2_125_3477_U714 ( .A(DP_OP_423J2_125_3477_n2767), .B(
        DP_OP_423J2_125_3477_n2151), .CI(DP_OP_423J2_125_3477_n2158), .CO(
        DP_OP_423J2_125_3477_n1114), .S(DP_OP_423J2_125_3477_n1115) );
  FADDX1_HVT DP_OP_423J2_125_3477_U713 ( .A(DP_OP_423J2_125_3477_n2737), .B(
        DP_OP_423J2_125_3477_n2165), .CI(DP_OP_423J2_125_3477_n2195), .CO(
        DP_OP_423J2_125_3477_n1112), .S(DP_OP_423J2_125_3477_n1113) );
  FADDX1_HVT DP_OP_423J2_125_3477_U712 ( .A(DP_OP_423J2_125_3477_n2730), .B(
        DP_OP_423J2_125_3477_n2202), .CI(DP_OP_423J2_125_3477_n2209), .CO(
        DP_OP_423J2_125_3477_n1110), .S(DP_OP_423J2_125_3477_n1111) );
  FADDX1_HVT DP_OP_423J2_125_3477_U711 ( .A(DP_OP_423J2_125_3477_n2723), .B(
        DP_OP_423J2_125_3477_n2341), .CI(DP_OP_423J2_125_3477_n2385), .CO(
        DP_OP_423J2_125_3477_n1108), .S(DP_OP_423J2_125_3477_n1109) );
  FADDX1_HVT DP_OP_423J2_125_3477_U710 ( .A(DP_OP_423J2_125_3477_n2693), .B(
        DP_OP_423J2_125_3477_n2415), .CI(DP_OP_423J2_125_3477_n2422), .CO(
        DP_OP_423J2_125_3477_n1106), .S(DP_OP_423J2_125_3477_n1107) );
  FADDX1_HVT DP_OP_423J2_125_3477_U709 ( .A(DP_OP_423J2_125_3477_n2686), .B(
        DP_OP_423J2_125_3477_n2429), .CI(DP_OP_423J2_125_3477_n2459), .CO(
        DP_OP_423J2_125_3477_n1104), .S(DP_OP_423J2_125_3477_n1105) );
  FADDX1_HVT DP_OP_423J2_125_3477_U708 ( .A(DP_OP_423J2_125_3477_n2679), .B(
        DP_OP_423J2_125_3477_n2466), .CI(DP_OP_423J2_125_3477_n2473), .CO(
        DP_OP_423J2_125_3477_n1102), .S(DP_OP_423J2_125_3477_n1103) );
  FADDX1_HVT DP_OP_423J2_125_3477_U707 ( .A(DP_OP_423J2_125_3477_n2649), .B(
        DP_OP_423J2_125_3477_n2503), .CI(DP_OP_423J2_125_3477_n2510), .CO(
        DP_OP_423J2_125_3477_n1100), .S(DP_OP_423J2_125_3477_n1101) );
  FADDX1_HVT DP_OP_423J2_125_3477_U706 ( .A(DP_OP_423J2_125_3477_n2642), .B(
        DP_OP_423J2_125_3477_n2517), .CI(DP_OP_423J2_125_3477_n2547), .CO(
        DP_OP_423J2_125_3477_n1098), .S(DP_OP_423J2_125_3477_n1099) );
  FADDX1_HVT DP_OP_423J2_125_3477_U705 ( .A(DP_OP_423J2_125_3477_n2635), .B(
        DP_OP_423J2_125_3477_n2554), .CI(DP_OP_423J2_125_3477_n2561), .CO(
        DP_OP_423J2_125_3477_n1096), .S(DP_OP_423J2_125_3477_n1097) );
  FADDX1_HVT DP_OP_423J2_125_3477_U704 ( .A(DP_OP_423J2_125_3477_n2591), .B(
        DP_OP_423J2_125_3477_n2598), .CI(DP_OP_423J2_125_3477_n2605), .CO(
        DP_OP_423J2_125_3477_n1094), .S(DP_OP_423J2_125_3477_n1095) );
  FADDX1_HVT DP_OP_423J2_125_3477_U703 ( .A(DP_OP_423J2_125_3477_n1348), .B(
        DP_OP_423J2_125_3477_n1336), .CI(DP_OP_423J2_125_3477_n1334), .CO(
        DP_OP_423J2_125_3477_n1092), .S(DP_OP_423J2_125_3477_n1093) );
  FADDX1_HVT DP_OP_423J2_125_3477_U702 ( .A(DP_OP_423J2_125_3477_n1332), .B(
        DP_OP_423J2_125_3477_n1338), .CI(DP_OP_423J2_125_3477_n1161), .CO(
        DP_OP_423J2_125_3477_n1090), .S(DP_OP_423J2_125_3477_n1091) );
  FADDX1_HVT DP_OP_423J2_125_3477_U701 ( .A(DP_OP_423J2_125_3477_n1342), .B(
        DP_OP_423J2_125_3477_n1346), .CI(DP_OP_423J2_125_3477_n1340), .CO(
        DP_OP_423J2_125_3477_n1088), .S(DP_OP_423J2_125_3477_n1089) );
  FADDX1_HVT DP_OP_423J2_125_3477_U700 ( .A(DP_OP_423J2_125_3477_n1344), .B(
        DP_OP_423J2_125_3477_n1308), .CI(DP_OP_423J2_125_3477_n1306), .CO(
        DP_OP_423J2_125_3477_n1086), .S(DP_OP_423J2_125_3477_n1087) );
  FADDX1_HVT DP_OP_423J2_125_3477_U699 ( .A(DP_OP_423J2_125_3477_n1310), .B(
        DP_OP_423J2_125_3477_n1282), .CI(DP_OP_423J2_125_3477_n1330), .CO(
        DP_OP_423J2_125_3477_n1084), .S(DP_OP_423J2_125_3477_n1085) );
  FADDX1_HVT DP_OP_423J2_125_3477_U698 ( .A(DP_OP_423J2_125_3477_n1302), .B(
        DP_OP_423J2_125_3477_n1284), .CI(DP_OP_423J2_125_3477_n1328), .CO(
        DP_OP_423J2_125_3477_n1082), .S(DP_OP_423J2_125_3477_n1083) );
  FADDX1_HVT DP_OP_423J2_125_3477_U697 ( .A(DP_OP_423J2_125_3477_n1300), .B(
        DP_OP_423J2_125_3477_n1286), .CI(DP_OP_423J2_125_3477_n1326), .CO(
        DP_OP_423J2_125_3477_n1080), .S(DP_OP_423J2_125_3477_n1081) );
  FADDX1_HVT DP_OP_423J2_125_3477_U696 ( .A(DP_OP_423J2_125_3477_n1296), .B(
        DP_OP_423J2_125_3477_n1324), .CI(DP_OP_423J2_125_3477_n1322), .CO(
        DP_OP_423J2_125_3477_n1078), .S(DP_OP_423J2_125_3477_n1079) );
  FADDX1_HVT DP_OP_423J2_125_3477_U695 ( .A(DP_OP_423J2_125_3477_n1290), .B(
        DP_OP_423J2_125_3477_n1320), .CI(DP_OP_423J2_125_3477_n1318), .CO(
        DP_OP_423J2_125_3477_n1076), .S(DP_OP_423J2_125_3477_n1077) );
  FADDX1_HVT DP_OP_423J2_125_3477_U694 ( .A(DP_OP_423J2_125_3477_n1298), .B(
        DP_OP_423J2_125_3477_n1316), .CI(DP_OP_423J2_125_3477_n1314), .CO(
        DP_OP_423J2_125_3477_n1074), .S(DP_OP_423J2_125_3477_n1075) );
  FADDX1_HVT DP_OP_423J2_125_3477_U693 ( .A(DP_OP_423J2_125_3477_n1292), .B(
        DP_OP_423J2_125_3477_n1312), .CI(DP_OP_423J2_125_3477_n1304), .CO(
        DP_OP_423J2_125_3477_n1072), .S(DP_OP_423J2_125_3477_n1073) );
  FADDX1_HVT DP_OP_423J2_125_3477_U692 ( .A(DP_OP_423J2_125_3477_n1294), .B(
        DP_OP_423J2_125_3477_n1288), .CI(DP_OP_423J2_125_3477_n1151), .CO(
        DP_OP_423J2_125_3477_n1070), .S(DP_OP_423J2_125_3477_n1071) );
  FADDX1_HVT DP_OP_423J2_125_3477_U691 ( .A(DP_OP_423J2_125_3477_n1147), .B(
        DP_OP_423J2_125_3477_n1145), .CI(DP_OP_423J2_125_3477_n1149), .CO(
        DP_OP_423J2_125_3477_n1068), .S(DP_OP_423J2_125_3477_n1069) );
  FADDX1_HVT DP_OP_423J2_125_3477_U690 ( .A(DP_OP_423J2_125_3477_n1157), .B(
        DP_OP_423J2_125_3477_n1155), .CI(DP_OP_423J2_125_3477_n1159), .CO(
        DP_OP_423J2_125_3477_n1066), .S(DP_OP_423J2_125_3477_n1067) );
  FADDX1_HVT DP_OP_423J2_125_3477_U689 ( .A(DP_OP_423J2_125_3477_n1153), .B(
        DP_OP_423J2_125_3477_n1101), .CI(DP_OP_423J2_125_3477_n1103), .CO(
        DP_OP_423J2_125_3477_n1064), .S(DP_OP_423J2_125_3477_n1065) );
  FADDX1_HVT DP_OP_423J2_125_3477_U688 ( .A(DP_OP_423J2_125_3477_n1099), .B(
        DP_OP_423J2_125_3477_n1135), .CI(DP_OP_423J2_125_3477_n1131), .CO(
        DP_OP_423J2_125_3477_n1062), .S(DP_OP_423J2_125_3477_n1063) );
  FADDX1_HVT DP_OP_423J2_125_3477_U687 ( .A(DP_OP_423J2_125_3477_n1137), .B(
        DP_OP_423J2_125_3477_n1121), .CI(DP_OP_423J2_125_3477_n1127), .CO(
        DP_OP_423J2_125_3477_n1060), .S(DP_OP_423J2_125_3477_n1061) );
  FADDX1_HVT DP_OP_423J2_125_3477_U686 ( .A(DP_OP_423J2_125_3477_n1125), .B(
        DP_OP_423J2_125_3477_n1123), .CI(DP_OP_423J2_125_3477_n1107), .CO(
        DP_OP_423J2_125_3477_n1058), .S(DP_OP_423J2_125_3477_n1059) );
  FADDX1_HVT DP_OP_423J2_125_3477_U685 ( .A(DP_OP_423J2_125_3477_n1129), .B(
        DP_OP_423J2_125_3477_n1097), .CI(DP_OP_423J2_125_3477_n1095), .CO(
        DP_OP_423J2_125_3477_n1056), .S(DP_OP_423J2_125_3477_n1057) );
  FADDX1_HVT DP_OP_423J2_125_3477_U684 ( .A(DP_OP_423J2_125_3477_n1133), .B(
        DP_OP_423J2_125_3477_n1115), .CI(DP_OP_423J2_125_3477_n1117), .CO(
        DP_OP_423J2_125_3477_n1054), .S(DP_OP_423J2_125_3477_n1055) );
  FADDX1_HVT DP_OP_423J2_125_3477_U683 ( .A(DP_OP_423J2_125_3477_n1113), .B(
        DP_OP_423J2_125_3477_n1111), .CI(DP_OP_423J2_125_3477_n1105), .CO(
        DP_OP_423J2_125_3477_n1052), .S(DP_OP_423J2_125_3477_n1053) );
  FADDX1_HVT DP_OP_423J2_125_3477_U682 ( .A(DP_OP_423J2_125_3477_n1109), .B(
        DP_OP_423J2_125_3477_n1143), .CI(DP_OP_423J2_125_3477_n1141), .CO(
        DP_OP_423J2_125_3477_n1050), .S(DP_OP_423J2_125_3477_n1051) );
  FADDX1_HVT DP_OP_423J2_125_3477_U681 ( .A(DP_OP_423J2_125_3477_n1139), .B(
        DP_OP_423J2_125_3477_n1119), .CI(DP_OP_423J2_125_3477_n1280), .CO(
        DP_OP_423J2_125_3477_n1048), .S(DP_OP_423J2_125_3477_n1049) );
  FADDX1_HVT DP_OP_423J2_125_3477_U680 ( .A(DP_OP_423J2_125_3477_n1278), .B(
        DP_OP_423J2_125_3477_n1276), .CI(DP_OP_423J2_125_3477_n1274), .CO(
        DP_OP_423J2_125_3477_n1046), .S(DP_OP_423J2_125_3477_n1047) );
  FADDX1_HVT DP_OP_423J2_125_3477_U679 ( .A(DP_OP_423J2_125_3477_n1272), .B(
        DP_OP_423J2_125_3477_n1260), .CI(DP_OP_423J2_125_3477_n1258), .CO(
        DP_OP_423J2_125_3477_n1044), .S(DP_OP_423J2_125_3477_n1045) );
  FADDX1_HVT DP_OP_423J2_125_3477_U678 ( .A(DP_OP_423J2_125_3477_n1264), .B(
        DP_OP_423J2_125_3477_n1262), .CI(DP_OP_423J2_125_3477_n1270), .CO(
        DP_OP_423J2_125_3477_n1042), .S(DP_OP_423J2_125_3477_n1043) );
  FADDX1_HVT DP_OP_423J2_125_3477_U677 ( .A(DP_OP_423J2_125_3477_n1268), .B(
        DP_OP_423J2_125_3477_n1266), .CI(DP_OP_423J2_125_3477_n1093), .CO(
        DP_OP_423J2_125_3477_n1040), .S(DP_OP_423J2_125_3477_n1041) );
  FADDX1_HVT DP_OP_423J2_125_3477_U676 ( .A(DP_OP_423J2_125_3477_n1256), .B(
        DP_OP_423J2_125_3477_n1254), .CI(DP_OP_423J2_125_3477_n1087), .CO(
        DP_OP_423J2_125_3477_n1038), .S(DP_OP_423J2_125_3477_n1039) );
  FADDX1_HVT DP_OP_423J2_125_3477_U675 ( .A(DP_OP_423J2_125_3477_n1091), .B(
        DP_OP_423J2_125_3477_n1089), .CI(DP_OP_423J2_125_3477_n1252), .CO(
        DP_OP_423J2_125_3477_n1036), .S(DP_OP_423J2_125_3477_n1037) );
  FADDX1_HVT DP_OP_423J2_125_3477_U674 ( .A(DP_OP_423J2_125_3477_n1240), .B(
        DP_OP_423J2_125_3477_n1085), .CI(DP_OP_423J2_125_3477_n1071), .CO(
        DP_OP_423J2_125_3477_n1034), .S(DP_OP_423J2_125_3477_n1035) );
  FADDX1_HVT DP_OP_423J2_125_3477_U673 ( .A(DP_OP_423J2_125_3477_n1238), .B(
        DP_OP_423J2_125_3477_n1081), .CI(DP_OP_423J2_125_3477_n1083), .CO(
        DP_OP_423J2_125_3477_n1032), .S(DP_OP_423J2_125_3477_n1033) );
  FADDX1_HVT DP_OP_423J2_125_3477_U672 ( .A(DP_OP_423J2_125_3477_n1242), .B(
        DP_OP_423J2_125_3477_n1079), .CI(DP_OP_423J2_125_3477_n1077), .CO(
        DP_OP_423J2_125_3477_n1030), .S(DP_OP_423J2_125_3477_n1031) );
  FADDX1_HVT DP_OP_423J2_125_3477_U671 ( .A(DP_OP_423J2_125_3477_n1250), .B(
        DP_OP_423J2_125_3477_n1073), .CI(DP_OP_423J2_125_3477_n1075), .CO(
        DP_OP_423J2_125_3477_n1028), .S(DP_OP_423J2_125_3477_n1029) );
  FADDX1_HVT DP_OP_423J2_125_3477_U670 ( .A(DP_OP_423J2_125_3477_n1248), .B(
        DP_OP_423J2_125_3477_n1244), .CI(DP_OP_423J2_125_3477_n1246), .CO(
        DP_OP_423J2_125_3477_n1026), .S(DP_OP_423J2_125_3477_n1027) );
  FADDX1_HVT DP_OP_423J2_125_3477_U669 ( .A(DP_OP_423J2_125_3477_n1067), .B(
        DP_OP_423J2_125_3477_n1236), .CI(DP_OP_423J2_125_3477_n1065), .CO(
        DP_OP_423J2_125_3477_n1024), .S(DP_OP_423J2_125_3477_n1025) );
  FADDX1_HVT DP_OP_423J2_125_3477_U668 ( .A(DP_OP_423J2_125_3477_n1069), .B(
        DP_OP_423J2_125_3477_n1059), .CI(DP_OP_423J2_125_3477_n1061), .CO(
        DP_OP_423J2_125_3477_n1022), .S(DP_OP_423J2_125_3477_n1023) );
  FADDX1_HVT DP_OP_423J2_125_3477_U667 ( .A(DP_OP_423J2_125_3477_n1057), .B(
        DP_OP_423J2_125_3477_n1051), .CI(DP_OP_423J2_125_3477_n1234), .CO(
        DP_OP_423J2_125_3477_n1020), .S(DP_OP_423J2_125_3477_n1021) );
  FADDX1_HVT DP_OP_423J2_125_3477_U666 ( .A(DP_OP_423J2_125_3477_n1053), .B(
        DP_OP_423J2_125_3477_n1063), .CI(DP_OP_423J2_125_3477_n1055), .CO(
        DP_OP_423J2_125_3477_n1018), .S(DP_OP_423J2_125_3477_n1019) );
  FADDX1_HVT DP_OP_423J2_125_3477_U665 ( .A(DP_OP_423J2_125_3477_n1049), .B(
        DP_OP_423J2_125_3477_n1232), .CI(DP_OP_423J2_125_3477_n1228), .CO(
        DP_OP_423J2_125_3477_n1016), .S(DP_OP_423J2_125_3477_n1017) );
  FADDX1_HVT DP_OP_423J2_125_3477_U664 ( .A(DP_OP_423J2_125_3477_n1230), .B(
        DP_OP_423J2_125_3477_n1226), .CI(DP_OP_423J2_125_3477_n1224), .CO(
        DP_OP_423J2_125_3477_n1014), .S(DP_OP_423J2_125_3477_n1015) );
  FADDX1_HVT DP_OP_423J2_125_3477_U663 ( .A(DP_OP_423J2_125_3477_n1047), .B(
        DP_OP_423J2_125_3477_n1222), .CI(DP_OP_423J2_125_3477_n1220), .CO(
        DP_OP_423J2_125_3477_n1012), .S(DP_OP_423J2_125_3477_n1013) );
  FADDX1_HVT DP_OP_423J2_125_3477_U662 ( .A(DP_OP_423J2_125_3477_n1218), .B(
        DP_OP_423J2_125_3477_n1043), .CI(DP_OP_423J2_125_3477_n1041), .CO(
        DP_OP_423J2_125_3477_n1010), .S(DP_OP_423J2_125_3477_n1011) );
  FADDX1_HVT DP_OP_423J2_125_3477_U661 ( .A(DP_OP_423J2_125_3477_n1216), .B(
        DP_OP_423J2_125_3477_n1214), .CI(DP_OP_423J2_125_3477_n1045), .CO(
        DP_OP_423J2_125_3477_n1008), .S(DP_OP_423J2_125_3477_n1009) );
  FADDX1_HVT DP_OP_423J2_125_3477_U660 ( .A(DP_OP_423J2_125_3477_n1037), .B(
        DP_OP_423J2_125_3477_n1212), .CI(DP_OP_423J2_125_3477_n1039), .CO(
        DP_OP_423J2_125_3477_n1006), .S(DP_OP_423J2_125_3477_n1007) );
  FADDX1_HVT DP_OP_423J2_125_3477_U659 ( .A(DP_OP_423J2_125_3477_n1031), .B(
        DP_OP_423J2_125_3477_n1035), .CI(DP_OP_423J2_125_3477_n1206), .CO(
        DP_OP_423J2_125_3477_n1004), .S(DP_OP_423J2_125_3477_n1005) );
  FADDX1_HVT DP_OP_423J2_125_3477_U658 ( .A(DP_OP_423J2_125_3477_n1210), .B(
        DP_OP_423J2_125_3477_n1029), .CI(DP_OP_423J2_125_3477_n1033), .CO(
        DP_OP_423J2_125_3477_n1002), .S(DP_OP_423J2_125_3477_n1003) );
  FADDX1_HVT DP_OP_423J2_125_3477_U657 ( .A(DP_OP_423J2_125_3477_n1208), .B(
        DP_OP_423J2_125_3477_n1027), .CI(DP_OP_423J2_125_3477_n1204), .CO(
        DP_OP_423J2_125_3477_n1000), .S(DP_OP_423J2_125_3477_n1001) );
  FADDX1_HVT DP_OP_423J2_125_3477_U656 ( .A(DP_OP_423J2_125_3477_n1025), .B(
        DP_OP_423J2_125_3477_n1023), .CI(DP_OP_423J2_125_3477_n1021), .CO(
        DP_OP_423J2_125_3477_n998), .S(DP_OP_423J2_125_3477_n999) );
  FADDX1_HVT DP_OP_423J2_125_3477_U655 ( .A(DP_OP_423J2_125_3477_n1019), .B(
        DP_OP_423J2_125_3477_n1202), .CI(DP_OP_423J2_125_3477_n1017), .CO(
        DP_OP_423J2_125_3477_n996), .S(DP_OP_423J2_125_3477_n997) );
  FADDX1_HVT DP_OP_423J2_125_3477_U654 ( .A(DP_OP_423J2_125_3477_n1200), .B(
        DP_OP_423J2_125_3477_n1198), .CI(DP_OP_423J2_125_3477_n1196), .CO(
        DP_OP_423J2_125_3477_n994), .S(DP_OP_423J2_125_3477_n995) );
  FADDX1_HVT DP_OP_423J2_125_3477_U653 ( .A(DP_OP_423J2_125_3477_n1015), .B(
        DP_OP_423J2_125_3477_n1194), .CI(DP_OP_423J2_125_3477_n1013), .CO(
        DP_OP_423J2_125_3477_n992), .S(DP_OP_423J2_125_3477_n993) );
  FADDX1_HVT DP_OP_423J2_125_3477_U652 ( .A(DP_OP_423J2_125_3477_n1192), .B(
        DP_OP_423J2_125_3477_n1009), .CI(DP_OP_423J2_125_3477_n1011), .CO(
        DP_OP_423J2_125_3477_n990), .S(DP_OP_423J2_125_3477_n991) );
  FADDX1_HVT DP_OP_423J2_125_3477_U651 ( .A(DP_OP_423J2_125_3477_n1190), .B(
        DP_OP_423J2_125_3477_n1188), .CI(DP_OP_423J2_125_3477_n1007), .CO(
        DP_OP_423J2_125_3477_n988), .S(DP_OP_423J2_125_3477_n989) );
  FADDX1_HVT DP_OP_423J2_125_3477_U650 ( .A(DP_OP_423J2_125_3477_n1186), .B(
        DP_OP_423J2_125_3477_n1003), .CI(DP_OP_423J2_125_3477_n1001), .CO(
        DP_OP_423J2_125_3477_n986), .S(DP_OP_423J2_125_3477_n987) );
  FADDX1_HVT DP_OP_423J2_125_3477_U649 ( .A(DP_OP_423J2_125_3477_n1005), .B(
        DP_OP_423J2_125_3477_n1184), .CI(DP_OP_423J2_125_3477_n999), .CO(
        DP_OP_423J2_125_3477_n984), .S(DP_OP_423J2_125_3477_n985) );
  FADDX1_HVT DP_OP_423J2_125_3477_U648 ( .A(DP_OP_423J2_125_3477_n1182), .B(
        DP_OP_423J2_125_3477_n997), .CI(DP_OP_423J2_125_3477_n1180), .CO(
        DP_OP_423J2_125_3477_n982), .S(DP_OP_423J2_125_3477_n983) );
  FADDX1_HVT DP_OP_423J2_125_3477_U647 ( .A(DP_OP_423J2_125_3477_n995), .B(
        DP_OP_423J2_125_3477_n1178), .CI(DP_OP_423J2_125_3477_n993), .CO(
        DP_OP_423J2_125_3477_n980), .S(DP_OP_423J2_125_3477_n981) );
  FADDX1_HVT DP_OP_423J2_125_3477_U646 ( .A(DP_OP_423J2_125_3477_n1176), .B(
        DP_OP_423J2_125_3477_n991), .CI(DP_OP_423J2_125_3477_n989), .CO(
        DP_OP_423J2_125_3477_n978), .S(DP_OP_423J2_125_3477_n979) );
  FADDX1_HVT DP_OP_423J2_125_3477_U645 ( .A(DP_OP_423J2_125_3477_n1174), .B(
        DP_OP_423J2_125_3477_n987), .CI(DP_OP_423J2_125_3477_n1172), .CO(
        DP_OP_423J2_125_3477_n976), .S(DP_OP_423J2_125_3477_n977) );
  FADDX1_HVT DP_OP_423J2_125_3477_U644 ( .A(DP_OP_423J2_125_3477_n985), .B(
        DP_OP_423J2_125_3477_n1170), .CI(DP_OP_423J2_125_3477_n983), .CO(
        DP_OP_423J2_125_3477_n974), .S(DP_OP_423J2_125_3477_n975) );
  FADDX1_HVT DP_OP_423J2_125_3477_U643 ( .A(DP_OP_423J2_125_3477_n981), .B(
        DP_OP_423J2_125_3477_n1168), .CI(DP_OP_423J2_125_3477_n979), .CO(
        DP_OP_423J2_125_3477_n972), .S(DP_OP_423J2_125_3477_n973) );
  FADDX1_HVT DP_OP_423J2_125_3477_U642 ( .A(DP_OP_423J2_125_3477_n1166), .B(
        DP_OP_423J2_125_3477_n977), .CI(DP_OP_423J2_125_3477_n975), .CO(
        DP_OP_423J2_125_3477_n970), .S(DP_OP_423J2_125_3477_n971) );
  FADDX1_HVT DP_OP_423J2_125_3477_U641 ( .A(DP_OP_423J2_125_3477_n1164), .B(
        DP_OP_423J2_125_3477_n973), .CI(DP_OP_423J2_125_3477_n1162), .CO(
        DP_OP_423J2_125_3477_n968), .S(DP_OP_423J2_125_3477_n969) );
  FADDX1_HVT DP_OP_423J2_125_3477_U640 ( .A(DP_OP_423J2_125_3477_n2978), .B(
        DP_OP_423J2_125_3477_n1923), .CI(DP_OP_423J2_125_3477_n1879), .CO(
        DP_OP_423J2_125_3477_n966), .S(DP_OP_423J2_125_3477_n967) );
  FADDX1_HVT DP_OP_423J2_125_3477_U639 ( .A(DP_OP_423J2_125_3477_n2803), .B(
        DP_OP_423J2_125_3477_n2120), .CI(DP_OP_423J2_125_3477_n2384), .CO(
        DP_OP_423J2_125_3477_n964), .S(DP_OP_423J2_125_3477_n965) );
  FADDX1_HVT DP_OP_423J2_125_3477_U638 ( .A(DP_OP_423J2_125_3477_n2011), .B(
        DP_OP_423J2_125_3477_n2428), .CI(DP_OP_423J2_125_3477_n1988), .CO(
        DP_OP_423J2_125_3477_n962), .S(DP_OP_423J2_125_3477_n963) );
  FADDX1_HVT DP_OP_423J2_125_3477_U637 ( .A(DP_OP_423J2_125_3477_n2319), .B(
        DP_OP_423J2_125_3477_n1944), .CI(DP_OP_423J2_125_3477_n2912), .CO(
        DP_OP_423J2_125_3477_n960), .S(DP_OP_423J2_125_3477_n961) );
  FADDX1_HVT DP_OP_423J2_125_3477_U636 ( .A(DP_OP_423J2_125_3477_n2275), .B(
        DP_OP_423J2_125_3477_n2252), .CI(DP_OP_423J2_125_3477_n2604), .CO(
        DP_OP_423J2_125_3477_n958), .S(DP_OP_423J2_125_3477_n959) );
  FADDX1_HVT DP_OP_423J2_125_3477_U635 ( .A(DP_OP_423J2_125_3477_n2187), .B(
        DP_OP_423J2_125_3477_n2296), .CI(DP_OP_423J2_125_3477_n2956), .CO(
        DP_OP_423J2_125_3477_n956), .S(DP_OP_423J2_125_3477_n957) );
  FADDX1_HVT DP_OP_423J2_125_3477_U634 ( .A(DP_OP_423J2_125_3477_n1967), .B(
        DP_OP_423J2_125_3477_n2032), .CI(DP_OP_423J2_125_3477_n2472), .CO(
        DP_OP_423J2_125_3477_n954), .S(DP_OP_423J2_125_3477_n955) );
  FADDX1_HVT DP_OP_423J2_125_3477_U633 ( .A(DP_OP_423J2_125_3477_n2055), .B(
        DP_OP_423J2_125_3477_n2736), .CI(DP_OP_423J2_125_3477_n2780), .CO(
        DP_OP_423J2_125_3477_n952), .S(DP_OP_423J2_125_3477_n953) );
  FADDX1_HVT DP_OP_423J2_125_3477_U632 ( .A(DP_OP_423J2_125_3477_n2143), .B(
        DP_OP_423J2_125_3477_n2692), .CI(DP_OP_423J2_125_3477_n2560), .CO(
        DP_OP_423J2_125_3477_n950), .S(DP_OP_423J2_125_3477_n951) );
  FADDX1_HVT DP_OP_423J2_125_3477_U631 ( .A(DP_OP_423J2_125_3477_n2495), .B(
        DP_OP_423J2_125_3477_n2340), .CI(DP_OP_423J2_125_3477_n2824), .CO(
        DP_OP_423J2_125_3477_n948), .S(DP_OP_423J2_125_3477_n949) );
  FADDX1_HVT DP_OP_423J2_125_3477_U630 ( .A(DP_OP_423J2_125_3477_n2891), .B(
        DP_OP_423J2_125_3477_n2164), .CI(DP_OP_423J2_125_3477_n2076), .CO(
        DP_OP_423J2_125_3477_n946), .S(DP_OP_423J2_125_3477_n947) );
  FADDX1_HVT DP_OP_423J2_125_3477_U629 ( .A(DP_OP_423J2_125_3477_n2627), .B(
        DP_OP_423J2_125_3477_n2868), .CI(DP_OP_423J2_125_3477_n2516), .CO(
        DP_OP_423J2_125_3477_n944), .S(DP_OP_423J2_125_3477_n945) );
  FADDX1_HVT DP_OP_423J2_125_3477_U628 ( .A(DP_OP_423J2_125_3477_n2407), .B(
        DP_OP_423J2_125_3477_n2998), .CI(DP_OP_423J2_125_3477_n2208), .CO(
        DP_OP_423J2_125_3477_n942), .S(DP_OP_423J2_125_3477_n943) );
  FADDX1_HVT DP_OP_423J2_125_3477_U627 ( .A(DP_OP_423J2_125_3477_n2099), .B(
        DP_OP_423J2_125_3477_n2363), .CI(DP_OP_423J2_125_3477_n2648), .CO(
        DP_OP_423J2_125_3477_n940), .S(DP_OP_423J2_125_3477_n941) );
  FADDX1_HVT DP_OP_423J2_125_3477_U626 ( .A(DP_OP_423J2_125_3477_n2715), .B(
        DP_OP_423J2_125_3477_n2759), .CI(DP_OP_423J2_125_3477_n2847), .CO(
        DP_OP_423J2_125_3477_n938), .S(DP_OP_423J2_125_3477_n939) );
  FADDX1_HVT DP_OP_423J2_125_3477_U625 ( .A(DP_OP_423J2_125_3477_n2451), .B(
        DP_OP_423J2_125_3477_n2539), .CI(DP_OP_423J2_125_3477_n2935), .CO(
        DP_OP_423J2_125_3477_n936), .S(DP_OP_423J2_125_3477_n937) );
  FADDX1_HVT DP_OP_423J2_125_3477_U624 ( .A(DP_OP_423J2_125_3477_n2583), .B(
        DP_OP_423J2_125_3477_n2231), .CI(DP_OP_423J2_125_3477_n2671), .CO(
        DP_OP_423J2_125_3477_n934), .S(DP_OP_423J2_125_3477_n935) );
  FADDX1_HVT DP_OP_423J2_125_3477_U623 ( .A(DP_OP_423J2_125_3477_n2991), .B(
        DP_OP_423J2_125_3477_n1937), .CI(DP_OP_423J2_125_3477_n1930), .CO(
        DP_OP_423J2_125_3477_n932), .S(DP_OP_423J2_125_3477_n933) );
  FADDX1_HVT DP_OP_423J2_125_3477_U622 ( .A(DP_OP_423J2_125_3477_n2984), .B(
        DP_OP_423J2_125_3477_n2949), .CI(DP_OP_423J2_125_3477_n2942), .CO(
        DP_OP_423J2_125_3477_n930), .S(DP_OP_423J2_125_3477_n931) );
  FADDX1_HVT DP_OP_423J2_125_3477_U621 ( .A(DP_OP_423J2_125_3477_n2465), .B(
        DP_OP_423J2_125_3477_n2905), .CI(DP_OP_423J2_125_3477_n2898), .CO(
        DP_OP_423J2_125_3477_n928), .S(DP_OP_423J2_125_3477_n929) );
  FADDX1_HVT DP_OP_423J2_125_3477_U620 ( .A(DP_OP_423J2_125_3477_n2861), .B(
        DP_OP_423J2_125_3477_n1974), .CI(DP_OP_423J2_125_3477_n1981), .CO(
        DP_OP_423J2_125_3477_n926), .S(DP_OP_423J2_125_3477_n927) );
  FADDX1_HVT DP_OP_423J2_125_3477_U619 ( .A(DP_OP_423J2_125_3477_n2854), .B(
        DP_OP_423J2_125_3477_n2018), .CI(DP_OP_423J2_125_3477_n2025), .CO(
        DP_OP_423J2_125_3477_n924), .S(DP_OP_423J2_125_3477_n925) );
  FADDX1_HVT DP_OP_423J2_125_3477_U618 ( .A(DP_OP_423J2_125_3477_n2817), .B(
        DP_OP_423J2_125_3477_n2062), .CI(DP_OP_423J2_125_3477_n2069), .CO(
        DP_OP_423J2_125_3477_n922), .S(DP_OP_423J2_125_3477_n923) );
  FADDX1_HVT DP_OP_423J2_125_3477_U617 ( .A(DP_OP_423J2_125_3477_n2810), .B(
        DP_OP_423J2_125_3477_n2106), .CI(DP_OP_423J2_125_3477_n2113), .CO(
        DP_OP_423J2_125_3477_n920), .S(DP_OP_423J2_125_3477_n921) );
  FADDX1_HVT DP_OP_423J2_125_3477_U616 ( .A(DP_OP_423J2_125_3477_n2773), .B(
        DP_OP_423J2_125_3477_n2150), .CI(DP_OP_423J2_125_3477_n2157), .CO(
        DP_OP_423J2_125_3477_n918), .S(DP_OP_423J2_125_3477_n919) );
  FADDX1_HVT DP_OP_423J2_125_3477_U615 ( .A(DP_OP_423J2_125_3477_n2766), .B(
        DP_OP_423J2_125_3477_n2194), .CI(DP_OP_423J2_125_3477_n2201), .CO(
        DP_OP_423J2_125_3477_n916), .S(DP_OP_423J2_125_3477_n917) );
  FADDX1_HVT DP_OP_423J2_125_3477_U614 ( .A(DP_OP_423J2_125_3477_n2729), .B(
        DP_OP_423J2_125_3477_n2238), .CI(DP_OP_423J2_125_3477_n2245), .CO(
        DP_OP_423J2_125_3477_n914), .S(DP_OP_423J2_125_3477_n915) );
  FADDX1_HVT DP_OP_423J2_125_3477_U613 ( .A(DP_OP_423J2_125_3477_n2722), .B(
        DP_OP_423J2_125_3477_n2282), .CI(DP_OP_423J2_125_3477_n2289), .CO(
        DP_OP_423J2_125_3477_n912), .S(DP_OP_423J2_125_3477_n913) );
  FADDX1_HVT DP_OP_423J2_125_3477_U612 ( .A(DP_OP_423J2_125_3477_n2685), .B(
        DP_OP_423J2_125_3477_n2326), .CI(DP_OP_423J2_125_3477_n2333), .CO(
        DP_OP_423J2_125_3477_n910), .S(DP_OP_423J2_125_3477_n911) );
  FADDX1_HVT DP_OP_423J2_125_3477_U611 ( .A(DP_OP_423J2_125_3477_n2678), .B(
        DP_OP_423J2_125_3477_n2370), .CI(DP_OP_423J2_125_3477_n2377), .CO(
        DP_OP_423J2_125_3477_n908), .S(DP_OP_423J2_125_3477_n909) );
  FADDX1_HVT DP_OP_423J2_125_3477_U610 ( .A(DP_OP_423J2_125_3477_n2641), .B(
        DP_OP_423J2_125_3477_n2414), .CI(DP_OP_423J2_125_3477_n2421), .CO(
        DP_OP_423J2_125_3477_n906), .S(DP_OP_423J2_125_3477_n907) );
  FADDX1_HVT DP_OP_423J2_125_3477_U609 ( .A(DP_OP_423J2_125_3477_n2634), .B(
        DP_OP_423J2_125_3477_n2458), .CI(DP_OP_423J2_125_3477_n2502), .CO(
        DP_OP_423J2_125_3477_n904), .S(DP_OP_423J2_125_3477_n905) );
  FADDX1_HVT DP_OP_423J2_125_3477_U608 ( .A(DP_OP_423J2_125_3477_n2597), .B(
        DP_OP_423J2_125_3477_n2509), .CI(DP_OP_423J2_125_3477_n2546), .CO(
        DP_OP_423J2_125_3477_n902), .S(DP_OP_423J2_125_3477_n903) );
  FADDX1_HVT DP_OP_423J2_125_3477_U607 ( .A(DP_OP_423J2_125_3477_n2590), .B(
        DP_OP_423J2_125_3477_n2553), .CI(DP_OP_423J2_125_3477_n1160), .CO(
        DP_OP_423J2_125_3477_n900), .S(DP_OP_423J2_125_3477_n901) );
  FADDX1_HVT DP_OP_423J2_125_3477_U606 ( .A(DP_OP_423J2_125_3477_n1148), .B(
        DP_OP_423J2_125_3477_n1144), .CI(DP_OP_423J2_125_3477_n1158), .CO(
        DP_OP_423J2_125_3477_n898), .S(DP_OP_423J2_125_3477_n899) );
  FADDX1_HVT DP_OP_423J2_125_3477_U605 ( .A(DP_OP_423J2_125_3477_n1156), .B(
        DP_OP_423J2_125_3477_n1146), .CI(DP_OP_423J2_125_3477_n1154), .CO(
        DP_OP_423J2_125_3477_n896), .S(DP_OP_423J2_125_3477_n897) );
  FADDX1_HVT DP_OP_423J2_125_3477_U604 ( .A(DP_OP_423J2_125_3477_n1152), .B(
        DP_OP_423J2_125_3477_n1150), .CI(DP_OP_423J2_125_3477_n1120), .CO(
        DP_OP_423J2_125_3477_n894), .S(DP_OP_423J2_125_3477_n895) );
  FADDX1_HVT DP_OP_423J2_125_3477_U603 ( .A(DP_OP_423J2_125_3477_n1118), .B(
        DP_OP_423J2_125_3477_n1094), .CI(DP_OP_423J2_125_3477_n1142), .CO(
        DP_OP_423J2_125_3477_n892), .S(DP_OP_423J2_125_3477_n893) );
  FADDX1_HVT DP_OP_423J2_125_3477_U602 ( .A(DP_OP_423J2_125_3477_n1116), .B(
        DP_OP_423J2_125_3477_n1140), .CI(DP_OP_423J2_125_3477_n1138), .CO(
        DP_OP_423J2_125_3477_n890), .S(DP_OP_423J2_125_3477_n891) );
  FADDX1_HVT DP_OP_423J2_125_3477_U601 ( .A(DP_OP_423J2_125_3477_n1110), .B(
        DP_OP_423J2_125_3477_n1136), .CI(DP_OP_423J2_125_3477_n1134), .CO(
        DP_OP_423J2_125_3477_n888), .S(DP_OP_423J2_125_3477_n889) );
  FADDX1_HVT DP_OP_423J2_125_3477_U600 ( .A(DP_OP_423J2_125_3477_n1132), .B(
        DP_OP_423J2_125_3477_n1130), .CI(DP_OP_423J2_125_3477_n1128), .CO(
        DP_OP_423J2_125_3477_n886), .S(DP_OP_423J2_125_3477_n887) );
  FADDX1_HVT DP_OP_423J2_125_3477_U599 ( .A(DP_OP_423J2_125_3477_n1100), .B(
        DP_OP_423J2_125_3477_n1126), .CI(DP_OP_423J2_125_3477_n1124), .CO(
        DP_OP_423J2_125_3477_n884), .S(DP_OP_423J2_125_3477_n885) );
  FADDX1_HVT DP_OP_423J2_125_3477_U598 ( .A(DP_OP_423J2_125_3477_n1106), .B(
        DP_OP_423J2_125_3477_n1122), .CI(DP_OP_423J2_125_3477_n1114), .CO(
        DP_OP_423J2_125_3477_n882), .S(DP_OP_423J2_125_3477_n883) );
  FADDX1_HVT DP_OP_423J2_125_3477_U597 ( .A(DP_OP_423J2_125_3477_n1098), .B(
        DP_OP_423J2_125_3477_n1112), .CI(DP_OP_423J2_125_3477_n1108), .CO(
        DP_OP_423J2_125_3477_n880), .S(DP_OP_423J2_125_3477_n881) );
  FADDX1_HVT DP_OP_423J2_125_3477_U596 ( .A(DP_OP_423J2_125_3477_n1102), .B(
        DP_OP_423J2_125_3477_n1096), .CI(DP_OP_423J2_125_3477_n1104), .CO(
        DP_OP_423J2_125_3477_n878), .S(DP_OP_423J2_125_3477_n879) );
  FADDX1_HVT DP_OP_423J2_125_3477_U595 ( .A(DP_OP_423J2_125_3477_n967), .B(
        DP_OP_423J2_125_3477_n953), .CI(DP_OP_423J2_125_3477_n955), .CO(
        DP_OP_423J2_125_3477_n876), .S(DP_OP_423J2_125_3477_n877) );
  FADDX1_HVT DP_OP_423J2_125_3477_U594 ( .A(DP_OP_423J2_125_3477_n959), .B(
        DP_OP_423J2_125_3477_n937), .CI(DP_OP_423J2_125_3477_n935), .CO(
        DP_OP_423J2_125_3477_n874), .S(DP_OP_423J2_125_3477_n875) );
  FADDX1_HVT DP_OP_423J2_125_3477_U593 ( .A(DP_OP_423J2_125_3477_n951), .B(
        DP_OP_423J2_125_3477_n949), .CI(DP_OP_423J2_125_3477_n945), .CO(
        DP_OP_423J2_125_3477_n872), .S(DP_OP_423J2_125_3477_n873) );
  FADDX1_HVT DP_OP_423J2_125_3477_U592 ( .A(DP_OP_423J2_125_3477_n957), .B(
        DP_OP_423J2_125_3477_n939), .CI(DP_OP_423J2_125_3477_n943), .CO(
        DP_OP_423J2_125_3477_n870), .S(DP_OP_423J2_125_3477_n871) );
  FADDX1_HVT DP_OP_423J2_125_3477_U591 ( .A(DP_OP_423J2_125_3477_n947), .B(
        DP_OP_423J2_125_3477_n965), .CI(DP_OP_423J2_125_3477_n961), .CO(
        DP_OP_423J2_125_3477_n868), .S(DP_OP_423J2_125_3477_n869) );
  FADDX1_HVT DP_OP_423J2_125_3477_U590 ( .A(DP_OP_423J2_125_3477_n941), .B(
        DP_OP_423J2_125_3477_n963), .CI(DP_OP_423J2_125_3477_n923), .CO(
        DP_OP_423J2_125_3477_n866), .S(DP_OP_423J2_125_3477_n867) );
  FADDX1_HVT DP_OP_423J2_125_3477_U589 ( .A(DP_OP_423J2_125_3477_n925), .B(
        DP_OP_423J2_125_3477_n907), .CI(DP_OP_423J2_125_3477_n901), .CO(
        DP_OP_423J2_125_3477_n864), .S(DP_OP_423J2_125_3477_n865) );
  FADDX1_HVT DP_OP_423J2_125_3477_U588 ( .A(DP_OP_423J2_125_3477_n927), .B(
        DP_OP_423J2_125_3477_n903), .CI(DP_OP_423J2_125_3477_n919), .CO(
        DP_OP_423J2_125_3477_n862), .S(DP_OP_423J2_125_3477_n863) );
  FADDX1_HVT DP_OP_423J2_125_3477_U587 ( .A(DP_OP_423J2_125_3477_n917), .B(
        DP_OP_423J2_125_3477_n915), .CI(DP_OP_423J2_125_3477_n905), .CO(
        DP_OP_423J2_125_3477_n860), .S(DP_OP_423J2_125_3477_n861) );
  FADDX1_HVT DP_OP_423J2_125_3477_U586 ( .A(DP_OP_423J2_125_3477_n921), .B(
        DP_OP_423J2_125_3477_n909), .CI(DP_OP_423J2_125_3477_n911), .CO(
        DP_OP_423J2_125_3477_n858), .S(DP_OP_423J2_125_3477_n859) );
  FADDX1_HVT DP_OP_423J2_125_3477_U585 ( .A(DP_OP_423J2_125_3477_n929), .B(
        DP_OP_423J2_125_3477_n933), .CI(DP_OP_423J2_125_3477_n931), .CO(
        DP_OP_423J2_125_3477_n856), .S(DP_OP_423J2_125_3477_n857) );
  FADDX1_HVT DP_OP_423J2_125_3477_U584 ( .A(DP_OP_423J2_125_3477_n913), .B(
        DP_OP_423J2_125_3477_n1092), .CI(DP_OP_423J2_125_3477_n1090), .CO(
        DP_OP_423J2_125_3477_n854), .S(DP_OP_423J2_125_3477_n855) );
  FADDX1_HVT DP_OP_423J2_125_3477_U583 ( .A(DP_OP_423J2_125_3477_n1088), .B(
        DP_OP_423J2_125_3477_n1086), .CI(DP_OP_423J2_125_3477_n1072), .CO(
        DP_OP_423J2_125_3477_n852), .S(DP_OP_423J2_125_3477_n853) );
  FADDX1_HVT DP_OP_423J2_125_3477_U582 ( .A(DP_OP_423J2_125_3477_n1084), .B(
        DP_OP_423J2_125_3477_n1082), .CI(DP_OP_423J2_125_3477_n1070), .CO(
        DP_OP_423J2_125_3477_n850), .S(DP_OP_423J2_125_3477_n851) );
  FADDX1_HVT DP_OP_423J2_125_3477_U581 ( .A(DP_OP_423J2_125_3477_n1080), .B(
        DP_OP_423J2_125_3477_n1074), .CI(DP_OP_423J2_125_3477_n1076), .CO(
        DP_OP_423J2_125_3477_n848), .S(DP_OP_423J2_125_3477_n849) );
  FADDX1_HVT DP_OP_423J2_125_3477_U580 ( .A(DP_OP_423J2_125_3477_n1078), .B(
        DP_OP_423J2_125_3477_n1068), .CI(DP_OP_423J2_125_3477_n1066), .CO(
        DP_OP_423J2_125_3477_n846), .S(DP_OP_423J2_125_3477_n847) );
  FADDX1_HVT DP_OP_423J2_125_3477_U579 ( .A(DP_OP_423J2_125_3477_n899), .B(
        DP_OP_423J2_125_3477_n895), .CI(DP_OP_423J2_125_3477_n1064), .CO(
        DP_OP_423J2_125_3477_n844), .S(DP_OP_423J2_125_3477_n845) );
  FADDX1_HVT DP_OP_423J2_125_3477_U578 ( .A(DP_OP_423J2_125_3477_n897), .B(
        DP_OP_423J2_125_3477_n1052), .CI(DP_OP_423J2_125_3477_n1050), .CO(
        DP_OP_423J2_125_3477_n842), .S(DP_OP_423J2_125_3477_n843) );
  FADDX1_HVT DP_OP_423J2_125_3477_U577 ( .A(DP_OP_423J2_125_3477_n1058), .B(
        DP_OP_423J2_125_3477_n893), .CI(DP_OP_423J2_125_3477_n1048), .CO(
        DP_OP_423J2_125_3477_n840), .S(DP_OP_423J2_125_3477_n841) );
  FADDX1_HVT DP_OP_423J2_125_3477_U576 ( .A(DP_OP_423J2_125_3477_n1056), .B(
        DP_OP_423J2_125_3477_n889), .CI(DP_OP_423J2_125_3477_n879), .CO(
        DP_OP_423J2_125_3477_n838), .S(DP_OP_423J2_125_3477_n839) );
  FADDX1_HVT DP_OP_423J2_125_3477_U575 ( .A(DP_OP_423J2_125_3477_n1062), .B(
        DP_OP_423J2_125_3477_n885), .CI(DP_OP_423J2_125_3477_n887), .CO(
        DP_OP_423J2_125_3477_n836), .S(DP_OP_423J2_125_3477_n837) );
  FADDX1_HVT DP_OP_423J2_125_3477_U574 ( .A(DP_OP_423J2_125_3477_n1060), .B(
        DP_OP_423J2_125_3477_n881), .CI(DP_OP_423J2_125_3477_n883), .CO(
        DP_OP_423J2_125_3477_n834), .S(DP_OP_423J2_125_3477_n835) );
  FADDX1_HVT DP_OP_423J2_125_3477_U573 ( .A(DP_OP_423J2_125_3477_n1054), .B(
        DP_OP_423J2_125_3477_n891), .CI(DP_OP_423J2_125_3477_n877), .CO(
        DP_OP_423J2_125_3477_n832), .S(DP_OP_423J2_125_3477_n833) );
  FADDX1_HVT DP_OP_423J2_125_3477_U572 ( .A(DP_OP_423J2_125_3477_n871), .B(
        DP_OP_423J2_125_3477_n875), .CI(DP_OP_423J2_125_3477_n867), .CO(
        DP_OP_423J2_125_3477_n830), .S(DP_OP_423J2_125_3477_n831) );
  FADDX1_HVT DP_OP_423J2_125_3477_U571 ( .A(DP_OP_423J2_125_3477_n869), .B(
        DP_OP_423J2_125_3477_n873), .CI(DP_OP_423J2_125_3477_n861), .CO(
        DP_OP_423J2_125_3477_n828), .S(DP_OP_423J2_125_3477_n829) );
  FADDX1_HVT DP_OP_423J2_125_3477_U570 ( .A(DP_OP_423J2_125_3477_n859), .B(
        DP_OP_423J2_125_3477_n865), .CI(DP_OP_423J2_125_3477_n1046), .CO(
        DP_OP_423J2_125_3477_n826), .S(DP_OP_423J2_125_3477_n827) );
  FADDX1_HVT DP_OP_423J2_125_3477_U569 ( .A(DP_OP_423J2_125_3477_n857), .B(
        DP_OP_423J2_125_3477_n863), .CI(DP_OP_423J2_125_3477_n1042), .CO(
        DP_OP_423J2_125_3477_n824), .S(DP_OP_423J2_125_3477_n825) );
  FADDX1_HVT DP_OP_423J2_125_3477_U568 ( .A(DP_OP_423J2_125_3477_n1044), .B(
        DP_OP_423J2_125_3477_n1040), .CI(DP_OP_423J2_125_3477_n855), .CO(
        DP_OP_423J2_125_3477_n822), .S(DP_OP_423J2_125_3477_n823) );
  FADDX1_HVT DP_OP_423J2_125_3477_U567 ( .A(DP_OP_423J2_125_3477_n1038), .B(
        DP_OP_423J2_125_3477_n1036), .CI(DP_OP_423J2_125_3477_n853), .CO(
        DP_OP_423J2_125_3477_n820), .S(DP_OP_423J2_125_3477_n821) );
  FADDX1_HVT DP_OP_423J2_125_3477_U566 ( .A(DP_OP_423J2_125_3477_n1034), .B(
        DP_OP_423J2_125_3477_n851), .CI(DP_OP_423J2_125_3477_n849), .CO(
        DP_OP_423J2_125_3477_n818), .S(DP_OP_423J2_125_3477_n819) );
  FADDX1_HVT DP_OP_423J2_125_3477_U565 ( .A(DP_OP_423J2_125_3477_n1032), .B(
        DP_OP_423J2_125_3477_n1026), .CI(DP_OP_423J2_125_3477_n1028), .CO(
        DP_OP_423J2_125_3477_n816), .S(DP_OP_423J2_125_3477_n817) );
  FADDX1_HVT DP_OP_423J2_125_3477_U564 ( .A(DP_OP_423J2_125_3477_n1030), .B(
        DP_OP_423J2_125_3477_n847), .CI(DP_OP_423J2_125_3477_n1024), .CO(
        DP_OP_423J2_125_3477_n814), .S(DP_OP_423J2_125_3477_n815) );
  FADDX1_HVT DP_OP_423J2_125_3477_U563 ( .A(DP_OP_423J2_125_3477_n845), .B(
        DP_OP_423J2_125_3477_n1022), .CI(DP_OP_423J2_125_3477_n843), .CO(
        DP_OP_423J2_125_3477_n812), .S(DP_OP_423J2_125_3477_n813) );
  FADDX1_HVT DP_OP_423J2_125_3477_U562 ( .A(DP_OP_423J2_125_3477_n1020), .B(
        DP_OP_423J2_125_3477_n837), .CI(DP_OP_423J2_125_3477_n833), .CO(
        DP_OP_423J2_125_3477_n810), .S(DP_OP_423J2_125_3477_n811) );
  FADDX1_HVT DP_OP_423J2_125_3477_U561 ( .A(DP_OP_423J2_125_3477_n1018), .B(
        DP_OP_423J2_125_3477_n841), .CI(DP_OP_423J2_125_3477_n839), .CO(
        DP_OP_423J2_125_3477_n808), .S(DP_OP_423J2_125_3477_n809) );
  FADDX1_HVT DP_OP_423J2_125_3477_U560 ( .A(DP_OP_423J2_125_3477_n835), .B(
        DP_OP_423J2_125_3477_n1016), .CI(DP_OP_423J2_125_3477_n831), .CO(
        DP_OP_423J2_125_3477_n806), .S(DP_OP_423J2_125_3477_n807) );
  FADDX1_HVT DP_OP_423J2_125_3477_U559 ( .A(DP_OP_423J2_125_3477_n829), .B(
        DP_OP_423J2_125_3477_n1014), .CI(DP_OP_423J2_125_3477_n827), .CO(
        DP_OP_423J2_125_3477_n804), .S(DP_OP_423J2_125_3477_n805) );
  FADDX1_HVT DP_OP_423J2_125_3477_U558 ( .A(DP_OP_423J2_125_3477_n825), .B(
        DP_OP_423J2_125_3477_n1012), .CI(DP_OP_423J2_125_3477_n1008), .CO(
        DP_OP_423J2_125_3477_n802), .S(DP_OP_423J2_125_3477_n803) );
  FADDX1_HVT DP_OP_423J2_125_3477_U557 ( .A(DP_OP_423J2_125_3477_n1010), .B(
        DP_OP_423J2_125_3477_n823), .CI(DP_OP_423J2_125_3477_n1006), .CO(
        DP_OP_423J2_125_3477_n800), .S(DP_OP_423J2_125_3477_n801) );
  FADDX1_HVT DP_OP_423J2_125_3477_U556 ( .A(DP_OP_423J2_125_3477_n821), .B(
        DP_OP_423J2_125_3477_n1004), .CI(DP_OP_423J2_125_3477_n1002), .CO(
        DP_OP_423J2_125_3477_n798), .S(DP_OP_423J2_125_3477_n799) );
  FADDX1_HVT DP_OP_423J2_125_3477_U555 ( .A(DP_OP_423J2_125_3477_n819), .B(
        DP_OP_423J2_125_3477_n1000), .CI(DP_OP_423J2_125_3477_n815), .CO(
        DP_OP_423J2_125_3477_n796), .S(DP_OP_423J2_125_3477_n797) );
  FADDX1_HVT DP_OP_423J2_125_3477_U554 ( .A(DP_OP_423J2_125_3477_n817), .B(
        DP_OP_423J2_125_3477_n998), .CI(DP_OP_423J2_125_3477_n813), .CO(
        DP_OP_423J2_125_3477_n794), .S(DP_OP_423J2_125_3477_n795) );
  FADDX1_HVT DP_OP_423J2_125_3477_U553 ( .A(DP_OP_423J2_125_3477_n996), .B(
        DP_OP_423J2_125_3477_n811), .CI(DP_OP_423J2_125_3477_n807), .CO(
        DP_OP_423J2_125_3477_n792), .S(DP_OP_423J2_125_3477_n793) );
  FADDX1_HVT DP_OP_423J2_125_3477_U552 ( .A(DP_OP_423J2_125_3477_n809), .B(
        DP_OP_423J2_125_3477_n994), .CI(DP_OP_423J2_125_3477_n805), .CO(
        DP_OP_423J2_125_3477_n790), .S(DP_OP_423J2_125_3477_n791) );
  FADDX1_HVT DP_OP_423J2_125_3477_U551 ( .A(DP_OP_423J2_125_3477_n992), .B(
        DP_OP_423J2_125_3477_n803), .CI(DP_OP_423J2_125_3477_n990), .CO(
        DP_OP_423J2_125_3477_n788), .S(DP_OP_423J2_125_3477_n789) );
  FADDX1_HVT DP_OP_423J2_125_3477_U550 ( .A(DP_OP_423J2_125_3477_n801), .B(
        DP_OP_423J2_125_3477_n988), .CI(DP_OP_423J2_125_3477_n799), .CO(
        DP_OP_423J2_125_3477_n786), .S(DP_OP_423J2_125_3477_n787) );
  FADDX1_HVT DP_OP_423J2_125_3477_U549 ( .A(DP_OP_423J2_125_3477_n986), .B(
        DP_OP_423J2_125_3477_n797), .CI(DP_OP_423J2_125_3477_n984), .CO(
        DP_OP_423J2_125_3477_n784), .S(DP_OP_423J2_125_3477_n785) );
  FADDX1_HVT DP_OP_423J2_125_3477_U548 ( .A(DP_OP_423J2_125_3477_n795), .B(
        DP_OP_423J2_125_3477_n793), .CI(DP_OP_423J2_125_3477_n982), .CO(
        DP_OP_423J2_125_3477_n782), .S(DP_OP_423J2_125_3477_n783) );
  FADDX1_HVT DP_OP_423J2_125_3477_U547 ( .A(DP_OP_423J2_125_3477_n791), .B(
        DP_OP_423J2_125_3477_n980), .CI(DP_OP_423J2_125_3477_n789), .CO(
        DP_OP_423J2_125_3477_n780), .S(DP_OP_423J2_125_3477_n781) );
  FADDX1_HVT DP_OP_423J2_125_3477_U546 ( .A(DP_OP_423J2_125_3477_n978), .B(
        DP_OP_423J2_125_3477_n787), .CI(DP_OP_423J2_125_3477_n976), .CO(
        DP_OP_423J2_125_3477_n778), .S(DP_OP_423J2_125_3477_n779) );
  FADDX1_HVT DP_OP_423J2_125_3477_U545 ( .A(DP_OP_423J2_125_3477_n785), .B(
        DP_OP_423J2_125_3477_n974), .CI(DP_OP_423J2_125_3477_n783), .CO(
        DP_OP_423J2_125_3477_n776), .S(DP_OP_423J2_125_3477_n777) );
  FADDX1_HVT DP_OP_423J2_125_3477_U544 ( .A(DP_OP_423J2_125_3477_n781), .B(
        DP_OP_423J2_125_3477_n972), .CI(DP_OP_423J2_125_3477_n779), .CO(
        DP_OP_423J2_125_3477_n774), .S(DP_OP_423J2_125_3477_n775) );
  FADDX1_HVT DP_OP_423J2_125_3477_U543 ( .A(DP_OP_423J2_125_3477_n970), .B(
        DP_OP_423J2_125_3477_n777), .CI(DP_OP_423J2_125_3477_n775), .CO(
        DP_OP_423J2_125_3477_n772), .S(DP_OP_423J2_125_3477_n773) );
  FADDX1_HVT DP_OP_423J2_125_3477_U541 ( .A(DP_OP_423J2_125_3477_n2186), .B(
        DP_OP_423J2_125_3477_n1922), .CI(DP_OP_423J2_125_3477_n1878), .CO(
        DP_OP_423J2_125_3477_n768), .S(DP_OP_423J2_125_3477_n769) );
  FADDX1_HVT DP_OP_423J2_125_3477_U540 ( .A(DP_OP_423J2_125_3477_n2758), .B(
        DP_OP_423J2_125_3477_n1980), .CI(DP_OP_423J2_125_3477_n2244), .CO(
        DP_OP_423J2_125_3477_n766), .S(DP_OP_423J2_125_3477_n767) );
  FADDX1_HVT DP_OP_423J2_125_3477_U539 ( .A(DP_OP_423J2_125_3477_n2230), .B(
        DP_OP_423J2_125_3477_n2990), .CI(DP_OP_423J2_125_3477_n2640), .CO(
        DP_OP_423J2_125_3477_n764), .S(DP_OP_423J2_125_3477_n765) );
  FADDX1_HVT DP_OP_423J2_125_3477_U538 ( .A(DP_OP_423J2_125_3477_n2450), .B(
        DP_OP_423J2_125_3477_n2024), .CI(DP_OP_423J2_125_3477_n2068), .CO(
        DP_OP_423J2_125_3477_n762), .S(DP_OP_423J2_125_3477_n763) );
  FADDX1_HVT DP_OP_423J2_125_3477_U537 ( .A(DP_OP_423J2_125_3477_n2010), .B(
        DP_OP_423J2_125_3477_n2112), .CI(DP_OP_423J2_125_3477_n2156), .CO(
        DP_OP_423J2_125_3477_n760), .S(DP_OP_423J2_125_3477_n761) );
  FADDX1_HVT DP_OP_423J2_125_3477_U536 ( .A(DP_OP_423J2_125_3477_n2714), .B(
        DP_OP_423J2_125_3477_n2816), .CI(DP_OP_423J2_125_3477_n2860), .CO(
        DP_OP_423J2_125_3477_n758), .S(DP_OP_423J2_125_3477_n759) );
  FADDX1_HVT DP_OP_423J2_125_3477_U535 ( .A(DP_OP_423J2_125_3477_n2054), .B(
        DP_OP_423J2_125_3477_n2772), .CI(DP_OP_423J2_125_3477_n2596), .CO(
        DP_OP_423J2_125_3477_n756), .S(DP_OP_423J2_125_3477_n757) );
  FADDX1_HVT DP_OP_423J2_125_3477_U534 ( .A(DP_OP_423J2_125_3477_n2142), .B(
        DP_OP_423J2_125_3477_n2420), .CI(DP_OP_423J2_125_3477_n2948), .CO(
        DP_OP_423J2_125_3477_n754), .S(DP_OP_423J2_125_3477_n755) );
  FADDX1_HVT DP_OP_423J2_125_3477_U533 ( .A(DP_OP_423J2_125_3477_n2670), .B(
        DP_OP_423J2_125_3477_n2904), .CI(DP_OP_423J2_125_3477_n2464), .CO(
        DP_OP_423J2_125_3477_n752), .S(DP_OP_423J2_125_3477_n753) );
  FADDX1_HVT DP_OP_423J2_125_3477_U532 ( .A(DP_OP_423J2_125_3477_n2626), .B(
        DP_OP_423J2_125_3477_n2376), .CI(DP_OP_423J2_125_3477_n2728), .CO(
        DP_OP_423J2_125_3477_n750), .S(DP_OP_423J2_125_3477_n751) );
  FADDX1_HVT DP_OP_423J2_125_3477_U531 ( .A(DP_OP_423J2_125_3477_n2846), .B(
        DP_OP_423J2_125_3477_n2508), .CI(DP_OP_423J2_125_3477_n2332), .CO(
        DP_OP_423J2_125_3477_n748), .S(DP_OP_423J2_125_3477_n749) );
  FADDX1_HVT DP_OP_423J2_125_3477_U530 ( .A(DP_OP_423J2_125_3477_n2318), .B(
        DP_OP_423J2_125_3477_n2288), .CI(DP_OP_423J2_125_3477_n1936), .CO(
        DP_OP_423J2_125_3477_n746), .S(DP_OP_423J2_125_3477_n747) );
  FADDX1_HVT DP_OP_423J2_125_3477_U529 ( .A(DP_OP_423J2_125_3477_n2538), .B(
        DP_OP_423J2_125_3477_n2200), .CI(DP_OP_423J2_125_3477_n2552), .CO(
        DP_OP_423J2_125_3477_n744), .S(DP_OP_423J2_125_3477_n745) );
  FADDX1_HVT DP_OP_423J2_125_3477_U528 ( .A(DP_OP_423J2_125_3477_n2494), .B(
        DP_OP_423J2_125_3477_n2362), .CI(DP_OP_423J2_125_3477_n2684), .CO(
        DP_OP_423J2_125_3477_n742), .S(DP_OP_423J2_125_3477_n743) );
  FADDX1_HVT DP_OP_423J2_125_3477_U527 ( .A(DP_OP_423J2_125_3477_n2802), .B(
        DP_OP_423J2_125_3477_n2098), .CI(DP_OP_423J2_125_3477_n2274), .CO(
        DP_OP_423J2_125_3477_n740), .S(DP_OP_423J2_125_3477_n741) );
  FADDX1_HVT DP_OP_423J2_125_3477_U526 ( .A(DP_OP_423J2_125_3477_n1966), .B(
        DP_OP_423J2_125_3477_n2582), .CI(DP_OP_423J2_125_3477_n2934), .CO(
        DP_OP_423J2_125_3477_n738), .S(DP_OP_423J2_125_3477_n739) );
  FADDX1_HVT DP_OP_423J2_125_3477_U525 ( .A(DP_OP_423J2_125_3477_n2890), .B(
        DP_OP_423J2_125_3477_n2406), .CI(DP_OP_423J2_125_3477_n771), .CO(
        DP_OP_423J2_125_3477_n736), .S(DP_OP_423J2_125_3477_n737) );
  FADDX1_HVT DP_OP_423J2_125_3477_U524 ( .A(DP_OP_423J2_125_3477_n2237), .B(
        DP_OP_423J2_125_3477_n1973), .CI(DP_OP_423J2_125_3477_n1929), .CO(
        DP_OP_423J2_125_3477_n734), .S(DP_OP_423J2_125_3477_n735) );
  FADDX1_HVT DP_OP_423J2_125_3477_U523 ( .A(DP_OP_423J2_125_3477_n2983), .B(
        DP_OP_423J2_125_3477_n2017), .CI(DP_OP_423J2_125_3477_n2061), .CO(
        DP_OP_423J2_125_3477_n732), .S(DP_OP_423J2_125_3477_n733) );
  FADDX1_HVT DP_OP_423J2_125_3477_U522 ( .A(DP_OP_423J2_125_3477_n2941), .B(
        DP_OP_423J2_125_3477_n2105), .CI(DP_OP_423J2_125_3477_n2149), .CO(
        DP_OP_423J2_125_3477_n730), .S(DP_OP_423J2_125_3477_n731) );
  FADDX1_HVT DP_OP_423J2_125_3477_U521 ( .A(DP_OP_423J2_125_3477_n2897), .B(
        DP_OP_423J2_125_3477_n2193), .CI(DP_OP_423J2_125_3477_n2281), .CO(
        DP_OP_423J2_125_3477_n728), .S(DP_OP_423J2_125_3477_n729) );
  FADDX1_HVT DP_OP_423J2_125_3477_U520 ( .A(DP_OP_423J2_125_3477_n2853), .B(
        DP_OP_423J2_125_3477_n2325), .CI(DP_OP_423J2_125_3477_n2369), .CO(
        DP_OP_423J2_125_3477_n726), .S(DP_OP_423J2_125_3477_n727) );
  FADDX1_HVT DP_OP_423J2_125_3477_U519 ( .A(DP_OP_423J2_125_3477_n2809), .B(
        DP_OP_423J2_125_3477_n2413), .CI(DP_OP_423J2_125_3477_n2457), .CO(
        DP_OP_423J2_125_3477_n724), .S(DP_OP_423J2_125_3477_n725) );
  FADDX1_HVT DP_OP_423J2_125_3477_U518 ( .A(DP_OP_423J2_125_3477_n2765), .B(
        DP_OP_423J2_125_3477_n2501), .CI(DP_OP_423J2_125_3477_n2545), .CO(
        DP_OP_423J2_125_3477_n722), .S(DP_OP_423J2_125_3477_n723) );
  FADDX1_HVT DP_OP_423J2_125_3477_U517 ( .A(DP_OP_423J2_125_3477_n2721), .B(
        DP_OP_423J2_125_3477_n2589), .CI(DP_OP_423J2_125_3477_n2633), .CO(
        DP_OP_423J2_125_3477_n720), .S(DP_OP_423J2_125_3477_n721) );
  FADDX1_HVT DP_OP_423J2_125_3477_U516 ( .A(DP_OP_423J2_125_3477_n2677), .B(
        DP_OP_423J2_125_3477_n966), .CI(DP_OP_423J2_125_3477_n964), .CO(
        DP_OP_423J2_125_3477_n718), .S(DP_OP_423J2_125_3477_n719) );
  FADDX1_HVT DP_OP_423J2_125_3477_U515 ( .A(DP_OP_423J2_125_3477_n962), .B(
        DP_OP_423J2_125_3477_n934), .CI(DP_OP_423J2_125_3477_n936), .CO(
        DP_OP_423J2_125_3477_n716), .S(DP_OP_423J2_125_3477_n717) );
  FADDX1_HVT DP_OP_423J2_125_3477_U514 ( .A(DP_OP_423J2_125_3477_n960), .B(
        DP_OP_423J2_125_3477_n938), .CI(DP_OP_423J2_125_3477_n940), .CO(
        DP_OP_423J2_125_3477_n714), .S(DP_OP_423J2_125_3477_n715) );
  FADDX1_HVT DP_OP_423J2_125_3477_U513 ( .A(DP_OP_423J2_125_3477_n958), .B(
        DP_OP_423J2_125_3477_n942), .CI(DP_OP_423J2_125_3477_n944), .CO(
        DP_OP_423J2_125_3477_n712), .S(DP_OP_423J2_125_3477_n713) );
  FADDX1_HVT DP_OP_423J2_125_3477_U512 ( .A(DP_OP_423J2_125_3477_n950), .B(
        DP_OP_423J2_125_3477_n956), .CI(DP_OP_423J2_125_3477_n946), .CO(
        DP_OP_423J2_125_3477_n710), .S(DP_OP_423J2_125_3477_n711) );
  FADDX1_HVT DP_OP_423J2_125_3477_U511 ( .A(DP_OP_423J2_125_3477_n948), .B(
        DP_OP_423J2_125_3477_n952), .CI(DP_OP_423J2_125_3477_n954), .CO(
        DP_OP_423J2_125_3477_n708), .S(DP_OP_423J2_125_3477_n709) );
  FADDX1_HVT DP_OP_423J2_125_3477_U510 ( .A(DP_OP_423J2_125_3477_n932), .B(
        DP_OP_423J2_125_3477_n930), .CI(DP_OP_423J2_125_3477_n900), .CO(
        DP_OP_423J2_125_3477_n706), .S(DP_OP_423J2_125_3477_n707) );
  FADDX1_HVT DP_OP_423J2_125_3477_U509 ( .A(DP_OP_423J2_125_3477_n914), .B(
        DP_OP_423J2_125_3477_n902), .CI(DP_OP_423J2_125_3477_n904), .CO(
        DP_OP_423J2_125_3477_n704), .S(DP_OP_423J2_125_3477_n705) );
  FADDX1_HVT DP_OP_423J2_125_3477_U508 ( .A(DP_OP_423J2_125_3477_n912), .B(
        DP_OP_423J2_125_3477_n906), .CI(DP_OP_423J2_125_3477_n908), .CO(
        DP_OP_423J2_125_3477_n702), .S(DP_OP_423J2_125_3477_n703) );
  FADDX1_HVT DP_OP_423J2_125_3477_U507 ( .A(DP_OP_423J2_125_3477_n910), .B(
        DP_OP_423J2_125_3477_n928), .CI(DP_OP_423J2_125_3477_n926), .CO(
        DP_OP_423J2_125_3477_n700), .S(DP_OP_423J2_125_3477_n701) );
  FADDX1_HVT DP_OP_423J2_125_3477_U506 ( .A(DP_OP_423J2_125_3477_n920), .B(
        DP_OP_423J2_125_3477_n916), .CI(DP_OP_423J2_125_3477_n918), .CO(
        DP_OP_423J2_125_3477_n698), .S(DP_OP_423J2_125_3477_n699) );
  FADDX1_HVT DP_OP_423J2_125_3477_U505 ( .A(DP_OP_423J2_125_3477_n924), .B(
        DP_OP_423J2_125_3477_n922), .CI(DP_OP_423J2_125_3477_n763), .CO(
        DP_OP_423J2_125_3477_n696), .S(DP_OP_423J2_125_3477_n697) );
  FADDX1_HVT DP_OP_423J2_125_3477_U504 ( .A(DP_OP_423J2_125_3477_n759), .B(
        DP_OP_423J2_125_3477_n755), .CI(DP_OP_423J2_125_3477_n737), .CO(
        DP_OP_423J2_125_3477_n694), .S(DP_OP_423J2_125_3477_n695) );
  FADDX1_HVT DP_OP_423J2_125_3477_U503 ( .A(DP_OP_423J2_125_3477_n761), .B(
        DP_OP_423J2_125_3477_n743), .CI(DP_OP_423J2_125_3477_n741), .CO(
        DP_OP_423J2_125_3477_n692), .S(DP_OP_423J2_125_3477_n693) );
  FADDX1_HVT DP_OP_423J2_125_3477_U502 ( .A(DP_OP_423J2_125_3477_n753), .B(
        DP_OP_423J2_125_3477_n757), .CI(DP_OP_423J2_125_3477_n749), .CO(
        DP_OP_423J2_125_3477_n690), .S(DP_OP_423J2_125_3477_n691) );
  FADDX1_HVT DP_OP_423J2_125_3477_U501 ( .A(DP_OP_423J2_125_3477_n765), .B(
        DP_OP_423J2_125_3477_n745), .CI(DP_OP_423J2_125_3477_n739), .CO(
        DP_OP_423J2_125_3477_n688), .S(DP_OP_423J2_125_3477_n689) );
  FADDX1_HVT DP_OP_423J2_125_3477_U500 ( .A(DP_OP_423J2_125_3477_n747), .B(
        DP_OP_423J2_125_3477_n769), .CI(DP_OP_423J2_125_3477_n767), .CO(
        DP_OP_423J2_125_3477_n686), .S(DP_OP_423J2_125_3477_n687) );
  FADDX1_HVT DP_OP_423J2_125_3477_U499 ( .A(DP_OP_423J2_125_3477_n751), .B(
        DP_OP_423J2_125_3477_n731), .CI(DP_OP_423J2_125_3477_n727), .CO(
        DP_OP_423J2_125_3477_n684), .S(DP_OP_423J2_125_3477_n685) );
  FADDX1_HVT DP_OP_423J2_125_3477_U498 ( .A(DP_OP_423J2_125_3477_n723), .B(
        DP_OP_423J2_125_3477_n721), .CI(DP_OP_423J2_125_3477_n733), .CO(
        DP_OP_423J2_125_3477_n682), .S(DP_OP_423J2_125_3477_n683) );
  FADDX1_HVT DP_OP_423J2_125_3477_U497 ( .A(DP_OP_423J2_125_3477_n729), .B(
        DP_OP_423J2_125_3477_n725), .CI(DP_OP_423J2_125_3477_n735), .CO(
        DP_OP_423J2_125_3477_n680), .S(DP_OP_423J2_125_3477_n681) );
  FADDX1_HVT DP_OP_423J2_125_3477_U496 ( .A(DP_OP_423J2_125_3477_n898), .B(
        DP_OP_423J2_125_3477_n894), .CI(DP_OP_423J2_125_3477_n896), .CO(
        DP_OP_423J2_125_3477_n678), .S(DP_OP_423J2_125_3477_n679) );
  FADDX1_HVT DP_OP_423J2_125_3477_U495 ( .A(DP_OP_423J2_125_3477_n892), .B(
        DP_OP_423J2_125_3477_n878), .CI(DP_OP_423J2_125_3477_n880), .CO(
        DP_OP_423J2_125_3477_n676), .S(DP_OP_423J2_125_3477_n677) );
  FADDX1_HVT DP_OP_423J2_125_3477_U494 ( .A(DP_OP_423J2_125_3477_n890), .B(
        DP_OP_423J2_125_3477_n882), .CI(DP_OP_423J2_125_3477_n888), .CO(
        DP_OP_423J2_125_3477_n674), .S(DP_OP_423J2_125_3477_n675) );
  FADDX1_HVT DP_OP_423J2_125_3477_U493 ( .A(DP_OP_423J2_125_3477_n886), .B(
        DP_OP_423J2_125_3477_n884), .CI(DP_OP_423J2_125_3477_n719), .CO(
        DP_OP_423J2_125_3477_n672), .S(DP_OP_423J2_125_3477_n673) );
  FADDX1_HVT DP_OP_423J2_125_3477_U492 ( .A(DP_OP_423J2_125_3477_n876), .B(
        DP_OP_423J2_125_3477_n717), .CI(DP_OP_423J2_125_3477_n715), .CO(
        DP_OP_423J2_125_3477_n670), .S(DP_OP_423J2_125_3477_n671) );
  FADDX1_HVT DP_OP_423J2_125_3477_U491 ( .A(DP_OP_423J2_125_3477_n874), .B(
        DP_OP_423J2_125_3477_n711), .CI(DP_OP_423J2_125_3477_n713), .CO(
        DP_OP_423J2_125_3477_n668), .S(DP_OP_423J2_125_3477_n669) );
  FADDX1_HVT DP_OP_423J2_125_3477_U490 ( .A(DP_OP_423J2_125_3477_n872), .B(
        DP_OP_423J2_125_3477_n709), .CI(DP_OP_423J2_125_3477_n866), .CO(
        DP_OP_423J2_125_3477_n666), .S(DP_OP_423J2_125_3477_n667) );
  FADDX1_HVT DP_OP_423J2_125_3477_U489 ( .A(DP_OP_423J2_125_3477_n870), .B(
        DP_OP_423J2_125_3477_n868), .CI(DP_OP_423J2_125_3477_n856), .CO(
        DP_OP_423J2_125_3477_n664), .S(DP_OP_423J2_125_3477_n665) );
  FADDX1_HVT DP_OP_423J2_125_3477_U488 ( .A(DP_OP_423J2_125_3477_n864), .B(
        DP_OP_423J2_125_3477_n707), .CI(DP_OP_423J2_125_3477_n697), .CO(
        DP_OP_423J2_125_3477_n662), .S(DP_OP_423J2_125_3477_n663) );
  FADDX1_HVT DP_OP_423J2_125_3477_U487 ( .A(DP_OP_423J2_125_3477_n862), .B(
        DP_OP_423J2_125_3477_n703), .CI(DP_OP_423J2_125_3477_n699), .CO(
        DP_OP_423J2_125_3477_n660), .S(DP_OP_423J2_125_3477_n661) );
  FADDX1_HVT DP_OP_423J2_125_3477_U486 ( .A(DP_OP_423J2_125_3477_n860), .B(
        DP_OP_423J2_125_3477_n705), .CI(DP_OP_423J2_125_3477_n701), .CO(
        DP_OP_423J2_125_3477_n658), .S(DP_OP_423J2_125_3477_n659) );
  FADDX1_HVT DP_OP_423J2_125_3477_U485 ( .A(DP_OP_423J2_125_3477_n858), .B(
        DP_OP_423J2_125_3477_n693), .CI(DP_OP_423J2_125_3477_n689), .CO(
        DP_OP_423J2_125_3477_n656), .S(DP_OP_423J2_125_3477_n657) );
  FADDX1_HVT DP_OP_423J2_125_3477_U484 ( .A(DP_OP_423J2_125_3477_n691), .B(
        DP_OP_423J2_125_3477_n854), .CI(DP_OP_423J2_125_3477_n685), .CO(
        DP_OP_423J2_125_3477_n654), .S(DP_OP_423J2_125_3477_n655) );
  FADDX1_HVT DP_OP_423J2_125_3477_U483 ( .A(DP_OP_423J2_125_3477_n687), .B(
        DP_OP_423J2_125_3477_n695), .CI(DP_OP_423J2_125_3477_n681), .CO(
        DP_OP_423J2_125_3477_n652), .S(DP_OP_423J2_125_3477_n653) );
  FADDX1_HVT DP_OP_423J2_125_3477_U482 ( .A(DP_OP_423J2_125_3477_n683), .B(
        DP_OP_423J2_125_3477_n852), .CI(DP_OP_423J2_125_3477_n850), .CO(
        DP_OP_423J2_125_3477_n650), .S(DP_OP_423J2_125_3477_n651) );
  FADDX1_HVT DP_OP_423J2_125_3477_U481 ( .A(DP_OP_423J2_125_3477_n848), .B(
        DP_OP_423J2_125_3477_n846), .CI(DP_OP_423J2_125_3477_n679), .CO(
        DP_OP_423J2_125_3477_n648), .S(DP_OP_423J2_125_3477_n649) );
  FADDX1_HVT DP_OP_423J2_125_3477_U480 ( .A(DP_OP_423J2_125_3477_n844), .B(
        DP_OP_423J2_125_3477_n842), .CI(DP_OP_423J2_125_3477_n840), .CO(
        DP_OP_423J2_125_3477_n646), .S(DP_OP_423J2_125_3477_n647) );
  FADDX1_HVT DP_OP_423J2_125_3477_U479 ( .A(DP_OP_423J2_125_3477_n838), .B(
        DP_OP_423J2_125_3477_n673), .CI(DP_OP_423J2_125_3477_n832), .CO(
        DP_OP_423J2_125_3477_n644), .S(DP_OP_423J2_125_3477_n645) );
  FADDX1_HVT DP_OP_423J2_125_3477_U478 ( .A(DP_OP_423J2_125_3477_n836), .B(
        DP_OP_423J2_125_3477_n675), .CI(DP_OP_423J2_125_3477_n677), .CO(
        DP_OP_423J2_125_3477_n642), .S(DP_OP_423J2_125_3477_n643) );
  FADDX1_HVT DP_OP_423J2_125_3477_U477 ( .A(DP_OP_423J2_125_3477_n834), .B(
        DP_OP_423J2_125_3477_n671), .CI(DP_OP_423J2_125_3477_n667), .CO(
        DP_OP_423J2_125_3477_n640), .S(DP_OP_423J2_125_3477_n641) );
  FADDX1_HVT DP_OP_423J2_125_3477_U476 ( .A(DP_OP_423J2_125_3477_n830), .B(
        DP_OP_423J2_125_3477_n669), .CI(DP_OP_423J2_125_3477_n665), .CO(
        DP_OP_423J2_125_3477_n638), .S(DP_OP_423J2_125_3477_n639) );
  FADDX1_HVT DP_OP_423J2_125_3477_U475 ( .A(DP_OP_423J2_125_3477_n828), .B(
        DP_OP_423J2_125_3477_n826), .CI(DP_OP_423J2_125_3477_n661), .CO(
        DP_OP_423J2_125_3477_n636), .S(DP_OP_423J2_125_3477_n637) );
  FADDX1_HVT DP_OP_423J2_125_3477_U474 ( .A(DP_OP_423J2_125_3477_n659), .B(
        DP_OP_423J2_125_3477_n663), .CI(DP_OP_423J2_125_3477_n824), .CO(
        DP_OP_423J2_125_3477_n634), .S(DP_OP_423J2_125_3477_n635) );
  FADDX1_HVT DP_OP_423J2_125_3477_U473 ( .A(DP_OP_423J2_125_3477_n657), .B(
        DP_OP_423J2_125_3477_n822), .CI(DP_OP_423J2_125_3477_n653), .CO(
        DP_OP_423J2_125_3477_n632), .S(DP_OP_423J2_125_3477_n633) );
  FADDX1_HVT DP_OP_423J2_125_3477_U472 ( .A(DP_OP_423J2_125_3477_n655), .B(
        DP_OP_423J2_125_3477_n820), .CI(DP_OP_423J2_125_3477_n651), .CO(
        DP_OP_423J2_125_3477_n630), .S(DP_OP_423J2_125_3477_n631) );
  FADDX1_HVT DP_OP_423J2_125_3477_U471 ( .A(DP_OP_423J2_125_3477_n818), .B(
        DP_OP_423J2_125_3477_n816), .CI(DP_OP_423J2_125_3477_n649), .CO(
        DP_OP_423J2_125_3477_n628), .S(DP_OP_423J2_125_3477_n629) );
  FADDX1_HVT DP_OP_423J2_125_3477_U470 ( .A(DP_OP_423J2_125_3477_n814), .B(
        DP_OP_423J2_125_3477_n812), .CI(DP_OP_423J2_125_3477_n647), .CO(
        DP_OP_423J2_125_3477_n626), .S(DP_OP_423J2_125_3477_n627) );
  FADDX1_HVT DP_OP_423J2_125_3477_U469 ( .A(DP_OP_423J2_125_3477_n810), .B(
        DP_OP_423J2_125_3477_n643), .CI(DP_OP_423J2_125_3477_n806), .CO(
        DP_OP_423J2_125_3477_n624), .S(DP_OP_423J2_125_3477_n625) );
  FADDX1_HVT DP_OP_423J2_125_3477_U468 ( .A(DP_OP_423J2_125_3477_n808), .B(
        DP_OP_423J2_125_3477_n645), .CI(DP_OP_423J2_125_3477_n641), .CO(
        DP_OP_423J2_125_3477_n622), .S(DP_OP_423J2_125_3477_n623) );
  FADDX1_HVT DP_OP_423J2_125_3477_U467 ( .A(DP_OP_423J2_125_3477_n639), .B(
        DP_OP_423J2_125_3477_n804), .CI(DP_OP_423J2_125_3477_n637), .CO(
        DP_OP_423J2_125_3477_n620), .S(DP_OP_423J2_125_3477_n621) );
  FADDX1_HVT DP_OP_423J2_125_3477_U466 ( .A(DP_OP_423J2_125_3477_n635), .B(
        DP_OP_423J2_125_3477_n802), .CI(DP_OP_423J2_125_3477_n633), .CO(
        DP_OP_423J2_125_3477_n618), .S(DP_OP_423J2_125_3477_n619) );
  FADDX1_HVT DP_OP_423J2_125_3477_U465 ( .A(DP_OP_423J2_125_3477_n800), .B(
        DP_OP_423J2_125_3477_n631), .CI(DP_OP_423J2_125_3477_n798), .CO(
        DP_OP_423J2_125_3477_n616), .S(DP_OP_423J2_125_3477_n617) );
  FADDX1_HVT DP_OP_423J2_125_3477_U464 ( .A(DP_OP_423J2_125_3477_n796), .B(
        DP_OP_423J2_125_3477_n629), .CI(DP_OP_423J2_125_3477_n794), .CO(
        DP_OP_423J2_125_3477_n614), .S(DP_OP_423J2_125_3477_n615) );
  FADDX1_HVT DP_OP_423J2_125_3477_U463 ( .A(DP_OP_423J2_125_3477_n627), .B(
        DP_OP_423J2_125_3477_n792), .CI(DP_OP_423J2_125_3477_n625), .CO(
        DP_OP_423J2_125_3477_n612), .S(DP_OP_423J2_125_3477_n613) );
  FADDX1_HVT DP_OP_423J2_125_3477_U462 ( .A(DP_OP_423J2_125_3477_n623), .B(
        DP_OP_423J2_125_3477_n790), .CI(DP_OP_423J2_125_3477_n621), .CO(
        DP_OP_423J2_125_3477_n610), .S(DP_OP_423J2_125_3477_n611) );
  FADDX1_HVT DP_OP_423J2_125_3477_U461 ( .A(DP_OP_423J2_125_3477_n788), .B(
        DP_OP_423J2_125_3477_n619), .CI(DP_OP_423J2_125_3477_n786), .CO(
        DP_OP_423J2_125_3477_n608), .S(DP_OP_423J2_125_3477_n609) );
  FADDX1_HVT DP_OP_423J2_125_3477_U460 ( .A(DP_OP_423J2_125_3477_n617), .B(
        DP_OP_423J2_125_3477_n784), .CI(DP_OP_423J2_125_3477_n615), .CO(
        DP_OP_423J2_125_3477_n606), .S(DP_OP_423J2_125_3477_n607) );
  FADDX1_HVT DP_OP_423J2_125_3477_U459 ( .A(DP_OP_423J2_125_3477_n782), .B(
        DP_OP_423J2_125_3477_n613), .CI(DP_OP_423J2_125_3477_n611), .CO(
        DP_OP_423J2_125_3477_n604), .S(DP_OP_423J2_125_3477_n605) );
  FADDX1_HVT DP_OP_423J2_125_3477_U458 ( .A(DP_OP_423J2_125_3477_n780), .B(
        DP_OP_423J2_125_3477_n609), .CI(DP_OP_423J2_125_3477_n778), .CO(
        DP_OP_423J2_125_3477_n602), .S(DP_OP_423J2_125_3477_n603) );
  FADDX1_HVT DP_OP_423J2_125_3477_U457 ( .A(DP_OP_423J2_125_3477_n607), .B(
        DP_OP_423J2_125_3477_n776), .CI(DP_OP_423J2_125_3477_n605), .CO(
        DP_OP_423J2_125_3477_n600), .S(DP_OP_423J2_125_3477_n601) );
  FADDX1_HVT DP_OP_423J2_125_3477_U456 ( .A(DP_OP_423J2_125_3477_n774), .B(
        DP_OP_423J2_125_3477_n603), .CI(DP_OP_423J2_125_3477_n601), .CO(
        DP_OP_423J2_125_3477_n598), .S(DP_OP_423J2_125_3477_n599) );
  FADDX1_HVT DP_OP_423J2_125_3477_U455 ( .A(DP_OP_423J2_125_3477_n2977), .B(
        DP_OP_423J2_125_3477_n1921), .CI(DP_OP_423J2_125_3477_n1877), .CO(
        DP_OP_423J2_125_3477_n596), .S(DP_OP_423J2_125_3477_n597) );
  FADDX1_HVT DP_OP_423J2_125_3477_U454 ( .A(DP_OP_423J2_125_3477_n770), .B(
        DP_OP_423J2_125_3477_n2236), .CI(DP_OP_423J2_125_3477_n1928), .CO(
        DP_OP_423J2_125_3477_n594), .S(DP_OP_423J2_125_3477_n595) );
  FADDX1_HVT DP_OP_423J2_125_3477_U453 ( .A(DP_OP_423J2_125_3477_n2317), .B(
        DP_OP_423J2_125_3477_n2982), .CI(DP_OP_423J2_125_3477_n2632), .CO(
        DP_OP_423J2_125_3477_n592), .S(DP_OP_423J2_125_3477_n593) );
  FADDX1_HVT DP_OP_423J2_125_3477_U452 ( .A(DP_OP_423J2_125_3477_n2009), .B(
        DP_OP_423J2_125_3477_n2544), .CI(DP_OP_423J2_125_3477_n2764), .CO(
        DP_OP_423J2_125_3477_n590), .S(DP_OP_423J2_125_3477_n591) );
  FADDX1_HVT DP_OP_423J2_125_3477_U451 ( .A(DP_OP_423J2_125_3477_n2229), .B(
        DP_OP_423J2_125_3477_n2324), .CI(DP_OP_423J2_125_3477_n2940), .CO(
        DP_OP_423J2_125_3477_n588), .S(DP_OP_423J2_125_3477_n589) );
  FADDX1_HVT DP_OP_423J2_125_3477_U450 ( .A(DP_OP_423J2_125_3477_n1965), .B(
        DP_OP_423J2_125_3477_n2852), .CI(DP_OP_423J2_125_3477_n2016), .CO(
        DP_OP_423J2_125_3477_n586), .S(DP_OP_423J2_125_3477_n587) );
  FADDX1_HVT DP_OP_423J2_125_3477_U449 ( .A(DP_OP_423J2_125_3477_n2097), .B(
        DP_OP_423J2_125_3477_n1972), .CI(DP_OP_423J2_125_3477_n2808), .CO(
        DP_OP_423J2_125_3477_n584), .S(DP_OP_423J2_125_3477_n585) );
  FADDX1_HVT DP_OP_423J2_125_3477_U448 ( .A(DP_OP_423J2_125_3477_n2933), .B(
        DP_OP_423J2_125_3477_n2368), .CI(DP_OP_423J2_125_3477_n2456), .CO(
        DP_OP_423J2_125_3477_n582), .S(DP_OP_423J2_125_3477_n583) );
  FADDX1_HVT DP_OP_423J2_125_3477_U447 ( .A(DP_OP_423J2_125_3477_n2449), .B(
        DP_OP_423J2_125_3477_n2500), .CI(DP_OP_423J2_125_3477_n2896), .CO(
        DP_OP_423J2_125_3477_n580), .S(DP_OP_423J2_125_3477_n581) );
  FADDX1_HVT DP_OP_423J2_125_3477_U446 ( .A(DP_OP_423J2_125_3477_n2713), .B(
        DP_OP_423J2_125_3477_n2192), .CI(DP_OP_423J2_125_3477_n2720), .CO(
        DP_OP_423J2_125_3477_n578), .S(DP_OP_423J2_125_3477_n579) );
  FADDX1_HVT DP_OP_423J2_125_3477_U445 ( .A(DP_OP_423J2_125_3477_n2889), .B(
        DP_OP_423J2_125_3477_n2412), .CI(DP_OP_423J2_125_3477_n2588), .CO(
        DP_OP_423J2_125_3477_n576), .S(DP_OP_423J2_125_3477_n577) );
  FADDX1_HVT DP_OP_423J2_125_3477_U444 ( .A(DP_OP_423J2_125_3477_n2185), .B(
        DP_OP_423J2_125_3477_n2060), .CI(DP_OP_423J2_125_3477_n2676), .CO(
        DP_OP_423J2_125_3477_n574), .S(DP_OP_423J2_125_3477_n575) );
  FADDX1_HVT DP_OP_423J2_125_3477_U443 ( .A(DP_OP_423J2_125_3477_n2141), .B(
        DP_OP_423J2_125_3477_n2280), .CI(DP_OP_423J2_125_3477_n2148), .CO(
        DP_OP_423J2_125_3477_n572), .S(DP_OP_423J2_125_3477_n573) );
  FADDX1_HVT DP_OP_423J2_125_3477_U442 ( .A(DP_OP_423J2_125_3477_n2537), .B(
        DP_OP_423J2_125_3477_n2361), .CI(DP_OP_423J2_125_3477_n2104), .CO(
        DP_OP_423J2_125_3477_n570), .S(DP_OP_423J2_125_3477_n571) );
  FADDX1_HVT DP_OP_423J2_125_3477_U441 ( .A(DP_OP_423J2_125_3477_n2845), .B(
        DP_OP_423J2_125_3477_n2053), .CI(DP_OP_423J2_125_3477_n2273), .CO(
        DP_OP_423J2_125_3477_n568), .S(DP_OP_423J2_125_3477_n569) );
  FADDX1_HVT DP_OP_423J2_125_3477_U440 ( .A(DP_OP_423J2_125_3477_n2801), .B(
        DP_OP_423J2_125_3477_n2405), .CI(DP_OP_423J2_125_3477_n2493), .CO(
        DP_OP_423J2_125_3477_n566), .S(DP_OP_423J2_125_3477_n567) );
  FADDX1_HVT DP_OP_423J2_125_3477_U439 ( .A(DP_OP_423J2_125_3477_n2757), .B(
        DP_OP_423J2_125_3477_n2581), .CI(DP_OP_423J2_125_3477_n2625), .CO(
        DP_OP_423J2_125_3477_n564), .S(DP_OP_423J2_125_3477_n565) );
  FADDX1_HVT DP_OP_423J2_125_3477_U438 ( .A(DP_OP_423J2_125_3477_n2669), .B(
        DP_OP_423J2_125_3477_n768), .CI(DP_OP_423J2_125_3477_n766), .CO(
        DP_OP_423J2_125_3477_n562), .S(DP_OP_423J2_125_3477_n563) );
  FADDX1_HVT DP_OP_423J2_125_3477_U437 ( .A(DP_OP_423J2_125_3477_n764), .B(
        DP_OP_423J2_125_3477_n736), .CI(DP_OP_423J2_125_3477_n738), .CO(
        DP_OP_423J2_125_3477_n560), .S(DP_OP_423J2_125_3477_n561) );
  FADDX1_HVT DP_OP_423J2_125_3477_U436 ( .A(DP_OP_423J2_125_3477_n762), .B(
        DP_OP_423J2_125_3477_n740), .CI(DP_OP_423J2_125_3477_n742), .CO(
        DP_OP_423J2_125_3477_n558), .S(DP_OP_423J2_125_3477_n559) );
  FADDX1_HVT DP_OP_423J2_125_3477_U435 ( .A(DP_OP_423J2_125_3477_n760), .B(
        DP_OP_423J2_125_3477_n744), .CI(DP_OP_423J2_125_3477_n746), .CO(
        DP_OP_423J2_125_3477_n556), .S(DP_OP_423J2_125_3477_n557) );
  FADDX1_HVT DP_OP_423J2_125_3477_U434 ( .A(DP_OP_423J2_125_3477_n758), .B(
        DP_OP_423J2_125_3477_n748), .CI(DP_OP_423J2_125_3477_n750), .CO(
        DP_OP_423J2_125_3477_n554), .S(DP_OP_423J2_125_3477_n555) );
  FADDX1_HVT DP_OP_423J2_125_3477_U433 ( .A(DP_OP_423J2_125_3477_n756), .B(
        DP_OP_423J2_125_3477_n752), .CI(DP_OP_423J2_125_3477_n754), .CO(
        DP_OP_423J2_125_3477_n552), .S(DP_OP_423J2_125_3477_n553) );
  FADDX1_HVT DP_OP_423J2_125_3477_U432 ( .A(DP_OP_423J2_125_3477_n734), .B(
        DP_OP_423J2_125_3477_n720), .CI(DP_OP_423J2_125_3477_n732), .CO(
        DP_OP_423J2_125_3477_n550), .S(DP_OP_423J2_125_3477_n551) );
  FADDX1_HVT DP_OP_423J2_125_3477_U431 ( .A(DP_OP_423J2_125_3477_n726), .B(
        DP_OP_423J2_125_3477_n722), .CI(DP_OP_423J2_125_3477_n724), .CO(
        DP_OP_423J2_125_3477_n548), .S(DP_OP_423J2_125_3477_n549) );
  FADDX1_HVT DP_OP_423J2_125_3477_U430 ( .A(DP_OP_423J2_125_3477_n730), .B(
        DP_OP_423J2_125_3477_n728), .CI(DP_OP_423J2_125_3477_n595), .CO(
        DP_OP_423J2_125_3477_n546), .S(DP_OP_423J2_125_3477_n547) );
  FADDX1_HVT DP_OP_423J2_125_3477_U429 ( .A(DP_OP_423J2_125_3477_n597), .B(
        DP_OP_423J2_125_3477_n583), .CI(DP_OP_423J2_125_3477_n589), .CO(
        DP_OP_423J2_125_3477_n544), .S(DP_OP_423J2_125_3477_n545) );
  FADDX1_HVT DP_OP_423J2_125_3477_U428 ( .A(DP_OP_423J2_125_3477_n565), .B(
        DP_OP_423J2_125_3477_n587), .CI(DP_OP_423J2_125_3477_n585), .CO(
        DP_OP_423J2_125_3477_n542), .S(DP_OP_423J2_125_3477_n543) );
  FADDX1_HVT DP_OP_423J2_125_3477_U427 ( .A(DP_OP_423J2_125_3477_n591), .B(
        DP_OP_423J2_125_3477_n573), .CI(DP_OP_423J2_125_3477_n575), .CO(
        DP_OP_423J2_125_3477_n540), .S(DP_OP_423J2_125_3477_n541) );
  FADDX1_HVT DP_OP_423J2_125_3477_U426 ( .A(DP_OP_423J2_125_3477_n577), .B(
        DP_OP_423J2_125_3477_n567), .CI(DP_OP_423J2_125_3477_n569), .CO(
        DP_OP_423J2_125_3477_n538), .S(DP_OP_423J2_125_3477_n539) );
  FADDX1_HVT DP_OP_423J2_125_3477_U425 ( .A(DP_OP_423J2_125_3477_n571), .B(
        DP_OP_423J2_125_3477_n593), .CI(DP_OP_423J2_125_3477_n581), .CO(
        DP_OP_423J2_125_3477_n536), .S(DP_OP_423J2_125_3477_n537) );
  FADDX1_HVT DP_OP_423J2_125_3477_U424 ( .A(DP_OP_423J2_125_3477_n579), .B(
        DP_OP_423J2_125_3477_n718), .CI(DP_OP_423J2_125_3477_n716), .CO(
        DP_OP_423J2_125_3477_n534), .S(DP_OP_423J2_125_3477_n535) );
  FADDX1_HVT DP_OP_423J2_125_3477_U423 ( .A(DP_OP_423J2_125_3477_n714), .B(
        DP_OP_423J2_125_3477_n708), .CI(DP_OP_423J2_125_3477_n710), .CO(
        DP_OP_423J2_125_3477_n532), .S(DP_OP_423J2_125_3477_n533) );
  FADDX1_HVT DP_OP_423J2_125_3477_U422 ( .A(DP_OP_423J2_125_3477_n712), .B(
        DP_OP_423J2_125_3477_n706), .CI(DP_OP_423J2_125_3477_n704), .CO(
        DP_OP_423J2_125_3477_n530), .S(DP_OP_423J2_125_3477_n531) );
  FADDX1_HVT DP_OP_423J2_125_3477_U421 ( .A(DP_OP_423J2_125_3477_n702), .B(
        DP_OP_423J2_125_3477_n698), .CI(DP_OP_423J2_125_3477_n696), .CO(
        DP_OP_423J2_125_3477_n528), .S(DP_OP_423J2_125_3477_n529) );
  FADDX1_HVT DP_OP_423J2_125_3477_U420 ( .A(DP_OP_423J2_125_3477_n700), .B(
        DP_OP_423J2_125_3477_n563), .CI(DP_OP_423J2_125_3477_n557), .CO(
        DP_OP_423J2_125_3477_n526), .S(DP_OP_423J2_125_3477_n527) );
  FADDX1_HVT DP_OP_423J2_125_3477_U419 ( .A(DP_OP_423J2_125_3477_n559), .B(
        DP_OP_423J2_125_3477_n553), .CI(DP_OP_423J2_125_3477_n684), .CO(
        DP_OP_423J2_125_3477_n524), .S(DP_OP_423J2_125_3477_n525) );
  FADDX1_HVT DP_OP_423J2_125_3477_U418 ( .A(DP_OP_423J2_125_3477_n694), .B(
        DP_OP_423J2_125_3477_n561), .CI(DP_OP_423J2_125_3477_n555), .CO(
        DP_OP_423J2_125_3477_n522), .S(DP_OP_423J2_125_3477_n523) );
  FADDX1_HVT DP_OP_423J2_125_3477_U417 ( .A(DP_OP_423J2_125_3477_n688), .B(
        DP_OP_423J2_125_3477_n692), .CI(DP_OP_423J2_125_3477_n686), .CO(
        DP_OP_423J2_125_3477_n520), .S(DP_OP_423J2_125_3477_n521) );
  FADDX1_HVT DP_OP_423J2_125_3477_U416 ( .A(DP_OP_423J2_125_3477_n690), .B(
        DP_OP_423J2_125_3477_n682), .CI(DP_OP_423J2_125_3477_n680), .CO(
        DP_OP_423J2_125_3477_n518), .S(DP_OP_423J2_125_3477_n519) );
  FADDX1_HVT DP_OP_423J2_125_3477_U415 ( .A(DP_OP_423J2_125_3477_n549), .B(
        DP_OP_423J2_125_3477_n551), .CI(DP_OP_423J2_125_3477_n547), .CO(
        DP_OP_423J2_125_3477_n516), .S(DP_OP_423J2_125_3477_n517) );
  FADDX1_HVT DP_OP_423J2_125_3477_U414 ( .A(DP_OP_423J2_125_3477_n545), .B(
        DP_OP_423J2_125_3477_n539), .CI(DP_OP_423J2_125_3477_n543), .CO(
        DP_OP_423J2_125_3477_n514), .S(DP_OP_423J2_125_3477_n515) );
  FADDX1_HVT DP_OP_423J2_125_3477_U413 ( .A(DP_OP_423J2_125_3477_n537), .B(
        DP_OP_423J2_125_3477_n541), .CI(DP_OP_423J2_125_3477_n678), .CO(
        DP_OP_423J2_125_3477_n512), .S(DP_OP_423J2_125_3477_n513) );
  FADDX1_HVT DP_OP_423J2_125_3477_U412 ( .A(DP_OP_423J2_125_3477_n676), .B(
        DP_OP_423J2_125_3477_n672), .CI(DP_OP_423J2_125_3477_n535), .CO(
        DP_OP_423J2_125_3477_n510), .S(DP_OP_423J2_125_3477_n511) );
  FADDX1_HVT DP_OP_423J2_125_3477_U411 ( .A(DP_OP_423J2_125_3477_n674), .B(
        DP_OP_423J2_125_3477_n670), .CI(DP_OP_423J2_125_3477_n668), .CO(
        DP_OP_423J2_125_3477_n508), .S(DP_OP_423J2_125_3477_n509) );
  FADDX1_HVT DP_OP_423J2_125_3477_U410 ( .A(DP_OP_423J2_125_3477_n666), .B(
        DP_OP_423J2_125_3477_n533), .CI(DP_OP_423J2_125_3477_n531), .CO(
        DP_OP_423J2_125_3477_n506), .S(DP_OP_423J2_125_3477_n507) );
  FADDX1_HVT DP_OP_423J2_125_3477_U409 ( .A(DP_OP_423J2_125_3477_n664), .B(
        DP_OP_423J2_125_3477_n662), .CI(DP_OP_423J2_125_3477_n660), .CO(
        DP_OP_423J2_125_3477_n504), .S(DP_OP_423J2_125_3477_n505) );
  FADDX1_HVT DP_OP_423J2_125_3477_U408 ( .A(DP_OP_423J2_125_3477_n658), .B(
        DP_OP_423J2_125_3477_n529), .CI(DP_OP_423J2_125_3477_n656), .CO(
        DP_OP_423J2_125_3477_n502), .S(DP_OP_423J2_125_3477_n503) );
  FADDX1_HVT DP_OP_423J2_125_3477_U407 ( .A(DP_OP_423J2_125_3477_n527), .B(
        DP_OP_423J2_125_3477_n654), .CI(DP_OP_423J2_125_3477_n525), .CO(
        DP_OP_423J2_125_3477_n500), .S(DP_OP_423J2_125_3477_n501) );
  FADDX1_HVT DP_OP_423J2_125_3477_U406 ( .A(DP_OP_423J2_125_3477_n652), .B(
        DP_OP_423J2_125_3477_n521), .CI(DP_OP_423J2_125_3477_n519), .CO(
        DP_OP_423J2_125_3477_n498), .S(DP_OP_423J2_125_3477_n499) );
  FADDX1_HVT DP_OP_423J2_125_3477_U405 ( .A(DP_OP_423J2_125_3477_n523), .B(
        DP_OP_423J2_125_3477_n517), .CI(DP_OP_423J2_125_3477_n650), .CO(
        DP_OP_423J2_125_3477_n496), .S(DP_OP_423J2_125_3477_n497) );
  FADDX1_HVT DP_OP_423J2_125_3477_U404 ( .A(DP_OP_423J2_125_3477_n515), .B(
        DP_OP_423J2_125_3477_n648), .CI(DP_OP_423J2_125_3477_n513), .CO(
        DP_OP_423J2_125_3477_n494), .S(DP_OP_423J2_125_3477_n495) );
  FADDX1_HVT DP_OP_423J2_125_3477_U403 ( .A(DP_OP_423J2_125_3477_n646), .B(
        DP_OP_423J2_125_3477_n644), .CI(DP_OP_423J2_125_3477_n642), .CO(
        DP_OP_423J2_125_3477_n492), .S(DP_OP_423J2_125_3477_n493) );
  FADDX1_HVT DP_OP_423J2_125_3477_U402 ( .A(DP_OP_423J2_125_3477_n511), .B(
        DP_OP_423J2_125_3477_n640), .CI(DP_OP_423J2_125_3477_n509), .CO(
        DP_OP_423J2_125_3477_n490), .S(DP_OP_423J2_125_3477_n491) );
  FADDX1_HVT DP_OP_423J2_125_3477_U401 ( .A(DP_OP_423J2_125_3477_n638), .B(
        DP_OP_423J2_125_3477_n507), .CI(DP_OP_423J2_125_3477_n505), .CO(
        DP_OP_423J2_125_3477_n488), .S(DP_OP_423J2_125_3477_n489) );
  FADDX1_HVT DP_OP_423J2_125_3477_U400 ( .A(DP_OP_423J2_125_3477_n636), .B(
        DP_OP_423J2_125_3477_n634), .CI(DP_OP_423J2_125_3477_n503), .CO(
        DP_OP_423J2_125_3477_n486), .S(DP_OP_423J2_125_3477_n487) );
  FADDX1_HVT DP_OP_423J2_125_3477_U399 ( .A(DP_OP_423J2_125_3477_n632), .B(
        DP_OP_423J2_125_3477_n501), .CI(DP_OP_423J2_125_3477_n499), .CO(
        DP_OP_423J2_125_3477_n484), .S(DP_OP_423J2_125_3477_n485) );
  FADDX1_HVT DP_OP_423J2_125_3477_U398 ( .A(DP_OP_423J2_125_3477_n630), .B(
        DP_OP_423J2_125_3477_n497), .CI(DP_OP_423J2_125_3477_n628), .CO(
        DP_OP_423J2_125_3477_n482), .S(DP_OP_423J2_125_3477_n483) );
  FADDX1_HVT DP_OP_423J2_125_3477_U397 ( .A(DP_OP_423J2_125_3477_n495), .B(
        DP_OP_423J2_125_3477_n626), .CI(DP_OP_423J2_125_3477_n493), .CO(
        DP_OP_423J2_125_3477_n480), .S(DP_OP_423J2_125_3477_n481) );
  FADDX1_HVT DP_OP_423J2_125_3477_U396 ( .A(DP_OP_423J2_125_3477_n624), .B(
        DP_OP_423J2_125_3477_n622), .CI(DP_OP_423J2_125_3477_n491), .CO(
        DP_OP_423J2_125_3477_n478), .S(DP_OP_423J2_125_3477_n479) );
  FADDX1_HVT DP_OP_423J2_125_3477_U395 ( .A(DP_OP_423J2_125_3477_n620), .B(
        DP_OP_423J2_125_3477_n489), .CI(DP_OP_423J2_125_3477_n487), .CO(
        DP_OP_423J2_125_3477_n476), .S(DP_OP_423J2_125_3477_n477) );
  FADDX1_HVT DP_OP_423J2_125_3477_U394 ( .A(DP_OP_423J2_125_3477_n618), .B(
        DP_OP_423J2_125_3477_n485), .CI(DP_OP_423J2_125_3477_n616), .CO(
        DP_OP_423J2_125_3477_n474), .S(DP_OP_423J2_125_3477_n475) );
  FADDX1_HVT DP_OP_423J2_125_3477_U393 ( .A(DP_OP_423J2_125_3477_n483), .B(
        DP_OP_423J2_125_3477_n614), .CI(DP_OP_423J2_125_3477_n481), .CO(
        DP_OP_423J2_125_3477_n472), .S(DP_OP_423J2_125_3477_n473) );
  FADDX1_HVT DP_OP_423J2_125_3477_U392 ( .A(DP_OP_423J2_125_3477_n612), .B(
        DP_OP_423J2_125_3477_n479), .CI(DP_OP_423J2_125_3477_n610), .CO(
        DP_OP_423J2_125_3477_n470), .S(DP_OP_423J2_125_3477_n471) );
  FADDX1_HVT DP_OP_423J2_125_3477_U391 ( .A(DP_OP_423J2_125_3477_n477), .B(
        DP_OP_423J2_125_3477_n608), .CI(DP_OP_423J2_125_3477_n475), .CO(
        DP_OP_423J2_125_3477_n468), .S(DP_OP_423J2_125_3477_n469) );
  FADDX1_HVT DP_OP_423J2_125_3477_U390 ( .A(DP_OP_423J2_125_3477_n606), .B(
        DP_OP_423J2_125_3477_n473), .CI(DP_OP_423J2_125_3477_n604), .CO(
        DP_OP_423J2_125_3477_n466), .S(DP_OP_423J2_125_3477_n467) );
  FADDX1_HVT DP_OP_423J2_125_3477_U389 ( .A(DP_OP_423J2_125_3477_n471), .B(
        DP_OP_423J2_125_3477_n469), .CI(DP_OP_423J2_125_3477_n602), .CO(
        DP_OP_423J2_125_3477_n464), .S(DP_OP_423J2_125_3477_n465) );
  FADDX1_HVT DP_OP_423J2_125_3477_U388 ( .A(DP_OP_423J2_125_3477_n600), .B(
        DP_OP_423J2_125_3477_n467), .CI(DP_OP_423J2_125_3477_n465), .CO(
        DP_OP_423J2_125_3477_n462), .S(DP_OP_423J2_125_3477_n463) );
  FADDX1_HVT DP_OP_423J2_125_3477_U386 ( .A(DP_OP_423J2_125_3477_n2976), .B(
        DP_OP_423J2_125_3477_n1920), .CI(DP_OP_423J2_125_3477_n461), .CO(
        DP_OP_423J2_125_3477_n458), .S(DP_OP_423J2_125_3477_n459) );
  FADDX1_HVT DP_OP_423J2_125_3477_U385 ( .A(DP_OP_423J2_125_3477_n2008), .B(
        DP_OP_423J2_125_3477_n2932), .CI(DP_OP_423J2_125_3477_n2360), .CO(
        DP_OP_423J2_125_3477_n456), .S(DP_OP_423J2_125_3477_n457) );
  FADDX1_HVT DP_OP_423J2_125_3477_U384 ( .A(DP_OP_423J2_125_3477_n2492), .B(
        DP_OP_423J2_125_3477_n2888), .CI(DP_OP_423J2_125_3477_n2844), .CO(
        DP_OP_423J2_125_3477_n454), .S(DP_OP_423J2_125_3477_n455) );
  FADDX1_HVT DP_OP_423J2_125_3477_U383 ( .A(DP_OP_423J2_125_3477_n2316), .B(
        DP_OP_423J2_125_3477_n2800), .CI(DP_OP_423J2_125_3477_n2756), .CO(
        DP_OP_423J2_125_3477_n452), .S(DP_OP_423J2_125_3477_n453) );
  FADDX1_HVT DP_OP_423J2_125_3477_U382 ( .A(DP_OP_423J2_125_3477_n2184), .B(
        DP_OP_423J2_125_3477_n1964), .CI(DP_OP_423J2_125_3477_n2712), .CO(
        DP_OP_423J2_125_3477_n450), .S(DP_OP_423J2_125_3477_n451) );
  FADDX1_HVT DP_OP_423J2_125_3477_U381 ( .A(DP_OP_423J2_125_3477_n2668), .B(
        DP_OP_423J2_125_3477_n2624), .CI(DP_OP_423J2_125_3477_n2580), .CO(
        DP_OP_423J2_125_3477_n448), .S(DP_OP_423J2_125_3477_n449) );
  FADDX1_HVT DP_OP_423J2_125_3477_U380 ( .A(DP_OP_423J2_125_3477_n2228), .B(
        DP_OP_423J2_125_3477_n2052), .CI(DP_OP_423J2_125_3477_n2096), .CO(
        DP_OP_423J2_125_3477_n446), .S(DP_OP_423J2_125_3477_n447) );
  FADDX1_HVT DP_OP_423J2_125_3477_U379 ( .A(DP_OP_423J2_125_3477_n2140), .B(
        DP_OP_423J2_125_3477_n2536), .CI(DP_OP_423J2_125_3477_n2448), .CO(
        DP_OP_423J2_125_3477_n444), .S(DP_OP_423J2_125_3477_n445) );
  FADDX1_HVT DP_OP_423J2_125_3477_U378 ( .A(DP_OP_423J2_125_3477_n2272), .B(
        DP_OP_423J2_125_3477_n2404), .CI(DP_OP_423J2_125_3477_n596), .CO(
        DP_OP_423J2_125_3477_n442), .S(DP_OP_423J2_125_3477_n443) );
  FADDX1_HVT DP_OP_423J2_125_3477_U377 ( .A(DP_OP_423J2_125_3477_n594), .B(
        DP_OP_423J2_125_3477_n564), .CI(DP_OP_423J2_125_3477_n592), .CO(
        DP_OP_423J2_125_3477_n440), .S(DP_OP_423J2_125_3477_n441) );
  FADDX1_HVT DP_OP_423J2_125_3477_U376 ( .A(DP_OP_423J2_125_3477_n590), .B(
        DP_OP_423J2_125_3477_n566), .CI(DP_OP_423J2_125_3477_n568), .CO(
        DP_OP_423J2_125_3477_n438), .S(DP_OP_423J2_125_3477_n439) );
  FADDX1_HVT DP_OP_423J2_125_3477_U375 ( .A(DP_OP_423J2_125_3477_n588), .B(
        DP_OP_423J2_125_3477_n570), .CI(DP_OP_423J2_125_3477_n572), .CO(
        DP_OP_423J2_125_3477_n436), .S(DP_OP_423J2_125_3477_n437) );
  FADDX1_HVT DP_OP_423J2_125_3477_U374 ( .A(DP_OP_423J2_125_3477_n586), .B(
        DP_OP_423J2_125_3477_n574), .CI(DP_OP_423J2_125_3477_n576), .CO(
        DP_OP_423J2_125_3477_n434), .S(DP_OP_423J2_125_3477_n435) );
  FADDX1_HVT DP_OP_423J2_125_3477_U373 ( .A(DP_OP_423J2_125_3477_n584), .B(
        DP_OP_423J2_125_3477_n578), .CI(DP_OP_423J2_125_3477_n580), .CO(
        DP_OP_423J2_125_3477_n432), .S(DP_OP_423J2_125_3477_n433) );
  FADDX1_HVT DP_OP_423J2_125_3477_U372 ( .A(DP_OP_423J2_125_3477_n582), .B(
        DP_OP_423J2_125_3477_n459), .CI(DP_OP_423J2_125_3477_n455), .CO(
        DP_OP_423J2_125_3477_n430), .S(DP_OP_423J2_125_3477_n431) );
  FADDX1_HVT DP_OP_423J2_125_3477_U371 ( .A(DP_OP_423J2_125_3477_n451), .B(
        DP_OP_423J2_125_3477_n445), .CI(DP_OP_423J2_125_3477_n447), .CO(
        DP_OP_423J2_125_3477_n428), .S(DP_OP_423J2_125_3477_n429) );
  FADDX1_HVT DP_OP_423J2_125_3477_U370 ( .A(DP_OP_423J2_125_3477_n449), .B(
        DP_OP_423J2_125_3477_n457), .CI(DP_OP_423J2_125_3477_n453), .CO(
        DP_OP_423J2_125_3477_n426), .S(DP_OP_423J2_125_3477_n427) );
  FADDX1_HVT DP_OP_423J2_125_3477_U369 ( .A(DP_OP_423J2_125_3477_n562), .B(
        DP_OP_423J2_125_3477_n560), .CI(DP_OP_423J2_125_3477_n552), .CO(
        DP_OP_423J2_125_3477_n424), .S(DP_OP_423J2_125_3477_n425) );
  FADDX1_HVT DP_OP_423J2_125_3477_U368 ( .A(DP_OP_423J2_125_3477_n558), .B(
        DP_OP_423J2_125_3477_n554), .CI(DP_OP_423J2_125_3477_n556), .CO(
        DP_OP_423J2_125_3477_n422), .S(DP_OP_423J2_125_3477_n423) );
  FADDX1_HVT DP_OP_423J2_125_3477_U367 ( .A(DP_OP_423J2_125_3477_n550), .B(
        DP_OP_423J2_125_3477_n546), .CI(DP_OP_423J2_125_3477_n443), .CO(
        DP_OP_423J2_125_3477_n420), .S(DP_OP_423J2_125_3477_n421) );
  FADDX1_HVT DP_OP_423J2_125_3477_U366 ( .A(DP_OP_423J2_125_3477_n548), .B(
        DP_OP_423J2_125_3477_n544), .CI(DP_OP_423J2_125_3477_n441), .CO(
        DP_OP_423J2_125_3477_n418), .S(DP_OP_423J2_125_3477_n419) );
  FADDX1_HVT DP_OP_423J2_125_3477_U365 ( .A(DP_OP_423J2_125_3477_n542), .B(
        DP_OP_423J2_125_3477_n435), .CI(DP_OP_423J2_125_3477_n437), .CO(
        DP_OP_423J2_125_3477_n416), .S(DP_OP_423J2_125_3477_n417) );
  FADDX1_HVT DP_OP_423J2_125_3477_U364 ( .A(DP_OP_423J2_125_3477_n540), .B(
        DP_OP_423J2_125_3477_n439), .CI(DP_OP_423J2_125_3477_n433), .CO(
        DP_OP_423J2_125_3477_n414), .S(DP_OP_423J2_125_3477_n415) );
  FADDX1_HVT DP_OP_423J2_125_3477_U363 ( .A(DP_OP_423J2_125_3477_n538), .B(
        DP_OP_423J2_125_3477_n536), .CI(DP_OP_423J2_125_3477_n534), .CO(
        DP_OP_423J2_125_3477_n412), .S(DP_OP_423J2_125_3477_n413) );
  FADDX1_HVT DP_OP_423J2_125_3477_U362 ( .A(DP_OP_423J2_125_3477_n431), .B(
        DP_OP_423J2_125_3477_n427), .CI(DP_OP_423J2_125_3477_n532), .CO(
        DP_OP_423J2_125_3477_n410), .S(DP_OP_423J2_125_3477_n411) );
  FADDX1_HVT DP_OP_423J2_125_3477_U361 ( .A(DP_OP_423J2_125_3477_n429), .B(
        DP_OP_423J2_125_3477_n530), .CI(DP_OP_423J2_125_3477_n528), .CO(
        DP_OP_423J2_125_3477_n408), .S(DP_OP_423J2_125_3477_n409) );
  FADDX1_HVT DP_OP_423J2_125_3477_U360 ( .A(DP_OP_423J2_125_3477_n526), .B(
        DP_OP_423J2_125_3477_n425), .CI(DP_OP_423J2_125_3477_n423), .CO(
        DP_OP_423J2_125_3477_n406), .S(DP_OP_423J2_125_3477_n407) );
  FADDX1_HVT DP_OP_423J2_125_3477_U359 ( .A(DP_OP_423J2_125_3477_n524), .B(
        DP_OP_423J2_125_3477_n520), .CI(DP_OP_423J2_125_3477_n518), .CO(
        DP_OP_423J2_125_3477_n404), .S(DP_OP_423J2_125_3477_n405) );
  FADDX1_HVT DP_OP_423J2_125_3477_U358 ( .A(DP_OP_423J2_125_3477_n522), .B(
        DP_OP_423J2_125_3477_n516), .CI(DP_OP_423J2_125_3477_n421), .CO(
        DP_OP_423J2_125_3477_n402), .S(DP_OP_423J2_125_3477_n403) );
  FADDX1_HVT DP_OP_423J2_125_3477_U357 ( .A(DP_OP_423J2_125_3477_n419), .B(
        DP_OP_423J2_125_3477_n514), .CI(DP_OP_423J2_125_3477_n512), .CO(
        DP_OP_423J2_125_3477_n400), .S(DP_OP_423J2_125_3477_n401) );
  FADDX1_HVT DP_OP_423J2_125_3477_U356 ( .A(DP_OP_423J2_125_3477_n417), .B(
        DP_OP_423J2_125_3477_n415), .CI(DP_OP_423J2_125_3477_n413), .CO(
        DP_OP_423J2_125_3477_n398), .S(DP_OP_423J2_125_3477_n399) );
  FADDX1_HVT DP_OP_423J2_125_3477_U355 ( .A(DP_OP_423J2_125_3477_n510), .B(
        DP_OP_423J2_125_3477_n508), .CI(DP_OP_423J2_125_3477_n411), .CO(
        DP_OP_423J2_125_3477_n396), .S(DP_OP_423J2_125_3477_n397) );
  FADDX1_HVT DP_OP_423J2_125_3477_U354 ( .A(DP_OP_423J2_125_3477_n506), .B(
        DP_OP_423J2_125_3477_n409), .CI(DP_OP_423J2_125_3477_n504), .CO(
        DP_OP_423J2_125_3477_n394), .S(DP_OP_423J2_125_3477_n395) );
  FADDX1_HVT DP_OP_423J2_125_3477_U353 ( .A(DP_OP_423J2_125_3477_n502), .B(
        DP_OP_423J2_125_3477_n407), .CI(DP_OP_423J2_125_3477_n500), .CO(
        DP_OP_423J2_125_3477_n392), .S(DP_OP_423J2_125_3477_n393) );
  FADDX1_HVT DP_OP_423J2_125_3477_U352 ( .A(DP_OP_423J2_125_3477_n498), .B(
        DP_OP_423J2_125_3477_n405), .CI(DP_OP_423J2_125_3477_n403), .CO(
        DP_OP_423J2_125_3477_n390), .S(DP_OP_423J2_125_3477_n391) );
  FADDX1_HVT DP_OP_423J2_125_3477_U351 ( .A(DP_OP_423J2_125_3477_n496), .B(
        DP_OP_423J2_125_3477_n401), .CI(DP_OP_423J2_125_3477_n494), .CO(
        DP_OP_423J2_125_3477_n388), .S(DP_OP_423J2_125_3477_n389) );
  FADDX1_HVT DP_OP_423J2_125_3477_U350 ( .A(DP_OP_423J2_125_3477_n399), .B(
        DP_OP_423J2_125_3477_n492), .CI(DP_OP_423J2_125_3477_n490), .CO(
        DP_OP_423J2_125_3477_n386), .S(DP_OP_423J2_125_3477_n387) );
  FADDX1_HVT DP_OP_423J2_125_3477_U349 ( .A(DP_OP_423J2_125_3477_n397), .B(
        DP_OP_423J2_125_3477_n488), .CI(DP_OP_423J2_125_3477_n395), .CO(
        DP_OP_423J2_125_3477_n384), .S(DP_OP_423J2_125_3477_n385) );
  FADDX1_HVT DP_OP_423J2_125_3477_U348 ( .A(DP_OP_423J2_125_3477_n486), .B(
        DP_OP_423J2_125_3477_n393), .CI(DP_OP_423J2_125_3477_n484), .CO(
        DP_OP_423J2_125_3477_n382), .S(DP_OP_423J2_125_3477_n383) );
  FADDX1_HVT DP_OP_423J2_125_3477_U347 ( .A(DP_OP_423J2_125_3477_n391), .B(
        DP_OP_423J2_125_3477_n482), .CI(DP_OP_423J2_125_3477_n389), .CO(
        DP_OP_423J2_125_3477_n380), .S(DP_OP_423J2_125_3477_n381) );
  FADDX1_HVT DP_OP_423J2_125_3477_U346 ( .A(DP_OP_423J2_125_3477_n480), .B(
        DP_OP_423J2_125_3477_n387), .CI(DP_OP_423J2_125_3477_n478), .CO(
        DP_OP_423J2_125_3477_n378), .S(DP_OP_423J2_125_3477_n379) );
  FADDX1_HVT DP_OP_423J2_125_3477_U345 ( .A(DP_OP_423J2_125_3477_n385), .B(
        DP_OP_423J2_125_3477_n476), .CI(DP_OP_423J2_125_3477_n383), .CO(
        DP_OP_423J2_125_3477_n376), .S(DP_OP_423J2_125_3477_n377) );
  FADDX1_HVT DP_OP_423J2_125_3477_U344 ( .A(DP_OP_423J2_125_3477_n474), .B(
        DP_OP_423J2_125_3477_n381), .CI(DP_OP_423J2_125_3477_n472), .CO(
        DP_OP_423J2_125_3477_n374), .S(DP_OP_423J2_125_3477_n375) );
  FADDX1_HVT DP_OP_423J2_125_3477_U343 ( .A(DP_OP_423J2_125_3477_n379), .B(
        DP_OP_423J2_125_3477_n470), .CI(DP_OP_423J2_125_3477_n377), .CO(
        DP_OP_423J2_125_3477_n372), .S(DP_OP_423J2_125_3477_n373) );
  FADDX1_HVT DP_OP_423J2_125_3477_U342 ( .A(DP_OP_423J2_125_3477_n468), .B(
        DP_OP_423J2_125_3477_n375), .CI(DP_OP_423J2_125_3477_n466), .CO(
        DP_OP_423J2_125_3477_n370), .S(DP_OP_423J2_125_3477_n371) );
  FADDX1_HVT DP_OP_423J2_125_3477_U341 ( .A(DP_OP_423J2_125_3477_n373), .B(
        DP_OP_423J2_125_3477_n464), .CI(DP_OP_423J2_125_3477_n371), .CO(
        DP_OP_423J2_125_3477_n368), .S(DP_OP_423J2_125_3477_n369) );
  FADDX1_HVT DP_OP_423J2_125_3477_U340 ( .A(DP_OP_423J2_125_3477_n1876), .B(
        DP_OP_423J2_125_3477_n460), .CI(DP_OP_423J2_125_3477_n458), .CO(
        DP_OP_423J2_125_3477_n366), .S(DP_OP_423J2_125_3477_n367) );
  FADDX1_HVT DP_OP_423J2_125_3477_U339 ( .A(DP_OP_423J2_125_3477_n448), .B(
        DP_OP_423J2_125_3477_n444), .CI(DP_OP_423J2_125_3477_n456), .CO(
        DP_OP_423J2_125_3477_n364), .S(DP_OP_423J2_125_3477_n365) );
  FADDX1_HVT DP_OP_423J2_125_3477_U338 ( .A(DP_OP_423J2_125_3477_n454), .B(
        DP_OP_423J2_125_3477_n452), .CI(DP_OP_423J2_125_3477_n450), .CO(
        DP_OP_423J2_125_3477_n362), .S(DP_OP_423J2_125_3477_n363) );
  FADDX1_HVT DP_OP_423J2_125_3477_U337 ( .A(DP_OP_423J2_125_3477_n446), .B(
        DP_OP_423J2_125_3477_n442), .CI(DP_OP_423J2_125_3477_n440), .CO(
        DP_OP_423J2_125_3477_n360), .S(DP_OP_423J2_125_3477_n361) );
  FADDX1_HVT DP_OP_423J2_125_3477_U336 ( .A(DP_OP_423J2_125_3477_n438), .B(
        DP_OP_423J2_125_3477_n436), .CI(DP_OP_423J2_125_3477_n434), .CO(
        DP_OP_423J2_125_3477_n358), .S(DP_OP_423J2_125_3477_n359) );
  FADDX1_HVT DP_OP_423J2_125_3477_U335 ( .A(DP_OP_423J2_125_3477_n432), .B(
        DP_OP_423J2_125_3477_n367), .CI(DP_OP_423J2_125_3477_n430), .CO(
        DP_OP_423J2_125_3477_n356), .S(DP_OP_423J2_125_3477_n357) );
  FADDX1_HVT DP_OP_423J2_125_3477_U334 ( .A(DP_OP_423J2_125_3477_n428), .B(
        DP_OP_423J2_125_3477_n363), .CI(DP_OP_423J2_125_3477_n365), .CO(
        DP_OP_423J2_125_3477_n354), .S(DP_OP_423J2_125_3477_n355) );
  FADDX1_HVT DP_OP_423J2_125_3477_U333 ( .A(DP_OP_423J2_125_3477_n426), .B(
        DP_OP_423J2_125_3477_n424), .CI(DP_OP_423J2_125_3477_n422), .CO(
        DP_OP_423J2_125_3477_n352), .S(DP_OP_423J2_125_3477_n353) );
  FADDX1_HVT DP_OP_423J2_125_3477_U332 ( .A(DP_OP_423J2_125_3477_n420), .B(
        DP_OP_423J2_125_3477_n361), .CI(DP_OP_423J2_125_3477_n418), .CO(
        DP_OP_423J2_125_3477_n350), .S(DP_OP_423J2_125_3477_n351) );
  FADDX1_HVT DP_OP_423J2_125_3477_U331 ( .A(DP_OP_423J2_125_3477_n416), .B(
        DP_OP_423J2_125_3477_n359), .CI(DP_OP_423J2_125_3477_n414), .CO(
        DP_OP_423J2_125_3477_n348), .S(DP_OP_423J2_125_3477_n349) );
  FADDX1_HVT DP_OP_423J2_125_3477_U330 ( .A(DP_OP_423J2_125_3477_n412), .B(
        DP_OP_423J2_125_3477_n357), .CI(DP_OP_423J2_125_3477_n410), .CO(
        DP_OP_423J2_125_3477_n346), .S(DP_OP_423J2_125_3477_n347) );
  FADDX1_HVT DP_OP_423J2_125_3477_U329 ( .A(DP_OP_423J2_125_3477_n355), .B(
        DP_OP_423J2_125_3477_n408), .CI(DP_OP_423J2_125_3477_n406), .CO(
        DP_OP_423J2_125_3477_n344), .S(DP_OP_423J2_125_3477_n345) );
  FADDX1_HVT DP_OP_423J2_125_3477_U328 ( .A(DP_OP_423J2_125_3477_n353), .B(
        DP_OP_423J2_125_3477_n404), .CI(DP_OP_423J2_125_3477_n402), .CO(
        DP_OP_423J2_125_3477_n342), .S(DP_OP_423J2_125_3477_n343) );
  FADDX1_HVT DP_OP_423J2_125_3477_U327 ( .A(DP_OP_423J2_125_3477_n351), .B(
        DP_OP_423J2_125_3477_n400), .CI(DP_OP_423J2_125_3477_n349), .CO(
        DP_OP_423J2_125_3477_n340), .S(DP_OP_423J2_125_3477_n341) );
  FADDX1_HVT DP_OP_423J2_125_3477_U326 ( .A(DP_OP_423J2_125_3477_n398), .B(
        DP_OP_423J2_125_3477_n347), .CI(DP_OP_423J2_125_3477_n396), .CO(
        DP_OP_423J2_125_3477_n338), .S(DP_OP_423J2_125_3477_n339) );
  FADDX1_HVT DP_OP_423J2_125_3477_U325 ( .A(DP_OP_423J2_125_3477_n394), .B(
        DP_OP_423J2_125_3477_n345), .CI(DP_OP_423J2_125_3477_n392), .CO(
        DP_OP_423J2_125_3477_n336), .S(DP_OP_423J2_125_3477_n337) );
  FADDX1_HVT DP_OP_423J2_125_3477_U324 ( .A(DP_OP_423J2_125_3477_n343), .B(
        DP_OP_423J2_125_3477_n390), .CI(DP_OP_423J2_125_3477_n388), .CO(
        DP_OP_423J2_125_3477_n334), .S(DP_OP_423J2_125_3477_n335) );
  FADDX1_HVT DP_OP_423J2_125_3477_U323 ( .A(DP_OP_423J2_125_3477_n341), .B(
        DP_OP_423J2_125_3477_n386), .CI(DP_OP_423J2_125_3477_n339), .CO(
        DP_OP_423J2_125_3477_n332), .S(DP_OP_423J2_125_3477_n333) );
  FADDX1_HVT DP_OP_423J2_125_3477_U322 ( .A(DP_OP_423J2_125_3477_n384), .B(
        DP_OP_423J2_125_3477_n337), .CI(DP_OP_423J2_125_3477_n382), .CO(
        DP_OP_423J2_125_3477_n330), .S(DP_OP_423J2_125_3477_n331) );
  FADDX1_HVT DP_OP_423J2_125_3477_U321 ( .A(DP_OP_423J2_125_3477_n380), .B(
        DP_OP_423J2_125_3477_n335), .CI(DP_OP_423J2_125_3477_n333), .CO(
        DP_OP_423J2_125_3477_n328), .S(DP_OP_423J2_125_3477_n329) );
  FADDX1_HVT DP_OP_423J2_125_3477_U320 ( .A(DP_OP_423J2_125_3477_n378), .B(
        DP_OP_423J2_125_3477_n331), .CI(DP_OP_423J2_125_3477_n376), .CO(
        DP_OP_423J2_125_3477_n326), .S(DP_OP_423J2_125_3477_n327) );
  FADDX1_HVT DP_OP_423J2_125_3477_U319 ( .A(DP_OP_423J2_125_3477_n374), .B(
        DP_OP_423J2_125_3477_n329), .CI(DP_OP_423J2_125_3477_n372), .CO(
        DP_OP_423J2_125_3477_n324), .S(DP_OP_423J2_125_3477_n325) );
  FADDX1_HVT DP_OP_423J2_125_3477_U318 ( .A(DP_OP_423J2_125_3477_n327), .B(
        DP_OP_423J2_125_3477_n370), .CI(DP_OP_423J2_125_3477_n325), .CO(
        DP_OP_423J2_125_3477_n322), .S(DP_OP_423J2_125_3477_n323) );
  FADDX1_HVT DP_OP_423J2_125_3477_U317 ( .A(DP_OP_423J2_125_3477_n1875), .B(
        DP_OP_423J2_125_3477_n366), .CI(DP_OP_423J2_125_3477_n364), .CO(
        DP_OP_423J2_125_3477_n320), .S(DP_OP_423J2_125_3477_n321) );
  FADDX1_HVT DP_OP_423J2_125_3477_U316 ( .A(DP_OP_423J2_125_3477_n362), .B(
        DP_OP_423J2_125_3477_n360), .CI(DP_OP_423J2_125_3477_n358), .CO(
        DP_OP_423J2_125_3477_n318), .S(DP_OP_423J2_125_3477_n319) );
  FADDX1_HVT DP_OP_423J2_125_3477_U315 ( .A(DP_OP_423J2_125_3477_n356), .B(
        DP_OP_423J2_125_3477_n321), .CI(DP_OP_423J2_125_3477_n354), .CO(
        DP_OP_423J2_125_3477_n316), .S(DP_OP_423J2_125_3477_n317) );
  FADDX1_HVT DP_OP_423J2_125_3477_U314 ( .A(DP_OP_423J2_125_3477_n352), .B(
        DP_OP_423J2_125_3477_n350), .CI(DP_OP_423J2_125_3477_n319), .CO(
        DP_OP_423J2_125_3477_n314), .S(DP_OP_423J2_125_3477_n315) );
  FADDX1_HVT DP_OP_423J2_125_3477_U313 ( .A(DP_OP_423J2_125_3477_n348), .B(
        DP_OP_423J2_125_3477_n346), .CI(DP_OP_423J2_125_3477_n317), .CO(
        DP_OP_423J2_125_3477_n312), .S(DP_OP_423J2_125_3477_n313) );
  FADDX1_HVT DP_OP_423J2_125_3477_U312 ( .A(DP_OP_423J2_125_3477_n344), .B(
        DP_OP_423J2_125_3477_n342), .CI(DP_OP_423J2_125_3477_n315), .CO(
        DP_OP_423J2_125_3477_n310), .S(DP_OP_423J2_125_3477_n311) );
  FADDX1_HVT DP_OP_423J2_125_3477_U311 ( .A(DP_OP_423J2_125_3477_n340), .B(
        DP_OP_423J2_125_3477_n313), .CI(DP_OP_423J2_125_3477_n338), .CO(
        DP_OP_423J2_125_3477_n308), .S(DP_OP_423J2_125_3477_n309) );
  FADDX1_HVT DP_OP_423J2_125_3477_U310 ( .A(DP_OP_423J2_125_3477_n336), .B(
        DP_OP_423J2_125_3477_n311), .CI(DP_OP_423J2_125_3477_n334), .CO(
        DP_OP_423J2_125_3477_n306), .S(DP_OP_423J2_125_3477_n307) );
  FADDX1_HVT DP_OP_423J2_125_3477_U309 ( .A(DP_OP_423J2_125_3477_n332), .B(
        DP_OP_423J2_125_3477_n309), .CI(DP_OP_423J2_125_3477_n330), .CO(
        DP_OP_423J2_125_3477_n304), .S(DP_OP_423J2_125_3477_n305) );
  FADDX1_HVT DP_OP_423J2_125_3477_U308 ( .A(DP_OP_423J2_125_3477_n307), .B(
        DP_OP_423J2_125_3477_n328), .CI(DP_OP_423J2_125_3477_n305), .CO(
        DP_OP_423J2_125_3477_n302), .S(DP_OP_423J2_125_3477_n303) );
  FADDX1_HVT DP_OP_423J2_125_3477_U307 ( .A(DP_OP_423J2_125_3477_n326), .B(
        DP_OP_423J2_125_3477_n324), .CI(DP_OP_423J2_125_3477_n303), .CO(
        DP_OP_423J2_125_3477_n300), .S(DP_OP_423J2_125_3477_n301) );
  FADDX1_HVT DP_OP_423J2_125_3477_U306 ( .A(DP_OP_423J2_125_3477_n1874), .B(
        DP_OP_423J2_125_3477_n320), .CI(DP_OP_423J2_125_3477_n318), .CO(
        DP_OP_423J2_125_3477_n298), .S(DP_OP_423J2_125_3477_n299) );
  FADDX1_HVT DP_OP_423J2_125_3477_U305 ( .A(DP_OP_423J2_125_3477_n316), .B(
        DP_OP_423J2_125_3477_n299), .CI(DP_OP_423J2_125_3477_n314), .CO(
        DP_OP_423J2_125_3477_n296), .S(DP_OP_423J2_125_3477_n297) );
  FADDX1_HVT DP_OP_423J2_125_3477_U304 ( .A(DP_OP_423J2_125_3477_n312), .B(
        DP_OP_423J2_125_3477_n310), .CI(DP_OP_423J2_125_3477_n297), .CO(
        DP_OP_423J2_125_3477_n294), .S(DP_OP_423J2_125_3477_n295) );
  FADDX1_HVT DP_OP_423J2_125_3477_U303 ( .A(DP_OP_423J2_125_3477_n308), .B(
        DP_OP_423J2_125_3477_n295), .CI(DP_OP_423J2_125_3477_n306), .CO(
        DP_OP_423J2_125_3477_n292), .S(DP_OP_423J2_125_3477_n293) );
  FADDX1_HVT DP_OP_423J2_125_3477_U302 ( .A(DP_OP_423J2_125_3477_n304), .B(
        DP_OP_423J2_125_3477_n293), .CI(DP_OP_423J2_125_3477_n302), .CO(
        DP_OP_423J2_125_3477_n290), .S(DP_OP_423J2_125_3477_n291) );
  FADDX1_HVT DP_OP_423J2_125_3477_U300 ( .A(DP_OP_423J2_125_3477_n289), .B(
        DP_OP_423J2_125_3477_n298), .CI(DP_OP_423J2_125_3477_n296), .CO(
        DP_OP_423J2_125_3477_n286), .S(DP_OP_423J2_125_3477_n287) );
  FADDX1_HVT DP_OP_423J2_125_3477_U299 ( .A(DP_OP_423J2_125_3477_n287), .B(
        DP_OP_423J2_125_3477_n294), .CI(DP_OP_423J2_125_3477_n292), .CO(
        DP_OP_423J2_125_3477_n284), .S(DP_OP_423J2_125_3477_n285) );
  FADDX1_HVT DP_OP_423J2_125_3477_U298 ( .A(DP_OP_423J2_125_3477_n1873), .B(
        DP_OP_423J2_125_3477_n288), .CI(DP_OP_423J2_125_3477_n286), .CO(
        DP_OP_423J2_125_3477_n282), .S(DP_OP_423J2_125_3477_n283) );
  FADDX1_HVT DP_OP_423J2_125_3477_U281 ( .A(DP_OP_423J2_125_3477_n1853), .B(
        DP_OP_423J2_125_3477_n1851), .CI(DP_OP_423J2_125_3477_n1849), .CO(
        DP_OP_423J2_125_3477_n219), .S(n_conv2_sum_b[0]) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U280 ( .A1(DP_OP_423J2_125_3477_n1787), 
        .A2(DP_OP_423J2_125_3477_n1789), .Y(DP_OP_423J2_125_3477_n218) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U279 ( .A1(DP_OP_423J2_125_3477_n1789), .A2(
        DP_OP_423J2_125_3477_n1787), .Y(DP_OP_423J2_125_3477_n217) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U273 ( .A1(DP_OP_423J2_125_3477_n1681), 
        .A2(DP_OP_423J2_125_3477_n1683), .Y(DP_OP_423J2_125_3477_n215) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U265 ( .A1(DP_OP_423J2_125_3477_n1527), 
        .A2(DP_OP_423J2_125_3477_n1529), .Y(DP_OP_423J2_125_3477_n210) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U264 ( .A1(DP_OP_423J2_125_3477_n1529), .A2(
        DP_OP_423J2_125_3477_n1527), .Y(DP_OP_423J2_125_3477_n209) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U259 ( .A1(DP_OP_423J2_125_3477_n1351), 
        .A2(DP_OP_423J2_125_3477_n1353), .Y(DP_OP_423J2_125_3477_n207) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U251 ( .A1(DP_OP_423J2_125_3477_n1163), 
        .A2(DP_OP_423J2_125_3477_n1165), .Y(DP_OP_423J2_125_3477_n202) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U250 ( .A1(DP_OP_423J2_125_3477_n1165), .A2(
        DP_OP_423J2_125_3477_n1163), .Y(DP_OP_423J2_125_3477_n201) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U245 ( .A1(DP_OP_423J2_125_3477_n969), .A2(
        DP_OP_423J2_125_3477_n971), .Y(DP_OP_423J2_125_3477_n199) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U237 ( .A1(DP_OP_423J2_125_3477_n773), .A2(
        DP_OP_423J2_125_3477_n968), .Y(DP_OP_423J2_125_3477_n194) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U236 ( .A1(DP_OP_423J2_125_3477_n968), .A2(
        DP_OP_423J2_125_3477_n773), .Y(DP_OP_423J2_125_3477_n193) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U230 ( .A1(DP_OP_423J2_125_3477_n599), .A2(
        DP_OP_423J2_125_3477_n772), .Y(DP_OP_423J2_125_3477_n190) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U229 ( .A1(DP_OP_423J2_125_3477_n772), .A2(
        DP_OP_423J2_125_3477_n599), .Y(DP_OP_423J2_125_3477_n189) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U224 ( .A1(DP_OP_423J2_125_3477_n463), .A2(
        DP_OP_423J2_125_3477_n598), .Y(DP_OP_423J2_125_3477_n187) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U223 ( .A1(DP_OP_423J2_125_3477_n598), .A2(
        DP_OP_423J2_125_3477_n463), .Y(DP_OP_423J2_125_3477_n186) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U219 ( .A1(DP_OP_423J2_125_3477_n189), .A2(
        DP_OP_423J2_125_3477_n186), .Y(DP_OP_423J2_125_3477_n184) );
  AOI21X1_HVT DP_OP_423J2_125_3477_U218 ( .A1(DP_OP_423J2_125_3477_n184), .A2(
        DP_OP_423J2_125_3477_n192), .A3(DP_OP_423J2_125_3477_n185), .Y(
        DP_OP_423J2_125_3477_n183) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U215 ( .A1(DP_OP_423J2_125_3477_n369), .A2(
        DP_OP_423J2_125_3477_n462), .Y(DP_OP_423J2_125_3477_n181) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U214 ( .A1(DP_OP_423J2_125_3477_n462), .A2(
        DP_OP_423J2_125_3477_n369), .Y(DP_OP_423J2_125_3477_n180) );
  AOI21X1_HVT DP_OP_423J2_125_3477_U209 ( .A1(DP_OP_423J2_125_3477_n182), .A2(
        DP_OP_423J2_125_3477_n241), .A3(DP_OP_423J2_125_3477_n179), .Y(
        DP_OP_423J2_125_3477_n177) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U207 ( .A1(DP_OP_423J2_125_3477_n323), .A2(
        DP_OP_423J2_125_3477_n368), .Y(DP_OP_423J2_125_3477_n176) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U206 ( .A1(DP_OP_423J2_125_3477_n368), .A2(
        DP_OP_423J2_125_3477_n323), .Y(DP_OP_423J2_125_3477_n175) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U204 ( .A1(DP_OP_423J2_125_3477_n240), .A2(
        DP_OP_423J2_125_3477_n176), .Y(DP_OP_423J2_125_3477_n25) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U202 ( .A1(DP_OP_423J2_125_3477_n175), .A2(
        DP_OP_423J2_125_3477_n180), .Y(DP_OP_423J2_125_3477_n173) );
  AOI21X1_HVT DP_OP_423J2_125_3477_U201 ( .A1(DP_OP_423J2_125_3477_n182), .A2(
        DP_OP_423J2_125_3477_n173), .A3(DP_OP_423J2_125_3477_n174), .Y(
        DP_OP_423J2_125_3477_n172) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U199 ( .A1(DP_OP_423J2_125_3477_n301), .A2(
        DP_OP_423J2_125_3477_n322), .Y(DP_OP_423J2_125_3477_n171) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U198 ( .A1(DP_OP_423J2_125_3477_n322), .A2(
        DP_OP_423J2_125_3477_n301), .Y(DP_OP_423J2_125_3477_n170) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U193 ( .A1(DP_OP_423J2_125_3477_n300), .A2(
        DP_OP_423J2_125_3477_n291), .Y(DP_OP_423J2_125_3477_n168) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U192 ( .A1(DP_OP_423J2_125_3477_n291), .A2(
        DP_OP_423J2_125_3477_n300), .Y(DP_OP_423J2_125_3477_n167) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U188 ( .A1(DP_OP_423J2_125_3477_n167), .A2(
        DP_OP_423J2_125_3477_n170), .Y(DP_OP_423J2_125_3477_n165) );
  AOI21X1_HVT DP_OP_423J2_125_3477_U187 ( .A1(DP_OP_423J2_125_3477_n174), .A2(
        DP_OP_423J2_125_3477_n165), .A3(DP_OP_423J2_125_3477_n166), .Y(
        DP_OP_423J2_125_3477_n164) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U186 ( .A1(DP_OP_423J2_125_3477_n173), .A2(
        DP_OP_423J2_125_3477_n165), .Y(DP_OP_423J2_125_3477_n163) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U182 ( .A1(DP_OP_423J2_125_3477_n290), .A2(
        DP_OP_423J2_125_3477_n285), .Y(DP_OP_423J2_125_3477_n152) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U181 ( .A1(DP_OP_423J2_125_3477_n285), .A2(
        DP_OP_423J2_125_3477_n290), .Y(DP_OP_423J2_125_3477_n151) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U168 ( .A1(DP_OP_423J2_125_3477_n284), .A2(
        DP_OP_423J2_125_3477_n283), .Y(DP_OP_423J2_125_3477_n149) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U167 ( .A1(DP_OP_423J2_125_3477_n283), .A2(
        DP_OP_423J2_125_3477_n284), .Y(DP_OP_423J2_125_3477_n148) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U161 ( .A1(DP_OP_423J2_125_3477_n237), .A2(
        DP_OP_423J2_125_3477_n236), .Y(DP_OP_423J2_125_3477_n144) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U156 ( .A1(DP_OP_423J2_125_3477_n282), .A2(
        DP_OP_423J2_125_3477_n281), .Y(DP_OP_423J2_125_3477_n140) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U153 ( .A1(DP_OP_423J2_125_3477_n235), .A2(
        DP_OP_423J2_125_3477_n140), .Y(DP_OP_423J2_125_3477_n20) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U146 ( .A1(DP_OP_423J2_125_3477_n279), .A2(
        DP_OP_423J2_125_3477_n280), .Y(DP_OP_423J2_125_3477_n133) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U145 ( .A1(DP_OP_423J2_125_3477_n280), .A2(
        DP_OP_423J2_125_3477_n279), .Y(DP_OP_423J2_125_3477_n132) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U143 ( .A1(DP_OP_423J2_125_3477_n234), .A2(
        DP_OP_423J2_125_3477_n133), .Y(DP_OP_423J2_125_3477_n19) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U140 ( .A1(DP_OP_423J2_125_3477_n277), .A2(
        DP_OP_423J2_125_3477_n278), .Y(DP_OP_423J2_125_3477_n130) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U139 ( .A1(DP_OP_423J2_125_3477_n278), .A2(
        DP_OP_423J2_125_3477_n277), .Y(DP_OP_423J2_125_3477_n129) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U137 ( .A1(DP_OP_423J2_125_3477_n233), .A2(
        DP_OP_423J2_125_3477_n130), .Y(DP_OP_423J2_125_3477_n18) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U135 ( .A1(DP_OP_423J2_125_3477_n129), .A2(
        DP_OP_423J2_125_3477_n132), .Y(DP_OP_423J2_125_3477_n127) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U130 ( .A1(DP_OP_423J2_125_3477_n275), .A2(
        DP_OP_423J2_125_3477_n276), .Y(DP_OP_423J2_125_3477_n123) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U127 ( .A1(n440), .A2(
        DP_OP_423J2_125_3477_n123), .Y(DP_OP_423J2_125_3477_n17) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U123 ( .A1(DP_OP_423J2_125_3477_n127), .A2(
        n440), .Y(DP_OP_423J2_125_3477_n118) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U120 ( .A1(DP_OP_423J2_125_3477_n273), .A2(
        DP_OP_423J2_125_3477_n274), .Y(DP_OP_423J2_125_3477_n116) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U119 ( .A1(DP_OP_423J2_125_3477_n274), .A2(
        DP_OP_423J2_125_3477_n273), .Y(DP_OP_423J2_125_3477_n115) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U110 ( .A1(DP_OP_423J2_125_3477_n271), .A2(
        DP_OP_423J2_125_3477_n272), .Y(DP_OP_423J2_125_3477_n109) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U103 ( .A1(DP_OP_423J2_125_3477_n113), .A2(
        n439), .Y(DP_OP_423J2_125_3477_n104) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U100 ( .A1(DP_OP_423J2_125_3477_n269), .A2(
        DP_OP_423J2_125_3477_n270), .Y(DP_OP_423J2_125_3477_n102) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U99 ( .A1(DP_OP_423J2_125_3477_n270), .A2(
        DP_OP_423J2_125_3477_n269), .Y(DP_OP_423J2_125_3477_n101) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U90 ( .A1(DP_OP_423J2_125_3477_n267), .A2(
        DP_OP_423J2_125_3477_n268), .Y(DP_OP_423J2_125_3477_n95) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U83 ( .A1(DP_OP_423J2_125_3477_n99), .A2(
        n435), .Y(DP_OP_423J2_125_3477_n90) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U80 ( .A1(DP_OP_423J2_125_3477_n265), .A2(
        DP_OP_423J2_125_3477_n266), .Y(DP_OP_423J2_125_3477_n88) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U79 ( .A1(DP_OP_423J2_125_3477_n266), .A2(
        DP_OP_423J2_125_3477_n265), .Y(DP_OP_423J2_125_3477_n87) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U70 ( .A1(DP_OP_423J2_125_3477_n263), .A2(
        DP_OP_423J2_125_3477_n264), .Y(DP_OP_423J2_125_3477_n81) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U63 ( .A1(DP_OP_423J2_125_3477_n85), .A2(
        n434), .Y(DP_OP_423J2_125_3477_n76) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U61 ( .A1(DP_OP_423J2_125_3477_n76), .A2(
        DP_OP_423J2_125_3477_n137), .Y(DP_OP_423J2_125_3477_n74) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U56 ( .A1(DP_OP_423J2_125_3477_n261), .A2(
        DP_OP_423J2_125_3477_n262), .Y(DP_OP_423J2_125_3477_n70) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U49 ( .A1(DP_OP_423J2_125_3477_n74), .A2(
        n433), .Y(DP_OP_423J2_125_3477_n65) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U45 ( .A1(DP_OP_423J2_125_3477_n237), .A2(
        DP_OP_423J2_125_3477_n63), .Y(DP_OP_423J2_125_3477_n61) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U42 ( .A1(DP_OP_423J2_125_3477_n259), .A2(
        DP_OP_423J2_125_3477_n260), .Y(DP_OP_423J2_125_3477_n59) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U41 ( .A1(DP_OP_423J2_125_3477_n260), .A2(
        DP_OP_423J2_125_3477_n259), .Y(DP_OP_423J2_125_3477_n58) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U32 ( .A1(DP_OP_423J2_125_3477_n257), .A2(
        DP_OP_423J2_125_3477_n258), .Y(DP_OP_423J2_125_3477_n52) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U25 ( .A1(DP_OP_423J2_125_3477_n56), .A2(
        n432), .Y(DP_OP_423J2_125_3477_n47) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U22 ( .A1(DP_OP_423J2_125_3477_n255), .A2(
        DP_OP_423J2_125_3477_n256), .Y(DP_OP_423J2_125_3477_n45) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U21 ( .A1(DP_OP_423J2_125_3477_n256), .A2(
        DP_OP_423J2_125_3477_n255), .Y(DP_OP_423J2_125_3477_n44) );
  AOI21X1_HVT DP_OP_423J2_125_3477_U16 ( .A1(DP_OP_423J2_125_3477_n162), .A2(
        DP_OP_423J2_125_3477_n42), .A3(DP_OP_423J2_125_3477_n43), .Y(
        DP_OP_423J2_125_3477_n41) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U14 ( .A1(DP_OP_423J2_125_3477_n253), .A2(
        DP_OP_423J2_125_3477_n254), .Y(DP_OP_423J2_125_3477_n40) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U13 ( .A1(DP_OP_423J2_125_3477_n254), .A2(
        DP_OP_423J2_125_3477_n253), .Y(DP_OP_423J2_125_3477_n39) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U8 ( .A1(n441), .A2(
        DP_OP_423J2_125_3477_n252), .Y(DP_OP_423J2_125_3477_n37) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U96 ( .A1(DP_OP_422J2_124_3477_n101), .A2(
        DP_OP_422J2_124_3477_n105), .A3(DP_OP_422J2_124_3477_n102), .Y(
        DP_OP_422J2_124_3477_n100) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U261 ( .A1(DP_OP_422J2_124_3477_n211), .A2(
        DP_OP_422J2_124_3477_n209), .A3(DP_OP_422J2_124_3477_n210), .Y(
        DP_OP_422J2_124_3477_n208) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U76 ( .A1(DP_OP_422J2_124_3477_n87), .A2(
        DP_OP_422J2_124_3477_n91), .A3(DP_OP_422J2_124_3477_n88), .Y(
        DP_OP_422J2_124_3477_n86) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U116 ( .A1(DP_OP_422J2_124_3477_n115), .A2(
        DP_OP_422J2_124_3477_n119), .A3(DP_OP_422J2_124_3477_n116), .Y(
        DP_OP_422J2_124_3477_n114) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U136 ( .A1(DP_OP_422J2_124_3477_n133), .A2(
        DP_OP_422J2_124_3477_n129), .A3(DP_OP_422J2_124_3477_n130), .Y(
        DP_OP_422J2_124_3477_n128) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U275 ( .A1(DP_OP_422J2_124_3477_n4), .A2(
        DP_OP_422J2_124_3477_n217), .A3(DP_OP_422J2_124_3477_n218), .Y(
        DP_OP_422J2_124_3477_n216) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1111 ( .A1(n496), .A2(
        DP_OP_423J2_125_3477_n2), .Y(DP_OP_422J2_124_3477_n288) );
  XNOR2X1_HVT DP_OP_422J2_124_3477_U737 ( .A1(DP_OP_422J2_124_3477_n2452), 
        .A2(DP_OP_422J2_124_3477_n2979), .Y(DP_OP_422J2_124_3477_n1161) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1109 ( .A1(n337), .A2(n390), .Y(
        DP_OP_422J2_124_3477_n280) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2239 ( .A1(DP_OP_422J2_124_3477_n3006), .A2(
        DP_OP_422J2_124_3477_n3017), .Y(DP_OP_422J2_124_3477_n2998) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2231 ( .A1(DP_OP_422J2_124_3477_n3006), .A2(
        DP_OP_422J2_124_3477_n3016), .Y(DP_OP_422J2_124_3477_n2990) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2223 ( .A1(DP_OP_422J2_124_3477_n3006), .A2(
        DP_OP_422J2_124_3477_n3015), .Y(DP_OP_422J2_124_3477_n2982) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2222 ( .A1(DP_OP_422J2_124_3477_n3013), .A2(
        DP_OP_422J2_124_3477_n3014), .Y(DP_OP_422J2_124_3477_n1678) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2221 ( .A1(DP_OP_422J2_124_3477_n3012), .A2(
        DP_OP_422J2_124_3477_n3014), .Y(DP_OP_422J2_124_3477_n2981) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2220 ( .A1(DP_OP_422J2_124_3477_n3011), .A2(
        DP_OP_422J2_124_3477_n3014), .Y(DP_OP_422J2_124_3477_n2980) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2219 ( .A1(DP_OP_422J2_124_3477_n3010), .A2(
        DP_OP_422J2_124_3477_n3014), .Y(DP_OP_422J2_124_3477_n2979) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2218 ( .A1(DP_OP_422J2_124_3477_n3009), .A2(
        DP_OP_422J2_124_3477_n3014), .Y(DP_OP_422J2_124_3477_n2978) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2217 ( .A1(DP_OP_422J2_124_3477_n3008), .A2(
        DP_OP_422J2_124_3477_n3014), .Y(DP_OP_422J2_124_3477_n770) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2216 ( .A1(DP_OP_422J2_124_3477_n3007), .A2(
        DP_OP_422J2_124_3477_n3014), .Y(DP_OP_422J2_124_3477_n2977) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2215 ( .A1(DP_OP_422J2_124_3477_n3006), 
        .A2(DP_OP_422J2_124_3477_n3014), .Y(DP_OP_422J2_124_3477_n2976) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2195 ( .A1(DP_OP_422J2_124_3477_n2964), .A2(
        DP_OP_422J2_124_3477_n2975), .Y(DP_OP_422J2_124_3477_n2956) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2187 ( .A1(DP_OP_422J2_124_3477_n2964), .A2(
        DP_OP_422J2_124_3477_n2974), .Y(DP_OP_422J2_124_3477_n2948) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2179 ( .A1(DP_OP_422J2_124_3477_n2964), .A2(
        DP_OP_422J2_124_3477_n2973), .Y(DP_OP_422J2_124_3477_n2940) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2178 ( .A1(DP_OP_422J2_124_3477_n2971), .A2(
        DP_OP_422J2_124_3477_n2972), .Y(DP_OP_422J2_124_3477_n2939) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2177 ( .A1(DP_OP_422J2_124_3477_n2970), .A2(
        DP_OP_422J2_124_3477_n2972), .Y(DP_OP_422J2_124_3477_n2938) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2176 ( .A1(DP_OP_422J2_124_3477_n2969), .A2(
        DP_OP_422J2_124_3477_n2972), .Y(DP_OP_422J2_124_3477_n2937) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2175 ( .A1(DP_OP_423J2_125_3477_n2000), .A2(
        DP_OP_422J2_124_3477_n2972), .Y(DP_OP_422J2_124_3477_n2936) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2174 ( .A1(DP_OP_424J2_126_3477_n2087), .A2(
        DP_OP_422J2_124_3477_n2972), .Y(DP_OP_422J2_124_3477_n2935) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2173 ( .A1(DP_OP_423J2_125_3477_n1998), .A2(
        DP_OP_422J2_124_3477_n2972), .Y(DP_OP_422J2_124_3477_n2934) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2172 ( .A1(DP_OP_423J2_125_3477_n1997), .A2(
        DP_OP_422J2_124_3477_n2972), .Y(DP_OP_422J2_124_3477_n2933) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2171 ( .A1(DP_OP_422J2_124_3477_n2964), 
        .A2(DP_OP_422J2_124_3477_n2972), .Y(DP_OP_422J2_124_3477_n2932) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2151 ( .A1(DP_OP_424J2_126_3477_n2128), .A2(
        DP_OP_422J2_124_3477_n2931), .Y(DP_OP_422J2_124_3477_n2912) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2143 ( .A1(DP_OP_424J2_126_3477_n2128), .A2(
        DP_OP_422J2_124_3477_n2930), .Y(DP_OP_422J2_124_3477_n2904) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2135 ( .A1(DP_OP_424J2_126_3477_n2128), .A2(
        DP_OP_422J2_124_3477_n2929), .Y(DP_OP_422J2_124_3477_n2896) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2134 ( .A1(DP_OP_422J2_124_3477_n2927), .A2(
        DP_OP_422J2_124_3477_n2928), .Y(DP_OP_422J2_124_3477_n2895) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2133 ( .A1(DP_OP_422J2_124_3477_n2926), .A2(
        DP_OP_422J2_124_3477_n2928), .Y(DP_OP_422J2_124_3477_n2894) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2132 ( .A1(DP_OP_424J2_126_3477_n2133), .A2(
        DP_OP_422J2_124_3477_n2928), .Y(DP_OP_422J2_124_3477_n2893) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2131 ( .A1(DP_OP_422J2_124_3477_n2924), .A2(
        DP_OP_422J2_124_3477_n2928), .Y(DP_OP_422J2_124_3477_n2892) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2130 ( .A1(DP_OP_422J2_124_3477_n2923), .A2(
        DP_OP_422J2_124_3477_n2928), .Y(DP_OP_422J2_124_3477_n2891) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2129 ( .A1(DP_OP_422J2_124_3477_n2922), .A2(
        DP_OP_422J2_124_3477_n2928), .Y(DP_OP_422J2_124_3477_n2890) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2128 ( .A1(DP_OP_422J2_124_3477_n2921), .A2(
        DP_OP_422J2_124_3477_n2928), .Y(DP_OP_422J2_124_3477_n2889) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2127 ( .A1(DP_OP_424J2_126_3477_n2128), 
        .A2(DP_OP_422J2_124_3477_n2928), .Y(DP_OP_422J2_124_3477_n2888) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2107 ( .A1(DP_OP_423J2_125_3477_n2084), .A2(
        DP_OP_422J2_124_3477_n2887), .Y(DP_OP_422J2_124_3477_n2868) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2099 ( .A1(DP_OP_423J2_125_3477_n2084), .A2(
        DP_OP_422J2_124_3477_n2886), .Y(DP_OP_422J2_124_3477_n2860) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2092 ( .A1(DP_OP_422J2_124_3477_n2877), 
        .A2(DP_OP_422J2_124_3477_n2885), .Y(DP_OP_422J2_124_3477_n2853) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2091 ( .A1(DP_OP_424J2_126_3477_n2172), .A2(
        DP_OP_422J2_124_3477_n2885), .Y(DP_OP_422J2_124_3477_n2852) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2090 ( .A1(DP_OP_422J2_124_3477_n2883), .A2(
        DP_OP_422J2_124_3477_n2884), .Y(DP_OP_422J2_124_3477_n2851) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2089 ( .A1(DP_OP_424J2_126_3477_n2178), .A2(
        DP_OP_422J2_124_3477_n2884), .Y(DP_OP_422J2_124_3477_n2850) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2088 ( .A1(DP_OP_424J2_126_3477_n2177), .A2(
        DP_OP_422J2_124_3477_n2884), .Y(DP_OP_422J2_124_3477_n2849) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2087 ( .A1(DP_OP_422J2_124_3477_n2880), .A2(
        DP_OP_422J2_124_3477_n2884), .Y(DP_OP_422J2_124_3477_n2848) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2086 ( .A1(DP_OP_423J2_125_3477_n2087), .A2(
        DP_OP_422J2_124_3477_n2884), .Y(DP_OP_422J2_124_3477_n2847) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2085 ( .A1(DP_OP_422J2_124_3477_n2878), .A2(
        DP_OP_422J2_124_3477_n2884), .Y(DP_OP_422J2_124_3477_n2846) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2084 ( .A1(DP_OP_422J2_124_3477_n2877), .A2(
        DP_OP_422J2_124_3477_n2884), .Y(DP_OP_422J2_124_3477_n2845) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2083 ( .A1(DP_OP_424J2_126_3477_n2172), 
        .A2(DP_OP_422J2_124_3477_n2884), .Y(DP_OP_422J2_124_3477_n2844) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2063 ( .A1(DP_OP_423J2_125_3477_n2128), .A2(
        DP_OP_422J2_124_3477_n2843), .Y(DP_OP_422J2_124_3477_n2824) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2055 ( .A1(DP_OP_425J2_127_3477_n2700), .A2(
        DP_OP_422J2_124_3477_n2842), .Y(DP_OP_422J2_124_3477_n2816) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2048 ( .A1(DP_OP_422J2_124_3477_n2833), 
        .A2(DP_OP_422J2_124_3477_n2841), .Y(DP_OP_422J2_124_3477_n2809) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2047 ( .A1(DP_OP_423J2_125_3477_n2128), .A2(
        DP_OP_423J2_125_3477_n2841), .Y(DP_OP_422J2_124_3477_n2808) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2046 ( .A1(DP_OP_425J2_127_3477_n2707), .A2(
        DP_OP_422J2_124_3477_n2840), .Y(DP_OP_422J2_124_3477_n2807) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2045 ( .A1(DP_OP_422J2_124_3477_n2838), .A2(
        DP_OP_422J2_124_3477_n2840), .Y(DP_OP_422J2_124_3477_n2806) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2044 ( .A1(DP_OP_422J2_124_3477_n2837), .A2(
        DP_OP_422J2_124_3477_n2840), .Y(DP_OP_422J2_124_3477_n2805) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2043 ( .A1(DP_OP_424J2_126_3477_n2220), .A2(
        DP_OP_422J2_124_3477_n2840), .Y(DP_OP_422J2_124_3477_n2804) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2042 ( .A1(DP_OP_422J2_124_3477_n2835), .A2(
        DP_OP_422J2_124_3477_n2840), .Y(DP_OP_422J2_124_3477_n2803) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2041 ( .A1(DP_OP_422J2_124_3477_n2834), .A2(
        DP_OP_422J2_124_3477_n2840), .Y(DP_OP_422J2_124_3477_n2802) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2040 ( .A1(DP_OP_422J2_124_3477_n2833), .A2(
        DP_OP_422J2_124_3477_n2840), .Y(DP_OP_422J2_124_3477_n2801) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2039 ( .A1(DP_OP_423J2_125_3477_n2128), 
        .A2(DP_OP_422J2_124_3477_n2840), .Y(DP_OP_422J2_124_3477_n2800) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2020 ( .A1(DP_OP_422J2_124_3477_n2789), 
        .A2(DP_OP_422J2_124_3477_n2799), .Y(DP_OP_422J2_124_3477_n2781) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2019 ( .A1(DP_OP_424J2_126_3477_n2260), .A2(
        DP_OP_422J2_124_3477_n2799), .Y(DP_OP_422J2_124_3477_n2780) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2011 ( .A1(DP_OP_423J2_125_3477_n2172), .A2(
        DP_OP_422J2_124_3477_n2798), .Y(DP_OP_422J2_124_3477_n2772) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2004 ( .A1(DP_OP_422J2_124_3477_n2789), 
        .A2(DP_OP_422J2_124_3477_n2797), .Y(DP_OP_422J2_124_3477_n2765) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2003 ( .A1(DP_OP_424J2_126_3477_n2260), .A2(
        DP_OP_422J2_124_3477_n2797), .Y(DP_OP_422J2_124_3477_n2764) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2002 ( .A1(DP_OP_422J2_124_3477_n2795), .A2(
        DP_OP_422J2_124_3477_n2796), .Y(DP_OP_422J2_124_3477_n2763) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2001 ( .A1(DP_OP_425J2_127_3477_n2662), .A2(
        DP_OP_422J2_124_3477_n2796), .Y(DP_OP_422J2_124_3477_n2762) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2000 ( .A1(DP_OP_422J2_124_3477_n2793), .A2(
        DP_OP_422J2_124_3477_n2796), .Y(DP_OP_422J2_124_3477_n2761) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1999 ( .A1(DP_OP_422J2_124_3477_n2792), .A2(
        DP_OP_422J2_124_3477_n2796), .Y(DP_OP_422J2_124_3477_n2760) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1998 ( .A1(DP_OP_422J2_124_3477_n2791), .A2(
        DP_OP_422J2_124_3477_n2796), .Y(DP_OP_422J2_124_3477_n2759) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1997 ( .A1(DP_OP_422J2_124_3477_n2790), .A2(
        DP_OP_422J2_124_3477_n2796), .Y(DP_OP_422J2_124_3477_n2758) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1996 ( .A1(DP_OP_422J2_124_3477_n2789), .A2(
        DP_OP_422J2_124_3477_n2796), .Y(DP_OP_422J2_124_3477_n2757) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1995 ( .A1(DP_OP_424J2_126_3477_n2260), 
        .A2(DP_OP_422J2_124_3477_n2796), .Y(DP_OP_422J2_124_3477_n2756) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1982 ( .A1(DP_OP_422J2_124_3477_n2751), 
        .A2(DP_OP_422J2_124_3477_n2755), .Y(DP_OP_422J2_124_3477_n2743) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1981 ( .A1(DP_OP_422J2_124_3477_n2750), 
        .A2(DP_OP_422J2_124_3477_n2755), .Y(DP_OP_422J2_124_3477_n2742) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1980 ( .A1(DP_OP_422J2_124_3477_n2749), 
        .A2(DP_OP_422J2_124_3477_n2755), .Y(DP_OP_422J2_124_3477_n2741) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1979 ( .A1(DP_OP_425J2_127_3477_n2616), 
        .A2(DP_OP_422J2_124_3477_n2755), .Y(DP_OP_422J2_124_3477_n2740) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1978 ( .A1(DP_OP_422J2_124_3477_n2747), 
        .A2(DP_OP_422J2_124_3477_n2755), .Y(DP_OP_422J2_124_3477_n2739) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1977 ( .A1(DP_OP_422J2_124_3477_n2746), 
        .A2(DP_OP_422J2_124_3477_n2755), .Y(DP_OP_422J2_124_3477_n2738) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1976 ( .A1(DP_OP_422J2_124_3477_n2745), 
        .A2(DP_OP_422J2_124_3477_n2755), .Y(DP_OP_422J2_124_3477_n2737) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1975 ( .A1(DP_OP_425J2_127_3477_n2612), .A2(
        DP_OP_422J2_124_3477_n2755), .Y(DP_OP_422J2_124_3477_n2736) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1968 ( .A1(DP_OP_422J2_124_3477_n2745), 
        .A2(DP_OP_422J2_124_3477_n2754), .Y(DP_OP_422J2_124_3477_n2729) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1967 ( .A1(DP_OP_425J2_127_3477_n2612), .A2(
        DP_OP_422J2_124_3477_n2754), .Y(DP_OP_422J2_124_3477_n2728) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1959 ( .A1(DP_OP_425J2_127_3477_n2612), .A2(
        DP_OP_422J2_124_3477_n2753), .Y(DP_OP_422J2_124_3477_n2720) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1958 ( .A1(DP_OP_422J2_124_3477_n2751), .A2(
        DP_OP_422J2_124_3477_n2752), .Y(DP_OP_422J2_124_3477_n2719) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1957 ( .A1(DP_OP_422J2_124_3477_n2750), .A2(
        DP_OP_422J2_124_3477_n2752), .Y(DP_OP_422J2_124_3477_n2718) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1956 ( .A1(DP_OP_422J2_124_3477_n2749), .A2(
        DP_OP_422J2_124_3477_n2752), .Y(DP_OP_422J2_124_3477_n2717) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1955 ( .A1(DP_OP_424J2_126_3477_n2308), .A2(
        DP_OP_422J2_124_3477_n2752), .Y(DP_OP_422J2_124_3477_n2716) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1954 ( .A1(DP_OP_422J2_124_3477_n2747), .A2(
        DP_OP_422J2_124_3477_n2752), .Y(DP_OP_422J2_124_3477_n2715) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1953 ( .A1(DP_OP_422J2_124_3477_n2746), .A2(
        DP_OP_422J2_124_3477_n2752), .Y(DP_OP_422J2_124_3477_n2714) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1952 ( .A1(DP_OP_422J2_124_3477_n2745), .A2(
        DP_OP_422J2_124_3477_n2752), .Y(DP_OP_422J2_124_3477_n2713) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1951 ( .A1(DP_OP_424J2_126_3477_n2304), 
        .A2(DP_OP_422J2_124_3477_n2752), .Y(DP_OP_422J2_124_3477_n2712) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1931 ( .A1(DP_OP_422J2_124_3477_n2700), .A2(
        DP_OP_422J2_124_3477_n2711), .Y(DP_OP_422J2_124_3477_n2692) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1923 ( .A1(DP_OP_422J2_124_3477_n2700), .A2(
        DP_OP_422J2_124_3477_n2710), .Y(DP_OP_422J2_124_3477_n2684) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1916 ( .A1(DP_OP_422J2_124_3477_n2701), 
        .A2(DP_OP_422J2_124_3477_n2709), .Y(DP_OP_422J2_124_3477_n2677) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1915 ( .A1(DP_OP_422J2_124_3477_n2700), .A2(
        DP_OP_422J2_124_3477_n2709), .Y(DP_OP_422J2_124_3477_n2676) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1914 ( .A1(DP_OP_422J2_124_3477_n2707), .A2(
        DP_OP_422J2_124_3477_n2708), .Y(DP_OP_422J2_124_3477_n2675) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1913 ( .A1(DP_OP_424J2_126_3477_n2354), .A2(
        DP_OP_422J2_124_3477_n2708), .Y(DP_OP_422J2_124_3477_n2674) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1912 ( .A1(DP_OP_424J2_126_3477_n2353), .A2(
        DP_OP_422J2_124_3477_n2708), .Y(DP_OP_422J2_124_3477_n2673) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1911 ( .A1(DP_OP_422J2_124_3477_n2704), .A2(
        DP_OP_422J2_124_3477_n2708), .Y(DP_OP_422J2_124_3477_n2672) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1910 ( .A1(DP_OP_424J2_126_3477_n2351), .A2(
        DP_OP_422J2_124_3477_n2708), .Y(DP_OP_422J2_124_3477_n2671) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1909 ( .A1(DP_OP_422J2_124_3477_n2702), .A2(
        DP_OP_422J2_124_3477_n2708), .Y(DP_OP_422J2_124_3477_n2670) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1908 ( .A1(DP_OP_422J2_124_3477_n2701), .A2(
        DP_OP_422J2_124_3477_n2708), .Y(DP_OP_422J2_124_3477_n2669) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1907 ( .A1(DP_OP_422J2_124_3477_n2700), 
        .A2(DP_OP_422J2_124_3477_n2708), .Y(DP_OP_422J2_124_3477_n2668) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1888 ( .A1(DP_OP_425J2_127_3477_n2525), 
        .A2(DP_OP_422J2_124_3477_n2667), .Y(DP_OP_422J2_124_3477_n2649) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1887 ( .A1(DP_OP_422J2_124_3477_n2656), .A2(
        DP_OP_422J2_124_3477_n2667), .Y(DP_OP_422J2_124_3477_n2648) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1879 ( .A1(DP_OP_422J2_124_3477_n2656), .A2(
        DP_OP_422J2_124_3477_n2666), .Y(DP_OP_422J2_124_3477_n2640) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1871 ( .A1(DP_OP_422J2_124_3477_n2656), .A2(
        DP_OP_423J2_125_3477_n2665), .Y(DP_OP_422J2_124_3477_n2632) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1870 ( .A1(DP_OP_422J2_124_3477_n2663), .A2(
        DP_OP_422J2_124_3477_n2664), .Y(DP_OP_422J2_124_3477_n2631) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1869 ( .A1(DP_OP_422J2_124_3477_n2662), .A2(
        DP_OP_422J2_124_3477_n2664), .Y(DP_OP_422J2_124_3477_n2630) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1868 ( .A1(DP_OP_424J2_126_3477_n2397), .A2(
        DP_OP_422J2_124_3477_n2664), .Y(DP_OP_422J2_124_3477_n2629) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1867 ( .A1(DP_OP_425J2_127_3477_n2528), .A2(
        DP_OP_422J2_124_3477_n2664), .Y(DP_OP_422J2_124_3477_n2628) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1866 ( .A1(DP_OP_422J2_124_3477_n2659), .A2(
        DP_OP_422J2_124_3477_n2664), .Y(DP_OP_422J2_124_3477_n2627) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1865 ( .A1(DP_OP_422J2_124_3477_n2658), .A2(
        DP_OP_422J2_124_3477_n2664), .Y(DP_OP_422J2_124_3477_n2626) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1864 ( .A1(DP_OP_425J2_127_3477_n2525), .A2(
        DP_OP_422J2_124_3477_n2664), .Y(DP_OP_422J2_124_3477_n2625) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1863 ( .A1(DP_OP_422J2_124_3477_n2656), 
        .A2(DP_OP_422J2_124_3477_n2664), .Y(DP_OP_422J2_124_3477_n2624) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1843 ( .A1(DP_OP_422J2_124_3477_n2612), .A2(
        DP_OP_422J2_124_3477_n2623), .Y(DP_OP_422J2_124_3477_n2604) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1842 ( .A1(DP_OP_422J2_124_3477_n2619), 
        .A2(DP_OP_422J2_124_3477_n2622), .Y(DP_OP_422J2_124_3477_n2603) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1841 ( .A1(DP_OP_424J2_126_3477_n2442), 
        .A2(DP_OP_422J2_124_3477_n2622), .Y(DP_OP_422J2_124_3477_n2602) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1840 ( .A1(DP_OP_422J2_124_3477_n2617), 
        .A2(DP_OP_422J2_124_3477_n2622), .Y(DP_OP_422J2_124_3477_n2601) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1839 ( .A1(DP_OP_422J2_124_3477_n2616), 
        .A2(DP_OP_422J2_124_3477_n2622), .Y(DP_OP_422J2_124_3477_n2600) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1838 ( .A1(DP_OP_423J2_125_3477_n2351), 
        .A2(DP_OP_422J2_124_3477_n2622), .Y(DP_OP_422J2_124_3477_n2599) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1837 ( .A1(DP_OP_423J2_125_3477_n2350), 
        .A2(DP_OP_422J2_124_3477_n2622), .Y(DP_OP_422J2_124_3477_n2598) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1836 ( .A1(DP_OP_422J2_124_3477_n2613), 
        .A2(DP_OP_422J2_124_3477_n2622), .Y(DP_OP_422J2_124_3477_n2597) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1835 ( .A1(DP_OP_422J2_124_3477_n2612), .A2(
        DP_OP_422J2_124_3477_n2622), .Y(DP_OP_422J2_124_3477_n2596) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1827 ( .A1(DP_OP_422J2_124_3477_n2612), .A2(
        DP_OP_422J2_124_3477_n2621), .Y(DP_OP_422J2_124_3477_n2588) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1826 ( .A1(DP_OP_422J2_124_3477_n2619), .A2(
        DP_OP_422J2_124_3477_n2620), .Y(DP_OP_422J2_124_3477_n2587) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1825 ( .A1(DP_OP_423J2_125_3477_n2354), .A2(
        DP_OP_422J2_124_3477_n2620), .Y(DP_OP_422J2_124_3477_n2586) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1824 ( .A1(DP_OP_422J2_124_3477_n2617), .A2(
        DP_OP_422J2_124_3477_n2620), .Y(DP_OP_422J2_124_3477_n2585) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1823 ( .A1(DP_OP_422J2_124_3477_n2616), .A2(
        DP_OP_422J2_124_3477_n2620), .Y(DP_OP_422J2_124_3477_n2584) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1822 ( .A1(DP_OP_424J2_126_3477_n2439), .A2(
        DP_OP_422J2_124_3477_n2620), .Y(DP_OP_422J2_124_3477_n2583) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1821 ( .A1(DP_OP_425J2_127_3477_n2482), .A2(
        DP_OP_422J2_124_3477_n2620), .Y(DP_OP_422J2_124_3477_n2582) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1820 ( .A1(DP_OP_422J2_124_3477_n2613), .A2(
        DP_OP_422J2_124_3477_n2620), .Y(DP_OP_422J2_124_3477_n2581) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1819 ( .A1(DP_OP_422J2_124_3477_n2612), 
        .A2(DP_OP_422J2_124_3477_n2620), .Y(DP_OP_422J2_124_3477_n2580) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1800 ( .A1(DP_OP_422J2_124_3477_n2569), 
        .A2(DP_OP_422J2_124_3477_n2579), .Y(DP_OP_422J2_124_3477_n2561) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1799 ( .A1(DP_OP_422J2_124_3477_n2568), .A2(
        DP_OP_422J2_124_3477_n2579), .Y(DP_OP_422J2_124_3477_n2560) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1791 ( .A1(DP_OP_422J2_124_3477_n2568), .A2(
        DP_OP_422J2_124_3477_n2578), .Y(DP_OP_422J2_124_3477_n2552) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1784 ( .A1(DP_OP_422J2_124_3477_n2569), 
        .A2(DP_OP_422J2_124_3477_n2577), .Y(DP_OP_422J2_124_3477_n2545) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1783 ( .A1(DP_OP_422J2_124_3477_n2568), .A2(
        DP_OP_422J2_124_3477_n2577), .Y(DP_OP_422J2_124_3477_n2544) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1782 ( .A1(DP_OP_422J2_124_3477_n2575), .A2(
        DP_OP_422J2_124_3477_n2576), .Y(DP_OP_422J2_124_3477_n2543) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1781 ( .A1(DP_OP_423J2_125_3477_n2398), .A2(
        DP_OP_422J2_124_3477_n2576), .Y(DP_OP_422J2_124_3477_n2542) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1780 ( .A1(DP_OP_423J2_125_3477_n2397), .A2(
        DP_OP_422J2_124_3477_n2576), .Y(DP_OP_422J2_124_3477_n2541) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1779 ( .A1(DP_OP_423J2_125_3477_n2396), .A2(
        DP_OP_422J2_124_3477_n2576), .Y(DP_OP_422J2_124_3477_n2540) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1778 ( .A1(DP_OP_422J2_124_3477_n2571), .A2(
        DP_OP_422J2_124_3477_n2576), .Y(DP_OP_422J2_124_3477_n2539) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1777 ( .A1(DP_OP_422J2_124_3477_n2570), .A2(
        DP_OP_422J2_124_3477_n2576), .Y(DP_OP_422J2_124_3477_n2538) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1776 ( .A1(DP_OP_422J2_124_3477_n2569), .A2(
        DP_OP_422J2_124_3477_n2576), .Y(DP_OP_422J2_124_3477_n2537) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1775 ( .A1(DP_OP_422J2_124_3477_n2568), 
        .A2(DP_OP_422J2_124_3477_n2576), .Y(DP_OP_422J2_124_3477_n2536) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1755 ( .A1(DP_OP_423J2_125_3477_n2436), .A2(
        DP_OP_422J2_124_3477_n2535), .Y(DP_OP_422J2_124_3477_n2516) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1747 ( .A1(DP_OP_423J2_125_3477_n2436), .A2(
        DP_OP_422J2_124_3477_n2534), .Y(DP_OP_422J2_124_3477_n2508) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1740 ( .A1(DP_OP_423J2_125_3477_n2437), 
        .A2(DP_OP_422J2_124_3477_n2533), .Y(DP_OP_422J2_124_3477_n2501) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1739 ( .A1(DP_OP_423J2_125_3477_n2436), .A2(
        DP_OP_422J2_124_3477_n2533), .Y(DP_OP_422J2_124_3477_n2500) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1738 ( .A1(DP_OP_422J2_124_3477_n2531), .A2(
        DP_OP_422J2_124_3477_n2532), .Y(DP_OP_422J2_124_3477_n2499) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1737 ( .A1(DP_OP_423J2_125_3477_n2442), .A2(
        DP_OP_422J2_124_3477_n2532), .Y(DP_OP_422J2_124_3477_n2498) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1736 ( .A1(DP_OP_423J2_125_3477_n2441), .A2(
        DP_OP_422J2_124_3477_n2532), .Y(DP_OP_422J2_124_3477_n2497) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1735 ( .A1(DP_OP_422J2_124_3477_n2528), .A2(
        DP_OP_422J2_124_3477_n2532), .Y(DP_OP_422J2_124_3477_n2496) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1734 ( .A1(DP_OP_423J2_125_3477_n2439), .A2(
        DP_OP_422J2_124_3477_n2532), .Y(DP_OP_422J2_124_3477_n2495) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1733 ( .A1(DP_OP_422J2_124_3477_n2526), .A2(
        DP_OP_422J2_124_3477_n2532), .Y(DP_OP_422J2_124_3477_n2494) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1732 ( .A1(DP_OP_423J2_125_3477_n2437), .A2(
        DP_OP_422J2_124_3477_n2532), .Y(DP_OP_422J2_124_3477_n2493) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1731 ( .A1(DP_OP_423J2_125_3477_n2436), 
        .A2(DP_OP_422J2_124_3477_n2532), .Y(DP_OP_422J2_124_3477_n2492) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1711 ( .A1(DP_OP_422J2_124_3477_n2480), .A2(
        DP_OP_422J2_124_3477_n2491), .Y(DP_OP_422J2_124_3477_n2472) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1703 ( .A1(DP_OP_422J2_124_3477_n2480), .A2(
        DP_OP_422J2_124_3477_n2490), .Y(DP_OP_422J2_124_3477_n2464) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1695 ( .A1(DP_OP_422J2_124_3477_n2480), .A2(
        DP_OP_422J2_124_3477_n2489), .Y(DP_OP_422J2_124_3477_n2456) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1694 ( .A1(DP_OP_422J2_124_3477_n2487), .A2(
        DP_OP_422J2_124_3477_n2488), .Y(DP_OP_422J2_124_3477_n2455) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1693 ( .A1(DP_OP_422J2_124_3477_n2486), .A2(
        DP_OP_422J2_124_3477_n2488), .Y(DP_OP_422J2_124_3477_n2454) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1692 ( .A1(DP_OP_422J2_124_3477_n2485), .A2(
        DP_OP_422J2_124_3477_n2488), .Y(DP_OP_422J2_124_3477_n2453) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1691 ( .A1(DP_OP_422J2_124_3477_n2484), .A2(
        DP_OP_422J2_124_3477_n2488), .Y(DP_OP_422J2_124_3477_n2452) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1690 ( .A1(DP_OP_422J2_124_3477_n2483), .A2(
        DP_OP_422J2_124_3477_n2488), .Y(DP_OP_422J2_124_3477_n2451) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1689 ( .A1(DP_OP_422J2_124_3477_n2482), .A2(
        DP_OP_422J2_124_3477_n2488), .Y(DP_OP_422J2_124_3477_n2450) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1688 ( .A1(DP_OP_422J2_124_3477_n2481), .A2(
        DP_OP_422J2_124_3477_n2488), .Y(DP_OP_422J2_124_3477_n2449) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1687 ( .A1(DP_OP_422J2_124_3477_n2480), 
        .A2(DP_OP_422J2_124_3477_n2488), .Y(DP_OP_422J2_124_3477_n2448) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1667 ( .A1(DP_OP_422J2_124_3477_n2436), .A2(
        DP_OP_422J2_124_3477_n2447), .Y(DP_OP_422J2_124_3477_n2428) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1659 ( .A1(DP_OP_422J2_124_3477_n2436), .A2(
        DP_OP_422J2_124_3477_n2446), .Y(DP_OP_422J2_124_3477_n2420) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1650 ( .A1(DP_OP_423J2_125_3477_n2487), .A2(
        DP_OP_422J2_124_3477_n2444), .Y(DP_OP_422J2_124_3477_n2411) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1649 ( .A1(DP_OP_422J2_124_3477_n2442), .A2(
        DP_OP_422J2_124_3477_n2444), .Y(DP_OP_422J2_124_3477_n2410) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1648 ( .A1(DP_OP_422J2_124_3477_n2441), .A2(
        DP_OP_422J2_124_3477_n2444), .Y(DP_OP_422J2_124_3477_n2409) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1647 ( .A1(DP_OP_423J2_125_3477_n2484), .A2(
        DP_OP_422J2_124_3477_n2444), .Y(DP_OP_422J2_124_3477_n2408) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1646 ( .A1(DP_OP_422J2_124_3477_n2439), .A2(
        DP_OP_422J2_124_3477_n2444), .Y(DP_OP_422J2_124_3477_n2407) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1645 ( .A1(DP_OP_423J2_125_3477_n2482), .A2(
        DP_OP_422J2_124_3477_n2444), .Y(DP_OP_422J2_124_3477_n2406) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1644 ( .A1(DP_OP_423J2_125_3477_n2481), .A2(
        DP_OP_422J2_124_3477_n2444), .Y(DP_OP_422J2_124_3477_n2405) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1643 ( .A1(DP_OP_422J2_124_3477_n2436), 
        .A2(DP_OP_422J2_124_3477_n2444), .Y(DP_OP_422J2_124_3477_n2404) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1623 ( .A1(DP_OP_422J2_124_3477_n2392), .A2(
        DP_OP_422J2_124_3477_n2403), .Y(DP_OP_422J2_124_3477_n2384) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1615 ( .A1(DP_OP_422J2_124_3477_n2392), .A2(
        DP_OP_423J2_125_3477_n2402), .Y(DP_OP_422J2_124_3477_n2376) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1607 ( .A1(DP_OP_422J2_124_3477_n2392), .A2(
        DP_OP_422J2_124_3477_n2401), .Y(DP_OP_422J2_124_3477_n2368) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1606 ( .A1(DP_OP_423J2_125_3477_n2531), .A2(
        DP_OP_422J2_124_3477_n2400), .Y(DP_OP_422J2_124_3477_n2367) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1605 ( .A1(DP_OP_423J2_125_3477_n2530), .A2(
        DP_OP_422J2_124_3477_n2400), .Y(DP_OP_422J2_124_3477_n2366) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1604 ( .A1(DP_OP_423J2_125_3477_n2529), .A2(
        DP_OP_422J2_124_3477_n2400), .Y(DP_OP_422J2_124_3477_n2365) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1603 ( .A1(DP_OP_423J2_125_3477_n2528), .A2(
        DP_OP_422J2_124_3477_n2400), .Y(DP_OP_422J2_124_3477_n2364) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1602 ( .A1(DP_OP_423J2_125_3477_n2527), .A2(
        DP_OP_422J2_124_3477_n2400), .Y(DP_OP_422J2_124_3477_n2363) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1601 ( .A1(DP_OP_423J2_125_3477_n2526), .A2(
        DP_OP_422J2_124_3477_n2400), .Y(DP_OP_422J2_124_3477_n2362) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1600 ( .A1(DP_OP_423J2_125_3477_n2525), .A2(
        DP_OP_422J2_124_3477_n2400), .Y(DP_OP_422J2_124_3477_n2361) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1599 ( .A1(DP_OP_422J2_124_3477_n2392), 
        .A2(DP_OP_422J2_124_3477_n2400), .Y(DP_OP_422J2_124_3477_n2360) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1579 ( .A1(DP_OP_422J2_124_3477_n2348), .A2(
        DP_OP_422J2_124_3477_n2359), .Y(DP_OP_422J2_124_3477_n2340) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1571 ( .A1(DP_OP_422J2_124_3477_n2348), .A2(
        DP_OP_422J2_124_3477_n2358), .Y(DP_OP_422J2_124_3477_n2332) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1563 ( .A1(DP_OP_422J2_124_3477_n2348), .A2(
        DP_OP_422J2_124_3477_n2357), .Y(DP_OP_422J2_124_3477_n2324) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1562 ( .A1(DP_OP_422J2_124_3477_n2355), .A2(
        DP_OP_422J2_124_3477_n2356), .Y(DP_OP_422J2_124_3477_n2323) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1561 ( .A1(DP_OP_422J2_124_3477_n2354), .A2(
        DP_OP_422J2_124_3477_n2356), .Y(DP_OP_422J2_124_3477_n2322) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1560 ( .A1(DP_OP_422J2_124_3477_n2353), .A2(
        DP_OP_422J2_124_3477_n2356), .Y(DP_OP_422J2_124_3477_n2321) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1559 ( .A1(DP_OP_424J2_126_3477_n2484), .A2(
        DP_OP_422J2_124_3477_n2356), .Y(DP_OP_422J2_124_3477_n2320) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1558 ( .A1(DP_OP_422J2_124_3477_n2351), .A2(
        DP_OP_422J2_124_3477_n2356), .Y(DP_OP_422J2_124_3477_n2319) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1557 ( .A1(DP_OP_424J2_126_3477_n2482), .A2(
        DP_OP_422J2_124_3477_n2356), .Y(DP_OP_422J2_124_3477_n2318) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1556 ( .A1(DP_OP_424J2_126_3477_n2481), .A2(
        DP_OP_422J2_124_3477_n2356), .Y(DP_OP_422J2_124_3477_n2317) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1555 ( .A1(DP_OP_422J2_124_3477_n2348), 
        .A2(DP_OP_422J2_124_3477_n2356), .Y(DP_OP_422J2_124_3477_n2316) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1536 ( .A1(DP_OP_422J2_124_3477_n2305), 
        .A2(DP_OP_422J2_124_3477_n2315), .Y(DP_OP_422J2_124_3477_n2297) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1535 ( .A1(DP_OP_422J2_124_3477_n2304), .A2(
        DP_OP_422J2_124_3477_n2315), .Y(DP_OP_422J2_124_3477_n2296) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1527 ( .A1(DP_OP_422J2_124_3477_n2304), .A2(
        DP_OP_424J2_126_3477_n2314), .Y(DP_OP_422J2_124_3477_n2288) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1519 ( .A1(DP_OP_422J2_124_3477_n2304), .A2(
        DP_OP_422J2_124_3477_n2313), .Y(DP_OP_422J2_124_3477_n2280) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1518 ( .A1(DP_OP_422J2_124_3477_n2311), .A2(
        DP_OP_422J2_124_3477_n2312), .Y(DP_OP_422J2_124_3477_n2279) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1517 ( .A1(DP_OP_424J2_126_3477_n2530), .A2(
        DP_OP_422J2_124_3477_n2312), .Y(DP_OP_422J2_124_3477_n2278) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1516 ( .A1(DP_OP_423J2_125_3477_n2617), .A2(
        DP_OP_422J2_124_3477_n2312), .Y(DP_OP_422J2_124_3477_n2277) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1515 ( .A1(DP_OP_422J2_124_3477_n2308), .A2(
        DP_OP_422J2_124_3477_n2312), .Y(DP_OP_422J2_124_3477_n2276) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1514 ( .A1(DP_OP_422J2_124_3477_n2307), .A2(
        DP_OP_422J2_124_3477_n2312), .Y(DP_OP_422J2_124_3477_n2275) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1513 ( .A1(DP_OP_424J2_126_3477_n2526), .A2(
        DP_OP_422J2_124_3477_n2312), .Y(DP_OP_422J2_124_3477_n2274) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1512 ( .A1(DP_OP_422J2_124_3477_n2305), .A2(
        DP_OP_422J2_124_3477_n2312), .Y(DP_OP_422J2_124_3477_n2273) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1511 ( .A1(DP_OP_422J2_124_3477_n2304), 
        .A2(DP_OP_422J2_124_3477_n2312), .Y(DP_OP_422J2_124_3477_n2272) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1492 ( .A1(DP_OP_422J2_124_3477_n2261), 
        .A2(DP_OP_422J2_124_3477_n2271), .Y(DP_OP_422J2_124_3477_n2253) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1491 ( .A1(DP_OP_422J2_124_3477_n2260), .A2(
        DP_OP_422J2_124_3477_n2271), .Y(DP_OP_422J2_124_3477_n2252) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1483 ( .A1(DP_OP_422J2_124_3477_n2260), .A2(
        DP_OP_422J2_124_3477_n2270), .Y(DP_OP_422J2_124_3477_n2244) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1475 ( .A1(DP_OP_422J2_124_3477_n2260), .A2(
        DP_OP_422J2_124_3477_n2269), .Y(DP_OP_422J2_124_3477_n2236) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1474 ( .A1(DP_OP_422J2_124_3477_n2267), .A2(
        DP_OP_422J2_124_3477_n2268), .Y(DP_OP_422J2_124_3477_n2235) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1473 ( .A1(DP_OP_425J2_127_3477_n2398), .A2(
        DP_OP_422J2_124_3477_n2268), .Y(DP_OP_422J2_124_3477_n2234) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1472 ( .A1(DP_OP_422J2_124_3477_n2265), .A2(
        DP_OP_422J2_124_3477_n2268), .Y(DP_OP_422J2_124_3477_n2233) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1471 ( .A1(DP_OP_425J2_127_3477_n2396), .A2(
        DP_OP_422J2_124_3477_n2268), .Y(DP_OP_422J2_124_3477_n2232) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1470 ( .A1(DP_OP_422J2_124_3477_n2263), .A2(
        DP_OP_422J2_124_3477_n2268), .Y(DP_OP_422J2_124_3477_n2231) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1469 ( .A1(DP_OP_422J2_124_3477_n2262), .A2(
        DP_OP_422J2_124_3477_n2268), .Y(DP_OP_422J2_124_3477_n2230) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1468 ( .A1(DP_OP_422J2_124_3477_n2261), .A2(
        DP_OP_422J2_124_3477_n2268), .Y(DP_OP_422J2_124_3477_n2229) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1467 ( .A1(DP_OP_422J2_124_3477_n2260), 
        .A2(DP_OP_422J2_124_3477_n2268), .Y(DP_OP_422J2_124_3477_n2228) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1448 ( .A1(DP_OP_422J2_124_3477_n2217), 
        .A2(DP_OP_422J2_124_3477_n2227), .Y(DP_OP_422J2_124_3477_n2209) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1447 ( .A1(DP_OP_424J2_126_3477_n2612), .A2(
        DP_OP_422J2_124_3477_n2227), .Y(DP_OP_422J2_124_3477_n2208) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1439 ( .A1(DP_OP_423J2_125_3477_n2700), .A2(
        DP_OP_424J2_126_3477_n2226), .Y(DP_OP_422J2_124_3477_n2200) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1432 ( .A1(DP_OP_422J2_124_3477_n2217), 
        .A2(DP_OP_422J2_124_3477_n2225), .Y(DP_OP_422J2_124_3477_n2193) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1431 ( .A1(DP_OP_424J2_126_3477_n2612), .A2(
        DP_OP_422J2_124_3477_n2225), .Y(DP_OP_422J2_124_3477_n2192) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1430 ( .A1(DP_OP_425J2_127_3477_n2355), .A2(
        DP_OP_422J2_124_3477_n2224), .Y(DP_OP_422J2_124_3477_n2191) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1429 ( .A1(DP_OP_424J2_126_3477_n2618), .A2(
        DP_OP_422J2_124_3477_n2224), .Y(DP_OP_422J2_124_3477_n2190) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1428 ( .A1(DP_OP_425J2_127_3477_n2353), .A2(
        DP_OP_422J2_124_3477_n2224), .Y(DP_OP_422J2_124_3477_n2189) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1427 ( .A1(DP_OP_422J2_124_3477_n2220), .A2(
        DP_OP_422J2_124_3477_n2224), .Y(DP_OP_422J2_124_3477_n2188) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1426 ( .A1(DP_OP_422J2_124_3477_n2219), .A2(
        DP_OP_422J2_124_3477_n2224), .Y(DP_OP_422J2_124_3477_n2187) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1425 ( .A1(DP_OP_422J2_124_3477_n2218), .A2(
        DP_OP_422J2_124_3477_n2224), .Y(DP_OP_422J2_124_3477_n2186) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1424 ( .A1(DP_OP_422J2_124_3477_n2217), .A2(
        DP_OP_422J2_124_3477_n2224), .Y(DP_OP_422J2_124_3477_n2185) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1423 ( .A1(DP_OP_424J2_126_3477_n2612), 
        .A2(DP_OP_422J2_124_3477_n2224), .Y(DP_OP_422J2_124_3477_n2184) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1403 ( .A1(DP_OP_422J2_124_3477_n2172), .A2(
        DP_OP_422J2_124_3477_n2183), .Y(DP_OP_422J2_124_3477_n2164) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1395 ( .A1(DP_OP_422J2_124_3477_n2172), .A2(
        DP_OP_422J2_124_3477_n2182), .Y(DP_OP_422J2_124_3477_n2156) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1387 ( .A1(DP_OP_422J2_124_3477_n2172), .A2(
        DP_OP_422J2_124_3477_n2181), .Y(DP_OP_422J2_124_3477_n2148) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1386 ( .A1(DP_OP_422J2_124_3477_n2179), .A2(
        DP_OP_422J2_124_3477_n2180), .Y(DP_OP_422J2_124_3477_n2147) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1385 ( .A1(DP_OP_422J2_124_3477_n2178), .A2(
        DP_OP_422J2_124_3477_n2180), .Y(DP_OP_422J2_124_3477_n2146) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1384 ( .A1(DP_OP_422J2_124_3477_n2177), .A2(
        DP_OP_422J2_124_3477_n2180), .Y(DP_OP_422J2_124_3477_n2145) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1383 ( .A1(DP_OP_423J2_125_3477_n2748), .A2(
        DP_OP_422J2_124_3477_n2180), .Y(DP_OP_422J2_124_3477_n2144) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1382 ( .A1(DP_OP_425J2_127_3477_n2307), .A2(
        DP_OP_422J2_124_3477_n2180), .Y(DP_OP_422J2_124_3477_n2143) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1381 ( .A1(DP_OP_423J2_125_3477_n2746), .A2(
        DP_OP_422J2_124_3477_n2180), .Y(DP_OP_422J2_124_3477_n2142) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1380 ( .A1(DP_OP_423J2_125_3477_n2745), .A2(
        DP_OP_422J2_124_3477_n2180), .Y(DP_OP_422J2_124_3477_n2141) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1379 ( .A1(DP_OP_422J2_124_3477_n2172), 
        .A2(DP_OP_422J2_124_3477_n2180), .Y(DP_OP_422J2_124_3477_n2140) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1359 ( .A1(DP_OP_424J2_126_3477_n2700), .A2(
        DP_OP_422J2_124_3477_n2139), .Y(DP_OP_422J2_124_3477_n2120) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1351 ( .A1(DP_OP_424J2_126_3477_n2700), .A2(
        DP_OP_422J2_124_3477_n2138), .Y(DP_OP_422J2_124_3477_n2112) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1344 ( .A1(DP_OP_422J2_124_3477_n2129), 
        .A2(DP_OP_422J2_124_3477_n2137), .Y(DP_OP_422J2_124_3477_n2105) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1343 ( .A1(DP_OP_424J2_126_3477_n2700), .A2(
        DP_OP_422J2_124_3477_n2137), .Y(DP_OP_422J2_124_3477_n2104) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1342 ( .A1(DP_OP_422J2_124_3477_n2135), .A2(
        DP_OP_422J2_124_3477_n2136), .Y(DP_OP_422J2_124_3477_n2103) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1341 ( .A1(DP_OP_422J2_124_3477_n2134), .A2(
        DP_OP_422J2_124_3477_n2136), .Y(DP_OP_422J2_124_3477_n2102) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1340 ( .A1(DP_OP_424J2_126_3477_n2705), .A2(
        DP_OP_422J2_124_3477_n2136), .Y(DP_OP_422J2_124_3477_n2101) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1339 ( .A1(DP_OP_422J2_124_3477_n2132), .A2(
        DP_OP_422J2_124_3477_n2136), .Y(DP_OP_422J2_124_3477_n2100) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1338 ( .A1(DP_OP_424J2_126_3477_n2703), .A2(
        DP_OP_422J2_124_3477_n2136), .Y(DP_OP_422J2_124_3477_n2099) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1337 ( .A1(DP_OP_422J2_124_3477_n2130), .A2(
        DP_OP_422J2_124_3477_n2136), .Y(DP_OP_422J2_124_3477_n2098) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1336 ( .A1(DP_OP_422J2_124_3477_n2129), .A2(
        DP_OP_422J2_124_3477_n2136), .Y(DP_OP_422J2_124_3477_n2097) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1335 ( .A1(DP_OP_424J2_126_3477_n2700), 
        .A2(DP_OP_422J2_124_3477_n2136), .Y(DP_OP_422J2_124_3477_n2096) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1322 ( .A1(DP_OP_422J2_124_3477_n2091), 
        .A2(DP_OP_422J2_124_3477_n2095), .Y(DP_OP_422J2_124_3477_n2083) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1321 ( .A1(DP_OP_422J2_124_3477_n2090), 
        .A2(DP_OP_422J2_124_3477_n2095), .Y(DP_OP_422J2_124_3477_n2082) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1320 ( .A1(DP_OP_423J2_125_3477_n2837), 
        .A2(DP_OP_422J2_124_3477_n2095), .Y(DP_OP_422J2_124_3477_n2081) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1319 ( .A1(DP_OP_422J2_124_3477_n2088), 
        .A2(DP_OP_422J2_124_3477_n2095), .Y(DP_OP_422J2_124_3477_n2080) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1318 ( .A1(DP_OP_424J2_126_3477_n2747), 
        .A2(DP_OP_422J2_124_3477_n2095), .Y(DP_OP_422J2_124_3477_n2079) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1317 ( .A1(DP_OP_425J2_127_3477_n2218), 
        .A2(DP_OP_422J2_124_3477_n2095), .Y(DP_OP_422J2_124_3477_n2078) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1316 ( .A1(DP_OP_425J2_127_3477_n2217), 
        .A2(DP_OP_422J2_124_3477_n2095), .Y(DP_OP_422J2_124_3477_n2077) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1315 ( .A1(DP_OP_422J2_124_3477_n2084), .A2(
        DP_OP_422J2_124_3477_n2095), .Y(DP_OP_422J2_124_3477_n2076) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1314 ( .A1(DP_OP_422J2_124_3477_n2091), 
        .A2(DP_OP_422J2_124_3477_n2094), .Y(DP_OP_422J2_124_3477_n2075) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1313 ( .A1(DP_OP_422J2_124_3477_n2090), 
        .A2(DP_OP_422J2_124_3477_n2094), .Y(DP_OP_422J2_124_3477_n2074) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1312 ( .A1(DP_OP_424J2_126_3477_n2749), 
        .A2(DP_OP_422J2_124_3477_n2094), .Y(DP_OP_422J2_124_3477_n2073) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1311 ( .A1(DP_OP_422J2_124_3477_n2088), 
        .A2(DP_OP_422J2_124_3477_n2094), .Y(DP_OP_422J2_124_3477_n2072) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1310 ( .A1(DP_OP_425J2_127_3477_n2219), 
        .A2(DP_OP_422J2_124_3477_n2094), .Y(DP_OP_422J2_124_3477_n2071) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1309 ( .A1(DP_OP_425J2_127_3477_n2218), 
        .A2(DP_OP_422J2_124_3477_n2094), .Y(DP_OP_422J2_124_3477_n2070) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1308 ( .A1(DP_OP_424J2_126_3477_n2745), 
        .A2(DP_OP_422J2_124_3477_n2094), .Y(DP_OP_422J2_124_3477_n2069) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1307 ( .A1(DP_OP_422J2_124_3477_n2084), .A2(
        DP_OP_422J2_124_3477_n2094), .Y(DP_OP_422J2_124_3477_n2068) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1299 ( .A1(DP_OP_422J2_124_3477_n2084), .A2(
        DP_OP_422J2_124_3477_n2093), .Y(DP_OP_422J2_124_3477_n2060) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1298 ( .A1(DP_OP_422J2_124_3477_n2091), .A2(
        DP_OP_422J2_124_3477_n2092), .Y(DP_OP_422J2_124_3477_n2059) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1297 ( .A1(DP_OP_422J2_124_3477_n2090), .A2(
        DP_OP_422J2_124_3477_n2092), .Y(DP_OP_422J2_124_3477_n2058) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1296 ( .A1(DP_OP_423J2_125_3477_n2837), .A2(
        DP_OP_422J2_124_3477_n2092), .Y(DP_OP_422J2_124_3477_n2057) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1295 ( .A1(DP_OP_422J2_124_3477_n2088), .A2(
        DP_OP_422J2_124_3477_n2092), .Y(DP_OP_422J2_124_3477_n2056) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1294 ( .A1(DP_OP_425J2_127_3477_n2219), .A2(
        DP_OP_422J2_124_3477_n2092), .Y(DP_OP_422J2_124_3477_n2055) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1293 ( .A1(DP_OP_425J2_127_3477_n2218), .A2(
        DP_OP_422J2_124_3477_n2092), .Y(DP_OP_422J2_124_3477_n2054) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1292 ( .A1(DP_OP_424J2_126_3477_n2745), .A2(
        DP_OP_422J2_124_3477_n2092), .Y(DP_OP_422J2_124_3477_n2053) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1291 ( .A1(DP_OP_422J2_124_3477_n2084), 
        .A2(DP_OP_422J2_124_3477_n2092), .Y(DP_OP_422J2_124_3477_n2052) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1278 ( .A1(DP_OP_422J2_124_3477_n2047), 
        .A2(DP_OP_422J2_124_3477_n2051), .Y(DP_OP_422J2_124_3477_n2039) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1277 ( .A1(DP_OP_425J2_127_3477_n2178), 
        .A2(DP_OP_422J2_124_3477_n2051), .Y(DP_OP_422J2_124_3477_n2038) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1276 ( .A1(DP_OP_422J2_124_3477_n2045), 
        .A2(DP_OP_422J2_124_3477_n2051), .Y(DP_OP_422J2_124_3477_n2037) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1275 ( .A1(DP_OP_422J2_124_3477_n2044), 
        .A2(DP_OP_422J2_124_3477_n2051), .Y(DP_OP_422J2_124_3477_n2036) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1274 ( .A1(DP_OP_424J2_126_3477_n2791), 
        .A2(DP_OP_422J2_124_3477_n2051), .Y(DP_OP_422J2_124_3477_n2035) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1273 ( .A1(DP_OP_424J2_126_3477_n2790), 
        .A2(DP_OP_422J2_124_3477_n2051), .Y(DP_OP_422J2_124_3477_n2034) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1272 ( .A1(DP_OP_424J2_126_3477_n2789), 
        .A2(DP_OP_422J2_124_3477_n2051), .Y(DP_OP_422J2_124_3477_n2033) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1271 ( .A1(DP_OP_422J2_124_3477_n2040), .A2(
        DP_OP_422J2_124_3477_n2051), .Y(DP_OP_422J2_124_3477_n2032) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1263 ( .A1(DP_OP_422J2_124_3477_n2040), .A2(
        DP_OP_422J2_124_3477_n2050), .Y(DP_OP_422J2_124_3477_n2024) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1255 ( .A1(DP_OP_422J2_124_3477_n2040), .A2(
        DP_OP_422J2_124_3477_n2049), .Y(DP_OP_422J2_124_3477_n2016) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1254 ( .A1(DP_OP_422J2_124_3477_n2047), .A2(
        DP_OP_422J2_124_3477_n2048), .Y(DP_OP_422J2_124_3477_n2015) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1253 ( .A1(DP_OP_424J2_126_3477_n2794), .A2(
        DP_OP_422J2_124_3477_n2048), .Y(DP_OP_422J2_124_3477_n2014) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1252 ( .A1(DP_OP_422J2_124_3477_n2045), .A2(
        DP_OP_422J2_124_3477_n2048), .Y(DP_OP_422J2_124_3477_n2013) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1251 ( .A1(DP_OP_422J2_124_3477_n2044), .A2(
        DP_OP_422J2_124_3477_n2048), .Y(DP_OP_422J2_124_3477_n2012) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1250 ( .A1(DP_OP_424J2_126_3477_n2791), .A2(
        DP_OP_422J2_124_3477_n2048), .Y(DP_OP_422J2_124_3477_n2011) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1249 ( .A1(DP_OP_423J2_125_3477_n2878), .A2(
        DP_OP_422J2_124_3477_n2048), .Y(DP_OP_422J2_124_3477_n2010) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1248 ( .A1(DP_OP_423J2_125_3477_n2877), .A2(
        DP_OP_422J2_124_3477_n2048), .Y(DP_OP_422J2_124_3477_n2009) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1247 ( .A1(DP_OP_422J2_124_3477_n2040), 
        .A2(DP_OP_422J2_124_3477_n2048), .Y(DP_OP_422J2_124_3477_n2008) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1227 ( .A1(DP_OP_423J2_125_3477_n2920), .A2(
        DP_OP_422J2_124_3477_n2007), .Y(DP_OP_422J2_124_3477_n1988) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1219 ( .A1(DP_OP_425J2_127_3477_n2128), .A2(
        DP_OP_422J2_124_3477_n2006), .Y(DP_OP_422J2_124_3477_n1980) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1212 ( .A1(DP_OP_423J2_125_3477_n2921), 
        .A2(DP_OP_422J2_124_3477_n2005), .Y(DP_OP_422J2_124_3477_n1973) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1211 ( .A1(DP_OP_423J2_125_3477_n2920), .A2(
        DP_OP_422J2_124_3477_n2005), .Y(DP_OP_422J2_124_3477_n1972) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1210 ( .A1(DP_OP_425J2_127_3477_n2135), .A2(
        DP_OP_422J2_124_3477_n2004), .Y(DP_OP_422J2_124_3477_n1971) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1209 ( .A1(DP_OP_425J2_127_3477_n2134), .A2(
        DP_OP_422J2_124_3477_n2004), .Y(DP_OP_422J2_124_3477_n1970) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1208 ( .A1(DP_OP_425J2_127_3477_n2133), .A2(
        DP_OP_422J2_124_3477_n2004), .Y(DP_OP_422J2_124_3477_n1969) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1207 ( .A1(DP_OP_422J2_124_3477_n2000), .A2(
        DP_OP_422J2_124_3477_n2004), .Y(DP_OP_422J2_124_3477_n1968) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1206 ( .A1(DP_OP_424J2_126_3477_n2835), .A2(
        DP_OP_422J2_124_3477_n2004), .Y(DP_OP_422J2_124_3477_n1967) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1205 ( .A1(DP_OP_423J2_125_3477_n2922), .A2(
        DP_OP_422J2_124_3477_n2004), .Y(DP_OP_422J2_124_3477_n1966) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1204 ( .A1(DP_OP_423J2_125_3477_n2921), .A2(
        DP_OP_422J2_124_3477_n2004), .Y(DP_OP_422J2_124_3477_n1965) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1203 ( .A1(DP_OP_423J2_125_3477_n2920), 
        .A2(DP_OP_422J2_124_3477_n2004), .Y(DP_OP_422J2_124_3477_n1964) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1184 ( .A1(DP_OP_424J2_126_3477_n2877), 
        .A2(DP_OP_422J2_124_3477_n1963), .Y(DP_OP_422J2_124_3477_n1945) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1183 ( .A1(DP_OP_423J2_125_3477_n2964), .A2(
        DP_OP_422J2_124_3477_n1963), .Y(DP_OP_422J2_124_3477_n1944) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1175 ( .A1(DP_OP_425J2_127_3477_n2084), .A2(
        DP_OP_422J2_124_3477_n1962), .Y(DP_OP_422J2_124_3477_n1936) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1167 ( .A1(DP_OP_423J2_125_3477_n2964), .A2(
        DP_OP_422J2_124_3477_n1961), .Y(DP_OP_422J2_124_3477_n1928) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1166 ( .A1(DP_OP_423J2_125_3477_n2971), .A2(
        DP_OP_422J2_124_3477_n1960), .Y(DP_OP_422J2_124_3477_n1927) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1165 ( .A1(DP_OP_422J2_124_3477_n1958), .A2(
        DP_OP_422J2_124_3477_n1960), .Y(DP_OP_422J2_124_3477_n1926) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1164 ( .A1(DP_OP_422J2_124_3477_n1957), .A2(
        DP_OP_422J2_124_3477_n1960), .Y(DP_OP_422J2_124_3477_n1925) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1163 ( .A1(DP_OP_425J2_127_3477_n2088), .A2(
        DP_OP_422J2_124_3477_n1960), .Y(DP_OP_422J2_124_3477_n1924) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1162 ( .A1(DP_OP_423J2_125_3477_n2967), .A2(
        DP_OP_422J2_124_3477_n1960), .Y(DP_OP_422J2_124_3477_n1923) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1161 ( .A1(DP_OP_425J2_127_3477_n2086), .A2(
        DP_OP_422J2_124_3477_n1960), .Y(DP_OP_422J2_124_3477_n1922) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1160 ( .A1(DP_OP_425J2_127_3477_n2085), .A2(
        DP_OP_422J2_124_3477_n1960), .Y(DP_OP_422J2_124_3477_n1921) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1159 ( .A1(DP_OP_425J2_127_3477_n2084), 
        .A2(DP_OP_422J2_124_3477_n1960), .Y(DP_OP_422J2_124_3477_n1920) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1112 ( .A1(n505), .A2(n388), .Y(
        DP_OP_422J2_124_3477_n1874) );
  HADDX1_HVT DP_OP_422J2_124_3477_U1093 ( .A0(DP_OP_422J2_124_3477_n1886), 
        .B0(DP_OP_422J2_124_3477_n1995), .C1(DP_OP_422J2_124_3477_n1870), .SO(
        DP_OP_422J2_124_3477_n1871) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1092 ( .A(DP_OP_422J2_124_3477_n2039), .B(
        DP_OP_422J2_124_3477_n1951), .CI(DP_OP_422J2_124_3477_n2083), .CO(
        DP_OP_422J2_124_3477_n1868), .S(DP_OP_422J2_124_3477_n1869) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1091 ( .A(DP_OP_422J2_124_3477_n2171), .B(
        DP_OP_422J2_124_3477_n2127), .CI(DP_OP_422J2_124_3477_n2215), .CO(
        DP_OP_422J2_124_3477_n1866), .S(DP_OP_422J2_124_3477_n1867) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1090 ( .A(DP_OP_422J2_124_3477_n2303), .B(
        DP_OP_422J2_124_3477_n2259), .CI(DP_OP_422J2_124_3477_n2347), .CO(
        DP_OP_422J2_124_3477_n1864), .S(DP_OP_422J2_124_3477_n1865) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1089 ( .A(DP_OP_422J2_124_3477_n2435), .B(
        DP_OP_422J2_124_3477_n2391), .CI(DP_OP_422J2_124_3477_n2479), .CO(
        DP_OP_422J2_124_3477_n1862), .S(DP_OP_422J2_124_3477_n1863) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1088 ( .A(DP_OP_422J2_124_3477_n2567), .B(
        DP_OP_422J2_124_3477_n2523), .CI(DP_OP_422J2_124_3477_n2611), .CO(
        DP_OP_422J2_124_3477_n1860), .S(DP_OP_422J2_124_3477_n1861) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1087 ( .A(DP_OP_422J2_124_3477_n2699), .B(
        DP_OP_422J2_124_3477_n2655), .CI(DP_OP_422J2_124_3477_n2743), .CO(
        DP_OP_422J2_124_3477_n1858), .S(DP_OP_422J2_124_3477_n1859) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1086 ( .A(DP_OP_422J2_124_3477_n3005), .B(
        DP_OP_422J2_124_3477_n2787), .CI(DP_OP_422J2_124_3477_n2831), .CO(
        DP_OP_422J2_124_3477_n1856), .S(DP_OP_422J2_124_3477_n1857) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1085 ( .A(DP_OP_422J2_124_3477_n2963), .B(
        DP_OP_422J2_124_3477_n2875), .CI(DP_OP_422J2_124_3477_n2919), .CO(
        DP_OP_422J2_124_3477_n1854), .S(DP_OP_422J2_124_3477_n1855) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1084 ( .A(DP_OP_422J2_124_3477_n1871), .B(
        DP_OP_422J2_124_3477_n1857), .CI(DP_OP_422J2_124_3477_n1859), .CO(
        DP_OP_422J2_124_3477_n1852), .S(DP_OP_422J2_124_3477_n1853) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1083 ( .A(DP_OP_422J2_124_3477_n1861), .B(
        DP_OP_422J2_124_3477_n1855), .CI(DP_OP_422J2_124_3477_n1863), .CO(
        DP_OP_422J2_124_3477_n1850), .S(DP_OP_422J2_124_3477_n1851) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1082 ( .A(DP_OP_422J2_124_3477_n1869), .B(
        DP_OP_422J2_124_3477_n1865), .CI(DP_OP_422J2_124_3477_n1867), .CO(
        DP_OP_422J2_124_3477_n1848), .S(DP_OP_422J2_124_3477_n1849) );
  HADDX1_HVT DP_OP_422J2_124_3477_U1081 ( .A0(DP_OP_422J2_124_3477_n1885), 
        .B0(DP_OP_422J2_124_3477_n1950), .C1(DP_OP_422J2_124_3477_n1846), .SO(
        DP_OP_422J2_124_3477_n1847) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1080 ( .A(DP_OP_422J2_124_3477_n1987), .B(
        DP_OP_422J2_124_3477_n1943), .CI(DP_OP_422J2_124_3477_n1994), .CO(
        DP_OP_422J2_124_3477_n1844), .S(DP_OP_422J2_124_3477_n1845) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1079 ( .A(DP_OP_422J2_124_3477_n2038), .B(
        DP_OP_422J2_124_3477_n2031), .CI(DP_OP_422J2_124_3477_n2075), .CO(
        DP_OP_422J2_124_3477_n1842), .S(DP_OP_422J2_124_3477_n1843) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1078 ( .A(DP_OP_422J2_124_3477_n2119), .B(
        DP_OP_422J2_124_3477_n2082), .CI(DP_OP_422J2_124_3477_n2126), .CO(
        DP_OP_422J2_124_3477_n1840), .S(DP_OP_422J2_124_3477_n1841) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1077 ( .A(DP_OP_422J2_124_3477_n2170), .B(
        DP_OP_422J2_124_3477_n2163), .CI(DP_OP_422J2_124_3477_n2207), .CO(
        DP_OP_422J2_124_3477_n1838), .S(DP_OP_422J2_124_3477_n1839) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1076 ( .A(DP_OP_422J2_124_3477_n2251), .B(
        DP_OP_422J2_124_3477_n2214), .CI(DP_OP_422J2_124_3477_n2258), .CO(
        DP_OP_422J2_124_3477_n1836), .S(DP_OP_422J2_124_3477_n1837) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1075 ( .A(DP_OP_422J2_124_3477_n2302), .B(
        DP_OP_422J2_124_3477_n2295), .CI(DP_OP_422J2_124_3477_n2339), .CO(
        DP_OP_422J2_124_3477_n1834), .S(DP_OP_422J2_124_3477_n1835) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1074 ( .A(DP_OP_422J2_124_3477_n2383), .B(
        DP_OP_422J2_124_3477_n2346), .CI(DP_OP_422J2_124_3477_n2390), .CO(
        DP_OP_422J2_124_3477_n1832), .S(DP_OP_422J2_124_3477_n1833) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1073 ( .A(DP_OP_422J2_124_3477_n2434), .B(
        DP_OP_422J2_124_3477_n2427), .CI(DP_OP_422J2_124_3477_n2471), .CO(
        DP_OP_422J2_124_3477_n1830), .S(DP_OP_422J2_124_3477_n1831) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1072 ( .A(DP_OP_422J2_124_3477_n2515), .B(
        DP_OP_422J2_124_3477_n2478), .CI(DP_OP_422J2_124_3477_n2522), .CO(
        DP_OP_422J2_124_3477_n1828), .S(DP_OP_422J2_124_3477_n1829) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1071 ( .A(DP_OP_422J2_124_3477_n3004), .B(
        DP_OP_422J2_124_3477_n2559), .CI(DP_OP_422J2_124_3477_n2997), .CO(
        DP_OP_422J2_124_3477_n1826), .S(DP_OP_422J2_124_3477_n1827) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1070 ( .A(DP_OP_422J2_124_3477_n2742), .B(
        DP_OP_422J2_124_3477_n2566), .CI(DP_OP_422J2_124_3477_n2603), .CO(
        DP_OP_422J2_124_3477_n1824), .S(DP_OP_422J2_124_3477_n1825) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1069 ( .A(DP_OP_422J2_124_3477_n2779), .B(
        DP_OP_422J2_124_3477_n2962), .CI(DP_OP_422J2_124_3477_n2955), .CO(
        DP_OP_422J2_124_3477_n1822), .S(DP_OP_422J2_124_3477_n1823) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1068 ( .A(DP_OP_422J2_124_3477_n2698), .B(
        DP_OP_422J2_124_3477_n2918), .CI(DP_OP_422J2_124_3477_n2911), .CO(
        DP_OP_422J2_124_3477_n1820), .S(DP_OP_422J2_124_3477_n1821) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1067 ( .A(DP_OP_422J2_124_3477_n2691), .B(
        DP_OP_422J2_124_3477_n2874), .CI(DP_OP_422J2_124_3477_n2610), .CO(
        DP_OP_422J2_124_3477_n1818), .S(DP_OP_422J2_124_3477_n1819) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1066 ( .A(DP_OP_422J2_124_3477_n2867), .B(
        DP_OP_422J2_124_3477_n2647), .CI(DP_OP_422J2_124_3477_n2654), .CO(
        DP_OP_422J2_124_3477_n1816), .S(DP_OP_422J2_124_3477_n1817) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1065 ( .A(DP_OP_422J2_124_3477_n2823), .B(
        DP_OP_422J2_124_3477_n2735), .CI(DP_OP_422J2_124_3477_n2786), .CO(
        DP_OP_422J2_124_3477_n1814), .S(DP_OP_422J2_124_3477_n1815) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1064 ( .A(DP_OP_422J2_124_3477_n2830), .B(
        DP_OP_422J2_124_3477_n1870), .CI(DP_OP_422J2_124_3477_n1847), .CO(
        DP_OP_422J2_124_3477_n1812), .S(DP_OP_422J2_124_3477_n1813) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1063 ( .A(DP_OP_422J2_124_3477_n1854), .B(
        DP_OP_422J2_124_3477_n1868), .CI(DP_OP_422J2_124_3477_n1866), .CO(
        DP_OP_422J2_124_3477_n1810), .S(DP_OP_422J2_124_3477_n1811) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1062 ( .A(DP_OP_422J2_124_3477_n1860), .B(
        DP_OP_422J2_124_3477_n1856), .CI(DP_OP_422J2_124_3477_n1864), .CO(
        DP_OP_422J2_124_3477_n1808), .S(DP_OP_422J2_124_3477_n1809) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1061 ( .A(DP_OP_422J2_124_3477_n1862), .B(
        DP_OP_422J2_124_3477_n1858), .CI(DP_OP_422J2_124_3477_n1815), .CO(
        DP_OP_422J2_124_3477_n1806), .S(DP_OP_422J2_124_3477_n1807) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1060 ( .A(DP_OP_422J2_124_3477_n1837), .B(
        DP_OP_422J2_124_3477_n1823), .CI(DP_OP_422J2_124_3477_n1821), .CO(
        DP_OP_422J2_124_3477_n1804), .S(DP_OP_422J2_124_3477_n1805) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1059 ( .A(DP_OP_422J2_124_3477_n1841), .B(
        DP_OP_422J2_124_3477_n1825), .CI(DP_OP_422J2_124_3477_n1829), .CO(
        DP_OP_422J2_124_3477_n1802), .S(DP_OP_422J2_124_3477_n1803) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1058 ( .A(DP_OP_422J2_124_3477_n1843), .B(
        DP_OP_422J2_124_3477_n1831), .CI(DP_OP_422J2_124_3477_n1827), .CO(
        DP_OP_422J2_124_3477_n1800), .S(DP_OP_422J2_124_3477_n1801) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1057 ( .A(DP_OP_422J2_124_3477_n1845), .B(
        DP_OP_422J2_124_3477_n1835), .CI(DP_OP_422J2_124_3477_n1819), .CO(
        DP_OP_422J2_124_3477_n1798), .S(DP_OP_422J2_124_3477_n1799) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1056 ( .A(DP_OP_422J2_124_3477_n1839), .B(
        DP_OP_422J2_124_3477_n1833), .CI(DP_OP_422J2_124_3477_n1817), .CO(
        DP_OP_422J2_124_3477_n1796), .S(DP_OP_422J2_124_3477_n1797) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1055 ( .A(DP_OP_422J2_124_3477_n1813), .B(
        DP_OP_422J2_124_3477_n1852), .CI(DP_OP_422J2_124_3477_n1850), .CO(
        DP_OP_422J2_124_3477_n1794), .S(DP_OP_422J2_124_3477_n1795) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1054 ( .A(DP_OP_422J2_124_3477_n1848), .B(
        DP_OP_422J2_124_3477_n1809), .CI(DP_OP_422J2_124_3477_n1811), .CO(
        DP_OP_422J2_124_3477_n1792), .S(DP_OP_422J2_124_3477_n1793) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1053 ( .A(DP_OP_422J2_124_3477_n1807), .B(
        DP_OP_422J2_124_3477_n1799), .CI(DP_OP_422J2_124_3477_n1801), .CO(
        DP_OP_422J2_124_3477_n1790), .S(DP_OP_422J2_124_3477_n1791) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1052 ( .A(DP_OP_422J2_124_3477_n1805), .B(
        DP_OP_422J2_124_3477_n1797), .CI(DP_OP_422J2_124_3477_n1803), .CO(
        DP_OP_422J2_124_3477_n1788), .S(DP_OP_422J2_124_3477_n1789) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1051 ( .A(DP_OP_422J2_124_3477_n1795), .B(
        DP_OP_422J2_124_3477_n1793), .CI(DP_OP_422J2_124_3477_n1791), .CO(
        DP_OP_422J2_124_3477_n1786), .S(DP_OP_422J2_124_3477_n1787) );
  HADDX1_HVT DP_OP_422J2_124_3477_U1050 ( .A0(DP_OP_422J2_124_3477_n1884), 
        .B0(DP_OP_422J2_124_3477_n1949), .C1(DP_OP_422J2_124_3477_n1784), .SO(
        DP_OP_422J2_124_3477_n1785) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1049 ( .A(DP_OP_422J2_124_3477_n1979), .B(
        DP_OP_422J2_124_3477_n1942), .CI(DP_OP_422J2_124_3477_n1935), .CO(
        DP_OP_422J2_124_3477_n1782), .S(DP_OP_422J2_124_3477_n1783) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1048 ( .A(DP_OP_422J2_124_3477_n1993), .B(
        DP_OP_422J2_124_3477_n1986), .CI(DP_OP_422J2_124_3477_n2023), .CO(
        DP_OP_422J2_124_3477_n1780), .S(DP_OP_422J2_124_3477_n1781) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1047 ( .A(DP_OP_422J2_124_3477_n2037), .B(
        DP_OP_422J2_124_3477_n2030), .CI(DP_OP_422J2_124_3477_n2067), .CO(
        DP_OP_422J2_124_3477_n1778), .S(DP_OP_422J2_124_3477_n1779) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1046 ( .A(DP_OP_422J2_124_3477_n2081), .B(
        DP_OP_422J2_124_3477_n2074), .CI(DP_OP_422J2_124_3477_n2111), .CO(
        DP_OP_422J2_124_3477_n1776), .S(DP_OP_422J2_124_3477_n1777) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1045 ( .A(DP_OP_422J2_124_3477_n2125), .B(
        DP_OP_422J2_124_3477_n2118), .CI(DP_OP_422J2_124_3477_n2155), .CO(
        DP_OP_422J2_124_3477_n1774), .S(DP_OP_422J2_124_3477_n1775) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1044 ( .A(DP_OP_422J2_124_3477_n2169), .B(
        DP_OP_422J2_124_3477_n2162), .CI(DP_OP_422J2_124_3477_n2199), .CO(
        DP_OP_422J2_124_3477_n1772), .S(DP_OP_422J2_124_3477_n1773) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1043 ( .A(DP_OP_422J2_124_3477_n2213), .B(
        DP_OP_422J2_124_3477_n2206), .CI(DP_OP_422J2_124_3477_n2243), .CO(
        DP_OP_422J2_124_3477_n1770), .S(DP_OP_422J2_124_3477_n1771) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1042 ( .A(DP_OP_422J2_124_3477_n2257), .B(
        DP_OP_422J2_124_3477_n2250), .CI(DP_OP_422J2_124_3477_n2287), .CO(
        DP_OP_422J2_124_3477_n1768), .S(DP_OP_422J2_124_3477_n1769) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1041 ( .A(DP_OP_422J2_124_3477_n2301), .B(
        DP_OP_422J2_124_3477_n2294), .CI(DP_OP_422J2_124_3477_n2331), .CO(
        DP_OP_422J2_124_3477_n1766), .S(DP_OP_422J2_124_3477_n1767) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1040 ( .A(DP_OP_422J2_124_3477_n2345), .B(
        DP_OP_422J2_124_3477_n2338), .CI(DP_OP_422J2_124_3477_n2375), .CO(
        DP_OP_422J2_124_3477_n1764), .S(DP_OP_422J2_124_3477_n1765) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1039 ( .A(DP_OP_422J2_124_3477_n2389), .B(
        DP_OP_422J2_124_3477_n2382), .CI(DP_OP_422J2_124_3477_n2419), .CO(
        DP_OP_422J2_124_3477_n1762), .S(DP_OP_422J2_124_3477_n1763) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1038 ( .A(DP_OP_422J2_124_3477_n2690), .B(
        DP_OP_422J2_124_3477_n3003), .CI(DP_OP_422J2_124_3477_n2996), .CO(
        DP_OP_422J2_124_3477_n1760), .S(DP_OP_422J2_124_3477_n1761) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1037 ( .A(DP_OP_422J2_124_3477_n2653), .B(
        DP_OP_422J2_124_3477_n2426), .CI(DP_OP_422J2_124_3477_n2989), .CO(
        DP_OP_422J2_124_3477_n1758), .S(DP_OP_422J2_124_3477_n1759) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1036 ( .A(DP_OP_422J2_124_3477_n2646), .B(
        DP_OP_422J2_124_3477_n2961), .CI(DP_OP_422J2_124_3477_n2433), .CO(
        DP_OP_422J2_124_3477_n1756), .S(DP_OP_422J2_124_3477_n1757) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1035 ( .A(DP_OP_422J2_124_3477_n2683), .B(
        DP_OP_422J2_124_3477_n2463), .CI(DP_OP_422J2_124_3477_n2470), .CO(
        DP_OP_422J2_124_3477_n1754), .S(DP_OP_422J2_124_3477_n1755) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1034 ( .A(DP_OP_422J2_124_3477_n2697), .B(
        DP_OP_422J2_124_3477_n2477), .CI(DP_OP_422J2_124_3477_n2954), .CO(
        DP_OP_422J2_124_3477_n1752), .S(DP_OP_422J2_124_3477_n1753) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1033 ( .A(DP_OP_422J2_124_3477_n2727), .B(
        DP_OP_422J2_124_3477_n2507), .CI(DP_OP_422J2_124_3477_n2947), .CO(
        DP_OP_422J2_124_3477_n1750), .S(DP_OP_422J2_124_3477_n1751) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1032 ( .A(DP_OP_422J2_124_3477_n2639), .B(
        DP_OP_422J2_124_3477_n2514), .CI(DP_OP_422J2_124_3477_n2917), .CO(
        DP_OP_422J2_124_3477_n1748), .S(DP_OP_422J2_124_3477_n1749) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1031 ( .A(DP_OP_422J2_124_3477_n2609), .B(
        DP_OP_422J2_124_3477_n2521), .CI(DP_OP_422J2_124_3477_n2910), .CO(
        DP_OP_422J2_124_3477_n1746), .S(DP_OP_422J2_124_3477_n1747) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1030 ( .A(DP_OP_422J2_124_3477_n2903), .B(
        DP_OP_422J2_124_3477_n2551), .CI(DP_OP_422J2_124_3477_n2558), .CO(
        DP_OP_422J2_124_3477_n1744), .S(DP_OP_422J2_124_3477_n1745) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1029 ( .A(DP_OP_422J2_124_3477_n2873), .B(
        DP_OP_422J2_124_3477_n2565), .CI(DP_OP_422J2_124_3477_n2595), .CO(
        DP_OP_422J2_124_3477_n1742), .S(DP_OP_422J2_124_3477_n1743) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1028 ( .A(DP_OP_422J2_124_3477_n2866), .B(
        DP_OP_422J2_124_3477_n2602), .CI(DP_OP_422J2_124_3477_n2734), .CO(
        DP_OP_422J2_124_3477_n1740), .S(DP_OP_422J2_124_3477_n1741) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1027 ( .A(DP_OP_422J2_124_3477_n2859), .B(
        DP_OP_422J2_124_3477_n2741), .CI(DP_OP_422J2_124_3477_n2771), .CO(
        DP_OP_422J2_124_3477_n1738), .S(DP_OP_422J2_124_3477_n1739) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1026 ( .A(DP_OP_422J2_124_3477_n2829), .B(
        DP_OP_422J2_124_3477_n2778), .CI(DP_OP_422J2_124_3477_n2785), .CO(
        DP_OP_422J2_124_3477_n1736), .S(DP_OP_422J2_124_3477_n1737) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1025 ( .A(DP_OP_422J2_124_3477_n2822), .B(
        DP_OP_422J2_124_3477_n2815), .CI(DP_OP_422J2_124_3477_n1846), .CO(
        DP_OP_422J2_124_3477_n1734), .S(DP_OP_422J2_124_3477_n1735) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1024 ( .A(DP_OP_422J2_124_3477_n1785), .B(
        DP_OP_422J2_124_3477_n1814), .CI(DP_OP_422J2_124_3477_n1816), .CO(
        DP_OP_422J2_124_3477_n1732), .S(DP_OP_422J2_124_3477_n1733) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1023 ( .A(DP_OP_422J2_124_3477_n1832), .B(
        DP_OP_422J2_124_3477_n1844), .CI(DP_OP_422J2_124_3477_n1818), .CO(
        DP_OP_422J2_124_3477_n1730), .S(DP_OP_422J2_124_3477_n1731) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1022 ( .A(DP_OP_422J2_124_3477_n1830), .B(
        DP_OP_422J2_124_3477_n1842), .CI(DP_OP_422J2_124_3477_n1820), .CO(
        DP_OP_422J2_124_3477_n1728), .S(DP_OP_422J2_124_3477_n1729) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1021 ( .A(DP_OP_422J2_124_3477_n1826), .B(
        DP_OP_422J2_124_3477_n1840), .CI(DP_OP_422J2_124_3477_n1822), .CO(
        DP_OP_422J2_124_3477_n1726), .S(DP_OP_422J2_124_3477_n1727) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1020 ( .A(DP_OP_422J2_124_3477_n1838), .B(
        DP_OP_422J2_124_3477_n1836), .CI(DP_OP_422J2_124_3477_n1834), .CO(
        DP_OP_422J2_124_3477_n1724), .S(DP_OP_422J2_124_3477_n1725) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1019 ( .A(DP_OP_422J2_124_3477_n1828), .B(
        DP_OP_422J2_124_3477_n1824), .CI(DP_OP_422J2_124_3477_n1757), .CO(
        DP_OP_422J2_124_3477_n1722), .S(DP_OP_422J2_124_3477_n1723) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1018 ( .A(DP_OP_422J2_124_3477_n1751), .B(
        DP_OP_422J2_124_3477_n1765), .CI(DP_OP_422J2_124_3477_n1769), .CO(
        DP_OP_422J2_124_3477_n1720), .S(DP_OP_422J2_124_3477_n1721) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1017 ( .A(DP_OP_422J2_124_3477_n1747), .B(
        DP_OP_422J2_124_3477_n1775), .CI(DP_OP_422J2_124_3477_n1777), .CO(
        DP_OP_422J2_124_3477_n1718), .S(DP_OP_422J2_124_3477_n1719) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1016 ( .A(DP_OP_422J2_124_3477_n1745), .B(
        DP_OP_422J2_124_3477_n1767), .CI(DP_OP_422J2_124_3477_n1781), .CO(
        DP_OP_422J2_124_3477_n1716), .S(DP_OP_422J2_124_3477_n1717) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1015 ( .A(DP_OP_422J2_124_3477_n1743), .B(
        DP_OP_422J2_124_3477_n1761), .CI(DP_OP_422J2_124_3477_n1779), .CO(
        DP_OP_422J2_124_3477_n1714), .S(DP_OP_422J2_124_3477_n1715) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1014 ( .A(DP_OP_422J2_124_3477_n1741), .B(
        DP_OP_422J2_124_3477_n1771), .CI(DP_OP_422J2_124_3477_n1759), .CO(
        DP_OP_422J2_124_3477_n1712), .S(DP_OP_422J2_124_3477_n1713) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1013 ( .A(DP_OP_422J2_124_3477_n1739), .B(
        DP_OP_422J2_124_3477_n1773), .CI(DP_OP_422J2_124_3477_n1783), .CO(
        DP_OP_422J2_124_3477_n1710), .S(DP_OP_422J2_124_3477_n1711) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1012 ( .A(DP_OP_422J2_124_3477_n1737), .B(
        DP_OP_422J2_124_3477_n1763), .CI(DP_OP_422J2_124_3477_n1749), .CO(
        DP_OP_422J2_124_3477_n1708), .S(DP_OP_422J2_124_3477_n1709) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1011 ( .A(DP_OP_422J2_124_3477_n1755), .B(
        DP_OP_422J2_124_3477_n1753), .CI(DP_OP_422J2_124_3477_n1812), .CO(
        DP_OP_422J2_124_3477_n1706), .S(DP_OP_422J2_124_3477_n1707) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1010 ( .A(DP_OP_422J2_124_3477_n1735), .B(
        DP_OP_422J2_124_3477_n1810), .CI(DP_OP_422J2_124_3477_n1808), .CO(
        DP_OP_422J2_124_3477_n1704), .S(DP_OP_422J2_124_3477_n1705) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1009 ( .A(DP_OP_422J2_124_3477_n1806), .B(
        DP_OP_422J2_124_3477_n1733), .CI(DP_OP_422J2_124_3477_n1800), .CO(
        DP_OP_422J2_124_3477_n1702), .S(DP_OP_422J2_124_3477_n1703) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1008 ( .A(DP_OP_422J2_124_3477_n1804), .B(
        DP_OP_422J2_124_3477_n1725), .CI(DP_OP_422J2_124_3477_n1731), .CO(
        DP_OP_422J2_124_3477_n1700), .S(DP_OP_422J2_124_3477_n1701) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1007 ( .A(DP_OP_422J2_124_3477_n1802), .B(
        DP_OP_422J2_124_3477_n1729), .CI(DP_OP_422J2_124_3477_n1727), .CO(
        DP_OP_422J2_124_3477_n1698), .S(DP_OP_422J2_124_3477_n1699) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1006 ( .A(DP_OP_422J2_124_3477_n1798), .B(
        DP_OP_422J2_124_3477_n1796), .CI(DP_OP_422J2_124_3477_n1723), .CO(
        DP_OP_422J2_124_3477_n1696), .S(DP_OP_422J2_124_3477_n1697) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1005 ( .A(DP_OP_422J2_124_3477_n1721), .B(
        DP_OP_422J2_124_3477_n1709), .CI(DP_OP_422J2_124_3477_n1707), .CO(
        DP_OP_422J2_124_3477_n1694), .S(DP_OP_422J2_124_3477_n1695) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1004 ( .A(DP_OP_422J2_124_3477_n1711), .B(
        DP_OP_422J2_124_3477_n1719), .CI(DP_OP_422J2_124_3477_n1717), .CO(
        DP_OP_422J2_124_3477_n1692), .S(DP_OP_422J2_124_3477_n1693) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1003 ( .A(DP_OP_422J2_124_3477_n1713), .B(
        DP_OP_422J2_124_3477_n1715), .CI(DP_OP_422J2_124_3477_n1794), .CO(
        DP_OP_422J2_124_3477_n1690), .S(DP_OP_422J2_124_3477_n1691) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1002 ( .A(DP_OP_422J2_124_3477_n1705), .B(
        DP_OP_422J2_124_3477_n1792), .CI(DP_OP_422J2_124_3477_n1703), .CO(
        DP_OP_422J2_124_3477_n1688), .S(DP_OP_422J2_124_3477_n1689) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1001 ( .A(DP_OP_422J2_124_3477_n1790), .B(
        DP_OP_422J2_124_3477_n1788), .CI(DP_OP_422J2_124_3477_n1699), .CO(
        DP_OP_422J2_124_3477_n1686), .S(DP_OP_422J2_124_3477_n1687) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1000 ( .A(DP_OP_422J2_124_3477_n1701), .B(
        DP_OP_422J2_124_3477_n1697), .CI(DP_OP_422J2_124_3477_n1695), .CO(
        DP_OP_422J2_124_3477_n1684), .S(DP_OP_422J2_124_3477_n1685) );
  FADDX1_HVT DP_OP_422J2_124_3477_U999 ( .A(DP_OP_422J2_124_3477_n1693), .B(
        DP_OP_422J2_124_3477_n1691), .CI(DP_OP_422J2_124_3477_n1689), .CO(
        DP_OP_422J2_124_3477_n1682), .S(DP_OP_422J2_124_3477_n1683) );
  FADDX1_HVT DP_OP_422J2_124_3477_U998 ( .A(DP_OP_422J2_124_3477_n1786), .B(
        DP_OP_422J2_124_3477_n1687), .CI(DP_OP_422J2_124_3477_n1685), .CO(
        DP_OP_422J2_124_3477_n1680), .S(DP_OP_422J2_124_3477_n1681) );
  FADDX1_HVT DP_OP_422J2_124_3477_U996 ( .A(DP_OP_422J2_124_3477_n2455), .B(
        DP_OP_422J2_124_3477_n1927), .CI(DP_OP_422J2_124_3477_n1883), .CO(
        DP_OP_422J2_124_3477_n1676), .S(DP_OP_422J2_124_3477_n1677) );
  FADDX1_HVT DP_OP_422J2_124_3477_U995 ( .A(DP_OP_422J2_124_3477_n2147), .B(
        DP_OP_422J2_124_3477_n2587), .CI(DP_OP_422J2_124_3477_n2367), .CO(
        DP_OP_422J2_124_3477_n1674), .S(DP_OP_422J2_124_3477_n1675) );
  FADDX1_HVT DP_OP_422J2_124_3477_U994 ( .A(DP_OP_422J2_124_3477_n2895), .B(
        DP_OP_422J2_124_3477_n2103), .CI(DP_OP_422J2_124_3477_n2323), .CO(
        DP_OP_422J2_124_3477_n1672), .S(DP_OP_422J2_124_3477_n1673) );
  FADDX1_HVT DP_OP_422J2_124_3477_U993 ( .A(DP_OP_422J2_124_3477_n2499), .B(
        DP_OP_422J2_124_3477_n2807), .CI(DP_OP_422J2_124_3477_n2411), .CO(
        DP_OP_422J2_124_3477_n1670), .S(DP_OP_422J2_124_3477_n1671) );
  FADDX1_HVT DP_OP_422J2_124_3477_U992 ( .A(DP_OP_422J2_124_3477_n2235), .B(
        DP_OP_422J2_124_3477_n2279), .CI(DP_OP_422J2_124_3477_n2059), .CO(
        DP_OP_422J2_124_3477_n1668), .S(DP_OP_422J2_124_3477_n1669) );
  FADDX1_HVT DP_OP_422J2_124_3477_U991 ( .A(DP_OP_422J2_124_3477_n2763), .B(
        DP_OP_422J2_124_3477_n2631), .CI(DP_OP_422J2_124_3477_n2675), .CO(
        DP_OP_422J2_124_3477_n1666), .S(DP_OP_422J2_124_3477_n1667) );
  FADDX1_HVT DP_OP_422J2_124_3477_U990 ( .A(DP_OP_422J2_124_3477_n2015), .B(
        DP_OP_422J2_124_3477_n2851), .CI(DP_OP_422J2_124_3477_n2719), .CO(
        DP_OP_422J2_124_3477_n1664), .S(DP_OP_422J2_124_3477_n1665) );
  FADDX1_HVT DP_OP_422J2_124_3477_U989 ( .A(DP_OP_422J2_124_3477_n2543), .B(
        DP_OP_422J2_124_3477_n2939), .CI(DP_OP_422J2_124_3477_n2191), .CO(
        DP_OP_422J2_124_3477_n1662), .S(DP_OP_422J2_124_3477_n1663) );
  FADDX1_HVT DP_OP_422J2_124_3477_U988 ( .A(DP_OP_422J2_124_3477_n1971), .B(
        DP_OP_422J2_124_3477_n1679), .CI(DP_OP_422J2_124_3477_n1948), .CO(
        DP_OP_422J2_124_3477_n1660), .S(DP_OP_422J2_124_3477_n1661) );
  FADDX1_HVT DP_OP_422J2_124_3477_U987 ( .A(DP_OP_422J2_124_3477_n1978), .B(
        DP_OP_422J2_124_3477_n1941), .CI(DP_OP_422J2_124_3477_n1934), .CO(
        DP_OP_422J2_124_3477_n1658), .S(DP_OP_422J2_124_3477_n1659) );
  FADDX1_HVT DP_OP_422J2_124_3477_U986 ( .A(DP_OP_422J2_124_3477_n1992), .B(
        DP_OP_422J2_124_3477_n1985), .CI(DP_OP_422J2_124_3477_n2022), .CO(
        DP_OP_422J2_124_3477_n1656), .S(DP_OP_422J2_124_3477_n1657) );
  FADDX1_HVT DP_OP_422J2_124_3477_U985 ( .A(DP_OP_422J2_124_3477_n2036), .B(
        DP_OP_422J2_124_3477_n2029), .CI(DP_OP_422J2_124_3477_n2066), .CO(
        DP_OP_422J2_124_3477_n1654), .S(DP_OP_422J2_124_3477_n1655) );
  FADDX1_HVT DP_OP_422J2_124_3477_U984 ( .A(DP_OP_422J2_124_3477_n3002), .B(
        DP_OP_422J2_124_3477_n2073), .CI(DP_OP_422J2_124_3477_n2080), .CO(
        DP_OP_422J2_124_3477_n1652), .S(DP_OP_422J2_124_3477_n1653) );
  FADDX1_HVT DP_OP_422J2_124_3477_U983 ( .A(DP_OP_422J2_124_3477_n2513), .B(
        DP_OP_422J2_124_3477_n2995), .CI(DP_OP_422J2_124_3477_n2988), .CO(
        DP_OP_422J2_124_3477_n1650), .S(DP_OP_422J2_124_3477_n1651) );
  FADDX1_HVT DP_OP_422J2_124_3477_U982 ( .A(DP_OP_422J2_124_3477_n2476), .B(
        DP_OP_422J2_124_3477_n2110), .CI(DP_OP_422J2_124_3477_n2960), .CO(
        DP_OP_422J2_124_3477_n1648), .S(DP_OP_422J2_124_3477_n1649) );
  FADDX1_HVT DP_OP_422J2_124_3477_U981 ( .A(DP_OP_422J2_124_3477_n2506), .B(
        DP_OP_422J2_124_3477_n2117), .CI(DP_OP_422J2_124_3477_n2953), .CO(
        DP_OP_422J2_124_3477_n1646), .S(DP_OP_422J2_124_3477_n1647) );
  FADDX1_HVT DP_OP_422J2_124_3477_U980 ( .A(DP_OP_422J2_124_3477_n2946), .B(
        DP_OP_422J2_124_3477_n2124), .CI(DP_OP_422J2_124_3477_n2154), .CO(
        DP_OP_422J2_124_3477_n1644), .S(DP_OP_422J2_124_3477_n1645) );
  FADDX1_HVT DP_OP_422J2_124_3477_U979 ( .A(DP_OP_422J2_124_3477_n2469), .B(
        DP_OP_422J2_124_3477_n2161), .CI(DP_OP_422J2_124_3477_n2168), .CO(
        DP_OP_422J2_124_3477_n1642), .S(DP_OP_422J2_124_3477_n1643) );
  FADDX1_HVT DP_OP_422J2_124_3477_U978 ( .A(DP_OP_422J2_124_3477_n2550), .B(
        DP_OP_422J2_124_3477_n2198), .CI(DP_OP_422J2_124_3477_n2205), .CO(
        DP_OP_422J2_124_3477_n1640), .S(DP_OP_422J2_124_3477_n1641) );
  FADDX1_HVT DP_OP_422J2_124_3477_U977 ( .A(DP_OP_422J2_124_3477_n2557), .B(
        DP_OP_422J2_124_3477_n2212), .CI(DP_OP_422J2_124_3477_n2242), .CO(
        DP_OP_422J2_124_3477_n1638), .S(DP_OP_422J2_124_3477_n1639) );
  FADDX1_HVT DP_OP_422J2_124_3477_U976 ( .A(DP_OP_422J2_124_3477_n2564), .B(
        DP_OP_422J2_124_3477_n2916), .CI(DP_OP_422J2_124_3477_n2249), .CO(
        DP_OP_422J2_124_3477_n1636), .S(DP_OP_422J2_124_3477_n1637) );
  FADDX1_HVT DP_OP_422J2_124_3477_U975 ( .A(DP_OP_422J2_124_3477_n2594), .B(
        DP_OP_422J2_124_3477_n2256), .CI(DP_OP_422J2_124_3477_n2909), .CO(
        DP_OP_422J2_124_3477_n1634), .S(DP_OP_422J2_124_3477_n1635) );
  FADDX1_HVT DP_OP_422J2_124_3477_U974 ( .A(DP_OP_422J2_124_3477_n2520), .B(
        DP_OP_422J2_124_3477_n2902), .CI(DP_OP_422J2_124_3477_n2872), .CO(
        DP_OP_422J2_124_3477_n1632), .S(DP_OP_422J2_124_3477_n1633) );
  FADDX1_HVT DP_OP_422J2_124_3477_U973 ( .A(DP_OP_422J2_124_3477_n2432), .B(
        DP_OP_422J2_124_3477_n2865), .CI(DP_OP_422J2_124_3477_n2286), .CO(
        DP_OP_422J2_124_3477_n1630), .S(DP_OP_422J2_124_3477_n1631) );
  FADDX1_HVT DP_OP_422J2_124_3477_U972 ( .A(DP_OP_422J2_124_3477_n2858), .B(
        DP_OP_422J2_124_3477_n2293), .CI(DP_OP_422J2_124_3477_n2828), .CO(
        DP_OP_422J2_124_3477_n1628), .S(DP_OP_422J2_124_3477_n1629) );
  FADDX1_HVT DP_OP_422J2_124_3477_U971 ( .A(DP_OP_422J2_124_3477_n2821), .B(
        DP_OP_422J2_124_3477_n2814), .CI(DP_OP_422J2_124_3477_n2300), .CO(
        DP_OP_422J2_124_3477_n1626), .S(DP_OP_422J2_124_3477_n1627) );
  FADDX1_HVT DP_OP_422J2_124_3477_U970 ( .A(DP_OP_422J2_124_3477_n2425), .B(
        DP_OP_422J2_124_3477_n2330), .CI(DP_OP_422J2_124_3477_n2784), .CO(
        DP_OP_422J2_124_3477_n1624), .S(DP_OP_422J2_124_3477_n1625) );
  FADDX1_HVT DP_OP_422J2_124_3477_U969 ( .A(DP_OP_422J2_124_3477_n2418), .B(
        DP_OP_422J2_124_3477_n2777), .CI(DP_OP_422J2_124_3477_n2770), .CO(
        DP_OP_422J2_124_3477_n1622), .S(DP_OP_422J2_124_3477_n1623) );
  FADDX1_HVT DP_OP_422J2_124_3477_U968 ( .A(DP_OP_422J2_124_3477_n2374), .B(
        DP_OP_422J2_124_3477_n2740), .CI(DP_OP_422J2_124_3477_n2733), .CO(
        DP_OP_422J2_124_3477_n1620), .S(DP_OP_422J2_124_3477_n1621) );
  FADDX1_HVT DP_OP_422J2_124_3477_U967 ( .A(DP_OP_422J2_124_3477_n2337), .B(
        DP_OP_422J2_124_3477_n2726), .CI(DP_OP_422J2_124_3477_n2696), .CO(
        DP_OP_422J2_124_3477_n1618), .S(DP_OP_422J2_124_3477_n1619) );
  FADDX1_HVT DP_OP_422J2_124_3477_U966 ( .A(DP_OP_422J2_124_3477_n2608), .B(
        DP_OP_422J2_124_3477_n2689), .CI(DP_OP_422J2_124_3477_n2344), .CO(
        DP_OP_422J2_124_3477_n1616), .S(DP_OP_422J2_124_3477_n1617) );
  FADDX1_HVT DP_OP_422J2_124_3477_U965 ( .A(DP_OP_422J2_124_3477_n2462), .B(
        DP_OP_422J2_124_3477_n2381), .CI(DP_OP_422J2_124_3477_n2682), .CO(
        DP_OP_422J2_124_3477_n1614), .S(DP_OP_422J2_124_3477_n1615) );
  FADDX1_HVT DP_OP_422J2_124_3477_U964 ( .A(DP_OP_422J2_124_3477_n2652), .B(
        DP_OP_422J2_124_3477_n2388), .CI(DP_OP_422J2_124_3477_n2601), .CO(
        DP_OP_422J2_124_3477_n1612), .S(DP_OP_422J2_124_3477_n1613) );
  FADDX1_HVT DP_OP_422J2_124_3477_U963 ( .A(DP_OP_422J2_124_3477_n2645), .B(
        DP_OP_422J2_124_3477_n2638), .CI(DP_OP_422J2_124_3477_n1784), .CO(
        DP_OP_422J2_124_3477_n1610), .S(DP_OP_422J2_124_3477_n1611) );
  FADDX1_HVT DP_OP_422J2_124_3477_U962 ( .A(DP_OP_422J2_124_3477_n1760), .B(
        DP_OP_422J2_124_3477_n1782), .CI(DP_OP_422J2_124_3477_n1736), .CO(
        DP_OP_422J2_124_3477_n1608), .S(DP_OP_422J2_124_3477_n1609) );
  FADDX1_HVT DP_OP_422J2_124_3477_U961 ( .A(DP_OP_422J2_124_3477_n1758), .B(
        DP_OP_422J2_124_3477_n1780), .CI(DP_OP_422J2_124_3477_n1778), .CO(
        DP_OP_422J2_124_3477_n1606), .S(DP_OP_422J2_124_3477_n1607) );
  FADDX1_HVT DP_OP_422J2_124_3477_U960 ( .A(DP_OP_422J2_124_3477_n1752), .B(
        DP_OP_422J2_124_3477_n1776), .CI(DP_OP_422J2_124_3477_n1774), .CO(
        DP_OP_422J2_124_3477_n1604), .S(DP_OP_422J2_124_3477_n1605) );
  FADDX1_HVT DP_OP_422J2_124_3477_U959 ( .A(DP_OP_422J2_124_3477_n1748), .B(
        DP_OP_422J2_124_3477_n1738), .CI(DP_OP_422J2_124_3477_n1740), .CO(
        DP_OP_422J2_124_3477_n1602), .S(DP_OP_422J2_124_3477_n1603) );
  FADDX1_HVT DP_OP_422J2_124_3477_U958 ( .A(DP_OP_422J2_124_3477_n1746), .B(
        DP_OP_422J2_124_3477_n1772), .CI(DP_OP_422J2_124_3477_n1742), .CO(
        DP_OP_422J2_124_3477_n1600), .S(DP_OP_422J2_124_3477_n1601) );
  FADDX1_HVT DP_OP_422J2_124_3477_U957 ( .A(DP_OP_422J2_124_3477_n1744), .B(
        DP_OP_422J2_124_3477_n1770), .CI(DP_OP_422J2_124_3477_n1768), .CO(
        DP_OP_422J2_124_3477_n1598), .S(DP_OP_422J2_124_3477_n1599) );
  FADDX1_HVT DP_OP_422J2_124_3477_U956 ( .A(DP_OP_422J2_124_3477_n1756), .B(
        DP_OP_422J2_124_3477_n1766), .CI(DP_OP_422J2_124_3477_n1750), .CO(
        DP_OP_422J2_124_3477_n1596), .S(DP_OP_422J2_124_3477_n1597) );
  FADDX1_HVT DP_OP_422J2_124_3477_U955 ( .A(DP_OP_422J2_124_3477_n1764), .B(
        DP_OP_422J2_124_3477_n1762), .CI(DP_OP_422J2_124_3477_n1754), .CO(
        DP_OP_422J2_124_3477_n1594), .S(DP_OP_422J2_124_3477_n1595) );
  FADDX1_HVT DP_OP_422J2_124_3477_U954 ( .A(DP_OP_422J2_124_3477_n1673), .B(
        DP_OP_422J2_124_3477_n1675), .CI(DP_OP_422J2_124_3477_n1661), .CO(
        DP_OP_422J2_124_3477_n1592), .S(DP_OP_422J2_124_3477_n1593) );
  FADDX1_HVT DP_OP_422J2_124_3477_U953 ( .A(DP_OP_422J2_124_3477_n1667), .B(
        DP_OP_422J2_124_3477_n1669), .CI(DP_OP_422J2_124_3477_n1734), .CO(
        DP_OP_422J2_124_3477_n1590), .S(DP_OP_422J2_124_3477_n1591) );
  FADDX1_HVT DP_OP_422J2_124_3477_U952 ( .A(DP_OP_422J2_124_3477_n1663), .B(
        DP_OP_422J2_124_3477_n1665), .CI(DP_OP_422J2_124_3477_n1671), .CO(
        DP_OP_422J2_124_3477_n1588), .S(DP_OP_422J2_124_3477_n1589) );
  FADDX1_HVT DP_OP_422J2_124_3477_U951 ( .A(DP_OP_422J2_124_3477_n1677), .B(
        DP_OP_422J2_124_3477_n1627), .CI(DP_OP_422J2_124_3477_n1625), .CO(
        DP_OP_422J2_124_3477_n1586), .S(DP_OP_422J2_124_3477_n1587) );
  FADDX1_HVT DP_OP_422J2_124_3477_U950 ( .A(DP_OP_422J2_124_3477_n1629), .B(
        DP_OP_422J2_124_3477_n1645), .CI(DP_OP_422J2_124_3477_n1653), .CO(
        DP_OP_422J2_124_3477_n1584), .S(DP_OP_422J2_124_3477_n1585) );
  FADDX1_HVT DP_OP_422J2_124_3477_U949 ( .A(DP_OP_422J2_124_3477_n1621), .B(
        DP_OP_422J2_124_3477_n1641), .CI(DP_OP_422J2_124_3477_n1639), .CO(
        DP_OP_422J2_124_3477_n1582), .S(DP_OP_422J2_124_3477_n1583) );
  FADDX1_HVT DP_OP_422J2_124_3477_U948 ( .A(DP_OP_422J2_124_3477_n1619), .B(
        DP_OP_422J2_124_3477_n1655), .CI(DP_OP_422J2_124_3477_n1643), .CO(
        DP_OP_422J2_124_3477_n1580), .S(DP_OP_422J2_124_3477_n1581) );
  FADDX1_HVT DP_OP_422J2_124_3477_U947 ( .A(DP_OP_422J2_124_3477_n1617), .B(
        DP_OP_422J2_124_3477_n1649), .CI(DP_OP_422J2_124_3477_n1651), .CO(
        DP_OP_422J2_124_3477_n1578), .S(DP_OP_422J2_124_3477_n1579) );
  FADDX1_HVT DP_OP_422J2_124_3477_U946 ( .A(DP_OP_422J2_124_3477_n1615), .B(
        DP_OP_422J2_124_3477_n1647), .CI(DP_OP_422J2_124_3477_n1659), .CO(
        DP_OP_422J2_124_3477_n1576), .S(DP_OP_422J2_124_3477_n1577) );
  FADDX1_HVT DP_OP_422J2_124_3477_U945 ( .A(DP_OP_422J2_124_3477_n1637), .B(
        DP_OP_422J2_124_3477_n1657), .CI(DP_OP_422J2_124_3477_n1613), .CO(
        DP_OP_422J2_124_3477_n1574), .S(DP_OP_422J2_124_3477_n1575) );
  FADDX1_HVT DP_OP_422J2_124_3477_U944 ( .A(DP_OP_422J2_124_3477_n1623), .B(
        DP_OP_422J2_124_3477_n1633), .CI(DP_OP_422J2_124_3477_n1635), .CO(
        DP_OP_422J2_124_3477_n1572), .S(DP_OP_422J2_124_3477_n1573) );
  FADDX1_HVT DP_OP_422J2_124_3477_U943 ( .A(DP_OP_422J2_124_3477_n1631), .B(
        DP_OP_422J2_124_3477_n1611), .CI(DP_OP_422J2_124_3477_n1732), .CO(
        DP_OP_422J2_124_3477_n1570), .S(DP_OP_422J2_124_3477_n1571) );
  FADDX1_HVT DP_OP_422J2_124_3477_U942 ( .A(DP_OP_422J2_124_3477_n1730), .B(
        DP_OP_422J2_124_3477_n1728), .CI(DP_OP_422J2_124_3477_n1726), .CO(
        DP_OP_422J2_124_3477_n1568), .S(DP_OP_422J2_124_3477_n1569) );
  FADDX1_HVT DP_OP_422J2_124_3477_U941 ( .A(DP_OP_422J2_124_3477_n1724), .B(
        DP_OP_422J2_124_3477_n1722), .CI(DP_OP_422J2_124_3477_n1710), .CO(
        DP_OP_422J2_124_3477_n1566), .S(DP_OP_422J2_124_3477_n1567) );
  FADDX1_HVT DP_OP_422J2_124_3477_U940 ( .A(DP_OP_422J2_124_3477_n1708), .B(
        DP_OP_422J2_124_3477_n1609), .CI(DP_OP_422J2_124_3477_n1706), .CO(
        DP_OP_422J2_124_3477_n1564), .S(DP_OP_422J2_124_3477_n1565) );
  FADDX1_HVT DP_OP_422J2_124_3477_U939 ( .A(DP_OP_422J2_124_3477_n1720), .B(
        DP_OP_422J2_124_3477_n1599), .CI(DP_OP_422J2_124_3477_n1607), .CO(
        DP_OP_422J2_124_3477_n1562), .S(DP_OP_422J2_124_3477_n1563) );
  FADDX1_HVT DP_OP_422J2_124_3477_U938 ( .A(DP_OP_422J2_124_3477_n1718), .B(
        DP_OP_422J2_124_3477_n1597), .CI(DP_OP_422J2_124_3477_n1601), .CO(
        DP_OP_422J2_124_3477_n1560), .S(DP_OP_422J2_124_3477_n1561) );
  FADDX1_HVT DP_OP_422J2_124_3477_U937 ( .A(DP_OP_422J2_124_3477_n1714), .B(
        DP_OP_422J2_124_3477_n1605), .CI(DP_OP_422J2_124_3477_n1603), .CO(
        DP_OP_422J2_124_3477_n1558), .S(DP_OP_422J2_124_3477_n1559) );
  FADDX1_HVT DP_OP_422J2_124_3477_U936 ( .A(DP_OP_422J2_124_3477_n1712), .B(
        DP_OP_422J2_124_3477_n1716), .CI(DP_OP_422J2_124_3477_n1595), .CO(
        DP_OP_422J2_124_3477_n1556), .S(DP_OP_422J2_124_3477_n1557) );
  FADDX1_HVT DP_OP_422J2_124_3477_U935 ( .A(DP_OP_422J2_124_3477_n1591), .B(
        DP_OP_422J2_124_3477_n1593), .CI(DP_OP_422J2_124_3477_n1587), .CO(
        DP_OP_422J2_124_3477_n1554), .S(DP_OP_422J2_124_3477_n1555) );
  FADDX1_HVT DP_OP_422J2_124_3477_U934 ( .A(DP_OP_422J2_124_3477_n1589), .B(
        DP_OP_422J2_124_3477_n1575), .CI(DP_OP_422J2_124_3477_n1577), .CO(
        DP_OP_422J2_124_3477_n1552), .S(DP_OP_422J2_124_3477_n1553) );
  FADDX1_HVT DP_OP_422J2_124_3477_U933 ( .A(DP_OP_422J2_124_3477_n1583), .B(
        DP_OP_422J2_124_3477_n1581), .CI(DP_OP_422J2_124_3477_n1704), .CO(
        DP_OP_422J2_124_3477_n1550), .S(DP_OP_422J2_124_3477_n1551) );
  FADDX1_HVT DP_OP_422J2_124_3477_U932 ( .A(DP_OP_422J2_124_3477_n1579), .B(
        DP_OP_422J2_124_3477_n1573), .CI(DP_OP_422J2_124_3477_n1585), .CO(
        DP_OP_422J2_124_3477_n1548), .S(DP_OP_422J2_124_3477_n1549) );
  FADDX1_HVT DP_OP_422J2_124_3477_U931 ( .A(DP_OP_422J2_124_3477_n1571), .B(
        DP_OP_422J2_124_3477_n1702), .CI(DP_OP_422J2_124_3477_n1698), .CO(
        DP_OP_422J2_124_3477_n1546), .S(DP_OP_422J2_124_3477_n1547) );
  FADDX1_HVT DP_OP_422J2_124_3477_U930 ( .A(DP_OP_422J2_124_3477_n1700), .B(
        DP_OP_422J2_124_3477_n1569), .CI(DP_OP_422J2_124_3477_n1696), .CO(
        DP_OP_422J2_124_3477_n1544), .S(DP_OP_422J2_124_3477_n1545) );
  FADDX1_HVT DP_OP_422J2_124_3477_U929 ( .A(DP_OP_422J2_124_3477_n1567), .B(
        DP_OP_422J2_124_3477_n1557), .CI(DP_OP_422J2_124_3477_n1559), .CO(
        DP_OP_422J2_124_3477_n1542), .S(DP_OP_422J2_124_3477_n1543) );
  FADDX1_HVT DP_OP_422J2_124_3477_U928 ( .A(DP_OP_422J2_124_3477_n1694), .B(
        DP_OP_422J2_124_3477_n1561), .CI(DP_OP_422J2_124_3477_n1692), .CO(
        DP_OP_422J2_124_3477_n1540), .S(DP_OP_422J2_124_3477_n1541) );
  FADDX1_HVT DP_OP_422J2_124_3477_U927 ( .A(DP_OP_422J2_124_3477_n1565), .B(
        DP_OP_422J2_124_3477_n1563), .CI(DP_OP_422J2_124_3477_n1555), .CO(
        DP_OP_422J2_124_3477_n1538), .S(DP_OP_422J2_124_3477_n1539) );
  FADDX1_HVT DP_OP_422J2_124_3477_U926 ( .A(DP_OP_422J2_124_3477_n1690), .B(
        DP_OP_422J2_124_3477_n1553), .CI(DP_OP_422J2_124_3477_n1549), .CO(
        DP_OP_422J2_124_3477_n1536), .S(DP_OP_422J2_124_3477_n1537) );
  FADDX1_HVT DP_OP_422J2_124_3477_U925 ( .A(DP_OP_422J2_124_3477_n1551), .B(
        DP_OP_422J2_124_3477_n1688), .CI(DP_OP_422J2_124_3477_n1547), .CO(
        DP_OP_422J2_124_3477_n1534), .S(DP_OP_422J2_124_3477_n1535) );
  FADDX1_HVT DP_OP_422J2_124_3477_U924 ( .A(DP_OP_422J2_124_3477_n1686), .B(
        DP_OP_422J2_124_3477_n1545), .CI(DP_OP_422J2_124_3477_n1684), .CO(
        DP_OP_422J2_124_3477_n1532), .S(DP_OP_422J2_124_3477_n1533) );
  FADDX1_HVT DP_OP_422J2_124_3477_U923 ( .A(DP_OP_422J2_124_3477_n1543), .B(
        DP_OP_422J2_124_3477_n1541), .CI(DP_OP_422J2_124_3477_n1539), .CO(
        DP_OP_422J2_124_3477_n1530), .S(DP_OP_422J2_124_3477_n1531) );
  FADDX1_HVT DP_OP_422J2_124_3477_U922 ( .A(DP_OP_422J2_124_3477_n1537), .B(
        DP_OP_422J2_124_3477_n1682), .CI(DP_OP_422J2_124_3477_n1535), .CO(
        DP_OP_422J2_124_3477_n1528), .S(DP_OP_422J2_124_3477_n1529) );
  FADDX1_HVT DP_OP_422J2_124_3477_U921 ( .A(DP_OP_422J2_124_3477_n1680), .B(
        DP_OP_422J2_124_3477_n1533), .CI(DP_OP_422J2_124_3477_n1531), .CO(
        DP_OP_422J2_124_3477_n1526), .S(DP_OP_422J2_124_3477_n1527) );
  FADDX1_HVT DP_OP_422J2_124_3477_U920 ( .A(DP_OP_422J2_124_3477_n1678), .B(
        DP_OP_422J2_124_3477_n1926), .CI(DP_OP_422J2_124_3477_n1882), .CO(
        DP_OP_422J2_124_3477_n1524), .S(DP_OP_422J2_124_3477_n1525) );
  FADDX1_HVT DP_OP_422J2_124_3477_U919 ( .A(DP_OP_422J2_124_3477_n2981), .B(
        DP_OP_422J2_124_3477_n2498), .CI(DP_OP_422J2_124_3477_n2366), .CO(
        DP_OP_422J2_124_3477_n1522), .S(DP_OP_422J2_124_3477_n1523) );
  FADDX1_HVT DP_OP_422J2_124_3477_U918 ( .A(DP_OP_422J2_124_3477_n2894), .B(
        DP_OP_422J2_124_3477_n2630), .CI(DP_OP_422J2_124_3477_n2278), .CO(
        DP_OP_422J2_124_3477_n1520), .S(DP_OP_422J2_124_3477_n1521) );
  FADDX1_HVT DP_OP_422J2_124_3477_U917 ( .A(DP_OP_422J2_124_3477_n2058), .B(
        DP_OP_422J2_124_3477_n2586), .CI(DP_OP_422J2_124_3477_n2806), .CO(
        DP_OP_422J2_124_3477_n1518), .S(DP_OP_422J2_124_3477_n1519) );
  FADDX1_HVT DP_OP_422J2_124_3477_U916 ( .A(DP_OP_422J2_124_3477_n2146), .B(
        DP_OP_422J2_124_3477_n2322), .CI(DP_OP_422J2_124_3477_n2410), .CO(
        DP_OP_422J2_124_3477_n1516), .S(DP_OP_422J2_124_3477_n1517) );
  FADDX1_HVT DP_OP_422J2_124_3477_U915 ( .A(DP_OP_422J2_124_3477_n2762), .B(
        DP_OP_422J2_124_3477_n2234), .CI(DP_OP_422J2_124_3477_n2850), .CO(
        DP_OP_422J2_124_3477_n1514), .S(DP_OP_422J2_124_3477_n1515) );
  FADDX1_HVT DP_OP_422J2_124_3477_U914 ( .A(DP_OP_422J2_124_3477_n2102), .B(
        DP_OP_422J2_124_3477_n2454), .CI(DP_OP_422J2_124_3477_n2542), .CO(
        DP_OP_422J2_124_3477_n1512), .S(DP_OP_422J2_124_3477_n1513) );
  FADDX1_HVT DP_OP_422J2_124_3477_U913 ( .A(DP_OP_422J2_124_3477_n2938), .B(
        DP_OP_422J2_124_3477_n2674), .CI(DP_OP_422J2_124_3477_n2718), .CO(
        DP_OP_422J2_124_3477_n1510), .S(DP_OP_422J2_124_3477_n1511) );
  FADDX1_HVT DP_OP_422J2_124_3477_U912 ( .A(DP_OP_422J2_124_3477_n2014), .B(
        DP_OP_422J2_124_3477_n2190), .CI(DP_OP_422J2_124_3477_n1970), .CO(
        DP_OP_422J2_124_3477_n1508), .S(DP_OP_422J2_124_3477_n1509) );
  FADDX1_HVT DP_OP_422J2_124_3477_U911 ( .A(DP_OP_422J2_124_3477_n2505), .B(
        DP_OP_422J2_124_3477_n1940), .CI(DP_OP_422J2_124_3477_n1933), .CO(
        DP_OP_422J2_124_3477_n1506), .S(DP_OP_422J2_124_3477_n1507) );
  FADDX1_HVT DP_OP_422J2_124_3477_U910 ( .A(DP_OP_422J2_124_3477_n3001), .B(
        DP_OP_422J2_124_3477_n1947), .CI(DP_OP_422J2_124_3477_n1977), .CO(
        DP_OP_422J2_124_3477_n1504), .S(DP_OP_422J2_124_3477_n1505) );
  FADDX1_HVT DP_OP_422J2_124_3477_U909 ( .A(DP_OP_422J2_124_3477_n2387), .B(
        DP_OP_422J2_124_3477_n2994), .CI(DP_OP_422J2_124_3477_n1984), .CO(
        DP_OP_422J2_124_3477_n1502), .S(DP_OP_422J2_124_3477_n1503) );
  FADDX1_HVT DP_OP_422J2_124_3477_U908 ( .A(DP_OP_422J2_124_3477_n2380), .B(
        DP_OP_422J2_124_3477_n2987), .CI(DP_OP_422J2_124_3477_n1991), .CO(
        DP_OP_422J2_124_3477_n1500), .S(DP_OP_422J2_124_3477_n1501) );
  FADDX1_HVT DP_OP_422J2_124_3477_U907 ( .A(DP_OP_422J2_124_3477_n2959), .B(
        DP_OP_422J2_124_3477_n2021), .CI(DP_OP_422J2_124_3477_n2028), .CO(
        DP_OP_422J2_124_3477_n1498), .S(DP_OP_422J2_124_3477_n1499) );
  FADDX1_HVT DP_OP_422J2_124_3477_U906 ( .A(DP_OP_422J2_124_3477_n2417), .B(
        DP_OP_422J2_124_3477_n2952), .CI(DP_OP_422J2_124_3477_n2945), .CO(
        DP_OP_422J2_124_3477_n1496), .S(DP_OP_422J2_124_3477_n1497) );
  FADDX1_HVT DP_OP_422J2_124_3477_U905 ( .A(DP_OP_422J2_124_3477_n2343), .B(
        DP_OP_422J2_124_3477_n2915), .CI(DP_OP_422J2_124_3477_n2908), .CO(
        DP_OP_422J2_124_3477_n1494), .S(DP_OP_422J2_124_3477_n1495) );
  FADDX1_HVT DP_OP_422J2_124_3477_U904 ( .A(DP_OP_422J2_124_3477_n2336), .B(
        DP_OP_422J2_124_3477_n2901), .CI(DP_OP_422J2_124_3477_n2035), .CO(
        DP_OP_422J2_124_3477_n1492), .S(DP_OP_422J2_124_3477_n1493) );
  FADDX1_HVT DP_OP_422J2_124_3477_U903 ( .A(DP_OP_422J2_124_3477_n2329), .B(
        DP_OP_422J2_124_3477_n2871), .CI(DP_OP_422J2_124_3477_n2864), .CO(
        DP_OP_422J2_124_3477_n1490), .S(DP_OP_422J2_124_3477_n1491) );
  FADDX1_HVT DP_OP_422J2_124_3477_U902 ( .A(DP_OP_422J2_124_3477_n2299), .B(
        DP_OP_422J2_124_3477_n2857), .CI(DP_OP_422J2_124_3477_n2065), .CO(
        DP_OP_422J2_124_3477_n1488), .S(DP_OP_422J2_124_3477_n1489) );
  FADDX1_HVT DP_OP_422J2_124_3477_U901 ( .A(DP_OP_422J2_124_3477_n2292), .B(
        DP_OP_422J2_124_3477_n2072), .CI(DP_OP_422J2_124_3477_n2079), .CO(
        DP_OP_422J2_124_3477_n1486), .S(DP_OP_422J2_124_3477_n1487) );
  FADDX1_HVT DP_OP_422J2_124_3477_U900 ( .A(DP_OP_422J2_124_3477_n2373), .B(
        DP_OP_422J2_124_3477_n2109), .CI(DP_OP_422J2_124_3477_n2827), .CO(
        DP_OP_422J2_124_3477_n1484), .S(DP_OP_422J2_124_3477_n1485) );
  FADDX1_HVT DP_OP_422J2_124_3477_U899 ( .A(DP_OP_422J2_124_3477_n2424), .B(
        DP_OP_422J2_124_3477_n2820), .CI(DP_OP_422J2_124_3477_n2813), .CO(
        DP_OP_422J2_124_3477_n1482), .S(DP_OP_422J2_124_3477_n1483) );
  FADDX1_HVT DP_OP_422J2_124_3477_U898 ( .A(DP_OP_422J2_124_3477_n2783), .B(
        DP_OP_422J2_124_3477_n2116), .CI(DP_OP_422J2_124_3477_n2123), .CO(
        DP_OP_422J2_124_3477_n1480), .S(DP_OP_422J2_124_3477_n1481) );
  FADDX1_HVT DP_OP_422J2_124_3477_U897 ( .A(DP_OP_422J2_124_3477_n2556), .B(
        DP_OP_422J2_124_3477_n2153), .CI(DP_OP_422J2_124_3477_n2160), .CO(
        DP_OP_422J2_124_3477_n1478), .S(DP_OP_422J2_124_3477_n1479) );
  FADDX1_HVT DP_OP_422J2_124_3477_U896 ( .A(DP_OP_422J2_124_3477_n2776), .B(
        DP_OP_422J2_124_3477_n2167), .CI(DP_OP_422J2_124_3477_n2197), .CO(
        DP_OP_422J2_124_3477_n1476), .S(DP_OP_422J2_124_3477_n1477) );
  FADDX1_HVT DP_OP_422J2_124_3477_U895 ( .A(DP_OP_422J2_124_3477_n2769), .B(
        DP_OP_422J2_124_3477_n2204), .CI(DP_OP_422J2_124_3477_n2211), .CO(
        DP_OP_422J2_124_3477_n1474), .S(DP_OP_422J2_124_3477_n1475) );
  FADDX1_HVT DP_OP_422J2_124_3477_U894 ( .A(DP_OP_422J2_124_3477_n2739), .B(
        DP_OP_422J2_124_3477_n2241), .CI(DP_OP_422J2_124_3477_n2248), .CO(
        DP_OP_422J2_124_3477_n1472), .S(DP_OP_422J2_124_3477_n1473) );
  FADDX1_HVT DP_OP_422J2_124_3477_U893 ( .A(DP_OP_422J2_124_3477_n2732), .B(
        DP_OP_422J2_124_3477_n2255), .CI(DP_OP_422J2_124_3477_n2285), .CO(
        DP_OP_422J2_124_3477_n1470), .S(DP_OP_422J2_124_3477_n1471) );
  FADDX1_HVT DP_OP_422J2_124_3477_U892 ( .A(DP_OP_422J2_124_3477_n2725), .B(
        DP_OP_422J2_124_3477_n2431), .CI(DP_OP_422J2_124_3477_n2461), .CO(
        DP_OP_422J2_124_3477_n1468), .S(DP_OP_422J2_124_3477_n1469) );
  FADDX1_HVT DP_OP_422J2_124_3477_U891 ( .A(DP_OP_422J2_124_3477_n2695), .B(
        DP_OP_422J2_124_3477_n2468), .CI(DP_OP_422J2_124_3477_n2688), .CO(
        DP_OP_422J2_124_3477_n1466), .S(DP_OP_422J2_124_3477_n1467) );
  FADDX1_HVT DP_OP_422J2_124_3477_U890 ( .A(DP_OP_422J2_124_3477_n2593), .B(
        DP_OP_422J2_124_3477_n2475), .CI(DP_OP_422J2_124_3477_n2512), .CO(
        DP_OP_422J2_124_3477_n1464), .S(DP_OP_422J2_124_3477_n1465) );
  FADDX1_HVT DP_OP_422J2_124_3477_U889 ( .A(DP_OP_422J2_124_3477_n2563), .B(
        DP_OP_422J2_124_3477_n2519), .CI(DP_OP_422J2_124_3477_n2681), .CO(
        DP_OP_422J2_124_3477_n1462), .S(DP_OP_422J2_124_3477_n1463) );
  FADDX1_HVT DP_OP_422J2_124_3477_U888 ( .A(DP_OP_422J2_124_3477_n2637), .B(
        DP_OP_422J2_124_3477_n2549), .CI(DP_OP_422J2_124_3477_n2651), .CO(
        DP_OP_422J2_124_3477_n1460), .S(DP_OP_422J2_124_3477_n1461) );
  FADDX1_HVT DP_OP_422J2_124_3477_U887 ( .A(DP_OP_422J2_124_3477_n2600), .B(
        DP_OP_422J2_124_3477_n2607), .CI(DP_OP_422J2_124_3477_n2644), .CO(
        DP_OP_422J2_124_3477_n1458), .S(DP_OP_422J2_124_3477_n1459) );
  FADDX1_HVT DP_OP_422J2_124_3477_U886 ( .A(DP_OP_422J2_124_3477_n1666), .B(
        DP_OP_422J2_124_3477_n1662), .CI(DP_OP_422J2_124_3477_n1660), .CO(
        DP_OP_422J2_124_3477_n1456), .S(DP_OP_422J2_124_3477_n1457) );
  FADDX1_HVT DP_OP_422J2_124_3477_U885 ( .A(DP_OP_422J2_124_3477_n1664), .B(
        DP_OP_422J2_124_3477_n1668), .CI(DP_OP_422J2_124_3477_n1670), .CO(
        DP_OP_422J2_124_3477_n1454), .S(DP_OP_422J2_124_3477_n1455) );
  FADDX1_HVT DP_OP_422J2_124_3477_U884 ( .A(DP_OP_422J2_124_3477_n1672), .B(
        DP_OP_422J2_124_3477_n1674), .CI(DP_OP_422J2_124_3477_n1676), .CO(
        DP_OP_422J2_124_3477_n1452), .S(DP_OP_422J2_124_3477_n1453) );
  FADDX1_HVT DP_OP_422J2_124_3477_U883 ( .A(DP_OP_422J2_124_3477_n1636), .B(
        DP_OP_422J2_124_3477_n1658), .CI(DP_OP_422J2_124_3477_n1656), .CO(
        DP_OP_422J2_124_3477_n1450), .S(DP_OP_422J2_124_3477_n1451) );
  FADDX1_HVT DP_OP_422J2_124_3477_U882 ( .A(DP_OP_422J2_124_3477_n1632), .B(
        DP_OP_422J2_124_3477_n1654), .CI(DP_OP_422J2_124_3477_n1652), .CO(
        DP_OP_422J2_124_3477_n1448), .S(DP_OP_422J2_124_3477_n1449) );
  FADDX1_HVT DP_OP_422J2_124_3477_U881 ( .A(DP_OP_422J2_124_3477_n1626), .B(
        DP_OP_422J2_124_3477_n1650), .CI(DP_OP_422J2_124_3477_n1648), .CO(
        DP_OP_422J2_124_3477_n1446), .S(DP_OP_422J2_124_3477_n1447) );
  FADDX1_HVT DP_OP_422J2_124_3477_U880 ( .A(DP_OP_422J2_124_3477_n1622), .B(
        DP_OP_422J2_124_3477_n1646), .CI(DP_OP_422J2_124_3477_n1612), .CO(
        DP_OP_422J2_124_3477_n1444), .S(DP_OP_422J2_124_3477_n1445) );
  FADDX1_HVT DP_OP_422J2_124_3477_U879 ( .A(DP_OP_422J2_124_3477_n1618), .B(
        DP_OP_422J2_124_3477_n1644), .CI(DP_OP_422J2_124_3477_n1642), .CO(
        DP_OP_422J2_124_3477_n1442), .S(DP_OP_422J2_124_3477_n1443) );
  FADDX1_HVT DP_OP_422J2_124_3477_U878 ( .A(DP_OP_422J2_124_3477_n1628), .B(
        DP_OP_422J2_124_3477_n1640), .CI(DP_OP_422J2_124_3477_n1638), .CO(
        DP_OP_422J2_124_3477_n1440), .S(DP_OP_422J2_124_3477_n1441) );
  FADDX1_HVT DP_OP_422J2_124_3477_U877 ( .A(DP_OP_422J2_124_3477_n1620), .B(
        DP_OP_422J2_124_3477_n1634), .CI(DP_OP_422J2_124_3477_n1630), .CO(
        DP_OP_422J2_124_3477_n1438), .S(DP_OP_422J2_124_3477_n1439) );
  FADDX1_HVT DP_OP_422J2_124_3477_U876 ( .A(DP_OP_422J2_124_3477_n1616), .B(
        DP_OP_422J2_124_3477_n1624), .CI(DP_OP_422J2_124_3477_n1614), .CO(
        DP_OP_422J2_124_3477_n1436), .S(DP_OP_422J2_124_3477_n1437) );
  FADDX1_HVT DP_OP_422J2_124_3477_U875 ( .A(DP_OP_422J2_124_3477_n1525), .B(
        DP_OP_422J2_124_3477_n1509), .CI(DP_OP_422J2_124_3477_n1610), .CO(
        DP_OP_422J2_124_3477_n1434), .S(DP_OP_422J2_124_3477_n1435) );
  FADDX1_HVT DP_OP_422J2_124_3477_U874 ( .A(DP_OP_422J2_124_3477_n1523), .B(
        DP_OP_422J2_124_3477_n1511), .CI(DP_OP_422J2_124_3477_n1513), .CO(
        DP_OP_422J2_124_3477_n1432), .S(DP_OP_422J2_124_3477_n1433) );
  FADDX1_HVT DP_OP_422J2_124_3477_U873 ( .A(DP_OP_422J2_124_3477_n1519), .B(
        DP_OP_422J2_124_3477_n1517), .CI(DP_OP_422J2_124_3477_n1521), .CO(
        DP_OP_422J2_124_3477_n1430), .S(DP_OP_422J2_124_3477_n1431) );
  FADDX1_HVT DP_OP_422J2_124_3477_U872 ( .A(DP_OP_422J2_124_3477_n1515), .B(
        DP_OP_422J2_124_3477_n1495), .CI(DP_OP_422J2_124_3477_n1499), .CO(
        DP_OP_422J2_124_3477_n1428), .S(DP_OP_422J2_124_3477_n1429) );
  FADDX1_HVT DP_OP_422J2_124_3477_U871 ( .A(DP_OP_422J2_124_3477_n1497), .B(
        DP_OP_422J2_124_3477_n1505), .CI(DP_OP_422J2_124_3477_n1503), .CO(
        DP_OP_422J2_124_3477_n1426), .S(DP_OP_422J2_124_3477_n1427) );
  FADDX1_HVT DP_OP_422J2_124_3477_U870 ( .A(DP_OP_422J2_124_3477_n1507), .B(
        DP_OP_422J2_124_3477_n1485), .CI(DP_OP_422J2_124_3477_n1479), .CO(
        DP_OP_422J2_124_3477_n1424), .S(DP_OP_422J2_124_3477_n1425) );
  FADDX1_HVT DP_OP_422J2_124_3477_U869 ( .A(DP_OP_422J2_124_3477_n1487), .B(
        DP_OP_422J2_124_3477_n1483), .CI(DP_OP_422J2_124_3477_n1477), .CO(
        DP_OP_422J2_124_3477_n1422), .S(DP_OP_422J2_124_3477_n1423) );
  FADDX1_HVT DP_OP_422J2_124_3477_U868 ( .A(DP_OP_422J2_124_3477_n1489), .B(
        DP_OP_422J2_124_3477_n1463), .CI(DP_OP_422J2_124_3477_n1461), .CO(
        DP_OP_422J2_124_3477_n1420), .S(DP_OP_422J2_124_3477_n1421) );
  FADDX1_HVT DP_OP_422J2_124_3477_U867 ( .A(DP_OP_422J2_124_3477_n1475), .B(
        DP_OP_422J2_124_3477_n1471), .CI(DP_OP_422J2_124_3477_n1473), .CO(
        DP_OP_422J2_124_3477_n1418), .S(DP_OP_422J2_124_3477_n1419) );
  FADDX1_HVT DP_OP_422J2_124_3477_U866 ( .A(DP_OP_422J2_124_3477_n1481), .B(
        DP_OP_422J2_124_3477_n1459), .CI(DP_OP_422J2_124_3477_n1467), .CO(
        DP_OP_422J2_124_3477_n1416), .S(DP_OP_422J2_124_3477_n1417) );
  FADDX1_HVT DP_OP_422J2_124_3477_U865 ( .A(DP_OP_422J2_124_3477_n1469), .B(
        DP_OP_422J2_124_3477_n1493), .CI(DP_OP_422J2_124_3477_n1501), .CO(
        DP_OP_422J2_124_3477_n1414), .S(DP_OP_422J2_124_3477_n1415) );
  FADDX1_HVT DP_OP_422J2_124_3477_U864 ( .A(DP_OP_422J2_124_3477_n1465), .B(
        DP_OP_422J2_124_3477_n1491), .CI(DP_OP_422J2_124_3477_n1608), .CO(
        DP_OP_422J2_124_3477_n1412), .S(DP_OP_422J2_124_3477_n1413) );
  FADDX1_HVT DP_OP_422J2_124_3477_U863 ( .A(DP_OP_422J2_124_3477_n1606), .B(
        DP_OP_422J2_124_3477_n1604), .CI(DP_OP_422J2_124_3477_n1602), .CO(
        DP_OP_422J2_124_3477_n1410), .S(DP_OP_422J2_124_3477_n1411) );
  FADDX1_HVT DP_OP_422J2_124_3477_U862 ( .A(DP_OP_422J2_124_3477_n1594), .B(
        DP_OP_422J2_124_3477_n1600), .CI(DP_OP_422J2_124_3477_n1596), .CO(
        DP_OP_422J2_124_3477_n1408), .S(DP_OP_422J2_124_3477_n1409) );
  FADDX1_HVT DP_OP_422J2_124_3477_U861 ( .A(DP_OP_422J2_124_3477_n1598), .B(
        DP_OP_422J2_124_3477_n1592), .CI(DP_OP_422J2_124_3477_n1453), .CO(
        DP_OP_422J2_124_3477_n1406), .S(DP_OP_422J2_124_3477_n1407) );
  FADDX1_HVT DP_OP_422J2_124_3477_U860 ( .A(DP_OP_422J2_124_3477_n1455), .B(
        DP_OP_422J2_124_3477_n1590), .CI(DP_OP_422J2_124_3477_n1586), .CO(
        DP_OP_422J2_124_3477_n1404), .S(DP_OP_422J2_124_3477_n1405) );
  FADDX1_HVT DP_OP_422J2_124_3477_U859 ( .A(DP_OP_422J2_124_3477_n1457), .B(
        DP_OP_422J2_124_3477_n1588), .CI(DP_OP_422J2_124_3477_n1584), .CO(
        DP_OP_422J2_124_3477_n1402), .S(DP_OP_422J2_124_3477_n1403) );
  FADDX1_HVT DP_OP_422J2_124_3477_U858 ( .A(DP_OP_422J2_124_3477_n1574), .B(
        DP_OP_422J2_124_3477_n1437), .CI(DP_OP_422J2_124_3477_n1449), .CO(
        DP_OP_422J2_124_3477_n1400), .S(DP_OP_422J2_124_3477_n1401) );
  FADDX1_HVT DP_OP_422J2_124_3477_U857 ( .A(DP_OP_422J2_124_3477_n1582), .B(
        DP_OP_422J2_124_3477_n1451), .CI(DP_OP_422J2_124_3477_n1447), .CO(
        DP_OP_422J2_124_3477_n1398), .S(DP_OP_422J2_124_3477_n1399) );
  FADDX1_HVT DP_OP_422J2_124_3477_U856 ( .A(DP_OP_422J2_124_3477_n1580), .B(
        DP_OP_422J2_124_3477_n1439), .CI(DP_OP_422J2_124_3477_n1441), .CO(
        DP_OP_422J2_124_3477_n1396), .S(DP_OP_422J2_124_3477_n1397) );
  FADDX1_HVT DP_OP_422J2_124_3477_U855 ( .A(DP_OP_422J2_124_3477_n1578), .B(
        DP_OP_422J2_124_3477_n1445), .CI(DP_OP_422J2_124_3477_n1443), .CO(
        DP_OP_422J2_124_3477_n1394), .S(DP_OP_422J2_124_3477_n1395) );
  FADDX1_HVT DP_OP_422J2_124_3477_U854 ( .A(DP_OP_422J2_124_3477_n1576), .B(
        DP_OP_422J2_124_3477_n1572), .CI(DP_OP_422J2_124_3477_n1433), .CO(
        DP_OP_422J2_124_3477_n1392), .S(DP_OP_422J2_124_3477_n1393) );
  FADDX1_HVT DP_OP_422J2_124_3477_U853 ( .A(DP_OP_422J2_124_3477_n1435), .B(
        DP_OP_422J2_124_3477_n1431), .CI(DP_OP_422J2_124_3477_n1429), .CO(
        DP_OP_422J2_124_3477_n1390), .S(DP_OP_422J2_124_3477_n1391) );
  FADDX1_HVT DP_OP_422J2_124_3477_U852 ( .A(DP_OP_422J2_124_3477_n1570), .B(
        DP_OP_422J2_124_3477_n1421), .CI(DP_OP_422J2_124_3477_n1419), .CO(
        DP_OP_422J2_124_3477_n1388), .S(DP_OP_422J2_124_3477_n1389) );
  FADDX1_HVT DP_OP_422J2_124_3477_U851 ( .A(DP_OP_422J2_124_3477_n1425), .B(
        DP_OP_422J2_124_3477_n1415), .CI(DP_OP_422J2_124_3477_n1417), .CO(
        DP_OP_422J2_124_3477_n1386), .S(DP_OP_422J2_124_3477_n1387) );
  FADDX1_HVT DP_OP_422J2_124_3477_U850 ( .A(DP_OP_422J2_124_3477_n1423), .B(
        DP_OP_422J2_124_3477_n1427), .CI(DP_OP_422J2_124_3477_n1568), .CO(
        DP_OP_422J2_124_3477_n1384), .S(DP_OP_422J2_124_3477_n1385) );
  FADDX1_HVT DP_OP_422J2_124_3477_U849 ( .A(DP_OP_422J2_124_3477_n1566), .B(
        DP_OP_422J2_124_3477_n1413), .CI(DP_OP_422J2_124_3477_n1564), .CO(
        DP_OP_422J2_124_3477_n1382), .S(DP_OP_422J2_124_3477_n1383) );
  FADDX1_HVT DP_OP_422J2_124_3477_U848 ( .A(DP_OP_422J2_124_3477_n1562), .B(
        DP_OP_422J2_124_3477_n1409), .CI(DP_OP_422J2_124_3477_n1411), .CO(
        DP_OP_422J2_124_3477_n1380), .S(DP_OP_422J2_124_3477_n1381) );
  FADDX1_HVT DP_OP_422J2_124_3477_U847 ( .A(DP_OP_422J2_124_3477_n1560), .B(
        DP_OP_422J2_124_3477_n1556), .CI(DP_OP_422J2_124_3477_n1558), .CO(
        DP_OP_422J2_124_3477_n1378), .S(DP_OP_422J2_124_3477_n1379) );
  FADDX1_HVT DP_OP_422J2_124_3477_U846 ( .A(DP_OP_422J2_124_3477_n1407), .B(
        DP_OP_422J2_124_3477_n1554), .CI(DP_OP_422J2_124_3477_n1552), .CO(
        DP_OP_422J2_124_3477_n1376), .S(DP_OP_422J2_124_3477_n1377) );
  FADDX1_HVT DP_OP_422J2_124_3477_U845 ( .A(DP_OP_422J2_124_3477_n1405), .B(
        DP_OP_422J2_124_3477_n1403), .CI(DP_OP_422J2_124_3477_n1399), .CO(
        DP_OP_422J2_124_3477_n1374), .S(DP_OP_422J2_124_3477_n1375) );
  FADDX1_HVT DP_OP_422J2_124_3477_U844 ( .A(DP_OP_422J2_124_3477_n1401), .B(
        DP_OP_422J2_124_3477_n1397), .CI(DP_OP_422J2_124_3477_n1393), .CO(
        DP_OP_422J2_124_3477_n1372), .S(DP_OP_422J2_124_3477_n1373) );
  FADDX1_HVT DP_OP_422J2_124_3477_U843 ( .A(DP_OP_422J2_124_3477_n1550), .B(
        DP_OP_422J2_124_3477_n1395), .CI(DP_OP_422J2_124_3477_n1548), .CO(
        DP_OP_422J2_124_3477_n1370), .S(DP_OP_422J2_124_3477_n1371) );
  FADDX1_HVT DP_OP_422J2_124_3477_U842 ( .A(DP_OP_422J2_124_3477_n1391), .B(
        DP_OP_422J2_124_3477_n1389), .CI(DP_OP_422J2_124_3477_n1387), .CO(
        DP_OP_422J2_124_3477_n1368), .S(DP_OP_422J2_124_3477_n1369) );
  FADDX1_HVT DP_OP_422J2_124_3477_U841 ( .A(DP_OP_422J2_124_3477_n1546), .B(
        DP_OP_422J2_124_3477_n1385), .CI(DP_OP_422J2_124_3477_n1544), .CO(
        DP_OP_422J2_124_3477_n1366), .S(DP_OP_422J2_124_3477_n1367) );
  FADDX1_HVT DP_OP_422J2_124_3477_U840 ( .A(DP_OP_422J2_124_3477_n1383), .B(
        DP_OP_422J2_124_3477_n1542), .CI(DP_OP_422J2_124_3477_n1540), .CO(
        DP_OP_422J2_124_3477_n1364), .S(DP_OP_422J2_124_3477_n1365) );
  FADDX1_HVT DP_OP_422J2_124_3477_U839 ( .A(DP_OP_422J2_124_3477_n1379), .B(
        DP_OP_422J2_124_3477_n1381), .CI(DP_OP_422J2_124_3477_n1538), .CO(
        DP_OP_422J2_124_3477_n1362), .S(DP_OP_422J2_124_3477_n1363) );
  FADDX1_HVT DP_OP_422J2_124_3477_U838 ( .A(DP_OP_422J2_124_3477_n1377), .B(
        DP_OP_422J2_124_3477_n1375), .CI(DP_OP_422J2_124_3477_n1536), .CO(
        DP_OP_422J2_124_3477_n1360), .S(DP_OP_422J2_124_3477_n1361) );
  FADDX1_HVT DP_OP_422J2_124_3477_U837 ( .A(DP_OP_422J2_124_3477_n1371), .B(
        DP_OP_422J2_124_3477_n1373), .CI(DP_OP_422J2_124_3477_n1534), .CO(
        DP_OP_422J2_124_3477_n1358), .S(DP_OP_422J2_124_3477_n1359) );
  FADDX1_HVT DP_OP_422J2_124_3477_U836 ( .A(DP_OP_422J2_124_3477_n1369), .B(
        DP_OP_422J2_124_3477_n1367), .CI(DP_OP_422J2_124_3477_n1532), .CO(
        DP_OP_422J2_124_3477_n1356), .S(DP_OP_422J2_124_3477_n1357) );
  FADDX1_HVT DP_OP_422J2_124_3477_U835 ( .A(DP_OP_422J2_124_3477_n1365), .B(
        DP_OP_422J2_124_3477_n1530), .CI(DP_OP_422J2_124_3477_n1363), .CO(
        DP_OP_422J2_124_3477_n1354), .S(DP_OP_422J2_124_3477_n1355) );
  FADDX1_HVT DP_OP_422J2_124_3477_U834 ( .A(DP_OP_422J2_124_3477_n1361), .B(
        DP_OP_422J2_124_3477_n1528), .CI(DP_OP_422J2_124_3477_n1359), .CO(
        DP_OP_422J2_124_3477_n1352), .S(DP_OP_422J2_124_3477_n1353) );
  FADDX1_HVT DP_OP_422J2_124_3477_U833 ( .A(DP_OP_422J2_124_3477_n1357), .B(
        DP_OP_422J2_124_3477_n1526), .CI(DP_OP_422J2_124_3477_n1355), .CO(
        DP_OP_422J2_124_3477_n1350), .S(DP_OP_422J2_124_3477_n1351) );
  HADDX1_HVT DP_OP_422J2_124_3477_U832 ( .A0(DP_OP_422J2_124_3477_n2980), .B0(
        DP_OP_422J2_124_3477_n1925), .C1(DP_OP_422J2_124_3477_n1348), .SO(
        DP_OP_422J2_124_3477_n1349) );
  FADDX1_HVT DP_OP_422J2_124_3477_U831 ( .A(DP_OP_422J2_124_3477_n2453), .B(
        DP_OP_422J2_124_3477_n2365), .CI(DP_OP_422J2_124_3477_n1881), .CO(
        DP_OP_422J2_124_3477_n1346), .S(DP_OP_422J2_124_3477_n1347) );
  FADDX1_HVT DP_OP_422J2_124_3477_U830 ( .A(DP_OP_422J2_124_3477_n2497), .B(
        DP_OP_422J2_124_3477_n2277), .CI(DP_OP_422J2_124_3477_n2321), .CO(
        DP_OP_422J2_124_3477_n1344), .S(DP_OP_422J2_124_3477_n1345) );
  FADDX1_HVT DP_OP_422J2_124_3477_U829 ( .A(DP_OP_422J2_124_3477_n2805), .B(
        DP_OP_422J2_124_3477_n1969), .CI(DP_OP_422J2_124_3477_n2057), .CO(
        DP_OP_422J2_124_3477_n1342), .S(DP_OP_422J2_124_3477_n1343) );
  FADDX1_HVT DP_OP_422J2_124_3477_U828 ( .A(DP_OP_422J2_124_3477_n2541), .B(
        DP_OP_422J2_124_3477_n2101), .CI(DP_OP_422J2_124_3477_n2629), .CO(
        DP_OP_422J2_124_3477_n1340), .S(DP_OP_422J2_124_3477_n1341) );
  FADDX1_HVT DP_OP_422J2_124_3477_U827 ( .A(DP_OP_422J2_124_3477_n2013), .B(
        DP_OP_422J2_124_3477_n2849), .CI(DP_OP_422J2_124_3477_n2145), .CO(
        DP_OP_422J2_124_3477_n1338), .S(DP_OP_422J2_124_3477_n1339) );
  FADDX1_HVT DP_OP_422J2_124_3477_U826 ( .A(DP_OP_422J2_124_3477_n2409), .B(
        DP_OP_422J2_124_3477_n2893), .CI(DP_OP_422J2_124_3477_n2717), .CO(
        DP_OP_422J2_124_3477_n1336), .S(DP_OP_422J2_124_3477_n1337) );
  FADDX1_HVT DP_OP_422J2_124_3477_U825 ( .A(DP_OP_422J2_124_3477_n2233), .B(
        DP_OP_422J2_124_3477_n2189), .CI(DP_OP_422J2_124_3477_n2673), .CO(
        DP_OP_422J2_124_3477_n1334), .S(DP_OP_422J2_124_3477_n1335) );
  FADDX1_HVT DP_OP_422J2_124_3477_U824 ( .A(DP_OP_422J2_124_3477_n2937), .B(
        DP_OP_422J2_124_3477_n2585), .CI(DP_OP_422J2_124_3477_n2761), .CO(
        DP_OP_422J2_124_3477_n1332), .S(DP_OP_422J2_124_3477_n1333) );
  FADDX1_HVT DP_OP_422J2_124_3477_U823 ( .A(DP_OP_422J2_124_3477_n2379), .B(
        DP_OP_422J2_124_3477_n3000), .CI(DP_OP_422J2_124_3477_n1932), .CO(
        DP_OP_422J2_124_3477_n1330), .S(DP_OP_422J2_124_3477_n1331) );
  FADDX1_HVT DP_OP_422J2_124_3477_U822 ( .A(DP_OP_422J2_124_3477_n2372), .B(
        DP_OP_422J2_124_3477_n1939), .CI(DP_OP_422J2_124_3477_n1946), .CO(
        DP_OP_422J2_124_3477_n1328), .S(DP_OP_422J2_124_3477_n1329) );
  FADDX1_HVT DP_OP_422J2_124_3477_U821 ( .A(DP_OP_422J2_124_3477_n2386), .B(
        DP_OP_422J2_124_3477_n1976), .CI(DP_OP_422J2_124_3477_n2993), .CO(
        DP_OP_422J2_124_3477_n1326), .S(DP_OP_422J2_124_3477_n1327) );
  FADDX1_HVT DP_OP_422J2_124_3477_U820 ( .A(DP_OP_422J2_124_3477_n2342), .B(
        DP_OP_422J2_124_3477_n2986), .CI(DP_OP_422J2_124_3477_n2958), .CO(
        DP_OP_422J2_124_3477_n1324), .S(DP_OP_422J2_124_3477_n1325) );
  FADDX1_HVT DP_OP_422J2_124_3477_U819 ( .A(DP_OP_422J2_124_3477_n2335), .B(
        DP_OP_422J2_124_3477_n2951), .CI(DP_OP_422J2_124_3477_n2944), .CO(
        DP_OP_422J2_124_3477_n1322), .S(DP_OP_422J2_124_3477_n1323) );
  FADDX1_HVT DP_OP_422J2_124_3477_U818 ( .A(DP_OP_422J2_124_3477_n2298), .B(
        DP_OP_422J2_124_3477_n2914), .CI(DP_OP_422J2_124_3477_n2907), .CO(
        DP_OP_422J2_124_3477_n1320), .S(DP_OP_422J2_124_3477_n1321) );
  FADDX1_HVT DP_OP_422J2_124_3477_U817 ( .A(DP_OP_422J2_124_3477_n2291), .B(
        DP_OP_422J2_124_3477_n1983), .CI(DP_OP_422J2_124_3477_n2900), .CO(
        DP_OP_422J2_124_3477_n1318), .S(DP_OP_422J2_124_3477_n1319) );
  FADDX1_HVT DP_OP_422J2_124_3477_U816 ( .A(DP_OP_422J2_124_3477_n2284), .B(
        DP_OP_422J2_124_3477_n2870), .CI(DP_OP_422J2_124_3477_n2863), .CO(
        DP_OP_422J2_124_3477_n1316), .S(DP_OP_422J2_124_3477_n1317) );
  FADDX1_HVT DP_OP_422J2_124_3477_U815 ( .A(DP_OP_422J2_124_3477_n2254), .B(
        DP_OP_422J2_124_3477_n2856), .CI(DP_OP_422J2_124_3477_n1990), .CO(
        DP_OP_422J2_124_3477_n1314), .S(DP_OP_422J2_124_3477_n1315) );
  FADDX1_HVT DP_OP_422J2_124_3477_U814 ( .A(DP_OP_422J2_124_3477_n2247), .B(
        DP_OP_422J2_124_3477_n2020), .CI(DP_OP_422J2_124_3477_n2027), .CO(
        DP_OP_422J2_124_3477_n1312), .S(DP_OP_422J2_124_3477_n1313) );
  FADDX1_HVT DP_OP_422J2_124_3477_U813 ( .A(DP_OP_422J2_124_3477_n2328), .B(
        DP_OP_422J2_124_3477_n2034), .CI(DP_OP_422J2_124_3477_n2826), .CO(
        DP_OP_422J2_124_3477_n1310), .S(DP_OP_422J2_124_3477_n1311) );
  FADDX1_HVT DP_OP_422J2_124_3477_U812 ( .A(DP_OP_422J2_124_3477_n2416), .B(
        DP_OP_422J2_124_3477_n2819), .CI(DP_OP_422J2_124_3477_n2064), .CO(
        DP_OP_422J2_124_3477_n1308), .S(DP_OP_422J2_124_3477_n1309) );
  FADDX1_HVT DP_OP_422J2_124_3477_U811 ( .A(DP_OP_422J2_124_3477_n2812), .B(
        DP_OP_422J2_124_3477_n2071), .CI(DP_OP_422J2_124_3477_n2078), .CO(
        DP_OP_422J2_124_3477_n1306), .S(DP_OP_422J2_124_3477_n1307) );
  FADDX1_HVT DP_OP_422J2_124_3477_U810 ( .A(DP_OP_422J2_124_3477_n2782), .B(
        DP_OP_422J2_124_3477_n2108), .CI(DP_OP_422J2_124_3477_n2115), .CO(
        DP_OP_422J2_124_3477_n1304), .S(DP_OP_422J2_124_3477_n1305) );
  FADDX1_HVT DP_OP_422J2_124_3477_U809 ( .A(DP_OP_422J2_124_3477_n2775), .B(
        DP_OP_422J2_124_3477_n2122), .CI(DP_OP_422J2_124_3477_n2152), .CO(
        DP_OP_422J2_124_3477_n1302), .S(DP_OP_422J2_124_3477_n1303) );
  FADDX1_HVT DP_OP_422J2_124_3477_U808 ( .A(DP_OP_422J2_124_3477_n2768), .B(
        DP_OP_422J2_124_3477_n2159), .CI(DP_OP_422J2_124_3477_n2166), .CO(
        DP_OP_422J2_124_3477_n1300), .S(DP_OP_422J2_124_3477_n1301) );
  FADDX1_HVT DP_OP_422J2_124_3477_U807 ( .A(DP_OP_422J2_124_3477_n2738), .B(
        DP_OP_422J2_124_3477_n2196), .CI(DP_OP_422J2_124_3477_n2203), .CO(
        DP_OP_422J2_124_3477_n1298), .S(DP_OP_422J2_124_3477_n1299) );
  FADDX1_HVT DP_OP_422J2_124_3477_U806 ( .A(DP_OP_422J2_124_3477_n2731), .B(
        DP_OP_422J2_124_3477_n2210), .CI(DP_OP_422J2_124_3477_n2240), .CO(
        DP_OP_422J2_124_3477_n1296), .S(DP_OP_422J2_124_3477_n1297) );
  FADDX1_HVT DP_OP_422J2_124_3477_U805 ( .A(DP_OP_422J2_124_3477_n2724), .B(
        DP_OP_422J2_124_3477_n2423), .CI(DP_OP_422J2_124_3477_n2430), .CO(
        DP_OP_422J2_124_3477_n1294), .S(DP_OP_422J2_124_3477_n1295) );
  FADDX1_HVT DP_OP_422J2_124_3477_U804 ( .A(DP_OP_422J2_124_3477_n2694), .B(
        DP_OP_422J2_124_3477_n2460), .CI(DP_OP_422J2_124_3477_n2467), .CO(
        DP_OP_422J2_124_3477_n1292), .S(DP_OP_422J2_124_3477_n1293) );
  FADDX1_HVT DP_OP_422J2_124_3477_U803 ( .A(DP_OP_422J2_124_3477_n2687), .B(
        DP_OP_422J2_124_3477_n2474), .CI(DP_OP_422J2_124_3477_n2504), .CO(
        DP_OP_422J2_124_3477_n1290), .S(DP_OP_422J2_124_3477_n1291) );
  FADDX1_HVT DP_OP_422J2_124_3477_U802 ( .A(DP_OP_422J2_124_3477_n2680), .B(
        DP_OP_422J2_124_3477_n2511), .CI(DP_OP_422J2_124_3477_n2518), .CO(
        DP_OP_422J2_124_3477_n1288), .S(DP_OP_422J2_124_3477_n1289) );
  FADDX1_HVT DP_OP_422J2_124_3477_U801 ( .A(DP_OP_422J2_124_3477_n2650), .B(
        DP_OP_422J2_124_3477_n2643), .CI(DP_OP_422J2_124_3477_n2636), .CO(
        DP_OP_422J2_124_3477_n1286), .S(DP_OP_422J2_124_3477_n1287) );
  FADDX1_HVT DP_OP_422J2_124_3477_U800 ( .A(DP_OP_422J2_124_3477_n2592), .B(
        DP_OP_422J2_124_3477_n2606), .CI(DP_OP_422J2_124_3477_n2548), .CO(
        DP_OP_422J2_124_3477_n1284), .S(DP_OP_422J2_124_3477_n1285) );
  FADDX1_HVT DP_OP_422J2_124_3477_U799 ( .A(DP_OP_422J2_124_3477_n2555), .B(
        DP_OP_422J2_124_3477_n2562), .CI(DP_OP_422J2_124_3477_n2599), .CO(
        DP_OP_422J2_124_3477_n1282), .S(DP_OP_422J2_124_3477_n1283) );
  FADDX1_HVT DP_OP_422J2_124_3477_U798 ( .A(DP_OP_422J2_124_3477_n1349), .B(
        DP_OP_422J2_124_3477_n1524), .CI(DP_OP_422J2_124_3477_n1514), .CO(
        DP_OP_422J2_124_3477_n1280), .S(DP_OP_422J2_124_3477_n1281) );
  FADDX1_HVT DP_OP_422J2_124_3477_U797 ( .A(DP_OP_422J2_124_3477_n1522), .B(
        DP_OP_422J2_124_3477_n1520), .CI(DP_OP_422J2_124_3477_n1518), .CO(
        DP_OP_422J2_124_3477_n1278), .S(DP_OP_422J2_124_3477_n1279) );
  FADDX1_HVT DP_OP_422J2_124_3477_U796 ( .A(DP_OP_422J2_124_3477_n1516), .B(
        DP_OP_422J2_124_3477_n1512), .CI(DP_OP_422J2_124_3477_n1508), .CO(
        DP_OP_422J2_124_3477_n1276), .S(DP_OP_422J2_124_3477_n1277) );
  FADDX1_HVT DP_OP_422J2_124_3477_U795 ( .A(DP_OP_422J2_124_3477_n1510), .B(
        DP_OP_422J2_124_3477_n1484), .CI(DP_OP_422J2_124_3477_n1482), .CO(
        DP_OP_422J2_124_3477_n1274), .S(DP_OP_422J2_124_3477_n1275) );
  FADDX1_HVT DP_OP_422J2_124_3477_U794 ( .A(DP_OP_422J2_124_3477_n1486), .B(
        DP_OP_422J2_124_3477_n1458), .CI(DP_OP_422J2_124_3477_n1506), .CO(
        DP_OP_422J2_124_3477_n1272), .S(DP_OP_422J2_124_3477_n1273) );
  FADDX1_HVT DP_OP_422J2_124_3477_U793 ( .A(DP_OP_422J2_124_3477_n1478), .B(
        DP_OP_422J2_124_3477_n1504), .CI(DP_OP_422J2_124_3477_n1502), .CO(
        DP_OP_422J2_124_3477_n1270), .S(DP_OP_422J2_124_3477_n1271) );
  FADDX1_HVT DP_OP_422J2_124_3477_U792 ( .A(DP_OP_422J2_124_3477_n1474), .B(
        DP_OP_422J2_124_3477_n1500), .CI(DP_OP_422J2_124_3477_n1498), .CO(
        DP_OP_422J2_124_3477_n1268), .S(DP_OP_422J2_124_3477_n1269) );
  FADDX1_HVT DP_OP_422J2_124_3477_U791 ( .A(DP_OP_422J2_124_3477_n1468), .B(
        DP_OP_422J2_124_3477_n1460), .CI(DP_OP_422J2_124_3477_n1462), .CO(
        DP_OP_422J2_124_3477_n1266), .S(DP_OP_422J2_124_3477_n1267) );
  FADDX1_HVT DP_OP_422J2_124_3477_U790 ( .A(DP_OP_422J2_124_3477_n1466), .B(
        DP_OP_422J2_124_3477_n1496), .CI(DP_OP_422J2_124_3477_n1494), .CO(
        DP_OP_422J2_124_3477_n1264), .S(DP_OP_422J2_124_3477_n1265) );
  FADDX1_HVT DP_OP_422J2_124_3477_U789 ( .A(DP_OP_422J2_124_3477_n1476), .B(
        DP_OP_422J2_124_3477_n1492), .CI(DP_OP_422J2_124_3477_n1464), .CO(
        DP_OP_422J2_124_3477_n1262), .S(DP_OP_422J2_124_3477_n1263) );
  FADDX1_HVT DP_OP_422J2_124_3477_U788 ( .A(DP_OP_422J2_124_3477_n1472), .B(
        DP_OP_422J2_124_3477_n1490), .CI(DP_OP_422J2_124_3477_n1488), .CO(
        DP_OP_422J2_124_3477_n1260), .S(DP_OP_422J2_124_3477_n1261) );
  FADDX1_HVT DP_OP_422J2_124_3477_U787 ( .A(DP_OP_422J2_124_3477_n1470), .B(
        DP_OP_422J2_124_3477_n1480), .CI(DP_OP_422J2_124_3477_n1339), .CO(
        DP_OP_422J2_124_3477_n1258), .S(DP_OP_422J2_124_3477_n1259) );
  FADDX1_HVT DP_OP_422J2_124_3477_U786 ( .A(DP_OP_422J2_124_3477_n1341), .B(
        DP_OP_422J2_124_3477_n1333), .CI(DP_OP_422J2_124_3477_n1335), .CO(
        DP_OP_422J2_124_3477_n1256), .S(DP_OP_422J2_124_3477_n1257) );
  FADDX1_HVT DP_OP_422J2_124_3477_U785 ( .A(DP_OP_422J2_124_3477_n1345), .B(
        DP_OP_422J2_124_3477_n1343), .CI(DP_OP_422J2_124_3477_n1347), .CO(
        DP_OP_422J2_124_3477_n1254), .S(DP_OP_422J2_124_3477_n1255) );
  FADDX1_HVT DP_OP_422J2_124_3477_U784 ( .A(DP_OP_422J2_124_3477_n1337), .B(
        DP_OP_422J2_124_3477_n1289), .CI(DP_OP_422J2_124_3477_n1287), .CO(
        DP_OP_422J2_124_3477_n1252), .S(DP_OP_422J2_124_3477_n1253) );
  FADDX1_HVT DP_OP_422J2_124_3477_U783 ( .A(DP_OP_422J2_124_3477_n1283), .B(
        DP_OP_422J2_124_3477_n1331), .CI(DP_OP_422J2_124_3477_n1329), .CO(
        DP_OP_422J2_124_3477_n1250), .S(DP_OP_422J2_124_3477_n1251) );
  FADDX1_HVT DP_OP_422J2_124_3477_U782 ( .A(DP_OP_422J2_124_3477_n1319), .B(
        DP_OP_422J2_124_3477_n1309), .CI(DP_OP_422J2_124_3477_n1315), .CO(
        DP_OP_422J2_124_3477_n1248), .S(DP_OP_422J2_124_3477_n1249) );
  FADDX1_HVT DP_OP_422J2_124_3477_U781 ( .A(DP_OP_422J2_124_3477_n1313), .B(
        DP_OP_422J2_124_3477_n1311), .CI(DP_OP_422J2_124_3477_n1295), .CO(
        DP_OP_422J2_124_3477_n1246), .S(DP_OP_422J2_124_3477_n1247) );
  FADDX1_HVT DP_OP_422J2_124_3477_U780 ( .A(DP_OP_422J2_124_3477_n1317), .B(
        DP_OP_422J2_124_3477_n1291), .CI(DP_OP_422J2_124_3477_n1285), .CO(
        DP_OP_422J2_124_3477_n1244), .S(DP_OP_422J2_124_3477_n1245) );
  FADDX1_HVT DP_OP_422J2_124_3477_U779 ( .A(DP_OP_422J2_124_3477_n1321), .B(
        DP_OP_422J2_124_3477_n1303), .CI(DP_OP_422J2_124_3477_n1305), .CO(
        DP_OP_422J2_124_3477_n1242), .S(DP_OP_422J2_124_3477_n1243) );
  FADDX1_HVT DP_OP_422J2_124_3477_U778 ( .A(DP_OP_422J2_124_3477_n1301), .B(
        DP_OP_422J2_124_3477_n1299), .CI(DP_OP_422J2_124_3477_n1293), .CO(
        DP_OP_422J2_124_3477_n1240), .S(DP_OP_422J2_124_3477_n1241) );
  FADDX1_HVT DP_OP_422J2_124_3477_U777 ( .A(DP_OP_422J2_124_3477_n1297), .B(
        DP_OP_422J2_124_3477_n1327), .CI(DP_OP_422J2_124_3477_n1323), .CO(
        DP_OP_422J2_124_3477_n1238), .S(DP_OP_422J2_124_3477_n1239) );
  FADDX1_HVT DP_OP_422J2_124_3477_U776 ( .A(DP_OP_422J2_124_3477_n1325), .B(
        DP_OP_422J2_124_3477_n1307), .CI(DP_OP_422J2_124_3477_n1456), .CO(
        DP_OP_422J2_124_3477_n1236), .S(DP_OP_422J2_124_3477_n1237) );
  FADDX1_HVT DP_OP_422J2_124_3477_U775 ( .A(DP_OP_422J2_124_3477_n1454), .B(
        DP_OP_422J2_124_3477_n1452), .CI(DP_OP_422J2_124_3477_n1450), .CO(
        DP_OP_422J2_124_3477_n1234), .S(DP_OP_422J2_124_3477_n1235) );
  FADDX1_HVT DP_OP_422J2_124_3477_U774 ( .A(DP_OP_422J2_124_3477_n1448), .B(
        DP_OP_422J2_124_3477_n1436), .CI(DP_OP_422J2_124_3477_n1438), .CO(
        DP_OP_422J2_124_3477_n1232), .S(DP_OP_422J2_124_3477_n1233) );
  FADDX1_HVT DP_OP_422J2_124_3477_U773 ( .A(DP_OP_422J2_124_3477_n1442), .B(
        DP_OP_422J2_124_3477_n1446), .CI(DP_OP_422J2_124_3477_n1440), .CO(
        DP_OP_422J2_124_3477_n1230), .S(DP_OP_422J2_124_3477_n1231) );
  FADDX1_HVT DP_OP_422J2_124_3477_U772 ( .A(DP_OP_422J2_124_3477_n1444), .B(
        DP_OP_422J2_124_3477_n1281), .CI(DP_OP_422J2_124_3477_n1434), .CO(
        DP_OP_422J2_124_3477_n1228), .S(DP_OP_422J2_124_3477_n1229) );
  FADDX1_HVT DP_OP_422J2_124_3477_U771 ( .A(DP_OP_422J2_124_3477_n1279), .B(
        DP_OP_422J2_124_3477_n1277), .CI(DP_OP_422J2_124_3477_n1275), .CO(
        DP_OP_422J2_124_3477_n1226), .S(DP_OP_422J2_124_3477_n1227) );
  FADDX1_HVT DP_OP_422J2_124_3477_U770 ( .A(DP_OP_422J2_124_3477_n1432), .B(
        DP_OP_422J2_124_3477_n1430), .CI(DP_OP_422J2_124_3477_n1428), .CO(
        DP_OP_422J2_124_3477_n1224), .S(DP_OP_422J2_124_3477_n1225) );
  FADDX1_HVT DP_OP_422J2_124_3477_U769 ( .A(DP_OP_422J2_124_3477_n1416), .B(
        DP_OP_422J2_124_3477_n1261), .CI(DP_OP_422J2_124_3477_n1259), .CO(
        DP_OP_422J2_124_3477_n1222), .S(DP_OP_422J2_124_3477_n1223) );
  FADDX1_HVT DP_OP_422J2_124_3477_U768 ( .A(DP_OP_422J2_124_3477_n1426), .B(
        DP_OP_422J2_124_3477_n1271), .CI(DP_OP_422J2_124_3477_n1273), .CO(
        DP_OP_422J2_124_3477_n1220), .S(DP_OP_422J2_124_3477_n1221) );
  FADDX1_HVT DP_OP_422J2_124_3477_U767 ( .A(DP_OP_422J2_124_3477_n1424), .B(
        DP_OP_422J2_124_3477_n1267), .CI(DP_OP_422J2_124_3477_n1263), .CO(
        DP_OP_422J2_124_3477_n1218), .S(DP_OP_422J2_124_3477_n1219) );
  FADDX1_HVT DP_OP_422J2_124_3477_U766 ( .A(DP_OP_422J2_124_3477_n1422), .B(
        DP_OP_422J2_124_3477_n1269), .CI(DP_OP_422J2_124_3477_n1265), .CO(
        DP_OP_422J2_124_3477_n1216), .S(DP_OP_422J2_124_3477_n1217) );
  FADDX1_HVT DP_OP_422J2_124_3477_U765 ( .A(DP_OP_422J2_124_3477_n1420), .B(
        DP_OP_422J2_124_3477_n1414), .CI(DP_OP_422J2_124_3477_n1418), .CO(
        DP_OP_422J2_124_3477_n1214), .S(DP_OP_422J2_124_3477_n1215) );
  FADDX1_HVT DP_OP_422J2_124_3477_U764 ( .A(DP_OP_422J2_124_3477_n1255), .B(
        DP_OP_422J2_124_3477_n1257), .CI(DP_OP_422J2_124_3477_n1253), .CO(
        DP_OP_422J2_124_3477_n1212), .S(DP_OP_422J2_124_3477_n1213) );
  FADDX1_HVT DP_OP_422J2_124_3477_U763 ( .A(DP_OP_422J2_124_3477_n1245), .B(
        DP_OP_422J2_124_3477_n1247), .CI(DP_OP_422J2_124_3477_n1412), .CO(
        DP_OP_422J2_124_3477_n1210), .S(DP_OP_422J2_124_3477_n1211) );
  FADDX1_HVT DP_OP_422J2_124_3477_U762 ( .A(DP_OP_422J2_124_3477_n1243), .B(
        DP_OP_422J2_124_3477_n1251), .CI(DP_OP_422J2_124_3477_n1249), .CO(
        DP_OP_422J2_124_3477_n1208), .S(DP_OP_422J2_124_3477_n1209) );
  FADDX1_HVT DP_OP_422J2_124_3477_U761 ( .A(DP_OP_422J2_124_3477_n1239), .B(
        DP_OP_422J2_124_3477_n1241), .CI(DP_OP_422J2_124_3477_n1408), .CO(
        DP_OP_422J2_124_3477_n1206), .S(DP_OP_422J2_124_3477_n1207) );
  FADDX1_HVT DP_OP_422J2_124_3477_U760 ( .A(DP_OP_422J2_124_3477_n1410), .B(
        DP_OP_422J2_124_3477_n1237), .CI(DP_OP_422J2_124_3477_n1406), .CO(
        DP_OP_422J2_124_3477_n1204), .S(DP_OP_422J2_124_3477_n1205) );
  FADDX1_HVT DP_OP_422J2_124_3477_U759 ( .A(DP_OP_422J2_124_3477_n1404), .B(
        DP_OP_422J2_124_3477_n1402), .CI(DP_OP_422J2_124_3477_n1235), .CO(
        DP_OP_422J2_124_3477_n1202), .S(DP_OP_422J2_124_3477_n1203) );
  FADDX1_HVT DP_OP_422J2_124_3477_U758 ( .A(DP_OP_422J2_124_3477_n1400), .B(
        DP_OP_422J2_124_3477_n1392), .CI(DP_OP_422J2_124_3477_n1229), .CO(
        DP_OP_422J2_124_3477_n1200), .S(DP_OP_422J2_124_3477_n1201) );
  FADDX1_HVT DP_OP_422J2_124_3477_U757 ( .A(DP_OP_422J2_124_3477_n1398), .B(
        DP_OP_422J2_124_3477_n1231), .CI(DP_OP_422J2_124_3477_n1233), .CO(
        DP_OP_422J2_124_3477_n1198), .S(DP_OP_422J2_124_3477_n1199) );
  FADDX1_HVT DP_OP_422J2_124_3477_U756 ( .A(DP_OP_422J2_124_3477_n1396), .B(
        DP_OP_422J2_124_3477_n1394), .CI(DP_OP_422J2_124_3477_n1390), .CO(
        DP_OP_422J2_124_3477_n1196), .S(DP_OP_422J2_124_3477_n1197) );
  FADDX1_HVT DP_OP_422J2_124_3477_U755 ( .A(DP_OP_422J2_124_3477_n1225), .B(
        DP_OP_422J2_124_3477_n1227), .CI(DP_OP_422J2_124_3477_n1388), .CO(
        DP_OP_422J2_124_3477_n1194), .S(DP_OP_422J2_124_3477_n1195) );
  FADDX1_HVT DP_OP_422J2_124_3477_U754 ( .A(DP_OP_422J2_124_3477_n1386), .B(
        DP_OP_422J2_124_3477_n1219), .CI(DP_OP_422J2_124_3477_n1384), .CO(
        DP_OP_422J2_124_3477_n1192), .S(DP_OP_422J2_124_3477_n1193) );
  FADDX1_HVT DP_OP_422J2_124_3477_U753 ( .A(DP_OP_422J2_124_3477_n1217), .B(
        DP_OP_422J2_124_3477_n1223), .CI(DP_OP_422J2_124_3477_n1221), .CO(
        DP_OP_422J2_124_3477_n1190), .S(DP_OP_422J2_124_3477_n1191) );
  FADDX1_HVT DP_OP_422J2_124_3477_U752 ( .A(DP_OP_422J2_124_3477_n1215), .B(
        DP_OP_422J2_124_3477_n1213), .CI(DP_OP_422J2_124_3477_n1209), .CO(
        DP_OP_422J2_124_3477_n1188), .S(DP_OP_422J2_124_3477_n1189) );
  FADDX1_HVT DP_OP_422J2_124_3477_U751 ( .A(DP_OP_422J2_124_3477_n1211), .B(
        DP_OP_422J2_124_3477_n1382), .CI(DP_OP_422J2_124_3477_n1207), .CO(
        DP_OP_422J2_124_3477_n1186), .S(DP_OP_422J2_124_3477_n1187) );
  FADDX1_HVT DP_OP_422J2_124_3477_U750 ( .A(DP_OP_422J2_124_3477_n1380), .B(
        DP_OP_422J2_124_3477_n1378), .CI(DP_OP_422J2_124_3477_n1205), .CO(
        DP_OP_422J2_124_3477_n1184), .S(DP_OP_422J2_124_3477_n1185) );
  FADDX1_HVT DP_OP_422J2_124_3477_U749 ( .A(DP_OP_422J2_124_3477_n1376), .B(
        DP_OP_422J2_124_3477_n1374), .CI(DP_OP_422J2_124_3477_n1203), .CO(
        DP_OP_422J2_124_3477_n1182), .S(DP_OP_422J2_124_3477_n1183) );
  FADDX1_HVT DP_OP_422J2_124_3477_U748 ( .A(DP_OP_422J2_124_3477_n1372), .B(
        DP_OP_422J2_124_3477_n1199), .CI(DP_OP_422J2_124_3477_n1197), .CO(
        DP_OP_422J2_124_3477_n1180), .S(DP_OP_422J2_124_3477_n1181) );
  FADDX1_HVT DP_OP_422J2_124_3477_U747 ( .A(DP_OP_422J2_124_3477_n1370), .B(
        DP_OP_422J2_124_3477_n1201), .CI(DP_OP_422J2_124_3477_n1195), .CO(
        DP_OP_422J2_124_3477_n1178), .S(DP_OP_422J2_124_3477_n1179) );
  FADDX1_HVT DP_OP_422J2_124_3477_U746 ( .A(DP_OP_422J2_124_3477_n1368), .B(
        DP_OP_422J2_124_3477_n1191), .CI(DP_OP_422J2_124_3477_n1366), .CO(
        DP_OP_422J2_124_3477_n1176), .S(DP_OP_422J2_124_3477_n1177) );
  FADDX1_HVT DP_OP_422J2_124_3477_U745 ( .A(DP_OP_422J2_124_3477_n1193), .B(
        DP_OP_422J2_124_3477_n1189), .CI(DP_OP_422J2_124_3477_n1187), .CO(
        DP_OP_422J2_124_3477_n1174), .S(DP_OP_422J2_124_3477_n1175) );
  FADDX1_HVT DP_OP_422J2_124_3477_U744 ( .A(DP_OP_422J2_124_3477_n1364), .B(
        DP_OP_422J2_124_3477_n1362), .CI(DP_OP_422J2_124_3477_n1185), .CO(
        DP_OP_422J2_124_3477_n1172), .S(DP_OP_422J2_124_3477_n1173) );
  FADDX1_HVT DP_OP_422J2_124_3477_U743 ( .A(DP_OP_422J2_124_3477_n1360), .B(
        DP_OP_422J2_124_3477_n1183), .CI(DP_OP_422J2_124_3477_n1181), .CO(
        DP_OP_422J2_124_3477_n1170), .S(DP_OP_422J2_124_3477_n1171) );
  FADDX1_HVT DP_OP_422J2_124_3477_U742 ( .A(DP_OP_422J2_124_3477_n1179), .B(
        DP_OP_422J2_124_3477_n1358), .CI(DP_OP_422J2_124_3477_n1177), .CO(
        DP_OP_422J2_124_3477_n1168), .S(DP_OP_422J2_124_3477_n1169) );
  FADDX1_HVT DP_OP_422J2_124_3477_U741 ( .A(DP_OP_422J2_124_3477_n1356), .B(
        DP_OP_422J2_124_3477_n1175), .CI(DP_OP_422J2_124_3477_n1354), .CO(
        DP_OP_422J2_124_3477_n1166), .S(DP_OP_422J2_124_3477_n1167) );
  FADDX1_HVT DP_OP_422J2_124_3477_U740 ( .A(DP_OP_422J2_124_3477_n1173), .B(
        DP_OP_422J2_124_3477_n1171), .CI(DP_OP_422J2_124_3477_n1352), .CO(
        DP_OP_422J2_124_3477_n1164), .S(DP_OP_422J2_124_3477_n1165) );
  FADDX1_HVT DP_OP_422J2_124_3477_U739 ( .A(DP_OP_422J2_124_3477_n1169), .B(
        DP_OP_422J2_124_3477_n1350), .CI(DP_OP_422J2_124_3477_n1167), .CO(
        DP_OP_422J2_124_3477_n1162), .S(DP_OP_422J2_124_3477_n1163) );
  OR2X1_HVT DP_OP_422J2_124_3477_U738 ( .A1(DP_OP_422J2_124_3477_n2979), .A2(
        DP_OP_422J2_124_3477_n2452), .Y(DP_OP_422J2_124_3477_n1160) );
  FADDX1_HVT DP_OP_422J2_124_3477_U736 ( .A(DP_OP_422J2_124_3477_n2144), .B(
        DP_OP_422J2_124_3477_n1924), .CI(DP_OP_422J2_124_3477_n1880), .CO(
        DP_OP_422J2_124_3477_n1158), .S(DP_OP_422J2_124_3477_n1159) );
  FADDX1_HVT DP_OP_422J2_124_3477_U735 ( .A(DP_OP_422J2_124_3477_n2584), .B(
        DP_OP_422J2_124_3477_n2012), .CI(DP_OP_422J2_124_3477_n2364), .CO(
        DP_OP_422J2_124_3477_n1156), .S(DP_OP_422J2_124_3477_n1157) );
  FADDX1_HVT DP_OP_422J2_124_3477_U734 ( .A(DP_OP_422J2_124_3477_n2804), .B(
        DP_OP_422J2_124_3477_n2628), .CI(DP_OP_422J2_124_3477_n2188), .CO(
        DP_OP_422J2_124_3477_n1154), .S(DP_OP_422J2_124_3477_n1155) );
  FADDX1_HVT DP_OP_422J2_124_3477_U733 ( .A(DP_OP_422J2_124_3477_n2276), .B(
        DP_OP_422J2_124_3477_n2100), .CI(DP_OP_422J2_124_3477_n2848), .CO(
        DP_OP_422J2_124_3477_n1152), .S(DP_OP_422J2_124_3477_n1153) );
  FADDX1_HVT DP_OP_422J2_124_3477_U732 ( .A(DP_OP_422J2_124_3477_n2408), .B(
        DP_OP_422J2_124_3477_n2892), .CI(DP_OP_422J2_124_3477_n2672), .CO(
        DP_OP_422J2_124_3477_n1150), .S(DP_OP_422J2_124_3477_n1151) );
  FADDX1_HVT DP_OP_422J2_124_3477_U731 ( .A(DP_OP_422J2_124_3477_n2496), .B(
        DP_OP_422J2_124_3477_n2716), .CI(DP_OP_422J2_124_3477_n2540), .CO(
        DP_OP_422J2_124_3477_n1148), .S(DP_OP_422J2_124_3477_n1149) );
  FADDX1_HVT DP_OP_422J2_124_3477_U730 ( .A(DP_OP_422J2_124_3477_n2232), .B(
        DP_OP_422J2_124_3477_n2056), .CI(DP_OP_422J2_124_3477_n2936), .CO(
        DP_OP_422J2_124_3477_n1146), .S(DP_OP_422J2_124_3477_n1147) );
  FADDX1_HVT DP_OP_422J2_124_3477_U729 ( .A(DP_OP_422J2_124_3477_n2760), .B(
        DP_OP_422J2_124_3477_n1968), .CI(DP_OP_422J2_124_3477_n2320), .CO(
        DP_OP_422J2_124_3477_n1144), .S(DP_OP_422J2_124_3477_n1145) );
  FADDX1_HVT DP_OP_422J2_124_3477_U728 ( .A(DP_OP_422J2_124_3477_n2371), .B(
        DP_OP_422J2_124_3477_n2999), .CI(DP_OP_422J2_124_3477_n1931), .CO(
        DP_OP_422J2_124_3477_n1142), .S(DP_OP_422J2_124_3477_n1143) );
  FADDX1_HVT DP_OP_422J2_124_3477_U727 ( .A(DP_OP_422J2_124_3477_n2378), .B(
        DP_OP_422J2_124_3477_n2992), .CI(DP_OP_422J2_124_3477_n2985), .CO(
        DP_OP_422J2_124_3477_n1140), .S(DP_OP_422J2_124_3477_n1141) );
  FADDX1_HVT DP_OP_422J2_124_3477_U726 ( .A(DP_OP_422J2_124_3477_n2334), .B(
        DP_OP_422J2_124_3477_n2957), .CI(DP_OP_422J2_124_3477_n2950), .CO(
        DP_OP_422J2_124_3477_n1138), .S(DP_OP_422J2_124_3477_n1139) );
  FADDX1_HVT DP_OP_422J2_124_3477_U725 ( .A(DP_OP_422J2_124_3477_n2297), .B(
        DP_OP_422J2_124_3477_n2943), .CI(DP_OP_422J2_124_3477_n2913), .CO(
        DP_OP_422J2_124_3477_n1136), .S(DP_OP_422J2_124_3477_n1137) );
  FADDX1_HVT DP_OP_422J2_124_3477_U724 ( .A(DP_OP_422J2_124_3477_n2290), .B(
        DP_OP_422J2_124_3477_n1938), .CI(DP_OP_422J2_124_3477_n2906), .CO(
        DP_OP_422J2_124_3477_n1134), .S(DP_OP_422J2_124_3477_n1135) );
  FADDX1_HVT DP_OP_422J2_124_3477_U723 ( .A(DP_OP_422J2_124_3477_n2327), .B(
        DP_OP_422J2_124_3477_n2899), .CI(DP_OP_422J2_124_3477_n1945), .CO(
        DP_OP_422J2_124_3477_n1132), .S(DP_OP_422J2_124_3477_n1133) );
  FADDX1_HVT DP_OP_422J2_124_3477_U722 ( .A(DP_OP_422J2_124_3477_n2283), .B(
        DP_OP_422J2_124_3477_n2869), .CI(DP_OP_422J2_124_3477_n1975), .CO(
        DP_OP_422J2_124_3477_n1130), .S(DP_OP_422J2_124_3477_n1131) );
  FADDX1_HVT DP_OP_422J2_124_3477_U721 ( .A(DP_OP_422J2_124_3477_n2253), .B(
        DP_OP_422J2_124_3477_n2862), .CI(DP_OP_422J2_124_3477_n2855), .CO(
        DP_OP_422J2_124_3477_n1128), .S(DP_OP_422J2_124_3477_n1129) );
  FADDX1_HVT DP_OP_422J2_124_3477_U720 ( .A(DP_OP_422J2_124_3477_n2246), .B(
        DP_OP_422J2_124_3477_n1982), .CI(DP_OP_422J2_124_3477_n2825), .CO(
        DP_OP_422J2_124_3477_n1126), .S(DP_OP_422J2_124_3477_n1127) );
  FADDX1_HVT DP_OP_422J2_124_3477_U719 ( .A(DP_OP_422J2_124_3477_n2239), .B(
        DP_OP_422J2_124_3477_n1989), .CI(DP_OP_422J2_124_3477_n2818), .CO(
        DP_OP_422J2_124_3477_n1124), .S(DP_OP_422J2_124_3477_n1125) );
  FADDX1_HVT DP_OP_422J2_124_3477_U718 ( .A(DP_OP_422J2_124_3477_n2019), .B(
        DP_OP_422J2_124_3477_n2026), .CI(DP_OP_422J2_124_3477_n2033), .CO(
        DP_OP_422J2_124_3477_n1122), .S(DP_OP_422J2_124_3477_n1123) );
  FADDX1_HVT DP_OP_422J2_124_3477_U717 ( .A(DP_OP_422J2_124_3477_n2811), .B(
        DP_OP_422J2_124_3477_n2063), .CI(DP_OP_422J2_124_3477_n2070), .CO(
        DP_OP_422J2_124_3477_n1120), .S(DP_OP_422J2_124_3477_n1121) );
  FADDX1_HVT DP_OP_422J2_124_3477_U716 ( .A(DP_OP_422J2_124_3477_n2781), .B(
        DP_OP_422J2_124_3477_n2077), .CI(DP_OP_422J2_124_3477_n2107), .CO(
        DP_OP_422J2_124_3477_n1118), .S(DP_OP_422J2_124_3477_n1119) );
  FADDX1_HVT DP_OP_422J2_124_3477_U715 ( .A(DP_OP_422J2_124_3477_n2774), .B(
        DP_OP_422J2_124_3477_n2114), .CI(DP_OP_422J2_124_3477_n2121), .CO(
        DP_OP_422J2_124_3477_n1116), .S(DP_OP_422J2_124_3477_n1117) );
  FADDX1_HVT DP_OP_422J2_124_3477_U714 ( .A(DP_OP_422J2_124_3477_n2767), .B(
        DP_OP_422J2_124_3477_n2151), .CI(DP_OP_422J2_124_3477_n2158), .CO(
        DP_OP_422J2_124_3477_n1114), .S(DP_OP_422J2_124_3477_n1115) );
  FADDX1_HVT DP_OP_422J2_124_3477_U713 ( .A(DP_OP_422J2_124_3477_n2737), .B(
        DP_OP_422J2_124_3477_n2165), .CI(DP_OP_422J2_124_3477_n2195), .CO(
        DP_OP_422J2_124_3477_n1112), .S(DP_OP_422J2_124_3477_n1113) );
  FADDX1_HVT DP_OP_422J2_124_3477_U712 ( .A(DP_OP_422J2_124_3477_n2730), .B(
        DP_OP_422J2_124_3477_n2202), .CI(DP_OP_422J2_124_3477_n2209), .CO(
        DP_OP_422J2_124_3477_n1110), .S(DP_OP_422J2_124_3477_n1111) );
  FADDX1_HVT DP_OP_422J2_124_3477_U711 ( .A(DP_OP_422J2_124_3477_n2723), .B(
        DP_OP_422J2_124_3477_n2341), .CI(DP_OP_422J2_124_3477_n2385), .CO(
        DP_OP_422J2_124_3477_n1108), .S(DP_OP_422J2_124_3477_n1109) );
  FADDX1_HVT DP_OP_422J2_124_3477_U710 ( .A(DP_OP_422J2_124_3477_n2693), .B(
        DP_OP_422J2_124_3477_n2415), .CI(DP_OP_422J2_124_3477_n2422), .CO(
        DP_OP_422J2_124_3477_n1106), .S(DP_OP_422J2_124_3477_n1107) );
  FADDX1_HVT DP_OP_422J2_124_3477_U709 ( .A(DP_OP_422J2_124_3477_n2686), .B(
        DP_OP_422J2_124_3477_n2429), .CI(DP_OP_422J2_124_3477_n2459), .CO(
        DP_OP_422J2_124_3477_n1104), .S(DP_OP_422J2_124_3477_n1105) );
  FADDX1_HVT DP_OP_422J2_124_3477_U708 ( .A(DP_OP_422J2_124_3477_n2679), .B(
        DP_OP_422J2_124_3477_n2466), .CI(DP_OP_422J2_124_3477_n2473), .CO(
        DP_OP_422J2_124_3477_n1102), .S(DP_OP_422J2_124_3477_n1103) );
  FADDX1_HVT DP_OP_422J2_124_3477_U707 ( .A(DP_OP_422J2_124_3477_n2649), .B(
        DP_OP_422J2_124_3477_n2503), .CI(DP_OP_422J2_124_3477_n2510), .CO(
        DP_OP_422J2_124_3477_n1100), .S(DP_OP_422J2_124_3477_n1101) );
  FADDX1_HVT DP_OP_422J2_124_3477_U706 ( .A(DP_OP_422J2_124_3477_n2642), .B(
        DP_OP_422J2_124_3477_n2517), .CI(DP_OP_422J2_124_3477_n2547), .CO(
        DP_OP_422J2_124_3477_n1098), .S(DP_OP_422J2_124_3477_n1099) );
  FADDX1_HVT DP_OP_422J2_124_3477_U705 ( .A(DP_OP_422J2_124_3477_n2635), .B(
        DP_OP_422J2_124_3477_n2554), .CI(DP_OP_422J2_124_3477_n2561), .CO(
        DP_OP_422J2_124_3477_n1096), .S(DP_OP_422J2_124_3477_n1097) );
  FADDX1_HVT DP_OP_422J2_124_3477_U704 ( .A(DP_OP_422J2_124_3477_n2591), .B(
        DP_OP_422J2_124_3477_n2598), .CI(DP_OP_422J2_124_3477_n2605), .CO(
        DP_OP_422J2_124_3477_n1094), .S(DP_OP_422J2_124_3477_n1095) );
  FADDX1_HVT DP_OP_422J2_124_3477_U703 ( .A(DP_OP_422J2_124_3477_n1348), .B(
        DP_OP_422J2_124_3477_n1336), .CI(DP_OP_422J2_124_3477_n1334), .CO(
        DP_OP_422J2_124_3477_n1092), .S(DP_OP_422J2_124_3477_n1093) );
  FADDX1_HVT DP_OP_422J2_124_3477_U702 ( .A(DP_OP_422J2_124_3477_n1332), .B(
        DP_OP_422J2_124_3477_n1338), .CI(DP_OP_422J2_124_3477_n1161), .CO(
        DP_OP_422J2_124_3477_n1090), .S(DP_OP_422J2_124_3477_n1091) );
  FADDX1_HVT DP_OP_422J2_124_3477_U701 ( .A(DP_OP_422J2_124_3477_n1342), .B(
        DP_OP_422J2_124_3477_n1346), .CI(DP_OP_422J2_124_3477_n1340), .CO(
        DP_OP_422J2_124_3477_n1088), .S(DP_OP_422J2_124_3477_n1089) );
  FADDX1_HVT DP_OP_422J2_124_3477_U700 ( .A(DP_OP_422J2_124_3477_n1344), .B(
        DP_OP_422J2_124_3477_n1308), .CI(DP_OP_422J2_124_3477_n1306), .CO(
        DP_OP_422J2_124_3477_n1086), .S(DP_OP_422J2_124_3477_n1087) );
  FADDX1_HVT DP_OP_422J2_124_3477_U699 ( .A(DP_OP_422J2_124_3477_n1310), .B(
        DP_OP_422J2_124_3477_n1282), .CI(DP_OP_422J2_124_3477_n1330), .CO(
        DP_OP_422J2_124_3477_n1084), .S(DP_OP_422J2_124_3477_n1085) );
  FADDX1_HVT DP_OP_422J2_124_3477_U698 ( .A(DP_OP_422J2_124_3477_n1302), .B(
        DP_OP_422J2_124_3477_n1284), .CI(DP_OP_422J2_124_3477_n1328), .CO(
        DP_OP_422J2_124_3477_n1082), .S(DP_OP_422J2_124_3477_n1083) );
  FADDX1_HVT DP_OP_422J2_124_3477_U697 ( .A(DP_OP_422J2_124_3477_n1300), .B(
        DP_OP_422J2_124_3477_n1286), .CI(DP_OP_422J2_124_3477_n1326), .CO(
        DP_OP_422J2_124_3477_n1080), .S(DP_OP_422J2_124_3477_n1081) );
  FADDX1_HVT DP_OP_422J2_124_3477_U696 ( .A(DP_OP_422J2_124_3477_n1296), .B(
        DP_OP_422J2_124_3477_n1324), .CI(DP_OP_422J2_124_3477_n1322), .CO(
        DP_OP_422J2_124_3477_n1078), .S(DP_OP_422J2_124_3477_n1079) );
  FADDX1_HVT DP_OP_422J2_124_3477_U695 ( .A(DP_OP_422J2_124_3477_n1290), .B(
        DP_OP_422J2_124_3477_n1320), .CI(DP_OP_422J2_124_3477_n1318), .CO(
        DP_OP_422J2_124_3477_n1076), .S(DP_OP_422J2_124_3477_n1077) );
  FADDX1_HVT DP_OP_422J2_124_3477_U694 ( .A(DP_OP_422J2_124_3477_n1298), .B(
        DP_OP_422J2_124_3477_n1316), .CI(DP_OP_422J2_124_3477_n1314), .CO(
        DP_OP_422J2_124_3477_n1074), .S(DP_OP_422J2_124_3477_n1075) );
  FADDX1_HVT DP_OP_422J2_124_3477_U693 ( .A(DP_OP_422J2_124_3477_n1292), .B(
        DP_OP_422J2_124_3477_n1312), .CI(DP_OP_422J2_124_3477_n1304), .CO(
        DP_OP_422J2_124_3477_n1072), .S(DP_OP_422J2_124_3477_n1073) );
  FADDX1_HVT DP_OP_422J2_124_3477_U692 ( .A(DP_OP_422J2_124_3477_n1294), .B(
        DP_OP_422J2_124_3477_n1288), .CI(DP_OP_422J2_124_3477_n1151), .CO(
        DP_OP_422J2_124_3477_n1070), .S(DP_OP_422J2_124_3477_n1071) );
  FADDX1_HVT DP_OP_422J2_124_3477_U691 ( .A(DP_OP_422J2_124_3477_n1147), .B(
        DP_OP_422J2_124_3477_n1145), .CI(DP_OP_422J2_124_3477_n1149), .CO(
        DP_OP_422J2_124_3477_n1068), .S(DP_OP_422J2_124_3477_n1069) );
  FADDX1_HVT DP_OP_422J2_124_3477_U690 ( .A(DP_OP_422J2_124_3477_n1157), .B(
        DP_OP_422J2_124_3477_n1155), .CI(DP_OP_422J2_124_3477_n1159), .CO(
        DP_OP_422J2_124_3477_n1066), .S(DP_OP_422J2_124_3477_n1067) );
  FADDX1_HVT DP_OP_422J2_124_3477_U689 ( .A(DP_OP_422J2_124_3477_n1153), .B(
        DP_OP_422J2_124_3477_n1101), .CI(DP_OP_422J2_124_3477_n1103), .CO(
        DP_OP_422J2_124_3477_n1064), .S(DP_OP_422J2_124_3477_n1065) );
  FADDX1_HVT DP_OP_422J2_124_3477_U688 ( .A(DP_OP_422J2_124_3477_n1099), .B(
        DP_OP_422J2_124_3477_n1135), .CI(DP_OP_422J2_124_3477_n1131), .CO(
        DP_OP_422J2_124_3477_n1062), .S(DP_OP_422J2_124_3477_n1063) );
  FADDX1_HVT DP_OP_422J2_124_3477_U687 ( .A(DP_OP_422J2_124_3477_n1137), .B(
        DP_OP_422J2_124_3477_n1121), .CI(DP_OP_422J2_124_3477_n1127), .CO(
        DP_OP_422J2_124_3477_n1060), .S(DP_OP_422J2_124_3477_n1061) );
  FADDX1_HVT DP_OP_422J2_124_3477_U686 ( .A(DP_OP_422J2_124_3477_n1125), .B(
        DP_OP_422J2_124_3477_n1123), .CI(DP_OP_422J2_124_3477_n1107), .CO(
        DP_OP_422J2_124_3477_n1058), .S(DP_OP_422J2_124_3477_n1059) );
  FADDX1_HVT DP_OP_422J2_124_3477_U685 ( .A(DP_OP_422J2_124_3477_n1129), .B(
        DP_OP_422J2_124_3477_n1097), .CI(DP_OP_422J2_124_3477_n1095), .CO(
        DP_OP_422J2_124_3477_n1056), .S(DP_OP_422J2_124_3477_n1057) );
  FADDX1_HVT DP_OP_422J2_124_3477_U684 ( .A(DP_OP_422J2_124_3477_n1133), .B(
        DP_OP_422J2_124_3477_n1115), .CI(DP_OP_422J2_124_3477_n1117), .CO(
        DP_OP_422J2_124_3477_n1054), .S(DP_OP_422J2_124_3477_n1055) );
  FADDX1_HVT DP_OP_422J2_124_3477_U683 ( .A(DP_OP_422J2_124_3477_n1113), .B(
        DP_OP_422J2_124_3477_n1111), .CI(DP_OP_422J2_124_3477_n1105), .CO(
        DP_OP_422J2_124_3477_n1052), .S(DP_OP_422J2_124_3477_n1053) );
  FADDX1_HVT DP_OP_422J2_124_3477_U682 ( .A(DP_OP_422J2_124_3477_n1109), .B(
        DP_OP_422J2_124_3477_n1143), .CI(DP_OP_422J2_124_3477_n1141), .CO(
        DP_OP_422J2_124_3477_n1050), .S(DP_OP_422J2_124_3477_n1051) );
  FADDX1_HVT DP_OP_422J2_124_3477_U681 ( .A(DP_OP_422J2_124_3477_n1139), .B(
        DP_OP_422J2_124_3477_n1119), .CI(DP_OP_422J2_124_3477_n1280), .CO(
        DP_OP_422J2_124_3477_n1048), .S(DP_OP_422J2_124_3477_n1049) );
  FADDX1_HVT DP_OP_422J2_124_3477_U680 ( .A(DP_OP_422J2_124_3477_n1278), .B(
        DP_OP_422J2_124_3477_n1276), .CI(DP_OP_422J2_124_3477_n1274), .CO(
        DP_OP_422J2_124_3477_n1046), .S(DP_OP_422J2_124_3477_n1047) );
  FADDX1_HVT DP_OP_422J2_124_3477_U679 ( .A(DP_OP_422J2_124_3477_n1272), .B(
        DP_OP_422J2_124_3477_n1260), .CI(DP_OP_422J2_124_3477_n1258), .CO(
        DP_OP_422J2_124_3477_n1044), .S(DP_OP_422J2_124_3477_n1045) );
  FADDX1_HVT DP_OP_422J2_124_3477_U678 ( .A(DP_OP_422J2_124_3477_n1264), .B(
        DP_OP_422J2_124_3477_n1262), .CI(DP_OP_422J2_124_3477_n1270), .CO(
        DP_OP_422J2_124_3477_n1042), .S(DP_OP_422J2_124_3477_n1043) );
  FADDX1_HVT DP_OP_422J2_124_3477_U677 ( .A(DP_OP_422J2_124_3477_n1268), .B(
        DP_OP_422J2_124_3477_n1266), .CI(DP_OP_422J2_124_3477_n1093), .CO(
        DP_OP_422J2_124_3477_n1040), .S(DP_OP_422J2_124_3477_n1041) );
  FADDX1_HVT DP_OP_422J2_124_3477_U676 ( .A(DP_OP_422J2_124_3477_n1256), .B(
        DP_OP_422J2_124_3477_n1254), .CI(DP_OP_422J2_124_3477_n1087), .CO(
        DP_OP_422J2_124_3477_n1038), .S(DP_OP_422J2_124_3477_n1039) );
  FADDX1_HVT DP_OP_422J2_124_3477_U675 ( .A(DP_OP_422J2_124_3477_n1091), .B(
        DP_OP_422J2_124_3477_n1089), .CI(DP_OP_422J2_124_3477_n1252), .CO(
        DP_OP_422J2_124_3477_n1036), .S(DP_OP_422J2_124_3477_n1037) );
  FADDX1_HVT DP_OP_422J2_124_3477_U674 ( .A(DP_OP_422J2_124_3477_n1240), .B(
        DP_OP_422J2_124_3477_n1085), .CI(DP_OP_422J2_124_3477_n1071), .CO(
        DP_OP_422J2_124_3477_n1034), .S(DP_OP_422J2_124_3477_n1035) );
  FADDX1_HVT DP_OP_422J2_124_3477_U673 ( .A(DP_OP_422J2_124_3477_n1238), .B(
        DP_OP_422J2_124_3477_n1081), .CI(DP_OP_422J2_124_3477_n1083), .CO(
        DP_OP_422J2_124_3477_n1032), .S(DP_OP_422J2_124_3477_n1033) );
  FADDX1_HVT DP_OP_422J2_124_3477_U672 ( .A(DP_OP_422J2_124_3477_n1242), .B(
        DP_OP_422J2_124_3477_n1079), .CI(DP_OP_422J2_124_3477_n1077), .CO(
        DP_OP_422J2_124_3477_n1030), .S(DP_OP_422J2_124_3477_n1031) );
  FADDX1_HVT DP_OP_422J2_124_3477_U671 ( .A(DP_OP_422J2_124_3477_n1250), .B(
        DP_OP_422J2_124_3477_n1073), .CI(DP_OP_422J2_124_3477_n1075), .CO(
        DP_OP_422J2_124_3477_n1028), .S(DP_OP_422J2_124_3477_n1029) );
  FADDX1_HVT DP_OP_422J2_124_3477_U670 ( .A(DP_OP_422J2_124_3477_n1248), .B(
        DP_OP_422J2_124_3477_n1244), .CI(DP_OP_422J2_124_3477_n1246), .CO(
        DP_OP_422J2_124_3477_n1026), .S(DP_OP_422J2_124_3477_n1027) );
  FADDX1_HVT DP_OP_422J2_124_3477_U669 ( .A(DP_OP_422J2_124_3477_n1067), .B(
        DP_OP_422J2_124_3477_n1236), .CI(DP_OP_422J2_124_3477_n1065), .CO(
        DP_OP_422J2_124_3477_n1024), .S(DP_OP_422J2_124_3477_n1025) );
  FADDX1_HVT DP_OP_422J2_124_3477_U668 ( .A(DP_OP_422J2_124_3477_n1069), .B(
        DP_OP_422J2_124_3477_n1059), .CI(DP_OP_422J2_124_3477_n1061), .CO(
        DP_OP_422J2_124_3477_n1022), .S(DP_OP_422J2_124_3477_n1023) );
  FADDX1_HVT DP_OP_422J2_124_3477_U667 ( .A(DP_OP_422J2_124_3477_n1057), .B(
        DP_OP_422J2_124_3477_n1051), .CI(DP_OP_422J2_124_3477_n1234), .CO(
        DP_OP_422J2_124_3477_n1020), .S(DP_OP_422J2_124_3477_n1021) );
  FADDX1_HVT DP_OP_422J2_124_3477_U666 ( .A(DP_OP_422J2_124_3477_n1053), .B(
        DP_OP_422J2_124_3477_n1063), .CI(DP_OP_422J2_124_3477_n1055), .CO(
        DP_OP_422J2_124_3477_n1018), .S(DP_OP_422J2_124_3477_n1019) );
  FADDX1_HVT DP_OP_422J2_124_3477_U665 ( .A(DP_OP_422J2_124_3477_n1049), .B(
        DP_OP_422J2_124_3477_n1232), .CI(DP_OP_422J2_124_3477_n1228), .CO(
        DP_OP_422J2_124_3477_n1016), .S(DP_OP_422J2_124_3477_n1017) );
  FADDX1_HVT DP_OP_422J2_124_3477_U664 ( .A(DP_OP_422J2_124_3477_n1230), .B(
        DP_OP_422J2_124_3477_n1226), .CI(DP_OP_422J2_124_3477_n1224), .CO(
        DP_OP_422J2_124_3477_n1014), .S(DP_OP_422J2_124_3477_n1015) );
  FADDX1_HVT DP_OP_422J2_124_3477_U663 ( .A(DP_OP_422J2_124_3477_n1047), .B(
        DP_OP_422J2_124_3477_n1222), .CI(DP_OP_422J2_124_3477_n1220), .CO(
        DP_OP_422J2_124_3477_n1012), .S(DP_OP_422J2_124_3477_n1013) );
  FADDX1_HVT DP_OP_422J2_124_3477_U662 ( .A(DP_OP_422J2_124_3477_n1218), .B(
        DP_OP_422J2_124_3477_n1043), .CI(DP_OP_422J2_124_3477_n1041), .CO(
        DP_OP_422J2_124_3477_n1010), .S(DP_OP_422J2_124_3477_n1011) );
  FADDX1_HVT DP_OP_422J2_124_3477_U661 ( .A(DP_OP_422J2_124_3477_n1216), .B(
        DP_OP_422J2_124_3477_n1214), .CI(DP_OP_422J2_124_3477_n1045), .CO(
        DP_OP_422J2_124_3477_n1008), .S(DP_OP_422J2_124_3477_n1009) );
  FADDX1_HVT DP_OP_422J2_124_3477_U660 ( .A(DP_OP_422J2_124_3477_n1037), .B(
        DP_OP_422J2_124_3477_n1212), .CI(DP_OP_422J2_124_3477_n1039), .CO(
        DP_OP_422J2_124_3477_n1006), .S(DP_OP_422J2_124_3477_n1007) );
  FADDX1_HVT DP_OP_422J2_124_3477_U659 ( .A(DP_OP_422J2_124_3477_n1031), .B(
        DP_OP_422J2_124_3477_n1035), .CI(DP_OP_422J2_124_3477_n1206), .CO(
        DP_OP_422J2_124_3477_n1004), .S(DP_OP_422J2_124_3477_n1005) );
  FADDX1_HVT DP_OP_422J2_124_3477_U658 ( .A(DP_OP_422J2_124_3477_n1210), .B(
        DP_OP_422J2_124_3477_n1029), .CI(DP_OP_422J2_124_3477_n1033), .CO(
        DP_OP_422J2_124_3477_n1002), .S(DP_OP_422J2_124_3477_n1003) );
  FADDX1_HVT DP_OP_422J2_124_3477_U657 ( .A(DP_OP_422J2_124_3477_n1208), .B(
        DP_OP_422J2_124_3477_n1027), .CI(DP_OP_422J2_124_3477_n1204), .CO(
        DP_OP_422J2_124_3477_n1000), .S(DP_OP_422J2_124_3477_n1001) );
  FADDX1_HVT DP_OP_422J2_124_3477_U656 ( .A(DP_OP_422J2_124_3477_n1025), .B(
        DP_OP_422J2_124_3477_n1023), .CI(DP_OP_422J2_124_3477_n1021), .CO(
        DP_OP_422J2_124_3477_n998), .S(DP_OP_422J2_124_3477_n999) );
  FADDX1_HVT DP_OP_422J2_124_3477_U655 ( .A(DP_OP_422J2_124_3477_n1019), .B(
        DP_OP_422J2_124_3477_n1202), .CI(DP_OP_422J2_124_3477_n1017), .CO(
        DP_OP_422J2_124_3477_n996), .S(DP_OP_422J2_124_3477_n997) );
  FADDX1_HVT DP_OP_422J2_124_3477_U654 ( .A(DP_OP_422J2_124_3477_n1200), .B(
        DP_OP_422J2_124_3477_n1198), .CI(DP_OP_422J2_124_3477_n1196), .CO(
        DP_OP_422J2_124_3477_n994), .S(DP_OP_422J2_124_3477_n995) );
  FADDX1_HVT DP_OP_422J2_124_3477_U653 ( .A(DP_OP_422J2_124_3477_n1015), .B(
        DP_OP_422J2_124_3477_n1194), .CI(DP_OP_422J2_124_3477_n1013), .CO(
        DP_OP_422J2_124_3477_n992), .S(DP_OP_422J2_124_3477_n993) );
  FADDX1_HVT DP_OP_422J2_124_3477_U652 ( .A(DP_OP_422J2_124_3477_n1192), .B(
        DP_OP_422J2_124_3477_n1009), .CI(DP_OP_422J2_124_3477_n1011), .CO(
        DP_OP_422J2_124_3477_n990), .S(DP_OP_422J2_124_3477_n991) );
  FADDX1_HVT DP_OP_422J2_124_3477_U651 ( .A(DP_OP_422J2_124_3477_n1190), .B(
        DP_OP_422J2_124_3477_n1188), .CI(DP_OP_422J2_124_3477_n1007), .CO(
        DP_OP_422J2_124_3477_n988), .S(DP_OP_422J2_124_3477_n989) );
  FADDX1_HVT DP_OP_422J2_124_3477_U650 ( .A(DP_OP_422J2_124_3477_n1186), .B(
        DP_OP_422J2_124_3477_n1003), .CI(DP_OP_422J2_124_3477_n1001), .CO(
        DP_OP_422J2_124_3477_n986), .S(DP_OP_422J2_124_3477_n987) );
  FADDX1_HVT DP_OP_422J2_124_3477_U649 ( .A(DP_OP_422J2_124_3477_n1005), .B(
        DP_OP_422J2_124_3477_n1184), .CI(DP_OP_422J2_124_3477_n999), .CO(
        DP_OP_422J2_124_3477_n984), .S(DP_OP_422J2_124_3477_n985) );
  FADDX1_HVT DP_OP_422J2_124_3477_U648 ( .A(DP_OP_422J2_124_3477_n1182), .B(
        DP_OP_422J2_124_3477_n997), .CI(DP_OP_422J2_124_3477_n1180), .CO(
        DP_OP_422J2_124_3477_n982), .S(DP_OP_422J2_124_3477_n983) );
  FADDX1_HVT DP_OP_422J2_124_3477_U647 ( .A(DP_OP_422J2_124_3477_n995), .B(
        DP_OP_422J2_124_3477_n1178), .CI(DP_OP_422J2_124_3477_n993), .CO(
        DP_OP_422J2_124_3477_n980), .S(DP_OP_422J2_124_3477_n981) );
  FADDX1_HVT DP_OP_422J2_124_3477_U646 ( .A(DP_OP_422J2_124_3477_n1176), .B(
        DP_OP_422J2_124_3477_n991), .CI(DP_OP_422J2_124_3477_n989), .CO(
        DP_OP_422J2_124_3477_n978), .S(DP_OP_422J2_124_3477_n979) );
  FADDX1_HVT DP_OP_422J2_124_3477_U645 ( .A(DP_OP_422J2_124_3477_n1174), .B(
        DP_OP_422J2_124_3477_n987), .CI(DP_OP_422J2_124_3477_n1172), .CO(
        DP_OP_422J2_124_3477_n976), .S(DP_OP_422J2_124_3477_n977) );
  FADDX1_HVT DP_OP_422J2_124_3477_U644 ( .A(DP_OP_422J2_124_3477_n985), .B(
        DP_OP_422J2_124_3477_n1170), .CI(DP_OP_422J2_124_3477_n983), .CO(
        DP_OP_422J2_124_3477_n974), .S(DP_OP_422J2_124_3477_n975) );
  FADDX1_HVT DP_OP_422J2_124_3477_U643 ( .A(DP_OP_422J2_124_3477_n981), .B(
        DP_OP_422J2_124_3477_n1168), .CI(DP_OP_422J2_124_3477_n979), .CO(
        DP_OP_422J2_124_3477_n972), .S(DP_OP_422J2_124_3477_n973) );
  FADDX1_HVT DP_OP_422J2_124_3477_U642 ( .A(DP_OP_422J2_124_3477_n1166), .B(
        DP_OP_422J2_124_3477_n977), .CI(DP_OP_422J2_124_3477_n975), .CO(
        DP_OP_422J2_124_3477_n970), .S(DP_OP_422J2_124_3477_n971) );
  FADDX1_HVT DP_OP_422J2_124_3477_U641 ( .A(DP_OP_422J2_124_3477_n1164), .B(
        DP_OP_422J2_124_3477_n973), .CI(DP_OP_422J2_124_3477_n1162), .CO(
        DP_OP_422J2_124_3477_n968), .S(DP_OP_422J2_124_3477_n969) );
  FADDX1_HVT DP_OP_422J2_124_3477_U640 ( .A(DP_OP_422J2_124_3477_n2978), .B(
        DP_OP_422J2_124_3477_n1923), .CI(DP_OP_422J2_124_3477_n1879), .CO(
        DP_OP_422J2_124_3477_n966), .S(DP_OP_422J2_124_3477_n967) );
  FADDX1_HVT DP_OP_422J2_124_3477_U639 ( .A(DP_OP_422J2_124_3477_n2803), .B(
        DP_OP_422J2_124_3477_n2120), .CI(DP_OP_422J2_124_3477_n2384), .CO(
        DP_OP_422J2_124_3477_n964), .S(DP_OP_422J2_124_3477_n965) );
  FADDX1_HVT DP_OP_422J2_124_3477_U638 ( .A(DP_OP_422J2_124_3477_n2011), .B(
        DP_OP_422J2_124_3477_n2428), .CI(DP_OP_422J2_124_3477_n1988), .CO(
        DP_OP_422J2_124_3477_n962), .S(DP_OP_422J2_124_3477_n963) );
  FADDX1_HVT DP_OP_422J2_124_3477_U637 ( .A(DP_OP_422J2_124_3477_n2319), .B(
        DP_OP_422J2_124_3477_n1944), .CI(DP_OP_422J2_124_3477_n2912), .CO(
        DP_OP_422J2_124_3477_n960), .S(DP_OP_422J2_124_3477_n961) );
  FADDX1_HVT DP_OP_422J2_124_3477_U636 ( .A(DP_OP_422J2_124_3477_n2275), .B(
        DP_OP_422J2_124_3477_n2252), .CI(DP_OP_422J2_124_3477_n2604), .CO(
        DP_OP_422J2_124_3477_n958), .S(DP_OP_422J2_124_3477_n959) );
  FADDX1_HVT DP_OP_422J2_124_3477_U635 ( .A(DP_OP_422J2_124_3477_n2187), .B(
        DP_OP_422J2_124_3477_n2296), .CI(DP_OP_422J2_124_3477_n2956), .CO(
        DP_OP_422J2_124_3477_n956), .S(DP_OP_422J2_124_3477_n957) );
  FADDX1_HVT DP_OP_422J2_124_3477_U634 ( .A(DP_OP_422J2_124_3477_n1967), .B(
        DP_OP_422J2_124_3477_n2032), .CI(DP_OP_422J2_124_3477_n2472), .CO(
        DP_OP_422J2_124_3477_n954), .S(DP_OP_422J2_124_3477_n955) );
  FADDX1_HVT DP_OP_422J2_124_3477_U633 ( .A(DP_OP_422J2_124_3477_n2055), .B(
        DP_OP_422J2_124_3477_n2736), .CI(DP_OP_422J2_124_3477_n2780), .CO(
        DP_OP_422J2_124_3477_n952), .S(DP_OP_422J2_124_3477_n953) );
  FADDX1_HVT DP_OP_422J2_124_3477_U632 ( .A(DP_OP_422J2_124_3477_n2143), .B(
        DP_OP_422J2_124_3477_n2692), .CI(DP_OP_422J2_124_3477_n2560), .CO(
        DP_OP_422J2_124_3477_n950), .S(DP_OP_422J2_124_3477_n951) );
  FADDX1_HVT DP_OP_422J2_124_3477_U631 ( .A(DP_OP_422J2_124_3477_n2495), .B(
        DP_OP_422J2_124_3477_n2340), .CI(DP_OP_422J2_124_3477_n2824), .CO(
        DP_OP_422J2_124_3477_n948), .S(DP_OP_422J2_124_3477_n949) );
  FADDX1_HVT DP_OP_422J2_124_3477_U630 ( .A(DP_OP_422J2_124_3477_n2891), .B(
        DP_OP_422J2_124_3477_n2164), .CI(DP_OP_422J2_124_3477_n2076), .CO(
        DP_OP_422J2_124_3477_n946), .S(DP_OP_422J2_124_3477_n947) );
  FADDX1_HVT DP_OP_422J2_124_3477_U629 ( .A(DP_OP_422J2_124_3477_n2627), .B(
        DP_OP_422J2_124_3477_n2868), .CI(DP_OP_422J2_124_3477_n2516), .CO(
        DP_OP_422J2_124_3477_n944), .S(DP_OP_422J2_124_3477_n945) );
  FADDX1_HVT DP_OP_422J2_124_3477_U628 ( .A(DP_OP_422J2_124_3477_n2407), .B(
        DP_OP_422J2_124_3477_n2998), .CI(DP_OP_422J2_124_3477_n2208), .CO(
        DP_OP_422J2_124_3477_n942), .S(DP_OP_422J2_124_3477_n943) );
  FADDX1_HVT DP_OP_422J2_124_3477_U627 ( .A(DP_OP_422J2_124_3477_n2099), .B(
        DP_OP_422J2_124_3477_n2363), .CI(DP_OP_422J2_124_3477_n2648), .CO(
        DP_OP_422J2_124_3477_n940), .S(DP_OP_422J2_124_3477_n941) );
  FADDX1_HVT DP_OP_422J2_124_3477_U626 ( .A(DP_OP_422J2_124_3477_n2715), .B(
        DP_OP_422J2_124_3477_n2759), .CI(DP_OP_422J2_124_3477_n2847), .CO(
        DP_OP_422J2_124_3477_n938), .S(DP_OP_422J2_124_3477_n939) );
  FADDX1_HVT DP_OP_422J2_124_3477_U625 ( .A(DP_OP_422J2_124_3477_n2451), .B(
        DP_OP_422J2_124_3477_n2539), .CI(DP_OP_422J2_124_3477_n2935), .CO(
        DP_OP_422J2_124_3477_n936), .S(DP_OP_422J2_124_3477_n937) );
  FADDX1_HVT DP_OP_422J2_124_3477_U624 ( .A(DP_OP_422J2_124_3477_n2583), .B(
        DP_OP_422J2_124_3477_n2231), .CI(DP_OP_422J2_124_3477_n2671), .CO(
        DP_OP_422J2_124_3477_n934), .S(DP_OP_422J2_124_3477_n935) );
  FADDX1_HVT DP_OP_422J2_124_3477_U623 ( .A(DP_OP_422J2_124_3477_n2991), .B(
        DP_OP_422J2_124_3477_n1937), .CI(DP_OP_422J2_124_3477_n1930), .CO(
        DP_OP_422J2_124_3477_n932), .S(DP_OP_422J2_124_3477_n933) );
  FADDX1_HVT DP_OP_422J2_124_3477_U622 ( .A(DP_OP_422J2_124_3477_n2984), .B(
        DP_OP_422J2_124_3477_n2949), .CI(DP_OP_422J2_124_3477_n2942), .CO(
        DP_OP_422J2_124_3477_n930), .S(DP_OP_422J2_124_3477_n931) );
  FADDX1_HVT DP_OP_422J2_124_3477_U621 ( .A(DP_OP_422J2_124_3477_n2465), .B(
        DP_OP_422J2_124_3477_n2905), .CI(DP_OP_422J2_124_3477_n2898), .CO(
        DP_OP_422J2_124_3477_n928), .S(DP_OP_422J2_124_3477_n929) );
  FADDX1_HVT DP_OP_422J2_124_3477_U620 ( .A(DP_OP_422J2_124_3477_n2861), .B(
        DP_OP_422J2_124_3477_n1974), .CI(DP_OP_422J2_124_3477_n1981), .CO(
        DP_OP_422J2_124_3477_n926), .S(DP_OP_422J2_124_3477_n927) );
  FADDX1_HVT DP_OP_422J2_124_3477_U619 ( .A(DP_OP_422J2_124_3477_n2854), .B(
        DP_OP_422J2_124_3477_n2018), .CI(DP_OP_422J2_124_3477_n2025), .CO(
        DP_OP_422J2_124_3477_n924), .S(DP_OP_422J2_124_3477_n925) );
  FADDX1_HVT DP_OP_422J2_124_3477_U618 ( .A(DP_OP_422J2_124_3477_n2817), .B(
        DP_OP_422J2_124_3477_n2062), .CI(DP_OP_422J2_124_3477_n2069), .CO(
        DP_OP_422J2_124_3477_n922), .S(DP_OP_422J2_124_3477_n923) );
  FADDX1_HVT DP_OP_422J2_124_3477_U617 ( .A(DP_OP_422J2_124_3477_n2810), .B(
        DP_OP_422J2_124_3477_n2106), .CI(DP_OP_422J2_124_3477_n2113), .CO(
        DP_OP_422J2_124_3477_n920), .S(DP_OP_422J2_124_3477_n921) );
  FADDX1_HVT DP_OP_422J2_124_3477_U616 ( .A(DP_OP_422J2_124_3477_n2773), .B(
        DP_OP_422J2_124_3477_n2150), .CI(DP_OP_422J2_124_3477_n2157), .CO(
        DP_OP_422J2_124_3477_n918), .S(DP_OP_422J2_124_3477_n919) );
  FADDX1_HVT DP_OP_422J2_124_3477_U615 ( .A(DP_OP_422J2_124_3477_n2766), .B(
        DP_OP_422J2_124_3477_n2194), .CI(DP_OP_422J2_124_3477_n2201), .CO(
        DP_OP_422J2_124_3477_n916), .S(DP_OP_422J2_124_3477_n917) );
  FADDX1_HVT DP_OP_422J2_124_3477_U614 ( .A(DP_OP_422J2_124_3477_n2729), .B(
        DP_OP_422J2_124_3477_n2238), .CI(DP_OP_422J2_124_3477_n2245), .CO(
        DP_OP_422J2_124_3477_n914), .S(DP_OP_422J2_124_3477_n915) );
  FADDX1_HVT DP_OP_422J2_124_3477_U613 ( .A(DP_OP_422J2_124_3477_n2722), .B(
        DP_OP_422J2_124_3477_n2282), .CI(DP_OP_422J2_124_3477_n2289), .CO(
        DP_OP_422J2_124_3477_n912), .S(DP_OP_422J2_124_3477_n913) );
  FADDX1_HVT DP_OP_422J2_124_3477_U612 ( .A(DP_OP_422J2_124_3477_n2685), .B(
        DP_OP_422J2_124_3477_n2326), .CI(DP_OP_422J2_124_3477_n2333), .CO(
        DP_OP_422J2_124_3477_n910), .S(DP_OP_422J2_124_3477_n911) );
  FADDX1_HVT DP_OP_422J2_124_3477_U611 ( .A(DP_OP_422J2_124_3477_n2678), .B(
        DP_OP_422J2_124_3477_n2370), .CI(DP_OP_422J2_124_3477_n2377), .CO(
        DP_OP_422J2_124_3477_n908), .S(DP_OP_422J2_124_3477_n909) );
  FADDX1_HVT DP_OP_422J2_124_3477_U610 ( .A(DP_OP_422J2_124_3477_n2641), .B(
        DP_OP_422J2_124_3477_n2414), .CI(DP_OP_422J2_124_3477_n2421), .CO(
        DP_OP_422J2_124_3477_n906), .S(DP_OP_422J2_124_3477_n907) );
  FADDX1_HVT DP_OP_422J2_124_3477_U609 ( .A(DP_OP_422J2_124_3477_n2634), .B(
        DP_OP_422J2_124_3477_n2458), .CI(DP_OP_422J2_124_3477_n2502), .CO(
        DP_OP_422J2_124_3477_n904), .S(DP_OP_422J2_124_3477_n905) );
  FADDX1_HVT DP_OP_422J2_124_3477_U608 ( .A(DP_OP_422J2_124_3477_n2597), .B(
        DP_OP_422J2_124_3477_n2509), .CI(DP_OP_422J2_124_3477_n2546), .CO(
        DP_OP_422J2_124_3477_n902), .S(DP_OP_422J2_124_3477_n903) );
  FADDX1_HVT DP_OP_422J2_124_3477_U607 ( .A(DP_OP_422J2_124_3477_n2590), .B(
        DP_OP_422J2_124_3477_n2553), .CI(DP_OP_422J2_124_3477_n1160), .CO(
        DP_OP_422J2_124_3477_n900), .S(DP_OP_422J2_124_3477_n901) );
  FADDX1_HVT DP_OP_422J2_124_3477_U606 ( .A(DP_OP_422J2_124_3477_n1148), .B(
        DP_OP_422J2_124_3477_n1144), .CI(DP_OP_422J2_124_3477_n1158), .CO(
        DP_OP_422J2_124_3477_n898), .S(DP_OP_422J2_124_3477_n899) );
  FADDX1_HVT DP_OP_422J2_124_3477_U605 ( .A(DP_OP_422J2_124_3477_n1156), .B(
        DP_OP_422J2_124_3477_n1146), .CI(DP_OP_422J2_124_3477_n1154), .CO(
        DP_OP_422J2_124_3477_n896), .S(DP_OP_422J2_124_3477_n897) );
  FADDX1_HVT DP_OP_422J2_124_3477_U604 ( .A(DP_OP_422J2_124_3477_n1152), .B(
        DP_OP_422J2_124_3477_n1150), .CI(DP_OP_422J2_124_3477_n1120), .CO(
        DP_OP_422J2_124_3477_n894), .S(DP_OP_422J2_124_3477_n895) );
  FADDX1_HVT DP_OP_422J2_124_3477_U603 ( .A(DP_OP_422J2_124_3477_n1118), .B(
        DP_OP_422J2_124_3477_n1094), .CI(DP_OP_422J2_124_3477_n1142), .CO(
        DP_OP_422J2_124_3477_n892), .S(DP_OP_422J2_124_3477_n893) );
  FADDX1_HVT DP_OP_422J2_124_3477_U602 ( .A(DP_OP_422J2_124_3477_n1116), .B(
        DP_OP_422J2_124_3477_n1140), .CI(DP_OP_422J2_124_3477_n1138), .CO(
        DP_OP_422J2_124_3477_n890), .S(DP_OP_422J2_124_3477_n891) );
  FADDX1_HVT DP_OP_422J2_124_3477_U601 ( .A(DP_OP_422J2_124_3477_n1110), .B(
        DP_OP_422J2_124_3477_n1136), .CI(DP_OP_422J2_124_3477_n1134), .CO(
        DP_OP_422J2_124_3477_n888), .S(DP_OP_422J2_124_3477_n889) );
  FADDX1_HVT DP_OP_422J2_124_3477_U600 ( .A(DP_OP_422J2_124_3477_n1132), .B(
        DP_OP_422J2_124_3477_n1130), .CI(DP_OP_422J2_124_3477_n1128), .CO(
        DP_OP_422J2_124_3477_n886), .S(DP_OP_422J2_124_3477_n887) );
  FADDX1_HVT DP_OP_422J2_124_3477_U599 ( .A(DP_OP_422J2_124_3477_n1100), .B(
        DP_OP_422J2_124_3477_n1126), .CI(DP_OP_422J2_124_3477_n1124), .CO(
        DP_OP_422J2_124_3477_n884), .S(DP_OP_422J2_124_3477_n885) );
  FADDX1_HVT DP_OP_422J2_124_3477_U598 ( .A(DP_OP_422J2_124_3477_n1106), .B(
        DP_OP_422J2_124_3477_n1122), .CI(DP_OP_422J2_124_3477_n1114), .CO(
        DP_OP_422J2_124_3477_n882), .S(DP_OP_422J2_124_3477_n883) );
  FADDX1_HVT DP_OP_422J2_124_3477_U597 ( .A(DP_OP_422J2_124_3477_n1098), .B(
        DP_OP_422J2_124_3477_n1112), .CI(DP_OP_422J2_124_3477_n1108), .CO(
        DP_OP_422J2_124_3477_n880), .S(DP_OP_422J2_124_3477_n881) );
  FADDX1_HVT DP_OP_422J2_124_3477_U596 ( .A(DP_OP_422J2_124_3477_n1102), .B(
        DP_OP_422J2_124_3477_n1096), .CI(DP_OP_422J2_124_3477_n1104), .CO(
        DP_OP_422J2_124_3477_n878), .S(DP_OP_422J2_124_3477_n879) );
  FADDX1_HVT DP_OP_422J2_124_3477_U595 ( .A(DP_OP_422J2_124_3477_n967), .B(
        DP_OP_422J2_124_3477_n953), .CI(DP_OP_422J2_124_3477_n955), .CO(
        DP_OP_422J2_124_3477_n876), .S(DP_OP_422J2_124_3477_n877) );
  FADDX1_HVT DP_OP_422J2_124_3477_U594 ( .A(DP_OP_422J2_124_3477_n959), .B(
        DP_OP_422J2_124_3477_n937), .CI(DP_OP_422J2_124_3477_n935), .CO(
        DP_OP_422J2_124_3477_n874), .S(DP_OP_422J2_124_3477_n875) );
  FADDX1_HVT DP_OP_422J2_124_3477_U593 ( .A(DP_OP_422J2_124_3477_n951), .B(
        DP_OP_422J2_124_3477_n949), .CI(DP_OP_422J2_124_3477_n945), .CO(
        DP_OP_422J2_124_3477_n872), .S(DP_OP_422J2_124_3477_n873) );
  FADDX1_HVT DP_OP_422J2_124_3477_U592 ( .A(DP_OP_422J2_124_3477_n957), .B(
        DP_OP_422J2_124_3477_n939), .CI(DP_OP_422J2_124_3477_n943), .CO(
        DP_OP_422J2_124_3477_n870), .S(DP_OP_422J2_124_3477_n871) );
  FADDX1_HVT DP_OP_422J2_124_3477_U591 ( .A(DP_OP_422J2_124_3477_n947), .B(
        DP_OP_422J2_124_3477_n965), .CI(DP_OP_422J2_124_3477_n961), .CO(
        DP_OP_422J2_124_3477_n868), .S(DP_OP_422J2_124_3477_n869) );
  FADDX1_HVT DP_OP_422J2_124_3477_U590 ( .A(DP_OP_422J2_124_3477_n941), .B(
        DP_OP_422J2_124_3477_n963), .CI(DP_OP_422J2_124_3477_n923), .CO(
        DP_OP_422J2_124_3477_n866), .S(DP_OP_422J2_124_3477_n867) );
  FADDX1_HVT DP_OP_422J2_124_3477_U589 ( .A(DP_OP_422J2_124_3477_n925), .B(
        DP_OP_422J2_124_3477_n907), .CI(DP_OP_422J2_124_3477_n901), .CO(
        DP_OP_422J2_124_3477_n864), .S(DP_OP_422J2_124_3477_n865) );
  FADDX1_HVT DP_OP_422J2_124_3477_U588 ( .A(DP_OP_422J2_124_3477_n927), .B(
        DP_OP_422J2_124_3477_n903), .CI(DP_OP_422J2_124_3477_n919), .CO(
        DP_OP_422J2_124_3477_n862), .S(DP_OP_422J2_124_3477_n863) );
  FADDX1_HVT DP_OP_422J2_124_3477_U587 ( .A(DP_OP_422J2_124_3477_n917), .B(
        DP_OP_422J2_124_3477_n915), .CI(DP_OP_422J2_124_3477_n905), .CO(
        DP_OP_422J2_124_3477_n860), .S(DP_OP_422J2_124_3477_n861) );
  FADDX1_HVT DP_OP_422J2_124_3477_U586 ( .A(DP_OP_422J2_124_3477_n921), .B(
        DP_OP_422J2_124_3477_n909), .CI(DP_OP_422J2_124_3477_n911), .CO(
        DP_OP_422J2_124_3477_n858), .S(DP_OP_422J2_124_3477_n859) );
  FADDX1_HVT DP_OP_422J2_124_3477_U585 ( .A(DP_OP_422J2_124_3477_n929), .B(
        DP_OP_422J2_124_3477_n933), .CI(DP_OP_422J2_124_3477_n931), .CO(
        DP_OP_422J2_124_3477_n856), .S(DP_OP_422J2_124_3477_n857) );
  FADDX1_HVT DP_OP_422J2_124_3477_U584 ( .A(DP_OP_422J2_124_3477_n913), .B(
        DP_OP_422J2_124_3477_n1092), .CI(DP_OP_422J2_124_3477_n1090), .CO(
        DP_OP_422J2_124_3477_n854), .S(DP_OP_422J2_124_3477_n855) );
  FADDX1_HVT DP_OP_422J2_124_3477_U583 ( .A(DP_OP_422J2_124_3477_n1088), .B(
        DP_OP_422J2_124_3477_n1086), .CI(DP_OP_422J2_124_3477_n1072), .CO(
        DP_OP_422J2_124_3477_n852), .S(DP_OP_422J2_124_3477_n853) );
  FADDX1_HVT DP_OP_422J2_124_3477_U582 ( .A(DP_OP_422J2_124_3477_n1084), .B(
        DP_OP_422J2_124_3477_n1082), .CI(DP_OP_422J2_124_3477_n1070), .CO(
        DP_OP_422J2_124_3477_n850), .S(DP_OP_422J2_124_3477_n851) );
  FADDX1_HVT DP_OP_422J2_124_3477_U581 ( .A(DP_OP_422J2_124_3477_n1080), .B(
        DP_OP_422J2_124_3477_n1074), .CI(DP_OP_422J2_124_3477_n1076), .CO(
        DP_OP_422J2_124_3477_n848), .S(DP_OP_422J2_124_3477_n849) );
  FADDX1_HVT DP_OP_422J2_124_3477_U580 ( .A(DP_OP_422J2_124_3477_n1078), .B(
        DP_OP_422J2_124_3477_n1068), .CI(DP_OP_422J2_124_3477_n1066), .CO(
        DP_OP_422J2_124_3477_n846), .S(DP_OP_422J2_124_3477_n847) );
  FADDX1_HVT DP_OP_422J2_124_3477_U579 ( .A(DP_OP_422J2_124_3477_n899), .B(
        DP_OP_422J2_124_3477_n895), .CI(DP_OP_422J2_124_3477_n1064), .CO(
        DP_OP_422J2_124_3477_n844), .S(DP_OP_422J2_124_3477_n845) );
  FADDX1_HVT DP_OP_422J2_124_3477_U578 ( .A(DP_OP_422J2_124_3477_n897), .B(
        DP_OP_422J2_124_3477_n1052), .CI(DP_OP_422J2_124_3477_n1050), .CO(
        DP_OP_422J2_124_3477_n842), .S(DP_OP_422J2_124_3477_n843) );
  FADDX1_HVT DP_OP_422J2_124_3477_U577 ( .A(DP_OP_422J2_124_3477_n1058), .B(
        DP_OP_422J2_124_3477_n893), .CI(DP_OP_422J2_124_3477_n1048), .CO(
        DP_OP_422J2_124_3477_n840), .S(DP_OP_422J2_124_3477_n841) );
  FADDX1_HVT DP_OP_422J2_124_3477_U576 ( .A(DP_OP_422J2_124_3477_n1056), .B(
        DP_OP_422J2_124_3477_n889), .CI(DP_OP_422J2_124_3477_n879), .CO(
        DP_OP_422J2_124_3477_n838), .S(DP_OP_422J2_124_3477_n839) );
  FADDX1_HVT DP_OP_422J2_124_3477_U575 ( .A(DP_OP_422J2_124_3477_n1062), .B(
        DP_OP_422J2_124_3477_n885), .CI(DP_OP_422J2_124_3477_n887), .CO(
        DP_OP_422J2_124_3477_n836), .S(DP_OP_422J2_124_3477_n837) );
  FADDX1_HVT DP_OP_422J2_124_3477_U574 ( .A(DP_OP_422J2_124_3477_n1060), .B(
        DP_OP_422J2_124_3477_n881), .CI(DP_OP_422J2_124_3477_n883), .CO(
        DP_OP_422J2_124_3477_n834), .S(DP_OP_422J2_124_3477_n835) );
  FADDX1_HVT DP_OP_422J2_124_3477_U573 ( .A(DP_OP_422J2_124_3477_n1054), .B(
        DP_OP_422J2_124_3477_n891), .CI(DP_OP_422J2_124_3477_n877), .CO(
        DP_OP_422J2_124_3477_n832), .S(DP_OP_422J2_124_3477_n833) );
  FADDX1_HVT DP_OP_422J2_124_3477_U572 ( .A(DP_OP_422J2_124_3477_n871), .B(
        DP_OP_422J2_124_3477_n875), .CI(DP_OP_422J2_124_3477_n867), .CO(
        DP_OP_422J2_124_3477_n830), .S(DP_OP_422J2_124_3477_n831) );
  FADDX1_HVT DP_OP_422J2_124_3477_U571 ( .A(DP_OP_422J2_124_3477_n869), .B(
        DP_OP_422J2_124_3477_n873), .CI(DP_OP_422J2_124_3477_n861), .CO(
        DP_OP_422J2_124_3477_n828), .S(DP_OP_422J2_124_3477_n829) );
  FADDX1_HVT DP_OP_422J2_124_3477_U570 ( .A(DP_OP_422J2_124_3477_n859), .B(
        DP_OP_422J2_124_3477_n865), .CI(DP_OP_422J2_124_3477_n1046), .CO(
        DP_OP_422J2_124_3477_n826), .S(DP_OP_422J2_124_3477_n827) );
  FADDX1_HVT DP_OP_422J2_124_3477_U569 ( .A(DP_OP_422J2_124_3477_n857), .B(
        DP_OP_422J2_124_3477_n863), .CI(DP_OP_422J2_124_3477_n1042), .CO(
        DP_OP_422J2_124_3477_n824), .S(DP_OP_422J2_124_3477_n825) );
  FADDX1_HVT DP_OP_422J2_124_3477_U568 ( .A(DP_OP_422J2_124_3477_n1044), .B(
        DP_OP_422J2_124_3477_n1040), .CI(DP_OP_422J2_124_3477_n855), .CO(
        DP_OP_422J2_124_3477_n822), .S(DP_OP_422J2_124_3477_n823) );
  FADDX1_HVT DP_OP_422J2_124_3477_U567 ( .A(DP_OP_422J2_124_3477_n1038), .B(
        DP_OP_422J2_124_3477_n1036), .CI(DP_OP_422J2_124_3477_n853), .CO(
        DP_OP_422J2_124_3477_n820), .S(DP_OP_422J2_124_3477_n821) );
  FADDX1_HVT DP_OP_422J2_124_3477_U566 ( .A(DP_OP_422J2_124_3477_n1034), .B(
        DP_OP_422J2_124_3477_n851), .CI(DP_OP_422J2_124_3477_n849), .CO(
        DP_OP_422J2_124_3477_n818), .S(DP_OP_422J2_124_3477_n819) );
  FADDX1_HVT DP_OP_422J2_124_3477_U565 ( .A(DP_OP_422J2_124_3477_n1032), .B(
        DP_OP_422J2_124_3477_n1026), .CI(DP_OP_422J2_124_3477_n1028), .CO(
        DP_OP_422J2_124_3477_n816), .S(DP_OP_422J2_124_3477_n817) );
  FADDX1_HVT DP_OP_422J2_124_3477_U564 ( .A(DP_OP_422J2_124_3477_n1030), .B(
        DP_OP_422J2_124_3477_n847), .CI(DP_OP_422J2_124_3477_n1024), .CO(
        DP_OP_422J2_124_3477_n814), .S(DP_OP_422J2_124_3477_n815) );
  FADDX1_HVT DP_OP_422J2_124_3477_U563 ( .A(DP_OP_422J2_124_3477_n845), .B(
        DP_OP_422J2_124_3477_n1022), .CI(DP_OP_422J2_124_3477_n843), .CO(
        DP_OP_422J2_124_3477_n812), .S(DP_OP_422J2_124_3477_n813) );
  FADDX1_HVT DP_OP_422J2_124_3477_U562 ( .A(DP_OP_422J2_124_3477_n1020), .B(
        DP_OP_422J2_124_3477_n837), .CI(DP_OP_422J2_124_3477_n833), .CO(
        DP_OP_422J2_124_3477_n810), .S(DP_OP_422J2_124_3477_n811) );
  FADDX1_HVT DP_OP_422J2_124_3477_U561 ( .A(DP_OP_422J2_124_3477_n1018), .B(
        DP_OP_422J2_124_3477_n841), .CI(DP_OP_422J2_124_3477_n839), .CO(
        DP_OP_422J2_124_3477_n808), .S(DP_OP_422J2_124_3477_n809) );
  FADDX1_HVT DP_OP_422J2_124_3477_U560 ( .A(DP_OP_422J2_124_3477_n835), .B(
        DP_OP_422J2_124_3477_n1016), .CI(DP_OP_422J2_124_3477_n831), .CO(
        DP_OP_422J2_124_3477_n806), .S(DP_OP_422J2_124_3477_n807) );
  FADDX1_HVT DP_OP_422J2_124_3477_U559 ( .A(DP_OP_422J2_124_3477_n829), .B(
        DP_OP_422J2_124_3477_n1014), .CI(DP_OP_422J2_124_3477_n827), .CO(
        DP_OP_422J2_124_3477_n804), .S(DP_OP_422J2_124_3477_n805) );
  FADDX1_HVT DP_OP_422J2_124_3477_U558 ( .A(DP_OP_422J2_124_3477_n825), .B(
        DP_OP_422J2_124_3477_n1012), .CI(DP_OP_422J2_124_3477_n1008), .CO(
        DP_OP_422J2_124_3477_n802), .S(DP_OP_422J2_124_3477_n803) );
  FADDX1_HVT DP_OP_422J2_124_3477_U557 ( .A(DP_OP_422J2_124_3477_n1010), .B(
        DP_OP_422J2_124_3477_n823), .CI(DP_OP_422J2_124_3477_n1006), .CO(
        DP_OP_422J2_124_3477_n800), .S(DP_OP_422J2_124_3477_n801) );
  FADDX1_HVT DP_OP_422J2_124_3477_U556 ( .A(DP_OP_422J2_124_3477_n821), .B(
        DP_OP_422J2_124_3477_n1004), .CI(DP_OP_422J2_124_3477_n1002), .CO(
        DP_OP_422J2_124_3477_n798), .S(DP_OP_422J2_124_3477_n799) );
  FADDX1_HVT DP_OP_422J2_124_3477_U555 ( .A(DP_OP_422J2_124_3477_n819), .B(
        DP_OP_422J2_124_3477_n1000), .CI(DP_OP_422J2_124_3477_n815), .CO(
        DP_OP_422J2_124_3477_n796), .S(DP_OP_422J2_124_3477_n797) );
  FADDX1_HVT DP_OP_422J2_124_3477_U554 ( .A(DP_OP_422J2_124_3477_n817), .B(
        DP_OP_422J2_124_3477_n998), .CI(DP_OP_422J2_124_3477_n813), .CO(
        DP_OP_422J2_124_3477_n794), .S(DP_OP_422J2_124_3477_n795) );
  FADDX1_HVT DP_OP_422J2_124_3477_U553 ( .A(DP_OP_422J2_124_3477_n996), .B(
        DP_OP_422J2_124_3477_n811), .CI(DP_OP_422J2_124_3477_n807), .CO(
        DP_OP_422J2_124_3477_n792), .S(DP_OP_422J2_124_3477_n793) );
  FADDX1_HVT DP_OP_422J2_124_3477_U552 ( .A(DP_OP_422J2_124_3477_n809), .B(
        DP_OP_422J2_124_3477_n994), .CI(DP_OP_422J2_124_3477_n805), .CO(
        DP_OP_422J2_124_3477_n790), .S(DP_OP_422J2_124_3477_n791) );
  FADDX1_HVT DP_OP_422J2_124_3477_U551 ( .A(DP_OP_422J2_124_3477_n992), .B(
        DP_OP_422J2_124_3477_n803), .CI(DP_OP_422J2_124_3477_n990), .CO(
        DP_OP_422J2_124_3477_n788), .S(DP_OP_422J2_124_3477_n789) );
  FADDX1_HVT DP_OP_422J2_124_3477_U550 ( .A(DP_OP_422J2_124_3477_n801), .B(
        DP_OP_422J2_124_3477_n988), .CI(DP_OP_422J2_124_3477_n799), .CO(
        DP_OP_422J2_124_3477_n786), .S(DP_OP_422J2_124_3477_n787) );
  FADDX1_HVT DP_OP_422J2_124_3477_U549 ( .A(DP_OP_422J2_124_3477_n986), .B(
        DP_OP_422J2_124_3477_n797), .CI(DP_OP_422J2_124_3477_n984), .CO(
        DP_OP_422J2_124_3477_n784), .S(DP_OP_422J2_124_3477_n785) );
  FADDX1_HVT DP_OP_422J2_124_3477_U548 ( .A(DP_OP_422J2_124_3477_n795), .B(
        DP_OP_422J2_124_3477_n793), .CI(DP_OP_422J2_124_3477_n982), .CO(
        DP_OP_422J2_124_3477_n782), .S(DP_OP_422J2_124_3477_n783) );
  FADDX1_HVT DP_OP_422J2_124_3477_U547 ( .A(DP_OP_422J2_124_3477_n791), .B(
        DP_OP_422J2_124_3477_n980), .CI(DP_OP_422J2_124_3477_n789), .CO(
        DP_OP_422J2_124_3477_n780), .S(DP_OP_422J2_124_3477_n781) );
  FADDX1_HVT DP_OP_422J2_124_3477_U546 ( .A(DP_OP_422J2_124_3477_n978), .B(
        DP_OP_422J2_124_3477_n787), .CI(DP_OP_422J2_124_3477_n976), .CO(
        DP_OP_422J2_124_3477_n778), .S(DP_OP_422J2_124_3477_n779) );
  FADDX1_HVT DP_OP_422J2_124_3477_U545 ( .A(DP_OP_422J2_124_3477_n785), .B(
        DP_OP_422J2_124_3477_n974), .CI(DP_OP_422J2_124_3477_n783), .CO(
        DP_OP_422J2_124_3477_n776), .S(DP_OP_422J2_124_3477_n777) );
  FADDX1_HVT DP_OP_422J2_124_3477_U544 ( .A(DP_OP_422J2_124_3477_n781), .B(
        DP_OP_422J2_124_3477_n972), .CI(DP_OP_422J2_124_3477_n779), .CO(
        DP_OP_422J2_124_3477_n774), .S(DP_OP_422J2_124_3477_n775) );
  FADDX1_HVT DP_OP_422J2_124_3477_U543 ( .A(DP_OP_422J2_124_3477_n970), .B(
        DP_OP_422J2_124_3477_n777), .CI(DP_OP_422J2_124_3477_n775), .CO(
        DP_OP_422J2_124_3477_n772), .S(DP_OP_422J2_124_3477_n773) );
  FADDX1_HVT DP_OP_422J2_124_3477_U541 ( .A(DP_OP_422J2_124_3477_n2186), .B(
        DP_OP_422J2_124_3477_n1922), .CI(DP_OP_422J2_124_3477_n1878), .CO(
        DP_OP_422J2_124_3477_n768), .S(DP_OP_422J2_124_3477_n769) );
  FADDX1_HVT DP_OP_422J2_124_3477_U540 ( .A(DP_OP_422J2_124_3477_n2758), .B(
        DP_OP_422J2_124_3477_n1980), .CI(DP_OP_422J2_124_3477_n2244), .CO(
        DP_OP_422J2_124_3477_n766), .S(DP_OP_422J2_124_3477_n767) );
  FADDX1_HVT DP_OP_422J2_124_3477_U539 ( .A(DP_OP_422J2_124_3477_n2230), .B(
        DP_OP_422J2_124_3477_n2990), .CI(DP_OP_422J2_124_3477_n2640), .CO(
        DP_OP_422J2_124_3477_n764), .S(DP_OP_422J2_124_3477_n765) );
  FADDX1_HVT DP_OP_422J2_124_3477_U538 ( .A(DP_OP_422J2_124_3477_n2450), .B(
        DP_OP_422J2_124_3477_n2024), .CI(DP_OP_422J2_124_3477_n2068), .CO(
        DP_OP_422J2_124_3477_n762), .S(DP_OP_422J2_124_3477_n763) );
  FADDX1_HVT DP_OP_422J2_124_3477_U537 ( .A(DP_OP_422J2_124_3477_n2010), .B(
        DP_OP_422J2_124_3477_n2112), .CI(DP_OP_422J2_124_3477_n2156), .CO(
        DP_OP_422J2_124_3477_n760), .S(DP_OP_422J2_124_3477_n761) );
  FADDX1_HVT DP_OP_422J2_124_3477_U536 ( .A(DP_OP_422J2_124_3477_n2714), .B(
        DP_OP_422J2_124_3477_n2816), .CI(DP_OP_422J2_124_3477_n2860), .CO(
        DP_OP_422J2_124_3477_n758), .S(DP_OP_422J2_124_3477_n759) );
  FADDX1_HVT DP_OP_422J2_124_3477_U535 ( .A(DP_OP_422J2_124_3477_n2054), .B(
        DP_OP_422J2_124_3477_n2772), .CI(DP_OP_422J2_124_3477_n2596), .CO(
        DP_OP_422J2_124_3477_n756), .S(DP_OP_422J2_124_3477_n757) );
  FADDX1_HVT DP_OP_422J2_124_3477_U534 ( .A(DP_OP_422J2_124_3477_n2142), .B(
        DP_OP_422J2_124_3477_n2420), .CI(DP_OP_422J2_124_3477_n2948), .CO(
        DP_OP_422J2_124_3477_n754), .S(DP_OP_422J2_124_3477_n755) );
  FADDX1_HVT DP_OP_422J2_124_3477_U533 ( .A(DP_OP_422J2_124_3477_n2670), .B(
        DP_OP_422J2_124_3477_n2904), .CI(DP_OP_422J2_124_3477_n2464), .CO(
        DP_OP_422J2_124_3477_n752), .S(DP_OP_422J2_124_3477_n753) );
  FADDX1_HVT DP_OP_422J2_124_3477_U532 ( .A(DP_OP_422J2_124_3477_n2626), .B(
        DP_OP_422J2_124_3477_n2376), .CI(DP_OP_422J2_124_3477_n2728), .CO(
        DP_OP_422J2_124_3477_n750), .S(DP_OP_422J2_124_3477_n751) );
  FADDX1_HVT DP_OP_422J2_124_3477_U531 ( .A(DP_OP_422J2_124_3477_n2846), .B(
        DP_OP_422J2_124_3477_n2508), .CI(DP_OP_422J2_124_3477_n2332), .CO(
        DP_OP_422J2_124_3477_n748), .S(DP_OP_422J2_124_3477_n749) );
  FADDX1_HVT DP_OP_422J2_124_3477_U530 ( .A(DP_OP_422J2_124_3477_n2318), .B(
        DP_OP_422J2_124_3477_n2288), .CI(DP_OP_422J2_124_3477_n1936), .CO(
        DP_OP_422J2_124_3477_n746), .S(DP_OP_422J2_124_3477_n747) );
  FADDX1_HVT DP_OP_422J2_124_3477_U529 ( .A(DP_OP_422J2_124_3477_n2538), .B(
        DP_OP_422J2_124_3477_n2200), .CI(DP_OP_422J2_124_3477_n2552), .CO(
        DP_OP_422J2_124_3477_n744), .S(DP_OP_422J2_124_3477_n745) );
  FADDX1_HVT DP_OP_422J2_124_3477_U528 ( .A(DP_OP_422J2_124_3477_n2494), .B(
        DP_OP_422J2_124_3477_n2362), .CI(DP_OP_422J2_124_3477_n2684), .CO(
        DP_OP_422J2_124_3477_n742), .S(DP_OP_422J2_124_3477_n743) );
  FADDX1_HVT DP_OP_422J2_124_3477_U527 ( .A(DP_OP_422J2_124_3477_n2802), .B(
        DP_OP_422J2_124_3477_n2098), .CI(DP_OP_422J2_124_3477_n2274), .CO(
        DP_OP_422J2_124_3477_n740), .S(DP_OP_422J2_124_3477_n741) );
  FADDX1_HVT DP_OP_422J2_124_3477_U526 ( .A(DP_OP_422J2_124_3477_n1966), .B(
        DP_OP_422J2_124_3477_n2582), .CI(DP_OP_422J2_124_3477_n2934), .CO(
        DP_OP_422J2_124_3477_n738), .S(DP_OP_422J2_124_3477_n739) );
  FADDX1_HVT DP_OP_422J2_124_3477_U525 ( .A(DP_OP_422J2_124_3477_n2890), .B(
        DP_OP_422J2_124_3477_n2406), .CI(DP_OP_422J2_124_3477_n771), .CO(
        DP_OP_422J2_124_3477_n736), .S(DP_OP_422J2_124_3477_n737) );
  FADDX1_HVT DP_OP_422J2_124_3477_U524 ( .A(DP_OP_422J2_124_3477_n2237), .B(
        DP_OP_422J2_124_3477_n1973), .CI(DP_OP_422J2_124_3477_n1929), .CO(
        DP_OP_422J2_124_3477_n734), .S(DP_OP_422J2_124_3477_n735) );
  FADDX1_HVT DP_OP_422J2_124_3477_U523 ( .A(DP_OP_422J2_124_3477_n2983), .B(
        DP_OP_422J2_124_3477_n2017), .CI(DP_OP_422J2_124_3477_n2061), .CO(
        DP_OP_422J2_124_3477_n732), .S(DP_OP_422J2_124_3477_n733) );
  FADDX1_HVT DP_OP_422J2_124_3477_U522 ( .A(DP_OP_422J2_124_3477_n2941), .B(
        DP_OP_422J2_124_3477_n2105), .CI(DP_OP_422J2_124_3477_n2149), .CO(
        DP_OP_422J2_124_3477_n730), .S(DP_OP_422J2_124_3477_n731) );
  FADDX1_HVT DP_OP_422J2_124_3477_U521 ( .A(DP_OP_422J2_124_3477_n2897), .B(
        DP_OP_422J2_124_3477_n2193), .CI(DP_OP_422J2_124_3477_n2281), .CO(
        DP_OP_422J2_124_3477_n728), .S(DP_OP_422J2_124_3477_n729) );
  FADDX1_HVT DP_OP_422J2_124_3477_U520 ( .A(DP_OP_422J2_124_3477_n2853), .B(
        DP_OP_422J2_124_3477_n2325), .CI(DP_OP_422J2_124_3477_n2369), .CO(
        DP_OP_422J2_124_3477_n726), .S(DP_OP_422J2_124_3477_n727) );
  FADDX1_HVT DP_OP_422J2_124_3477_U519 ( .A(DP_OP_422J2_124_3477_n2809), .B(
        DP_OP_422J2_124_3477_n2413), .CI(DP_OP_422J2_124_3477_n2457), .CO(
        DP_OP_422J2_124_3477_n724), .S(DP_OP_422J2_124_3477_n725) );
  FADDX1_HVT DP_OP_422J2_124_3477_U518 ( .A(DP_OP_422J2_124_3477_n2765), .B(
        DP_OP_422J2_124_3477_n2501), .CI(DP_OP_422J2_124_3477_n2545), .CO(
        DP_OP_422J2_124_3477_n722), .S(DP_OP_422J2_124_3477_n723) );
  FADDX1_HVT DP_OP_422J2_124_3477_U517 ( .A(DP_OP_422J2_124_3477_n2721), .B(
        DP_OP_422J2_124_3477_n2589), .CI(DP_OP_422J2_124_3477_n2633), .CO(
        DP_OP_422J2_124_3477_n720), .S(DP_OP_422J2_124_3477_n721) );
  FADDX1_HVT DP_OP_422J2_124_3477_U516 ( .A(DP_OP_422J2_124_3477_n2677), .B(
        DP_OP_422J2_124_3477_n966), .CI(DP_OP_422J2_124_3477_n964), .CO(
        DP_OP_422J2_124_3477_n718), .S(DP_OP_422J2_124_3477_n719) );
  FADDX1_HVT DP_OP_422J2_124_3477_U515 ( .A(DP_OP_422J2_124_3477_n962), .B(
        DP_OP_422J2_124_3477_n934), .CI(DP_OP_422J2_124_3477_n936), .CO(
        DP_OP_422J2_124_3477_n716), .S(DP_OP_422J2_124_3477_n717) );
  FADDX1_HVT DP_OP_422J2_124_3477_U514 ( .A(DP_OP_422J2_124_3477_n960), .B(
        DP_OP_422J2_124_3477_n938), .CI(DP_OP_422J2_124_3477_n940), .CO(
        DP_OP_422J2_124_3477_n714), .S(DP_OP_422J2_124_3477_n715) );
  FADDX1_HVT DP_OP_422J2_124_3477_U513 ( .A(DP_OP_422J2_124_3477_n958), .B(
        DP_OP_422J2_124_3477_n942), .CI(DP_OP_422J2_124_3477_n944), .CO(
        DP_OP_422J2_124_3477_n712), .S(DP_OP_422J2_124_3477_n713) );
  FADDX1_HVT DP_OP_422J2_124_3477_U512 ( .A(DP_OP_422J2_124_3477_n950), .B(
        DP_OP_422J2_124_3477_n956), .CI(DP_OP_422J2_124_3477_n946), .CO(
        DP_OP_422J2_124_3477_n710), .S(DP_OP_422J2_124_3477_n711) );
  FADDX1_HVT DP_OP_422J2_124_3477_U511 ( .A(DP_OP_422J2_124_3477_n948), .B(
        DP_OP_422J2_124_3477_n952), .CI(DP_OP_422J2_124_3477_n954), .CO(
        DP_OP_422J2_124_3477_n708), .S(DP_OP_422J2_124_3477_n709) );
  FADDX1_HVT DP_OP_422J2_124_3477_U510 ( .A(DP_OP_422J2_124_3477_n932), .B(
        DP_OP_422J2_124_3477_n930), .CI(DP_OP_422J2_124_3477_n900), .CO(
        DP_OP_422J2_124_3477_n706), .S(DP_OP_422J2_124_3477_n707) );
  FADDX1_HVT DP_OP_422J2_124_3477_U509 ( .A(DP_OP_422J2_124_3477_n914), .B(
        DP_OP_422J2_124_3477_n902), .CI(DP_OP_422J2_124_3477_n904), .CO(
        DP_OP_422J2_124_3477_n704), .S(DP_OP_422J2_124_3477_n705) );
  FADDX1_HVT DP_OP_422J2_124_3477_U508 ( .A(DP_OP_422J2_124_3477_n912), .B(
        DP_OP_422J2_124_3477_n906), .CI(DP_OP_422J2_124_3477_n908), .CO(
        DP_OP_422J2_124_3477_n702), .S(DP_OP_422J2_124_3477_n703) );
  FADDX1_HVT DP_OP_422J2_124_3477_U507 ( .A(DP_OP_422J2_124_3477_n910), .B(
        DP_OP_422J2_124_3477_n928), .CI(DP_OP_422J2_124_3477_n926), .CO(
        DP_OP_422J2_124_3477_n700), .S(DP_OP_422J2_124_3477_n701) );
  FADDX1_HVT DP_OP_422J2_124_3477_U506 ( .A(DP_OP_422J2_124_3477_n920), .B(
        DP_OP_422J2_124_3477_n916), .CI(DP_OP_422J2_124_3477_n918), .CO(
        DP_OP_422J2_124_3477_n698), .S(DP_OP_422J2_124_3477_n699) );
  FADDX1_HVT DP_OP_422J2_124_3477_U505 ( .A(DP_OP_422J2_124_3477_n924), .B(
        DP_OP_422J2_124_3477_n922), .CI(DP_OP_422J2_124_3477_n763), .CO(
        DP_OP_422J2_124_3477_n696), .S(DP_OP_422J2_124_3477_n697) );
  FADDX1_HVT DP_OP_422J2_124_3477_U504 ( .A(DP_OP_422J2_124_3477_n759), .B(
        DP_OP_422J2_124_3477_n755), .CI(DP_OP_422J2_124_3477_n737), .CO(
        DP_OP_422J2_124_3477_n694), .S(DP_OP_422J2_124_3477_n695) );
  FADDX1_HVT DP_OP_422J2_124_3477_U503 ( .A(DP_OP_422J2_124_3477_n761), .B(
        DP_OP_422J2_124_3477_n743), .CI(DP_OP_422J2_124_3477_n741), .CO(
        DP_OP_422J2_124_3477_n692), .S(DP_OP_422J2_124_3477_n693) );
  FADDX1_HVT DP_OP_422J2_124_3477_U502 ( .A(DP_OP_422J2_124_3477_n753), .B(
        DP_OP_422J2_124_3477_n757), .CI(DP_OP_422J2_124_3477_n749), .CO(
        DP_OP_422J2_124_3477_n690), .S(DP_OP_422J2_124_3477_n691) );
  FADDX1_HVT DP_OP_422J2_124_3477_U501 ( .A(DP_OP_422J2_124_3477_n765), .B(
        DP_OP_422J2_124_3477_n745), .CI(DP_OP_422J2_124_3477_n739), .CO(
        DP_OP_422J2_124_3477_n688), .S(DP_OP_422J2_124_3477_n689) );
  FADDX1_HVT DP_OP_422J2_124_3477_U500 ( .A(DP_OP_422J2_124_3477_n747), .B(
        DP_OP_422J2_124_3477_n769), .CI(DP_OP_422J2_124_3477_n767), .CO(
        DP_OP_422J2_124_3477_n686), .S(DP_OP_422J2_124_3477_n687) );
  FADDX1_HVT DP_OP_422J2_124_3477_U499 ( .A(DP_OP_422J2_124_3477_n751), .B(
        DP_OP_422J2_124_3477_n731), .CI(DP_OP_422J2_124_3477_n727), .CO(
        DP_OP_422J2_124_3477_n684), .S(DP_OP_422J2_124_3477_n685) );
  FADDX1_HVT DP_OP_422J2_124_3477_U498 ( .A(DP_OP_422J2_124_3477_n723), .B(
        DP_OP_422J2_124_3477_n721), .CI(DP_OP_422J2_124_3477_n733), .CO(
        DP_OP_422J2_124_3477_n682), .S(DP_OP_422J2_124_3477_n683) );
  FADDX1_HVT DP_OP_422J2_124_3477_U497 ( .A(DP_OP_422J2_124_3477_n729), .B(
        DP_OP_422J2_124_3477_n725), .CI(DP_OP_422J2_124_3477_n735), .CO(
        DP_OP_422J2_124_3477_n680), .S(DP_OP_422J2_124_3477_n681) );
  FADDX1_HVT DP_OP_422J2_124_3477_U496 ( .A(DP_OP_422J2_124_3477_n898), .B(
        DP_OP_422J2_124_3477_n894), .CI(DP_OP_422J2_124_3477_n896), .CO(
        DP_OP_422J2_124_3477_n678), .S(DP_OP_422J2_124_3477_n679) );
  FADDX1_HVT DP_OP_422J2_124_3477_U495 ( .A(DP_OP_422J2_124_3477_n892), .B(
        DP_OP_422J2_124_3477_n878), .CI(DP_OP_422J2_124_3477_n880), .CO(
        DP_OP_422J2_124_3477_n676), .S(DP_OP_422J2_124_3477_n677) );
  FADDX1_HVT DP_OP_422J2_124_3477_U494 ( .A(DP_OP_422J2_124_3477_n890), .B(
        DP_OP_422J2_124_3477_n882), .CI(DP_OP_422J2_124_3477_n888), .CO(
        DP_OP_422J2_124_3477_n674), .S(DP_OP_422J2_124_3477_n675) );
  FADDX1_HVT DP_OP_422J2_124_3477_U493 ( .A(DP_OP_422J2_124_3477_n886), .B(
        DP_OP_422J2_124_3477_n884), .CI(DP_OP_422J2_124_3477_n719), .CO(
        DP_OP_422J2_124_3477_n672), .S(DP_OP_422J2_124_3477_n673) );
  FADDX1_HVT DP_OP_422J2_124_3477_U492 ( .A(DP_OP_422J2_124_3477_n876), .B(
        DP_OP_422J2_124_3477_n717), .CI(DP_OP_422J2_124_3477_n715), .CO(
        DP_OP_422J2_124_3477_n670), .S(DP_OP_422J2_124_3477_n671) );
  FADDX1_HVT DP_OP_422J2_124_3477_U491 ( .A(DP_OP_422J2_124_3477_n874), .B(
        DP_OP_422J2_124_3477_n711), .CI(DP_OP_422J2_124_3477_n713), .CO(
        DP_OP_422J2_124_3477_n668), .S(DP_OP_422J2_124_3477_n669) );
  FADDX1_HVT DP_OP_422J2_124_3477_U490 ( .A(DP_OP_422J2_124_3477_n872), .B(
        DP_OP_422J2_124_3477_n709), .CI(DP_OP_422J2_124_3477_n866), .CO(
        DP_OP_422J2_124_3477_n666), .S(DP_OP_422J2_124_3477_n667) );
  FADDX1_HVT DP_OP_422J2_124_3477_U489 ( .A(DP_OP_422J2_124_3477_n870), .B(
        DP_OP_422J2_124_3477_n868), .CI(DP_OP_422J2_124_3477_n856), .CO(
        DP_OP_422J2_124_3477_n664), .S(DP_OP_422J2_124_3477_n665) );
  FADDX1_HVT DP_OP_422J2_124_3477_U488 ( .A(DP_OP_422J2_124_3477_n864), .B(
        DP_OP_422J2_124_3477_n707), .CI(DP_OP_422J2_124_3477_n697), .CO(
        DP_OP_422J2_124_3477_n662), .S(DP_OP_422J2_124_3477_n663) );
  FADDX1_HVT DP_OP_422J2_124_3477_U487 ( .A(DP_OP_422J2_124_3477_n862), .B(
        DP_OP_422J2_124_3477_n703), .CI(DP_OP_422J2_124_3477_n699), .CO(
        DP_OP_422J2_124_3477_n660), .S(DP_OP_422J2_124_3477_n661) );
  FADDX1_HVT DP_OP_422J2_124_3477_U486 ( .A(DP_OP_422J2_124_3477_n860), .B(
        DP_OP_422J2_124_3477_n705), .CI(DP_OP_422J2_124_3477_n701), .CO(
        DP_OP_422J2_124_3477_n658), .S(DP_OP_422J2_124_3477_n659) );
  FADDX1_HVT DP_OP_422J2_124_3477_U485 ( .A(DP_OP_422J2_124_3477_n858), .B(
        DP_OP_422J2_124_3477_n693), .CI(DP_OP_422J2_124_3477_n689), .CO(
        DP_OP_422J2_124_3477_n656), .S(DP_OP_422J2_124_3477_n657) );
  FADDX1_HVT DP_OP_422J2_124_3477_U484 ( .A(DP_OP_422J2_124_3477_n691), .B(
        DP_OP_422J2_124_3477_n854), .CI(DP_OP_422J2_124_3477_n685), .CO(
        DP_OP_422J2_124_3477_n654), .S(DP_OP_422J2_124_3477_n655) );
  FADDX1_HVT DP_OP_422J2_124_3477_U483 ( .A(DP_OP_422J2_124_3477_n687), .B(
        DP_OP_422J2_124_3477_n695), .CI(DP_OP_422J2_124_3477_n681), .CO(
        DP_OP_422J2_124_3477_n652), .S(DP_OP_422J2_124_3477_n653) );
  FADDX1_HVT DP_OP_422J2_124_3477_U482 ( .A(DP_OP_422J2_124_3477_n683), .B(
        DP_OP_422J2_124_3477_n852), .CI(DP_OP_422J2_124_3477_n850), .CO(
        DP_OP_422J2_124_3477_n650), .S(DP_OP_422J2_124_3477_n651) );
  FADDX1_HVT DP_OP_422J2_124_3477_U481 ( .A(DP_OP_422J2_124_3477_n848), .B(
        DP_OP_422J2_124_3477_n846), .CI(DP_OP_422J2_124_3477_n679), .CO(
        DP_OP_422J2_124_3477_n648), .S(DP_OP_422J2_124_3477_n649) );
  FADDX1_HVT DP_OP_422J2_124_3477_U480 ( .A(DP_OP_422J2_124_3477_n844), .B(
        DP_OP_422J2_124_3477_n842), .CI(DP_OP_422J2_124_3477_n840), .CO(
        DP_OP_422J2_124_3477_n646), .S(DP_OP_422J2_124_3477_n647) );
  FADDX1_HVT DP_OP_422J2_124_3477_U479 ( .A(DP_OP_422J2_124_3477_n838), .B(
        DP_OP_422J2_124_3477_n673), .CI(DP_OP_422J2_124_3477_n832), .CO(
        DP_OP_422J2_124_3477_n644), .S(DP_OP_422J2_124_3477_n645) );
  FADDX1_HVT DP_OP_422J2_124_3477_U478 ( .A(DP_OP_422J2_124_3477_n836), .B(
        DP_OP_422J2_124_3477_n675), .CI(DP_OP_422J2_124_3477_n677), .CO(
        DP_OP_422J2_124_3477_n642), .S(DP_OP_422J2_124_3477_n643) );
  FADDX1_HVT DP_OP_422J2_124_3477_U477 ( .A(DP_OP_422J2_124_3477_n834), .B(
        DP_OP_422J2_124_3477_n671), .CI(DP_OP_422J2_124_3477_n667), .CO(
        DP_OP_422J2_124_3477_n640), .S(DP_OP_422J2_124_3477_n641) );
  FADDX1_HVT DP_OP_422J2_124_3477_U476 ( .A(DP_OP_422J2_124_3477_n830), .B(
        DP_OP_422J2_124_3477_n669), .CI(DP_OP_422J2_124_3477_n665), .CO(
        DP_OP_422J2_124_3477_n638), .S(DP_OP_422J2_124_3477_n639) );
  FADDX1_HVT DP_OP_422J2_124_3477_U475 ( .A(DP_OP_422J2_124_3477_n828), .B(
        DP_OP_422J2_124_3477_n826), .CI(DP_OP_422J2_124_3477_n661), .CO(
        DP_OP_422J2_124_3477_n636), .S(DP_OP_422J2_124_3477_n637) );
  FADDX1_HVT DP_OP_422J2_124_3477_U474 ( .A(DP_OP_422J2_124_3477_n659), .B(
        DP_OP_422J2_124_3477_n663), .CI(DP_OP_422J2_124_3477_n824), .CO(
        DP_OP_422J2_124_3477_n634), .S(DP_OP_422J2_124_3477_n635) );
  FADDX1_HVT DP_OP_422J2_124_3477_U473 ( .A(DP_OP_422J2_124_3477_n657), .B(
        DP_OP_422J2_124_3477_n822), .CI(DP_OP_422J2_124_3477_n653), .CO(
        DP_OP_422J2_124_3477_n632), .S(DP_OP_422J2_124_3477_n633) );
  FADDX1_HVT DP_OP_422J2_124_3477_U472 ( .A(DP_OP_422J2_124_3477_n655), .B(
        DP_OP_422J2_124_3477_n820), .CI(DP_OP_422J2_124_3477_n651), .CO(
        DP_OP_422J2_124_3477_n630), .S(DP_OP_422J2_124_3477_n631) );
  FADDX1_HVT DP_OP_422J2_124_3477_U471 ( .A(DP_OP_422J2_124_3477_n818), .B(
        DP_OP_422J2_124_3477_n816), .CI(DP_OP_422J2_124_3477_n649), .CO(
        DP_OP_422J2_124_3477_n628), .S(DP_OP_422J2_124_3477_n629) );
  FADDX1_HVT DP_OP_422J2_124_3477_U470 ( .A(DP_OP_422J2_124_3477_n814), .B(
        DP_OP_422J2_124_3477_n812), .CI(DP_OP_422J2_124_3477_n647), .CO(
        DP_OP_422J2_124_3477_n626), .S(DP_OP_422J2_124_3477_n627) );
  FADDX1_HVT DP_OP_422J2_124_3477_U469 ( .A(DP_OP_422J2_124_3477_n810), .B(
        DP_OP_422J2_124_3477_n643), .CI(DP_OP_422J2_124_3477_n806), .CO(
        DP_OP_422J2_124_3477_n624), .S(DP_OP_422J2_124_3477_n625) );
  FADDX1_HVT DP_OP_422J2_124_3477_U468 ( .A(DP_OP_422J2_124_3477_n808), .B(
        DP_OP_422J2_124_3477_n645), .CI(DP_OP_422J2_124_3477_n641), .CO(
        DP_OP_422J2_124_3477_n622), .S(DP_OP_422J2_124_3477_n623) );
  FADDX1_HVT DP_OP_422J2_124_3477_U467 ( .A(DP_OP_422J2_124_3477_n639), .B(
        DP_OP_422J2_124_3477_n804), .CI(DP_OP_422J2_124_3477_n637), .CO(
        DP_OP_422J2_124_3477_n620), .S(DP_OP_422J2_124_3477_n621) );
  FADDX1_HVT DP_OP_422J2_124_3477_U466 ( .A(DP_OP_422J2_124_3477_n635), .B(
        DP_OP_422J2_124_3477_n802), .CI(DP_OP_422J2_124_3477_n633), .CO(
        DP_OP_422J2_124_3477_n618), .S(DP_OP_422J2_124_3477_n619) );
  FADDX1_HVT DP_OP_422J2_124_3477_U465 ( .A(DP_OP_422J2_124_3477_n800), .B(
        DP_OP_422J2_124_3477_n631), .CI(DP_OP_422J2_124_3477_n798), .CO(
        DP_OP_422J2_124_3477_n616), .S(DP_OP_422J2_124_3477_n617) );
  FADDX1_HVT DP_OP_422J2_124_3477_U464 ( .A(DP_OP_422J2_124_3477_n796), .B(
        DP_OP_422J2_124_3477_n629), .CI(DP_OP_422J2_124_3477_n794), .CO(
        DP_OP_422J2_124_3477_n614), .S(DP_OP_422J2_124_3477_n615) );
  FADDX1_HVT DP_OP_422J2_124_3477_U463 ( .A(DP_OP_422J2_124_3477_n627), .B(
        DP_OP_422J2_124_3477_n792), .CI(DP_OP_422J2_124_3477_n625), .CO(
        DP_OP_422J2_124_3477_n612), .S(DP_OP_422J2_124_3477_n613) );
  FADDX1_HVT DP_OP_422J2_124_3477_U462 ( .A(DP_OP_422J2_124_3477_n623), .B(
        DP_OP_422J2_124_3477_n790), .CI(DP_OP_422J2_124_3477_n621), .CO(
        DP_OP_422J2_124_3477_n610), .S(DP_OP_422J2_124_3477_n611) );
  FADDX1_HVT DP_OP_422J2_124_3477_U461 ( .A(DP_OP_422J2_124_3477_n788), .B(
        DP_OP_422J2_124_3477_n619), .CI(DP_OP_422J2_124_3477_n786), .CO(
        DP_OP_422J2_124_3477_n608), .S(DP_OP_422J2_124_3477_n609) );
  FADDX1_HVT DP_OP_422J2_124_3477_U460 ( .A(DP_OP_422J2_124_3477_n617), .B(
        DP_OP_422J2_124_3477_n784), .CI(DP_OP_422J2_124_3477_n615), .CO(
        DP_OP_422J2_124_3477_n606), .S(DP_OP_422J2_124_3477_n607) );
  FADDX1_HVT DP_OP_422J2_124_3477_U459 ( .A(DP_OP_422J2_124_3477_n782), .B(
        DP_OP_422J2_124_3477_n613), .CI(DP_OP_422J2_124_3477_n611), .CO(
        DP_OP_422J2_124_3477_n604), .S(DP_OP_422J2_124_3477_n605) );
  FADDX1_HVT DP_OP_422J2_124_3477_U458 ( .A(DP_OP_422J2_124_3477_n780), .B(
        DP_OP_422J2_124_3477_n609), .CI(DP_OP_422J2_124_3477_n778), .CO(
        DP_OP_422J2_124_3477_n602), .S(DP_OP_422J2_124_3477_n603) );
  FADDX1_HVT DP_OP_422J2_124_3477_U457 ( .A(DP_OP_422J2_124_3477_n607), .B(
        DP_OP_422J2_124_3477_n776), .CI(DP_OP_422J2_124_3477_n605), .CO(
        DP_OP_422J2_124_3477_n600), .S(DP_OP_422J2_124_3477_n601) );
  FADDX1_HVT DP_OP_422J2_124_3477_U456 ( .A(DP_OP_422J2_124_3477_n774), .B(
        DP_OP_422J2_124_3477_n603), .CI(DP_OP_422J2_124_3477_n601), .CO(
        DP_OP_422J2_124_3477_n598), .S(DP_OP_422J2_124_3477_n599) );
  FADDX1_HVT DP_OP_422J2_124_3477_U455 ( .A(DP_OP_422J2_124_3477_n2977), .B(
        DP_OP_422J2_124_3477_n1921), .CI(DP_OP_422J2_124_3477_n1877), .CO(
        DP_OP_422J2_124_3477_n596), .S(DP_OP_422J2_124_3477_n597) );
  FADDX1_HVT DP_OP_422J2_124_3477_U454 ( .A(DP_OP_422J2_124_3477_n770), .B(
        DP_OP_422J2_124_3477_n2236), .CI(DP_OP_422J2_124_3477_n1928), .CO(
        DP_OP_422J2_124_3477_n594), .S(DP_OP_422J2_124_3477_n595) );
  FADDX1_HVT DP_OP_422J2_124_3477_U453 ( .A(DP_OP_422J2_124_3477_n2317), .B(
        DP_OP_422J2_124_3477_n2982), .CI(DP_OP_422J2_124_3477_n2632), .CO(
        DP_OP_422J2_124_3477_n592), .S(DP_OP_422J2_124_3477_n593) );
  FADDX1_HVT DP_OP_422J2_124_3477_U452 ( .A(DP_OP_422J2_124_3477_n2009), .B(
        DP_OP_422J2_124_3477_n2544), .CI(DP_OP_422J2_124_3477_n2764), .CO(
        DP_OP_422J2_124_3477_n590), .S(DP_OP_422J2_124_3477_n591) );
  FADDX1_HVT DP_OP_422J2_124_3477_U451 ( .A(DP_OP_422J2_124_3477_n2229), .B(
        DP_OP_422J2_124_3477_n2324), .CI(DP_OP_422J2_124_3477_n2940), .CO(
        DP_OP_422J2_124_3477_n588), .S(DP_OP_422J2_124_3477_n589) );
  FADDX1_HVT DP_OP_422J2_124_3477_U450 ( .A(DP_OP_422J2_124_3477_n1965), .B(
        DP_OP_422J2_124_3477_n2852), .CI(DP_OP_422J2_124_3477_n2016), .CO(
        DP_OP_422J2_124_3477_n586), .S(DP_OP_422J2_124_3477_n587) );
  FADDX1_HVT DP_OP_422J2_124_3477_U449 ( .A(DP_OP_422J2_124_3477_n2097), .B(
        DP_OP_422J2_124_3477_n1972), .CI(DP_OP_422J2_124_3477_n2808), .CO(
        DP_OP_422J2_124_3477_n584), .S(DP_OP_422J2_124_3477_n585) );
  FADDX1_HVT DP_OP_422J2_124_3477_U448 ( .A(DP_OP_422J2_124_3477_n2933), .B(
        DP_OP_422J2_124_3477_n2368), .CI(DP_OP_422J2_124_3477_n2456), .CO(
        DP_OP_422J2_124_3477_n582), .S(DP_OP_422J2_124_3477_n583) );
  FADDX1_HVT DP_OP_422J2_124_3477_U447 ( .A(DP_OP_422J2_124_3477_n2449), .B(
        DP_OP_422J2_124_3477_n2500), .CI(DP_OP_422J2_124_3477_n2896), .CO(
        DP_OP_422J2_124_3477_n580), .S(DP_OP_422J2_124_3477_n581) );
  FADDX1_HVT DP_OP_422J2_124_3477_U446 ( .A(DP_OP_422J2_124_3477_n2713), .B(
        DP_OP_422J2_124_3477_n2192), .CI(DP_OP_422J2_124_3477_n2720), .CO(
        DP_OP_422J2_124_3477_n578), .S(DP_OP_422J2_124_3477_n579) );
  FADDX1_HVT DP_OP_422J2_124_3477_U445 ( .A(DP_OP_422J2_124_3477_n2889), .B(
        DP_OP_422J2_124_3477_n2412), .CI(DP_OP_422J2_124_3477_n2588), .CO(
        DP_OP_422J2_124_3477_n576), .S(DP_OP_422J2_124_3477_n577) );
  FADDX1_HVT DP_OP_422J2_124_3477_U444 ( .A(DP_OP_422J2_124_3477_n2185), .B(
        DP_OP_422J2_124_3477_n2060), .CI(DP_OP_422J2_124_3477_n2676), .CO(
        DP_OP_422J2_124_3477_n574), .S(DP_OP_422J2_124_3477_n575) );
  FADDX1_HVT DP_OP_422J2_124_3477_U443 ( .A(DP_OP_422J2_124_3477_n2141), .B(
        DP_OP_422J2_124_3477_n2280), .CI(DP_OP_422J2_124_3477_n2148), .CO(
        DP_OP_422J2_124_3477_n572), .S(DP_OP_422J2_124_3477_n573) );
  FADDX1_HVT DP_OP_422J2_124_3477_U442 ( .A(DP_OP_422J2_124_3477_n2537), .B(
        DP_OP_422J2_124_3477_n2361), .CI(DP_OP_422J2_124_3477_n2104), .CO(
        DP_OP_422J2_124_3477_n570), .S(DP_OP_422J2_124_3477_n571) );
  FADDX1_HVT DP_OP_422J2_124_3477_U441 ( .A(DP_OP_422J2_124_3477_n2845), .B(
        DP_OP_422J2_124_3477_n2053), .CI(DP_OP_422J2_124_3477_n2273), .CO(
        DP_OP_422J2_124_3477_n568), .S(DP_OP_422J2_124_3477_n569) );
  FADDX1_HVT DP_OP_422J2_124_3477_U440 ( .A(DP_OP_422J2_124_3477_n2801), .B(
        DP_OP_422J2_124_3477_n2405), .CI(DP_OP_422J2_124_3477_n2493), .CO(
        DP_OP_422J2_124_3477_n566), .S(DP_OP_422J2_124_3477_n567) );
  FADDX1_HVT DP_OP_422J2_124_3477_U439 ( .A(DP_OP_422J2_124_3477_n2757), .B(
        DP_OP_422J2_124_3477_n2581), .CI(DP_OP_422J2_124_3477_n2625), .CO(
        DP_OP_422J2_124_3477_n564), .S(DP_OP_422J2_124_3477_n565) );
  FADDX1_HVT DP_OP_422J2_124_3477_U438 ( .A(DP_OP_422J2_124_3477_n2669), .B(
        DP_OP_422J2_124_3477_n768), .CI(DP_OP_422J2_124_3477_n766), .CO(
        DP_OP_422J2_124_3477_n562), .S(DP_OP_422J2_124_3477_n563) );
  FADDX1_HVT DP_OP_422J2_124_3477_U437 ( .A(DP_OP_422J2_124_3477_n764), .B(
        DP_OP_422J2_124_3477_n736), .CI(DP_OP_422J2_124_3477_n738), .CO(
        DP_OP_422J2_124_3477_n560), .S(DP_OP_422J2_124_3477_n561) );
  FADDX1_HVT DP_OP_422J2_124_3477_U436 ( .A(DP_OP_422J2_124_3477_n762), .B(
        DP_OP_422J2_124_3477_n740), .CI(DP_OP_422J2_124_3477_n742), .CO(
        DP_OP_422J2_124_3477_n558), .S(DP_OP_422J2_124_3477_n559) );
  FADDX1_HVT DP_OP_422J2_124_3477_U435 ( .A(DP_OP_422J2_124_3477_n760), .B(
        DP_OP_422J2_124_3477_n744), .CI(DP_OP_422J2_124_3477_n746), .CO(
        DP_OP_422J2_124_3477_n556), .S(DP_OP_422J2_124_3477_n557) );
  FADDX1_HVT DP_OP_422J2_124_3477_U434 ( .A(DP_OP_422J2_124_3477_n758), .B(
        DP_OP_422J2_124_3477_n748), .CI(DP_OP_422J2_124_3477_n750), .CO(
        DP_OP_422J2_124_3477_n554), .S(DP_OP_422J2_124_3477_n555) );
  FADDX1_HVT DP_OP_422J2_124_3477_U433 ( .A(DP_OP_422J2_124_3477_n756), .B(
        DP_OP_422J2_124_3477_n752), .CI(DP_OP_422J2_124_3477_n754), .CO(
        DP_OP_422J2_124_3477_n552), .S(DP_OP_422J2_124_3477_n553) );
  FADDX1_HVT DP_OP_422J2_124_3477_U432 ( .A(DP_OP_422J2_124_3477_n734), .B(
        DP_OP_422J2_124_3477_n720), .CI(DP_OP_422J2_124_3477_n732), .CO(
        DP_OP_422J2_124_3477_n550), .S(DP_OP_422J2_124_3477_n551) );
  FADDX1_HVT DP_OP_422J2_124_3477_U431 ( .A(DP_OP_422J2_124_3477_n726), .B(
        DP_OP_422J2_124_3477_n722), .CI(DP_OP_422J2_124_3477_n724), .CO(
        DP_OP_422J2_124_3477_n548), .S(DP_OP_422J2_124_3477_n549) );
  FADDX1_HVT DP_OP_422J2_124_3477_U430 ( .A(DP_OP_422J2_124_3477_n730), .B(
        DP_OP_422J2_124_3477_n728), .CI(DP_OP_422J2_124_3477_n595), .CO(
        DP_OP_422J2_124_3477_n546), .S(DP_OP_422J2_124_3477_n547) );
  FADDX1_HVT DP_OP_422J2_124_3477_U429 ( .A(DP_OP_422J2_124_3477_n597), .B(
        DP_OP_422J2_124_3477_n583), .CI(DP_OP_422J2_124_3477_n589), .CO(
        DP_OP_422J2_124_3477_n544), .S(DP_OP_422J2_124_3477_n545) );
  FADDX1_HVT DP_OP_422J2_124_3477_U428 ( .A(DP_OP_422J2_124_3477_n565), .B(
        DP_OP_422J2_124_3477_n587), .CI(DP_OP_422J2_124_3477_n585), .CO(
        DP_OP_422J2_124_3477_n542), .S(DP_OP_422J2_124_3477_n543) );
  FADDX1_HVT DP_OP_422J2_124_3477_U427 ( .A(DP_OP_422J2_124_3477_n591), .B(
        DP_OP_422J2_124_3477_n573), .CI(DP_OP_422J2_124_3477_n575), .CO(
        DP_OP_422J2_124_3477_n540), .S(DP_OP_422J2_124_3477_n541) );
  FADDX1_HVT DP_OP_422J2_124_3477_U426 ( .A(DP_OP_422J2_124_3477_n577), .B(
        DP_OP_422J2_124_3477_n567), .CI(DP_OP_422J2_124_3477_n569), .CO(
        DP_OP_422J2_124_3477_n538), .S(DP_OP_422J2_124_3477_n539) );
  FADDX1_HVT DP_OP_422J2_124_3477_U425 ( .A(DP_OP_422J2_124_3477_n571), .B(
        DP_OP_422J2_124_3477_n593), .CI(DP_OP_422J2_124_3477_n581), .CO(
        DP_OP_422J2_124_3477_n536), .S(DP_OP_422J2_124_3477_n537) );
  FADDX1_HVT DP_OP_422J2_124_3477_U424 ( .A(DP_OP_422J2_124_3477_n579), .B(
        DP_OP_422J2_124_3477_n718), .CI(DP_OP_422J2_124_3477_n716), .CO(
        DP_OP_422J2_124_3477_n534), .S(DP_OP_422J2_124_3477_n535) );
  FADDX1_HVT DP_OP_422J2_124_3477_U423 ( .A(DP_OP_422J2_124_3477_n714), .B(
        DP_OP_422J2_124_3477_n708), .CI(DP_OP_422J2_124_3477_n710), .CO(
        DP_OP_422J2_124_3477_n532), .S(DP_OP_422J2_124_3477_n533) );
  FADDX1_HVT DP_OP_422J2_124_3477_U422 ( .A(DP_OP_422J2_124_3477_n712), .B(
        DP_OP_422J2_124_3477_n706), .CI(DP_OP_422J2_124_3477_n704), .CO(
        DP_OP_422J2_124_3477_n530), .S(DP_OP_422J2_124_3477_n531) );
  FADDX1_HVT DP_OP_422J2_124_3477_U421 ( .A(DP_OP_422J2_124_3477_n702), .B(
        DP_OP_422J2_124_3477_n698), .CI(DP_OP_422J2_124_3477_n696), .CO(
        DP_OP_422J2_124_3477_n528), .S(DP_OP_422J2_124_3477_n529) );
  FADDX1_HVT DP_OP_422J2_124_3477_U420 ( .A(DP_OP_422J2_124_3477_n700), .B(
        DP_OP_422J2_124_3477_n563), .CI(DP_OP_422J2_124_3477_n557), .CO(
        DP_OP_422J2_124_3477_n526), .S(DP_OP_422J2_124_3477_n527) );
  FADDX1_HVT DP_OP_422J2_124_3477_U419 ( .A(DP_OP_422J2_124_3477_n559), .B(
        DP_OP_422J2_124_3477_n553), .CI(DP_OP_422J2_124_3477_n684), .CO(
        DP_OP_422J2_124_3477_n524), .S(DP_OP_422J2_124_3477_n525) );
  FADDX1_HVT DP_OP_422J2_124_3477_U418 ( .A(DP_OP_422J2_124_3477_n694), .B(
        DP_OP_422J2_124_3477_n561), .CI(DP_OP_422J2_124_3477_n555), .CO(
        DP_OP_422J2_124_3477_n522), .S(DP_OP_422J2_124_3477_n523) );
  FADDX1_HVT DP_OP_422J2_124_3477_U417 ( .A(DP_OP_422J2_124_3477_n688), .B(
        DP_OP_422J2_124_3477_n692), .CI(DP_OP_422J2_124_3477_n686), .CO(
        DP_OP_422J2_124_3477_n520), .S(DP_OP_422J2_124_3477_n521) );
  FADDX1_HVT DP_OP_422J2_124_3477_U416 ( .A(DP_OP_422J2_124_3477_n690), .B(
        DP_OP_422J2_124_3477_n682), .CI(DP_OP_422J2_124_3477_n680), .CO(
        DP_OP_422J2_124_3477_n518), .S(DP_OP_422J2_124_3477_n519) );
  FADDX1_HVT DP_OP_422J2_124_3477_U415 ( .A(DP_OP_422J2_124_3477_n549), .B(
        DP_OP_422J2_124_3477_n551), .CI(DP_OP_422J2_124_3477_n547), .CO(
        DP_OP_422J2_124_3477_n516), .S(DP_OP_422J2_124_3477_n517) );
  FADDX1_HVT DP_OP_422J2_124_3477_U414 ( .A(DP_OP_422J2_124_3477_n545), .B(
        DP_OP_422J2_124_3477_n539), .CI(DP_OP_422J2_124_3477_n543), .CO(
        DP_OP_422J2_124_3477_n514), .S(DP_OP_422J2_124_3477_n515) );
  FADDX1_HVT DP_OP_422J2_124_3477_U413 ( .A(DP_OP_422J2_124_3477_n537), .B(
        DP_OP_422J2_124_3477_n541), .CI(DP_OP_422J2_124_3477_n678), .CO(
        DP_OP_422J2_124_3477_n512), .S(DP_OP_422J2_124_3477_n513) );
  FADDX1_HVT DP_OP_422J2_124_3477_U412 ( .A(DP_OP_422J2_124_3477_n676), .B(
        DP_OP_422J2_124_3477_n672), .CI(DP_OP_422J2_124_3477_n535), .CO(
        DP_OP_422J2_124_3477_n510), .S(DP_OP_422J2_124_3477_n511) );
  FADDX1_HVT DP_OP_422J2_124_3477_U411 ( .A(DP_OP_422J2_124_3477_n674), .B(
        DP_OP_422J2_124_3477_n670), .CI(DP_OP_422J2_124_3477_n668), .CO(
        DP_OP_422J2_124_3477_n508), .S(DP_OP_422J2_124_3477_n509) );
  FADDX1_HVT DP_OP_422J2_124_3477_U410 ( .A(DP_OP_422J2_124_3477_n666), .B(
        DP_OP_422J2_124_3477_n533), .CI(DP_OP_422J2_124_3477_n531), .CO(
        DP_OP_422J2_124_3477_n506), .S(DP_OP_422J2_124_3477_n507) );
  FADDX1_HVT DP_OP_422J2_124_3477_U409 ( .A(DP_OP_422J2_124_3477_n664), .B(
        DP_OP_422J2_124_3477_n662), .CI(DP_OP_422J2_124_3477_n660), .CO(
        DP_OP_422J2_124_3477_n504), .S(DP_OP_422J2_124_3477_n505) );
  FADDX1_HVT DP_OP_422J2_124_3477_U408 ( .A(DP_OP_422J2_124_3477_n658), .B(
        DP_OP_422J2_124_3477_n529), .CI(DP_OP_422J2_124_3477_n656), .CO(
        DP_OP_422J2_124_3477_n502), .S(DP_OP_422J2_124_3477_n503) );
  FADDX1_HVT DP_OP_422J2_124_3477_U407 ( .A(DP_OP_422J2_124_3477_n527), .B(
        DP_OP_422J2_124_3477_n654), .CI(DP_OP_422J2_124_3477_n525), .CO(
        DP_OP_422J2_124_3477_n500), .S(DP_OP_422J2_124_3477_n501) );
  FADDX1_HVT DP_OP_422J2_124_3477_U406 ( .A(DP_OP_422J2_124_3477_n652), .B(
        DP_OP_422J2_124_3477_n521), .CI(DP_OP_422J2_124_3477_n519), .CO(
        DP_OP_422J2_124_3477_n498), .S(DP_OP_422J2_124_3477_n499) );
  FADDX1_HVT DP_OP_422J2_124_3477_U405 ( .A(DP_OP_422J2_124_3477_n523), .B(
        DP_OP_422J2_124_3477_n517), .CI(DP_OP_422J2_124_3477_n650), .CO(
        DP_OP_422J2_124_3477_n496), .S(DP_OP_422J2_124_3477_n497) );
  FADDX1_HVT DP_OP_422J2_124_3477_U404 ( .A(DP_OP_422J2_124_3477_n515), .B(
        DP_OP_422J2_124_3477_n648), .CI(DP_OP_422J2_124_3477_n513), .CO(
        DP_OP_422J2_124_3477_n494), .S(DP_OP_422J2_124_3477_n495) );
  FADDX1_HVT DP_OP_422J2_124_3477_U403 ( .A(DP_OP_422J2_124_3477_n646), .B(
        DP_OP_422J2_124_3477_n644), .CI(DP_OP_422J2_124_3477_n642), .CO(
        DP_OP_422J2_124_3477_n492), .S(DP_OP_422J2_124_3477_n493) );
  FADDX1_HVT DP_OP_422J2_124_3477_U402 ( .A(DP_OP_422J2_124_3477_n511), .B(
        DP_OP_422J2_124_3477_n640), .CI(DP_OP_422J2_124_3477_n509), .CO(
        DP_OP_422J2_124_3477_n490), .S(DP_OP_422J2_124_3477_n491) );
  FADDX1_HVT DP_OP_422J2_124_3477_U401 ( .A(DP_OP_422J2_124_3477_n638), .B(
        DP_OP_422J2_124_3477_n507), .CI(DP_OP_422J2_124_3477_n505), .CO(
        DP_OP_422J2_124_3477_n488), .S(DP_OP_422J2_124_3477_n489) );
  FADDX1_HVT DP_OP_422J2_124_3477_U400 ( .A(DP_OP_422J2_124_3477_n636), .B(
        DP_OP_422J2_124_3477_n634), .CI(DP_OP_422J2_124_3477_n503), .CO(
        DP_OP_422J2_124_3477_n486), .S(DP_OP_422J2_124_3477_n487) );
  FADDX1_HVT DP_OP_422J2_124_3477_U399 ( .A(DP_OP_422J2_124_3477_n632), .B(
        DP_OP_422J2_124_3477_n501), .CI(DP_OP_422J2_124_3477_n499), .CO(
        DP_OP_422J2_124_3477_n484), .S(DP_OP_422J2_124_3477_n485) );
  FADDX1_HVT DP_OP_422J2_124_3477_U398 ( .A(DP_OP_422J2_124_3477_n630), .B(
        DP_OP_422J2_124_3477_n497), .CI(DP_OP_422J2_124_3477_n628), .CO(
        DP_OP_422J2_124_3477_n482), .S(DP_OP_422J2_124_3477_n483) );
  FADDX1_HVT DP_OP_422J2_124_3477_U397 ( .A(DP_OP_422J2_124_3477_n495), .B(
        DP_OP_422J2_124_3477_n626), .CI(DP_OP_422J2_124_3477_n493), .CO(
        DP_OP_422J2_124_3477_n480), .S(DP_OP_422J2_124_3477_n481) );
  FADDX1_HVT DP_OP_422J2_124_3477_U396 ( .A(DP_OP_422J2_124_3477_n624), .B(
        DP_OP_422J2_124_3477_n622), .CI(DP_OP_422J2_124_3477_n491), .CO(
        DP_OP_422J2_124_3477_n478), .S(DP_OP_422J2_124_3477_n479) );
  FADDX1_HVT DP_OP_422J2_124_3477_U395 ( .A(DP_OP_422J2_124_3477_n620), .B(
        DP_OP_422J2_124_3477_n489), .CI(DP_OP_422J2_124_3477_n487), .CO(
        DP_OP_422J2_124_3477_n476), .S(DP_OP_422J2_124_3477_n477) );
  FADDX1_HVT DP_OP_422J2_124_3477_U394 ( .A(DP_OP_422J2_124_3477_n618), .B(
        DP_OP_422J2_124_3477_n485), .CI(DP_OP_422J2_124_3477_n616), .CO(
        DP_OP_422J2_124_3477_n474), .S(DP_OP_422J2_124_3477_n475) );
  FADDX1_HVT DP_OP_422J2_124_3477_U393 ( .A(DP_OP_422J2_124_3477_n483), .B(
        DP_OP_422J2_124_3477_n614), .CI(DP_OP_422J2_124_3477_n481), .CO(
        DP_OP_422J2_124_3477_n472), .S(DP_OP_422J2_124_3477_n473) );
  FADDX1_HVT DP_OP_422J2_124_3477_U392 ( .A(DP_OP_422J2_124_3477_n612), .B(
        DP_OP_422J2_124_3477_n479), .CI(DP_OP_422J2_124_3477_n610), .CO(
        DP_OP_422J2_124_3477_n470), .S(DP_OP_422J2_124_3477_n471) );
  FADDX1_HVT DP_OP_422J2_124_3477_U391 ( .A(DP_OP_422J2_124_3477_n477), .B(
        DP_OP_422J2_124_3477_n608), .CI(DP_OP_422J2_124_3477_n475), .CO(
        DP_OP_422J2_124_3477_n468), .S(DP_OP_422J2_124_3477_n469) );
  FADDX1_HVT DP_OP_422J2_124_3477_U390 ( .A(DP_OP_422J2_124_3477_n606), .B(
        DP_OP_422J2_124_3477_n473), .CI(DP_OP_422J2_124_3477_n604), .CO(
        DP_OP_422J2_124_3477_n466), .S(DP_OP_422J2_124_3477_n467) );
  FADDX1_HVT DP_OP_422J2_124_3477_U389 ( .A(DP_OP_422J2_124_3477_n471), .B(
        DP_OP_422J2_124_3477_n469), .CI(DP_OP_422J2_124_3477_n602), .CO(
        DP_OP_422J2_124_3477_n464), .S(DP_OP_422J2_124_3477_n465) );
  FADDX1_HVT DP_OP_422J2_124_3477_U388 ( .A(DP_OP_422J2_124_3477_n600), .B(
        DP_OP_422J2_124_3477_n467), .CI(DP_OP_422J2_124_3477_n465), .CO(
        DP_OP_422J2_124_3477_n462), .S(DP_OP_422J2_124_3477_n463) );
  FADDX1_HVT DP_OP_422J2_124_3477_U386 ( .A(DP_OP_422J2_124_3477_n2976), .B(
        DP_OP_422J2_124_3477_n1920), .CI(DP_OP_422J2_124_3477_n461), .CO(
        DP_OP_422J2_124_3477_n458), .S(DP_OP_422J2_124_3477_n459) );
  FADDX1_HVT DP_OP_422J2_124_3477_U385 ( .A(DP_OP_422J2_124_3477_n2008), .B(
        DP_OP_422J2_124_3477_n2932), .CI(DP_OP_422J2_124_3477_n2360), .CO(
        DP_OP_422J2_124_3477_n456), .S(DP_OP_422J2_124_3477_n457) );
  FADDX1_HVT DP_OP_422J2_124_3477_U384 ( .A(DP_OP_422J2_124_3477_n2492), .B(
        DP_OP_422J2_124_3477_n2888), .CI(DP_OP_422J2_124_3477_n2844), .CO(
        DP_OP_422J2_124_3477_n454), .S(DP_OP_422J2_124_3477_n455) );
  FADDX1_HVT DP_OP_422J2_124_3477_U383 ( .A(DP_OP_422J2_124_3477_n2316), .B(
        DP_OP_422J2_124_3477_n2800), .CI(DP_OP_422J2_124_3477_n2756), .CO(
        DP_OP_422J2_124_3477_n452), .S(DP_OP_422J2_124_3477_n453) );
  FADDX1_HVT DP_OP_422J2_124_3477_U382 ( .A(DP_OP_422J2_124_3477_n2184), .B(
        DP_OP_422J2_124_3477_n1964), .CI(DP_OP_422J2_124_3477_n2712), .CO(
        DP_OP_422J2_124_3477_n450), .S(DP_OP_422J2_124_3477_n451) );
  FADDX1_HVT DP_OP_422J2_124_3477_U381 ( .A(DP_OP_422J2_124_3477_n2668), .B(
        DP_OP_422J2_124_3477_n2624), .CI(DP_OP_422J2_124_3477_n2580), .CO(
        DP_OP_422J2_124_3477_n448), .S(DP_OP_422J2_124_3477_n449) );
  FADDX1_HVT DP_OP_422J2_124_3477_U380 ( .A(DP_OP_422J2_124_3477_n2228), .B(
        DP_OP_422J2_124_3477_n2052), .CI(DP_OP_422J2_124_3477_n2096), .CO(
        DP_OP_422J2_124_3477_n446), .S(DP_OP_422J2_124_3477_n447) );
  FADDX1_HVT DP_OP_422J2_124_3477_U379 ( .A(DP_OP_422J2_124_3477_n2140), .B(
        DP_OP_422J2_124_3477_n2536), .CI(DP_OP_422J2_124_3477_n2448), .CO(
        DP_OP_422J2_124_3477_n444), .S(DP_OP_422J2_124_3477_n445) );
  FADDX1_HVT DP_OP_422J2_124_3477_U378 ( .A(DP_OP_422J2_124_3477_n2272), .B(
        DP_OP_422J2_124_3477_n2404), .CI(DP_OP_422J2_124_3477_n596), .CO(
        DP_OP_422J2_124_3477_n442), .S(DP_OP_422J2_124_3477_n443) );
  FADDX1_HVT DP_OP_422J2_124_3477_U377 ( .A(DP_OP_422J2_124_3477_n594), .B(
        DP_OP_422J2_124_3477_n564), .CI(DP_OP_422J2_124_3477_n592), .CO(
        DP_OP_422J2_124_3477_n440), .S(DP_OP_422J2_124_3477_n441) );
  FADDX1_HVT DP_OP_422J2_124_3477_U376 ( .A(DP_OP_422J2_124_3477_n590), .B(
        DP_OP_422J2_124_3477_n566), .CI(DP_OP_422J2_124_3477_n568), .CO(
        DP_OP_422J2_124_3477_n438), .S(DP_OP_422J2_124_3477_n439) );
  FADDX1_HVT DP_OP_422J2_124_3477_U375 ( .A(DP_OP_422J2_124_3477_n588), .B(
        DP_OP_422J2_124_3477_n570), .CI(DP_OP_422J2_124_3477_n572), .CO(
        DP_OP_422J2_124_3477_n436), .S(DP_OP_422J2_124_3477_n437) );
  FADDX1_HVT DP_OP_422J2_124_3477_U374 ( .A(DP_OP_422J2_124_3477_n586), .B(
        DP_OP_422J2_124_3477_n574), .CI(DP_OP_422J2_124_3477_n576), .CO(
        DP_OP_422J2_124_3477_n434), .S(DP_OP_422J2_124_3477_n435) );
  FADDX1_HVT DP_OP_422J2_124_3477_U373 ( .A(DP_OP_422J2_124_3477_n584), .B(
        DP_OP_422J2_124_3477_n578), .CI(DP_OP_422J2_124_3477_n580), .CO(
        DP_OP_422J2_124_3477_n432), .S(DP_OP_422J2_124_3477_n433) );
  FADDX1_HVT DP_OP_422J2_124_3477_U372 ( .A(DP_OP_422J2_124_3477_n582), .B(
        DP_OP_422J2_124_3477_n459), .CI(DP_OP_422J2_124_3477_n455), .CO(
        DP_OP_422J2_124_3477_n430), .S(DP_OP_422J2_124_3477_n431) );
  FADDX1_HVT DP_OP_422J2_124_3477_U371 ( .A(DP_OP_422J2_124_3477_n451), .B(
        DP_OP_422J2_124_3477_n445), .CI(DP_OP_422J2_124_3477_n447), .CO(
        DP_OP_422J2_124_3477_n428), .S(DP_OP_422J2_124_3477_n429) );
  FADDX1_HVT DP_OP_422J2_124_3477_U370 ( .A(DP_OP_422J2_124_3477_n449), .B(
        DP_OP_422J2_124_3477_n457), .CI(DP_OP_422J2_124_3477_n453), .CO(
        DP_OP_422J2_124_3477_n426), .S(DP_OP_422J2_124_3477_n427) );
  FADDX1_HVT DP_OP_422J2_124_3477_U369 ( .A(DP_OP_422J2_124_3477_n562), .B(
        DP_OP_422J2_124_3477_n560), .CI(DP_OP_422J2_124_3477_n552), .CO(
        DP_OP_422J2_124_3477_n424), .S(DP_OP_422J2_124_3477_n425) );
  FADDX1_HVT DP_OP_422J2_124_3477_U368 ( .A(DP_OP_422J2_124_3477_n558), .B(
        DP_OP_422J2_124_3477_n554), .CI(DP_OP_422J2_124_3477_n556), .CO(
        DP_OP_422J2_124_3477_n422), .S(DP_OP_422J2_124_3477_n423) );
  FADDX1_HVT DP_OP_422J2_124_3477_U367 ( .A(DP_OP_422J2_124_3477_n550), .B(
        DP_OP_422J2_124_3477_n546), .CI(DP_OP_422J2_124_3477_n443), .CO(
        DP_OP_422J2_124_3477_n420), .S(DP_OP_422J2_124_3477_n421) );
  FADDX1_HVT DP_OP_422J2_124_3477_U366 ( .A(DP_OP_422J2_124_3477_n548), .B(
        DP_OP_422J2_124_3477_n544), .CI(DP_OP_422J2_124_3477_n441), .CO(
        DP_OP_422J2_124_3477_n418), .S(DP_OP_422J2_124_3477_n419) );
  FADDX1_HVT DP_OP_422J2_124_3477_U365 ( .A(DP_OP_422J2_124_3477_n542), .B(
        DP_OP_422J2_124_3477_n435), .CI(DP_OP_422J2_124_3477_n437), .CO(
        DP_OP_422J2_124_3477_n416), .S(DP_OP_422J2_124_3477_n417) );
  FADDX1_HVT DP_OP_422J2_124_3477_U364 ( .A(DP_OP_422J2_124_3477_n540), .B(
        DP_OP_422J2_124_3477_n439), .CI(DP_OP_422J2_124_3477_n433), .CO(
        DP_OP_422J2_124_3477_n414), .S(DP_OP_422J2_124_3477_n415) );
  FADDX1_HVT DP_OP_422J2_124_3477_U363 ( .A(DP_OP_422J2_124_3477_n538), .B(
        DP_OP_422J2_124_3477_n536), .CI(DP_OP_422J2_124_3477_n534), .CO(
        DP_OP_422J2_124_3477_n412), .S(DP_OP_422J2_124_3477_n413) );
  FADDX1_HVT DP_OP_422J2_124_3477_U362 ( .A(DP_OP_422J2_124_3477_n431), .B(
        DP_OP_422J2_124_3477_n427), .CI(DP_OP_422J2_124_3477_n532), .CO(
        DP_OP_422J2_124_3477_n410), .S(DP_OP_422J2_124_3477_n411) );
  FADDX1_HVT DP_OP_422J2_124_3477_U361 ( .A(DP_OP_422J2_124_3477_n429), .B(
        DP_OP_422J2_124_3477_n530), .CI(DP_OP_422J2_124_3477_n528), .CO(
        DP_OP_422J2_124_3477_n408), .S(DP_OP_422J2_124_3477_n409) );
  FADDX1_HVT DP_OP_422J2_124_3477_U360 ( .A(DP_OP_422J2_124_3477_n526), .B(
        DP_OP_422J2_124_3477_n425), .CI(DP_OP_422J2_124_3477_n423), .CO(
        DP_OP_422J2_124_3477_n406), .S(DP_OP_422J2_124_3477_n407) );
  FADDX1_HVT DP_OP_422J2_124_3477_U359 ( .A(DP_OP_422J2_124_3477_n524), .B(
        DP_OP_422J2_124_3477_n520), .CI(DP_OP_422J2_124_3477_n518), .CO(
        DP_OP_422J2_124_3477_n404), .S(DP_OP_422J2_124_3477_n405) );
  FADDX1_HVT DP_OP_422J2_124_3477_U358 ( .A(DP_OP_422J2_124_3477_n522), .B(
        DP_OP_422J2_124_3477_n516), .CI(DP_OP_422J2_124_3477_n421), .CO(
        DP_OP_422J2_124_3477_n402), .S(DP_OP_422J2_124_3477_n403) );
  FADDX1_HVT DP_OP_422J2_124_3477_U357 ( .A(DP_OP_422J2_124_3477_n419), .B(
        DP_OP_422J2_124_3477_n514), .CI(DP_OP_422J2_124_3477_n512), .CO(
        DP_OP_422J2_124_3477_n400), .S(DP_OP_422J2_124_3477_n401) );
  FADDX1_HVT DP_OP_422J2_124_3477_U356 ( .A(DP_OP_422J2_124_3477_n417), .B(
        DP_OP_422J2_124_3477_n415), .CI(DP_OP_422J2_124_3477_n413), .CO(
        DP_OP_422J2_124_3477_n398), .S(DP_OP_422J2_124_3477_n399) );
  FADDX1_HVT DP_OP_422J2_124_3477_U355 ( .A(DP_OP_422J2_124_3477_n510), .B(
        DP_OP_422J2_124_3477_n508), .CI(DP_OP_422J2_124_3477_n411), .CO(
        DP_OP_422J2_124_3477_n396), .S(DP_OP_422J2_124_3477_n397) );
  FADDX1_HVT DP_OP_422J2_124_3477_U354 ( .A(DP_OP_422J2_124_3477_n506), .B(
        DP_OP_422J2_124_3477_n409), .CI(DP_OP_422J2_124_3477_n504), .CO(
        DP_OP_422J2_124_3477_n394), .S(DP_OP_422J2_124_3477_n395) );
  FADDX1_HVT DP_OP_422J2_124_3477_U353 ( .A(DP_OP_422J2_124_3477_n502), .B(
        DP_OP_422J2_124_3477_n407), .CI(DP_OP_422J2_124_3477_n500), .CO(
        DP_OP_422J2_124_3477_n392), .S(DP_OP_422J2_124_3477_n393) );
  FADDX1_HVT DP_OP_422J2_124_3477_U352 ( .A(DP_OP_422J2_124_3477_n498), .B(
        DP_OP_422J2_124_3477_n405), .CI(DP_OP_422J2_124_3477_n403), .CO(
        DP_OP_422J2_124_3477_n390), .S(DP_OP_422J2_124_3477_n391) );
  FADDX1_HVT DP_OP_422J2_124_3477_U351 ( .A(DP_OP_422J2_124_3477_n496), .B(
        DP_OP_422J2_124_3477_n401), .CI(DP_OP_422J2_124_3477_n494), .CO(
        DP_OP_422J2_124_3477_n388), .S(DP_OP_422J2_124_3477_n389) );
  FADDX1_HVT DP_OP_422J2_124_3477_U350 ( .A(DP_OP_422J2_124_3477_n399), .B(
        DP_OP_422J2_124_3477_n492), .CI(DP_OP_422J2_124_3477_n490), .CO(
        DP_OP_422J2_124_3477_n386), .S(DP_OP_422J2_124_3477_n387) );
  FADDX1_HVT DP_OP_422J2_124_3477_U349 ( .A(DP_OP_422J2_124_3477_n397), .B(
        DP_OP_422J2_124_3477_n488), .CI(DP_OP_422J2_124_3477_n395), .CO(
        DP_OP_422J2_124_3477_n384), .S(DP_OP_422J2_124_3477_n385) );
  FADDX1_HVT DP_OP_422J2_124_3477_U348 ( .A(DP_OP_422J2_124_3477_n486), .B(
        DP_OP_422J2_124_3477_n393), .CI(DP_OP_422J2_124_3477_n484), .CO(
        DP_OP_422J2_124_3477_n382), .S(DP_OP_422J2_124_3477_n383) );
  FADDX1_HVT DP_OP_422J2_124_3477_U347 ( .A(DP_OP_422J2_124_3477_n391), .B(
        DP_OP_422J2_124_3477_n482), .CI(DP_OP_422J2_124_3477_n389), .CO(
        DP_OP_422J2_124_3477_n380), .S(DP_OP_422J2_124_3477_n381) );
  FADDX1_HVT DP_OP_422J2_124_3477_U346 ( .A(DP_OP_422J2_124_3477_n480), .B(
        DP_OP_422J2_124_3477_n387), .CI(DP_OP_422J2_124_3477_n478), .CO(
        DP_OP_422J2_124_3477_n378), .S(DP_OP_422J2_124_3477_n379) );
  FADDX1_HVT DP_OP_422J2_124_3477_U345 ( .A(DP_OP_422J2_124_3477_n385), .B(
        DP_OP_422J2_124_3477_n476), .CI(DP_OP_422J2_124_3477_n383), .CO(
        DP_OP_422J2_124_3477_n376), .S(DP_OP_422J2_124_3477_n377) );
  FADDX1_HVT DP_OP_422J2_124_3477_U344 ( .A(DP_OP_422J2_124_3477_n474), .B(
        DP_OP_422J2_124_3477_n381), .CI(DP_OP_422J2_124_3477_n472), .CO(
        DP_OP_422J2_124_3477_n374), .S(DP_OP_422J2_124_3477_n375) );
  FADDX1_HVT DP_OP_422J2_124_3477_U343 ( .A(DP_OP_422J2_124_3477_n379), .B(
        DP_OP_422J2_124_3477_n470), .CI(DP_OP_422J2_124_3477_n377), .CO(
        DP_OP_422J2_124_3477_n372), .S(DP_OP_422J2_124_3477_n373) );
  FADDX1_HVT DP_OP_422J2_124_3477_U342 ( .A(DP_OP_422J2_124_3477_n468), .B(
        DP_OP_422J2_124_3477_n375), .CI(DP_OP_422J2_124_3477_n466), .CO(
        DP_OP_422J2_124_3477_n370), .S(DP_OP_422J2_124_3477_n371) );
  FADDX1_HVT DP_OP_422J2_124_3477_U341 ( .A(DP_OP_422J2_124_3477_n373), .B(
        DP_OP_422J2_124_3477_n464), .CI(DP_OP_422J2_124_3477_n371), .CO(
        DP_OP_422J2_124_3477_n368), .S(DP_OP_422J2_124_3477_n369) );
  FADDX1_HVT DP_OP_422J2_124_3477_U340 ( .A(DP_OP_422J2_124_3477_n1876), .B(
        DP_OP_422J2_124_3477_n460), .CI(DP_OP_422J2_124_3477_n458), .CO(
        DP_OP_422J2_124_3477_n366), .S(DP_OP_422J2_124_3477_n367) );
  FADDX1_HVT DP_OP_422J2_124_3477_U339 ( .A(DP_OP_422J2_124_3477_n448), .B(
        DP_OP_422J2_124_3477_n444), .CI(DP_OP_422J2_124_3477_n456), .CO(
        DP_OP_422J2_124_3477_n364), .S(DP_OP_422J2_124_3477_n365) );
  FADDX1_HVT DP_OP_422J2_124_3477_U338 ( .A(DP_OP_422J2_124_3477_n454), .B(
        DP_OP_422J2_124_3477_n452), .CI(DP_OP_422J2_124_3477_n450), .CO(
        DP_OP_422J2_124_3477_n362), .S(DP_OP_422J2_124_3477_n363) );
  FADDX1_HVT DP_OP_422J2_124_3477_U337 ( .A(DP_OP_422J2_124_3477_n446), .B(
        DP_OP_422J2_124_3477_n442), .CI(DP_OP_422J2_124_3477_n440), .CO(
        DP_OP_422J2_124_3477_n360), .S(DP_OP_422J2_124_3477_n361) );
  FADDX1_HVT DP_OP_422J2_124_3477_U336 ( .A(DP_OP_422J2_124_3477_n438), .B(
        DP_OP_422J2_124_3477_n436), .CI(DP_OP_422J2_124_3477_n434), .CO(
        DP_OP_422J2_124_3477_n358), .S(DP_OP_422J2_124_3477_n359) );
  FADDX1_HVT DP_OP_422J2_124_3477_U335 ( .A(DP_OP_422J2_124_3477_n432), .B(
        DP_OP_422J2_124_3477_n367), .CI(DP_OP_422J2_124_3477_n430), .CO(
        DP_OP_422J2_124_3477_n356), .S(DP_OP_422J2_124_3477_n357) );
  FADDX1_HVT DP_OP_422J2_124_3477_U334 ( .A(DP_OP_422J2_124_3477_n428), .B(
        DP_OP_422J2_124_3477_n363), .CI(DP_OP_422J2_124_3477_n365), .CO(
        DP_OP_422J2_124_3477_n354), .S(DP_OP_422J2_124_3477_n355) );
  FADDX1_HVT DP_OP_422J2_124_3477_U333 ( .A(DP_OP_422J2_124_3477_n426), .B(
        DP_OP_422J2_124_3477_n424), .CI(DP_OP_422J2_124_3477_n422), .CO(
        DP_OP_422J2_124_3477_n352), .S(DP_OP_422J2_124_3477_n353) );
  FADDX1_HVT DP_OP_422J2_124_3477_U332 ( .A(DP_OP_422J2_124_3477_n420), .B(
        DP_OP_422J2_124_3477_n361), .CI(DP_OP_422J2_124_3477_n418), .CO(
        DP_OP_422J2_124_3477_n350), .S(DP_OP_422J2_124_3477_n351) );
  FADDX1_HVT DP_OP_422J2_124_3477_U331 ( .A(DP_OP_422J2_124_3477_n416), .B(
        DP_OP_422J2_124_3477_n359), .CI(DP_OP_422J2_124_3477_n414), .CO(
        DP_OP_422J2_124_3477_n348), .S(DP_OP_422J2_124_3477_n349) );
  FADDX1_HVT DP_OP_422J2_124_3477_U330 ( .A(DP_OP_422J2_124_3477_n412), .B(
        DP_OP_422J2_124_3477_n357), .CI(DP_OP_422J2_124_3477_n410), .CO(
        DP_OP_422J2_124_3477_n346), .S(DP_OP_422J2_124_3477_n347) );
  FADDX1_HVT DP_OP_422J2_124_3477_U329 ( .A(DP_OP_422J2_124_3477_n355), .B(
        DP_OP_422J2_124_3477_n408), .CI(DP_OP_422J2_124_3477_n406), .CO(
        DP_OP_422J2_124_3477_n344), .S(DP_OP_422J2_124_3477_n345) );
  FADDX1_HVT DP_OP_422J2_124_3477_U328 ( .A(DP_OP_422J2_124_3477_n353), .B(
        DP_OP_422J2_124_3477_n404), .CI(DP_OP_422J2_124_3477_n402), .CO(
        DP_OP_422J2_124_3477_n342), .S(DP_OP_422J2_124_3477_n343) );
  FADDX1_HVT DP_OP_422J2_124_3477_U327 ( .A(DP_OP_422J2_124_3477_n351), .B(
        DP_OP_422J2_124_3477_n400), .CI(DP_OP_422J2_124_3477_n349), .CO(
        DP_OP_422J2_124_3477_n340), .S(DP_OP_422J2_124_3477_n341) );
  FADDX1_HVT DP_OP_422J2_124_3477_U326 ( .A(DP_OP_422J2_124_3477_n398), .B(
        DP_OP_422J2_124_3477_n347), .CI(DP_OP_422J2_124_3477_n396), .CO(
        DP_OP_422J2_124_3477_n338), .S(DP_OP_422J2_124_3477_n339) );
  FADDX1_HVT DP_OP_422J2_124_3477_U325 ( .A(DP_OP_422J2_124_3477_n394), .B(
        DP_OP_422J2_124_3477_n345), .CI(DP_OP_422J2_124_3477_n392), .CO(
        DP_OP_422J2_124_3477_n336), .S(DP_OP_422J2_124_3477_n337) );
  FADDX1_HVT DP_OP_422J2_124_3477_U324 ( .A(DP_OP_422J2_124_3477_n343), .B(
        DP_OP_422J2_124_3477_n390), .CI(DP_OP_422J2_124_3477_n388), .CO(
        DP_OP_422J2_124_3477_n334), .S(DP_OP_422J2_124_3477_n335) );
  FADDX1_HVT DP_OP_422J2_124_3477_U323 ( .A(DP_OP_422J2_124_3477_n341), .B(
        DP_OP_422J2_124_3477_n386), .CI(DP_OP_422J2_124_3477_n339), .CO(
        DP_OP_422J2_124_3477_n332), .S(DP_OP_422J2_124_3477_n333) );
  FADDX1_HVT DP_OP_422J2_124_3477_U322 ( .A(DP_OP_422J2_124_3477_n384), .B(
        DP_OP_422J2_124_3477_n337), .CI(DP_OP_422J2_124_3477_n382), .CO(
        DP_OP_422J2_124_3477_n330), .S(DP_OP_422J2_124_3477_n331) );
  FADDX1_HVT DP_OP_422J2_124_3477_U321 ( .A(DP_OP_422J2_124_3477_n380), .B(
        DP_OP_422J2_124_3477_n335), .CI(DP_OP_422J2_124_3477_n333), .CO(
        DP_OP_422J2_124_3477_n328), .S(DP_OP_422J2_124_3477_n329) );
  FADDX1_HVT DP_OP_422J2_124_3477_U320 ( .A(DP_OP_422J2_124_3477_n378), .B(
        DP_OP_422J2_124_3477_n331), .CI(DP_OP_422J2_124_3477_n376), .CO(
        DP_OP_422J2_124_3477_n326), .S(DP_OP_422J2_124_3477_n327) );
  FADDX1_HVT DP_OP_422J2_124_3477_U319 ( .A(DP_OP_422J2_124_3477_n374), .B(
        DP_OP_422J2_124_3477_n329), .CI(DP_OP_422J2_124_3477_n372), .CO(
        DP_OP_422J2_124_3477_n324), .S(DP_OP_422J2_124_3477_n325) );
  FADDX1_HVT DP_OP_422J2_124_3477_U318 ( .A(DP_OP_422J2_124_3477_n327), .B(
        DP_OP_422J2_124_3477_n370), .CI(DP_OP_422J2_124_3477_n325), .CO(
        DP_OP_422J2_124_3477_n322), .S(DP_OP_422J2_124_3477_n323) );
  FADDX1_HVT DP_OP_422J2_124_3477_U317 ( .A(DP_OP_422J2_124_3477_n1875), .B(
        DP_OP_422J2_124_3477_n366), .CI(DP_OP_422J2_124_3477_n364), .CO(
        DP_OP_422J2_124_3477_n320), .S(DP_OP_422J2_124_3477_n321) );
  FADDX1_HVT DP_OP_422J2_124_3477_U316 ( .A(DP_OP_422J2_124_3477_n362), .B(
        DP_OP_422J2_124_3477_n360), .CI(DP_OP_422J2_124_3477_n358), .CO(
        DP_OP_422J2_124_3477_n318), .S(DP_OP_422J2_124_3477_n319) );
  FADDX1_HVT DP_OP_422J2_124_3477_U315 ( .A(DP_OP_422J2_124_3477_n356), .B(
        DP_OP_422J2_124_3477_n321), .CI(DP_OP_422J2_124_3477_n354), .CO(
        DP_OP_422J2_124_3477_n316), .S(DP_OP_422J2_124_3477_n317) );
  FADDX1_HVT DP_OP_422J2_124_3477_U314 ( .A(DP_OP_422J2_124_3477_n352), .B(
        DP_OP_422J2_124_3477_n350), .CI(DP_OP_422J2_124_3477_n319), .CO(
        DP_OP_422J2_124_3477_n314), .S(DP_OP_422J2_124_3477_n315) );
  FADDX1_HVT DP_OP_422J2_124_3477_U313 ( .A(DP_OP_422J2_124_3477_n348), .B(
        DP_OP_422J2_124_3477_n346), .CI(DP_OP_422J2_124_3477_n317), .CO(
        DP_OP_422J2_124_3477_n312), .S(DP_OP_422J2_124_3477_n313) );
  FADDX1_HVT DP_OP_422J2_124_3477_U312 ( .A(DP_OP_422J2_124_3477_n344), .B(
        DP_OP_422J2_124_3477_n342), .CI(DP_OP_422J2_124_3477_n315), .CO(
        DP_OP_422J2_124_3477_n310), .S(DP_OP_422J2_124_3477_n311) );
  FADDX1_HVT DP_OP_422J2_124_3477_U311 ( .A(DP_OP_422J2_124_3477_n340), .B(
        DP_OP_422J2_124_3477_n313), .CI(DP_OP_422J2_124_3477_n338), .CO(
        DP_OP_422J2_124_3477_n308), .S(DP_OP_422J2_124_3477_n309) );
  FADDX1_HVT DP_OP_422J2_124_3477_U310 ( .A(DP_OP_422J2_124_3477_n336), .B(
        DP_OP_422J2_124_3477_n311), .CI(DP_OP_422J2_124_3477_n334), .CO(
        DP_OP_422J2_124_3477_n306), .S(DP_OP_422J2_124_3477_n307) );
  FADDX1_HVT DP_OP_422J2_124_3477_U309 ( .A(DP_OP_422J2_124_3477_n332), .B(
        DP_OP_422J2_124_3477_n309), .CI(DP_OP_422J2_124_3477_n330), .CO(
        DP_OP_422J2_124_3477_n304), .S(DP_OP_422J2_124_3477_n305) );
  FADDX1_HVT DP_OP_422J2_124_3477_U308 ( .A(DP_OP_422J2_124_3477_n307), .B(
        DP_OP_422J2_124_3477_n328), .CI(DP_OP_422J2_124_3477_n305), .CO(
        DP_OP_422J2_124_3477_n302), .S(DP_OP_422J2_124_3477_n303) );
  FADDX1_HVT DP_OP_422J2_124_3477_U307 ( .A(DP_OP_422J2_124_3477_n326), .B(
        DP_OP_422J2_124_3477_n324), .CI(DP_OP_422J2_124_3477_n303), .CO(
        DP_OP_422J2_124_3477_n300), .S(DP_OP_422J2_124_3477_n301) );
  FADDX1_HVT DP_OP_422J2_124_3477_U306 ( .A(DP_OP_422J2_124_3477_n1874), .B(
        DP_OP_422J2_124_3477_n320), .CI(DP_OP_422J2_124_3477_n318), .CO(
        DP_OP_422J2_124_3477_n298), .S(DP_OP_422J2_124_3477_n299) );
  FADDX1_HVT DP_OP_422J2_124_3477_U305 ( .A(DP_OP_422J2_124_3477_n316), .B(
        DP_OP_422J2_124_3477_n299), .CI(DP_OP_422J2_124_3477_n314), .CO(
        DP_OP_422J2_124_3477_n296), .S(DP_OP_422J2_124_3477_n297) );
  FADDX1_HVT DP_OP_422J2_124_3477_U304 ( .A(DP_OP_422J2_124_3477_n312), .B(
        DP_OP_422J2_124_3477_n310), .CI(DP_OP_422J2_124_3477_n297), .CO(
        DP_OP_422J2_124_3477_n294), .S(DP_OP_422J2_124_3477_n295) );
  FADDX1_HVT DP_OP_422J2_124_3477_U303 ( .A(DP_OP_422J2_124_3477_n308), .B(
        DP_OP_422J2_124_3477_n295), .CI(DP_OP_422J2_124_3477_n306), .CO(
        DP_OP_422J2_124_3477_n292), .S(DP_OP_422J2_124_3477_n293) );
  FADDX1_HVT DP_OP_422J2_124_3477_U302 ( .A(DP_OP_422J2_124_3477_n304), .B(
        DP_OP_422J2_124_3477_n293), .CI(DP_OP_422J2_124_3477_n302), .CO(
        DP_OP_422J2_124_3477_n290), .S(DP_OP_422J2_124_3477_n291) );
  FADDX1_HVT DP_OP_422J2_124_3477_U300 ( .A(DP_OP_422J2_124_3477_n289), .B(
        DP_OP_422J2_124_3477_n298), .CI(DP_OP_422J2_124_3477_n296), .CO(
        DP_OP_422J2_124_3477_n286), .S(DP_OP_422J2_124_3477_n287) );
  FADDX1_HVT DP_OP_422J2_124_3477_U299 ( .A(DP_OP_422J2_124_3477_n287), .B(
        DP_OP_422J2_124_3477_n294), .CI(DP_OP_422J2_124_3477_n292), .CO(
        DP_OP_422J2_124_3477_n284), .S(DP_OP_422J2_124_3477_n285) );
  FADDX1_HVT DP_OP_422J2_124_3477_U298 ( .A(DP_OP_422J2_124_3477_n1873), .B(
        DP_OP_422J2_124_3477_n288), .CI(DP_OP_422J2_124_3477_n286), .CO(
        DP_OP_422J2_124_3477_n282), .S(DP_OP_422J2_124_3477_n283) );
  FADDX1_HVT DP_OP_422J2_124_3477_U281 ( .A(DP_OP_422J2_124_3477_n1853), .B(
        DP_OP_422J2_124_3477_n1851), .CI(DP_OP_422J2_124_3477_n1849), .CO(
        DP_OP_422J2_124_3477_n219), .S(n_conv2_sum_a[0]) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U280 ( .A1(DP_OP_422J2_124_3477_n1787), 
        .A2(DP_OP_422J2_124_3477_n1789), .Y(DP_OP_422J2_124_3477_n218) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U279 ( .A1(DP_OP_422J2_124_3477_n1789), .A2(
        DP_OP_422J2_124_3477_n1787), .Y(DP_OP_422J2_124_3477_n217) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U273 ( .A1(DP_OP_422J2_124_3477_n1681), 
        .A2(DP_OP_422J2_124_3477_n1683), .Y(DP_OP_422J2_124_3477_n215) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U265 ( .A1(DP_OP_422J2_124_3477_n1527), 
        .A2(DP_OP_422J2_124_3477_n1529), .Y(DP_OP_422J2_124_3477_n210) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U264 ( .A1(DP_OP_422J2_124_3477_n1529), .A2(
        DP_OP_422J2_124_3477_n1527), .Y(DP_OP_422J2_124_3477_n209) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U259 ( .A1(DP_OP_422J2_124_3477_n1351), 
        .A2(DP_OP_422J2_124_3477_n1353), .Y(DP_OP_422J2_124_3477_n207) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U251 ( .A1(DP_OP_422J2_124_3477_n1163), 
        .A2(DP_OP_422J2_124_3477_n1165), .Y(DP_OP_422J2_124_3477_n202) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U250 ( .A1(DP_OP_422J2_124_3477_n1165), .A2(
        DP_OP_422J2_124_3477_n1163), .Y(DP_OP_422J2_124_3477_n201) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U245 ( .A1(DP_OP_422J2_124_3477_n969), .A2(
        DP_OP_422J2_124_3477_n971), .Y(DP_OP_422J2_124_3477_n199) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U237 ( .A1(DP_OP_422J2_124_3477_n773), .A2(
        DP_OP_422J2_124_3477_n968), .Y(DP_OP_422J2_124_3477_n194) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U236 ( .A1(DP_OP_422J2_124_3477_n968), .A2(
        DP_OP_422J2_124_3477_n773), .Y(DP_OP_422J2_124_3477_n193) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U230 ( .A1(DP_OP_422J2_124_3477_n599), .A2(
        DP_OP_422J2_124_3477_n772), .Y(DP_OP_422J2_124_3477_n190) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U229 ( .A1(DP_OP_422J2_124_3477_n772), .A2(
        DP_OP_422J2_124_3477_n599), .Y(DP_OP_422J2_124_3477_n189) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U224 ( .A1(DP_OP_422J2_124_3477_n463), .A2(
        DP_OP_422J2_124_3477_n598), .Y(DP_OP_422J2_124_3477_n187) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U223 ( .A1(DP_OP_422J2_124_3477_n598), .A2(
        DP_OP_422J2_124_3477_n463), .Y(DP_OP_422J2_124_3477_n186) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U219 ( .A1(DP_OP_422J2_124_3477_n189), .A2(
        DP_OP_422J2_124_3477_n186), .Y(DP_OP_422J2_124_3477_n184) );
  AOI21X1_HVT DP_OP_422J2_124_3477_U218 ( .A1(DP_OP_422J2_124_3477_n184), .A2(
        DP_OP_422J2_124_3477_n192), .A3(DP_OP_422J2_124_3477_n185), .Y(
        DP_OP_422J2_124_3477_n183) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U215 ( .A1(DP_OP_422J2_124_3477_n369), .A2(
        DP_OP_422J2_124_3477_n462), .Y(DP_OP_422J2_124_3477_n181) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U214 ( .A1(DP_OP_422J2_124_3477_n462), .A2(
        DP_OP_422J2_124_3477_n369), .Y(DP_OP_422J2_124_3477_n180) );
  AOI21X1_HVT DP_OP_422J2_124_3477_U209 ( .A1(DP_OP_422J2_124_3477_n182), .A2(
        DP_OP_422J2_124_3477_n241), .A3(DP_OP_422J2_124_3477_n179), .Y(
        DP_OP_422J2_124_3477_n177) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U207 ( .A1(DP_OP_422J2_124_3477_n323), .A2(
        DP_OP_422J2_124_3477_n368), .Y(DP_OP_422J2_124_3477_n176) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U206 ( .A1(DP_OP_422J2_124_3477_n368), .A2(
        DP_OP_422J2_124_3477_n323), .Y(DP_OP_422J2_124_3477_n175) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U204 ( .A1(DP_OP_422J2_124_3477_n240), .A2(
        DP_OP_422J2_124_3477_n176), .Y(DP_OP_422J2_124_3477_n25) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U202 ( .A1(DP_OP_422J2_124_3477_n175), .A2(
        DP_OP_422J2_124_3477_n180), .Y(DP_OP_422J2_124_3477_n173) );
  AOI21X1_HVT DP_OP_422J2_124_3477_U201 ( .A1(DP_OP_422J2_124_3477_n182), .A2(
        DP_OP_422J2_124_3477_n173), .A3(DP_OP_422J2_124_3477_n174), .Y(
        DP_OP_422J2_124_3477_n172) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U199 ( .A1(DP_OP_422J2_124_3477_n301), .A2(
        DP_OP_422J2_124_3477_n322), .Y(DP_OP_422J2_124_3477_n171) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U198 ( .A1(DP_OP_422J2_124_3477_n322), .A2(
        DP_OP_422J2_124_3477_n301), .Y(DP_OP_422J2_124_3477_n170) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U193 ( .A1(DP_OP_422J2_124_3477_n300), .A2(
        DP_OP_422J2_124_3477_n291), .Y(DP_OP_422J2_124_3477_n168) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U192 ( .A1(DP_OP_422J2_124_3477_n291), .A2(
        DP_OP_422J2_124_3477_n300), .Y(DP_OP_422J2_124_3477_n167) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U188 ( .A1(DP_OP_422J2_124_3477_n167), .A2(
        DP_OP_422J2_124_3477_n170), .Y(DP_OP_422J2_124_3477_n165) );
  AOI21X1_HVT DP_OP_422J2_124_3477_U187 ( .A1(DP_OP_422J2_124_3477_n174), .A2(
        DP_OP_422J2_124_3477_n165), .A3(DP_OP_422J2_124_3477_n166), .Y(
        DP_OP_422J2_124_3477_n164) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U186 ( .A1(DP_OP_422J2_124_3477_n173), .A2(
        DP_OP_422J2_124_3477_n165), .Y(DP_OP_422J2_124_3477_n163) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U182 ( .A1(DP_OP_422J2_124_3477_n290), .A2(
        DP_OP_422J2_124_3477_n285), .Y(DP_OP_422J2_124_3477_n152) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U181 ( .A1(DP_OP_422J2_124_3477_n285), .A2(
        DP_OP_422J2_124_3477_n290), .Y(DP_OP_422J2_124_3477_n151) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U179 ( .A1(DP_OP_422J2_124_3477_n237), .A2(
        DP_OP_422J2_124_3477_n152), .Y(DP_OP_422J2_124_3477_n22) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U168 ( .A1(DP_OP_422J2_124_3477_n284), .A2(
        DP_OP_422J2_124_3477_n283), .Y(DP_OP_422J2_124_3477_n149) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U167 ( .A1(DP_OP_422J2_124_3477_n283), .A2(
        DP_OP_422J2_124_3477_n284), .Y(DP_OP_422J2_124_3477_n148) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U165 ( .A1(DP_OP_422J2_124_3477_n236), .A2(
        DP_OP_422J2_124_3477_n149), .Y(DP_OP_422J2_124_3477_n21) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U161 ( .A1(DP_OP_422J2_124_3477_n237), .A2(
        DP_OP_422J2_124_3477_n236), .Y(DP_OP_422J2_124_3477_n144) );
  AOI21X1_HVT DP_OP_422J2_124_3477_U158 ( .A1(DP_OP_422J2_124_3477_n162), .A2(
        DP_OP_422J2_124_3477_n142), .A3(DP_OP_422J2_124_3477_n143), .Y(
        DP_OP_422J2_124_3477_n141) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U156 ( .A1(DP_OP_422J2_124_3477_n282), .A2(
        DP_OP_422J2_124_3477_n281), .Y(DP_OP_422J2_124_3477_n140) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U146 ( .A1(DP_OP_422J2_124_3477_n279), .A2(
        DP_OP_422J2_124_3477_n280), .Y(DP_OP_422J2_124_3477_n133) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U145 ( .A1(DP_OP_422J2_124_3477_n280), .A2(
        DP_OP_422J2_124_3477_n279), .Y(DP_OP_422J2_124_3477_n132) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U140 ( .A1(DP_OP_422J2_124_3477_n277), .A2(
        DP_OP_422J2_124_3477_n278), .Y(DP_OP_422J2_124_3477_n130) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U139 ( .A1(DP_OP_422J2_124_3477_n278), .A2(
        DP_OP_422J2_124_3477_n277), .Y(DP_OP_422J2_124_3477_n129) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U135 ( .A1(DP_OP_422J2_124_3477_n129), .A2(
        DP_OP_422J2_124_3477_n132), .Y(DP_OP_422J2_124_3477_n127) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U130 ( .A1(DP_OP_422J2_124_3477_n275), .A2(
        DP_OP_422J2_124_3477_n276), .Y(DP_OP_422J2_124_3477_n123) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U123 ( .A1(DP_OP_422J2_124_3477_n127), .A2(
        n430), .Y(DP_OP_422J2_124_3477_n118) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U120 ( .A1(DP_OP_422J2_124_3477_n273), .A2(
        DP_OP_422J2_124_3477_n274), .Y(DP_OP_422J2_124_3477_n116) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U119 ( .A1(DP_OP_422J2_124_3477_n274), .A2(
        DP_OP_422J2_124_3477_n273), .Y(DP_OP_422J2_124_3477_n115) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U110 ( .A1(DP_OP_422J2_124_3477_n271), .A2(
        DP_OP_422J2_124_3477_n272), .Y(DP_OP_422J2_124_3477_n109) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U103 ( .A1(DP_OP_422J2_124_3477_n113), .A2(
        n429), .Y(DP_OP_422J2_124_3477_n104) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U100 ( .A1(DP_OP_422J2_124_3477_n269), .A2(
        DP_OP_422J2_124_3477_n270), .Y(DP_OP_422J2_124_3477_n102) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U99 ( .A1(DP_OP_422J2_124_3477_n270), .A2(
        DP_OP_422J2_124_3477_n269), .Y(DP_OP_422J2_124_3477_n101) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U90 ( .A1(DP_OP_422J2_124_3477_n267), .A2(
        DP_OP_422J2_124_3477_n268), .Y(DP_OP_422J2_124_3477_n95) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U83 ( .A1(DP_OP_422J2_124_3477_n99), .A2(
        n425), .Y(DP_OP_422J2_124_3477_n90) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U80 ( .A1(DP_OP_422J2_124_3477_n265), .A2(
        DP_OP_422J2_124_3477_n266), .Y(DP_OP_422J2_124_3477_n88) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U79 ( .A1(DP_OP_422J2_124_3477_n266), .A2(
        DP_OP_422J2_124_3477_n265), .Y(DP_OP_422J2_124_3477_n87) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U70 ( .A1(DP_OP_422J2_124_3477_n263), .A2(
        DP_OP_422J2_124_3477_n264), .Y(DP_OP_422J2_124_3477_n81) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U63 ( .A1(DP_OP_422J2_124_3477_n85), .A2(
        n424), .Y(DP_OP_422J2_124_3477_n76) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U61 ( .A1(DP_OP_422J2_124_3477_n76), .A2(
        DP_OP_422J2_124_3477_n137), .Y(DP_OP_422J2_124_3477_n74) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U56 ( .A1(DP_OP_422J2_124_3477_n261), .A2(
        DP_OP_422J2_124_3477_n262), .Y(DP_OP_422J2_124_3477_n70) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U49 ( .A1(DP_OP_422J2_124_3477_n74), .A2(
        n423), .Y(DP_OP_422J2_124_3477_n65) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U45 ( .A1(DP_OP_422J2_124_3477_n237), .A2(
        DP_OP_422J2_124_3477_n63), .Y(DP_OP_422J2_124_3477_n61) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U42 ( .A1(DP_OP_422J2_124_3477_n259), .A2(
        DP_OP_422J2_124_3477_n260), .Y(DP_OP_422J2_124_3477_n59) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U41 ( .A1(DP_OP_422J2_124_3477_n260), .A2(
        DP_OP_422J2_124_3477_n259), .Y(DP_OP_422J2_124_3477_n58) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U32 ( .A1(DP_OP_422J2_124_3477_n257), .A2(
        DP_OP_422J2_124_3477_n258), .Y(DP_OP_422J2_124_3477_n52) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U25 ( .A1(DP_OP_422J2_124_3477_n56), .A2(
        n422), .Y(DP_OP_422J2_124_3477_n47) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U22 ( .A1(DP_OP_422J2_124_3477_n255), .A2(
        DP_OP_422J2_124_3477_n256), .Y(DP_OP_422J2_124_3477_n45) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U21 ( .A1(DP_OP_422J2_124_3477_n256), .A2(
        DP_OP_422J2_124_3477_n255), .Y(DP_OP_422J2_124_3477_n44) );
  AOI21X1_HVT DP_OP_422J2_124_3477_U16 ( .A1(DP_OP_422J2_124_3477_n162), .A2(
        DP_OP_422J2_124_3477_n42), .A3(DP_OP_422J2_124_3477_n43), .Y(
        DP_OP_422J2_124_3477_n41) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U14 ( .A1(DP_OP_422J2_124_3477_n253), .A2(
        DP_OP_422J2_124_3477_n254), .Y(DP_OP_422J2_124_3477_n40) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U13 ( .A1(DP_OP_422J2_124_3477_n254), .A2(
        DP_OP_422J2_124_3477_n253), .Y(DP_OP_422J2_124_3477_n39) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U8 ( .A1(n421), .A2(
        DP_OP_422J2_124_3477_n252), .Y(DP_OP_422J2_124_3477_n37) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1969 ( .A1(DP_OP_425J2_127_3477_n2218), 
        .A2(DP_OP_423J2_125_3477_n2754), .Y(DP_OP_424J2_126_3477_n2730) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1441 ( .A1(DP_OP_424J2_126_3477_n2218), 
        .A2(DP_OP_424J2_126_3477_n2226), .Y(DP_OP_424J2_126_3477_n2202) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1803 ( .A1(DP_OP_424J2_126_3477_n2572), 
        .A2(DP_OP_422J2_124_3477_n2579), .Y(DP_OP_424J2_126_3477_n2564) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1187 ( .A1(DP_OP_424J2_126_3477_n2044), 
        .A2(DP_OP_423J2_125_3477_n1963), .Y(DP_OP_423J2_125_3477_n1948) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1529 ( .A1(DP_OP_422J2_124_3477_n2746), 
        .A2(DP_OP_424J2_126_3477_n2314), .Y(DP_OP_424J2_126_3477_n2290) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1534 ( .A1(DP_OP_422J2_124_3477_n2311), 
        .A2(DP_OP_423J2_125_3477_n2314), .Y(DP_OP_422J2_124_3477_n2295) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1531 ( .A1(DP_OP_424J2_126_3477_n2308), 
        .A2(DP_OP_424J2_126_3477_n2314), .Y(DP_OP_424J2_126_3477_n2292) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1530 ( .A1(DP_OP_423J2_125_3477_n2219), 
        .A2(DP_OP_424J2_126_3477_n2314), .Y(DP_OP_424J2_126_3477_n2291) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1971 ( .A1(DP_OP_422J2_124_3477_n2880), 
        .A2(DP_OP_425J2_127_3477_n2754), .Y(DP_OP_425J2_127_3477_n2732) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1190 ( .A1(DP_OP_424J2_126_3477_n3013), 
        .A2(DP_OP_425J2_127_3477_n1963), .Y(DP_OP_425J2_127_3477_n1951) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1186 ( .A1(DP_OP_425J2_127_3477_n2967), 
        .A2(DP_OP_423J2_125_3477_n1963), .Y(DP_OP_424J2_126_3477_n1947) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1189 ( .A1(DP_OP_424J2_126_3477_n1958), 
        .A2(DP_OP_425J2_127_3477_n1963), .Y(DP_OP_424J2_126_3477_n1950) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1187 ( .A1(DP_OP_424J2_126_3477_n1956), 
        .A2(DP_OP_423J2_125_3477_n1963), .Y(DP_OP_424J2_126_3477_n1948) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1973 ( .A1(DP_OP_423J2_125_3477_n2750), 
        .A2(DP_OP_423J2_125_3477_n2754), .Y(DP_OP_423J2_125_3477_n2734) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1186 ( .A1(DP_OP_423J2_125_3477_n2967), 
        .A2(DP_OP_422J2_124_3477_n1963), .Y(DP_OP_422J2_124_3477_n1947) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1801 ( .A1(DP_OP_423J2_125_3477_n2262), 
        .A2(DP_OP_425J2_127_3477_n2579), .Y(DP_OP_425J2_127_3477_n2562) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1974 ( .A1(DP_OP_422J2_124_3477_n2179), 
        .A2(DP_OP_423J2_125_3477_n2754), .Y(DP_OP_423J2_125_3477_n2735) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1529 ( .A1(DP_OP_424J2_126_3477_n2526), 
        .A2(DP_OP_424J2_126_3477_n2314), .Y(DP_OP_422J2_124_3477_n2290) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1970 ( .A1(DP_OP_424J2_126_3477_n2747), 
        .A2(DP_OP_423J2_125_3477_n2754), .Y(DP_OP_424J2_126_3477_n2731) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1185 ( .A1(DP_OP_424J2_126_3477_n1954), 
        .A2(DP_OP_422J2_124_3477_n1963), .Y(DP_OP_424J2_126_3477_n1946) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1806 ( .A1(DP_OP_422J2_124_3477_n2575), 
        .A2(DP_OP_422J2_124_3477_n2579), .Y(DP_OP_422J2_124_3477_n2567) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1445 ( .A1(DP_OP_422J2_124_3477_n2750), 
        .A2(DP_OP_423J2_125_3477_n2226), .Y(DP_OP_423J2_125_3477_n2206) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1528 ( .A1(DP_OP_422J2_124_3477_n2305), 
        .A2(DP_OP_425J2_127_3477_n2314), .Y(DP_OP_422J2_124_3477_n2289) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2007 ( .A1(DP_OP_422J2_124_3477_n2044), 
        .A2(DP_OP_424J2_126_3477_n2797), .Y(DP_OP_424J2_126_3477_n2768) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1532 ( .A1(DP_OP_423J2_125_3477_n2617), 
        .A2(DP_OP_425J2_127_3477_n2314), .Y(DP_OP_422J2_124_3477_n2293) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1532 ( .A1(DP_OP_425J2_127_3477_n2617), 
        .A2(DP_OP_424J2_126_3477_n2314), .Y(DP_OP_424J2_126_3477_n2293) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1444 ( .A1(DP_OP_422J2_124_3477_n2837), 
        .A2(DP_OP_424J2_126_3477_n2226), .Y(DP_OP_424J2_126_3477_n2205) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2007 ( .A1(DP_OP_425J2_127_3477_n2264), 
        .A2(DP_OP_424J2_126_3477_n2797), .Y(DP_OP_423J2_125_3477_n2768) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1442 ( .A1(DP_OP_425J2_127_3477_n2219), 
        .A2(DP_OP_425J2_127_3477_n2226), .Y(DP_OP_425J2_127_3477_n2203) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1442 ( .A1(DP_OP_424J2_126_3477_n2219), 
        .A2(DP_OP_424J2_126_3477_n2226), .Y(DP_OP_424J2_126_3477_n2203) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1802 ( .A1(DP_OP_422J2_124_3477_n2263), 
        .A2(DP_OP_423J2_125_3477_n2579), .Y(DP_OP_424J2_126_3477_n2563) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1530 ( .A1(DP_OP_422J2_124_3477_n2307), 
        .A2(DP_OP_423J2_125_3477_n2314), .Y(DP_OP_422J2_124_3477_n2291) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1804 ( .A1(DP_OP_423J2_125_3477_n2573), 
        .A2(DP_OP_423J2_125_3477_n2579), .Y(DP_OP_423J2_125_3477_n2565) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1531 ( .A1(DP_OP_423J2_125_3477_n2308), 
        .A2(DP_OP_423J2_125_3477_n2314), .Y(DP_OP_423J2_125_3477_n2292) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1533 ( .A1(DP_OP_422J2_124_3477_n2178), 
        .A2(DP_OP_425J2_127_3477_n2314), .Y(DP_OP_425J2_127_3477_n2294) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1187 ( .A1(DP_OP_424J2_126_3477_n2880), 
        .A2(DP_OP_422J2_124_3477_n1963), .Y(DP_OP_422J2_124_3477_n1948) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2010 ( .A1(DP_OP_422J2_124_3477_n2795), 
        .A2(DP_OP_422J2_124_3477_n2797), .Y(DP_OP_422J2_124_3477_n2771) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1801 ( .A1(DP_OP_422J2_124_3477_n2570), 
        .A2(DP_OP_422J2_124_3477_n2579), .Y(DP_OP_422J2_124_3477_n2562) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1530 ( .A1(DP_OP_425J2_127_3477_n2307), 
        .A2(DP_OP_425J2_127_3477_n2314), .Y(DP_OP_425J2_127_3477_n2291) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1803 ( .A1(DP_OP_423J2_125_3477_n2396), 
        .A2(DP_OP_422J2_124_3477_n2579), .Y(DP_OP_422J2_124_3477_n2564) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1188 ( .A1(DP_OP_423J2_125_3477_n1957), 
        .A2(DP_OP_423J2_125_3477_n1963), .Y(DP_OP_423J2_125_3477_n1949) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1970 ( .A1(DP_OP_425J2_127_3477_n2747), 
        .A2(DP_OP_425J2_127_3477_n2754), .Y(DP_OP_425J2_127_3477_n2731) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1805 ( .A1(DP_OP_423J2_125_3477_n2574), 
        .A2(DP_OP_423J2_125_3477_n2579), .Y(DP_OP_423J2_125_3477_n2566) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1531 ( .A1(DP_OP_425J2_127_3477_n2308), 
        .A2(DP_OP_425J2_127_3477_n2314), .Y(DP_OP_425J2_127_3477_n2292) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1185 ( .A1(DP_OP_424J2_126_3477_n3008), 
        .A2(DP_OP_425J2_127_3477_n1963), .Y(DP_OP_425J2_127_3477_n1946) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1974 ( .A1(DP_OP_422J2_124_3477_n2751), 
        .A2(DP_OP_422J2_124_3477_n2754), .Y(DP_OP_422J2_124_3477_n2735) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1441 ( .A1(DP_OP_422J2_124_3477_n2218), 
        .A2(DP_OP_424J2_126_3477_n2226), .Y(DP_OP_422J2_124_3477_n2202) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1971 ( .A1(DP_OP_423J2_125_3477_n2748), 
        .A2(DP_OP_423J2_125_3477_n2754), .Y(DP_OP_423J2_125_3477_n2732) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2006 ( .A1(DP_OP_424J2_126_3477_n2791), 
        .A2(DP_OP_424J2_126_3477_n2797), .Y(DP_OP_424J2_126_3477_n2767) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1969 ( .A1(DP_OP_422J2_124_3477_n2746), 
        .A2(DP_OP_422J2_124_3477_n2754), .Y(DP_OP_422J2_124_3477_n2730) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1804 ( .A1(DP_OP_423J2_125_3477_n2397), 
        .A2(DP_OP_422J2_124_3477_n2579), .Y(DP_OP_422J2_124_3477_n2565) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1969 ( .A1(DP_OP_423J2_125_3477_n2746), 
        .A2(DP_OP_423J2_125_3477_n2754), .Y(DP_OP_423J2_125_3477_n2730) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1443 ( .A1(DP_OP_425J2_127_3477_n2616), 
        .A2(DP_OP_423J2_125_3477_n2226), .Y(DP_OP_423J2_125_3477_n2204) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2006 ( .A1(DP_OP_423J2_125_3477_n2791), 
        .A2(DP_OP_422J2_124_3477_n2797), .Y(DP_OP_423J2_125_3477_n2767) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2006 ( .A1(DP_OP_422J2_124_3477_n2791), 
        .A2(DP_OP_422J2_124_3477_n2797), .Y(DP_OP_422J2_124_3477_n2767) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1444 ( .A1(DP_OP_422J2_124_3477_n2749), 
        .A2(DP_OP_423J2_125_3477_n2226), .Y(DP_OP_423J2_125_3477_n2205) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1972 ( .A1(DP_OP_424J2_126_3477_n2749), 
        .A2(DP_OP_425J2_127_3477_n2754), .Y(DP_OP_424J2_126_3477_n2733) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1185 ( .A1(DP_OP_425J2_127_3477_n2878), 
        .A2(DP_OP_423J2_125_3477_n1963), .Y(DP_OP_423J2_125_3477_n1946) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1971 ( .A1(DP_OP_425J2_127_3477_n2220), 
        .A2(DP_OP_422J2_124_3477_n2754), .Y(DP_OP_424J2_126_3477_n2732) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2005 ( .A1(DP_OP_422J2_124_3477_n2790), 
        .A2(DP_OP_422J2_124_3477_n2797), .Y(DP_OP_422J2_124_3477_n2766) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1804 ( .A1(DP_OP_423J2_125_3477_n2265), 
        .A2(DP_OP_425J2_127_3477_n2579), .Y(DP_OP_425J2_127_3477_n2565) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2009 ( .A1(DP_OP_424J2_126_3477_n2794), 
        .A2(DP_OP_424J2_126_3477_n2797), .Y(DP_OP_424J2_126_3477_n2770) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1444 ( .A1(DP_OP_423J2_125_3477_n2705), 
        .A2(DP_OP_425J2_127_3477_n2226), .Y(DP_OP_422J2_124_3477_n2205) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1185 ( .A1(DP_OP_424J2_126_3477_n2878), 
        .A2(DP_OP_422J2_124_3477_n1963), .Y(DP_OP_422J2_124_3477_n1946) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1973 ( .A1(DP_OP_422J2_124_3477_n2750), 
        .A2(DP_OP_422J2_124_3477_n2754), .Y(DP_OP_422J2_124_3477_n2734) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2007 ( .A1(DP_OP_423J2_125_3477_n2044), 
        .A2(DP_OP_425J2_127_3477_n2797), .Y(DP_OP_425J2_127_3477_n2768) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1189 ( .A1(DP_OP_423J2_125_3477_n1958), 
        .A2(DP_OP_423J2_125_3477_n1963), .Y(DP_OP_423J2_125_3477_n1950) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1188 ( .A1(DP_OP_424J2_126_3477_n1957), 
        .A2(DP_OP_422J2_124_3477_n1963), .Y(DP_OP_424J2_126_3477_n1949) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1186 ( .A1(DP_OP_424J2_126_3477_n3009), 
        .A2(DP_OP_425J2_127_3477_n1963), .Y(DP_OP_425J2_127_3477_n1947) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2009 ( .A1(DP_OP_423J2_125_3477_n2794), 
        .A2(DP_OP_422J2_124_3477_n2797), .Y(DP_OP_423J2_125_3477_n2770) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2008 ( .A1(DP_OP_423J2_125_3477_n2793), 
        .A2(DP_OP_422J2_124_3477_n2797), .Y(DP_OP_423J2_125_3477_n2769) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1440 ( .A1(DP_OP_422J2_124_3477_n2217), 
        .A2(DP_OP_423J2_125_3477_n2226), .Y(DP_OP_422J2_124_3477_n2201) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1188 ( .A1(DP_OP_422J2_124_3477_n1957), 
        .A2(DP_OP_422J2_124_3477_n1963), .Y(DP_OP_422J2_124_3477_n1949) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2008 ( .A1(DP_OP_424J2_126_3477_n2793), 
        .A2(DP_OP_424J2_126_3477_n2797), .Y(DP_OP_424J2_126_3477_n2769) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2005 ( .A1(DP_OP_425J2_127_3477_n2790), 
        .A2(DP_OP_425J2_127_3477_n2797), .Y(DP_OP_425J2_127_3477_n2766) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1533 ( .A1(DP_OP_425J2_127_3477_n2442), 
        .A2(DP_OP_424J2_126_3477_n2314), .Y(DP_OP_422J2_124_3477_n2294) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1443 ( .A1(DP_OP_424J2_126_3477_n2220), 
        .A2(DP_OP_424J2_126_3477_n2226), .Y(DP_OP_424J2_126_3477_n2204) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1441 ( .A1(DP_OP_425J2_127_3477_n2218), 
        .A2(DP_OP_425J2_127_3477_n2226), .Y(DP_OP_425J2_127_3477_n2202) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1970 ( .A1(DP_OP_423J2_125_3477_n2747), 
        .A2(DP_OP_423J2_125_3477_n2754), .Y(DP_OP_423J2_125_3477_n2731) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1189 ( .A1(DP_OP_422J2_124_3477_n1958), 
        .A2(DP_OP_422J2_124_3477_n1963), .Y(DP_OP_422J2_124_3477_n1950) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1974 ( .A1(DP_OP_424J2_126_3477_n2751), 
        .A2(DP_OP_425J2_127_3477_n2754), .Y(DP_OP_424J2_126_3477_n2735) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1188 ( .A1(DP_OP_424J2_126_3477_n3011), 
        .A2(DP_OP_425J2_127_3477_n1963), .Y(DP_OP_425J2_127_3477_n1949) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1971 ( .A1(DP_OP_425J2_127_3477_n2616), 
        .A2(DP_OP_422J2_124_3477_n2754), .Y(DP_OP_422J2_124_3477_n2732) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1531 ( .A1(DP_OP_422J2_124_3477_n2308), 
        .A2(DP_OP_423J2_125_3477_n2314), .Y(DP_OP_422J2_124_3477_n2292) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1446 ( .A1(DP_OP_425J2_127_3477_n2619), 
        .A2(DP_OP_423J2_125_3477_n2226), .Y(DP_OP_423J2_125_3477_n2207) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1803 ( .A1(DP_OP_425J2_127_3477_n2572), 
        .A2(DP_OP_425J2_127_3477_n2579), .Y(DP_OP_425J2_127_3477_n2564) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1445 ( .A1(DP_OP_424J2_126_3477_n2618), 
        .A2(DP_OP_425J2_127_3477_n2226), .Y(DP_OP_422J2_124_3477_n2206) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1801 ( .A1(DP_OP_423J2_125_3477_n2570), 
        .A2(DP_OP_423J2_125_3477_n2579), .Y(DP_OP_423J2_125_3477_n2562) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2007 ( .A1(DP_OP_422J2_124_3477_n2792), 
        .A2(DP_OP_422J2_124_3477_n2797), .Y(DP_OP_422J2_124_3477_n2768) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1533 ( .A1(DP_OP_422J2_124_3477_n2662), 
        .A2(DP_OP_423J2_125_3477_n2314), .Y(DP_OP_423J2_125_3477_n2294) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1190 ( .A1(DP_OP_424J2_126_3477_n2047), 
        .A2(DP_OP_423J2_125_3477_n1963), .Y(DP_OP_423J2_125_3477_n1951) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1805 ( .A1(DP_OP_423J2_125_3477_n2398), 
        .A2(DP_OP_422J2_124_3477_n2579), .Y(DP_OP_422J2_124_3477_n2566) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1446 ( .A1(DP_OP_425J2_127_3477_n2707), 
        .A2(DP_OP_424J2_126_3477_n2226), .Y(DP_OP_424J2_126_3477_n2207) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1534 ( .A1(DP_OP_425J2_127_3477_n2619), 
        .A2(DP_OP_424J2_126_3477_n2314), .Y(DP_OP_424J2_126_3477_n2295) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2008 ( .A1(DP_OP_422J2_124_3477_n2793), 
        .A2(DP_OP_422J2_124_3477_n2797), .Y(DP_OP_422J2_124_3477_n2769) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1805 ( .A1(DP_OP_423J2_125_3477_n2662), 
        .A2(DP_OP_425J2_127_3477_n2579), .Y(DP_OP_424J2_126_3477_n2566) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1443 ( .A1(DP_OP_422J2_124_3477_n2220), 
        .A2(DP_OP_425J2_127_3477_n2226), .Y(DP_OP_422J2_124_3477_n2204) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1802 ( .A1(DP_OP_423J2_125_3477_n2571), 
        .A2(DP_OP_423J2_125_3477_n2579), .Y(DP_OP_423J2_125_3477_n2563) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1442 ( .A1(DP_OP_423J2_125_3477_n2219), 
        .A2(DP_OP_423J2_125_3477_n2226), .Y(DP_OP_423J2_125_3477_n2203) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1972 ( .A1(DP_OP_422J2_124_3477_n2749), 
        .A2(DP_OP_422J2_124_3477_n2754), .Y(DP_OP_422J2_124_3477_n2733) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1532 ( .A1(DP_OP_422J2_124_3477_n2177), 
        .A2(DP_OP_425J2_127_3477_n2314), .Y(DP_OP_425J2_127_3477_n2293) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1446 ( .A1(DP_OP_425J2_127_3477_n2355), 
        .A2(DP_OP_424J2_126_3477_n2226), .Y(DP_OP_422J2_124_3477_n2207) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1445 ( .A1(DP_OP_424J2_126_3477_n2750), 
        .A2(DP_OP_425J2_127_3477_n2226), .Y(DP_OP_425J2_127_3477_n2206) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1802 ( .A1(DP_OP_423J2_125_3477_n2263), 
        .A2(DP_OP_425J2_127_3477_n2579), .Y(DP_OP_425J2_127_3477_n2563) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1444 ( .A1(DP_OP_424J2_126_3477_n2749), 
        .A2(DP_OP_425J2_127_3477_n2226), .Y(DP_OP_425J2_127_3477_n2205) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2005 ( .A1(DP_OP_423J2_125_3477_n2790), 
        .A2(DP_OP_425J2_127_3477_n2797), .Y(DP_OP_423J2_125_3477_n2766) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1442 ( .A1(DP_OP_422J2_124_3477_n2219), 
        .A2(DP_OP_423J2_125_3477_n2226), .Y(DP_OP_422J2_124_3477_n2203) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1529 ( .A1(DP_OP_425J2_127_3477_n2526), 
        .A2(DP_OP_423J2_125_3477_n2314), .Y(DP_OP_423J2_125_3477_n2290) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1803 ( .A1(DP_OP_423J2_125_3477_n2572), 
        .A2(DP_OP_423J2_125_3477_n2579), .Y(DP_OP_423J2_125_3477_n2564) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1972 ( .A1(DP_OP_425J2_127_3477_n2749), 
        .A2(DP_OP_425J2_127_3477_n2754), .Y(DP_OP_425J2_127_3477_n2733) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1974 ( .A1(DP_OP_422J2_124_3477_n2883), 
        .A2(DP_OP_425J2_127_3477_n2754), .Y(DP_OP_425J2_127_3477_n2735) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1806 ( .A1(DP_OP_423J2_125_3477_n2575), 
        .A2(DP_OP_423J2_125_3477_n2579), .Y(DP_OP_423J2_125_3477_n2567) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1190 ( .A1(DP_OP_425J2_127_3477_n2971), 
        .A2(DP_OP_423J2_125_3477_n1963), .Y(DP_OP_424J2_126_3477_n1951) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1189 ( .A1(DP_OP_424J2_126_3477_n3012), 
        .A2(DP_OP_425J2_127_3477_n1963), .Y(DP_OP_425J2_127_3477_n1950) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1806 ( .A1(DP_OP_423J2_125_3477_n2663), 
        .A2(DP_OP_422J2_124_3477_n2579), .Y(DP_OP_424J2_126_3477_n2567) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1530 ( .A1(DP_OP_423J2_125_3477_n2307), 
        .A2(DP_OP_423J2_125_3477_n2314), .Y(DP_OP_423J2_125_3477_n2291) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2009 ( .A1(DP_OP_425J2_127_3477_n2794), 
        .A2(DP_OP_425J2_127_3477_n2797), .Y(DP_OP_425J2_127_3477_n2770) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2006 ( .A1(DP_OP_425J2_127_3477_n2791), 
        .A2(DP_OP_425J2_127_3477_n2797), .Y(DP_OP_425J2_127_3477_n2767) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2005 ( .A1(DP_OP_424J2_126_3477_n2790), 
        .A2(DP_OP_424J2_126_3477_n2797), .Y(DP_OP_424J2_126_3477_n2766) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1969 ( .A1(DP_OP_423J2_125_3477_n2086), 
        .A2(DP_OP_425J2_127_3477_n2754), .Y(DP_OP_425J2_127_3477_n2730) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1443 ( .A1(DP_OP_425J2_127_3477_n2220), 
        .A2(DP_OP_425J2_127_3477_n2226), .Y(DP_OP_425J2_127_3477_n2204) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1534 ( .A1(DP_OP_423J2_125_3477_n2311), 
        .A2(DP_OP_423J2_125_3477_n2314), .Y(DP_OP_423J2_125_3477_n2295) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1973 ( .A1(DP_OP_424J2_126_3477_n2750), 
        .A2(DP_OP_422J2_124_3477_n2754), .Y(DP_OP_424J2_126_3477_n2734) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1973 ( .A1(DP_OP_425J2_127_3477_n2750), 
        .A2(DP_OP_425J2_127_3477_n2754), .Y(DP_OP_425J2_127_3477_n2734) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1806 ( .A1(DP_OP_423J2_125_3477_n2267), 
        .A2(DP_OP_425J2_127_3477_n2579), .Y(DP_OP_425J2_127_3477_n2567) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1972 ( .A1(DP_OP_423J2_125_3477_n2749), 
        .A2(DP_OP_423J2_125_3477_n2754), .Y(DP_OP_423J2_125_3477_n2733) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1190 ( .A1(DP_OP_423J2_125_3477_n2971), 
        .A2(DP_OP_422J2_124_3477_n1963), .Y(DP_OP_422J2_124_3477_n1951) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2009 ( .A1(DP_OP_425J2_127_3477_n2662), 
        .A2(DP_OP_422J2_124_3477_n2797), .Y(DP_OP_422J2_124_3477_n2770) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2010 ( .A1(DP_OP_424J2_126_3477_n2795), 
        .A2(DP_OP_424J2_126_3477_n2797), .Y(DP_OP_424J2_126_3477_n2771) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1804 ( .A1(DP_OP_425J2_127_3477_n2397), 
        .A2(DP_OP_422J2_124_3477_n2579), .Y(DP_OP_424J2_126_3477_n2565) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2010 ( .A1(DP_OP_425J2_127_3477_n2795), 
        .A2(DP_OP_425J2_127_3477_n2797), .Y(DP_OP_425J2_127_3477_n2771) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2008 ( .A1(DP_OP_425J2_127_3477_n2793), 
        .A2(DP_OP_425J2_127_3477_n2797), .Y(DP_OP_425J2_127_3477_n2769) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1970 ( .A1(DP_OP_422J2_124_3477_n2747), 
        .A2(DP_OP_422J2_124_3477_n2754), .Y(DP_OP_422J2_124_3477_n2731) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1534 ( .A1(DP_OP_424J2_126_3477_n2663), 
        .A2(DP_OP_425J2_127_3477_n2314), .Y(DP_OP_425J2_127_3477_n2295) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1532 ( .A1(DP_OP_424J2_126_3477_n2397), 
        .A2(DP_OP_423J2_125_3477_n2314), .Y(DP_OP_423J2_125_3477_n2293) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1533 ( .A1(DP_OP_424J2_126_3477_n2310), 
        .A2(DP_OP_424J2_126_3477_n2314), .Y(DP_OP_424J2_126_3477_n2294) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1441 ( .A1(DP_OP_423J2_125_3477_n2218), 
        .A2(DP_OP_423J2_125_3477_n2226), .Y(DP_OP_423J2_125_3477_n2202) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1805 ( .A1(DP_OP_423J2_125_3477_n2266), 
        .A2(DP_OP_425J2_127_3477_n2579), .Y(DP_OP_425J2_127_3477_n2566) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1446 ( .A1(DP_OP_422J2_124_3477_n2091), 
        .A2(DP_OP_425J2_127_3477_n2226), .Y(DP_OP_425J2_127_3477_n2207) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1187 ( .A1(DP_OP_424J2_126_3477_n3010), 
        .A2(DP_OP_425J2_127_3477_n1963), .Y(DP_OP_425J2_127_3477_n1948) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1801 ( .A1(DP_OP_423J2_125_3477_n2658), 
        .A2(DP_OP_423J2_125_3477_n2579), .Y(DP_OP_424J2_126_3477_n2562) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2010 ( .A1(DP_OP_423J2_125_3477_n2795), 
        .A2(DP_OP_425J2_127_3477_n2797), .Y(DP_OP_423J2_125_3477_n2771) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1445 ( .A1(DP_OP_422J2_124_3477_n2838), 
        .A2(DP_OP_424J2_126_3477_n2226), .Y(DP_OP_424J2_126_3477_n2206) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1528 ( .A1(DP_OP_423J2_125_3477_n2305), 
        .A2(DP_OP_423J2_125_3477_n2314), .Y(DP_OP_423J2_125_3477_n2289) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1186 ( .A1(DP_OP_425J2_127_3477_n2879), 
        .A2(DP_OP_423J2_125_3477_n1963), .Y(DP_OP_423J2_125_3477_n1947) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1802 ( .A1(DP_OP_422J2_124_3477_n2571), 
        .A2(DP_OP_422J2_124_3477_n2579), .Y(DP_OP_422J2_124_3477_n2563) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1104 ( .A1(n509), .A2(n385), .Y(
        DP_OP_422J2_124_3477_n270) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1103 ( .A1(n498), .A2(
        DP_OP_424J2_126_3477_n2), .Y(DP_OP_422J2_124_3477_n268) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1095 ( .A1(n527), .A2(n388), .Y(
        DP_OP_422J2_124_3477_n252) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1124 ( .A1(n543), .A2(n386), .Y(
        DP_OP_425J2_127_3477_n1885) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1120 ( .A1(n474), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_424J2_126_3477_n1881) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1105 ( .A1(n497), .A2(n387), .Y(
        DP_OP_422J2_124_3477_n272) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1117 ( .A1(n332), .A2(n390), .Y(
        DP_OP_424J2_126_3477_n1878) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1098 ( .A1(n523), .A2(n391), .Y(
        DP_OP_422J2_124_3477_n258) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1115 ( .A1(n483), .A2(n387), .Y(
        DP_OP_422J2_124_3477_n460) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1108 ( .A1(n507), .A2(
        DP_OP_423J2_125_3477_n2), .Y(DP_OP_422J2_124_3477_n278) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1121 ( .A1(n328), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_425J2_127_3477_n1882) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1114 ( .A1(n476), .A2(
        DP_OP_423J2_125_3477_n2), .Y(DP_OP_424J2_126_3477_n1876) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1100 ( .A1(n511), .A2(
        DP_OP_424J2_126_3477_n2), .Y(DP_OP_422J2_124_3477_n262) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1112 ( .A1(n512), .A2(n387), .Y(
        DP_OP_424J2_126_3477_n1874) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1099 ( .A1(n519), .A2(
        DP_OP_424J2_126_3477_n2), .Y(DP_OP_422J2_124_3477_n260) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1123 ( .A1(n335), .A2(n391), .Y(
        DP_OP_425J2_127_3477_n1884) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1096 ( .A1(n524), .A2(n386), .Y(
        DP_OP_422J2_124_3477_n254) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1102 ( .A1(n510), .A2(
        DP_OP_425J2_127_3477_n2), .Y(DP_OP_422J2_124_3477_n266) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1106 ( .A1(n508), .A2(n391), .Y(
        DP_OP_422J2_124_3477_n274) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1119 ( .A1(n487), .A2(n390), .Y(
        DP_OP_424J2_126_3477_n1880) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1097 ( .A1(n520), .A2(n391), .Y(
        DP_OP_422J2_124_3477_n256) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1107 ( .A1(n482), .A2(
        DP_OP_425J2_127_3477_n2), .Y(DP_OP_422J2_124_3477_n276) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1124 ( .A1(n546), .A2(n389), .Y(
        DP_OP_423J2_125_3477_n1885) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1101 ( .A1(n499), .A2(n388), .Y(
        DP_OP_422J2_124_3477_n264) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1122 ( .A1(n538), .A2(
        DP_OP_425J2_127_3477_n2), .Y(DP_OP_425J2_127_3477_n1883) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1125 ( .A1(n344), .A2(n387), .Y(
        DP_OP_423J2_125_3477_n1886) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1104 ( .A1(n362), .A2(
        DP_OP_424J2_126_3477_n2), .Y(DP_OP_423J2_125_3477_n270) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1098 ( .A1(n525), .A2(n385), .Y(
        DP_OP_424J2_126_3477_n258) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1097 ( .A1(n522), .A2(
        DP_OP_424J2_126_3477_n2), .Y(DP_OP_424J2_126_3477_n256) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1105 ( .A1(n358), .A2(n386), .Y(
        DP_OP_423J2_125_3477_n272) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1096 ( .A1(n526), .A2(
        DP_OP_424J2_126_3477_n2), .Y(DP_OP_424J2_126_3477_n254) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1106 ( .A1(n348), .A2(
        DP_OP_423J2_125_3477_n2), .Y(DP_OP_423J2_125_3477_n274) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1095 ( .A1(n528), .A2(n391), .Y(
        DP_OP_424J2_126_3477_n252) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1123 ( .A1(n326), .A2(
        DP_OP_424J2_126_3477_n2), .Y(DP_OP_423J2_125_3477_n1884) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1107 ( .A1(n325), .A2(
        DP_OP_423J2_125_3477_n2), .Y(DP_OP_423J2_125_3477_n276) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1108 ( .A1(n333), .A2(n388), .Y(
        DP_OP_423J2_125_3477_n278) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1117 ( .A1(n477), .A2(n387), .Y(
        DP_OP_423J2_125_3477_n1878) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1109 ( .A1(n493), .A2(n387), .Y(
        DP_OP_423J2_125_3477_n280) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1118 ( .A1(n319), .A2(n390), .Y(
        DP_OP_423J2_125_3477_n1879) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1105 ( .A1(n502), .A2(n390), .Y(
        DP_OP_424J2_126_3477_n272) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1104 ( .A1(n516), .A2(
        DP_OP_423J2_125_3477_n2), .Y(DP_OP_424J2_126_3477_n270) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1100 ( .A1(n361), .A2(n391), .Y(
        DP_OP_423J2_125_3477_n262) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1103 ( .A1(n503), .A2(
        DP_OP_425J2_127_3477_n2), .Y(DP_OP_424J2_126_3477_n268) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1101 ( .A1(n357), .A2(
        DP_OP_424J2_126_3477_n2), .Y(DP_OP_423J2_125_3477_n264) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1101 ( .A1(n504), .A2(
        DP_OP_423J2_125_3477_n2), .Y(DP_OP_424J2_126_3477_n264) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1102 ( .A1(n347), .A2(n391), .Y(
        DP_OP_423J2_125_3477_n266) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1125 ( .A1(n342), .A2(n386), .Y(
        DP_OP_424J2_126_3477_n1886) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1120 ( .A1(n321), .A2(
        DP_OP_425J2_127_3477_n2), .Y(DP_OP_425J2_127_3477_n1881) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1100 ( .A1(n518), .A2(n386), .Y(
        DP_OP_424J2_126_3477_n262) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1103 ( .A1(n354), .A2(
        DP_OP_423J2_125_3477_n2), .Y(DP_OP_423J2_125_3477_n268) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1099 ( .A1(n521), .A2(n387), .Y(
        DP_OP_424J2_126_3477_n260) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1116 ( .A1(n340), .A2(n390), .Y(
        DP_OP_425J2_127_3477_n1877) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1113 ( .A1(n366), .A2(n388), .Y(
        DP_OP_423J2_125_3477_n1875) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1114 ( .A1(n323), .A2(n389), .Y(
        DP_OP_425J2_127_3477_n1876) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1110 ( .A1(n506), .A2(n385), .Y(
        DP_OP_422J2_124_3477_n1873) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1119 ( .A1(n484), .A2(
        DP_OP_425J2_127_3477_n2), .Y(DP_OP_422J2_124_3477_n1880) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1125 ( .A1(n341), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_422J2_124_3477_n1886) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1122 ( .A1(n490), .A2(n388), .Y(
        DP_OP_424J2_126_3477_n1883) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1122 ( .A1(n545), .A2(n390), .Y(
        DP_OP_422J2_124_3477_n1883) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1117 ( .A1(n478), .A2(n389), .Y(
        DP_OP_425J2_127_3477_n1878) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1125 ( .A1(n343), .A2(n390), .Y(
        DP_OP_425J2_127_3477_n1886) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1124 ( .A1(n544), .A2(n389), .Y(
        DP_OP_424J2_126_3477_n1885) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1121 ( .A1(n480), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_424J2_126_3477_n1882) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1123 ( .A1(n488), .A2(n385), .Y(
        DP_OP_422J2_124_3477_n1884) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1119 ( .A1(n330), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_425J2_127_3477_n1880) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1118 ( .A1(n473), .A2(n388), .Y(
        DP_OP_422J2_124_3477_n1879) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1117 ( .A1(n331), .A2(n390), .Y(
        DP_OP_422J2_124_3477_n1878) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1123 ( .A1(n481), .A2(
        DP_OP_423J2_125_3477_n2), .Y(DP_OP_424J2_126_3477_n1884) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1110 ( .A1(n350), .A2(n385), .Y(
        DP_OP_425J2_127_3477_n1873) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1121 ( .A1(n479), .A2(
        DP_OP_425J2_127_3477_n2), .Y(DP_OP_422J2_124_3477_n1882) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1106 ( .A1(n515), .A2(n389), .Y(
        DP_OP_424J2_126_3477_n274) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1096 ( .A1(n376), .A2(
        DP_OP_424J2_126_3477_n2), .Y(DP_OP_425J2_127_3477_n254) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1097 ( .A1(n374), .A2(n387), .Y(
        DP_OP_425J2_127_3477_n256) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1098 ( .A1(n370), .A2(
        DP_OP_424J2_126_3477_n2), .Y(DP_OP_425J2_127_3477_n258) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1099 ( .A1(n372), .A2(n385), .Y(
        DP_OP_425J2_127_3477_n260) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1100 ( .A1(n360), .A2(n387), .Y(
        DP_OP_425J2_127_3477_n262) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1101 ( .A1(n356), .A2(
        DP_OP_425J2_127_3477_n2), .Y(DP_OP_425J2_127_3477_n264) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1102 ( .A1(n349), .A2(n389), .Y(
        DP_OP_425J2_127_3477_n266) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1103 ( .A1(n353), .A2(n385), .Y(
        DP_OP_425J2_127_3477_n268) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1121 ( .A1(n327), .A2(
        DP_OP_423J2_125_3477_n2), .Y(DP_OP_423J2_125_3477_n1882) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1104 ( .A1(n359), .A2(
        DP_OP_423J2_125_3477_n2), .Y(DP_OP_425J2_127_3477_n270) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1105 ( .A1(n355), .A2(
        DP_OP_425J2_127_3477_n2), .Y(DP_OP_425J2_127_3477_n272) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1116 ( .A1(n548), .A2(n389), .Y(
        DP_OP_423J2_125_3477_n1877) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1119 ( .A1(n329), .A2(n388), .Y(
        DP_OP_423J2_125_3477_n1880) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1116 ( .A1(n549), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_422J2_124_3477_n1877) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1122 ( .A1(n466), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_423J2_125_3477_n1883) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1116 ( .A1(n489), .A2(n387), .Y(
        DP_OP_424J2_126_3477_n1877) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1124 ( .A1(n345), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_422J2_124_3477_n1885) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1120 ( .A1(n472), .A2(n389), .Y(
        DP_OP_422J2_124_3477_n1881) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1095 ( .A1(n380), .A2(n385), .Y(
        DP_OP_425J2_127_3477_n252) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1118 ( .A1(n318), .A2(n390), .Y(
        DP_OP_425J2_127_3477_n1879) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1096 ( .A1(n375), .A2(n385), .Y(
        DP_OP_423J2_125_3477_n254) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1097 ( .A1(n373), .A2(n385), .Y(
        DP_OP_423J2_125_3477_n256) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1095 ( .A1(n379), .A2(
        DP_OP_424J2_126_3477_n2), .Y(DP_OP_423J2_125_3477_n252) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1108 ( .A1(n514), .A2(n386), .Y(
        DP_OP_424J2_126_3477_n278) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1120 ( .A1(n320), .A2(n386), .Y(
        DP_OP_423J2_125_3477_n1881) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1098 ( .A1(n369), .A2(n388), .Y(
        DP_OP_423J2_125_3477_n258) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1118 ( .A1(n475), .A2(n387), .Y(
        DP_OP_424J2_126_3477_n1879) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1106 ( .A1(n352), .A2(
        DP_OP_425J2_127_3477_n2), .Y(DP_OP_425J2_127_3477_n274) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1108 ( .A1(n339), .A2(n391), .Y(
        DP_OP_425J2_127_3477_n278) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1107 ( .A1(n324), .A2(n389), .Y(
        DP_OP_425J2_127_3477_n276) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1489 ( .A1(DP_OP_423J2_125_3477_n2662), 
        .A2(DP_OP_422J2_124_3477_n2270), .Y(DP_OP_422J2_124_3477_n2250) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1305 ( .A1(DP_OP_422J2_124_3477_n2090), 
        .A2(DP_OP_422J2_124_3477_n2093), .Y(DP_OP_422J2_124_3477_n2066) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1664 ( .A1(DP_OP_422J2_124_3477_n2441), 
        .A2(DP_OP_422J2_124_3477_n2446), .Y(DP_OP_422J2_124_3477_n2425) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1407 ( .A1(DP_OP_423J2_125_3477_n2748), 
        .A2(DP_OP_422J2_124_3477_n2183), .Y(DP_OP_422J2_124_3477_n2168) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1743 ( .A1(DP_OP_422J2_124_3477_n2528), 
        .A2(DP_OP_422J2_124_3477_n2533), .Y(DP_OP_422J2_124_3477_n2504) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2199 ( .A1(DP_OP_423J2_125_3477_n2000), 
        .A2(DP_OP_422J2_124_3477_n2975), .Y(DP_OP_422J2_124_3477_n2960) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1178 ( .A1(DP_OP_423J2_125_3477_n2967), 
        .A2(DP_OP_422J2_124_3477_n1962), .Y(DP_OP_422J2_124_3477_n1939) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2104 ( .A1(DP_OP_425J2_127_3477_n2749), 
        .A2(DP_OP_422J2_124_3477_n2886), .Y(DP_OP_422J2_124_3477_n2865) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1618 ( .A1(DP_OP_423J2_125_3477_n2527), 
        .A2(DP_OP_425J2_127_3477_n2402), .Y(DP_OP_422J2_124_3477_n2379) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1172 ( .A1(DP_OP_422J2_124_3477_n1957), 
        .A2(DP_OP_422J2_124_3477_n1961), .Y(DP_OP_422J2_124_3477_n1933) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1265 ( .A1(DP_OP_423J2_125_3477_n2878), 
        .A2(DP_OP_422J2_124_3477_n2050), .Y(DP_OP_422J2_124_3477_n2026) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1671 ( .A1(DP_OP_423J2_125_3477_n2484), 
        .A2(DP_OP_422J2_124_3477_n2447), .Y(DP_OP_422J2_124_3477_n2432) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1611 ( .A1(DP_OP_423J2_125_3477_n2528), 
        .A2(DP_OP_422J2_124_3477_n2401), .Y(DP_OP_422J2_124_3477_n2372) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1660 ( .A1(DP_OP_423J2_125_3477_n2481), 
        .A2(DP_OP_422J2_124_3477_n2446), .Y(DP_OP_422J2_124_3477_n2421) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1521 ( .A1(DP_OP_425J2_127_3477_n2438), 
        .A2(DP_OP_422J2_124_3477_n2313), .Y(DP_OP_422J2_124_3477_n2282) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1890 ( .A1(DP_OP_422J2_124_3477_n2659), 
        .A2(DP_OP_422J2_124_3477_n2667), .Y(DP_OP_422J2_124_3477_n2651) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1269 ( .A1(DP_OP_424J2_126_3477_n2794), 
        .A2(DP_OP_422J2_124_3477_n2050), .Y(DP_OP_422J2_124_3477_n2030) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1845 ( .A1(DP_OP_425J2_127_3477_n2482), 
        .A2(DP_OP_422J2_124_3477_n2623), .Y(DP_OP_422J2_124_3477_n2606) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1179 ( .A1(DP_OP_424J2_126_3477_n2880), 
        .A2(DP_OP_422J2_124_3477_n1962), .Y(DP_OP_422J2_124_3477_n1940) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2182 ( .A1(DP_OP_425J2_127_3477_n2835), 
        .A2(DP_OP_422J2_124_3477_n2973), .Y(DP_OP_422J2_124_3477_n2943) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2070 ( .A1(DP_OP_424J2_126_3477_n2751), 
        .A2(DP_OP_423J2_125_3477_n2843), .Y(DP_OP_423J2_125_3477_n2831) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1961 ( .A1(DP_OP_422J2_124_3477_n2746), 
        .A2(DP_OP_422J2_124_3477_n2753), .Y(DP_OP_422J2_124_3477_n2722) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1831 ( .A1(DP_OP_422J2_124_3477_n2616), 
        .A2(DP_OP_422J2_124_3477_n2621), .Y(DP_OP_422J2_124_3477_n2592) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1400 ( .A1(DP_OP_422J2_124_3477_n2177), 
        .A2(DP_OP_422J2_124_3477_n2182), .Y(DP_OP_422J2_124_3477_n2161) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1390 ( .A1(DP_OP_425J2_127_3477_n2307), 
        .A2(DP_OP_422J2_124_3477_n2181), .Y(DP_OP_422J2_124_3477_n2151) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1261 ( .A1(DP_OP_424J2_126_3477_n2794), 
        .A2(DP_OP_422J2_124_3477_n2049), .Y(DP_OP_422J2_124_3477_n2022) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1537 ( .A1(DP_OP_425J2_127_3477_n2438), 
        .A2(DP_OP_422J2_124_3477_n2315), .Y(DP_OP_422J2_124_3477_n2298) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1391 ( .A1(DP_OP_423J2_125_3477_n2748), 
        .A2(DP_OP_422J2_124_3477_n2181), .Y(DP_OP_422J2_124_3477_n2152) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2146 ( .A1(DP_OP_422J2_124_3477_n2923), 
        .A2(DP_OP_422J2_124_3477_n2930), .Y(DP_OP_422J2_124_3477_n2907) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1920 ( .A1(DP_OP_424J2_126_3477_n2353), 
        .A2(DP_OP_422J2_124_3477_n2709), .Y(DP_OP_422J2_124_3477_n2681) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1744 ( .A1(DP_OP_423J2_125_3477_n2441), 
        .A2(DP_OP_422J2_124_3477_n2533), .Y(DP_OP_422J2_124_3477_n2505) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1526 ( .A1(DP_OP_422J2_124_3477_n2311), 
        .A2(DP_OP_422J2_124_3477_n2313), .Y(DP_OP_422J2_124_3477_n2287) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1171 ( .A1(DP_OP_425J2_127_3477_n2088), 
        .A2(DP_OP_422J2_124_3477_n1961), .Y(DP_OP_422J2_124_3477_n1932) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1884 ( .A1(DP_OP_424J2_126_3477_n2397), 
        .A2(DP_OP_422J2_124_3477_n2666), .Y(DP_OP_422J2_124_3477_n2645) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1708 ( .A1(DP_OP_422J2_124_3477_n2485), 
        .A2(DP_OP_422J2_124_3477_n2490), .Y(DP_OP_422J2_124_3477_n2469) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1880 ( .A1(DP_OP_425J2_127_3477_n2525), 
        .A2(DP_OP_422J2_124_3477_n2666), .Y(DP_OP_422J2_124_3477_n2641) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1397 ( .A1(DP_OP_423J2_125_3477_n2746), 
        .A2(DP_OP_422J2_124_3477_n2182), .Y(DP_OP_422J2_124_3477_n2158) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2112 ( .A1(DP_OP_425J2_127_3477_n2749), 
        .A2(DP_OP_422J2_124_3477_n2887), .Y(DP_OP_422J2_124_3477_n2873) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1525 ( .A1(DP_OP_424J2_126_3477_n2530), 
        .A2(DP_OP_422J2_124_3477_n2313), .Y(DP_OP_422J2_124_3477_n2286) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1846 ( .A1(DP_OP_423J2_125_3477_n2351), 
        .A2(DP_OP_422J2_124_3477_n2623), .Y(DP_OP_422J2_124_3477_n2607) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1306 ( .A1(DP_OP_422J2_124_3477_n2091), 
        .A2(DP_OP_422J2_124_3477_n2093), .Y(DP_OP_422J2_124_3477_n2067) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2069 ( .A1(DP_OP_422J2_124_3477_n2838), 
        .A2(DP_OP_422J2_124_3477_n2843), .Y(DP_OP_422J2_124_3477_n2830) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2153 ( .A1(DP_OP_422J2_124_3477_n2922), 
        .A2(DP_OP_422J2_124_3477_n2931), .Y(DP_OP_422J2_124_3477_n2914) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1570 ( .A1(DP_OP_422J2_124_3477_n2355), 
        .A2(DP_OP_422J2_124_3477_n2357), .Y(DP_OP_422J2_124_3477_n2331) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1883 ( .A1(DP_OP_425J2_127_3477_n2528), 
        .A2(DP_OP_422J2_124_3477_n2666), .Y(DP_OP_422J2_124_3477_n2644) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1758 ( .A1(DP_OP_423J2_125_3477_n2439), 
        .A2(DP_OP_422J2_124_3477_n2535), .Y(DP_OP_422J2_124_3477_n2519) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2014 ( .A1(DP_OP_422J2_124_3477_n2791), 
        .A2(DP_OP_422J2_124_3477_n2798), .Y(DP_OP_422J2_124_3477_n2775) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1523 ( .A1(DP_OP_422J2_124_3477_n2308), 
        .A2(DP_OP_422J2_124_3477_n2313), .Y(DP_OP_422J2_124_3477_n2284) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1450 ( .A1(DP_OP_422J2_124_3477_n2219), 
        .A2(DP_OP_422J2_124_3477_n2227), .Y(DP_OP_422J2_124_3477_n2211) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2181 ( .A1(DP_OP_423J2_125_3477_n1998), 
        .A2(DP_OP_422J2_124_3477_n2973), .Y(DP_OP_422J2_124_3477_n2942) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1829 ( .A1(DP_OP_425J2_127_3477_n2482), 
        .A2(DP_OP_422J2_124_3477_n2621), .Y(DP_OP_422J2_124_3477_n2590) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1435 ( .A1(DP_OP_422J2_124_3477_n2220), 
        .A2(DP_OP_422J2_124_3477_n2225), .Y(DP_OP_422J2_124_3477_n2196) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1665 ( .A1(DP_OP_422J2_124_3477_n2442), 
        .A2(DP_OP_422J2_124_3477_n2446), .Y(DP_OP_422J2_124_3477_n2426) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1892 ( .A1(DP_OP_425J2_127_3477_n2529), 
        .A2(DP_OP_422J2_124_3477_n2667), .Y(DP_OP_422J2_124_3477_n2653) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1586 ( .A1(DP_OP_423J2_125_3477_n2355), 
        .A2(DP_OP_423J2_125_3477_n2359), .Y(DP_OP_423J2_125_3477_n2347) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2109 ( .A1(DP_OP_422J2_124_3477_n2878), 
        .A2(DP_OP_422J2_124_3477_n2887), .Y(DP_OP_422J2_124_3477_n2870) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1797 ( .A1(DP_OP_423J2_125_3477_n2398), 
        .A2(DP_OP_422J2_124_3477_n2578), .Y(DP_OP_422J2_124_3477_n2558) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2200 ( .A1(DP_OP_422J2_124_3477_n2969), 
        .A2(DP_OP_422J2_124_3477_n2975), .Y(DP_OP_422J2_124_3477_n2961) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1619 ( .A1(DP_OP_423J2_125_3477_n2528), 
        .A2(DP_OP_423J2_125_3477_n2402), .Y(DP_OP_422J2_124_3477_n2380) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1792 ( .A1(DP_OP_422J2_124_3477_n2569), 
        .A2(DP_OP_422J2_124_3477_n2578), .Y(DP_OP_422J2_124_3477_n2553) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2230 ( .A1(DP_OP_422J2_124_3477_n3013), 
        .A2(DP_OP_422J2_124_3477_n3015), .Y(DP_OP_422J2_124_3477_n2989) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2234 ( .A1(DP_OP_422J2_124_3477_n3009), 
        .A2(DP_OP_422J2_124_3477_n3016), .Y(DP_OP_422J2_124_3477_n2993) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2102 ( .A1(DP_OP_423J2_125_3477_n2087), 
        .A2(DP_OP_422J2_124_3477_n2886), .Y(DP_OP_422J2_124_3477_n2863) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2228 ( .A1(DP_OP_422J2_124_3477_n3011), 
        .A2(DP_OP_422J2_124_3477_n3015), .Y(DP_OP_422J2_124_3477_n2987) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1539 ( .A1(DP_OP_422J2_124_3477_n2308), 
        .A2(DP_OP_422J2_124_3477_n2315), .Y(DP_OP_422J2_124_3477_n2300) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1215 ( .A1(DP_OP_422J2_124_3477_n2000), 
        .A2(DP_OP_422J2_124_3477_n2005), .Y(DP_OP_422J2_124_3477_n1976) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1625 ( .A1(DP_OP_423J2_125_3477_n2526), 
        .A2(DP_OP_422J2_124_3477_n2403), .Y(DP_OP_422J2_124_3477_n2386) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1613 ( .A1(DP_OP_423J2_125_3477_n2530), 
        .A2(DP_OP_422J2_124_3477_n2401), .Y(DP_OP_422J2_124_3477_n2374) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1452 ( .A1(DP_OP_423J2_125_3477_n2705), 
        .A2(DP_OP_422J2_124_3477_n2227), .Y(DP_OP_422J2_124_3477_n2213) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2225 ( .A1(DP_OP_422J2_124_3477_n3008), 
        .A2(DP_OP_422J2_124_3477_n3015), .Y(DP_OP_422J2_124_3477_n2984) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1232 ( .A1(DP_OP_425J2_127_3477_n2133), 
        .A2(DP_OP_422J2_124_3477_n2007), .Y(DP_OP_422J2_124_3477_n1993) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1493 ( .A1(DP_OP_422J2_124_3477_n2262), 
        .A2(DP_OP_422J2_124_3477_n2271), .Y(DP_OP_422J2_124_3477_n2254) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1875 ( .A1(DP_OP_423J2_125_3477_n2308), 
        .A2(DP_OP_425J2_127_3477_n2665), .Y(DP_OP_422J2_124_3477_n2636) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1355 ( .A1(DP_OP_422J2_124_3477_n2132), 
        .A2(DP_OP_422J2_124_3477_n2138), .Y(DP_OP_422J2_124_3477_n2116) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1672 ( .A1(DP_OP_422J2_124_3477_n2441), 
        .A2(DP_OP_422J2_124_3477_n2447), .Y(DP_OP_422J2_124_3477_n2433) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1230 ( .A1(DP_OP_424J2_126_3477_n2835), 
        .A2(DP_OP_422J2_124_3477_n2007), .Y(DP_OP_422J2_124_3477_n1991) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1882 ( .A1(DP_OP_422J2_124_3477_n2659), 
        .A2(DP_OP_422J2_124_3477_n2666), .Y(DP_OP_422J2_124_3477_n2643) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2022 ( .A1(DP_OP_422J2_124_3477_n2791), 
        .A2(DP_OP_422J2_124_3477_n2799), .Y(DP_OP_422J2_124_3477_n2783) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1217 ( .A1(DP_OP_425J2_127_3477_n2134), 
        .A2(DP_OP_422J2_124_3477_n2005), .Y(DP_OP_422J2_124_3477_n1978) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1224 ( .A1(DP_OP_425J2_127_3477_n2133), 
        .A2(DP_OP_422J2_124_3477_n2006), .Y(DP_OP_422J2_124_3477_n1985) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1889 ( .A1(DP_OP_422J2_124_3477_n2658), 
        .A2(DP_OP_422J2_124_3477_n2667), .Y(DP_OP_422J2_124_3477_n2650) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2198 ( .A1(DP_OP_425J2_127_3477_n2835), 
        .A2(DP_OP_422J2_124_3477_n2975), .Y(DP_OP_422J2_124_3477_n2959) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1498 ( .A1(DP_OP_423J2_125_3477_n2267), 
        .A2(DP_OP_424J2_126_3477_n2271), .Y(DP_OP_423J2_125_3477_n2259) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1229 ( .A1(DP_OP_423J2_125_3477_n2922), 
        .A2(DP_OP_422J2_124_3477_n2007), .Y(DP_OP_422J2_124_3477_n1990) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1405 ( .A1(DP_OP_424J2_126_3477_n2658), 
        .A2(DP_OP_422J2_124_3477_n2183), .Y(DP_OP_422J2_124_3477_n2166) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2053 ( .A1(DP_OP_422J2_124_3477_n2838), 
        .A2(DP_OP_424J2_126_3477_n2841), .Y(DP_OP_422J2_124_3477_n2814) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1169 ( .A1(DP_OP_425J2_127_3477_n2086), 
        .A2(DP_OP_422J2_124_3477_n1961), .Y(DP_OP_422J2_124_3477_n1930) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1260 ( .A1(DP_OP_422J2_124_3477_n2045), 
        .A2(DP_OP_422J2_124_3477_n2049), .Y(DP_OP_422J2_124_3477_n2021) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1752 ( .A1(DP_OP_423J2_125_3477_n2441), 
        .A2(DP_OP_422J2_124_3477_n2534), .Y(DP_OP_422J2_124_3477_n2513) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1524 ( .A1(DP_OP_423J2_125_3477_n2617), 
        .A2(DP_OP_422J2_124_3477_n2313), .Y(DP_OP_422J2_124_3477_n2285) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1225 ( .A1(DP_OP_425J2_127_3477_n2134), 
        .A2(DP_OP_422J2_124_3477_n2006), .Y(DP_OP_422J2_124_3477_n1986) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1885 ( .A1(DP_OP_422J2_124_3477_n2662), 
        .A2(DP_OP_422J2_124_3477_n2666), .Y(DP_OP_422J2_124_3477_n2646) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1494 ( .A1(DP_OP_422J2_124_3477_n2263), 
        .A2(DP_OP_422J2_124_3477_n2271), .Y(DP_OP_422J2_124_3477_n2255) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1477 ( .A1(DP_OP_422J2_124_3477_n2262), 
        .A2(DP_OP_422J2_124_3477_n2269), .Y(DP_OP_422J2_124_3477_n2238) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1877 ( .A1(DP_OP_422J2_124_3477_n2662), 
        .A2(DP_OP_424J2_126_3477_n2665), .Y(DP_OP_422J2_124_3477_n2638) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1267 ( .A1(DP_OP_422J2_124_3477_n2044), 
        .A2(DP_OP_422J2_124_3477_n2050), .Y(DP_OP_422J2_124_3477_n2028) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1484 ( .A1(DP_OP_422J2_124_3477_n2261), 
        .A2(DP_OP_422J2_124_3477_n2270), .Y(DP_OP_422J2_124_3477_n2245) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2060 ( .A1(DP_OP_422J2_124_3477_n2837), 
        .A2(DP_OP_422J2_124_3477_n2842), .Y(DP_OP_422J2_124_3477_n2821) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1488 ( .A1(DP_OP_422J2_124_3477_n2265), 
        .A2(DP_OP_422J2_124_3477_n2270), .Y(DP_OP_422J2_124_3477_n2249) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1304 ( .A1(DP_OP_424J2_126_3477_n2749), 
        .A2(DP_OP_422J2_124_3477_n2093), .Y(DP_OP_422J2_124_3477_n2065) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1701 ( .A1(DP_OP_422J2_124_3477_n2486), 
        .A2(DP_OP_422J2_124_3477_n2489), .Y(DP_OP_422J2_124_3477_n2462) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1540 ( .A1(DP_OP_425J2_127_3477_n2441), 
        .A2(DP_OP_422J2_124_3477_n2315), .Y(DP_OP_422J2_124_3477_n2301) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1482 ( .A1(DP_OP_422J2_124_3477_n2267), 
        .A2(DP_OP_422J2_124_3477_n2269), .Y(DP_OP_422J2_124_3477_n2243) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2236 ( .A1(DP_OP_422J2_124_3477_n3011), 
        .A2(DP_OP_422J2_124_3477_n3016), .Y(DP_OP_422J2_124_3477_n2995) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2229 ( .A1(DP_OP_422J2_124_3477_n3012), 
        .A2(DP_OP_422J2_124_3477_n3015), .Y(DP_OP_422J2_124_3477_n2988) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1538 ( .A1(DP_OP_422J2_124_3477_n2307), 
        .A2(DP_OP_422J2_124_3477_n2315), .Y(DP_OP_422J2_124_3477_n2299) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2142 ( .A1(DP_OP_422J2_124_3477_n2927), 
        .A2(DP_OP_422J2_124_3477_n2929), .Y(DP_OP_422J2_124_3477_n2903) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1833 ( .A1(DP_OP_423J2_125_3477_n2354), 
        .A2(DP_OP_422J2_124_3477_n2621), .Y(DP_OP_422J2_124_3477_n2594) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1926 ( .A1(DP_OP_424J2_126_3477_n2351), 
        .A2(DP_OP_422J2_124_3477_n2710), .Y(DP_OP_422J2_124_3477_n2687) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1964 ( .A1(DP_OP_422J2_124_3477_n2749), 
        .A2(DP_OP_422J2_124_3477_n2753), .Y(DP_OP_422J2_124_3477_n2725) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2111 ( .A1(DP_OP_422J2_124_3477_n2880), 
        .A2(DP_OP_422J2_124_3477_n2887), .Y(DP_OP_422J2_124_3477_n2872) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1748 ( .A1(DP_OP_423J2_125_3477_n2437), 
        .A2(DP_OP_422J2_124_3477_n2534), .Y(DP_OP_422J2_124_3477_n2509) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1757 ( .A1(DP_OP_422J2_124_3477_n2526), 
        .A2(DP_OP_422J2_124_3477_n2535), .Y(DP_OP_422J2_124_3477_n2518) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1542 ( .A1(DP_OP_423J2_125_3477_n2311), 
        .A2(DP_OP_423J2_125_3477_n2315), .Y(DP_OP_423J2_125_3477_n2303) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2103 ( .A1(DP_OP_422J2_124_3477_n2880), 
        .A2(DP_OP_422J2_124_3477_n2886), .Y(DP_OP_422J2_124_3477_n2864) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1670 ( .A1(DP_OP_422J2_124_3477_n2439), 
        .A2(DP_OP_422J2_124_3477_n2447), .Y(DP_OP_422J2_124_3477_n2431) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2110 ( .A1(DP_OP_423J2_125_3477_n2087), 
        .A2(DP_OP_422J2_124_3477_n2887), .Y(DP_OP_422J2_124_3477_n2871) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1750 ( .A1(DP_OP_423J2_125_3477_n2439), 
        .A2(DP_OP_422J2_124_3477_n2534), .Y(DP_OP_422J2_124_3477_n2511) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1495 ( .A1(DP_OP_424J2_126_3477_n2572), 
        .A2(DP_OP_422J2_124_3477_n2271), .Y(DP_OP_422J2_124_3477_n2256) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1715 ( .A1(DP_OP_422J2_124_3477_n2484), 
        .A2(DP_OP_422J2_124_3477_n2491), .Y(DP_OP_422J2_124_3477_n2476) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1919 ( .A1(DP_OP_422J2_124_3477_n2704), 
        .A2(DP_OP_422J2_124_3477_n2709), .Y(DP_OP_422J2_124_3477_n2680) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1568 ( .A1(DP_OP_422J2_124_3477_n2353), 
        .A2(DP_OP_422J2_124_3477_n2357), .Y(DP_OP_422J2_124_3477_n2329) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1700 ( .A1(DP_OP_422J2_124_3477_n2485), 
        .A2(DP_OP_422J2_124_3477_n2489), .Y(DP_OP_422J2_124_3477_n2461) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1496 ( .A1(DP_OP_422J2_124_3477_n2265), 
        .A2(DP_OP_422J2_124_3477_n2271), .Y(DP_OP_422J2_124_3477_n2257) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2148 ( .A1(DP_OP_424J2_126_3477_n2133), 
        .A2(DP_OP_422J2_124_3477_n2930), .Y(DP_OP_422J2_124_3477_n2909) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1669 ( .A1(DP_OP_423J2_125_3477_n2482), 
        .A2(DP_OP_422J2_124_3477_n2447), .Y(DP_OP_422J2_124_3477_n2430) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1262 ( .A1(DP_OP_422J2_124_3477_n2047), 
        .A2(DP_OP_422J2_124_3477_n2049), .Y(DP_OP_422J2_124_3477_n2023) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1834 ( .A1(DP_OP_422J2_124_3477_n2619), 
        .A2(DP_OP_422J2_124_3477_n2621), .Y(DP_OP_422J2_124_3477_n2595) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1873 ( .A1(DP_OP_422J2_124_3477_n2658), 
        .A2(DP_OP_423J2_125_3477_n2665), .Y(DP_OP_422J2_124_3477_n2634) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1662 ( .A1(DP_OP_422J2_124_3477_n2439), 
        .A2(DP_OP_422J2_124_3477_n2446), .Y(DP_OP_422J2_124_3477_n2423) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1487 ( .A1(DP_OP_425J2_127_3477_n2396), 
        .A2(DP_OP_422J2_124_3477_n2270), .Y(DP_OP_422J2_124_3477_n2248) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1697 ( .A1(DP_OP_422J2_124_3477_n2482), 
        .A2(DP_OP_422J2_124_3477_n2489), .Y(DP_OP_422J2_124_3477_n2458) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1963 ( .A1(DP_OP_425J2_127_3477_n2616), 
        .A2(DP_OP_422J2_124_3477_n2753), .Y(DP_OP_422J2_124_3477_n2724) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1876 ( .A1(DP_OP_425J2_127_3477_n2529), 
        .A2(DP_OP_425J2_127_3477_n2665), .Y(DP_OP_422J2_124_3477_n2637) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1480 ( .A1(DP_OP_422J2_124_3477_n2265), 
        .A2(DP_OP_422J2_124_3477_n2269), .Y(DP_OP_422J2_124_3477_n2241) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1713 ( .A1(DP_OP_422J2_124_3477_n2482), 
        .A2(DP_OP_422J2_124_3477_n2491), .Y(DP_OP_422J2_124_3477_n2474) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2145 ( .A1(DP_OP_422J2_124_3477_n2922), 
        .A2(DP_OP_422J2_124_3477_n2930), .Y(DP_OP_422J2_124_3477_n2906) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1349 ( .A1(DP_OP_422J2_124_3477_n2134), 
        .A2(DP_OP_422J2_124_3477_n2137), .Y(DP_OP_422J2_124_3477_n2110) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1741 ( .A1(DP_OP_422J2_124_3477_n2526), 
        .A2(DP_OP_422J2_124_3477_n2533), .Y(DP_OP_422J2_124_3477_n2502) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1398 ( .A1(DP_OP_423J2_125_3477_n2747), 
        .A2(DP_OP_422J2_124_3477_n2182), .Y(DP_OP_422J2_124_3477_n2159) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1393 ( .A1(DP_OP_422J2_124_3477_n2178), 
        .A2(DP_OP_422J2_124_3477_n2181), .Y(DP_OP_422J2_124_3477_n2154) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1346 ( .A1(DP_OP_424J2_126_3477_n2703), 
        .A2(DP_OP_422J2_124_3477_n2137), .Y(DP_OP_422J2_124_3477_n2107) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1742 ( .A1(DP_OP_423J2_125_3477_n2439), 
        .A2(DP_OP_422J2_124_3477_n2533), .Y(DP_OP_422J2_124_3477_n2503) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1575 ( .A1(DP_OP_424J2_126_3477_n2484), 
        .A2(DP_OP_422J2_124_3477_n2358), .Y(DP_OP_422J2_124_3477_n2336) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2186 ( .A1(DP_OP_422J2_124_3477_n2971), 
        .A2(DP_OP_422J2_124_3477_n2973), .Y(DP_OP_422J2_124_3477_n2947) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1760 ( .A1(DP_OP_423J2_125_3477_n2441), 
        .A2(DP_OP_422J2_124_3477_n2535), .Y(DP_OP_422J2_124_3477_n2521) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1569 ( .A1(DP_OP_422J2_124_3477_n2354), 
        .A2(DP_OP_422J2_124_3477_n2357), .Y(DP_OP_422J2_124_3477_n2330) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1436 ( .A1(DP_OP_423J2_125_3477_n2705), 
        .A2(DP_OP_422J2_124_3477_n2225), .Y(DP_OP_422J2_124_3477_n2197) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1627 ( .A1(DP_OP_423J2_125_3477_n2528), 
        .A2(DP_OP_422J2_124_3477_n2403), .Y(DP_OP_422J2_124_3477_n2388) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2155 ( .A1(DP_OP_422J2_124_3477_n2924), 
        .A2(DP_OP_422J2_124_3477_n2931), .Y(DP_OP_422J2_124_3477_n2916) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1830 ( .A1(DP_OP_424J2_126_3477_n2439), 
        .A2(DP_OP_422J2_124_3477_n2621), .Y(DP_OP_422J2_124_3477_n2591) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1357 ( .A1(DP_OP_422J2_124_3477_n2134), 
        .A2(DP_OP_422J2_124_3477_n2138), .Y(DP_OP_422J2_124_3477_n2118) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1181 ( .A1(DP_OP_422J2_124_3477_n1958), 
        .A2(DP_OP_422J2_124_3477_n1962), .Y(DP_OP_422J2_124_3477_n1942) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1257 ( .A1(DP_OP_423J2_125_3477_n2878), 
        .A2(DP_OP_422J2_124_3477_n2049), .Y(DP_OP_422J2_124_3477_n2018) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2026 ( .A1(DP_OP_423J2_125_3477_n2795), 
        .A2(DP_OP_422J2_124_3477_n2799), .Y(DP_OP_423J2_125_3477_n2787) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1406 ( .A1(DP_OP_425J2_127_3477_n2307), 
        .A2(DP_OP_422J2_124_3477_n2183), .Y(DP_OP_422J2_124_3477_n2167) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2015 ( .A1(DP_OP_422J2_124_3477_n2792), 
        .A2(DP_OP_422J2_124_3477_n2798), .Y(DP_OP_422J2_124_3477_n2776) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1214 ( .A1(DP_OP_423J2_125_3477_n2923), 
        .A2(DP_OP_422J2_124_3477_n2005), .Y(DP_OP_422J2_124_3477_n1975) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1394 ( .A1(DP_OP_422J2_124_3477_n2179), 
        .A2(DP_OP_422J2_124_3477_n2181), .Y(DP_OP_422J2_124_3477_n2155) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1218 ( .A1(DP_OP_425J2_127_3477_n2135), 
        .A2(DP_OP_422J2_124_3477_n2005), .Y(DP_OP_422J2_124_3477_n1979) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1844 ( .A1(DP_OP_422J2_124_3477_n2613), 
        .A2(DP_OP_422J2_124_3477_n2623), .Y(DP_OP_422J2_124_3477_n2605) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1848 ( .A1(DP_OP_422J2_124_3477_n2617), 
        .A2(DP_OP_422J2_124_3477_n2623), .Y(DP_OP_422J2_124_3477_n2609) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1522 ( .A1(DP_OP_422J2_124_3477_n2307), 
        .A2(DP_OP_422J2_124_3477_n2313), .Y(DP_OP_422J2_124_3477_n2283) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2056 ( .A1(DP_OP_422J2_124_3477_n2833), 
        .A2(DP_OP_422J2_124_3477_n2842), .Y(DP_OP_422J2_124_3477_n2817) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2105 ( .A1(DP_OP_425J2_127_3477_n2750), 
        .A2(DP_OP_422J2_124_3477_n2886), .Y(DP_OP_422J2_124_3477_n2866) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2202 ( .A1(DP_OP_423J2_125_3477_n2971), 
        .A2(DP_OP_422J2_124_3477_n2975), .Y(DP_OP_423J2_125_3477_n2963) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2147 ( .A1(DP_OP_422J2_124_3477_n2924), 
        .A2(DP_OP_422J2_124_3477_n2930), .Y(DP_OP_422J2_124_3477_n2908) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1759 ( .A1(DP_OP_422J2_124_3477_n2528), 
        .A2(DP_OP_422J2_124_3477_n2535), .Y(DP_OP_422J2_124_3477_n2520) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1301 ( .A1(DP_OP_423J2_125_3477_n2834), 
        .A2(DP_OP_422J2_124_3477_n2093), .Y(DP_OP_422J2_124_3477_n2062) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2237 ( .A1(DP_OP_422J2_124_3477_n3012), 
        .A2(DP_OP_422J2_124_3477_n3016), .Y(DP_OP_422J2_124_3477_n2996) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2154 ( .A1(DP_OP_422J2_124_3477_n2923), 
        .A2(DP_OP_422J2_124_3477_n2931), .Y(DP_OP_422J2_124_3477_n2915) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2138 ( .A1(DP_OP_422J2_124_3477_n2923), 
        .A2(DP_OP_422J2_124_3477_n2929), .Y(DP_OP_422J2_124_3477_n2899) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1610 ( .A1(DP_OP_423J2_125_3477_n2527), 
        .A2(DP_OP_422J2_124_3477_n2401), .Y(DP_OP_422J2_124_3477_n2371) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1891 ( .A1(DP_OP_425J2_127_3477_n2528), 
        .A2(DP_OP_422J2_124_3477_n2667), .Y(DP_OP_422J2_124_3477_n2652) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1574 ( .A1(DP_OP_422J2_124_3477_n2351), 
        .A2(DP_OP_422J2_124_3477_n2358), .Y(DP_OP_422J2_124_3477_n2335) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1566 ( .A1(DP_OP_422J2_124_3477_n2351), 
        .A2(DP_OP_422J2_124_3477_n2357), .Y(DP_OP_422J2_124_3477_n2327) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2016 ( .A1(DP_OP_422J2_124_3477_n2793), 
        .A2(DP_OP_422J2_124_3477_n2798), .Y(DP_OP_422J2_124_3477_n2777) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1582 ( .A1(DP_OP_422J2_124_3477_n2351), 
        .A2(DP_OP_422J2_124_3477_n2359), .Y(DP_OP_422J2_124_3477_n2343) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1584 ( .A1(DP_OP_422J2_124_3477_n2353), 
        .A2(DP_OP_422J2_124_3477_n2359), .Y(DP_OP_422J2_124_3477_n2345) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1796 ( .A1(DP_OP_423J2_125_3477_n2397), 
        .A2(DP_OP_422J2_124_3477_n2578), .Y(DP_OP_422J2_124_3477_n2557) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1624 ( .A1(DP_OP_423J2_125_3477_n2525), 
        .A2(DP_OP_422J2_124_3477_n2403), .Y(DP_OP_422J2_124_3477_n2385) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1577 ( .A1(DP_OP_422J2_124_3477_n2354), 
        .A2(DP_OP_422J2_124_3477_n2358), .Y(DP_OP_422J2_124_3477_n2338) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1878 ( .A1(DP_OP_422J2_124_3477_n2663), 
        .A2(DP_OP_423J2_125_3477_n2665), .Y(DP_OP_422J2_124_3477_n2639) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2184 ( .A1(DP_OP_422J2_124_3477_n2969), 
        .A2(DP_OP_422J2_124_3477_n2973), .Y(DP_OP_422J2_124_3477_n2945) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1170 ( .A1(DP_OP_423J2_125_3477_n2967), 
        .A2(DP_OP_422J2_124_3477_n1961), .Y(DP_OP_422J2_124_3477_n1931) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2191 ( .A1(DP_OP_423J2_125_3477_n2000), 
        .A2(DP_OP_422J2_124_3477_n2974), .Y(DP_OP_422J2_124_3477_n2952) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1580 ( .A1(DP_OP_424J2_126_3477_n2481), 
        .A2(DP_OP_422J2_124_3477_n2359), .Y(DP_OP_422J2_124_3477_n2341) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2244 ( .A1(DP_OP_422J2_124_3477_n3011), 
        .A2(DP_OP_422J2_124_3477_n3017), .Y(DP_OP_422J2_124_3477_n3003) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1614 ( .A1(DP_OP_423J2_125_3477_n2531), 
        .A2(DP_OP_422J2_124_3477_n2401), .Y(DP_OP_422J2_124_3477_n2375) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1173 ( .A1(DP_OP_422J2_124_3477_n1958), 
        .A2(DP_OP_422J2_124_3477_n1961), .Y(DP_OP_422J2_124_3477_n1934) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2190 ( .A1(DP_OP_424J2_126_3477_n2087), 
        .A2(DP_OP_422J2_124_3477_n2974), .Y(DP_OP_422J2_124_3477_n2951) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1962 ( .A1(DP_OP_422J2_124_3477_n2747), 
        .A2(DP_OP_422J2_124_3477_n2753), .Y(DP_OP_422J2_124_3477_n2723) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2246 ( .A1(DP_OP_425J2_127_3477_n2047), 
        .A2(DP_OP_423J2_125_3477_n3017), .Y(DP_OP_423J2_125_3477_n3005) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1481 ( .A1(DP_OP_425J2_127_3477_n2398), 
        .A2(DP_OP_422J2_124_3477_n2269), .Y(DP_OP_422J2_124_3477_n2242) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1628 ( .A1(DP_OP_423J2_125_3477_n2529), 
        .A2(DP_OP_422J2_124_3477_n2403), .Y(DP_OP_422J2_124_3477_n2389) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1709 ( .A1(DP_OP_422J2_124_3477_n2486), 
        .A2(DP_OP_422J2_124_3477_n2490), .Y(DP_OP_422J2_124_3477_n2470) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1434 ( .A1(DP_OP_422J2_124_3477_n2219), 
        .A2(DP_OP_422J2_124_3477_n2225), .Y(DP_OP_422J2_124_3477_n2195) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1753 ( .A1(DP_OP_423J2_125_3477_n2442), 
        .A2(DP_OP_422J2_124_3477_n2534), .Y(DP_OP_422J2_124_3477_n2514) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1929 ( .A1(DP_OP_424J2_126_3477_n2354), 
        .A2(DP_OP_422J2_124_3477_n2710), .Y(DP_OP_422J2_124_3477_n2690) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1565 ( .A1(DP_OP_424J2_126_3477_n2482), 
        .A2(DP_OP_422J2_124_3477_n2357), .Y(DP_OP_422J2_124_3477_n2326) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1621 ( .A1(DP_OP_423J2_125_3477_n2530), 
        .A2(DP_OP_425J2_127_3477_n2402), .Y(DP_OP_422J2_124_3477_n2382) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1927 ( .A1(DP_OP_422J2_124_3477_n2704), 
        .A2(DP_OP_422J2_124_3477_n2710), .Y(DP_OP_422J2_124_3477_n2688) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2183 ( .A1(DP_OP_423J2_125_3477_n2000), 
        .A2(DP_OP_422J2_124_3477_n2973), .Y(DP_OP_422J2_124_3477_n2944) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1918 ( .A1(DP_OP_424J2_126_3477_n2351), 
        .A2(DP_OP_422J2_124_3477_n2709), .Y(DP_OP_422J2_124_3477_n2679) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1707 ( .A1(DP_OP_422J2_124_3477_n2484), 
        .A2(DP_OP_422J2_124_3477_n2490), .Y(DP_OP_422J2_124_3477_n2468) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1705 ( .A1(DP_OP_422J2_124_3477_n2482), 
        .A2(DP_OP_422J2_124_3477_n2490), .Y(DP_OP_422J2_124_3477_n2466) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1934 ( .A1(DP_OP_424J2_126_3477_n2351), 
        .A2(DP_OP_422J2_124_3477_n2711), .Y(DP_OP_422J2_124_3477_n2695) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2156 ( .A1(DP_OP_424J2_126_3477_n2133), 
        .A2(DP_OP_422J2_124_3477_n2931), .Y(DP_OP_422J2_124_3477_n2917) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1745 ( .A1(DP_OP_423J2_125_3477_n2442), 
        .A2(DP_OP_422J2_124_3477_n2533), .Y(DP_OP_422J2_124_3477_n2506) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1921 ( .A1(DP_OP_424J2_126_3477_n2354), 
        .A2(DP_OP_422J2_124_3477_n2709), .Y(DP_OP_422J2_124_3477_n2682) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1712 ( .A1(DP_OP_422J2_124_3477_n2481), 
        .A2(DP_OP_422J2_124_3477_n2491), .Y(DP_OP_422J2_124_3477_n2473) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1612 ( .A1(DP_OP_423J2_125_3477_n2529), 
        .A2(DP_OP_422J2_124_3477_n2401), .Y(DP_OP_422J2_124_3477_n2373) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1702 ( .A1(DP_OP_422J2_124_3477_n2487), 
        .A2(DP_OP_422J2_124_3477_n2489), .Y(DP_OP_422J2_124_3477_n2463) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1881 ( .A1(DP_OP_422J2_124_3477_n2658), 
        .A2(DP_OP_422J2_124_3477_n2666), .Y(DP_OP_422J2_124_3477_n2642) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1356 ( .A1(DP_OP_424J2_126_3477_n2705), 
        .A2(DP_OP_422J2_124_3477_n2138), .Y(DP_OP_422J2_124_3477_n2117) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1348 ( .A1(DP_OP_424J2_126_3477_n2705), 
        .A2(DP_OP_422J2_124_3477_n2137), .Y(DP_OP_422J2_124_3477_n2109) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2137 ( .A1(DP_OP_422J2_124_3477_n2922), 
        .A2(DP_OP_422J2_124_3477_n2929), .Y(DP_OP_422J2_124_3477_n2898) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1451 ( .A1(DP_OP_422J2_124_3477_n2220), 
        .A2(DP_OP_422J2_124_3477_n2227), .Y(DP_OP_422J2_124_3477_n2212) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1698 ( .A1(DP_OP_422J2_124_3477_n2483), 
        .A2(DP_OP_422J2_124_3477_n2489), .Y(DP_OP_422J2_124_3477_n2459) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2066 ( .A1(DP_OP_422J2_124_3477_n2835), 
        .A2(DP_OP_422J2_124_3477_n2843), .Y(DP_OP_422J2_124_3477_n2827) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1874 ( .A1(DP_OP_422J2_124_3477_n2659), 
        .A2(DP_OP_424J2_126_3477_n2665), .Y(DP_OP_422J2_124_3477_n2635) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1663 ( .A1(DP_OP_423J2_125_3477_n2484), 
        .A2(DP_OP_422J2_124_3477_n2446), .Y(DP_OP_422J2_124_3477_n2424) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1925 ( .A1(DP_OP_422J2_124_3477_n2702), 
        .A2(DP_OP_422J2_124_3477_n2710), .Y(DP_OP_422J2_124_3477_n2686) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2059 ( .A1(DP_OP_425J2_127_3477_n2704), 
        .A2(DP_OP_422J2_124_3477_n2842), .Y(DP_OP_422J2_124_3477_n2820) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1220 ( .A1(DP_OP_424J2_126_3477_n2833), 
        .A2(DP_OP_422J2_124_3477_n2006), .Y(DP_OP_422J2_124_3477_n1981) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2192 ( .A1(DP_OP_422J2_124_3477_n2969), 
        .A2(DP_OP_422J2_124_3477_n2974), .Y(DP_OP_422J2_124_3477_n2953) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1213 ( .A1(DP_OP_424J2_126_3477_n2834), 
        .A2(DP_OP_422J2_124_3477_n2005), .Y(DP_OP_422J2_124_3477_n1974) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1850 ( .A1(DP_OP_423J2_125_3477_n2619), 
        .A2(DP_OP_423J2_125_3477_n2623), .Y(DP_OP_423J2_125_3477_n2611) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1922 ( .A1(DP_OP_422J2_124_3477_n2707), 
        .A2(DP_OP_422J2_124_3477_n2709), .Y(DP_OP_422J2_124_3477_n2683) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2052 ( .A1(DP_OP_422J2_124_3477_n2837), 
        .A2(DP_OP_422J2_124_3477_n2841), .Y(DP_OP_422J2_124_3477_n2813) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1258 ( .A1(DP_OP_424J2_126_3477_n2791), 
        .A2(DP_OP_422J2_124_3477_n2049), .Y(DP_OP_422J2_124_3477_n2019) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1794 ( .A1(DP_OP_422J2_124_3477_n2571), 
        .A2(DP_OP_422J2_124_3477_n2578), .Y(DP_OP_422J2_124_3477_n2555) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1438 ( .A1(DP_OP_425J2_127_3477_n2355), 
        .A2(DP_OP_422J2_124_3477_n2225), .Y(DP_OP_422J2_124_3477_n2199) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1936 ( .A1(DP_OP_424J2_126_3477_n2353), 
        .A2(DP_OP_422J2_124_3477_n2711), .Y(DP_OP_422J2_124_3477_n2697) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1222 ( .A1(DP_OP_424J2_126_3477_n2835), 
        .A2(DP_OP_422J2_124_3477_n2006), .Y(DP_OP_422J2_124_3477_n1983) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1917 ( .A1(DP_OP_422J2_124_3477_n2702), 
        .A2(DP_OP_422J2_124_3477_n2709), .Y(DP_OP_422J2_124_3477_n2678) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1661 ( .A1(DP_OP_423J2_125_3477_n2482), 
        .A2(DP_OP_422J2_124_3477_n2446), .Y(DP_OP_422J2_124_3477_n2422) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2065 ( .A1(DP_OP_422J2_124_3477_n2834), 
        .A2(DP_OP_422J2_124_3477_n2843), .Y(DP_OP_422J2_124_3477_n2826) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1762 ( .A1(DP_OP_423J2_125_3477_n2531), 
        .A2(DP_OP_423J2_125_3477_n2535), .Y(DP_OP_423J2_125_3477_n2523) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2141 ( .A1(DP_OP_422J2_124_3477_n2926), 
        .A2(DP_OP_422J2_124_3477_n2929), .Y(DP_OP_422J2_124_3477_n2902) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1966 ( .A1(DP_OP_422J2_124_3477_n2751), 
        .A2(DP_OP_422J2_124_3477_n2753), .Y(DP_OP_422J2_124_3477_n2727) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1567 ( .A1(DP_OP_424J2_126_3477_n2484), 
        .A2(DP_OP_422J2_124_3477_n2357), .Y(DP_OP_422J2_124_3477_n2328) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1716 ( .A1(DP_OP_422J2_124_3477_n2485), 
        .A2(DP_OP_422J2_124_3477_n2491), .Y(DP_OP_422J2_124_3477_n2477) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2024 ( .A1(DP_OP_422J2_124_3477_n2793), 
        .A2(DP_OP_422J2_124_3477_n2799), .Y(DP_OP_422J2_124_3477_n2785) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1268 ( .A1(DP_OP_422J2_124_3477_n2045), 
        .A2(DP_OP_422J2_124_3477_n2050), .Y(DP_OP_422J2_124_3477_n2029) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1609 ( .A1(DP_OP_423J2_125_3477_n2526), 
        .A2(DP_OP_422J2_124_3477_n2401), .Y(DP_OP_422J2_124_3477_n2370) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1354 ( .A1(DP_OP_424J2_126_3477_n2703), 
        .A2(DP_OP_422J2_124_3477_n2138), .Y(DP_OP_422J2_124_3477_n2115) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2189 ( .A1(DP_OP_423J2_125_3477_n1998), 
        .A2(DP_OP_422J2_124_3477_n2974), .Y(DP_OP_422J2_124_3477_n2950) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1223 ( .A1(DP_OP_422J2_124_3477_n2000), 
        .A2(DP_OP_422J2_124_3477_n2006), .Y(DP_OP_422J2_124_3477_n1984) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2139 ( .A1(DP_OP_422J2_124_3477_n2924), 
        .A2(DP_OP_422J2_124_3477_n2929), .Y(DP_OP_422J2_124_3477_n2900) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1347 ( .A1(DP_OP_422J2_124_3477_n2132), 
        .A2(DP_OP_422J2_124_3477_n2137), .Y(DP_OP_422J2_124_3477_n2108) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2185 ( .A1(DP_OP_422J2_124_3477_n2970), 
        .A2(DP_OP_422J2_124_3477_n2973), .Y(DP_OP_422J2_124_3477_n2946) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2021 ( .A1(DP_OP_422J2_124_3477_n2790), 
        .A2(DP_OP_422J2_124_3477_n2799), .Y(DP_OP_422J2_124_3477_n2782) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2193 ( .A1(DP_OP_422J2_124_3477_n2970), 
        .A2(DP_OP_422J2_124_3477_n2974), .Y(DP_OP_422J2_124_3477_n2954) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2235 ( .A1(DP_OP_422J2_124_3477_n3010), 
        .A2(DP_OP_422J2_124_3477_n3016), .Y(DP_OP_422J2_124_3477_n2994) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2226 ( .A1(DP_OP_422J2_124_3477_n3009), 
        .A2(DP_OP_422J2_124_3477_n3015), .Y(DP_OP_422J2_124_3477_n2985) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1626 ( .A1(DP_OP_423J2_125_3477_n2527), 
        .A2(DP_OP_422J2_124_3477_n2403), .Y(DP_OP_422J2_124_3477_n2387) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1266 ( .A1(DP_OP_424J2_126_3477_n2791), 
        .A2(DP_OP_422J2_124_3477_n2050), .Y(DP_OP_422J2_124_3477_n2027) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1401 ( .A1(DP_OP_422J2_124_3477_n2178), 
        .A2(DP_OP_422J2_124_3477_n2182), .Y(DP_OP_422J2_124_3477_n2162) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1935 ( .A1(DP_OP_422J2_124_3477_n2704), 
        .A2(DP_OP_422J2_124_3477_n2711), .Y(DP_OP_422J2_124_3477_n2696) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1259 ( .A1(DP_OP_422J2_124_3477_n2044), 
        .A2(DP_OP_422J2_124_3477_n2049), .Y(DP_OP_422J2_124_3477_n2020) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2233 ( .A1(DP_OP_422J2_124_3477_n3008), 
        .A2(DP_OP_422J2_124_3477_n3016), .Y(DP_OP_422J2_124_3477_n2992) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1216 ( .A1(DP_OP_424J2_126_3477_n2837), 
        .A2(DP_OP_422J2_124_3477_n2005), .Y(DP_OP_422J2_124_3477_n1977) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2049 ( .A1(DP_OP_422J2_124_3477_n2834), 
        .A2(DP_OP_425J2_127_3477_n2841), .Y(DP_OP_422J2_124_3477_n2810) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1486 ( .A1(DP_OP_422J2_124_3477_n2263), 
        .A2(DP_OP_422J2_124_3477_n2270), .Y(DP_OP_422J2_124_3477_n2247) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1965 ( .A1(DP_OP_422J2_124_3477_n2750), 
        .A2(DP_OP_422J2_124_3477_n2753), .Y(DP_OP_422J2_124_3477_n2726) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1345 ( .A1(DP_OP_422J2_124_3477_n2130), 
        .A2(DP_OP_422J2_124_3477_n2137), .Y(DP_OP_422J2_124_3477_n2106) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1706 ( .A1(DP_OP_422J2_124_3477_n2483), 
        .A2(DP_OP_422J2_124_3477_n2490), .Y(DP_OP_422J2_124_3477_n2467) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1353 ( .A1(DP_OP_422J2_124_3477_n2130), 
        .A2(DP_OP_422J2_124_3477_n2138), .Y(DP_OP_422J2_124_3477_n2114) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2017 ( .A1(DP_OP_423J2_125_3477_n2178), 
        .A2(DP_OP_422J2_124_3477_n2798), .Y(DP_OP_422J2_124_3477_n2778) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1699 ( .A1(DP_OP_422J2_124_3477_n2484), 
        .A2(DP_OP_422J2_124_3477_n2489), .Y(DP_OP_422J2_124_3477_n2460) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2242 ( .A1(DP_OP_422J2_124_3477_n3009), 
        .A2(DP_OP_422J2_124_3477_n3017), .Y(DP_OP_422J2_124_3477_n3001) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2013 ( .A1(DP_OP_422J2_124_3477_n2790), 
        .A2(DP_OP_422J2_124_3477_n2798), .Y(DP_OP_422J2_124_3477_n2774) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1933 ( .A1(DP_OP_422J2_124_3477_n2702), 
        .A2(DP_OP_422J2_124_3477_n2711), .Y(DP_OP_422J2_124_3477_n2694) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1352 ( .A1(DP_OP_422J2_124_3477_n2129), 
        .A2(DP_OP_422J2_124_3477_n2138), .Y(DP_OP_422J2_124_3477_n2113) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1847 ( .A1(DP_OP_422J2_124_3477_n2616), 
        .A2(DP_OP_422J2_124_3477_n2623), .Y(DP_OP_422J2_124_3477_n2608) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1454 ( .A1(DP_OP_422J2_124_3477_n2751), 
        .A2(DP_OP_425J2_127_3477_n2227), .Y(DP_OP_423J2_125_3477_n2215) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1399 ( .A1(DP_OP_423J2_125_3477_n2748), 
        .A2(DP_OP_422J2_124_3477_n2182), .Y(DP_OP_422J2_124_3477_n2160) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1410 ( .A1(DP_OP_425J2_127_3477_n2663), 
        .A2(DP_OP_423J2_125_3477_n2183), .Y(DP_OP_423J2_125_3477_n2171) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2068 ( .A1(DP_OP_422J2_124_3477_n2837), 
        .A2(DP_OP_422J2_124_3477_n2843), .Y(DP_OP_422J2_124_3477_n2829) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2158 ( .A1(DP_OP_423J2_125_3477_n2927), 
        .A2(DP_OP_423J2_125_3477_n2931), .Y(DP_OP_423J2_125_3477_n2919) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1746 ( .A1(DP_OP_422J2_124_3477_n2531), 
        .A2(DP_OP_422J2_124_3477_n2533), .Y(DP_OP_422J2_124_3477_n2507) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1392 ( .A1(DP_OP_422J2_124_3477_n2177), 
        .A2(DP_OP_422J2_124_3477_n2181), .Y(DP_OP_422J2_124_3477_n2153) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2051 ( .A1(DP_OP_425J2_127_3477_n2704), 
        .A2(DP_OP_424J2_126_3477_n2841), .Y(DP_OP_422J2_124_3477_n2812) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1479 ( .A1(DP_OP_425J2_127_3477_n2396), 
        .A2(DP_OP_422J2_124_3477_n2269), .Y(DP_OP_422J2_124_3477_n2240) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1408 ( .A1(DP_OP_422J2_124_3477_n2177), 
        .A2(DP_OP_422J2_124_3477_n2183), .Y(DP_OP_422J2_124_3477_n2169) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1795 ( .A1(DP_OP_423J2_125_3477_n2396), 
        .A2(DP_OP_422J2_124_3477_n2578), .Y(DP_OP_422J2_124_3477_n2556) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2057 ( .A1(DP_OP_422J2_124_3477_n2834), 
        .A2(DP_OP_422J2_124_3477_n2842), .Y(DP_OP_422J2_124_3477_n2818) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1303 ( .A1(DP_OP_422J2_124_3477_n2088), 
        .A2(DP_OP_422J2_124_3477_n2093), .Y(DP_OP_422J2_124_3477_n2064) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1234 ( .A1(DP_OP_425J2_127_3477_n2135), 
        .A2(DP_OP_422J2_124_3477_n2007), .Y(DP_OP_422J2_124_3477_n1995) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1928 ( .A1(DP_OP_424J2_126_3477_n2353), 
        .A2(DP_OP_422J2_124_3477_n2710), .Y(DP_OP_422J2_124_3477_n2689) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1433 ( .A1(DP_OP_422J2_124_3477_n2218), 
        .A2(DP_OP_422J2_124_3477_n2225), .Y(DP_OP_422J2_124_3477_n2194) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2058 ( .A1(DP_OP_422J2_124_3477_n2835), 
        .A2(DP_OP_422J2_124_3477_n2842), .Y(DP_OP_422J2_124_3477_n2819) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2067 ( .A1(DP_OP_424J2_126_3477_n2220), 
        .A2(DP_OP_422J2_124_3477_n2843), .Y(DP_OP_422J2_124_3477_n2828) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1478 ( .A1(DP_OP_422J2_124_3477_n2263), 
        .A2(DP_OP_422J2_124_3477_n2269), .Y(DP_OP_422J2_124_3477_n2239) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1350 ( .A1(DP_OP_422J2_124_3477_n2135), 
        .A2(DP_OP_422J2_124_3477_n2137), .Y(DP_OP_422J2_124_3477_n2111) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1751 ( .A1(DP_OP_422J2_124_3477_n2528), 
        .A2(DP_OP_422J2_124_3477_n2534), .Y(DP_OP_422J2_124_3477_n2512) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2012 ( .A1(DP_OP_422J2_124_3477_n2789), 
        .A2(DP_OP_422J2_124_3477_n2798), .Y(DP_OP_422J2_124_3477_n2773) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1714 ( .A1(DP_OP_422J2_124_3477_n2483), 
        .A2(DP_OP_422J2_124_3477_n2491), .Y(DP_OP_422J2_124_3477_n2475) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1620 ( .A1(DP_OP_423J2_125_3477_n2529), 
        .A2(DP_OP_425J2_127_3477_n2402), .Y(DP_OP_422J2_124_3477_n2381) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2023 ( .A1(DP_OP_422J2_124_3477_n2792), 
        .A2(DP_OP_422J2_124_3477_n2799), .Y(DP_OP_422J2_124_3477_n2784) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1302 ( .A1(DP_OP_425J2_127_3477_n2219), 
        .A2(DP_OP_422J2_124_3477_n2093), .Y(DP_OP_422J2_124_3477_n2063) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1174 ( .A1(DP_OP_424J2_126_3477_n2883), 
        .A2(DP_OP_422J2_124_3477_n1961), .Y(DP_OP_422J2_124_3477_n1935) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1832 ( .A1(DP_OP_422J2_124_3477_n2617), 
        .A2(DP_OP_422J2_124_3477_n2621), .Y(DP_OP_422J2_124_3477_n2593) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1437 ( .A1(DP_OP_425J2_127_3477_n2354), 
        .A2(DP_OP_422J2_124_3477_n2225), .Y(DP_OP_422J2_124_3477_n2198) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1389 ( .A1(DP_OP_424J2_126_3477_n2658), 
        .A2(DP_OP_422J2_124_3477_n2181), .Y(DP_OP_422J2_124_3477_n2150) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1221 ( .A1(DP_OP_424J2_126_3477_n2834), 
        .A2(DP_OP_422J2_124_3477_n2006), .Y(DP_OP_422J2_124_3477_n1982) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2054 ( .A1(DP_OP_425J2_127_3477_n2707), 
        .A2(DP_OP_422J2_124_3477_n2841), .Y(DP_OP_422J2_124_3477_n2815) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2227 ( .A1(DP_OP_422J2_124_3477_n3010), 
        .A2(DP_OP_422J2_124_3477_n3015), .Y(DP_OP_422J2_124_3477_n2986) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2149 ( .A1(DP_OP_422J2_124_3477_n2926), 
        .A2(DP_OP_422J2_124_3477_n2930), .Y(DP_OP_422J2_124_3477_n2910) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1583 ( .A1(DP_OP_424J2_126_3477_n2484), 
        .A2(DP_OP_422J2_124_3477_n2359), .Y(DP_OP_422J2_124_3477_n2344) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2140 ( .A1(DP_OP_424J2_126_3477_n2133), 
        .A2(DP_OP_422J2_124_3477_n2929), .Y(DP_OP_422J2_124_3477_n2901) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1576 ( .A1(DP_OP_422J2_124_3477_n2353), 
        .A2(DP_OP_422J2_124_3477_n2358), .Y(DP_OP_422J2_124_3477_n2337) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2061 ( .A1(DP_OP_422J2_124_3477_n2838), 
        .A2(DP_OP_422J2_124_3477_n2842), .Y(DP_OP_422J2_124_3477_n2822) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1396 ( .A1(DP_OP_425J2_127_3477_n2305), 
        .A2(DP_OP_422J2_124_3477_n2182), .Y(DP_OP_422J2_124_3477_n2157) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2243 ( .A1(DP_OP_422J2_124_3477_n3010), 
        .A2(DP_OP_422J2_124_3477_n3017), .Y(DP_OP_422J2_124_3477_n3002) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1485 ( .A1(DP_OP_422J2_124_3477_n2262), 
        .A2(DP_OP_422J2_124_3477_n2270), .Y(DP_OP_422J2_124_3477_n2246) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2050 ( .A1(DP_OP_422J2_124_3477_n2835), 
        .A2(DP_OP_422J2_124_3477_n2841), .Y(DP_OP_422J2_124_3477_n2811) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2114 ( .A1(DP_OP_424J2_126_3477_n2795), 
        .A2(DP_OP_425J2_127_3477_n2887), .Y(DP_OP_423J2_125_3477_n2875) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1749 ( .A1(DP_OP_422J2_124_3477_n2526), 
        .A2(DP_OP_422J2_124_3477_n2534), .Y(DP_OP_422J2_124_3477_n2510) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1180 ( .A1(DP_OP_422J2_124_3477_n1957), 
        .A2(DP_OP_422J2_124_3477_n1962), .Y(DP_OP_422J2_124_3477_n1941) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1231 ( .A1(DP_OP_422J2_124_3477_n2000), 
        .A2(DP_OP_422J2_124_3477_n2007), .Y(DP_OP_422J2_124_3477_n1992) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1357 ( .A1(DP_OP_422J2_124_3477_n2926), 
        .A2(DP_OP_422J2_124_3477_n2138), .Y(DP_OP_424J2_126_3477_n2118) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1394 ( .A1(DP_OP_424J2_126_3477_n2179), 
        .A2(DP_OP_423J2_125_3477_n2181), .Y(DP_OP_424J2_126_3477_n2155) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1878 ( .A1(DP_OP_424J2_126_3477_n2663), 
        .A2(DP_OP_424J2_126_3477_n2665), .Y(DP_OP_424J2_126_3477_n2639) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1753 ( .A1(DP_OP_424J2_126_3477_n2530), 
        .A2(DP_OP_422J2_124_3477_n2534), .Y(DP_OP_424J2_126_3477_n2514) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2156 ( .A1(DP_OP_424J2_126_3477_n2925), 
        .A2(DP_OP_425J2_127_3477_n2931), .Y(DP_OP_424J2_126_3477_n2917) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2105 ( .A1(DP_OP_423J2_125_3477_n2970), 
        .A2(DP_OP_424J2_126_3477_n2886), .Y(DP_OP_424J2_126_3477_n2866) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2142 ( .A1(DP_OP_424J2_126_3477_n2927), 
        .A2(DP_OP_424J2_126_3477_n2929), .Y(DP_OP_424J2_126_3477_n2903) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2067 ( .A1(DP_OP_425J2_127_3477_n2220), 
        .A2(DP_OP_423J2_125_3477_n2843), .Y(DP_OP_423J2_125_3477_n2828) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1797 ( .A1(DP_OP_423J2_125_3477_n2662), 
        .A2(DP_OP_424J2_126_3477_n2578), .Y(DP_OP_424J2_126_3477_n2558) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1452 ( .A1(DP_OP_425J2_127_3477_n2705), 
        .A2(DP_OP_424J2_126_3477_n2227), .Y(DP_OP_424J2_126_3477_n2213) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1482 ( .A1(DP_OP_422J2_124_3477_n2795), 
        .A2(DP_OP_424J2_126_3477_n2269), .Y(DP_OP_424J2_126_3477_n2243) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1496 ( .A1(DP_OP_424J2_126_3477_n2265), 
        .A2(DP_OP_424J2_126_3477_n2271), .Y(DP_OP_424J2_126_3477_n2257) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1489 ( .A1(DP_OP_425J2_127_3477_n2662), 
        .A2(DP_OP_424J2_126_3477_n2270), .Y(DP_OP_424J2_126_3477_n2250) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1526 ( .A1(DP_OP_422J2_124_3477_n2751), 
        .A2(DP_OP_425J2_127_3477_n2313), .Y(DP_OP_424J2_126_3477_n2287) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2061 ( .A1(DP_OP_423J2_125_3477_n2926), 
        .A2(DP_OP_425J2_127_3477_n2842), .Y(DP_OP_424J2_126_3477_n2822) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2054 ( .A1(DP_OP_425J2_127_3477_n2135), 
        .A2(DP_OP_422J2_124_3477_n2841), .Y(DP_OP_424J2_126_3477_n2815) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1751 ( .A1(DP_OP_423J2_125_3477_n2528), 
        .A2(DP_OP_423J2_125_3477_n2534), .Y(DP_OP_423J2_125_3477_n2512) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1934 ( .A1(DP_OP_425J2_127_3477_n2351), 
        .A2(DP_OP_425J2_127_3477_n2711), .Y(DP_OP_423J2_125_3477_n2695) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2155 ( .A1(DP_OP_424J2_126_3477_n2924), 
        .A2(DP_OP_422J2_124_3477_n2931), .Y(DP_OP_424J2_126_3477_n2916) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1488 ( .A1(DP_OP_424J2_126_3477_n2265), 
        .A2(DP_OP_424J2_126_3477_n2270), .Y(DP_OP_424J2_126_3477_n2249) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1217 ( .A1(DP_OP_425J2_127_3477_n2926), 
        .A2(DP_OP_425J2_127_3477_n2005), .Y(DP_OP_424J2_126_3477_n1978) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1180 ( .A1(DP_OP_424J2_126_3477_n1957), 
        .A2(DP_OP_424J2_126_3477_n1962), .Y(DP_OP_424J2_126_3477_n1941) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1173 ( .A1(DP_OP_424J2_126_3477_n1958), 
        .A2(DP_OP_424J2_126_3477_n1961), .Y(DP_OP_424J2_126_3477_n1934) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1231 ( .A1(DP_OP_425J2_127_3477_n2924), 
        .A2(DP_OP_422J2_124_3477_n2007), .Y(DP_OP_424J2_126_3477_n1992) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1224 ( .A1(DP_OP_424J2_126_3477_n2001), 
        .A2(DP_OP_423J2_125_3477_n2006), .Y(DP_OP_424J2_126_3477_n1985) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1261 ( .A1(DP_OP_422J2_124_3477_n3012), 
        .A2(DP_OP_424J2_126_3477_n2049), .Y(DP_OP_424J2_126_3477_n2022) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1759 ( .A1(DP_OP_424J2_126_3477_n2528), 
        .A2(DP_OP_422J2_124_3477_n2535), .Y(DP_OP_424J2_126_3477_n2520) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1437 ( .A1(DP_OP_422J2_124_3477_n2750), 
        .A2(DP_OP_423J2_125_3477_n2225), .Y(DP_OP_423J2_125_3477_n2198) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2141 ( .A1(DP_OP_424J2_126_3477_n2926), 
        .A2(DP_OP_424J2_126_3477_n2929), .Y(DP_OP_424J2_126_3477_n2902) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2111 ( .A1(DP_OP_424J2_126_3477_n2880), 
        .A2(DP_OP_424J2_126_3477_n2887), .Y(DP_OP_424J2_126_3477_n2872) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2243 ( .A1(DP_OP_424J2_126_3477_n3010), 
        .A2(DP_OP_422J2_124_3477_n3017), .Y(DP_OP_424J2_126_3477_n3002) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1350 ( .A1(DP_OP_422J2_124_3477_n2927), 
        .A2(DP_OP_424J2_126_3477_n2137), .Y(DP_OP_424J2_126_3477_n2111) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1715 ( .A1(DP_OP_423J2_125_3477_n2484), 
        .A2(DP_OP_423J2_125_3477_n2491), .Y(DP_OP_423J2_125_3477_n2476) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1717 ( .A1(DP_OP_422J2_124_3477_n2354), 
        .A2(DP_OP_423J2_125_3477_n2491), .Y(DP_OP_424J2_126_3477_n2478) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1761 ( .A1(DP_OP_424J2_126_3477_n2530), 
        .A2(DP_OP_422J2_124_3477_n2535), .Y(DP_OP_424J2_126_3477_n2522) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1349 ( .A1(DP_OP_423J2_125_3477_n2134), 
        .A2(DP_OP_422J2_124_3477_n2137), .Y(DP_OP_423J2_125_3477_n2110) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2069 ( .A1(DP_OP_425J2_127_3477_n2134), 
        .A2(DP_OP_423J2_125_3477_n2843), .Y(DP_OP_424J2_126_3477_n2830) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1234 ( .A1(DP_OP_425J2_127_3477_n2927), 
        .A2(DP_OP_425J2_127_3477_n2007), .Y(DP_OP_424J2_126_3477_n1995) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2199 ( .A1(DP_OP_424J2_126_3477_n2880), 
        .A2(DP_OP_422J2_124_3477_n2975), .Y(DP_OP_423J2_125_3477_n2960) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2242 ( .A1(DP_OP_423J2_125_3477_n3009), 
        .A2(DP_OP_423J2_125_3477_n3017), .Y(DP_OP_423J2_125_3477_n3001) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1584 ( .A1(DP_OP_424J2_126_3477_n2353), 
        .A2(DP_OP_423J2_125_3477_n2359), .Y(DP_OP_424J2_126_3477_n2345) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1577 ( .A1(DP_OP_424J2_126_3477_n2354), 
        .A2(DP_OP_424J2_126_3477_n2358), .Y(DP_OP_424J2_126_3477_n2338) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1614 ( .A1(DP_OP_422J2_124_3477_n2663), 
        .A2(DP_OP_424J2_126_3477_n2401), .Y(DP_OP_424J2_126_3477_n2375) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1628 ( .A1(DP_OP_424J2_126_3477_n2397), 
        .A2(DP_OP_422J2_124_3477_n2403), .Y(DP_OP_424J2_126_3477_n2389) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1621 ( .A1(DP_OP_422J2_124_3477_n2662), 
        .A2(DP_OP_424J2_126_3477_n2402), .Y(DP_OP_424J2_126_3477_n2382) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1658 ( .A1(DP_OP_422J2_124_3477_n2619), 
        .A2(DP_OP_424J2_126_3477_n2445), .Y(DP_OP_424J2_126_3477_n2419) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1168 ( .A1(DP_OP_422J2_124_3477_n3007), 
        .A2(DP_OP_424J2_126_3477_n1961), .Y(DP_OP_423J2_125_3477_n1929) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1922 ( .A1(DP_OP_422J2_124_3477_n2135), 
        .A2(DP_OP_425J2_127_3477_n2709), .Y(DP_OP_424J2_126_3477_n2683) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1702 ( .A1(DP_OP_422J2_124_3477_n2355), 
        .A2(DP_OP_424J2_126_3477_n2489), .Y(DP_OP_424J2_126_3477_n2463) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1709 ( .A1(DP_OP_422J2_124_3477_n2354), 
        .A2(DP_OP_425J2_127_3477_n2490), .Y(DP_OP_424J2_126_3477_n2470) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1848 ( .A1(DP_OP_423J2_125_3477_n2705), 
        .A2(DP_OP_424J2_126_3477_n2623), .Y(DP_OP_424J2_126_3477_n2609) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1760 ( .A1(DP_OP_425J2_127_3477_n2441), 
        .A2(DP_OP_423J2_125_3477_n2535), .Y(DP_OP_424J2_126_3477_n2521) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2149 ( .A1(DP_OP_424J2_126_3477_n2926), 
        .A2(DP_OP_423J2_125_3477_n2930), .Y(DP_OP_424J2_126_3477_n2910) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1399 ( .A1(DP_OP_422J2_124_3477_n2792), 
        .A2(DP_OP_425J2_127_3477_n2182), .Y(DP_OP_423J2_125_3477_n2160) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1408 ( .A1(DP_OP_424J2_126_3477_n2177), 
        .A2(DP_OP_424J2_126_3477_n2183), .Y(DP_OP_424J2_126_3477_n2169) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1401 ( .A1(DP_OP_424J2_126_3477_n2178), 
        .A2(DP_OP_424J2_126_3477_n2182), .Y(DP_OP_424J2_126_3477_n2162) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1438 ( .A1(DP_OP_425J2_127_3477_n2707), 
        .A2(DP_OP_424J2_126_3477_n2225), .Y(DP_OP_424J2_126_3477_n2199) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1392 ( .A1(DP_OP_424J2_126_3477_n2265), 
        .A2(DP_OP_423J2_125_3477_n2181), .Y(DP_OP_423J2_125_3477_n2153) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2112 ( .A1(DP_OP_423J2_125_3477_n2969), 
        .A2(DP_OP_424J2_126_3477_n2887), .Y(DP_OP_424J2_126_3477_n2873) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1834 ( .A1(DP_OP_423J2_125_3477_n2707), 
        .A2(DP_OP_425J2_127_3477_n2621), .Y(DP_OP_424J2_126_3477_n2595) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1885 ( .A1(DP_OP_422J2_124_3477_n2178), 
        .A2(DP_OP_424J2_126_3477_n2666), .Y(DP_OP_424J2_126_3477_n2646) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2200 ( .A1(DP_OP_424J2_126_3477_n2969), 
        .A2(DP_OP_424J2_126_3477_n2975), .Y(DP_OP_424J2_126_3477_n2961) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1672 ( .A1(DP_OP_422J2_124_3477_n2617), 
        .A2(DP_OP_424J2_126_3477_n2447), .Y(DP_OP_424J2_126_3477_n2433) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1540 ( .A1(DP_OP_422J2_124_3477_n2749), 
        .A2(DP_OP_424J2_126_3477_n2315), .Y(DP_OP_424J2_126_3477_n2301) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1570 ( .A1(DP_OP_422J2_124_3477_n2707), 
        .A2(DP_OP_424J2_126_3477_n2357), .Y(DP_OP_424J2_126_3477_n2331) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1966 ( .A1(DP_OP_424J2_126_3477_n2751), 
        .A2(DP_OP_424J2_126_3477_n2753), .Y(DP_OP_424J2_126_3477_n2727) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1746 ( .A1(DP_OP_422J2_124_3477_n2311), 
        .A2(DP_OP_424J2_126_3477_n2533), .Y(DP_OP_424J2_126_3477_n2507) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2186 ( .A1(DP_OP_425J2_127_3477_n2003), 
        .A2(DP_OP_425J2_127_3477_n2973), .Y(DP_OP_424J2_126_3477_n2947) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1929 ( .A1(DP_OP_422J2_124_3477_n2134), 
        .A2(DP_OP_423J2_125_3477_n2710), .Y(DP_OP_424J2_126_3477_n2690) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2244 ( .A1(DP_OP_424J2_126_3477_n3011), 
        .A2(DP_OP_423J2_125_3477_n3017), .Y(DP_OP_424J2_126_3477_n3003) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2237 ( .A1(DP_OP_424J2_126_3477_n3012), 
        .A2(DP_OP_424J2_126_3477_n3016), .Y(DP_OP_424J2_126_3477_n2996) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1218 ( .A1(DP_OP_425J2_127_3477_n2927), 
        .A2(DP_OP_422J2_124_3477_n2005), .Y(DP_OP_424J2_126_3477_n1979) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1795 ( .A1(DP_OP_423J2_125_3477_n2572), 
        .A2(DP_OP_422J2_124_3477_n2578), .Y(DP_OP_423J2_125_3477_n2556) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1181 ( .A1(DP_OP_424J2_126_3477_n1958), 
        .A2(DP_OP_424J2_126_3477_n1962), .Y(DP_OP_424J2_126_3477_n1942) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1174 ( .A1(DP_OP_425J2_127_3477_n2971), 
        .A2(DP_OP_424J2_126_3477_n1961), .Y(DP_OP_424J2_126_3477_n1935) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2068 ( .A1(DP_OP_424J2_126_3477_n2837), 
        .A2(DP_OP_422J2_124_3477_n2843), .Y(DP_OP_424J2_126_3477_n2829) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2017 ( .A1(DP_OP_424J2_126_3477_n2794), 
        .A2(DP_OP_423J2_125_3477_n2798), .Y(DP_OP_424J2_126_3477_n2778) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2024 ( .A1(DP_OP_424J2_126_3477_n2793), 
        .A2(DP_OP_424J2_126_3477_n2799), .Y(DP_OP_424J2_126_3477_n2785) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1892 ( .A1(DP_OP_423J2_125_3477_n2749), 
        .A2(DP_OP_425J2_127_3477_n2667), .Y(DP_OP_424J2_126_3477_n2653) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1665 ( .A1(DP_OP_424J2_126_3477_n2442), 
        .A2(DP_OP_424J2_126_3477_n2446), .Y(DP_OP_424J2_126_3477_n2426) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2230 ( .A1(DP_OP_424J2_126_3477_n3013), 
        .A2(DP_OP_424J2_126_3477_n3015), .Y(DP_OP_424J2_126_3477_n2989) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1232 ( .A1(DP_OP_424J2_126_3477_n2001), 
        .A2(DP_OP_425J2_127_3477_n2007), .Y(DP_OP_424J2_126_3477_n1993) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1225 ( .A1(DP_OP_425J2_127_3477_n2926), 
        .A2(DP_OP_425J2_127_3477_n2006), .Y(DP_OP_424J2_126_3477_n1986) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1262 ( .A1(DP_OP_424J2_126_3477_n2047), 
        .A2(DP_OP_424J2_126_3477_n2049), .Y(DP_OP_424J2_126_3477_n2023) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1269 ( .A1(DP_OP_423J2_125_3477_n1958), 
        .A2(DP_OP_422J2_124_3477_n2050), .Y(DP_OP_424J2_126_3477_n2030) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1306 ( .A1(DP_OP_423J2_125_3477_n2003), 
        .A2(DP_OP_422J2_124_3477_n2093), .Y(DP_OP_424J2_126_3477_n2067) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1936 ( .A1(DP_OP_424J2_126_3477_n2705), 
        .A2(DP_OP_424J2_126_3477_n2711), .Y(DP_OP_424J2_126_3477_n2697) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1716 ( .A1(DP_OP_422J2_124_3477_n2353), 
        .A2(DP_OP_422J2_124_3477_n2491), .Y(DP_OP_424J2_126_3477_n2477) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2193 ( .A1(DP_OP_424J2_126_3477_n2970), 
        .A2(DP_OP_423J2_125_3477_n2974), .Y(DP_OP_424J2_126_3477_n2954) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1664 ( .A1(DP_OP_422J2_124_3477_n2617), 
        .A2(DP_OP_424J2_126_3477_n2446), .Y(DP_OP_424J2_126_3477_n2425) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1477 ( .A1(DP_OP_423J2_125_3477_n2262), 
        .A2(DP_OP_422J2_124_3477_n2269), .Y(DP_OP_423J2_125_3477_n2238) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1612 ( .A1(DP_OP_424J2_126_3477_n2397), 
        .A2(DP_OP_424J2_126_3477_n2401), .Y(DP_OP_424J2_126_3477_n2373) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1348 ( .A1(DP_OP_424J2_126_3477_n2133), 
        .A2(DP_OP_424J2_126_3477_n2137), .Y(DP_OP_424J2_126_3477_n2109) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2066 ( .A1(DP_OP_424J2_126_3477_n2835), 
        .A2(DP_OP_425J2_127_3477_n2843), .Y(DP_OP_424J2_126_3477_n2827) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1480 ( .A1(DP_OP_424J2_126_3477_n2265), 
        .A2(DP_OP_424J2_126_3477_n2269), .Y(DP_OP_424J2_126_3477_n2241) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1748 ( .A1(DP_OP_423J2_125_3477_n2525), 
        .A2(DP_OP_423J2_125_3477_n2534), .Y(DP_OP_423J2_125_3477_n2509) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1663 ( .A1(DP_OP_425J2_127_3477_n2484), 
        .A2(DP_OP_424J2_126_3477_n2446), .Y(DP_OP_424J2_126_3477_n2424) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2059 ( .A1(DP_OP_423J2_125_3477_n2924), 
        .A2(DP_OP_422J2_124_3477_n2842), .Y(DP_OP_424J2_126_3477_n2820) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2052 ( .A1(DP_OP_424J2_126_3477_n2837), 
        .A2(DP_OP_423J2_125_3477_n2841), .Y(DP_OP_424J2_126_3477_n2813) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1934 ( .A1(DP_OP_424J2_126_3477_n2703), 
        .A2(DP_OP_424J2_126_3477_n2711), .Y(DP_OP_424J2_126_3477_n2695) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1707 ( .A1(DP_OP_424J2_126_3477_n2484), 
        .A2(DP_OP_425J2_127_3477_n2490), .Y(DP_OP_424J2_126_3477_n2468) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1927 ( .A1(DP_OP_422J2_124_3477_n2132), 
        .A2(DP_OP_425J2_127_3477_n2710), .Y(DP_OP_424J2_126_3477_n2688) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1656 ( .A1(DP_OP_422J2_124_3477_n2617), 
        .A2(DP_OP_424J2_126_3477_n2445), .Y(DP_OP_424J2_126_3477_n2417) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2191 ( .A1(DP_OP_425J2_127_3477_n2000), 
        .A2(DP_OP_422J2_124_3477_n2974), .Y(DP_OP_424J2_126_3477_n2952) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2184 ( .A1(DP_OP_424J2_126_3477_n2969), 
        .A2(DP_OP_422J2_124_3477_n2973), .Y(DP_OP_424J2_126_3477_n2945) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1582 ( .A1(DP_OP_424J2_126_3477_n2351), 
        .A2(DP_OP_422J2_124_3477_n2359), .Y(DP_OP_424J2_126_3477_n2343) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2154 ( .A1(DP_OP_424J2_126_3477_n2923), 
        .A2(DP_OP_423J2_125_3477_n2931), .Y(DP_OP_424J2_126_3477_n2915) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2147 ( .A1(DP_OP_424J2_126_3477_n2924), 
        .A2(DP_OP_422J2_124_3477_n2930), .Y(DP_OP_424J2_126_3477_n2908) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2015 ( .A1(DP_OP_423J2_125_3477_n2880), 
        .A2(DP_OP_425J2_127_3477_n2798), .Y(DP_OP_424J2_126_3477_n2776) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1406 ( .A1(DP_OP_425J2_127_3477_n2747), 
        .A2(DP_OP_424J2_126_3477_n2183), .Y(DP_OP_424J2_126_3477_n2167) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1436 ( .A1(DP_OP_422J2_124_3477_n2837), 
        .A2(DP_OP_424J2_126_3477_n2225), .Y(DP_OP_424J2_126_3477_n2197) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1575 ( .A1(DP_OP_422J2_124_3477_n2704), 
        .A2(DP_OP_424J2_126_3477_n2358), .Y(DP_OP_424J2_126_3477_n2336) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1873 ( .A1(DP_OP_423J2_125_3477_n2658), 
        .A2(DP_OP_423J2_125_3477_n2665), .Y(DP_OP_423J2_125_3477_n2634) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2140 ( .A1(DP_OP_424J2_126_3477_n2925), 
        .A2(DP_OP_424J2_126_3477_n2929), .Y(DP_OP_424J2_126_3477_n2901) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1832 ( .A1(DP_OP_425J2_127_3477_n2353), 
        .A2(DP_OP_422J2_124_3477_n2621), .Y(DP_OP_424J2_126_3477_n2593) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1714 ( .A1(DP_OP_422J2_124_3477_n2351), 
        .A2(DP_OP_425J2_127_3477_n2491), .Y(DP_OP_424J2_126_3477_n2475) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1751 ( .A1(DP_OP_424J2_126_3477_n2528), 
        .A2(DP_OP_425J2_127_3477_n2534), .Y(DP_OP_424J2_126_3477_n2512) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1795 ( .A1(DP_OP_424J2_126_3477_n2572), 
        .A2(DP_OP_424J2_126_3477_n2578), .Y(DP_OP_424J2_126_3477_n2556) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1392 ( .A1(DP_OP_424J2_126_3477_n2177), 
        .A2(DP_OP_422J2_124_3477_n2181), .Y(DP_OP_424J2_126_3477_n2153) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1399 ( .A1(DP_OP_422J2_124_3477_n2880), 
        .A2(DP_OP_424J2_126_3477_n2182), .Y(DP_OP_424J2_126_3477_n2160) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2242 ( .A1(DP_OP_424J2_126_3477_n3009), 
        .A2(DP_OP_425J2_127_3477_n3017), .Y(DP_OP_424J2_126_3477_n3001) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1216 ( .A1(DP_OP_424J2_126_3477_n2001), 
        .A2(DP_OP_422J2_124_3477_n2005), .Y(DP_OP_424J2_126_3477_n1977) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1626 ( .A1(DP_OP_422J2_124_3477_n2659), 
        .A2(DP_OP_425J2_127_3477_n2403), .Y(DP_OP_424J2_126_3477_n2387) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2235 ( .A1(DP_OP_424J2_126_3477_n3010), 
        .A2(DP_OP_424J2_126_3477_n3016), .Y(DP_OP_424J2_126_3477_n2994) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1223 ( .A1(DP_OP_425J2_127_3477_n2924), 
        .A2(DP_OP_423J2_125_3477_n2006), .Y(DP_OP_424J2_126_3477_n1984) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1846 ( .A1(DP_OP_422J2_124_3477_n2219), 
        .A2(DP_OP_424J2_126_3477_n2623), .Y(DP_OP_424J2_126_3477_n2607) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1883 ( .A1(DP_OP_423J2_125_3477_n2748), 
        .A2(DP_OP_424J2_126_3477_n2666), .Y(DP_OP_424J2_126_3477_n2644) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1744 ( .A1(DP_OP_425J2_127_3477_n2441), 
        .A2(DP_OP_424J2_126_3477_n2533), .Y(DP_OP_424J2_126_3477_n2505) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1697 ( .A1(DP_OP_423J2_125_3477_n2482), 
        .A2(DP_OP_423J2_125_3477_n2489), .Y(DP_OP_423J2_125_3477_n2458) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1179 ( .A1(DP_OP_424J2_126_3477_n1956), 
        .A2(DP_OP_424J2_126_3477_n1962), .Y(DP_OP_424J2_126_3477_n1940) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1172 ( .A1(DP_OP_424J2_126_3477_n1957), 
        .A2(DP_OP_424J2_126_3477_n1961), .Y(DP_OP_424J2_126_3477_n1933) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1569 ( .A1(DP_OP_424J2_126_3477_n2354), 
        .A2(DP_OP_424J2_126_3477_n2357), .Y(DP_OP_424J2_126_3477_n2330) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2023 ( .A1(DP_OP_423J2_125_3477_n2880), 
        .A2(DP_OP_424J2_126_3477_n2799), .Y(DP_OP_424J2_126_3477_n2784) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1701 ( .A1(DP_OP_422J2_124_3477_n2354), 
        .A2(DP_OP_424J2_126_3477_n2489), .Y(DP_OP_424J2_126_3477_n2462) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1620 ( .A1(DP_OP_424J2_126_3477_n2397), 
        .A2(DP_OP_424J2_126_3477_n2402), .Y(DP_OP_424J2_126_3477_n2381) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1921 ( .A1(DP_OP_422J2_124_3477_n2134), 
        .A2(DP_OP_423J2_125_3477_n2709), .Y(DP_OP_424J2_126_3477_n2682) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1268 ( .A1(DP_OP_423J2_125_3477_n1957), 
        .A2(DP_OP_422J2_124_3477_n2050), .Y(DP_OP_424J2_126_3477_n2029) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1305 ( .A1(DP_OP_424J2_126_3477_n2090), 
        .A2(DP_OP_422J2_124_3477_n2093), .Y(DP_OP_424J2_126_3477_n2066) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1613 ( .A1(DP_OP_422J2_124_3477_n2662), 
        .A2(DP_OP_424J2_126_3477_n2401), .Y(DP_OP_424J2_126_3477_n2374) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1833 ( .A1(DP_OP_424J2_126_3477_n2618), 
        .A2(DP_OP_422J2_124_3477_n2621), .Y(DP_OP_424J2_126_3477_n2594) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1495 ( .A1(DP_OP_424J2_126_3477_n2264), 
        .A2(DP_OP_424J2_126_3477_n2271), .Y(DP_OP_424J2_126_3477_n2256) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2148 ( .A1(DP_OP_424J2_126_3477_n2925), 
        .A2(DP_OP_425J2_127_3477_n2930), .Y(DP_OP_424J2_126_3477_n2909) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1671 ( .A1(DP_OP_422J2_124_3477_n2616), 
        .A2(DP_OP_424J2_126_3477_n2447), .Y(DP_OP_424J2_126_3477_n2432) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2104 ( .A1(DP_OP_423J2_125_3477_n2969), 
        .A2(DP_OP_424J2_126_3477_n2886), .Y(DP_OP_424J2_126_3477_n2865) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1525 ( .A1(DP_OP_424J2_126_3477_n2310), 
        .A2(DP_OP_422J2_124_3477_n2313), .Y(DP_OP_424J2_126_3477_n2286) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1847 ( .A1(DP_OP_424J2_126_3477_n2616), 
        .A2(DP_OP_424J2_126_3477_n2623), .Y(DP_OP_424J2_126_3477_n2608) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1928 ( .A1(DP_OP_424J2_126_3477_n2705), 
        .A2(DP_OP_422J2_124_3477_n2710), .Y(DP_OP_424J2_126_3477_n2689) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1583 ( .A1(DP_OP_422J2_124_3477_n2704), 
        .A2(DP_OP_425J2_127_3477_n2359), .Y(DP_OP_424J2_126_3477_n2344) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1714 ( .A1(DP_OP_422J2_124_3477_n2439), 
        .A2(DP_OP_423J2_125_3477_n2491), .Y(DP_OP_423J2_125_3477_n2475) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1657 ( .A1(DP_OP_424J2_126_3477_n2442), 
        .A2(DP_OP_424J2_126_3477_n2445), .Y(DP_OP_424J2_126_3477_n2418) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2016 ( .A1(DP_OP_424J2_126_3477_n2793), 
        .A2(DP_OP_422J2_124_3477_n2798), .Y(DP_OP_424J2_126_3477_n2777) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1745 ( .A1(DP_OP_424J2_126_3477_n2530), 
        .A2(DP_OP_424J2_126_3477_n2533), .Y(DP_OP_424J2_126_3477_n2506) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1356 ( .A1(DP_OP_424J2_126_3477_n2133), 
        .A2(DP_OP_423J2_125_3477_n2138), .Y(DP_OP_424J2_126_3477_n2117) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2192 ( .A1(DP_OP_424J2_126_3477_n2969), 
        .A2(DP_OP_423J2_125_3477_n2974), .Y(DP_OP_424J2_126_3477_n2953) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1891 ( .A1(DP_OP_423J2_125_3477_n2748), 
        .A2(DP_OP_422J2_124_3477_n2667), .Y(DP_OP_424J2_126_3477_n2652) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1627 ( .A1(DP_OP_423J2_125_3477_n2308), 
        .A2(DP_OP_425J2_127_3477_n2403), .Y(DP_OP_424J2_126_3477_n2388) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1884 ( .A1(DP_OP_422J2_124_3477_n2177), 
        .A2(DP_OP_424J2_126_3477_n2666), .Y(DP_OP_424J2_126_3477_n2645) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1877 ( .A1(DP_OP_423J2_125_3477_n2750), 
        .A2(DP_OP_424J2_126_3477_n2665), .Y(DP_OP_424J2_126_3477_n2638) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1576 ( .A1(DP_OP_424J2_126_3477_n2353), 
        .A2(DP_OP_424J2_126_3477_n2358), .Y(DP_OP_424J2_126_3477_n2337) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1965 ( .A1(DP_OP_424J2_126_3477_n2750), 
        .A2(DP_OP_424J2_126_3477_n2753), .Y(DP_OP_424J2_126_3477_n2726) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1935 ( .A1(DP_OP_422J2_124_3477_n2132), 
        .A2(DP_OP_424J2_126_3477_n2711), .Y(DP_OP_424J2_126_3477_n2696) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2185 ( .A1(DP_OP_424J2_126_3477_n2970), 
        .A2(DP_OP_422J2_124_3477_n2973), .Y(DP_OP_424J2_126_3477_n2946) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1393 ( .A1(DP_OP_424J2_126_3477_n2178), 
        .A2(DP_OP_422J2_124_3477_n2181), .Y(DP_OP_424J2_126_3477_n2154) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1708 ( .A1(DP_OP_422J2_124_3477_n2353), 
        .A2(DP_OP_423J2_125_3477_n2490), .Y(DP_OP_424J2_126_3477_n2469) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1400 ( .A1(DP_OP_424J2_126_3477_n2177), 
        .A2(DP_OP_424J2_126_3477_n2182), .Y(DP_OP_424J2_126_3477_n2161) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1407 ( .A1(DP_OP_422J2_124_3477_n2880), 
        .A2(DP_OP_424J2_126_3477_n2183), .Y(DP_OP_424J2_126_3477_n2168) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2060 ( .A1(DP_OP_424J2_126_3477_n2837), 
        .A2(DP_OP_422J2_124_3477_n2842), .Y(DP_OP_424J2_126_3477_n2821) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2053 ( .A1(DP_OP_425J2_127_3477_n2134), 
        .A2(DP_OP_424J2_126_3477_n2841), .Y(DP_OP_424J2_126_3477_n2814) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1539 ( .A1(DP_OP_424J2_126_3477_n2308), 
        .A2(DP_OP_424J2_126_3477_n2315), .Y(DP_OP_424J2_126_3477_n2300) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1752 ( .A1(DP_OP_423J2_125_3477_n2617), 
        .A2(DP_OP_422J2_124_3477_n2534), .Y(DP_OP_424J2_126_3477_n2513) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2236 ( .A1(DP_OP_424J2_126_3477_n3011), 
        .A2(DP_OP_424J2_126_3477_n3016), .Y(DP_OP_424J2_126_3477_n2995) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1169 ( .A1(DP_OP_425J2_127_3477_n2878), 
        .A2(DP_OP_422J2_124_3477_n1961), .Y(DP_OP_423J2_125_3477_n1930) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2229 ( .A1(DP_OP_424J2_126_3477_n3012), 
        .A2(DP_OP_424J2_126_3477_n3015), .Y(DP_OP_424J2_126_3477_n2988) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1796 ( .A1(DP_OP_423J2_125_3477_n2573), 
        .A2(DP_OP_425J2_127_3477_n2578), .Y(DP_OP_423J2_125_3477_n2557) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1715 ( .A1(DP_OP_424J2_126_3477_n2484), 
        .A2(DP_OP_423J2_125_3477_n2491), .Y(DP_OP_424J2_126_3477_n2476) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1349 ( .A1(DP_OP_422J2_124_3477_n2926), 
        .A2(DP_OP_424J2_126_3477_n2137), .Y(DP_OP_424J2_126_3477_n2110) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2199 ( .A1(DP_OP_425J2_127_3477_n2000), 
        .A2(DP_OP_424J2_126_3477_n2975), .Y(DP_OP_424J2_126_3477_n2960) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1451 ( .A1(DP_OP_425J2_127_3477_n2616), 
        .A2(DP_OP_424J2_126_3477_n2227), .Y(DP_OP_423J2_125_3477_n2212) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2067 ( .A1(DP_OP_422J2_124_3477_n2000), 
        .A2(DP_OP_423J2_125_3477_n2843), .Y(DP_OP_424J2_126_3477_n2828) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2225 ( .A1(DP_OP_423J2_125_3477_n3008), 
        .A2(DP_OP_422J2_124_3477_n3015), .Y(DP_OP_423J2_125_3477_n2984) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1437 ( .A1(DP_OP_423J2_125_3477_n2134), 
        .A2(DP_OP_424J2_126_3477_n2225), .Y(DP_OP_424J2_126_3477_n2198) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1796 ( .A1(DP_OP_425J2_127_3477_n2397), 
        .A2(DP_OP_424J2_126_3477_n2578), .Y(DP_OP_424J2_126_3477_n2557) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1451 ( .A1(DP_OP_424J2_126_3477_n2220), 
        .A2(DP_OP_424J2_126_3477_n2227), .Y(DP_OP_424J2_126_3477_n2212) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1481 ( .A1(DP_OP_425J2_127_3477_n2662), 
        .A2(DP_OP_424J2_126_3477_n2269), .Y(DP_OP_424J2_126_3477_n2242) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2181 ( .A1(DP_OP_425J2_127_3477_n2086), 
        .A2(DP_OP_423J2_125_3477_n2973), .Y(DP_OP_423J2_125_3477_n2942) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1829 ( .A1(DP_OP_425J2_127_3477_n2438), 
        .A2(DP_OP_423J2_125_3477_n2621), .Y(DP_OP_423J2_125_3477_n2590) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1792 ( .A1(DP_OP_423J2_125_3477_n2569), 
        .A2(DP_OP_424J2_126_3477_n2578), .Y(DP_OP_423J2_125_3477_n2553) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1832 ( .A1(DP_OP_423J2_125_3477_n2617), 
        .A2(DP_OP_423J2_125_3477_n2621), .Y(DP_OP_423J2_125_3477_n2593) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1481 ( .A1(DP_OP_423J2_125_3477_n2266), 
        .A2(DP_OP_422J2_124_3477_n2269), .Y(DP_OP_423J2_125_3477_n2242) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1754 ( .A1(DP_OP_423J2_125_3477_n2619), 
        .A2(DP_OP_423J2_125_3477_n2534), .Y(DP_OP_424J2_126_3477_n2515) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1168 ( .A1(DP_OP_424J2_126_3477_n3007), 
        .A2(DP_OP_425J2_127_3477_n1961), .Y(DP_OP_425J2_127_3477_n1929) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1520 ( .A1(DP_OP_425J2_127_3477_n2305), 
        .A2(DP_OP_425J2_127_3477_n2313), .Y(DP_OP_425J2_127_3477_n2281) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1223 ( .A1(DP_OP_423J2_125_3477_n2000), 
        .A2(DP_OP_423J2_125_3477_n2006), .Y(DP_OP_423J2_125_3477_n1984) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2235 ( .A1(DP_OP_423J2_125_3477_n3010), 
        .A2(DP_OP_423J2_125_3477_n3016), .Y(DP_OP_423J2_125_3477_n2994) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1393 ( .A1(DP_OP_423J2_125_3477_n2178), 
        .A2(DP_OP_423J2_125_3477_n2181), .Y(DP_OP_423J2_125_3477_n2154) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1626 ( .A1(DP_OP_422J2_124_3477_n2571), 
        .A2(DP_OP_423J2_125_3477_n2403), .Y(DP_OP_423J2_125_3477_n2387) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1216 ( .A1(DP_OP_422J2_124_3477_n2969), 
        .A2(DP_OP_423J2_125_3477_n2005), .Y(DP_OP_423J2_125_3477_n1977) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1179 ( .A1(DP_OP_424J2_126_3477_n2044), 
        .A2(DP_OP_423J2_125_3477_n1962), .Y(DP_OP_423J2_125_3477_n1940) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1744 ( .A1(DP_OP_423J2_125_3477_n2529), 
        .A2(DP_OP_423J2_125_3477_n2533), .Y(DP_OP_423J2_125_3477_n2505) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1935 ( .A1(DP_OP_422J2_124_3477_n2220), 
        .A2(DP_OP_422J2_124_3477_n2711), .Y(DP_OP_423J2_125_3477_n2696) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1883 ( .A1(DP_OP_424J2_126_3477_n2572), 
        .A2(DP_OP_425J2_127_3477_n2666), .Y(DP_OP_423J2_125_3477_n2644) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1846 ( .A1(DP_OP_425J2_127_3477_n2439), 
        .A2(DP_OP_423J2_125_3477_n2623), .Y(DP_OP_423J2_125_3477_n2607) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2185 ( .A1(DP_OP_423J2_125_3477_n2970), 
        .A2(DP_OP_423J2_125_3477_n2973), .Y(DP_OP_423J2_125_3477_n2946) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2114 ( .A1(DP_OP_424J2_126_3477_n2883), 
        .A2(DP_OP_424J2_126_3477_n2887), .Y(DP_OP_424J2_126_3477_n2875) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2158 ( .A1(DP_OP_424J2_126_3477_n2927), 
        .A2(DP_OP_425J2_127_3477_n2931), .Y(DP_OP_424J2_126_3477_n2919) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1410 ( .A1(DP_OP_424J2_126_3477_n2179), 
        .A2(DP_OP_424J2_126_3477_n2183), .Y(DP_OP_424J2_126_3477_n2171) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1454 ( .A1(DP_OP_423J2_125_3477_n2135), 
        .A2(DP_OP_424J2_126_3477_n2227), .Y(DP_OP_424J2_126_3477_n2215) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1762 ( .A1(DP_OP_423J2_125_3477_n2619), 
        .A2(DP_OP_425J2_127_3477_n2535), .Y(DP_OP_424J2_126_3477_n2523) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1850 ( .A1(DP_OP_425J2_127_3477_n2355), 
        .A2(DP_OP_424J2_126_3477_n2623), .Y(DP_OP_424J2_126_3477_n2611) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2246 ( .A1(DP_OP_424J2_126_3477_n3013), 
        .A2(DP_OP_423J2_125_3477_n3017), .Y(DP_OP_424J2_126_3477_n3005) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2026 ( .A1(DP_OP_424J2_126_3477_n2795), 
        .A2(DP_OP_424J2_126_3477_n2799), .Y(DP_OP_424J2_126_3477_n2787) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2070 ( .A1(DP_OP_423J2_125_3477_n2927), 
        .A2(DP_OP_425J2_127_3477_n2843), .Y(DP_OP_424J2_126_3477_n2831) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1542 ( .A1(DP_OP_422J2_124_3477_n2751), 
        .A2(DP_OP_424J2_126_3477_n2315), .Y(DP_OP_424J2_126_3477_n2303) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1498 ( .A1(DP_OP_425J2_127_3477_n2663), 
        .A2(DP_OP_424J2_126_3477_n2271), .Y(DP_OP_424J2_126_3477_n2259) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1586 ( .A1(DP_OP_422J2_124_3477_n2707), 
        .A2(DP_OP_423J2_125_3477_n2359), .Y(DP_OP_424J2_126_3477_n2347) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1674 ( .A1(DP_OP_422J2_124_3477_n2619), 
        .A2(DP_OP_424J2_126_3477_n2447), .Y(DP_OP_424J2_126_3477_n2435) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1630 ( .A1(DP_OP_423J2_125_3477_n2311), 
        .A2(DP_OP_423J2_125_3477_n2403), .Y(DP_OP_424J2_126_3477_n2391) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1718 ( .A1(DP_OP_422J2_124_3477_n2355), 
        .A2(DP_OP_423J2_125_3477_n2491), .Y(DP_OP_424J2_126_3477_n2479) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1938 ( .A1(DP_OP_422J2_124_3477_n2135), 
        .A2(DP_OP_424J2_126_3477_n2711), .Y(DP_OP_424J2_126_3477_n2699) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1894 ( .A1(DP_OP_424J2_126_3477_n2663), 
        .A2(DP_OP_422J2_124_3477_n2667), .Y(DP_OP_424J2_126_3477_n2655) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1539 ( .A1(DP_OP_423J2_125_3477_n2308), 
        .A2(DP_OP_423J2_125_3477_n2315), .Y(DP_OP_423J2_125_3477_n2300) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1752 ( .A1(DP_OP_423J2_125_3477_n2529), 
        .A2(DP_OP_423J2_125_3477_n2534), .Y(DP_OP_423J2_125_3477_n2513) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2062 ( .A1(DP_OP_423J2_125_3477_n2927), 
        .A2(DP_OP_422J2_124_3477_n2842), .Y(DP_OP_424J2_126_3477_n2823) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2025 ( .A1(DP_OP_424J2_126_3477_n2794), 
        .A2(DP_OP_424J2_126_3477_n2799), .Y(DP_OP_424J2_126_3477_n2786) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2106 ( .A1(DP_OP_424J2_126_3477_n2883), 
        .A2(DP_OP_424J2_126_3477_n2886), .Y(DP_OP_424J2_126_3477_n2867) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1886 ( .A1(DP_OP_424J2_126_3477_n2663), 
        .A2(DP_OP_424J2_126_3477_n2666), .Y(DP_OP_424J2_126_3477_n2647) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1893 ( .A1(DP_OP_422J2_124_3477_n2178), 
        .A2(DP_OP_423J2_125_3477_n2667), .Y(DP_OP_424J2_126_3477_n2654) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1578 ( .A1(DP_OP_422J2_124_3477_n2707), 
        .A2(DP_OP_424J2_126_3477_n2358), .Y(DP_OP_424J2_126_3477_n2339) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2236 ( .A1(DP_OP_423J2_125_3477_n3011), 
        .A2(DP_OP_423J2_125_3477_n3016), .Y(DP_OP_423J2_125_3477_n2995) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1622 ( .A1(DP_OP_423J2_125_3477_n2311), 
        .A2(DP_OP_424J2_126_3477_n2402), .Y(DP_OP_424J2_126_3477_n2383) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1585 ( .A1(DP_OP_424J2_126_3477_n2354), 
        .A2(DP_OP_422J2_124_3477_n2359), .Y(DP_OP_424J2_126_3477_n2346) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1629 ( .A1(DP_OP_425J2_127_3477_n2530), 
        .A2(DP_OP_422J2_124_3477_n2403), .Y(DP_OP_424J2_126_3477_n2390) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2229 ( .A1(DP_OP_423J2_125_3477_n3012), 
        .A2(DP_OP_422J2_124_3477_n3015), .Y(DP_OP_423J2_125_3477_n2988) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1226 ( .A1(DP_OP_425J2_127_3477_n2927), 
        .A2(DP_OP_422J2_124_3477_n2006), .Y(DP_OP_424J2_126_3477_n1987) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1182 ( .A1(DP_OP_425J2_127_3477_n2971), 
        .A2(DP_OP_424J2_126_3477_n1962), .Y(DP_OP_424J2_126_3477_n1943) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1233 ( .A1(DP_OP_425J2_127_3477_n2926), 
        .A2(DP_OP_422J2_124_3477_n2007), .Y(DP_OP_424J2_126_3477_n1994) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1930 ( .A1(DP_OP_422J2_124_3477_n2135), 
        .A2(DP_OP_423J2_125_3477_n2710), .Y(DP_OP_424J2_126_3477_n2691) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2113 ( .A1(DP_OP_423J2_125_3477_n2970), 
        .A2(DP_OP_424J2_126_3477_n2887), .Y(DP_OP_424J2_126_3477_n2874) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1849 ( .A1(DP_OP_424J2_126_3477_n2618), 
        .A2(DP_OP_424J2_126_3477_n2623), .Y(DP_OP_424J2_126_3477_n2610) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1673 ( .A1(DP_OP_424J2_126_3477_n2442), 
        .A2(DP_OP_424J2_126_3477_n2447), .Y(DP_OP_424J2_126_3477_n2434) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1666 ( .A1(DP_OP_422J2_124_3477_n2619), 
        .A2(DP_OP_424J2_126_3477_n2446), .Y(DP_OP_424J2_126_3477_n2427) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1710 ( .A1(DP_OP_422J2_124_3477_n2355), 
        .A2(DP_OP_425J2_127_3477_n2490), .Y(DP_OP_424J2_126_3477_n2471) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1270 ( .A1(DP_OP_424J2_126_3477_n2047), 
        .A2(DP_OP_423J2_125_3477_n2050), .Y(DP_OP_424J2_126_3477_n2031) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1937 ( .A1(DP_OP_422J2_124_3477_n2134), 
        .A2(DP_OP_424J2_126_3477_n2711), .Y(DP_OP_424J2_126_3477_n2698) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2157 ( .A1(DP_OP_424J2_126_3477_n2926), 
        .A2(DP_OP_422J2_124_3477_n2931), .Y(DP_OP_424J2_126_3477_n2918) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2150 ( .A1(DP_OP_424J2_126_3477_n2927), 
        .A2(DP_OP_423J2_125_3477_n2930), .Y(DP_OP_424J2_126_3477_n2911) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2245 ( .A1(DP_OP_424J2_126_3477_n3012), 
        .A2(DP_OP_425J2_127_3477_n3017), .Y(DP_OP_424J2_126_3477_n3004) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1798 ( .A1(DP_OP_423J2_125_3477_n2663), 
        .A2(DP_OP_424J2_126_3477_n2578), .Y(DP_OP_424J2_126_3477_n2559) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2238 ( .A1(DP_OP_424J2_126_3477_n3013), 
        .A2(DP_OP_424J2_126_3477_n3016), .Y(DP_OP_424J2_126_3477_n2997) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1358 ( .A1(DP_OP_422J2_124_3477_n2927), 
        .A2(DP_OP_425J2_127_3477_n2138), .Y(DP_OP_424J2_126_3477_n2119) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2018 ( .A1(DP_OP_424J2_126_3477_n2795), 
        .A2(DP_OP_422J2_124_3477_n2798), .Y(DP_OP_424J2_126_3477_n2779) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2201 ( .A1(DP_OP_424J2_126_3477_n2970), 
        .A2(DP_OP_424J2_126_3477_n2975), .Y(DP_OP_424J2_126_3477_n2962) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2194 ( .A1(DP_OP_425J2_127_3477_n2003), 
        .A2(DP_OP_422J2_124_3477_n2974), .Y(DP_OP_424J2_126_3477_n2955) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1409 ( .A1(DP_OP_424J2_126_3477_n2178), 
        .A2(DP_OP_424J2_126_3477_n2183), .Y(DP_OP_424J2_126_3477_n2170) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1402 ( .A1(DP_OP_424J2_126_3477_n2179), 
        .A2(DP_OP_424J2_126_3477_n2182), .Y(DP_OP_424J2_126_3477_n2163) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1490 ( .A1(DP_OP_425J2_127_3477_n2663), 
        .A2(DP_OP_424J2_126_3477_n2270), .Y(DP_OP_424J2_126_3477_n2251) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1453 ( .A1(DP_OP_422J2_124_3477_n2838), 
        .A2(DP_OP_424J2_126_3477_n2227), .Y(DP_OP_424J2_126_3477_n2214) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1497 ( .A1(DP_OP_423J2_125_3477_n2178), 
        .A2(DP_OP_424J2_126_3477_n2271), .Y(DP_OP_424J2_126_3477_n2258) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1541 ( .A1(DP_OP_424J2_126_3477_n2310), 
        .A2(DP_OP_424J2_126_3477_n2315), .Y(DP_OP_424J2_126_3477_n2302) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1708 ( .A1(DP_OP_422J2_124_3477_n2441), 
        .A2(DP_OP_423J2_125_3477_n2490), .Y(DP_OP_423J2_125_3477_n2469) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1400 ( .A1(DP_OP_422J2_124_3477_n2793), 
        .A2(DP_OP_422J2_124_3477_n2182), .Y(DP_OP_423J2_125_3477_n2161) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1407 ( .A1(DP_OP_424J2_126_3477_n2264), 
        .A2(DP_OP_423J2_125_3477_n2183), .Y(DP_OP_423J2_125_3477_n2168) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2060 ( .A1(DP_OP_423J2_125_3477_n2837), 
        .A2(DP_OP_423J2_125_3477_n2842), .Y(DP_OP_423J2_125_3477_n2821) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2053 ( .A1(DP_OP_424J2_126_3477_n2750), 
        .A2(DP_OP_422J2_124_3477_n2841), .Y(DP_OP_423J2_125_3477_n2814) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2202 ( .A1(DP_OP_425J2_127_3477_n2003), 
        .A2(DP_OP_424J2_126_3477_n2975), .Y(DP_OP_424J2_126_3477_n2963) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1487 ( .A1(DP_OP_424J2_126_3477_n2264), 
        .A2(DP_OP_424J2_126_3477_n2270), .Y(DP_OP_424J2_126_3477_n2248) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1391 ( .A1(DP_OP_424J2_126_3477_n2264), 
        .A2(DP_OP_423J2_125_3477_n2181), .Y(DP_OP_423J2_125_3477_n2152) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2014 ( .A1(DP_OP_423J2_125_3477_n2791), 
        .A2(DP_OP_423J2_125_3477_n2798), .Y(DP_OP_423J2_125_3477_n2775) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1171 ( .A1(DP_OP_424J2_126_3477_n2044), 
        .A2(DP_OP_422J2_124_3477_n1961), .Y(DP_OP_423J2_125_3477_n1932) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2241 ( .A1(DP_OP_423J2_125_3477_n3008), 
        .A2(DP_OP_423J2_125_3477_n3017), .Y(DP_OP_423J2_125_3477_n3000) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1618 ( .A1(DP_OP_422J2_124_3477_n2571), 
        .A2(DP_OP_423J2_125_3477_n2402), .Y(DP_OP_423J2_125_3477_n2379) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1565 ( .A1(DP_OP_423J2_125_3477_n2350), 
        .A2(DP_OP_423J2_125_3477_n2357), .Y(DP_OP_423J2_125_3477_n2326) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1794 ( .A1(DP_OP_423J2_125_3477_n2571), 
        .A2(DP_OP_424J2_126_3477_n2578), .Y(DP_OP_423J2_125_3477_n2555) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1259 ( .A1(DP_OP_423J2_125_3477_n2044), 
        .A2(DP_OP_425J2_127_3477_n2049), .Y(DP_OP_423J2_125_3477_n2020) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2065 ( .A1(DP_OP_423J2_125_3477_n2834), 
        .A2(DP_OP_423J2_125_3477_n2843), .Y(DP_OP_423J2_125_3477_n2826) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1572 ( .A1(DP_OP_422J2_124_3477_n2613), 
        .A2(DP_OP_423J2_125_3477_n2358), .Y(DP_OP_423J2_125_3477_n2333) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1567 ( .A1(DP_OP_422J2_124_3477_n2616), 
        .A2(DP_OP_423J2_125_3477_n2357), .Y(DP_OP_423J2_125_3477_n2328) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1354 ( .A1(DP_OP_422J2_124_3477_n2835), 
        .A2(DP_OP_423J2_125_3477_n2138), .Y(DP_OP_423J2_125_3477_n2115) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1347 ( .A1(DP_OP_425J2_127_3477_n2704), 
        .A2(DP_OP_422J2_124_3477_n2137), .Y(DP_OP_423J2_125_3477_n2108) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2021 ( .A1(DP_OP_423J2_125_3477_n2790), 
        .A2(DP_OP_424J2_126_3477_n2799), .Y(DP_OP_423J2_125_3477_n2782) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1476 ( .A1(DP_OP_424J2_126_3477_n2261), 
        .A2(DP_OP_424J2_126_3477_n2269), .Y(DP_OP_424J2_126_3477_n2237) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1266 ( .A1(DP_OP_425J2_127_3477_n2791), 
        .A2(DP_OP_423J2_125_3477_n2050), .Y(DP_OP_423J2_125_3477_n2027) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1960 ( .A1(DP_OP_424J2_126_3477_n2745), 
        .A2(DP_OP_424J2_126_3477_n2753), .Y(DP_OP_424J2_126_3477_n2721) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1872 ( .A1(DP_OP_425J2_127_3477_n2305), 
        .A2(DP_OP_424J2_126_3477_n2665), .Y(DP_OP_424J2_126_3477_n2633) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1405 ( .A1(DP_OP_425J2_127_3477_n2658), 
        .A2(DP_OP_423J2_125_3477_n2183), .Y(DP_OP_423J2_125_3477_n2166) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1875 ( .A1(DP_OP_423J2_125_3477_n2748), 
        .A2(DP_OP_424J2_126_3477_n2665), .Y(DP_OP_424J2_126_3477_n2636) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1625 ( .A1(DP_OP_425J2_127_3477_n2526), 
        .A2(DP_OP_423J2_125_3477_n2403), .Y(DP_OP_424J2_126_3477_n2386) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1215 ( .A1(DP_OP_425J2_127_3477_n2924), 
        .A2(DP_OP_423J2_125_3477_n2005), .Y(DP_OP_424J2_126_3477_n1976) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2234 ( .A1(DP_OP_424J2_126_3477_n3009), 
        .A2(DP_OP_424J2_126_3477_n3016), .Y(DP_OP_424J2_126_3477_n2993) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1398 ( .A1(DP_OP_423J2_125_3477_n2175), 
        .A2(DP_OP_424J2_126_3477_n2182), .Y(DP_OP_423J2_125_3477_n2159) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1301 ( .A1(DP_OP_423J2_125_3477_n2086), 
        .A2(DP_OP_423J2_125_3477_n2093), .Y(DP_OP_423J2_125_3477_n2062) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1435 ( .A1(DP_OP_424J2_126_3477_n2220), 
        .A2(DP_OP_424J2_126_3477_n2225), .Y(DP_OP_424J2_126_3477_n2196) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1523 ( .A1(DP_OP_424J2_126_3477_n2308), 
        .A2(DP_OP_423J2_125_3477_n2313), .Y(DP_OP_424J2_126_3477_n2284) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2109 ( .A1(DP_OP_424J2_126_3477_n2878), 
        .A2(DP_OP_424J2_126_3477_n2887), .Y(DP_OP_424J2_126_3477_n2870) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2102 ( .A1(DP_OP_425J2_127_3477_n2087), 
        .A2(DP_OP_424J2_126_3477_n2886), .Y(DP_OP_424J2_126_3477_n2863) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1493 ( .A1(DP_OP_425J2_127_3477_n2658), 
        .A2(DP_OP_424J2_126_3477_n2271), .Y(DP_OP_424J2_126_3477_n2254) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1229 ( .A1(DP_OP_425J2_127_3477_n2922), 
        .A2(DP_OP_423J2_125_3477_n2007), .Y(DP_OP_424J2_126_3477_n1990) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1926 ( .A1(DP_OP_424J2_126_3477_n2703), 
        .A2(DP_OP_422J2_124_3477_n2710), .Y(DP_OP_424J2_126_3477_n2687) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1713 ( .A1(DP_OP_424J2_126_3477_n2482), 
        .A2(DP_OP_425J2_127_3477_n2491), .Y(DP_OP_424J2_126_3477_n2474) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1743 ( .A1(DP_OP_424J2_126_3477_n2528), 
        .A2(DP_OP_424J2_126_3477_n2533), .Y(DP_OP_424J2_126_3477_n2504) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1537 ( .A1(DP_OP_422J2_124_3477_n2746), 
        .A2(DP_OP_424J2_126_3477_n2315), .Y(DP_OP_424J2_126_3477_n2298) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2153 ( .A1(DP_OP_424J2_126_3477_n2922), 
        .A2(DP_OP_422J2_124_3477_n2931), .Y(DP_OP_424J2_126_3477_n2914) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2146 ( .A1(DP_OP_424J2_126_3477_n2923), 
        .A2(DP_OP_423J2_125_3477_n2930), .Y(DP_OP_424J2_126_3477_n2907) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1222 ( .A1(DP_OP_425J2_127_3477_n2923), 
        .A2(DP_OP_425J2_127_3477_n2006), .Y(DP_OP_424J2_126_3477_n1983) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2139 ( .A1(DP_OP_424J2_126_3477_n2924), 
        .A2(DP_OP_424J2_126_3477_n2929), .Y(DP_OP_424J2_126_3477_n2900) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1449 ( .A1(DP_OP_424J2_126_3477_n2218), 
        .A2(DP_OP_424J2_126_3477_n2227), .Y(DP_OP_424J2_126_3477_n2210) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1479 ( .A1(DP_OP_424J2_126_3477_n2264), 
        .A2(DP_OP_424J2_126_3477_n2269), .Y(DP_OP_424J2_126_3477_n2240) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1581 ( .A1(DP_OP_422J2_124_3477_n2702), 
        .A2(DP_OP_425J2_127_3477_n2359), .Y(DP_OP_424J2_126_3477_n2342) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2227 ( .A1(DP_OP_424J2_126_3477_n3010), 
        .A2(DP_OP_424J2_126_3477_n3015), .Y(DP_OP_424J2_126_3477_n2986) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2197 ( .A1(DP_OP_425J2_127_3477_n1998), 
        .A2(DP_OP_424J2_126_3477_n2975), .Y(DP_OP_424J2_126_3477_n2958) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1574 ( .A1(DP_OP_424J2_126_3477_n2351), 
        .A2(DP_OP_424J2_126_3477_n2358), .Y(DP_OP_424J2_126_3477_n2335) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2190 ( .A1(DP_OP_424J2_126_3477_n2967), 
        .A2(DP_OP_425J2_127_3477_n2974), .Y(DP_OP_424J2_126_3477_n2951) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2183 ( .A1(DP_OP_425J2_127_3477_n2000), 
        .A2(DP_OP_422J2_124_3477_n2973), .Y(DP_OP_424J2_126_3477_n2944) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1757 ( .A1(DP_OP_423J2_125_3477_n2526), 
        .A2(DP_OP_423J2_125_3477_n2535), .Y(DP_OP_423J2_125_3477_n2518) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1750 ( .A1(DP_OP_423J2_125_3477_n2527), 
        .A2(DP_OP_423J2_125_3477_n2534), .Y(DP_OP_423J2_125_3477_n2511) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1406 ( .A1(DP_OP_423J2_125_3477_n2175), 
        .A2(DP_OP_423J2_125_3477_n2183), .Y(DP_OP_423J2_125_3477_n2167) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1919 ( .A1(DP_OP_424J2_126_3477_n2616), 
        .A2(DP_OP_423J2_125_3477_n2709), .Y(DP_OP_423J2_125_3477_n2680) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1669 ( .A1(DP_OP_422J2_124_3477_n2526), 
        .A2(DP_OP_422J2_124_3477_n2447), .Y(DP_OP_423J2_125_3477_n2430) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1662 ( .A1(DP_OP_423J2_125_3477_n2439), 
        .A2(DP_OP_423J2_125_3477_n2446), .Y(DP_OP_423J2_125_3477_n2423) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1963 ( .A1(DP_OP_423J2_125_3477_n2748), 
        .A2(DP_OP_423J2_125_3477_n2753), .Y(DP_OP_423J2_125_3477_n2724) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2050 ( .A1(DP_OP_424J2_126_3477_n2835), 
        .A2(DP_OP_422J2_124_3477_n2841), .Y(DP_OP_424J2_126_3477_n2811) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1302 ( .A1(DP_OP_424J2_126_3477_n2087), 
        .A2(DP_OP_425J2_127_3477_n2093), .Y(DP_OP_424J2_126_3477_n2063) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1178 ( .A1(DP_OP_422J2_124_3477_n3009), 
        .A2(DP_OP_423J2_125_3477_n1962), .Y(DP_OP_423J2_125_3477_n1939) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2015 ( .A1(DP_OP_425J2_127_3477_n2264), 
        .A2(DP_OP_423J2_125_3477_n2798), .Y(DP_OP_423J2_125_3477_n2776) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1611 ( .A1(DP_OP_423J2_125_3477_n2396), 
        .A2(DP_OP_423J2_125_3477_n2401), .Y(DP_OP_423J2_125_3477_n2372) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1845 ( .A1(DP_OP_424J2_126_3477_n2526), 
        .A2(DP_OP_423J2_125_3477_n2623), .Y(DP_OP_423J2_125_3477_n2606) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1831 ( .A1(DP_OP_424J2_126_3477_n2528), 
        .A2(DP_OP_423J2_125_3477_n2621), .Y(DP_OP_423J2_125_3477_n2592) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2154 ( .A1(DP_OP_423J2_125_3477_n2923), 
        .A2(DP_OP_423J2_125_3477_n2931), .Y(DP_OP_423J2_125_3477_n2915) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1582 ( .A1(DP_OP_423J2_125_3477_n2351), 
        .A2(DP_OP_423J2_125_3477_n2359), .Y(DP_OP_423J2_125_3477_n2343) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2184 ( .A1(DP_OP_423J2_125_3477_n2969), 
        .A2(DP_OP_423J2_125_3477_n2973), .Y(DP_OP_423J2_125_3477_n2945) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2191 ( .A1(DP_OP_424J2_126_3477_n2880), 
        .A2(DP_OP_423J2_125_3477_n2974), .Y(DP_OP_423J2_125_3477_n2952) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1656 ( .A1(DP_OP_423J2_125_3477_n2441), 
        .A2(DP_OP_423J2_125_3477_n2445), .Y(DP_OP_423J2_125_3477_n2417) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1927 ( .A1(DP_OP_422J2_124_3477_n2220), 
        .A2(DP_OP_423J2_125_3477_n2710), .Y(DP_OP_423J2_125_3477_n2688) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1612 ( .A1(DP_OP_423J2_125_3477_n2397), 
        .A2(DP_OP_423J2_125_3477_n2401), .Y(DP_OP_423J2_125_3477_n2373) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1348 ( .A1(DP_OP_422J2_124_3477_n2837), 
        .A2(DP_OP_422J2_124_3477_n2137), .Y(DP_OP_423J2_125_3477_n2109) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2066 ( .A1(DP_OP_424J2_126_3477_n2747), 
        .A2(DP_OP_423J2_125_3477_n2843), .Y(DP_OP_423J2_125_3477_n2827) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1707 ( .A1(DP_OP_423J2_125_3477_n2484), 
        .A2(DP_OP_423J2_125_3477_n2490), .Y(DP_OP_423J2_125_3477_n2468) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1663 ( .A1(DP_OP_422J2_124_3477_n2528), 
        .A2(DP_OP_423J2_125_3477_n2446), .Y(DP_OP_423J2_125_3477_n2424) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2059 ( .A1(DP_OP_422J2_124_3477_n2088), 
        .A2(DP_OP_423J2_125_3477_n2842), .Y(DP_OP_423J2_125_3477_n2820) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2052 ( .A1(DP_OP_423J2_125_3477_n2837), 
        .A2(DP_OP_422J2_124_3477_n2841), .Y(DP_OP_423J2_125_3477_n2813) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1256 ( .A1(DP_OP_422J2_124_3477_n3007), 
        .A2(DP_OP_424J2_126_3477_n2049), .Y(DP_OP_424J2_126_3477_n2017) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1486 ( .A1(DP_OP_423J2_125_3477_n2263), 
        .A2(DP_OP_423J2_125_3477_n2270), .Y(DP_OP_423J2_125_3477_n2247) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1706 ( .A1(DP_OP_422J2_124_3477_n2439), 
        .A2(DP_OP_423J2_125_3477_n2490), .Y(DP_OP_423J2_125_3477_n2467) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1564 ( .A1(DP_OP_422J2_124_3477_n2701), 
        .A2(DP_OP_424J2_126_3477_n2357), .Y(DP_OP_424J2_126_3477_n2325) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1699 ( .A1(DP_OP_423J2_125_3477_n2484), 
        .A2(DP_OP_423J2_125_3477_n2489), .Y(DP_OP_423J2_125_3477_n2460) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1696 ( .A1(DP_OP_424J2_126_3477_n2481), 
        .A2(DP_OP_424J2_126_3477_n2489), .Y(DP_OP_424J2_126_3477_n2457) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1933 ( .A1(DP_OP_423J2_125_3477_n2702), 
        .A2(DP_OP_424J2_126_3477_n2711), .Y(DP_OP_423J2_125_3477_n2694) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2137 ( .A1(DP_OP_423J2_125_3477_n2922), 
        .A2(DP_OP_423J2_125_3477_n2929), .Y(DP_OP_423J2_125_3477_n2898) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2051 ( .A1(DP_OP_422J2_124_3477_n2088), 
        .A2(DP_OP_423J2_125_3477_n2841), .Y(DP_OP_423J2_125_3477_n2812) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1303 ( .A1(DP_OP_423J2_125_3477_n2088), 
        .A2(DP_OP_423J2_125_3477_n2093), .Y(DP_OP_423J2_125_3477_n2064) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2058 ( .A1(DP_OP_425J2_127_3477_n2219), 
        .A2(DP_OP_423J2_125_3477_n2842), .Y(DP_OP_423J2_125_3477_n2819) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1655 ( .A1(DP_OP_422J2_124_3477_n2528), 
        .A2(DP_OP_423J2_125_3477_n2445), .Y(DP_OP_423J2_125_3477_n2416) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1213 ( .A1(DP_OP_423J2_125_3477_n1998), 
        .A2(DP_OP_423J2_125_3477_n2005), .Y(DP_OP_423J2_125_3477_n1974) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2147 ( .A1(DP_OP_423J2_125_3477_n2924), 
        .A2(DP_OP_423J2_125_3477_n2930), .Y(DP_OP_423J2_125_3477_n2908) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1568 ( .A1(DP_OP_424J2_126_3477_n2353), 
        .A2(DP_OP_424J2_126_3477_n2357), .Y(DP_OP_424J2_126_3477_n2329) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2013 ( .A1(DP_OP_424J2_126_3477_n2790), 
        .A2(DP_OP_422J2_124_3477_n2798), .Y(DP_OP_424J2_126_3477_n2774) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2233 ( .A1(DP_OP_424J2_126_3477_n3008), 
        .A2(DP_OP_424J2_126_3477_n3016), .Y(DP_OP_424J2_126_3477_n2992) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2226 ( .A1(DP_OP_424J2_126_3477_n3009), 
        .A2(DP_OP_424J2_126_3477_n3015), .Y(DP_OP_424J2_126_3477_n2985) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1573 ( .A1(DP_OP_422J2_124_3477_n2702), 
        .A2(DP_OP_424J2_126_3477_n2358), .Y(DP_OP_424J2_126_3477_n2334) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2196 ( .A1(DP_OP_425J2_127_3477_n1997), 
        .A2(DP_OP_424J2_126_3477_n2975), .Y(DP_OP_424J2_126_3477_n2957) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2189 ( .A1(DP_OP_425J2_127_3477_n1998), 
        .A2(DP_OP_425J2_127_3477_n2974), .Y(DP_OP_424J2_126_3477_n2950) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1660 ( .A1(DP_OP_423J2_125_3477_n2437), 
        .A2(DP_OP_423J2_125_3477_n2446), .Y(DP_OP_423J2_125_3477_n2421) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1654 ( .A1(DP_OP_424J2_126_3477_n2439), 
        .A2(DP_OP_424J2_126_3477_n2445), .Y(DP_OP_424J2_126_3477_n2415) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1661 ( .A1(DP_OP_423J2_125_3477_n2350), 
        .A2(DP_OP_424J2_126_3477_n2446), .Y(DP_OP_424J2_126_3477_n2422) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1258 ( .A1(DP_OP_425J2_127_3477_n2879), 
        .A2(DP_OP_424J2_126_3477_n2049), .Y(DP_OP_424J2_126_3477_n2019) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1265 ( .A1(DP_OP_422J2_124_3477_n3008), 
        .A2(DP_OP_423J2_125_3477_n2050), .Y(DP_OP_424J2_126_3477_n2026) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1390 ( .A1(DP_OP_425J2_127_3477_n2747), 
        .A2(DP_OP_423J2_125_3477_n2181), .Y(DP_OP_424J2_126_3477_n2151) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1397 ( .A1(DP_OP_423J2_125_3477_n2086), 
        .A2(DP_OP_424J2_126_3477_n2182), .Y(DP_OP_424J2_126_3477_n2158) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1302 ( .A1(DP_OP_423J2_125_3477_n2087), 
        .A2(DP_OP_423J2_125_3477_n2093), .Y(DP_OP_423J2_125_3477_n2063) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1917 ( .A1(DP_OP_423J2_125_3477_n2702), 
        .A2(DP_OP_423J2_125_3477_n2709), .Y(DP_OP_423J2_125_3477_n2678) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2182 ( .A1(DP_OP_424J2_126_3477_n2967), 
        .A2(DP_OP_425J2_127_3477_n2973), .Y(DP_OP_424J2_126_3477_n2943) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2152 ( .A1(DP_OP_424J2_126_3477_n2921), 
        .A2(DP_OP_423J2_125_3477_n2931), .Y(DP_OP_424J2_126_3477_n2913) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2050 ( .A1(DP_OP_424J2_126_3477_n2747), 
        .A2(DP_OP_423J2_125_3477_n2841), .Y(DP_OP_423J2_125_3477_n2811) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1177 ( .A1(DP_OP_424J2_126_3477_n1954), 
        .A2(DP_OP_424J2_126_3477_n1962), .Y(DP_OP_424J2_126_3477_n1938) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2145 ( .A1(DP_OP_424J2_126_3477_n2922), 
        .A2(DP_OP_422J2_124_3477_n2930), .Y(DP_OP_424J2_126_3477_n2906) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1609 ( .A1(DP_OP_422J2_124_3477_n2570), 
        .A2(DP_OP_423J2_125_3477_n2401), .Y(DP_OP_423J2_125_3477_n2370) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1616 ( .A1(DP_OP_422J2_124_3477_n2569), 
        .A2(DP_OP_423J2_125_3477_n2402), .Y(DP_OP_423J2_125_3477_n2377) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1575 ( .A1(DP_OP_422J2_124_3477_n2616), 
        .A2(DP_OP_423J2_125_3477_n2358), .Y(DP_OP_423J2_125_3477_n2336) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2049 ( .A1(DP_OP_423J2_125_3477_n2834), 
        .A2(DP_OP_425J2_127_3477_n2841), .Y(DP_OP_423J2_125_3477_n2810) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1345 ( .A1(DP_OP_422J2_124_3477_n2834), 
        .A2(DP_OP_425J2_127_3477_n2137), .Y(DP_OP_423J2_125_3477_n2106) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1352 ( .A1(DP_OP_422J2_124_3477_n2833), 
        .A2(DP_OP_423J2_125_3477_n2138), .Y(DP_OP_423J2_125_3477_n2113) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2110 ( .A1(DP_OP_423J2_125_3477_n2967), 
        .A2(DP_OP_424J2_126_3477_n2887), .Y(DP_OP_424J2_126_3477_n2871) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2103 ( .A1(DP_OP_424J2_126_3477_n2880), 
        .A2(DP_OP_424J2_126_3477_n2886), .Y(DP_OP_424J2_126_3477_n2864) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1538 ( .A1(DP_OP_423J2_125_3477_n2219), 
        .A2(DP_OP_424J2_126_3477_n2315), .Y(DP_OP_424J2_126_3477_n2299) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1304 ( .A1(DP_OP_422J2_124_3477_n2969), 
        .A2(DP_OP_423J2_125_3477_n2093), .Y(DP_OP_424J2_126_3477_n2065) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1741 ( .A1(DP_OP_423J2_125_3477_n2526), 
        .A2(DP_OP_423J2_125_3477_n2533), .Y(DP_OP_423J2_125_3477_n2502) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1494 ( .A1(DP_OP_423J2_125_3477_n2175), 
        .A2(DP_OP_424J2_126_3477_n2271), .Y(DP_OP_424J2_126_3477_n2255) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1524 ( .A1(DP_OP_425J2_127_3477_n2617), 
        .A2(DP_OP_425J2_127_3477_n2313), .Y(DP_OP_424J2_126_3477_n2285) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2022 ( .A1(DP_OP_424J2_126_3477_n2791), 
        .A2(DP_OP_424J2_126_3477_n2799), .Y(DP_OP_424J2_126_3477_n2783) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1355 ( .A1(DP_OP_422J2_124_3477_n2924), 
        .A2(DP_OP_422J2_124_3477_n2138), .Y(DP_OP_424J2_126_3477_n2116) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1450 ( .A1(DP_OP_424J2_126_3477_n2219), 
        .A2(DP_OP_424J2_126_3477_n2227), .Y(DP_OP_424J2_126_3477_n2211) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1619 ( .A1(DP_OP_423J2_125_3477_n2308), 
        .A2(DP_OP_424J2_126_3477_n2402), .Y(DP_OP_424J2_126_3477_n2380) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2228 ( .A1(DP_OP_424J2_126_3477_n3011), 
        .A2(DP_OP_424J2_126_3477_n3015), .Y(DP_OP_424J2_126_3477_n2987) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1230 ( .A1(DP_OP_425J2_127_3477_n2923), 
        .A2(DP_OP_423J2_125_3477_n2007), .Y(DP_OP_424J2_126_3477_n1991) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2198 ( .A1(DP_OP_424J2_126_3477_n2967), 
        .A2(DP_OP_424J2_126_3477_n2975), .Y(DP_OP_424J2_126_3477_n2959) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1260 ( .A1(DP_OP_422J2_124_3477_n3011), 
        .A2(DP_OP_424J2_126_3477_n2049), .Y(DP_OP_424J2_126_3477_n2021) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2140 ( .A1(DP_OP_425J2_127_3477_n2133), 
        .A2(DP_OP_423J2_125_3477_n2929), .Y(DP_OP_423J2_125_3477_n2901) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1267 ( .A1(DP_OP_424J2_126_3477_n2044), 
        .A2(DP_OP_422J2_124_3477_n2050), .Y(DP_OP_424J2_126_3477_n2028) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1964 ( .A1(DP_OP_424J2_126_3477_n2749), 
        .A2(DP_OP_424J2_126_3477_n2753), .Y(DP_OP_424J2_126_3477_n2725) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1670 ( .A1(DP_OP_424J2_126_3477_n2439), 
        .A2(DP_OP_424J2_126_3477_n2447), .Y(DP_OP_424J2_126_3477_n2431) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1700 ( .A1(DP_OP_422J2_124_3477_n2353), 
        .A2(DP_OP_424J2_126_3477_n2489), .Y(DP_OP_424J2_126_3477_n2461) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1876 ( .A1(DP_OP_422J2_124_3477_n2177), 
        .A2(DP_OP_424J2_126_3477_n2665), .Y(DP_OP_424J2_126_3477_n2637) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1890 ( .A1(DP_OP_425J2_127_3477_n2307), 
        .A2(DP_OP_423J2_125_3477_n2667), .Y(DP_OP_424J2_126_3477_n2651) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1758 ( .A1(DP_OP_425J2_127_3477_n2439), 
        .A2(DP_OP_422J2_124_3477_n2535), .Y(DP_OP_424J2_126_3477_n2519) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1920 ( .A1(DP_OP_424J2_126_3477_n2705), 
        .A2(DP_OP_423J2_125_3477_n2709), .Y(DP_OP_424J2_126_3477_n2681) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1961 ( .A1(DP_OP_423J2_125_3477_n2746), 
        .A2(DP_OP_423J2_125_3477_n2753), .Y(DP_OP_423J2_125_3477_n2722) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1346 ( .A1(DP_OP_422J2_124_3477_n2923), 
        .A2(DP_OP_424J2_126_3477_n2137), .Y(DP_OP_424J2_126_3477_n2107) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1830 ( .A1(DP_OP_422J2_124_3477_n2219), 
        .A2(DP_OP_425J2_127_3477_n2621), .Y(DP_OP_424J2_126_3477_n2591) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1610 ( .A1(DP_OP_422J2_124_3477_n2659), 
        .A2(DP_OP_424J2_126_3477_n2401), .Y(DP_OP_424J2_126_3477_n2371) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1653 ( .A1(DP_OP_422J2_124_3477_n2526), 
        .A2(DP_OP_423J2_125_3477_n2445), .Y(DP_OP_423J2_125_3477_n2414) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2240 ( .A1(DP_OP_424J2_126_3477_n3007), 
        .A2(DP_OP_422J2_124_3477_n3017), .Y(DP_OP_424J2_126_3477_n2999) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1170 ( .A1(DP_OP_425J2_127_3477_n2967), 
        .A2(DP_OP_424J2_126_3477_n1961), .Y(DP_OP_424J2_126_3477_n1931) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1918 ( .A1(DP_OP_424J2_126_3477_n2703), 
        .A2(DP_OP_425J2_127_3477_n2709), .Y(DP_OP_424J2_126_3477_n2679) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1705 ( .A1(DP_OP_424J2_126_3477_n2482), 
        .A2(DP_OP_423J2_125_3477_n2490), .Y(DP_OP_424J2_126_3477_n2466) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1712 ( .A1(DP_OP_424J2_126_3477_n2481), 
        .A2(DP_OP_422J2_124_3477_n2491), .Y(DP_OP_424J2_126_3477_n2473) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1874 ( .A1(DP_OP_425J2_127_3477_n2307), 
        .A2(DP_OP_424J2_126_3477_n2665), .Y(DP_OP_424J2_126_3477_n2635) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1793 ( .A1(DP_OP_423J2_125_3477_n2658), 
        .A2(DP_OP_424J2_126_3477_n2578), .Y(DP_OP_424J2_126_3477_n2554) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1925 ( .A1(DP_OP_422J2_124_3477_n2130), 
        .A2(DP_OP_422J2_124_3477_n2710), .Y(DP_OP_424J2_126_3477_n2686) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1521 ( .A1(DP_OP_425J2_127_3477_n2526), 
        .A2(DP_OP_423J2_125_3477_n2313), .Y(DP_OP_423J2_125_3477_n2282) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1698 ( .A1(DP_OP_422J2_124_3477_n2351), 
        .A2(DP_OP_424J2_126_3477_n2489), .Y(DP_OP_424J2_126_3477_n2459) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1881 ( .A1(DP_OP_424J2_126_3477_n2658), 
        .A2(DP_OP_424J2_126_3477_n2666), .Y(DP_OP_424J2_126_3477_n2642) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1434 ( .A1(DP_OP_424J2_126_3477_n2219), 
        .A2(DP_OP_424J2_126_3477_n2225), .Y(DP_OP_424J2_126_3477_n2195) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1962 ( .A1(DP_OP_424J2_126_3477_n2747), 
        .A2(DP_OP_424J2_126_3477_n2753), .Y(DP_OP_424J2_126_3477_n2723) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1580 ( .A1(DP_OP_422J2_124_3477_n2701), 
        .A2(DP_OP_422J2_124_3477_n2359), .Y(DP_OP_424J2_126_3477_n2341) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1624 ( .A1(DP_OP_425J2_127_3477_n2525), 
        .A2(DP_OP_422J2_124_3477_n2403), .Y(DP_OP_424J2_126_3477_n2385) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1566 ( .A1(DP_OP_424J2_126_3477_n2351), 
        .A2(DP_OP_424J2_126_3477_n2357), .Y(DP_OP_424J2_126_3477_n2327) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1880 ( .A1(DP_OP_422J2_124_3477_n2261), 
        .A2(DP_OP_425J2_127_3477_n2666), .Y(DP_OP_423J2_125_3477_n2641) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2138 ( .A1(DP_OP_424J2_126_3477_n2923), 
        .A2(DP_OP_424J2_126_3477_n2929), .Y(DP_OP_424J2_126_3477_n2899) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1522 ( .A1(DP_OP_422J2_124_3477_n2747), 
        .A2(DP_OP_422J2_124_3477_n2313), .Y(DP_OP_424J2_126_3477_n2283) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1214 ( .A1(DP_OP_425J2_127_3477_n2923), 
        .A2(DP_OP_425J2_127_3477_n2005), .Y(DP_OP_424J2_126_3477_n1975) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2101 ( .A1(DP_OP_424J2_126_3477_n2878), 
        .A2(DP_OP_424J2_126_3477_n2886), .Y(DP_OP_424J2_126_3477_n2862) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1742 ( .A1(DP_OP_425J2_127_3477_n2439), 
        .A2(DP_OP_424J2_126_3477_n2533), .Y(DP_OP_424J2_126_3477_n2503) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1749 ( .A1(DP_OP_424J2_126_3477_n2526), 
        .A2(DP_OP_423J2_125_3477_n2534), .Y(DP_OP_424J2_126_3477_n2510) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1485 ( .A1(DP_OP_425J2_127_3477_n2658), 
        .A2(DP_OP_424J2_126_3477_n2270), .Y(DP_OP_424J2_126_3477_n2246) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1221 ( .A1(DP_OP_425J2_127_3477_n2922), 
        .A2(DP_OP_423J2_125_3477_n2006), .Y(DP_OP_424J2_126_3477_n1982) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2064 ( .A1(DP_OP_424J2_126_3477_n2833), 
        .A2(DP_OP_422J2_124_3477_n2843), .Y(DP_OP_424J2_126_3477_n2825) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1478 ( .A1(DP_OP_422J2_124_3477_n2791), 
        .A2(DP_OP_424J2_126_3477_n2269), .Y(DP_OP_424J2_126_3477_n2239) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2057 ( .A1(DP_OP_424J2_126_3477_n2834), 
        .A2(DP_OP_423J2_125_3477_n2842), .Y(DP_OP_424J2_126_3477_n2818) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1882 ( .A1(DP_OP_423J2_125_3477_n2747), 
        .A2(DP_OP_424J2_126_3477_n2666), .Y(DP_OP_424J2_126_3477_n2643) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1704 ( .A1(DP_OP_424J2_126_3477_n2481), 
        .A2(DP_OP_422J2_124_3477_n2490), .Y(DP_OP_424J2_126_3477_n2465) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2137 ( .A1(DP_OP_424J2_126_3477_n2922), 
        .A2(DP_OP_424J2_126_3477_n2929), .Y(DP_OP_424J2_126_3477_n2898) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1537 ( .A1(DP_OP_425J2_127_3477_n2526), 
        .A2(DP_OP_423J2_125_3477_n2315), .Y(DP_OP_423J2_125_3477_n2298) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2100 ( .A1(DP_OP_424J2_126_3477_n2877), 
        .A2(DP_OP_424J2_126_3477_n2886), .Y(DP_OP_424J2_126_3477_n2861) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1213 ( .A1(DP_OP_425J2_127_3477_n2922), 
        .A2(DP_OP_422J2_124_3477_n2005), .Y(DP_OP_424J2_126_3477_n1974) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1220 ( .A1(DP_OP_425J2_127_3477_n2921), 
        .A2(DP_OP_422J2_124_3477_n2006), .Y(DP_OP_424J2_126_3477_n1981) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1743 ( .A1(DP_OP_423J2_125_3477_n2528), 
        .A2(DP_OP_423J2_125_3477_n2533), .Y(DP_OP_423J2_125_3477_n2504) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1436 ( .A1(DP_OP_425J2_127_3477_n2617), 
        .A2(DP_OP_423J2_125_3477_n2225), .Y(DP_OP_423J2_125_3477_n2197) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1713 ( .A1(DP_OP_423J2_125_3477_n2482), 
        .A2(DP_OP_423J2_125_3477_n2491), .Y(DP_OP_423J2_125_3477_n2474) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1926 ( .A1(DP_OP_425J2_127_3477_n2351), 
        .A2(DP_OP_423J2_125_3477_n2710), .Y(DP_OP_423J2_125_3477_n2687) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1229 ( .A1(DP_OP_423J2_125_3477_n1998), 
        .A2(DP_OP_423J2_125_3477_n2007), .Y(DP_OP_423J2_125_3477_n1990) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1493 ( .A1(DP_OP_423J2_125_3477_n2262), 
        .A2(DP_OP_422J2_124_3477_n2271), .Y(DP_OP_423J2_125_3477_n2254) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2102 ( .A1(DP_OP_425J2_127_3477_n2175), 
        .A2(DP_OP_423J2_125_3477_n2886), .Y(DP_OP_423J2_125_3477_n2863) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1655 ( .A1(DP_OP_425J2_127_3477_n2484), 
        .A2(DP_OP_424J2_126_3477_n2445), .Y(DP_OP_424J2_126_3477_n2416) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2109 ( .A1(DP_OP_423J2_125_3477_n2878), 
        .A2(DP_OP_424J2_126_3477_n2887), .Y(DP_OP_423J2_125_3477_n2870) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2058 ( .A1(DP_OP_424J2_126_3477_n2835), 
        .A2(DP_OP_423J2_125_3477_n2842), .Y(DP_OP_424J2_126_3477_n2819) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1303 ( .A1(DP_OP_424J2_126_3477_n2088), 
        .A2(DP_OP_423J2_125_3477_n2093), .Y(DP_OP_424J2_126_3477_n2064) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2051 ( .A1(DP_OP_422J2_124_3477_n2000), 
        .A2(DP_OP_423J2_125_3477_n2841), .Y(DP_OP_424J2_126_3477_n2812) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1523 ( .A1(DP_OP_423J2_125_3477_n2308), 
        .A2(DP_OP_423J2_125_3477_n2313), .Y(DP_OP_423J2_125_3477_n2284) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1933 ( .A1(DP_OP_422J2_124_3477_n2130), 
        .A2(DP_OP_424J2_126_3477_n2711), .Y(DP_OP_424J2_126_3477_n2694) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1699 ( .A1(DP_OP_424J2_126_3477_n2484), 
        .A2(DP_OP_424J2_126_3477_n2489), .Y(DP_OP_424J2_126_3477_n2460) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1889 ( .A1(DP_OP_424J2_126_3477_n2658), 
        .A2(DP_OP_423J2_125_3477_n2667), .Y(DP_OP_424J2_126_3477_n2650) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1706 ( .A1(DP_OP_422J2_124_3477_n2351), 
        .A2(DP_OP_422J2_124_3477_n2490), .Y(DP_OP_424J2_126_3477_n2467) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1486 ( .A1(DP_OP_422J2_124_3477_n2791), 
        .A2(DP_OP_424J2_126_3477_n2270), .Y(DP_OP_424J2_126_3477_n2247) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1259 ( .A1(DP_OP_424J2_126_3477_n2044), 
        .A2(DP_OP_424J2_126_3477_n2049), .Y(DP_OP_424J2_126_3477_n2020) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1435 ( .A1(DP_OP_424J2_126_3477_n2308), 
        .A2(DP_OP_423J2_125_3477_n2225), .Y(DP_OP_423J2_125_3477_n2196) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1266 ( .A1(DP_OP_422J2_124_3477_n3009), 
        .A2(DP_OP_425J2_127_3477_n2050), .Y(DP_OP_424J2_126_3477_n2027) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1257 ( .A1(DP_OP_425J2_127_3477_n2790), 
        .A2(DP_OP_422J2_124_3477_n2049), .Y(DP_OP_423J2_125_3477_n2018) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2021 ( .A1(DP_OP_424J2_126_3477_n2790), 
        .A2(DP_OP_424J2_126_3477_n2799), .Y(DP_OP_424J2_126_3477_n2782) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1347 ( .A1(DP_OP_422J2_124_3477_n2924), 
        .A2(DP_OP_424J2_126_3477_n2137), .Y(DP_OP_424J2_126_3477_n2108) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1354 ( .A1(DP_OP_422J2_124_3477_n2923), 
        .A2(DP_OP_425J2_127_3477_n2138), .Y(DP_OP_424J2_126_3477_n2115) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1567 ( .A1(DP_OP_422J2_124_3477_n2704), 
        .A2(DP_OP_424J2_126_3477_n2357), .Y(DP_OP_424J2_126_3477_n2328) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2065 ( .A1(DP_OP_424J2_126_3477_n2834), 
        .A2(DP_OP_423J2_125_3477_n2843), .Y(DP_OP_424J2_126_3477_n2826) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1794 ( .A1(DP_OP_423J2_125_3477_n2659), 
        .A2(DP_OP_424J2_126_3477_n2578), .Y(DP_OP_424J2_126_3477_n2555) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1618 ( .A1(DP_OP_423J2_125_3477_n2307), 
        .A2(DP_OP_424J2_126_3477_n2402), .Y(DP_OP_424J2_126_3477_n2379) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2234 ( .A1(DP_OP_423J2_125_3477_n3009), 
        .A2(DP_OP_423J2_125_3477_n3016), .Y(DP_OP_423J2_125_3477_n2993) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1171 ( .A1(DP_OP_424J2_126_3477_n1956), 
        .A2(DP_OP_424J2_126_3477_n1961), .Y(DP_OP_424J2_126_3477_n1932) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2014 ( .A1(DP_OP_424J2_126_3477_n2791), 
        .A2(DP_OP_423J2_125_3477_n2798), .Y(DP_OP_424J2_126_3477_n2775) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1215 ( .A1(DP_OP_423J2_125_3477_n2000), 
        .A2(DP_OP_423J2_125_3477_n2005), .Y(DP_OP_423J2_125_3477_n1976) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1391 ( .A1(DP_OP_423J2_125_3477_n2088), 
        .A2(DP_OP_422J2_124_3477_n2181), .Y(DP_OP_424J2_126_3477_n2152) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1831 ( .A1(DP_OP_424J2_126_3477_n2616), 
        .A2(DP_OP_423J2_125_3477_n2621), .Y(DP_OP_424J2_126_3477_n2592) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1845 ( .A1(DP_OP_422J2_124_3477_n2218), 
        .A2(DP_OP_424J2_126_3477_n2623), .Y(DP_OP_424J2_126_3477_n2606) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1625 ( .A1(DP_OP_422J2_124_3477_n2570), 
        .A2(DP_OP_423J2_125_3477_n2403), .Y(DP_OP_423J2_125_3477_n2386) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1611 ( .A1(DP_OP_423J2_125_3477_n2308), 
        .A2(DP_OP_424J2_126_3477_n2401), .Y(DP_OP_424J2_126_3477_n2372) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1178 ( .A1(DP_OP_425J2_127_3477_n2967), 
        .A2(DP_OP_424J2_126_3477_n1962), .Y(DP_OP_424J2_126_3477_n1939) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1963 ( .A1(DP_OP_425J2_127_3477_n2220), 
        .A2(DP_OP_424J2_126_3477_n2753), .Y(DP_OP_424J2_126_3477_n2724) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1875 ( .A1(DP_OP_424J2_126_3477_n2572), 
        .A2(DP_OP_423J2_125_3477_n2665), .Y(DP_OP_423J2_125_3477_n2636) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1662 ( .A1(DP_OP_424J2_126_3477_n2439), 
        .A2(DP_OP_424J2_126_3477_n2446), .Y(DP_OP_424J2_126_3477_n2423) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1669 ( .A1(DP_OP_423J2_125_3477_n2350), 
        .A2(DP_OP_424J2_126_3477_n2447), .Y(DP_OP_424J2_126_3477_n2430) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1919 ( .A1(DP_OP_422J2_124_3477_n2132), 
        .A2(DP_OP_422J2_124_3477_n2709), .Y(DP_OP_424J2_126_3477_n2680) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1750 ( .A1(DP_OP_422J2_124_3477_n2307), 
        .A2(DP_OP_422J2_124_3477_n2534), .Y(DP_OP_424J2_126_3477_n2511) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1757 ( .A1(DP_OP_424J2_126_3477_n2526), 
        .A2(DP_OP_423J2_125_3477_n2535), .Y(DP_OP_424J2_126_3477_n2518) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1882 ( .A1(DP_OP_423J2_125_3477_n2659), 
        .A2(DP_OP_422J2_124_3477_n2666), .Y(DP_OP_423J2_125_3477_n2643) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1889 ( .A1(DP_OP_423J2_125_3477_n2658), 
        .A2(DP_OP_423J2_125_3477_n2667), .Y(DP_OP_423J2_125_3477_n2650) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1398 ( .A1(DP_OP_423J2_125_3477_n2087), 
        .A2(DP_OP_424J2_126_3477_n2182), .Y(DP_OP_424J2_126_3477_n2159) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1405 ( .A1(DP_OP_422J2_124_3477_n2878), 
        .A2(DP_OP_424J2_126_3477_n2183), .Y(DP_OP_424J2_126_3477_n2166) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1433 ( .A1(DP_OP_423J2_125_3477_n2218), 
        .A2(DP_OP_423J2_125_3477_n2225), .Y(DP_OP_423J2_125_3477_n2194) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2183 ( .A1(DP_OP_424J2_126_3477_n2880), 
        .A2(DP_OP_423J2_125_3477_n2973), .Y(DP_OP_423J2_125_3477_n2944) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2190 ( .A1(DP_OP_423J2_125_3477_n2967), 
        .A2(DP_OP_423J2_125_3477_n2974), .Y(DP_OP_423J2_125_3477_n2951) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2012 ( .A1(DP_OP_425J2_127_3477_n2261), 
        .A2(DP_OP_423J2_125_3477_n2798), .Y(DP_OP_423J2_125_3477_n2773) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1574 ( .A1(DP_OP_423J2_125_3477_n2351), 
        .A2(DP_OP_423J2_125_3477_n2358), .Y(DP_OP_423J2_125_3477_n2335) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2232 ( .A1(DP_OP_424J2_126_3477_n3007), 
        .A2(DP_OP_424J2_126_3477_n3016), .Y(DP_OP_424J2_126_3477_n2991) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1169 ( .A1(DP_OP_424J2_126_3477_n1954), 
        .A2(DP_OP_424J2_126_3477_n1961), .Y(DP_OP_424J2_126_3477_n1930) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2225 ( .A1(DP_OP_424J2_126_3477_n3008), 
        .A2(DP_OP_424J2_126_3477_n3015), .Y(DP_OP_424J2_126_3477_n2984) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2197 ( .A1(DP_OP_424J2_126_3477_n2878), 
        .A2(DP_OP_424J2_126_3477_n2975), .Y(DP_OP_423J2_125_3477_n2958) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2188 ( .A1(DP_OP_425J2_127_3477_n1997), 
        .A2(DP_OP_422J2_124_3477_n2974), .Y(DP_OP_424J2_126_3477_n2949) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2181 ( .A1(DP_OP_425J2_127_3477_n1998), 
        .A2(DP_OP_423J2_125_3477_n2973), .Y(DP_OP_424J2_126_3477_n2942) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1829 ( .A1(DP_OP_422J2_124_3477_n2218), 
        .A2(DP_OP_423J2_125_3477_n2621), .Y(DP_OP_424J2_126_3477_n2590) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1792 ( .A1(DP_OP_424J2_126_3477_n2569), 
        .A2(DP_OP_424J2_126_3477_n2578), .Y(DP_OP_424J2_126_3477_n2553) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2227 ( .A1(DP_OP_423J2_125_3477_n3010), 
        .A2(DP_OP_422J2_124_3477_n3015), .Y(DP_OP_423J2_125_3477_n2986) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1477 ( .A1(DP_OP_425J2_127_3477_n2658), 
        .A2(DP_OP_424J2_126_3477_n2269), .Y(DP_OP_424J2_126_3477_n2238) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1484 ( .A1(DP_OP_424J2_126_3477_n2261), 
        .A2(DP_OP_424J2_126_3477_n2270), .Y(DP_OP_424J2_126_3477_n2245) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1581 ( .A1(DP_OP_423J2_125_3477_n2350), 
        .A2(DP_OP_423J2_125_3477_n2359), .Y(DP_OP_423J2_125_3477_n2342) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1873 ( .A1(DP_OP_424J2_126_3477_n2658), 
        .A2(DP_OP_424J2_126_3477_n2665), .Y(DP_OP_424J2_126_3477_n2634) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1697 ( .A1(DP_OP_424J2_126_3477_n2482), 
        .A2(DP_OP_424J2_126_3477_n2489), .Y(DP_OP_424J2_126_3477_n2458) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1479 ( .A1(DP_OP_425J2_127_3477_n2572), 
        .A2(DP_OP_425J2_127_3477_n2269), .Y(DP_OP_423J2_125_3477_n2240) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1741 ( .A1(DP_OP_424J2_126_3477_n2526), 
        .A2(DP_OP_424J2_126_3477_n2533), .Y(DP_OP_424J2_126_3477_n2502) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1389 ( .A1(DP_OP_422J2_124_3477_n2790), 
        .A2(DP_OP_423J2_125_3477_n2181), .Y(DP_OP_423J2_125_3477_n2150) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1961 ( .A1(DP_OP_423J2_125_3477_n2834), 
        .A2(DP_OP_424J2_126_3477_n2753), .Y(DP_OP_424J2_126_3477_n2722) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1521 ( .A1(DP_OP_422J2_124_3477_n2746), 
        .A2(DP_OP_423J2_125_3477_n2313), .Y(DP_OP_424J2_126_3477_n2282) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1880 ( .A1(DP_OP_425J2_127_3477_n2305), 
        .A2(DP_OP_424J2_126_3477_n2666), .Y(DP_OP_424J2_126_3477_n2641) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1449 ( .A1(DP_OP_423J2_125_3477_n2218), 
        .A2(DP_OP_422J2_124_3477_n2227), .Y(DP_OP_423J2_125_3477_n2210) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1653 ( .A1(DP_OP_423J2_125_3477_n2350), 
        .A2(DP_OP_424J2_126_3477_n2445), .Y(DP_OP_424J2_126_3477_n2414) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1660 ( .A1(DP_OP_425J2_127_3477_n2481), 
        .A2(DP_OP_424J2_126_3477_n2446), .Y(DP_OP_424J2_126_3477_n2421) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1917 ( .A1(DP_OP_422J2_124_3477_n2130), 
        .A2(DP_OP_422J2_124_3477_n2709), .Y(DP_OP_424J2_126_3477_n2678) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1609 ( .A1(DP_OP_425J2_127_3477_n2526), 
        .A2(DP_OP_424J2_126_3477_n2401), .Y(DP_OP_424J2_126_3477_n2370) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1616 ( .A1(DP_OP_423J2_125_3477_n2305), 
        .A2(DP_OP_424J2_126_3477_n2402), .Y(DP_OP_424J2_126_3477_n2377) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2049 ( .A1(DP_OP_424J2_126_3477_n2834), 
        .A2(DP_OP_425J2_127_3477_n2841), .Y(DP_OP_424J2_126_3477_n2810) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1345 ( .A1(DP_OP_422J2_124_3477_n2922), 
        .A2(DP_OP_424J2_126_3477_n2137), .Y(DP_OP_424J2_126_3477_n2106) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2139 ( .A1(DP_OP_423J2_125_3477_n2924), 
        .A2(DP_OP_423J2_125_3477_n2929), .Y(DP_OP_423J2_125_3477_n2900) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1352 ( .A1(DP_OP_422J2_124_3477_n2921), 
        .A2(DP_OP_425J2_127_3477_n2138), .Y(DP_OP_424J2_126_3477_n2113) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1433 ( .A1(DP_OP_424J2_126_3477_n2218), 
        .A2(DP_OP_424J2_126_3477_n2225), .Y(DP_OP_424J2_126_3477_n2194) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1222 ( .A1(DP_OP_425J2_127_3477_n2835), 
        .A2(DP_OP_423J2_125_3477_n2006), .Y(DP_OP_423J2_125_3477_n1983) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2012 ( .A1(DP_OP_424J2_126_3477_n2789), 
        .A2(DP_OP_425J2_127_3477_n2798), .Y(DP_OP_424J2_126_3477_n2773) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1389 ( .A1(DP_OP_423J2_125_3477_n2086), 
        .A2(DP_OP_425J2_127_3477_n2181), .Y(DP_OP_424J2_126_3477_n2150) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1396 ( .A1(DP_OP_425J2_127_3477_n2745), 
        .A2(DP_OP_424J2_126_3477_n2182), .Y(DP_OP_424J2_126_3477_n2157) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1257 ( .A1(DP_OP_422J2_124_3477_n3008), 
        .A2(DP_OP_424J2_126_3477_n2049), .Y(DP_OP_424J2_126_3477_n2018) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2056 ( .A1(DP_OP_424J2_126_3477_n2833), 
        .A2(DP_OP_425J2_127_3477_n2842), .Y(DP_OP_424J2_126_3477_n2817) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2146 ( .A1(DP_OP_423J2_125_3477_n2923), 
        .A2(DP_OP_423J2_125_3477_n2930), .Y(DP_OP_423J2_125_3477_n2907) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1301 ( .A1(DP_OP_423J2_125_3477_n1998), 
        .A2(DP_OP_425J2_127_3477_n2093), .Y(DP_OP_424J2_126_3477_n2062) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1924 ( .A1(DP_OP_422J2_124_3477_n2129), 
        .A2(DP_OP_425J2_127_3477_n2710), .Y(DP_OP_424J2_126_3477_n2685) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1565 ( .A1(DP_OP_422J2_124_3477_n2702), 
        .A2(DP_OP_424J2_126_3477_n2357), .Y(DP_OP_424J2_126_3477_n2326) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2153 ( .A1(DP_OP_423J2_125_3477_n2922), 
        .A2(DP_OP_423J2_125_3477_n2931), .Y(DP_OP_423J2_125_3477_n2914) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1572 ( .A1(DP_OP_422J2_124_3477_n2701), 
        .A2(DP_OP_424J2_126_3477_n2358), .Y(DP_OP_424J2_126_3477_n2333) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1397 ( .A1(DP_OP_425J2_127_3477_n2658), 
        .A2(DP_OP_422J2_124_3477_n2182), .Y(DP_OP_423J2_125_3477_n2158) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1658 ( .A1(DP_OP_422J2_124_3477_n2531), 
        .A2(DP_OP_423J2_125_3477_n2445), .Y(DP_OP_423J2_125_3477_n2419) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1621 ( .A1(DP_OP_423J2_125_3477_n2398), 
        .A2(DP_OP_423J2_125_3477_n2402), .Y(DP_OP_423J2_125_3477_n2382) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1628 ( .A1(DP_OP_423J2_125_3477_n2397), 
        .A2(DP_OP_423J2_125_3477_n2403), .Y(DP_OP_423J2_125_3477_n2389) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1390 ( .A1(DP_OP_423J2_125_3477_n2175), 
        .A2(DP_OP_423J2_125_3477_n2181), .Y(DP_OP_423J2_125_3477_n2151) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1614 ( .A1(DP_OP_422J2_124_3477_n2575), 
        .A2(DP_OP_423J2_125_3477_n2401), .Y(DP_OP_423J2_125_3477_n2375) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2054 ( .A1(DP_OP_422J2_124_3477_n2971), 
        .A2(DP_OP_423J2_125_3477_n2841), .Y(DP_OP_425J2_127_3477_n2815) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2061 ( .A1(DP_OP_424J2_126_3477_n2090), 
        .A2(DP_OP_425J2_127_3477_n2842), .Y(DP_OP_425J2_127_3477_n2822) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1577 ( .A1(DP_OP_423J2_125_3477_n2354), 
        .A2(DP_OP_423J2_125_3477_n2358), .Y(DP_OP_423J2_125_3477_n2338) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1584 ( .A1(DP_OP_423J2_125_3477_n2353), 
        .A2(DP_OP_423J2_125_3477_n2359), .Y(DP_OP_423J2_125_3477_n2345) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1265 ( .A1(DP_OP_425J2_127_3477_n2790), 
        .A2(DP_OP_423J2_125_3477_n2050), .Y(DP_OP_423J2_125_3477_n2026) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2202 ( .A1(DP_OP_422J2_124_3477_n2971), 
        .A2(DP_OP_422J2_124_3477_n2975), .Y(DP_OP_422J2_124_3477_n2963) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1526 ( .A1(DP_OP_424J2_126_3477_n2663), 
        .A2(DP_OP_425J2_127_3477_n2313), .Y(DP_OP_425J2_127_3477_n2287) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1489 ( .A1(DP_OP_423J2_125_3477_n2794), 
        .A2(DP_OP_425J2_127_3477_n2270), .Y(DP_OP_425J2_127_3477_n2250) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2114 ( .A1(DP_OP_422J2_124_3477_n2883), 
        .A2(DP_OP_422J2_124_3477_n2887), .Y(DP_OP_422J2_124_3477_n2875) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1496 ( .A1(DP_OP_423J2_125_3477_n2793), 
        .A2(DP_OP_425J2_127_3477_n2271), .Y(DP_OP_425J2_127_3477_n2257) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1482 ( .A1(DP_OP_423J2_125_3477_n2795), 
        .A2(DP_OP_425J2_127_3477_n2269), .Y(DP_OP_425J2_127_3477_n2243) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1258 ( .A1(DP_OP_425J2_127_3477_n2791), 
        .A2(DP_OP_424J2_126_3477_n2049), .Y(DP_OP_423J2_125_3477_n2019) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1452 ( .A1(DP_OP_424J2_126_3477_n2749), 
        .A2(DP_OP_425J2_127_3477_n2227), .Y(DP_OP_425J2_127_3477_n2213) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2158 ( .A1(DP_OP_422J2_124_3477_n2927), 
        .A2(DP_OP_422J2_124_3477_n2931), .Y(DP_OP_422J2_124_3477_n2919) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1797 ( .A1(DP_OP_423J2_125_3477_n2266), 
        .A2(DP_OP_425J2_127_3477_n2578), .Y(DP_OP_425J2_127_3477_n2558) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2142 ( .A1(DP_OP_425J2_127_3477_n2927), 
        .A2(DP_OP_425J2_127_3477_n2929), .Y(DP_OP_425J2_127_3477_n2903) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2105 ( .A1(DP_OP_423J2_125_3477_n1958), 
        .A2(DP_OP_424J2_126_3477_n2886), .Y(DP_OP_425J2_127_3477_n2866) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2156 ( .A1(DP_OP_424J2_126_3477_n2001), 
        .A2(DP_OP_425J2_127_3477_n2931), .Y(DP_OP_425J2_127_3477_n2917) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1753 ( .A1(DP_OP_425J2_127_3477_n2530), 
        .A2(DP_OP_425J2_127_3477_n2534), .Y(DP_OP_425J2_127_3477_n2514) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1878 ( .A1(DP_OP_425J2_127_3477_n2663), 
        .A2(DP_OP_425J2_127_3477_n2665), .Y(DP_OP_425J2_127_3477_n2639) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1661 ( .A1(DP_OP_422J2_124_3477_n2526), 
        .A2(DP_OP_423J2_125_3477_n2446), .Y(DP_OP_423J2_125_3477_n2422) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1394 ( .A1(DP_OP_424J2_126_3477_n2795), 
        .A2(DP_OP_425J2_127_3477_n2181), .Y(DP_OP_425J2_127_3477_n2155) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1410 ( .A1(DP_OP_422J2_124_3477_n2179), 
        .A2(DP_OP_422J2_124_3477_n2183), .Y(DP_OP_422J2_124_3477_n2171) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1357 ( .A1(DP_OP_425J2_127_3477_n2134), 
        .A2(DP_OP_425J2_127_3477_n2138), .Y(DP_OP_425J2_127_3477_n2118) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1350 ( .A1(DP_OP_425J2_127_3477_n2135), 
        .A2(DP_OP_425J2_127_3477_n2137), .Y(DP_OP_425J2_127_3477_n2111) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2193 ( .A1(DP_OP_424J2_126_3477_n1958), 
        .A2(DP_OP_425J2_127_3477_n2974), .Y(DP_OP_425J2_127_3477_n2954) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1454 ( .A1(DP_OP_425J2_127_3477_n2355), 
        .A2(DP_OP_422J2_124_3477_n2227), .Y(DP_OP_422J2_124_3477_n2215) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1716 ( .A1(DP_OP_422J2_124_3477_n2617), 
        .A2(DP_OP_425J2_127_3477_n2491), .Y(DP_OP_425J2_127_3477_n2477) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1936 ( .A1(DP_OP_425J2_127_3477_n2705), 
        .A2(DP_OP_425J2_127_3477_n2711), .Y(DP_OP_425J2_127_3477_n2697) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1306 ( .A1(DP_OP_423J2_125_3477_n2971), 
        .A2(DP_OP_425J2_127_3477_n2093), .Y(DP_OP_425J2_127_3477_n2067) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1269 ( .A1(DP_OP_423J2_125_3477_n3012), 
        .A2(DP_OP_425J2_127_3477_n2050), .Y(DP_OP_425J2_127_3477_n2030) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1654 ( .A1(DP_OP_423J2_125_3477_n2439), 
        .A2(DP_OP_423J2_125_3477_n2445), .Y(DP_OP_423J2_125_3477_n2415) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1262 ( .A1(DP_OP_425J2_127_3477_n2047), 
        .A2(DP_OP_425J2_127_3477_n2049), .Y(DP_OP_425J2_127_3477_n2023) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1762 ( .A1(DP_OP_422J2_124_3477_n2531), 
        .A2(DP_OP_422J2_124_3477_n2535), .Y(DP_OP_422J2_124_3477_n2523) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1225 ( .A1(DP_OP_424J2_126_3477_n2970), 
        .A2(DP_OP_425J2_127_3477_n2006), .Y(DP_OP_425J2_127_3477_n1986) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1232 ( .A1(DP_OP_424J2_126_3477_n2969), 
        .A2(DP_OP_425J2_127_3477_n2007), .Y(DP_OP_425J2_127_3477_n1993) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2230 ( .A1(DP_OP_425J2_127_3477_n3013), 
        .A2(DP_OP_425J2_127_3477_n3015), .Y(DP_OP_425J2_127_3477_n2989) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1850 ( .A1(DP_OP_422J2_124_3477_n2619), 
        .A2(DP_OP_422J2_124_3477_n2623), .Y(DP_OP_422J2_124_3477_n2611) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1665 ( .A1(DP_OP_425J2_127_3477_n2442), 
        .A2(DP_OP_425J2_127_3477_n2446), .Y(DP_OP_425J2_127_3477_n2426) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1892 ( .A1(DP_OP_424J2_126_3477_n2265), 
        .A2(DP_OP_425J2_127_3477_n2667), .Y(DP_OP_425J2_127_3477_n2653) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2024 ( .A1(DP_OP_425J2_127_3477_n2793), 
        .A2(DP_OP_425J2_127_3477_n2799), .Y(DP_OP_425J2_127_3477_n2785) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2246 ( .A1(DP_OP_422J2_124_3477_n3013), 
        .A2(DP_OP_422J2_124_3477_n3017), .Y(DP_OP_422J2_124_3477_n3005) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2017 ( .A1(DP_OP_425J2_127_3477_n2794), 
        .A2(DP_OP_425J2_127_3477_n2798), .Y(DP_OP_425J2_127_3477_n2778) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2068 ( .A1(DP_OP_425J2_127_3477_n2837), 
        .A2(DP_OP_425J2_127_3477_n2843), .Y(DP_OP_425J2_127_3477_n2829) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1174 ( .A1(DP_OP_424J2_126_3477_n3013), 
        .A2(DP_OP_425J2_127_3477_n1961), .Y(DP_OP_425J2_127_3477_n1935) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2026 ( .A1(DP_OP_422J2_124_3477_n2795), 
        .A2(DP_OP_422J2_124_3477_n2799), .Y(DP_OP_422J2_124_3477_n2787) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1181 ( .A1(DP_OP_424J2_126_3477_n3012), 
        .A2(DP_OP_424J2_126_3477_n1962), .Y(DP_OP_425J2_127_3477_n1942) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1218 ( .A1(DP_OP_425J2_127_3477_n2003), 
        .A2(DP_OP_425J2_127_3477_n2005), .Y(DP_OP_425J2_127_3477_n1979) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2237 ( .A1(DP_OP_425J2_127_3477_n3012), 
        .A2(DP_OP_423J2_125_3477_n3016), .Y(DP_OP_425J2_127_3477_n2996) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2070 ( .A1(DP_OP_423J2_125_3477_n2135), 
        .A2(DP_OP_422J2_124_3477_n2843), .Y(DP_OP_422J2_124_3477_n2831) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2244 ( .A1(DP_OP_425J2_127_3477_n3011), 
        .A2(DP_OP_425J2_127_3477_n3017), .Y(DP_OP_425J2_127_3477_n3003) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1929 ( .A1(DP_OP_422J2_124_3477_n2838), 
        .A2(DP_OP_425J2_127_3477_n2710), .Y(DP_OP_425J2_127_3477_n2690) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2189 ( .A1(DP_OP_424J2_126_3477_n2878), 
        .A2(DP_OP_423J2_125_3477_n2974), .Y(DP_OP_423J2_125_3477_n2950) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1542 ( .A1(DP_OP_422J2_124_3477_n2311), 
        .A2(DP_OP_422J2_124_3477_n2315), .Y(DP_OP_422J2_124_3477_n2303) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2186 ( .A1(DP_OP_425J2_127_3477_n2971), 
        .A2(DP_OP_425J2_127_3477_n2973), .Y(DP_OP_425J2_127_3477_n2947) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1746 ( .A1(DP_OP_423J2_125_3477_n2311), 
        .A2(DP_OP_424J2_126_3477_n2533), .Y(DP_OP_425J2_127_3477_n2507) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1966 ( .A1(DP_OP_424J2_126_3477_n2179), 
        .A2(DP_OP_424J2_126_3477_n2753), .Y(DP_OP_425J2_127_3477_n2727) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1498 ( .A1(DP_OP_422J2_124_3477_n2267), 
        .A2(DP_OP_422J2_124_3477_n2271), .Y(DP_OP_422J2_124_3477_n2259) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1570 ( .A1(DP_OP_425J2_127_3477_n2355), 
        .A2(DP_OP_425J2_127_3477_n2357), .Y(DP_OP_425J2_127_3477_n2331) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1540 ( .A1(DP_OP_422J2_124_3477_n2177), 
        .A2(DP_OP_425J2_127_3477_n2315), .Y(DP_OP_425J2_127_3477_n2301) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1710 ( .A1(DP_OP_423J2_125_3477_n2355), 
        .A2(DP_OP_425J2_127_3477_n2490), .Y(DP_OP_425J2_127_3477_n2471) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1586 ( .A1(DP_OP_422J2_124_3477_n2355), 
        .A2(DP_OP_422J2_124_3477_n2359), .Y(DP_OP_422J2_124_3477_n2347) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1672 ( .A1(DP_OP_425J2_127_3477_n2441), 
        .A2(DP_OP_425J2_127_3477_n2447), .Y(DP_OP_425J2_127_3477_n2433) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2200 ( .A1(DP_OP_424J2_126_3477_n1957), 
        .A2(DP_OP_425J2_127_3477_n2975), .Y(DP_OP_425J2_127_3477_n2961) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1885 ( .A1(DP_OP_425J2_127_3477_n2662), 
        .A2(DP_OP_425J2_127_3477_n2666), .Y(DP_OP_425J2_127_3477_n2646) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1834 ( .A1(DP_OP_425J2_127_3477_n2619), 
        .A2(DP_OP_425J2_127_3477_n2621), .Y(DP_OP_425J2_127_3477_n2595) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2112 ( .A1(DP_OP_423J2_125_3477_n1957), 
        .A2(DP_OP_425J2_127_3477_n2887), .Y(DP_OP_425J2_127_3477_n2873) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1234 ( .A1(DP_OP_423J2_125_3477_n2003), 
        .A2(DP_OP_423J2_125_3477_n2007), .Y(DP_OP_423J2_125_3477_n1995) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1438 ( .A1(DP_OP_424J2_126_3477_n2751), 
        .A2(DP_OP_423J2_125_3477_n2225), .Y(DP_OP_425J2_127_3477_n2199) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1401 ( .A1(DP_OP_425J2_127_3477_n2178), 
        .A2(DP_OP_425J2_127_3477_n2182), .Y(DP_OP_425J2_127_3477_n2162) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1408 ( .A1(DP_OP_424J2_126_3477_n2793), 
        .A2(DP_OP_423J2_125_3477_n2183), .Y(DP_OP_425J2_127_3477_n2169) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2149 ( .A1(DP_OP_425J2_127_3477_n2926), 
        .A2(DP_OP_425J2_127_3477_n2930), .Y(DP_OP_425J2_127_3477_n2910) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1760 ( .A1(DP_OP_425J2_127_3477_n2529), 
        .A2(DP_OP_425J2_127_3477_n2535), .Y(DP_OP_425J2_127_3477_n2521) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1848 ( .A1(DP_OP_425J2_127_3477_n2617), 
        .A2(DP_OP_425J2_127_3477_n2623), .Y(DP_OP_425J2_127_3477_n2609) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1709 ( .A1(DP_OP_423J2_125_3477_n2354), 
        .A2(DP_OP_425J2_127_3477_n2490), .Y(DP_OP_425J2_127_3477_n2470) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1702 ( .A1(DP_OP_423J2_125_3477_n2355), 
        .A2(DP_OP_425J2_127_3477_n2489), .Y(DP_OP_425J2_127_3477_n2463) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1922 ( .A1(DP_OP_425J2_127_3477_n2707), 
        .A2(DP_OP_425J2_127_3477_n2709), .Y(DP_OP_425J2_127_3477_n2683) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1658 ( .A1(DP_OP_423J2_125_3477_n2619), 
        .A2(DP_OP_425J2_127_3477_n2445), .Y(DP_OP_425J2_127_3477_n2419) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2069 ( .A1(DP_OP_422J2_124_3477_n2090), 
        .A2(DP_OP_423J2_125_3477_n2843), .Y(DP_OP_423J2_125_3477_n2830) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1621 ( .A1(DP_OP_425J2_127_3477_n2398), 
        .A2(DP_OP_425J2_127_3477_n2402), .Y(DP_OP_425J2_127_3477_n2382) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1573 ( .A1(DP_OP_423J2_125_3477_n2350), 
        .A2(DP_OP_423J2_125_3477_n2358), .Y(DP_OP_423J2_125_3477_n2334) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1628 ( .A1(DP_OP_425J2_127_3477_n2397), 
        .A2(DP_OP_425J2_127_3477_n2403), .Y(DP_OP_425J2_127_3477_n2389) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1614 ( .A1(DP_OP_422J2_124_3477_n2267), 
        .A2(DP_OP_425J2_127_3477_n2401), .Y(DP_OP_425J2_127_3477_n2375) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1577 ( .A1(DP_OP_425J2_127_3477_n2354), 
        .A2(DP_OP_425J2_127_3477_n2358), .Y(DP_OP_425J2_127_3477_n2338) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1584 ( .A1(DP_OP_425J2_127_3477_n2353), 
        .A2(DP_OP_425J2_127_3477_n2359), .Y(DP_OP_425J2_127_3477_n2345) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1674 ( .A1(DP_OP_423J2_125_3477_n2487), 
        .A2(DP_OP_422J2_124_3477_n2447), .Y(DP_OP_422J2_124_3477_n2435) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2226 ( .A1(DP_OP_423J2_125_3477_n3009), 
        .A2(DP_OP_424J2_126_3477_n3015), .Y(DP_OP_423J2_125_3477_n2985) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1630 ( .A1(DP_OP_423J2_125_3477_n2531), 
        .A2(DP_OP_422J2_124_3477_n2403), .Y(DP_OP_422J2_124_3477_n2391) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1718 ( .A1(DP_OP_422J2_124_3477_n2487), 
        .A2(DP_OP_422J2_124_3477_n2491), .Y(DP_OP_422J2_124_3477_n2479) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1938 ( .A1(DP_OP_422J2_124_3477_n2707), 
        .A2(DP_OP_422J2_124_3477_n2711), .Y(DP_OP_422J2_124_3477_n2699) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1894 ( .A1(DP_OP_422J2_124_3477_n2663), 
        .A2(DP_OP_422J2_124_3477_n2667), .Y(DP_OP_422J2_124_3477_n2655) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1761 ( .A1(DP_OP_423J2_125_3477_n2530), 
        .A2(DP_OP_423J2_125_3477_n2535), .Y(DP_OP_423J2_125_3477_n2522) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1717 ( .A1(DP_OP_422J2_124_3477_n2442), 
        .A2(DP_OP_423J2_125_3477_n2491), .Y(DP_OP_423J2_125_3477_n2478) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1234 ( .A1(DP_OP_425J2_127_3477_n2003), 
        .A2(DP_OP_425J2_127_3477_n2007), .Y(DP_OP_425J2_127_3477_n1995) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2069 ( .A1(DP_OP_422J2_124_3477_n2970), 
        .A2(DP_OP_425J2_127_3477_n2843), .Y(DP_OP_425J2_127_3477_n2830) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1754 ( .A1(DP_OP_423J2_125_3477_n2531), 
        .A2(DP_OP_423J2_125_3477_n2534), .Y(DP_OP_423J2_125_3477_n2515) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1346 ( .A1(DP_OP_422J2_124_3477_n2835), 
        .A2(DP_OP_425J2_127_3477_n2137), .Y(DP_OP_423J2_125_3477_n2107) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1578 ( .A1(DP_OP_423J2_125_3477_n2355), 
        .A2(DP_OP_423J2_125_3477_n2358), .Y(DP_OP_423J2_125_3477_n2339) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1761 ( .A1(DP_OP_425J2_127_3477_n2530), 
        .A2(DP_OP_425J2_127_3477_n2535), .Y(DP_OP_425J2_127_3477_n2522) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1541 ( .A1(DP_OP_422J2_124_3477_n2662), 
        .A2(DP_OP_423J2_125_3477_n2315), .Y(DP_OP_423J2_125_3477_n2302) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1717 ( .A1(DP_OP_424J2_126_3477_n2442), 
        .A2(DP_OP_425J2_127_3477_n2491), .Y(DP_OP_425J2_127_3477_n2478) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1754 ( .A1(DP_OP_423J2_125_3477_n2311), 
        .A2(DP_OP_425J2_127_3477_n2534), .Y(DP_OP_425J2_127_3477_n2515) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1578 ( .A1(DP_OP_425J2_127_3477_n2355), 
        .A2(DP_OP_425J2_127_3477_n2358), .Y(DP_OP_425J2_127_3477_n2339) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1497 ( .A1(DP_OP_423J2_125_3477_n2266), 
        .A2(DP_OP_425J2_127_3477_n2271), .Y(DP_OP_423J2_125_3477_n2258) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1541 ( .A1(DP_OP_423J2_125_3477_n2750), 
        .A2(DP_OP_425J2_127_3477_n2315), .Y(DP_OP_425J2_127_3477_n2302) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1353 ( .A1(DP_OP_424J2_126_3477_n2218), 
        .A2(DP_OP_423J2_125_3477_n2138), .Y(DP_OP_423J2_125_3477_n2114) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1497 ( .A1(DP_OP_423J2_125_3477_n2794), 
        .A2(DP_OP_425J2_127_3477_n2271), .Y(DP_OP_425J2_127_3477_n2258) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1453 ( .A1(DP_OP_422J2_124_3477_n2090), 
        .A2(DP_OP_425J2_127_3477_n2227), .Y(DP_OP_425J2_127_3477_n2214) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1453 ( .A1(DP_OP_424J2_126_3477_n2310), 
        .A2(DP_OP_422J2_124_3477_n2227), .Y(DP_OP_423J2_125_3477_n2214) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1490 ( .A1(DP_OP_423J2_125_3477_n2795), 
        .A2(DP_OP_425J2_127_3477_n2270), .Y(DP_OP_425J2_127_3477_n2251) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1402 ( .A1(DP_OP_422J2_124_3477_n2047), 
        .A2(DP_OP_425J2_127_3477_n2182), .Y(DP_OP_425J2_127_3477_n2163) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1409 ( .A1(DP_OP_425J2_127_3477_n2178), 
        .A2(DP_OP_422J2_124_3477_n2183), .Y(DP_OP_425J2_127_3477_n2170) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1490 ( .A1(DP_OP_423J2_125_3477_n2267), 
        .A2(DP_OP_423J2_125_3477_n2270), .Y(DP_OP_423J2_125_3477_n2251) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2194 ( .A1(DP_OP_425J2_127_3477_n2971), 
        .A2(DP_OP_425J2_127_3477_n2974), .Y(DP_OP_425J2_127_3477_n2955) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2201 ( .A1(DP_OP_424J2_126_3477_n1958), 
        .A2(DP_OP_425J2_127_3477_n2975), .Y(DP_OP_425J2_127_3477_n2962) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2018 ( .A1(DP_OP_425J2_127_3477_n2795), 
        .A2(DP_OP_425J2_127_3477_n2798), .Y(DP_OP_425J2_127_3477_n2779) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1358 ( .A1(DP_OP_425J2_127_3477_n2135), 
        .A2(DP_OP_425J2_127_3477_n2138), .Y(DP_OP_425J2_127_3477_n2119) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1402 ( .A1(DP_OP_422J2_124_3477_n2795), 
        .A2(DP_OP_425J2_127_3477_n2182), .Y(DP_OP_423J2_125_3477_n2163) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2238 ( .A1(DP_OP_425J2_127_3477_n3013), 
        .A2(DP_OP_423J2_125_3477_n3016), .Y(DP_OP_425J2_127_3477_n2997) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1798 ( .A1(DP_OP_423J2_125_3477_n2267), 
        .A2(DP_OP_425J2_127_3477_n2578), .Y(DP_OP_425J2_127_3477_n2559) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2245 ( .A1(DP_OP_425J2_127_3477_n3012), 
        .A2(DP_OP_425J2_127_3477_n3017), .Y(DP_OP_425J2_127_3477_n3004) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1409 ( .A1(DP_OP_423J2_125_3477_n2178), 
        .A2(DP_OP_423J2_125_3477_n2183), .Y(DP_OP_423J2_125_3477_n2170) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1830 ( .A1(DP_OP_422J2_124_3477_n2307), 
        .A2(DP_OP_423J2_125_3477_n2621), .Y(DP_OP_423J2_125_3477_n2591) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2150 ( .A1(DP_OP_425J2_127_3477_n2927), 
        .A2(DP_OP_425J2_127_3477_n2930), .Y(DP_OP_425J2_127_3477_n2911) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2157 ( .A1(DP_OP_425J2_127_3477_n2926), 
        .A2(DP_OP_425J2_127_3477_n2931), .Y(DP_OP_425J2_127_3477_n2918) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1937 ( .A1(DP_OP_423J2_125_3477_n2134), 
        .A2(DP_OP_425J2_127_3477_n2711), .Y(DP_OP_425J2_127_3477_n2698) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2194 ( .A1(DP_OP_423J2_125_3477_n2971), 
        .A2(DP_OP_423J2_125_3477_n2974), .Y(DP_OP_423J2_125_3477_n2955) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1270 ( .A1(DP_OP_425J2_127_3477_n2047), 
        .A2(DP_OP_425J2_127_3477_n2050), .Y(DP_OP_425J2_127_3477_n2031) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2201 ( .A1(DP_OP_423J2_125_3477_n2970), 
        .A2(DP_OP_425J2_127_3477_n2975), .Y(DP_OP_423J2_125_3477_n2962) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1922 ( .A1(DP_OP_423J2_125_3477_n2707), 
        .A2(DP_OP_423J2_125_3477_n2709), .Y(DP_OP_423J2_125_3477_n2683) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2198 ( .A1(DP_OP_423J2_125_3477_n2967), 
        .A2(DP_OP_422J2_124_3477_n2975), .Y(DP_OP_423J2_125_3477_n2959) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2156 ( .A1(DP_OP_424J2_126_3477_n2837), 
        .A2(DP_OP_423J2_125_3477_n2931), .Y(DP_OP_423J2_125_3477_n2917) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1753 ( .A1(DP_OP_423J2_125_3477_n2530), 
        .A2(DP_OP_423J2_125_3477_n2534), .Y(DP_OP_423J2_125_3477_n2514) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1260 ( .A1(DP_OP_425J2_127_3477_n2793), 
        .A2(DP_OP_425J2_127_3477_n2049), .Y(DP_OP_423J2_125_3477_n2021) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1878 ( .A1(DP_OP_423J2_125_3477_n2663), 
        .A2(DP_OP_423J2_125_3477_n2665), .Y(DP_OP_423J2_125_3477_n2639) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1394 ( .A1(DP_OP_425J2_127_3477_n2663), 
        .A2(DP_OP_423J2_125_3477_n2181), .Y(DP_OP_423J2_125_3477_n2155) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1267 ( .A1(DP_OP_423J2_125_3477_n2044), 
        .A2(DP_OP_423J2_125_3477_n2050), .Y(DP_OP_423J2_125_3477_n2028) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1481 ( .A1(DP_OP_423J2_125_3477_n2794), 
        .A2(DP_OP_425J2_127_3477_n2269), .Y(DP_OP_425J2_127_3477_n2242) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1357 ( .A1(DP_OP_423J2_125_3477_n2134), 
        .A2(DP_OP_423J2_125_3477_n2138), .Y(DP_OP_423J2_125_3477_n2118) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1451 ( .A1(DP_OP_425J2_127_3477_n2220), 
        .A2(DP_OP_425J2_127_3477_n2227), .Y(DP_OP_425J2_127_3477_n2212) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1796 ( .A1(DP_OP_423J2_125_3477_n2265), 
        .A2(DP_OP_425J2_127_3477_n2578), .Y(DP_OP_425J2_127_3477_n2557) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1437 ( .A1(DP_OP_422J2_124_3477_n2090), 
        .A2(DP_OP_424J2_126_3477_n2225), .Y(DP_OP_425J2_127_3477_n2198) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2067 ( .A1(DP_OP_423J2_125_3477_n2000), 
        .A2(DP_OP_425J2_127_3477_n2843), .Y(DP_OP_425J2_127_3477_n2828) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1350 ( .A1(DP_OP_423J2_125_3477_n2135), 
        .A2(DP_OP_424J2_126_3477_n2137), .Y(DP_OP_423J2_125_3477_n2111) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2199 ( .A1(DP_OP_424J2_126_3477_n1956), 
        .A2(DP_OP_425J2_127_3477_n2975), .Y(DP_OP_425J2_127_3477_n2960) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1349 ( .A1(DP_OP_425J2_127_3477_n2134), 
        .A2(DP_OP_425J2_127_3477_n2137), .Y(DP_OP_425J2_127_3477_n2110) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1715 ( .A1(DP_OP_425J2_127_3477_n2484), 
        .A2(DP_OP_425J2_127_3477_n2491), .Y(DP_OP_425J2_127_3477_n2476) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1964 ( .A1(DP_OP_423J2_125_3477_n2749), 
        .A2(DP_OP_423J2_125_3477_n2753), .Y(DP_OP_423J2_125_3477_n2725) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2229 ( .A1(DP_OP_425J2_127_3477_n3012), 
        .A2(DP_OP_425J2_127_3477_n3015), .Y(DP_OP_425J2_127_3477_n2988) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2236 ( .A1(DP_OP_425J2_127_3477_n3011), 
        .A2(DP_OP_424J2_126_3477_n3016), .Y(DP_OP_425J2_127_3477_n2995) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1752 ( .A1(DP_OP_425J2_127_3477_n2529), 
        .A2(DP_OP_425J2_127_3477_n2534), .Y(DP_OP_425J2_127_3477_n2513) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1539 ( .A1(DP_OP_425J2_127_3477_n2308), 
        .A2(DP_OP_425J2_127_3477_n2315), .Y(DP_OP_425J2_127_3477_n2300) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2053 ( .A1(DP_OP_424J2_126_3477_n2090), 
        .A2(DP_OP_423J2_125_3477_n2841), .Y(DP_OP_425J2_127_3477_n2814) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2060 ( .A1(DP_OP_425J2_127_3477_n2837), 
        .A2(DP_OP_425J2_127_3477_n2842), .Y(DP_OP_425J2_127_3477_n2821) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2193 ( .A1(DP_OP_423J2_125_3477_n2970), 
        .A2(DP_OP_423J2_125_3477_n2974), .Y(DP_OP_423J2_125_3477_n2954) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1670 ( .A1(DP_OP_423J2_125_3477_n2439), 
        .A2(DP_OP_425J2_127_3477_n2447), .Y(DP_OP_423J2_125_3477_n2431) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1407 ( .A1(DP_OP_422J2_124_3477_n2044), 
        .A2(DP_OP_422J2_124_3477_n2183), .Y(DP_OP_425J2_127_3477_n2168) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1400 ( .A1(DP_OP_424J2_126_3477_n2793), 
        .A2(DP_OP_425J2_127_3477_n2182), .Y(DP_OP_425J2_127_3477_n2161) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1708 ( .A1(DP_OP_422J2_124_3477_n2617), 
        .A2(DP_OP_425J2_127_3477_n2490), .Y(DP_OP_425J2_127_3477_n2469) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1716 ( .A1(DP_OP_422J2_124_3477_n2441), 
        .A2(DP_OP_423J2_125_3477_n2491), .Y(DP_OP_423J2_125_3477_n2477) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1393 ( .A1(DP_OP_425J2_127_3477_n2178), 
        .A2(DP_OP_425J2_127_3477_n2181), .Y(DP_OP_425J2_127_3477_n2154) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2185 ( .A1(DP_OP_424J2_126_3477_n1958), 
        .A2(DP_OP_425J2_127_3477_n2973), .Y(DP_OP_425J2_127_3477_n2946) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1936 ( .A1(DP_OP_423J2_125_3477_n2705), 
        .A2(DP_OP_422J2_124_3477_n2711), .Y(DP_OP_423J2_125_3477_n2697) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1935 ( .A1(DP_OP_425J2_127_3477_n2704), 
        .A2(DP_OP_425J2_127_3477_n2711), .Y(DP_OP_425J2_127_3477_n2696) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1965 ( .A1(DP_OP_425J2_127_3477_n2750), 
        .A2(DP_OP_423J2_125_3477_n2753), .Y(DP_OP_425J2_127_3477_n2726) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1576 ( .A1(DP_OP_425J2_127_3477_n2353), 
        .A2(DP_OP_425J2_127_3477_n2358), .Y(DP_OP_425J2_127_3477_n2337) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1306 ( .A1(DP_OP_424J2_126_3477_n2179), 
        .A2(DP_OP_423J2_125_3477_n2093), .Y(DP_OP_423J2_125_3477_n2067) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1700 ( .A1(DP_OP_422J2_124_3477_n2441), 
        .A2(DP_OP_423J2_125_3477_n2489), .Y(DP_OP_423J2_125_3477_n2461) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1269 ( .A1(DP_OP_425J2_127_3477_n2794), 
        .A2(DP_OP_423J2_125_3477_n2050), .Y(DP_OP_423J2_125_3477_n2030) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1877 ( .A1(DP_OP_425J2_127_3477_n2662), 
        .A2(DP_OP_425J2_127_3477_n2665), .Y(DP_OP_425J2_127_3477_n2638) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1876 ( .A1(DP_OP_425J2_127_3477_n2397), 
        .A2(DP_OP_423J2_125_3477_n2665), .Y(DP_OP_423J2_125_3477_n2637) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1884 ( .A1(DP_OP_422J2_124_3477_n2793), 
        .A2(DP_OP_425J2_127_3477_n2666), .Y(DP_OP_425J2_127_3477_n2645) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1262 ( .A1(DP_OP_425J2_127_3477_n2795), 
        .A2(DP_OP_424J2_126_3477_n2049), .Y(DP_OP_423J2_125_3477_n2023) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1627 ( .A1(DP_OP_425J2_127_3477_n2396), 
        .A2(DP_OP_425J2_127_3477_n2403), .Y(DP_OP_425J2_127_3477_n2388) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1891 ( .A1(DP_OP_422J2_124_3477_n2792), 
        .A2(DP_OP_425J2_127_3477_n2667), .Y(DP_OP_425J2_127_3477_n2652) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1225 ( .A1(DP_OP_424J2_126_3477_n2090), 
        .A2(DP_OP_423J2_125_3477_n2006), .Y(DP_OP_423J2_125_3477_n1986) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2192 ( .A1(DP_OP_424J2_126_3477_n1957), 
        .A2(DP_OP_425J2_127_3477_n2974), .Y(DP_OP_425J2_127_3477_n2953) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1356 ( .A1(DP_OP_425J2_127_3477_n2133), 
        .A2(DP_OP_425J2_127_3477_n2138), .Y(DP_OP_425J2_127_3477_n2117) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1745 ( .A1(DP_OP_425J2_127_3477_n2530), 
        .A2(DP_OP_423J2_125_3477_n2533), .Y(DP_OP_425J2_127_3477_n2506) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1232 ( .A1(DP_OP_422J2_124_3477_n2969), 
        .A2(DP_OP_423J2_125_3477_n2007), .Y(DP_OP_423J2_125_3477_n1993) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2016 ( .A1(DP_OP_425J2_127_3477_n2793), 
        .A2(DP_OP_425J2_127_3477_n2798), .Y(DP_OP_425J2_127_3477_n2777) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1657 ( .A1(DP_OP_425J2_127_3477_n2442), 
        .A2(DP_OP_425J2_127_3477_n2445), .Y(DP_OP_425J2_127_3477_n2418) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2230 ( .A1(DP_OP_425J2_127_3477_n2047), 
        .A2(DP_OP_424J2_126_3477_n3015), .Y(DP_OP_423J2_125_3477_n2989) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1890 ( .A1(DP_OP_423J2_125_3477_n2659), 
        .A2(DP_OP_423J2_125_3477_n2667), .Y(DP_OP_423J2_125_3477_n2651) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1583 ( .A1(DP_OP_422J2_124_3477_n2220), 
        .A2(DP_OP_425J2_127_3477_n2359), .Y(DP_OP_425J2_127_3477_n2344) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1665 ( .A1(DP_OP_423J2_125_3477_n2442), 
        .A2(DP_OP_423J2_125_3477_n2446), .Y(DP_OP_423J2_125_3477_n2426) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1928 ( .A1(DP_OP_425J2_127_3477_n2705), 
        .A2(DP_OP_425J2_127_3477_n2710), .Y(DP_OP_425J2_127_3477_n2689) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1847 ( .A1(DP_OP_425J2_127_3477_n2616), 
        .A2(DP_OP_425J2_127_3477_n2623), .Y(DP_OP_425J2_127_3477_n2608) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1892 ( .A1(DP_OP_425J2_127_3477_n2397), 
        .A2(DP_OP_423J2_125_3477_n2667), .Y(DP_OP_423J2_125_3477_n2653) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1525 ( .A1(DP_OP_423J2_125_3477_n2750), 
        .A2(DP_OP_425J2_127_3477_n2313), .Y(DP_OP_425J2_127_3477_n2286) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2104 ( .A1(DP_OP_423J2_125_3477_n1957), 
        .A2(DP_OP_423J2_125_3477_n2886), .Y(DP_OP_425J2_127_3477_n2865) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1671 ( .A1(DP_OP_422J2_124_3477_n2308), 
        .A2(DP_OP_425J2_127_3477_n2447), .Y(DP_OP_425J2_127_3477_n2432) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2024 ( .A1(DP_OP_423J2_125_3477_n2793), 
        .A2(DP_OP_425J2_127_3477_n2799), .Y(DP_OP_423J2_125_3477_n2785) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2148 ( .A1(DP_OP_424J2_126_3477_n2001), 
        .A2(DP_OP_425J2_127_3477_n2930), .Y(DP_OP_425J2_127_3477_n2909) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1758 ( .A1(DP_OP_423J2_125_3477_n2527), 
        .A2(DP_OP_423J2_125_3477_n2535), .Y(DP_OP_423J2_125_3477_n2519) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1495 ( .A1(DP_OP_425J2_127_3477_n2264), 
        .A2(DP_OP_425J2_127_3477_n2271), .Y(DP_OP_425J2_127_3477_n2256) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1833 ( .A1(DP_OP_424J2_126_3477_n2310), 
        .A2(DP_OP_425J2_127_3477_n2621), .Y(DP_OP_425J2_127_3477_n2594) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2017 ( .A1(DP_OP_423J2_125_3477_n2794), 
        .A2(DP_OP_423J2_125_3477_n2798), .Y(DP_OP_423J2_125_3477_n2778) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1613 ( .A1(DP_OP_425J2_127_3477_n2398), 
        .A2(DP_OP_425J2_127_3477_n2401), .Y(DP_OP_425J2_127_3477_n2374) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2068 ( .A1(DP_OP_423J2_125_3477_n2837), 
        .A2(DP_OP_423J2_125_3477_n2843), .Y(DP_OP_423J2_125_3477_n2829) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1305 ( .A1(DP_OP_423J2_125_3477_n2970), 
        .A2(DP_OP_425J2_127_3477_n2093), .Y(DP_OP_425J2_127_3477_n2066) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1268 ( .A1(DP_OP_423J2_125_3477_n3011), 
        .A2(DP_OP_425J2_127_3477_n2050), .Y(DP_OP_425J2_127_3477_n2029) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1174 ( .A1(DP_OP_424J2_126_3477_n2047), 
        .A2(DP_OP_422J2_124_3477_n1961), .Y(DP_OP_423J2_125_3477_n1935) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1920 ( .A1(DP_OP_423J2_125_3477_n2705), 
        .A2(DP_OP_423J2_125_3477_n2709), .Y(DP_OP_423J2_125_3477_n2681) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1921 ( .A1(DP_OP_423J2_125_3477_n2134), 
        .A2(DP_OP_425J2_127_3477_n2709), .Y(DP_OP_425J2_127_3477_n2682) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1181 ( .A1(DP_OP_423J2_125_3477_n1958), 
        .A2(DP_OP_423J2_125_3477_n1962), .Y(DP_OP_423J2_125_3477_n1942) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1620 ( .A1(DP_OP_425J2_127_3477_n2397), 
        .A2(DP_OP_425J2_127_3477_n2402), .Y(DP_OP_425J2_127_3477_n2381) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1701 ( .A1(DP_OP_424J2_126_3477_n2442), 
        .A2(DP_OP_425J2_127_3477_n2489), .Y(DP_OP_425J2_127_3477_n2462) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2023 ( .A1(DP_OP_423J2_125_3477_n2044), 
        .A2(DP_OP_425J2_127_3477_n2799), .Y(DP_OP_425J2_127_3477_n2784) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1218 ( .A1(DP_OP_423J2_125_3477_n2003), 
        .A2(DP_OP_423J2_125_3477_n2005), .Y(DP_OP_423J2_125_3477_n1979) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1569 ( .A1(DP_OP_425J2_127_3477_n2354), 
        .A2(DP_OP_425J2_127_3477_n2357), .Y(DP_OP_425J2_127_3477_n2330) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1664 ( .A1(DP_OP_425J2_127_3477_n2441), 
        .A2(DP_OP_425J2_127_3477_n2446), .Y(DP_OP_425J2_127_3477_n2425) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2237 ( .A1(DP_OP_423J2_125_3477_n3012), 
        .A2(DP_OP_423J2_125_3477_n3016), .Y(DP_OP_423J2_125_3477_n2996) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2243 ( .A1(DP_OP_425J2_127_3477_n3010), 
        .A2(DP_OP_425J2_127_3477_n3017), .Y(DP_OP_425J2_127_3477_n3002) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2244 ( .A1(DP_OP_423J2_125_3477_n3011), 
        .A2(DP_OP_423J2_125_3477_n3017), .Y(DP_OP_423J2_125_3477_n3003) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2111 ( .A1(DP_OP_424J2_126_3477_n2044), 
        .A2(DP_OP_425J2_127_3477_n2887), .Y(DP_OP_425J2_127_3477_n2872) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2141 ( .A1(DP_OP_425J2_127_3477_n2926), 
        .A2(DP_OP_425J2_127_3477_n2929), .Y(DP_OP_425J2_127_3477_n2902) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1759 ( .A1(DP_OP_425J2_127_3477_n2528), 
        .A2(DP_OP_425J2_127_3477_n2535), .Y(DP_OP_425J2_127_3477_n2520) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1929 ( .A1(DP_OP_424J2_126_3477_n2618), 
        .A2(DP_OP_423J2_125_3477_n2710), .Y(DP_OP_423J2_125_3477_n2690) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2145 ( .A1(DP_OP_423J2_125_3477_n2922), 
        .A2(DP_OP_423J2_125_3477_n2930), .Y(DP_OP_423J2_125_3477_n2906) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2186 ( .A1(DP_OP_423J2_125_3477_n2971), 
        .A2(DP_OP_423J2_125_3477_n2973), .Y(DP_OP_423J2_125_3477_n2947) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1261 ( .A1(DP_OP_423J2_125_3477_n3012), 
        .A2(DP_OP_425J2_127_3477_n2049), .Y(DP_OP_425J2_127_3477_n2022) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1224 ( .A1(DP_OP_424J2_126_3477_n2969), 
        .A2(DP_OP_425J2_127_3477_n2006), .Y(DP_OP_425J2_127_3477_n1985) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1231 ( .A1(DP_OP_425J2_127_3477_n2000), 
        .A2(DP_OP_425J2_127_3477_n2007), .Y(DP_OP_425J2_127_3477_n1992) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1746 ( .A1(DP_OP_423J2_125_3477_n2531), 
        .A2(DP_OP_423J2_125_3477_n2533), .Y(DP_OP_423J2_125_3477_n2507) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1173 ( .A1(DP_OP_424J2_126_3477_n3012), 
        .A2(DP_OP_425J2_127_3477_n1961), .Y(DP_OP_425J2_127_3477_n1934) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1180 ( .A1(DP_OP_424J2_126_3477_n3011), 
        .A2(DP_OP_423J2_125_3477_n1962), .Y(DP_OP_425J2_127_3477_n1941) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1217 ( .A1(DP_OP_424J2_126_3477_n2970), 
        .A2(DP_OP_425J2_127_3477_n2005), .Y(DP_OP_425J2_127_3477_n1978) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1966 ( .A1(DP_OP_422J2_124_3477_n2179), 
        .A2(DP_OP_423J2_125_3477_n2753), .Y(DP_OP_423J2_125_3477_n2727) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1488 ( .A1(DP_OP_423J2_125_3477_n2793), 
        .A2(DP_OP_425J2_127_3477_n2270), .Y(DP_OP_425J2_127_3477_n2249) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2155 ( .A1(DP_OP_425J2_127_3477_n2924), 
        .A2(DP_OP_425J2_127_3477_n2931), .Y(DP_OP_425J2_127_3477_n2916) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1570 ( .A1(DP_OP_423J2_125_3477_n2355), 
        .A2(DP_OP_423J2_125_3477_n2357), .Y(DP_OP_423J2_125_3477_n2331) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1540 ( .A1(DP_OP_424J2_126_3477_n2397), 
        .A2(DP_OP_423J2_125_3477_n2315), .Y(DP_OP_423J2_125_3477_n2301) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1672 ( .A1(DP_OP_423J2_125_3477_n2441), 
        .A2(DP_OP_422J2_124_3477_n2447), .Y(DP_OP_423J2_125_3477_n2433) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2200 ( .A1(DP_OP_423J2_125_3477_n2969), 
        .A2(DP_OP_425J2_127_3477_n2975), .Y(DP_OP_423J2_125_3477_n2961) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1885 ( .A1(DP_OP_423J2_125_3477_n2662), 
        .A2(DP_OP_424J2_126_3477_n2666), .Y(DP_OP_423J2_125_3477_n2646) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2182 ( .A1(DP_OP_423J2_125_3477_n2967), 
        .A2(DP_OP_423J2_125_3477_n2973), .Y(DP_OP_423J2_125_3477_n2943) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1834 ( .A1(DP_OP_423J2_125_3477_n2619), 
        .A2(DP_OP_423J2_125_3477_n2621), .Y(DP_OP_423J2_125_3477_n2595) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2112 ( .A1(DP_OP_422J2_124_3477_n2045), 
        .A2(DP_OP_425J2_127_3477_n2887), .Y(DP_OP_423J2_125_3477_n2873) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1438 ( .A1(DP_OP_425J2_127_3477_n2619), 
        .A2(DP_OP_423J2_125_3477_n2225), .Y(DP_OP_423J2_125_3477_n2199) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1401 ( .A1(DP_OP_423J2_125_3477_n2178), 
        .A2(DP_OP_424J2_126_3477_n2182), .Y(DP_OP_423J2_125_3477_n2162) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1408 ( .A1(DP_OP_424J2_126_3477_n2265), 
        .A2(DP_OP_423J2_125_3477_n2183), .Y(DP_OP_423J2_125_3477_n2169) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2149 ( .A1(DP_OP_423J2_125_3477_n2926), 
        .A2(DP_OP_423J2_125_3477_n2930), .Y(DP_OP_423J2_125_3477_n2910) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1760 ( .A1(DP_OP_423J2_125_3477_n2529), 
        .A2(DP_OP_423J2_125_3477_n2535), .Y(DP_OP_423J2_125_3477_n2521) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1848 ( .A1(DP_OP_423J2_125_3477_n2617), 
        .A2(DP_OP_423J2_125_3477_n2623), .Y(DP_OP_423J2_125_3477_n2609) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1709 ( .A1(DP_OP_422J2_124_3477_n2442), 
        .A2(DP_OP_423J2_125_3477_n2490), .Y(DP_OP_423J2_125_3477_n2470) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1702 ( .A1(DP_OP_423J2_125_3477_n2487), 
        .A2(DP_OP_423J2_125_3477_n2489), .Y(DP_OP_423J2_125_3477_n2463) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1666 ( .A1(DP_OP_422J2_124_3477_n2311), 
        .A2(DP_OP_425J2_127_3477_n2446), .Y(DP_OP_425J2_127_3477_n2427) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1182 ( .A1(DP_OP_423J2_125_3477_n2971), 
        .A2(DP_OP_422J2_124_3477_n1962), .Y(DP_OP_422J2_124_3477_n1943) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1233 ( .A1(DP_OP_425J2_127_3477_n2134), 
        .A2(DP_OP_422J2_124_3477_n2007), .Y(DP_OP_422J2_124_3477_n1994) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2138 ( .A1(DP_OP_423J2_125_3477_n2923), 
        .A2(DP_OP_423J2_125_3477_n2929), .Y(DP_OP_423J2_125_3477_n2899) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1930 ( .A1(DP_OP_422J2_124_3477_n2707), 
        .A2(DP_OP_422J2_124_3477_n2710), .Y(DP_OP_422J2_124_3477_n2691) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2113 ( .A1(DP_OP_425J2_127_3477_n2750), 
        .A2(DP_OP_422J2_124_3477_n2887), .Y(DP_OP_422J2_124_3477_n2874) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1849 ( .A1(DP_OP_423J2_125_3477_n2354), 
        .A2(DP_OP_422J2_124_3477_n2623), .Y(DP_OP_422J2_124_3477_n2610) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2025 ( .A1(DP_OP_423J2_125_3477_n2794), 
        .A2(DP_OP_425J2_127_3477_n2799), .Y(DP_OP_423J2_125_3477_n2786) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1566 ( .A1(DP_OP_423J2_125_3477_n2351), 
        .A2(DP_OP_423J2_125_3477_n2357), .Y(DP_OP_423J2_125_3477_n2327) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1673 ( .A1(DP_OP_422J2_124_3477_n2442), 
        .A2(DP_OP_422J2_124_3477_n2447), .Y(DP_OP_422J2_124_3477_n2434) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1610 ( .A1(DP_OP_422J2_124_3477_n2571), 
        .A2(DP_OP_423J2_125_3477_n2401), .Y(DP_OP_423J2_125_3477_n2371) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1666 ( .A1(DP_OP_423J2_125_3477_n2487), 
        .A2(DP_OP_422J2_124_3477_n2446), .Y(DP_OP_422J2_124_3477_n2427) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1710 ( .A1(DP_OP_422J2_124_3477_n2487), 
        .A2(DP_OP_422J2_124_3477_n2490), .Y(DP_OP_422J2_124_3477_n2471) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1270 ( .A1(DP_OP_422J2_124_3477_n2047), 
        .A2(DP_OP_422J2_124_3477_n2050), .Y(DP_OP_422J2_124_3477_n2031) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1937 ( .A1(DP_OP_424J2_126_3477_n2354), 
        .A2(DP_OP_422J2_124_3477_n2711), .Y(DP_OP_422J2_124_3477_n2698) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2157 ( .A1(DP_OP_422J2_124_3477_n2926), 
        .A2(DP_OP_422J2_124_3477_n2931), .Y(DP_OP_422J2_124_3477_n2918) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1962 ( .A1(DP_OP_423J2_125_3477_n2747), 
        .A2(DP_OP_423J2_125_3477_n2753), .Y(DP_OP_423J2_125_3477_n2723) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2150 ( .A1(DP_OP_422J2_124_3477_n2927), 
        .A2(DP_OP_422J2_124_3477_n2930), .Y(DP_OP_422J2_124_3477_n2911) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2245 ( .A1(DP_OP_422J2_124_3477_n3012), 
        .A2(DP_OP_422J2_124_3477_n3017), .Y(DP_OP_422J2_124_3477_n3004) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1798 ( .A1(DP_OP_422J2_124_3477_n2575), 
        .A2(DP_OP_422J2_124_3477_n2578), .Y(DP_OP_422J2_124_3477_n2559) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1434 ( .A1(DP_OP_423J2_125_3477_n2219), 
        .A2(DP_OP_423J2_125_3477_n2225), .Y(DP_OP_423J2_125_3477_n2195) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2238 ( .A1(DP_OP_422J2_124_3477_n3013), 
        .A2(DP_OP_422J2_124_3477_n3016), .Y(DP_OP_422J2_124_3477_n2997) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1404 ( .A1(DP_OP_424J2_126_3477_n2261), 
        .A2(DP_OP_423J2_125_3477_n2183), .Y(DP_OP_423J2_125_3477_n2165) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1358 ( .A1(DP_OP_422J2_124_3477_n2135), 
        .A2(DP_OP_422J2_124_3477_n2138), .Y(DP_OP_422J2_124_3477_n2119) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2062 ( .A1(DP_OP_422J2_124_3477_n2091), 
        .A2(DP_OP_423J2_125_3477_n2842), .Y(DP_OP_423J2_125_3477_n2823) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2018 ( .A1(DP_OP_422J2_124_3477_n2795), 
        .A2(DP_OP_422J2_124_3477_n2798), .Y(DP_OP_422J2_124_3477_n2779) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2201 ( .A1(DP_OP_422J2_124_3477_n2970), 
        .A2(DP_OP_422J2_124_3477_n2975), .Y(DP_OP_422J2_124_3477_n2962) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2194 ( .A1(DP_OP_422J2_124_3477_n2971), 
        .A2(DP_OP_422J2_124_3477_n2974), .Y(DP_OP_422J2_124_3477_n2955) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1894 ( .A1(DP_OP_423J2_125_3477_n2663), 
        .A2(DP_OP_423J2_125_3477_n2667), .Y(DP_OP_423J2_125_3477_n2655) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1696 ( .A1(DP_OP_422J2_124_3477_n2481), 
        .A2(DP_OP_422J2_124_3477_n2489), .Y(DP_OP_422J2_124_3477_n2457) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1881 ( .A1(DP_OP_423J2_125_3477_n2658), 
        .A2(DP_OP_422J2_124_3477_n2666), .Y(DP_OP_423J2_125_3477_n2642) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1938 ( .A1(DP_OP_423J2_125_3477_n2707), 
        .A2(DP_OP_425J2_127_3477_n2711), .Y(DP_OP_423J2_125_3477_n2699) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1608 ( .A1(DP_OP_423J2_125_3477_n2525), 
        .A2(DP_OP_422J2_124_3477_n2401), .Y(DP_OP_422J2_124_3477_n2369) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1409 ( .A1(DP_OP_422J2_124_3477_n2178), 
        .A2(DP_OP_422J2_124_3477_n2183), .Y(DP_OP_422J2_124_3477_n2170) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1170 ( .A1(DP_OP_425J2_127_3477_n2879), 
        .A2(DP_OP_424J2_126_3477_n1961), .Y(DP_OP_423J2_125_3477_n1931) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1520 ( .A1(DP_OP_422J2_124_3477_n2305), 
        .A2(DP_OP_422J2_124_3477_n2313), .Y(DP_OP_422J2_124_3477_n2281) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1402 ( .A1(DP_OP_422J2_124_3477_n2179), 
        .A2(DP_OP_422J2_124_3477_n2182), .Y(DP_OP_422J2_124_3477_n2163) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2136 ( .A1(DP_OP_422J2_124_3477_n2921), 
        .A2(DP_OP_422J2_124_3477_n2929), .Y(DP_OP_422J2_124_3477_n2897) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1388 ( .A1(DP_OP_425J2_127_3477_n2305), 
        .A2(DP_OP_422J2_124_3477_n2181), .Y(DP_OP_422J2_124_3477_n2149) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1718 ( .A1(DP_OP_423J2_125_3477_n2487), 
        .A2(DP_OP_423J2_125_3477_n2491), .Y(DP_OP_423J2_125_3477_n2479) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1300 ( .A1(DP_OP_424J2_126_3477_n2745), 
        .A2(DP_OP_422J2_124_3477_n2093), .Y(DP_OP_422J2_124_3477_n2061) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1698 ( .A1(DP_OP_422J2_124_3477_n2439), 
        .A2(DP_OP_423J2_125_3477_n2489), .Y(DP_OP_423J2_125_3477_n2459) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1490 ( .A1(DP_OP_422J2_124_3477_n2267), 
        .A2(DP_OP_422J2_124_3477_n2270), .Y(DP_OP_422J2_124_3477_n2251) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1828 ( .A1(DP_OP_422J2_124_3477_n2613), 
        .A2(DP_OP_422J2_124_3477_n2621), .Y(DP_OP_422J2_124_3477_n2589) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1453 ( .A1(DP_OP_424J2_126_3477_n2618), 
        .A2(DP_OP_422J2_124_3477_n2227), .Y(DP_OP_422J2_124_3477_n2214) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1960 ( .A1(DP_OP_422J2_124_3477_n2745), 
        .A2(DP_OP_422J2_124_3477_n2753), .Y(DP_OP_422J2_124_3477_n2721) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1168 ( .A1(DP_OP_425J2_127_3477_n2085), 
        .A2(DP_OP_422J2_124_3477_n1961), .Y(DP_OP_422J2_124_3477_n1929) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1497 ( .A1(DP_OP_423J2_125_3477_n2662), 
        .A2(DP_OP_422J2_124_3477_n2271), .Y(DP_OP_422J2_124_3477_n2258) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1925 ( .A1(DP_OP_423J2_125_3477_n2702), 
        .A2(DP_OP_423J2_125_3477_n2710), .Y(DP_OP_423J2_125_3477_n2686) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1541 ( .A1(DP_OP_424J2_126_3477_n2530), 
        .A2(DP_OP_422J2_124_3477_n2315), .Y(DP_OP_422J2_124_3477_n2302) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1578 ( .A1(DP_OP_422J2_124_3477_n2355), 
        .A2(DP_OP_422J2_124_3477_n2358), .Y(DP_OP_422J2_124_3477_n2339) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1793 ( .A1(DP_OP_423J2_125_3477_n2570), 
        .A2(DP_OP_422J2_124_3477_n2578), .Y(DP_OP_423J2_125_3477_n2554) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1630 ( .A1(DP_OP_422J2_124_3477_n2575), 
        .A2(DP_OP_423J2_125_3477_n2403), .Y(DP_OP_423J2_125_3477_n2391) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1754 ( .A1(DP_OP_422J2_124_3477_n2531), 
        .A2(DP_OP_422J2_124_3477_n2534), .Y(DP_OP_422J2_124_3477_n2515) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1874 ( .A1(DP_OP_423J2_125_3477_n2659), 
        .A2(DP_OP_423J2_125_3477_n2665), .Y(DP_OP_423J2_125_3477_n2635) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1717 ( .A1(DP_OP_422J2_124_3477_n2486), 
        .A2(DP_OP_422J2_124_3477_n2491), .Y(DP_OP_422J2_124_3477_n2478) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1712 ( .A1(DP_OP_423J2_125_3477_n2481), 
        .A2(DP_OP_423J2_125_3477_n2491), .Y(DP_OP_423J2_125_3477_n2473) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1761 ( .A1(DP_OP_423J2_125_3477_n2442), 
        .A2(DP_OP_422J2_124_3477_n2535), .Y(DP_OP_422J2_124_3477_n2522) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1705 ( .A1(DP_OP_423J2_125_3477_n2482), 
        .A2(DP_OP_423J2_125_3477_n2490), .Y(DP_OP_423J2_125_3477_n2466) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1674 ( .A1(DP_OP_422J2_124_3477_n2531), 
        .A2(DP_OP_425J2_127_3477_n2447), .Y(DP_OP_423J2_125_3477_n2435) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1673 ( .A1(DP_OP_425J2_127_3477_n2442), 
        .A2(DP_OP_425J2_127_3477_n2447), .Y(DP_OP_425J2_127_3477_n2434) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2018 ( .A1(DP_OP_423J2_125_3477_n2795), 
        .A2(DP_OP_423J2_125_3477_n2798), .Y(DP_OP_423J2_125_3477_n2779) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2057 ( .A1(DP_OP_423J2_125_3477_n2834), 
        .A2(DP_OP_423J2_125_3477_n2842), .Y(DP_OP_423J2_125_3477_n2818) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1849 ( .A1(DP_OP_424J2_126_3477_n2310), 
        .A2(DP_OP_425J2_127_3477_n2623), .Y(DP_OP_425J2_127_3477_n2610) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2113 ( .A1(DP_OP_423J2_125_3477_n1958), 
        .A2(DP_OP_425J2_127_3477_n2887), .Y(DP_OP_425J2_127_3477_n2874) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1930 ( .A1(DP_OP_425J2_127_3477_n2707), 
        .A2(DP_OP_425J2_127_3477_n2710), .Y(DP_OP_425J2_127_3477_n2691) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1233 ( .A1(DP_OP_424J2_126_3477_n2970), 
        .A2(DP_OP_425J2_127_3477_n2007), .Y(DP_OP_425J2_127_3477_n1994) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1182 ( .A1(DP_OP_424J2_126_3477_n3013), 
        .A2(DP_OP_422J2_124_3477_n1962), .Y(DP_OP_425J2_127_3477_n1943) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1226 ( .A1(DP_OP_425J2_127_3477_n2003), 
        .A2(DP_OP_425J2_127_3477_n2006), .Y(DP_OP_425J2_127_3477_n1987) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1629 ( .A1(DP_OP_425J2_127_3477_n2398), 
        .A2(DP_OP_425J2_127_3477_n2403), .Y(DP_OP_425J2_127_3477_n2390) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1585 ( .A1(DP_OP_425J2_127_3477_n2354), 
        .A2(DP_OP_425J2_127_3477_n2359), .Y(DP_OP_425J2_127_3477_n2346) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1622 ( .A1(DP_OP_422J2_124_3477_n2267), 
        .A2(DP_OP_425J2_127_3477_n2402), .Y(DP_OP_425J2_127_3477_n2383) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1358 ( .A1(DP_OP_423J2_125_3477_n2135), 
        .A2(DP_OP_423J2_125_3477_n2138), .Y(DP_OP_423J2_125_3477_n2119) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1893 ( .A1(DP_OP_425J2_127_3477_n2662), 
        .A2(DP_OP_425J2_127_3477_n2667), .Y(DP_OP_425J2_127_3477_n2654) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1886 ( .A1(DP_OP_425J2_127_3477_n2663), 
        .A2(DP_OP_425J2_127_3477_n2666), .Y(DP_OP_425J2_127_3477_n2647) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2106 ( .A1(DP_OP_422J2_124_3477_n3013), 
        .A2(DP_OP_424J2_126_3477_n2886), .Y(DP_OP_425J2_127_3477_n2867) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2238 ( .A1(DP_OP_425J2_127_3477_n2047), 
        .A2(DP_OP_423J2_125_3477_n3016), .Y(DP_OP_423J2_125_3477_n2997) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1478 ( .A1(DP_OP_423J2_125_3477_n2263), 
        .A2(DP_OP_424J2_126_3477_n2269), .Y(DP_OP_423J2_125_3477_n2239) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2025 ( .A1(DP_OP_425J2_127_3477_n2794), 
        .A2(DP_OP_425J2_127_3477_n2799), .Y(DP_OP_425J2_127_3477_n2786) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2062 ( .A1(DP_OP_422J2_124_3477_n2971), 
        .A2(DP_OP_425J2_127_3477_n2842), .Y(DP_OP_425J2_127_3477_n2823) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1798 ( .A1(DP_OP_423J2_125_3477_n2575), 
        .A2(DP_OP_425J2_127_3477_n2578), .Y(DP_OP_423J2_125_3477_n2559) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2245 ( .A1(DP_OP_423J2_125_3477_n3012), 
        .A2(DP_OP_423J2_125_3477_n3017), .Y(DP_OP_423J2_125_3477_n3004) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2150 ( .A1(DP_OP_423J2_125_3477_n2927), 
        .A2(DP_OP_423J2_125_3477_n2930), .Y(DP_OP_423J2_125_3477_n2911) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2064 ( .A1(DP_OP_424J2_126_3477_n2745), 
        .A2(DP_OP_423J2_125_3477_n2843), .Y(DP_OP_423J2_125_3477_n2825) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2157 ( .A1(DP_OP_423J2_125_3477_n2926), 
        .A2(DP_OP_423J2_125_3477_n2931), .Y(DP_OP_423J2_125_3477_n2918) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1937 ( .A1(DP_OP_425J2_127_3477_n2354), 
        .A2(DP_OP_422J2_124_3477_n2711), .Y(DP_OP_423J2_125_3477_n2698) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1221 ( .A1(DP_OP_423J2_125_3477_n1998), 
        .A2(DP_OP_423J2_125_3477_n2006), .Y(DP_OP_423J2_125_3477_n1982) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1270 ( .A1(DP_OP_425J2_127_3477_n2795), 
        .A2(DP_OP_423J2_125_3477_n2050), .Y(DP_OP_423J2_125_3477_n2031) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1894 ( .A1(DP_OP_425J2_127_3477_n2663), 
        .A2(DP_OP_425J2_127_3477_n2667), .Y(DP_OP_425J2_127_3477_n2655) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1938 ( .A1(DP_OP_425J2_127_3477_n2707), 
        .A2(DP_OP_425J2_127_3477_n2711), .Y(DP_OP_425J2_127_3477_n2699) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1710 ( .A1(DP_OP_423J2_125_3477_n2487), 
        .A2(DP_OP_423J2_125_3477_n2490), .Y(DP_OP_423J2_125_3477_n2471) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1718 ( .A1(DP_OP_422J2_124_3477_n2619), 
        .A2(DP_OP_425J2_127_3477_n2491), .Y(DP_OP_425J2_127_3477_n2479) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1485 ( .A1(DP_OP_423J2_125_3477_n2262), 
        .A2(DP_OP_423J2_125_3477_n2270), .Y(DP_OP_423J2_125_3477_n2246) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1630 ( .A1(DP_OP_422J2_124_3477_n2267), 
        .A2(DP_OP_425J2_127_3477_n2403), .Y(DP_OP_425J2_127_3477_n2391) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1674 ( .A1(DP_OP_422J2_124_3477_n2311), 
        .A2(DP_OP_425J2_127_3477_n2447), .Y(DP_OP_425J2_127_3477_n2435) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1666 ( .A1(DP_OP_422J2_124_3477_n2531), 
        .A2(DP_OP_423J2_125_3477_n2446), .Y(DP_OP_423J2_125_3477_n2427) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1586 ( .A1(DP_OP_425J2_127_3477_n2355), 
        .A2(DP_OP_425J2_127_3477_n2359), .Y(DP_OP_425J2_127_3477_n2347) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1673 ( .A1(DP_OP_423J2_125_3477_n2442), 
        .A2(DP_OP_424J2_126_3477_n2447), .Y(DP_OP_423J2_125_3477_n2434) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1498 ( .A1(DP_OP_423J2_125_3477_n2795), 
        .A2(DP_OP_425J2_127_3477_n2271), .Y(DP_OP_425J2_127_3477_n2259) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1542 ( .A1(DP_OP_422J2_124_3477_n2179), 
        .A2(DP_OP_425J2_127_3477_n2315), .Y(DP_OP_425J2_127_3477_n2303) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2070 ( .A1(DP_OP_423J2_125_3477_n2003), 
        .A2(DP_OP_425J2_127_3477_n2843), .Y(DP_OP_425J2_127_3477_n2831) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2026 ( .A1(DP_OP_425J2_127_3477_n2795), 
        .A2(DP_OP_425J2_127_3477_n2799), .Y(DP_OP_425J2_127_3477_n2787) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1849 ( .A1(DP_OP_424J2_126_3477_n2530), 
        .A2(DP_OP_423J2_125_3477_n2623), .Y(DP_OP_423J2_125_3477_n2610) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2246 ( .A1(DP_OP_425J2_127_3477_n3013), 
        .A2(DP_OP_425J2_127_3477_n3017), .Y(DP_OP_425J2_127_3477_n3005) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1850 ( .A1(DP_OP_425J2_127_3477_n2619), 
        .A2(DP_OP_425J2_127_3477_n2623), .Y(DP_OP_425J2_127_3477_n2611) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1762 ( .A1(DP_OP_422J2_124_3477_n2663), 
        .A2(DP_OP_425J2_127_3477_n2535), .Y(DP_OP_425J2_127_3477_n2523) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2113 ( .A1(DP_OP_424J2_126_3477_n2794), 
        .A2(DP_OP_424J2_126_3477_n2887), .Y(DP_OP_423J2_125_3477_n2874) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1749 ( .A1(DP_OP_423J2_125_3477_n2526), 
        .A2(DP_OP_423J2_125_3477_n2534), .Y(DP_OP_423J2_125_3477_n2510) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1454 ( .A1(DP_OP_422J2_124_3477_n2091), 
        .A2(DP_OP_425J2_127_3477_n2227), .Y(DP_OP_425J2_127_3477_n2215) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1410 ( .A1(DP_OP_424J2_126_3477_n2795), 
        .A2(DP_OP_423J2_125_3477_n2183), .Y(DP_OP_425J2_127_3477_n2171) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1930 ( .A1(DP_OP_423J2_125_3477_n2707), 
        .A2(DP_OP_423J2_125_3477_n2710), .Y(DP_OP_423J2_125_3477_n2691) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1233 ( .A1(DP_OP_424J2_126_3477_n2090), 
        .A2(DP_OP_423J2_125_3477_n2007), .Y(DP_OP_423J2_125_3477_n1994) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2158 ( .A1(DP_OP_425J2_127_3477_n2927), 
        .A2(DP_OP_425J2_127_3477_n2931), .Y(DP_OP_425J2_127_3477_n2919) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1742 ( .A1(DP_OP_423J2_125_3477_n2527), 
        .A2(DP_OP_423J2_125_3477_n2533), .Y(DP_OP_423J2_125_3477_n2503) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2114 ( .A1(DP_OP_424J2_126_3477_n2047), 
        .A2(DP_OP_425J2_127_3477_n2887), .Y(DP_OP_425J2_127_3477_n2875) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2202 ( .A1(DP_OP_425J2_127_3477_n2971), 
        .A2(DP_OP_425J2_127_3477_n2975), .Y(DP_OP_425J2_127_3477_n2963) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1182 ( .A1(DP_OP_422J2_124_3477_n3013), 
        .A2(DP_OP_423J2_125_3477_n1962), .Y(DP_OP_423J2_125_3477_n1943) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2062 ( .A1(DP_OP_423J2_125_3477_n2135), 
        .A2(DP_OP_422J2_124_3477_n2842), .Y(DP_OP_422J2_124_3477_n2823) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1226 ( .A1(DP_OP_425J2_127_3477_n2135), 
        .A2(DP_OP_422J2_124_3477_n2006), .Y(DP_OP_422J2_124_3477_n1987) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2025 ( .A1(DP_OP_425J2_127_3477_n2662), 
        .A2(DP_OP_422J2_124_3477_n2799), .Y(DP_OP_422J2_124_3477_n2786) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2106 ( .A1(DP_OP_422J2_124_3477_n2883), 
        .A2(DP_OP_422J2_124_3477_n2886), .Y(DP_OP_422J2_124_3477_n2867) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1886 ( .A1(DP_OP_422J2_124_3477_n2663), 
        .A2(DP_OP_422J2_124_3477_n2666), .Y(DP_OP_422J2_124_3477_n2647) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1893 ( .A1(DP_OP_422J2_124_3477_n2662), 
        .A2(DP_OP_422J2_124_3477_n2667), .Y(DP_OP_422J2_124_3477_n2654) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1226 ( .A1(DP_OP_423J2_125_3477_n2003), 
        .A2(DP_OP_423J2_125_3477_n2006), .Y(DP_OP_423J2_125_3477_n1987) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1629 ( .A1(DP_OP_423J2_125_3477_n2398), 
        .A2(DP_OP_423J2_125_3477_n2403), .Y(DP_OP_423J2_125_3477_n2390) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2101 ( .A1(DP_OP_423J2_125_3477_n2878), 
        .A2(DP_OP_423J2_125_3477_n2886), .Y(DP_OP_423J2_125_3477_n2862) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1585 ( .A1(DP_OP_423J2_125_3477_n2354), 
        .A2(DP_OP_423J2_125_3477_n2359), .Y(DP_OP_423J2_125_3477_n2346) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1622 ( .A1(DP_OP_422J2_124_3477_n2575), 
        .A2(DP_OP_423J2_125_3477_n2402), .Y(DP_OP_423J2_125_3477_n2383) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1893 ( .A1(DP_OP_423J2_125_3477_n2662), 
        .A2(DP_OP_423J2_125_3477_n2667), .Y(DP_OP_423J2_125_3477_n2654) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1886 ( .A1(DP_OP_423J2_125_3477_n2663), 
        .A2(DP_OP_425J2_127_3477_n2666), .Y(DP_OP_423J2_125_3477_n2647) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1214 ( .A1(DP_OP_425J2_127_3477_n2835), 
        .A2(DP_OP_423J2_125_3477_n2005), .Y(DP_OP_423J2_125_3477_n1975) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2106 ( .A1(DP_OP_422J2_124_3477_n2047), 
        .A2(DP_OP_423J2_125_3477_n2886), .Y(DP_OP_423J2_125_3477_n2867) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1622 ( .A1(DP_OP_423J2_125_3477_n2531), 
        .A2(DP_OP_424J2_126_3477_n2402), .Y(DP_OP_422J2_124_3477_n2383) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1585 ( .A1(DP_OP_422J2_124_3477_n2354), 
        .A2(DP_OP_422J2_124_3477_n2359), .Y(DP_OP_422J2_124_3477_n2346) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1522 ( .A1(DP_OP_423J2_125_3477_n2307), 
        .A2(DP_OP_423J2_125_3477_n2313), .Y(DP_OP_423J2_125_3477_n2283) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1629 ( .A1(DP_OP_423J2_125_3477_n2530), 
        .A2(DP_OP_422J2_124_3477_n2403), .Y(DP_OP_422J2_124_3477_n2390) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1389 ( .A1(DP_OP_423J2_125_3477_n2878), 
        .A2(DP_OP_425J2_127_3477_n2181), .Y(DP_OP_425J2_127_3477_n2150) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1433 ( .A1(DP_OP_425J2_127_3477_n2218), 
        .A2(DP_OP_422J2_124_3477_n2225), .Y(DP_OP_425J2_127_3477_n2194) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1345 ( .A1(DP_OP_424J2_126_3477_n2834), 
        .A2(DP_OP_425J2_127_3477_n2137), .Y(DP_OP_425J2_127_3477_n2106) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2049 ( .A1(DP_OP_425J2_127_3477_n2834), 
        .A2(DP_OP_425J2_127_3477_n2841), .Y(DP_OP_425J2_127_3477_n2810) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1609 ( .A1(DP_OP_422J2_124_3477_n2262), 
        .A2(DP_OP_425J2_127_3477_n2401), .Y(DP_OP_425J2_127_3477_n2370) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1917 ( .A1(DP_OP_424J2_126_3477_n2218), 
        .A2(DP_OP_425J2_127_3477_n2709), .Y(DP_OP_425J2_127_3477_n2678) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1653 ( .A1(DP_OP_425J2_127_3477_n2438), 
        .A2(DP_OP_425J2_127_3477_n2445), .Y(DP_OP_425J2_127_3477_n2414) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2103 ( .A1(DP_OP_423J2_125_3477_n2880), 
        .A2(DP_OP_423J2_125_3477_n2886), .Y(DP_OP_423J2_125_3477_n2864) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1521 ( .A1(DP_OP_423J2_125_3477_n2746), 
        .A2(DP_OP_425J2_127_3477_n2313), .Y(DP_OP_425J2_127_3477_n2282) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1961 ( .A1(DP_OP_422J2_124_3477_n2878), 
        .A2(DP_OP_424J2_126_3477_n2753), .Y(DP_OP_425J2_127_3477_n2722) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2016 ( .A1(DP_OP_423J2_125_3477_n2793), 
        .A2(DP_OP_423J2_125_3477_n2798), .Y(DP_OP_423J2_125_3477_n2777) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1741 ( .A1(DP_OP_425J2_127_3477_n2526), 
        .A2(DP_OP_422J2_124_3477_n2533), .Y(DP_OP_425J2_127_3477_n2502) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1697 ( .A1(DP_OP_425J2_127_3477_n2482), 
        .A2(DP_OP_425J2_127_3477_n2489), .Y(DP_OP_425J2_127_3477_n2458) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1873 ( .A1(DP_OP_425J2_127_3477_n2658), 
        .A2(DP_OP_425J2_127_3477_n2665), .Y(DP_OP_425J2_127_3477_n2634) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1538 ( .A1(DP_OP_423J2_125_3477_n2307), 
        .A2(DP_OP_423J2_125_3477_n2315), .Y(DP_OP_423J2_125_3477_n2299) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1477 ( .A1(DP_OP_423J2_125_3477_n2790), 
        .A2(DP_OP_425J2_127_3477_n2269), .Y(DP_OP_425J2_127_3477_n2238) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1829 ( .A1(DP_OP_422J2_124_3477_n2746), 
        .A2(DP_OP_425J2_127_3477_n2621), .Y(DP_OP_425J2_127_3477_n2590) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2181 ( .A1(DP_OP_424J2_126_3477_n1954), 
        .A2(DP_OP_425J2_127_3477_n2973), .Y(DP_OP_425J2_127_3477_n2942) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2225 ( .A1(DP_OP_425J2_127_3477_n3008), 
        .A2(DP_OP_425J2_127_3477_n3015), .Y(DP_OP_425J2_127_3477_n2984) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1169 ( .A1(DP_OP_424J2_126_3477_n3008), 
        .A2(DP_OP_425J2_127_3477_n1961), .Y(DP_OP_425J2_127_3477_n1930) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1918 ( .A1(DP_OP_422J2_124_3477_n2219), 
        .A2(DP_OP_423J2_125_3477_n2709), .Y(DP_OP_423J2_125_3477_n2679) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1657 ( .A1(DP_OP_423J2_125_3477_n2442), 
        .A2(DP_OP_423J2_125_3477_n2445), .Y(DP_OP_423J2_125_3477_n2418) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1583 ( .A1(DP_OP_422J2_124_3477_n2616), 
        .A2(DP_OP_423J2_125_3477_n2359), .Y(DP_OP_423J2_125_3477_n2344) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1928 ( .A1(DP_OP_423J2_125_3477_n2705), 
        .A2(DP_OP_423J2_125_3477_n2710), .Y(DP_OP_423J2_125_3477_n2689) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1847 ( .A1(DP_OP_422J2_124_3477_n2308), 
        .A2(DP_OP_423J2_125_3477_n2623), .Y(DP_OP_423J2_125_3477_n2608) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1525 ( .A1(DP_OP_425J2_127_3477_n2530), 
        .A2(DP_OP_423J2_125_3477_n2313), .Y(DP_OP_423J2_125_3477_n2286) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2104 ( .A1(DP_OP_422J2_124_3477_n2045), 
        .A2(DP_OP_423J2_125_3477_n2886), .Y(DP_OP_423J2_125_3477_n2865) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1671 ( .A1(DP_OP_422J2_124_3477_n2528), 
        .A2(DP_OP_422J2_124_3477_n2447), .Y(DP_OP_423J2_125_3477_n2432) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2148 ( .A1(DP_OP_424J2_126_3477_n2837), 
        .A2(DP_OP_423J2_125_3477_n2930), .Y(DP_OP_423J2_125_3477_n2909) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1495 ( .A1(DP_OP_425J2_127_3477_n2572), 
        .A2(DP_OP_425J2_127_3477_n2271), .Y(DP_OP_423J2_125_3477_n2256) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1833 ( .A1(DP_OP_424J2_126_3477_n2530), 
        .A2(DP_OP_423J2_125_3477_n2621), .Y(DP_OP_423J2_125_3477_n2594) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1613 ( .A1(DP_OP_423J2_125_3477_n2398), 
        .A2(DP_OP_423J2_125_3477_n2401), .Y(DP_OP_423J2_125_3477_n2374) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1305 ( .A1(DP_OP_425J2_127_3477_n2750), 
        .A2(DP_OP_423J2_125_3477_n2093), .Y(DP_OP_423J2_125_3477_n2066) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1268 ( .A1(DP_OP_425J2_127_3477_n2793), 
        .A2(DP_OP_423J2_125_3477_n2050), .Y(DP_OP_423J2_125_3477_n2029) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1921 ( .A1(DP_OP_425J2_127_3477_n2354), 
        .A2(DP_OP_423J2_125_3477_n2709), .Y(DP_OP_423J2_125_3477_n2682) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1620 ( .A1(DP_OP_423J2_125_3477_n2397), 
        .A2(DP_OP_423J2_125_3477_n2402), .Y(DP_OP_423J2_125_3477_n2381) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1701 ( .A1(DP_OP_422J2_124_3477_n2442), 
        .A2(DP_OP_423J2_125_3477_n2489), .Y(DP_OP_423J2_125_3477_n2462) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2023 ( .A1(DP_OP_425J2_127_3477_n2264), 
        .A2(DP_OP_424J2_126_3477_n2799), .Y(DP_OP_423J2_125_3477_n2784) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1569 ( .A1(DP_OP_423J2_125_3477_n2354), 
        .A2(DP_OP_423J2_125_3477_n2357), .Y(DP_OP_423J2_125_3477_n2330) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1304 ( .A1(DP_OP_424J2_126_3477_n2177), 
        .A2(DP_OP_423J2_125_3477_n2093), .Y(DP_OP_423J2_125_3477_n2065) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1664 ( .A1(DP_OP_423J2_125_3477_n2441), 
        .A2(DP_OP_423J2_125_3477_n2446), .Y(DP_OP_423J2_125_3477_n2425) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2243 ( .A1(DP_OP_423J2_125_3477_n3010), 
        .A2(DP_OP_423J2_125_3477_n3017), .Y(DP_OP_423J2_125_3477_n3002) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2111 ( .A1(DP_OP_423J2_125_3477_n2880), 
        .A2(DP_OP_422J2_124_3477_n2887), .Y(DP_OP_423J2_125_3477_n2872) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2141 ( .A1(DP_OP_423J2_125_3477_n2926), 
        .A2(DP_OP_423J2_125_3477_n2929), .Y(DP_OP_423J2_125_3477_n2902) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1759 ( .A1(DP_OP_423J2_125_3477_n2528), 
        .A2(DP_OP_423J2_125_3477_n2535), .Y(DP_OP_423J2_125_3477_n2520) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1302 ( .A1(DP_OP_425J2_127_3477_n2087), 
        .A2(DP_OP_425J2_127_3477_n2093), .Y(DP_OP_425J2_127_3477_n2063) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2050 ( .A1(DP_OP_425J2_127_3477_n2835), 
        .A2(DP_OP_424J2_126_3477_n2841), .Y(DP_OP_425J2_127_3477_n2811) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1172 ( .A1(DP_OP_423J2_125_3477_n1957), 
        .A2(DP_OP_425J2_127_3477_n1961), .Y(DP_OP_423J2_125_3477_n1933) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1965 ( .A1(DP_OP_423J2_125_3477_n2750), 
        .A2(DP_OP_423J2_125_3477_n2753), .Y(DP_OP_423J2_125_3477_n2726) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1480 ( .A1(DP_OP_423J2_125_3477_n2265), 
        .A2(DP_OP_425J2_127_3477_n2269), .Y(DP_OP_423J2_125_3477_n2241) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1487 ( .A1(DP_OP_425J2_127_3477_n2572), 
        .A2(DP_OP_423J2_125_3477_n2270), .Y(DP_OP_423J2_125_3477_n2248) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2183 ( .A1(DP_OP_424J2_126_3477_n1956), 
        .A2(DP_OP_425J2_127_3477_n2973), .Y(DP_OP_425J2_127_3477_n2944) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2190 ( .A1(DP_OP_425J2_127_3477_n2967), 
        .A2(DP_OP_425J2_127_3477_n2974), .Y(DP_OP_425J2_127_3477_n2951) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1574 ( .A1(DP_OP_425J2_127_3477_n2351), 
        .A2(DP_OP_425J2_127_3477_n2358), .Y(DP_OP_425J2_127_3477_n2335) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1576 ( .A1(DP_OP_423J2_125_3477_n2353), 
        .A2(DP_OP_423J2_125_3477_n2358), .Y(DP_OP_423J2_125_3477_n2337) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2197 ( .A1(DP_OP_424J2_126_3477_n1954), 
        .A2(DP_OP_425J2_127_3477_n2975), .Y(DP_OP_425J2_127_3477_n2958) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2227 ( .A1(DP_OP_425J2_127_3477_n3010), 
        .A2(DP_OP_425J2_127_3477_n3015), .Y(DP_OP_425J2_127_3477_n2986) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1581 ( .A1(DP_OP_423J2_125_3477_n2702), 
        .A2(DP_OP_425J2_127_3477_n2359), .Y(DP_OP_425J2_127_3477_n2342) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1479 ( .A1(DP_OP_425J2_127_3477_n2264), 
        .A2(DP_OP_425J2_127_3477_n2269), .Y(DP_OP_425J2_127_3477_n2240) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1449 ( .A1(DP_OP_425J2_127_3477_n2218), 
        .A2(DP_OP_425J2_127_3477_n2227), .Y(DP_OP_425J2_127_3477_n2210) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2139 ( .A1(DP_OP_425J2_127_3477_n2924), 
        .A2(DP_OP_425J2_127_3477_n2929), .Y(DP_OP_425J2_127_3477_n2900) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1222 ( .A1(DP_OP_424J2_126_3477_n2967), 
        .A2(DP_OP_425J2_127_3477_n2006), .Y(DP_OP_425J2_127_3477_n1983) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2146 ( .A1(DP_OP_425J2_127_3477_n2923), 
        .A2(DP_OP_425J2_127_3477_n2930), .Y(DP_OP_425J2_127_3477_n2907) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2153 ( .A1(DP_OP_425J2_127_3477_n2922), 
        .A2(DP_OP_425J2_127_3477_n2931), .Y(DP_OP_425J2_127_3477_n2914) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1537 ( .A1(DP_OP_423J2_125_3477_n2746), 
        .A2(DP_OP_425J2_127_3477_n2315), .Y(DP_OP_425J2_127_3477_n2298) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1743 ( .A1(DP_OP_425J2_127_3477_n2528), 
        .A2(DP_OP_424J2_126_3477_n2533), .Y(DP_OP_425J2_127_3477_n2504) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1713 ( .A1(DP_OP_425J2_127_3477_n2482), 
        .A2(DP_OP_425J2_127_3477_n2491), .Y(DP_OP_425J2_127_3477_n2474) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1926 ( .A1(DP_OP_422J2_124_3477_n2835), 
        .A2(DP_OP_425J2_127_3477_n2710), .Y(DP_OP_425J2_127_3477_n2687) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1229 ( .A1(DP_OP_425J2_127_3477_n1998), 
        .A2(DP_OP_425J2_127_3477_n2007), .Y(DP_OP_425J2_127_3477_n1990) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1493 ( .A1(DP_OP_423J2_125_3477_n2790), 
        .A2(DP_OP_425J2_127_3477_n2271), .Y(DP_OP_425J2_127_3477_n2254) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2102 ( .A1(DP_OP_425J2_127_3477_n2879), 
        .A2(DP_OP_422J2_124_3477_n2886), .Y(DP_OP_425J2_127_3477_n2863) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2109 ( .A1(DP_OP_425J2_127_3477_n2878), 
        .A2(DP_OP_425J2_127_3477_n2887), .Y(DP_OP_425J2_127_3477_n2870) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1523 ( .A1(DP_OP_425J2_127_3477_n2308), 
        .A2(DP_OP_425J2_127_3477_n2313), .Y(DP_OP_425J2_127_3477_n2284) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1435 ( .A1(DP_OP_425J2_127_3477_n2220), 
        .A2(DP_OP_423J2_125_3477_n2225), .Y(DP_OP_425J2_127_3477_n2196) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2234 ( .A1(DP_OP_425J2_127_3477_n3009), 
        .A2(DP_OP_424J2_126_3477_n3016), .Y(DP_OP_425J2_127_3477_n2993) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1215 ( .A1(DP_OP_425J2_127_3477_n2000), 
        .A2(DP_OP_425J2_127_3477_n2005), .Y(DP_OP_425J2_127_3477_n1976) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1625 ( .A1(DP_OP_422J2_124_3477_n2262), 
        .A2(DP_OP_425J2_127_3477_n2403), .Y(DP_OP_425J2_127_3477_n2386) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1875 ( .A1(DP_OP_424J2_126_3477_n2264), 
        .A2(DP_OP_425J2_127_3477_n2665), .Y(DP_OP_425J2_127_3477_n2636) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1882 ( .A1(DP_OP_423J2_125_3477_n2175), 
        .A2(DP_OP_425J2_127_3477_n2666), .Y(DP_OP_425J2_127_3477_n2643) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1889 ( .A1(DP_OP_425J2_127_3477_n2658), 
        .A2(DP_OP_425J2_127_3477_n2667), .Y(DP_OP_425J2_127_3477_n2650) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1405 ( .A1(DP_OP_423J2_125_3477_n2878), 
        .A2(DP_OP_423J2_125_3477_n2183), .Y(DP_OP_425J2_127_3477_n2166) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1398 ( .A1(DP_OP_425J2_127_3477_n2175), 
        .A2(DP_OP_425J2_127_3477_n2182), .Y(DP_OP_425J2_127_3477_n2159) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1877 ( .A1(DP_OP_423J2_125_3477_n2662), 
        .A2(DP_OP_423J2_125_3477_n2665), .Y(DP_OP_423J2_125_3477_n2638) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1757 ( .A1(DP_OP_425J2_127_3477_n2526), 
        .A2(DP_OP_425J2_127_3477_n2535), .Y(DP_OP_425J2_127_3477_n2518) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1750 ( .A1(DP_OP_422J2_124_3477_n2659), 
        .A2(DP_OP_425J2_127_3477_n2534), .Y(DP_OP_425J2_127_3477_n2511) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1919 ( .A1(DP_OP_425J2_127_3477_n2704), 
        .A2(DP_OP_425J2_127_3477_n2709), .Y(DP_OP_425J2_127_3477_n2680) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1669 ( .A1(DP_OP_425J2_127_3477_n2438), 
        .A2(DP_OP_425J2_127_3477_n2447), .Y(DP_OP_425J2_127_3477_n2430) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1662 ( .A1(DP_OP_425J2_127_3477_n2439), 
        .A2(DP_OP_425J2_127_3477_n2446), .Y(DP_OP_425J2_127_3477_n2423) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1963 ( .A1(DP_OP_422J2_124_3477_n2880), 
        .A2(DP_OP_422J2_124_3477_n2753), .Y(DP_OP_425J2_127_3477_n2724) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1178 ( .A1(DP_OP_424J2_126_3477_n3009), 
        .A2(DP_OP_423J2_125_3477_n1962), .Y(DP_OP_425J2_127_3477_n1939) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1611 ( .A1(DP_OP_425J2_127_3477_n2396), 
        .A2(DP_OP_425J2_127_3477_n2401), .Y(DP_OP_425J2_127_3477_n2372) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1845 ( .A1(DP_OP_422J2_124_3477_n2746), 
        .A2(DP_OP_425J2_127_3477_n2623), .Y(DP_OP_425J2_127_3477_n2606) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1831 ( .A1(DP_OP_425J2_127_3477_n2616), 
        .A2(DP_OP_425J2_127_3477_n2621), .Y(DP_OP_425J2_127_3477_n2592) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1391 ( .A1(DP_OP_422J2_124_3477_n2044), 
        .A2(DP_OP_425J2_127_3477_n2181), .Y(DP_OP_425J2_127_3477_n2152) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2014 ( .A1(DP_OP_425J2_127_3477_n2791), 
        .A2(DP_OP_425J2_127_3477_n2798), .Y(DP_OP_425J2_127_3477_n2775) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1884 ( .A1(DP_OP_425J2_127_3477_n2397), 
        .A2(DP_OP_424J2_126_3477_n2666), .Y(DP_OP_423J2_125_3477_n2645) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1171 ( .A1(DP_OP_424J2_126_3477_n3010), 
        .A2(DP_OP_425J2_127_3477_n1961), .Y(DP_OP_425J2_127_3477_n1932) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2241 ( .A1(DP_OP_425J2_127_3477_n3008), 
        .A2(DP_OP_425J2_127_3477_n3017), .Y(DP_OP_425J2_127_3477_n3000) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1618 ( .A1(DP_OP_423J2_125_3477_n2659), 
        .A2(DP_OP_425J2_127_3477_n2402), .Y(DP_OP_425J2_127_3477_n2379) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1794 ( .A1(DP_OP_423J2_125_3477_n2263), 
        .A2(DP_OP_425J2_127_3477_n2578), .Y(DP_OP_425J2_127_3477_n2555) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2065 ( .A1(DP_OP_425J2_127_3477_n2834), 
        .A2(DP_OP_425J2_127_3477_n2843), .Y(DP_OP_425J2_127_3477_n2826) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1567 ( .A1(DP_OP_424J2_126_3477_n2616), 
        .A2(DP_OP_425J2_127_3477_n2357), .Y(DP_OP_425J2_127_3477_n2328) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1354 ( .A1(DP_OP_423J2_125_3477_n2923), 
        .A2(DP_OP_425J2_127_3477_n2138), .Y(DP_OP_425J2_127_3477_n2115) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1347 ( .A1(DP_OP_423J2_125_3477_n2924), 
        .A2(DP_OP_425J2_127_3477_n2137), .Y(DP_OP_425J2_127_3477_n2108) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2021 ( .A1(DP_OP_425J2_127_3477_n2790), 
        .A2(DP_OP_425J2_127_3477_n2799), .Y(DP_OP_425J2_127_3477_n2782) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1266 ( .A1(DP_OP_423J2_125_3477_n3009), 
        .A2(DP_OP_425J2_127_3477_n2050), .Y(DP_OP_425J2_127_3477_n2027) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1259 ( .A1(DP_OP_423J2_125_3477_n3010), 
        .A2(DP_OP_425J2_127_3477_n2049), .Y(DP_OP_425J2_127_3477_n2020) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1486 ( .A1(DP_OP_423J2_125_3477_n2791), 
        .A2(DP_OP_425J2_127_3477_n2270), .Y(DP_OP_425J2_127_3477_n2247) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1706 ( .A1(DP_OP_424J2_126_3477_n2439), 
        .A2(DP_OP_425J2_127_3477_n2490), .Y(DP_OP_425J2_127_3477_n2467) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1699 ( .A1(DP_OP_425J2_127_3477_n2484), 
        .A2(DP_OP_425J2_127_3477_n2489), .Y(DP_OP_425J2_127_3477_n2460) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1933 ( .A1(DP_OP_422J2_124_3477_n2834), 
        .A2(DP_OP_425J2_127_3477_n2711), .Y(DP_OP_425J2_127_3477_n2694) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2051 ( .A1(DP_OP_424J2_126_3477_n2088), 
        .A2(DP_OP_424J2_126_3477_n2841), .Y(DP_OP_425J2_127_3477_n2812) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1303 ( .A1(DP_OP_425J2_127_3477_n2088), 
        .A2(DP_OP_425J2_127_3477_n2093), .Y(DP_OP_425J2_127_3477_n2064) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1568 ( .A1(DP_OP_423J2_125_3477_n2353), 
        .A2(DP_OP_423J2_125_3477_n2357), .Y(DP_OP_423J2_125_3477_n2329) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2058 ( .A1(DP_OP_425J2_127_3477_n2835), 
        .A2(DP_OP_425J2_127_3477_n2842), .Y(DP_OP_425J2_127_3477_n2819) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1655 ( .A1(DP_OP_424J2_126_3477_n2528), 
        .A2(DP_OP_425J2_127_3477_n2445), .Y(DP_OP_425J2_127_3477_n2416) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1627 ( .A1(DP_OP_423J2_125_3477_n2396), 
        .A2(DP_OP_423J2_125_3477_n2403), .Y(DP_OP_423J2_125_3477_n2388) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1891 ( .A1(DP_OP_424J2_126_3477_n2572), 
        .A2(DP_OP_423J2_125_3477_n2667), .Y(DP_OP_423J2_125_3477_n2652) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2192 ( .A1(DP_OP_423J2_125_3477_n2969), 
        .A2(DP_OP_423J2_125_3477_n2974), .Y(DP_OP_423J2_125_3477_n2953) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1356 ( .A1(DP_OP_425J2_127_3477_n2705), 
        .A2(DP_OP_423J2_125_3477_n2138), .Y(DP_OP_423J2_125_3477_n2117) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1213 ( .A1(DP_OP_425J2_127_3477_n1998), 
        .A2(DP_OP_425J2_127_3477_n2005), .Y(DP_OP_425J2_127_3477_n1974) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2100 ( .A1(DP_OP_425J2_127_3477_n2877), 
        .A2(DP_OP_423J2_125_3477_n2886), .Y(DP_OP_425J2_127_3477_n2861) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2137 ( .A1(DP_OP_425J2_127_3477_n2922), 
        .A2(DP_OP_425J2_127_3477_n2929), .Y(DP_OP_425J2_127_3477_n2898) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1572 ( .A1(DP_OP_424J2_126_3477_n2613), 
        .A2(DP_OP_425J2_127_3477_n2358), .Y(DP_OP_425J2_127_3477_n2333) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1565 ( .A1(DP_OP_423J2_125_3477_n2702), 
        .A2(DP_OP_425J2_127_3477_n2357), .Y(DP_OP_425J2_127_3477_n2326) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1301 ( .A1(DP_OP_425J2_127_3477_n2086), 
        .A2(DP_OP_425J2_127_3477_n2093), .Y(DP_OP_425J2_127_3477_n2062) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2056 ( .A1(DP_OP_425J2_127_3477_n2833), 
        .A2(DP_OP_425J2_127_3477_n2842), .Y(DP_OP_425J2_127_3477_n2817) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1745 ( .A1(DP_OP_423J2_125_3477_n2530), 
        .A2(DP_OP_423J2_125_3477_n2533), .Y(DP_OP_423J2_125_3477_n2506) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2110 ( .A1(DP_OP_425J2_127_3477_n2175), 
        .A2(DP_OP_424J2_126_3477_n2887), .Y(DP_OP_423J2_125_3477_n2871) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1257 ( .A1(DP_OP_423J2_125_3477_n3008), 
        .A2(DP_OP_425J2_127_3477_n2049), .Y(DP_OP_425J2_127_3477_n2018) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1925 ( .A1(DP_OP_422J2_124_3477_n2834), 
        .A2(DP_OP_425J2_127_3477_n2710), .Y(DP_OP_425J2_127_3477_n2686) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1793 ( .A1(DP_OP_423J2_125_3477_n2262), 
        .A2(DP_OP_425J2_127_3477_n2578), .Y(DP_OP_425J2_127_3477_n2554) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2015 ( .A1(DP_OP_423J2_125_3477_n2044), 
        .A2(DP_OP_425J2_127_3477_n2798), .Y(DP_OP_425J2_127_3477_n2776) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1874 ( .A1(DP_OP_422J2_124_3477_n2791), 
        .A2(DP_OP_425J2_127_3477_n2665), .Y(DP_OP_425J2_127_3477_n2635) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1712 ( .A1(DP_OP_425J2_127_3477_n2481), 
        .A2(DP_OP_425J2_127_3477_n2491), .Y(DP_OP_425J2_127_3477_n2473) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2054 ( .A1(DP_OP_422J2_124_3477_n2091), 
        .A2(DP_OP_424J2_126_3477_n2841), .Y(DP_OP_423J2_125_3477_n2815) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1705 ( .A1(DP_OP_425J2_127_3477_n2482), 
        .A2(DP_OP_425J2_127_3477_n2490), .Y(DP_OP_425J2_127_3477_n2466) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1406 ( .A1(DP_OP_425J2_127_3477_n2175), 
        .A2(DP_OP_424J2_126_3477_n2183), .Y(DP_OP_425J2_127_3477_n2167) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1918 ( .A1(DP_OP_422J2_124_3477_n2835), 
        .A2(DP_OP_425J2_127_3477_n2709), .Y(DP_OP_425J2_127_3477_n2679) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1170 ( .A1(DP_OP_424J2_126_3477_n3009), 
        .A2(DP_OP_425J2_127_3477_n1961), .Y(DP_OP_425J2_127_3477_n1931) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1610 ( .A1(DP_OP_422J2_124_3477_n2263), 
        .A2(DP_OP_425J2_127_3477_n2401), .Y(DP_OP_425J2_127_3477_n2371) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1619 ( .A1(DP_OP_423J2_125_3477_n2396), 
        .A2(DP_OP_423J2_125_3477_n2402), .Y(DP_OP_423J2_125_3477_n2380) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2022 ( .A1(DP_OP_423J2_125_3477_n2791), 
        .A2(DP_OP_422J2_124_3477_n2799), .Y(DP_OP_423J2_125_3477_n2783) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1830 ( .A1(DP_OP_423J2_125_3477_n2219), 
        .A2(DP_OP_425J2_127_3477_n2621), .Y(DP_OP_425J2_127_3477_n2591) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1346 ( .A1(DP_OP_424J2_126_3477_n2835), 
        .A2(DP_OP_425J2_127_3477_n2137), .Y(DP_OP_425J2_127_3477_n2107) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1436 ( .A1(DP_OP_423J2_125_3477_n2837), 
        .A2(DP_OP_422J2_124_3477_n2225), .Y(DP_OP_425J2_127_3477_n2197) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1575 ( .A1(DP_OP_424J2_126_3477_n2616), 
        .A2(DP_OP_425J2_127_3477_n2358), .Y(DP_OP_425J2_127_3477_n2336) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1920 ( .A1(DP_OP_425J2_127_3477_n2705), 
        .A2(DP_OP_425J2_127_3477_n2709), .Y(DP_OP_425J2_127_3477_n2681) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2140 ( .A1(DP_OP_424J2_126_3477_n2001), 
        .A2(DP_OP_425J2_127_3477_n2929), .Y(DP_OP_425J2_127_3477_n2901) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1758 ( .A1(DP_OP_423J2_125_3477_n2307), 
        .A2(DP_OP_425J2_127_3477_n2535), .Y(DP_OP_425J2_127_3477_n2519) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1890 ( .A1(DP_OP_423J2_125_3477_n2175), 
        .A2(DP_OP_425J2_127_3477_n2667), .Y(DP_OP_425J2_127_3477_n2651) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1876 ( .A1(DP_OP_424J2_126_3477_n2265), 
        .A2(DP_OP_425J2_127_3477_n2665), .Y(DP_OP_425J2_127_3477_n2637) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1700 ( .A1(DP_OP_422J2_124_3477_n2617), 
        .A2(DP_OP_425J2_127_3477_n2489), .Y(DP_OP_425J2_127_3477_n2461) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1670 ( .A1(DP_OP_425J2_127_3477_n2439), 
        .A2(DP_OP_425J2_127_3477_n2447), .Y(DP_OP_425J2_127_3477_n2431) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1964 ( .A1(DP_OP_425J2_127_3477_n2749), 
        .A2(DP_OP_422J2_124_3477_n2753), .Y(DP_OP_425J2_127_3477_n2725) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1267 ( .A1(DP_OP_423J2_125_3477_n3010), 
        .A2(DP_OP_425J2_127_3477_n2050), .Y(DP_OP_425J2_127_3477_n2028) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1832 ( .A1(DP_OP_425J2_127_3477_n2617), 
        .A2(DP_OP_425J2_127_3477_n2621), .Y(DP_OP_425J2_127_3477_n2593) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1260 ( .A1(DP_OP_423J2_125_3477_n3011), 
        .A2(DP_OP_425J2_127_3477_n2049), .Y(DP_OP_425J2_127_3477_n2021) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2198 ( .A1(DP_OP_425J2_127_3477_n2967), 
        .A2(DP_OP_425J2_127_3477_n2975), .Y(DP_OP_425J2_127_3477_n2959) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1230 ( .A1(DP_OP_424J2_126_3477_n2967), 
        .A2(DP_OP_425J2_127_3477_n2007), .Y(DP_OP_425J2_127_3477_n1991) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2228 ( .A1(DP_OP_425J2_127_3477_n3011), 
        .A2(DP_OP_425J2_127_3477_n3015), .Y(DP_OP_425J2_127_3477_n2987) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1355 ( .A1(DP_OP_425J2_127_3477_n2704), 
        .A2(DP_OP_423J2_125_3477_n2138), .Y(DP_OP_423J2_125_3477_n2116) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1619 ( .A1(DP_OP_425J2_127_3477_n2396), 
        .A2(DP_OP_425J2_127_3477_n2402), .Y(DP_OP_425J2_127_3477_n2380) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1450 ( .A1(DP_OP_425J2_127_3477_n2219), 
        .A2(DP_OP_425J2_127_3477_n2227), .Y(DP_OP_425J2_127_3477_n2211) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1714 ( .A1(DP_OP_424J2_126_3477_n2439), 
        .A2(DP_OP_425J2_127_3477_n2491), .Y(DP_OP_425J2_127_3477_n2475) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1751 ( .A1(DP_OP_425J2_127_3477_n2528), 
        .A2(DP_OP_425J2_127_3477_n2534), .Y(DP_OP_425J2_127_3477_n2512) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1355 ( .A1(DP_OP_423J2_125_3477_n2924), 
        .A2(DP_OP_425J2_127_3477_n2138), .Y(DP_OP_425J2_127_3477_n2116) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2022 ( .A1(DP_OP_425J2_127_3477_n2791), 
        .A2(DP_OP_425J2_127_3477_n2799), .Y(DP_OP_425J2_127_3477_n2783) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1524 ( .A1(DP_OP_423J2_125_3477_n2749), 
        .A2(DP_OP_425J2_127_3477_n2313), .Y(DP_OP_425J2_127_3477_n2285) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1494 ( .A1(DP_OP_423J2_125_3477_n2791), 
        .A2(DP_OP_425J2_127_3477_n2271), .Y(DP_OP_425J2_127_3477_n2255) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1304 ( .A1(DP_OP_423J2_125_3477_n2969), 
        .A2(DP_OP_425J2_127_3477_n2093), .Y(DP_OP_425J2_127_3477_n2065) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1795 ( .A1(DP_OP_425J2_127_3477_n2572), 
        .A2(DP_OP_425J2_127_3477_n2578), .Y(DP_OP_425J2_127_3477_n2556) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1538 ( .A1(DP_OP_425J2_127_3477_n2307), 
        .A2(DP_OP_425J2_127_3477_n2315), .Y(DP_OP_425J2_127_3477_n2299) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2103 ( .A1(DP_OP_424J2_126_3477_n2044), 
        .A2(DP_OP_424J2_126_3477_n2886), .Y(DP_OP_425J2_127_3477_n2864) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2110 ( .A1(DP_OP_425J2_127_3477_n2879), 
        .A2(DP_OP_425J2_127_3477_n2887), .Y(DP_OP_425J2_127_3477_n2871) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1568 ( .A1(DP_OP_425J2_127_3477_n2353), 
        .A2(DP_OP_425J2_127_3477_n2357), .Y(DP_OP_425J2_127_3477_n2329) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1392 ( .A1(DP_OP_424J2_126_3477_n2793), 
        .A2(DP_OP_425J2_127_3477_n2181), .Y(DP_OP_425J2_127_3477_n2153) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1487 ( .A1(DP_OP_425J2_127_3477_n2264), 
        .A2(DP_OP_425J2_127_3477_n2270), .Y(DP_OP_425J2_127_3477_n2248) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1480 ( .A1(DP_OP_423J2_125_3477_n2793), 
        .A2(DP_OP_425J2_127_3477_n2269), .Y(DP_OP_425J2_127_3477_n2241) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1172 ( .A1(DP_OP_424J2_126_3477_n3011), 
        .A2(DP_OP_425J2_127_3477_n1961), .Y(DP_OP_425J2_127_3477_n1933) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1179 ( .A1(DP_OP_424J2_126_3477_n3010), 
        .A2(DP_OP_422J2_124_3477_n1962), .Y(DP_OP_425J2_127_3477_n1940) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1744 ( .A1(DP_OP_425J2_127_3477_n2529), 
        .A2(DP_OP_422J2_124_3477_n2533), .Y(DP_OP_425J2_127_3477_n2505) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1883 ( .A1(DP_OP_422J2_124_3477_n2792), 
        .A2(DP_OP_425J2_127_3477_n2666), .Y(DP_OP_425J2_127_3477_n2644) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1846 ( .A1(DP_OP_422J2_124_3477_n2747), 
        .A2(DP_OP_425J2_127_3477_n2623), .Y(DP_OP_425J2_127_3477_n2607) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1399 ( .A1(DP_OP_423J2_125_3477_n2880), 
        .A2(DP_OP_425J2_127_3477_n2182), .Y(DP_OP_425J2_127_3477_n2160) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1450 ( .A1(DP_OP_423J2_125_3477_n2219), 
        .A2(DP_OP_425J2_127_3477_n2227), .Y(DP_OP_423J2_125_3477_n2211) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1223 ( .A1(DP_OP_425J2_127_3477_n2000), 
        .A2(DP_OP_425J2_127_3477_n2006), .Y(DP_OP_425J2_127_3477_n1984) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2235 ( .A1(DP_OP_425J2_127_3477_n3010), 
        .A2(DP_OP_422J2_124_3477_n3016), .Y(DP_OP_425J2_127_3477_n2994) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1626 ( .A1(DP_OP_422J2_124_3477_n2263), 
        .A2(DP_OP_425J2_127_3477_n2403), .Y(DP_OP_425J2_127_3477_n2387) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1216 ( .A1(DP_OP_424J2_126_3477_n2969), 
        .A2(DP_OP_425J2_127_3477_n2005), .Y(DP_OP_425J2_127_3477_n1977) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1261 ( .A1(DP_OP_425J2_127_3477_n2794), 
        .A2(DP_OP_422J2_124_3477_n2049), .Y(DP_OP_423J2_125_3477_n2022) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2052 ( .A1(DP_OP_425J2_127_3477_n2837), 
        .A2(DP_OP_424J2_126_3477_n2841), .Y(DP_OP_425J2_127_3477_n2813) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2059 ( .A1(DP_OP_423J2_125_3477_n2000), 
        .A2(DP_OP_425J2_127_3477_n2842), .Y(DP_OP_425J2_127_3477_n2820) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2145 ( .A1(DP_OP_425J2_127_3477_n2922), 
        .A2(DP_OP_425J2_127_3477_n2930), .Y(DP_OP_425J2_127_3477_n2906) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1230 ( .A1(DP_OP_425J2_127_3477_n2835), 
        .A2(DP_OP_423J2_125_3477_n2007), .Y(DP_OP_423J2_125_3477_n1991) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1177 ( .A1(DP_OP_424J2_126_3477_n3008), 
        .A2(DP_OP_422J2_124_3477_n1962), .Y(DP_OP_425J2_127_3477_n1938) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2105 ( .A1(DP_OP_424J2_126_3477_n2794), 
        .A2(DP_OP_423J2_125_3477_n2886), .Y(DP_OP_423J2_125_3477_n2866) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1224 ( .A1(DP_OP_422J2_124_3477_n2969), 
        .A2(DP_OP_423J2_125_3477_n2006), .Y(DP_OP_423J2_125_3477_n1985) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1663 ( .A1(DP_OP_424J2_126_3477_n2528), 
        .A2(DP_OP_425J2_127_3477_n2446), .Y(DP_OP_425J2_127_3477_n2424) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2152 ( .A1(DP_OP_425J2_127_3477_n2921), 
        .A2(DP_OP_425J2_127_3477_n2931), .Y(DP_OP_425J2_127_3477_n2913) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2182 ( .A1(DP_OP_425J2_127_3477_n2967), 
        .A2(DP_OP_425J2_127_3477_n2973), .Y(DP_OP_425J2_127_3477_n2943) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1231 ( .A1(DP_OP_423J2_125_3477_n2000), 
        .A2(DP_OP_423J2_125_3477_n2007), .Y(DP_OP_423J2_125_3477_n1992) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2066 ( .A1(DP_OP_425J2_127_3477_n2835), 
        .A2(DP_OP_425J2_127_3477_n2843), .Y(DP_OP_425J2_127_3477_n2827) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1494 ( .A1(DP_OP_423J2_125_3477_n2263), 
        .A2(DP_OP_424J2_126_3477_n2271), .Y(DP_OP_423J2_125_3477_n2255) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1397 ( .A1(DP_OP_423J2_125_3477_n2878), 
        .A2(DP_OP_425J2_127_3477_n2182), .Y(DP_OP_425J2_127_3477_n2158) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1390 ( .A1(DP_OP_425J2_127_3477_n2175), 
        .A2(DP_OP_425J2_127_3477_n2181), .Y(DP_OP_425J2_127_3477_n2151) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1173 ( .A1(DP_OP_423J2_125_3477_n1958), 
        .A2(DP_OP_425J2_127_3477_n1961), .Y(DP_OP_423J2_125_3477_n1934) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1265 ( .A1(DP_OP_423J2_125_3477_n3008), 
        .A2(DP_OP_425J2_127_3477_n2050), .Y(DP_OP_425J2_127_3477_n2026) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1258 ( .A1(DP_OP_423J2_125_3477_n3009), 
        .A2(DP_OP_425J2_127_3477_n2049), .Y(DP_OP_425J2_127_3477_n2019) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1661 ( .A1(DP_OP_425J2_127_3477_n2438), 
        .A2(DP_OP_425J2_127_3477_n2446), .Y(DP_OP_425J2_127_3477_n2422) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2142 ( .A1(DP_OP_423J2_125_3477_n2927), 
        .A2(DP_OP_423J2_125_3477_n2929), .Y(DP_OP_423J2_125_3477_n2903) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1654 ( .A1(DP_OP_425J2_127_3477_n2439), 
        .A2(DP_OP_425J2_127_3477_n2445), .Y(DP_OP_425J2_127_3477_n2415) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1348 ( .A1(DP_OP_425J2_127_3477_n2133), 
        .A2(DP_OP_425J2_127_3477_n2137), .Y(DP_OP_425J2_127_3477_n2109) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1180 ( .A1(DP_OP_423J2_125_3477_n1957), 
        .A2(DP_OP_423J2_125_3477_n1962), .Y(DP_OP_423J2_125_3477_n1941) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1612 ( .A1(DP_OP_425J2_127_3477_n2397), 
        .A2(DP_OP_425J2_127_3477_n2401), .Y(DP_OP_425J2_127_3477_n2373) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2189 ( .A1(DP_OP_424J2_126_3477_n1954), 
        .A2(DP_OP_425J2_127_3477_n2974), .Y(DP_OP_425J2_127_3477_n2950) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1573 ( .A1(DP_OP_423J2_125_3477_n2702), 
        .A2(DP_OP_425J2_127_3477_n2358), .Y(DP_OP_425J2_127_3477_n2334) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1217 ( .A1(DP_OP_422J2_124_3477_n2970), 
        .A2(DP_OP_423J2_125_3477_n2005), .Y(DP_OP_423J2_125_3477_n1978) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1934 ( .A1(DP_OP_422J2_124_3477_n2835), 
        .A2(DP_OP_425J2_127_3477_n2711), .Y(DP_OP_425J2_127_3477_n2695) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2226 ( .A1(DP_OP_425J2_127_3477_n3009), 
        .A2(DP_OP_425J2_127_3477_n3015), .Y(DP_OP_425J2_127_3477_n2985) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2233 ( .A1(DP_OP_425J2_127_3477_n3008), 
        .A2(DP_OP_422J2_124_3477_n3016), .Y(DP_OP_425J2_127_3477_n2992) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1707 ( .A1(DP_OP_425J2_127_3477_n2484), 
        .A2(DP_OP_425J2_127_3477_n2490), .Y(DP_OP_425J2_127_3477_n2468) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1617 ( .A1(DP_OP_422J2_124_3477_n2262), 
        .A2(DP_OP_425J2_127_3477_n2402), .Y(DP_OP_425J2_127_3477_n2378) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1927 ( .A1(DP_OP_425J2_127_3477_n2704), 
        .A2(DP_OP_425J2_127_3477_n2710), .Y(DP_OP_425J2_127_3477_n2688) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1353 ( .A1(DP_OP_423J2_125_3477_n2922), 
        .A2(DP_OP_425J2_127_3477_n2138), .Y(DP_OP_425J2_127_3477_n2114) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1797 ( .A1(DP_OP_423J2_125_3477_n2574), 
        .A2(DP_OP_422J2_124_3477_n2578), .Y(DP_OP_423J2_125_3477_n2558) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1488 ( .A1(DP_OP_423J2_125_3477_n2265), 
        .A2(DP_OP_423J2_125_3477_n2270), .Y(DP_OP_423J2_125_3477_n2249) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2013 ( .A1(DP_OP_425J2_127_3477_n2790), 
        .A2(DP_OP_425J2_127_3477_n2798), .Y(DP_OP_425J2_127_3477_n2774) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1656 ( .A1(DP_OP_425J2_127_3477_n2441), 
        .A2(DP_OP_425J2_127_3477_n2445), .Y(DP_OP_425J2_127_3477_n2417) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1214 ( .A1(DP_OP_424J2_126_3477_n2967), 
        .A2(DP_OP_425J2_127_3477_n2005), .Y(DP_OP_425J2_127_3477_n1975) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2057 ( .A1(DP_OP_425J2_127_3477_n2834), 
        .A2(DP_OP_425J2_127_3477_n2842), .Y(DP_OP_425J2_127_3477_n2818) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2155 ( .A1(DP_OP_423J2_125_3477_n2924), 
        .A2(DP_OP_423J2_125_3477_n2931), .Y(DP_OP_423J2_125_3477_n2916) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1452 ( .A1(DP_OP_422J2_124_3477_n2749), 
        .A2(DP_OP_425J2_127_3477_n2227), .Y(DP_OP_423J2_125_3477_n2213) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1478 ( .A1(DP_OP_423J2_125_3477_n2791), 
        .A2(DP_OP_425J2_127_3477_n2269), .Y(DP_OP_425J2_127_3477_n2239) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2191 ( .A1(DP_OP_424J2_126_3477_n1956), 
        .A2(DP_OP_425J2_127_3477_n2974), .Y(DP_OP_425J2_127_3477_n2952) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1522 ( .A1(DP_OP_425J2_127_3477_n2307), 
        .A2(DP_OP_425J2_127_3477_n2313), .Y(DP_OP_425J2_127_3477_n2283) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2064 ( .A1(DP_OP_425J2_127_3477_n2833), 
        .A2(DP_OP_425J2_127_3477_n2843), .Y(DP_OP_425J2_127_3477_n2825) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2184 ( .A1(DP_OP_424J2_126_3477_n1957), 
        .A2(DP_OP_425J2_127_3477_n2973), .Y(DP_OP_425J2_127_3477_n2945) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1582 ( .A1(DP_OP_425J2_127_3477_n2351), 
        .A2(DP_OP_425J2_127_3477_n2359), .Y(DP_OP_425J2_127_3477_n2343) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1221 ( .A1(DP_OP_425J2_127_3477_n1998), 
        .A2(DP_OP_425J2_127_3477_n2006), .Y(DP_OP_425J2_127_3477_n1982) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1485 ( .A1(DP_OP_423J2_125_3477_n2790), 
        .A2(DP_OP_425J2_127_3477_n2270), .Y(DP_OP_425J2_127_3477_n2246) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1749 ( .A1(DP_OP_425J2_127_3477_n2526), 
        .A2(DP_OP_425J2_127_3477_n2534), .Y(DP_OP_425J2_127_3477_n2510) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1742 ( .A1(DP_OP_422J2_124_3477_n2659), 
        .A2(DP_OP_422J2_124_3477_n2533), .Y(DP_OP_425J2_127_3477_n2503) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1962 ( .A1(DP_OP_425J2_127_3477_n2747), 
        .A2(DP_OP_422J2_124_3477_n2753), .Y(DP_OP_425J2_127_3477_n2723) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1489 ( .A1(DP_OP_423J2_125_3477_n2266), 
        .A2(DP_OP_423J2_125_3477_n2270), .Y(DP_OP_423J2_125_3477_n2250) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1566 ( .A1(DP_OP_425J2_127_3477_n2351), 
        .A2(DP_OP_425J2_127_3477_n2357), .Y(DP_OP_425J2_127_3477_n2327) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1482 ( .A1(DP_OP_423J2_125_3477_n2267), 
        .A2(DP_OP_424J2_126_3477_n2269), .Y(DP_OP_423J2_125_3477_n2243) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2101 ( .A1(DP_OP_425J2_127_3477_n2878), 
        .A2(DP_OP_424J2_126_3477_n2886), .Y(DP_OP_425J2_127_3477_n2862) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1580 ( .A1(DP_OP_424J2_126_3477_n2613), 
        .A2(DP_OP_425J2_127_3477_n2359), .Y(DP_OP_425J2_127_3477_n2341) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2061 ( .A1(DP_OP_424J2_126_3477_n2750), 
        .A2(DP_OP_423J2_125_3477_n2842), .Y(DP_OP_423J2_125_3477_n2822) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1404 ( .A1(DP_OP_424J2_126_3477_n2789), 
        .A2(DP_OP_424J2_126_3477_n2183), .Y(DP_OP_425J2_127_3477_n2165) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2138 ( .A1(DP_OP_425J2_127_3477_n2923), 
        .A2(DP_OP_425J2_127_3477_n2929), .Y(DP_OP_425J2_127_3477_n2899) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1496 ( .A1(DP_OP_423J2_125_3477_n2265), 
        .A2(DP_OP_424J2_126_3477_n2271), .Y(DP_OP_423J2_125_3477_n2257) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2228 ( .A1(DP_OP_423J2_125_3477_n3011), 
        .A2(DP_OP_425J2_127_3477_n3015), .Y(DP_OP_423J2_125_3477_n2987) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2154 ( .A1(DP_OP_425J2_127_3477_n2923), 
        .A2(DP_OP_425J2_127_3477_n2931), .Y(DP_OP_425J2_127_3477_n2915) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1624 ( .A1(DP_OP_422J2_124_3477_n2261), 
        .A2(DP_OP_425J2_127_3477_n2403), .Y(DP_OP_425J2_127_3477_n2385) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1698 ( .A1(DP_OP_424J2_126_3477_n2439), 
        .A2(DP_OP_425J2_127_3477_n2489), .Y(DP_OP_425J2_127_3477_n2459) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2147 ( .A1(DP_OP_425J2_127_3477_n2924), 
        .A2(DP_OP_425J2_127_3477_n2930), .Y(DP_OP_425J2_127_3477_n2908) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1881 ( .A1(DP_OP_425J2_127_3477_n2658), 
        .A2(DP_OP_425J2_127_3477_n2666), .Y(DP_OP_425J2_127_3477_n2642) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1434 ( .A1(DP_OP_425J2_127_3477_n2219), 
        .A2(DP_OP_424J2_126_3477_n2225), .Y(DP_OP_425J2_127_3477_n2195) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2242 ( .A1(DP_OP_425J2_127_3477_n3009), 
        .A2(DP_OP_425J2_127_3477_n3017), .Y(DP_OP_425J2_127_3477_n3001) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1526 ( .A1(DP_OP_423J2_125_3477_n2311), 
        .A2(DP_OP_423J2_125_3477_n2313), .Y(DP_OP_423J2_125_3477_n2287) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1524 ( .A1(DP_OP_424J2_126_3477_n2397), 
        .A2(DP_OP_423J2_125_3477_n2313), .Y(DP_OP_423J2_125_3477_n2285) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1756 ( .A1(DP_OP_425J2_127_3477_n2525), 
        .A2(DP_OP_425J2_127_3477_n2535), .Y(DP_OP_425J2_127_3477_n2517) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U115 ( .A1(DP_OP_425J2_127_3477_n115), .A2(
        DP_OP_425J2_127_3477_n118), .Y(DP_OP_425J2_127_3477_n113) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U115 ( .A1(DP_OP_424J2_126_3477_n115), .A2(
        DP_OP_424J2_126_3477_n118), .Y(DP_OP_424J2_126_3477_n113) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U115 ( .A1(DP_OP_423J2_125_3477_n115), .A2(
        DP_OP_423J2_125_3477_n118), .Y(DP_OP_423J2_125_3477_n113) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U115 ( .A1(DP_OP_422J2_124_3477_n115), .A2(
        DP_OP_422J2_124_3477_n118), .Y(DP_OP_422J2_124_3477_n113) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U95 ( .A1(DP_OP_425J2_127_3477_n101), .A2(
        DP_OP_425J2_127_3477_n104), .Y(DP_OP_425J2_127_3477_n99) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U95 ( .A1(DP_OP_423J2_125_3477_n101), .A2(
        DP_OP_423J2_125_3477_n104), .Y(DP_OP_423J2_125_3477_n99) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U75 ( .A1(DP_OP_423J2_125_3477_n87), .A2(
        DP_OP_423J2_125_3477_n90), .Y(DP_OP_423J2_125_3477_n85) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U75 ( .A1(DP_OP_425J2_127_3477_n87), .A2(
        DP_OP_425J2_127_3477_n90), .Y(DP_OP_425J2_127_3477_n85) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U247 ( .A1(DP_OP_422J2_124_3477_n203), .A2(
        DP_OP_422J2_124_3477_n201), .A3(DP_OP_422J2_124_3477_n202), .Y(
        DP_OP_422J2_124_3477_n200) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U47 ( .A1(DP_OP_425J2_127_3477_n65), .A2(
        DP_OP_425J2_127_3477_n148), .Y(DP_OP_425J2_127_3477_n63) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U47 ( .A1(DP_OP_423J2_125_3477_n65), .A2(
        DP_OP_423J2_125_3477_n148), .Y(DP_OP_423J2_125_3477_n63) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U247 ( .A1(DP_OP_423J2_125_3477_n203), .A2(
        DP_OP_423J2_125_3477_n201), .A3(DP_OP_423J2_125_3477_n202), .Y(
        DP_OP_423J2_125_3477_n200) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U47 ( .A1(DP_OP_422J2_124_3477_n65), .A2(
        DP_OP_422J2_124_3477_n148), .Y(DP_OP_422J2_124_3477_n63) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U247 ( .A1(DP_OP_425J2_127_3477_n203), .A2(
        DP_OP_425J2_127_3477_n201), .A3(DP_OP_425J2_127_3477_n202), .Y(
        DP_OP_425J2_127_3477_n200) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U247 ( .A1(DP_OP_424J2_126_3477_n203), .A2(
        DP_OP_424J2_126_3477_n201), .A3(DP_OP_424J2_126_3477_n202), .Y(
        DP_OP_424J2_126_3477_n200) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U47 ( .A1(DP_OP_424J2_126_3477_n65), .A2(
        DP_OP_424J2_126_3477_n148), .Y(DP_OP_424J2_126_3477_n63) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U220 ( .A1(DP_OP_423J2_125_3477_n190), .A2(
        DP_OP_423J2_125_3477_n186), .A3(DP_OP_423J2_125_3477_n187), .Y(
        DP_OP_423J2_125_3477_n185) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U233 ( .A1(DP_OP_424J2_126_3477_n193), .A2(
        DP_OP_424J2_126_3477_n195), .A3(DP_OP_424J2_126_3477_n194), .Y(
        DP_OP_424J2_126_3477_n192) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U220 ( .A1(DP_OP_425J2_127_3477_n190), .A2(
        DP_OP_425J2_127_3477_n186), .A3(DP_OP_425J2_127_3477_n187), .Y(
        DP_OP_425J2_127_3477_n185) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U189 ( .A1(DP_OP_422J2_124_3477_n167), .A2(
        DP_OP_422J2_124_3477_n171), .A3(DP_OP_422J2_124_3477_n168), .Y(
        DP_OP_422J2_124_3477_n166) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U189 ( .A1(DP_OP_423J2_125_3477_n167), .A2(
        DP_OP_423J2_125_3477_n171), .A3(DP_OP_423J2_125_3477_n168), .Y(
        DP_OP_423J2_125_3477_n166) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U220 ( .A1(DP_OP_424J2_126_3477_n190), .A2(
        DP_OP_424J2_126_3477_n186), .A3(DP_OP_424J2_126_3477_n187), .Y(
        DP_OP_424J2_126_3477_n185) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U233 ( .A1(DP_OP_425J2_127_3477_n193), .A2(
        DP_OP_425J2_127_3477_n195), .A3(DP_OP_425J2_127_3477_n194), .Y(
        DP_OP_425J2_127_3477_n192) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U220 ( .A1(DP_OP_422J2_124_3477_n190), .A2(
        DP_OP_422J2_124_3477_n186), .A3(DP_OP_422J2_124_3477_n187), .Y(
        DP_OP_422J2_124_3477_n185) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U189 ( .A1(DP_OP_425J2_127_3477_n167), .A2(
        DP_OP_425J2_127_3477_n171), .A3(DP_OP_425J2_127_3477_n168), .Y(
        DP_OP_425J2_127_3477_n166) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U189 ( .A1(DP_OP_424J2_126_3477_n167), .A2(
        DP_OP_424J2_126_3477_n171), .A3(DP_OP_424J2_126_3477_n168), .Y(
        DP_OP_424J2_126_3477_n166) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U233 ( .A1(DP_OP_423J2_125_3477_n193), .A2(
        DP_OP_423J2_125_3477_n195), .A3(DP_OP_423J2_125_3477_n194), .Y(
        DP_OP_423J2_125_3477_n192) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U233 ( .A1(DP_OP_422J2_124_3477_n193), .A2(
        DP_OP_422J2_124_3477_n195), .A3(DP_OP_422J2_124_3477_n194), .Y(
        DP_OP_422J2_124_3477_n192) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U150 ( .A1(DP_OP_425J2_127_3477_n137), .A2(
        DP_OP_425J2_127_3477_n145), .A3(DP_OP_425J2_127_3477_n140), .Y(
        DP_OP_425J2_127_3477_n136) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U38 ( .A1(DP_OP_422J2_124_3477_n58), .A2(
        DP_OP_422J2_124_3477_n62), .A3(DP_OP_422J2_124_3477_n59), .Y(
        DP_OP_422J2_124_3477_n57) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U150 ( .A1(DP_OP_422J2_124_3477_n137), .A2(
        DP_OP_422J2_124_3477_n145), .A3(DP_OP_422J2_124_3477_n140), .Y(
        DP_OP_422J2_124_3477_n136) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U37 ( .A1(DP_OP_422J2_124_3477_n58), .A2(
        DP_OP_422J2_124_3477_n61), .Y(DP_OP_422J2_124_3477_n56) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U150 ( .A1(DP_OP_424J2_126_3477_n137), .A2(
        DP_OP_424J2_126_3477_n145), .A3(DP_OP_424J2_126_3477_n140), .Y(
        DP_OP_424J2_126_3477_n136) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U37 ( .A1(DP_OP_423J2_125_3477_n58), .A2(
        DP_OP_423J2_125_3477_n61), .Y(DP_OP_423J2_125_3477_n56) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U150 ( .A1(DP_OP_423J2_125_3477_n137), .A2(
        DP_OP_423J2_125_3477_n145), .A3(DP_OP_423J2_125_3477_n140), .Y(
        DP_OP_423J2_125_3477_n136) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U37 ( .A1(DP_OP_424J2_126_3477_n58), .A2(
        DP_OP_424J2_126_3477_n61), .Y(DP_OP_424J2_126_3477_n56) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U38 ( .A1(DP_OP_423J2_125_3477_n58), .A2(
        DP_OP_423J2_125_3477_n62), .A3(DP_OP_423J2_125_3477_n59), .Y(
        DP_OP_423J2_125_3477_n57) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U38 ( .A1(DP_OP_424J2_126_3477_n58), .A2(
        DP_OP_424J2_126_3477_n62), .A3(DP_OP_424J2_126_3477_n59), .Y(
        DP_OP_424J2_126_3477_n57) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U38 ( .A1(DP_OP_425J2_127_3477_n58), .A2(
        DP_OP_425J2_127_3477_n62), .A3(DP_OP_425J2_127_3477_n59), .Y(
        DP_OP_425J2_127_3477_n57) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U37 ( .A1(DP_OP_425J2_127_3477_n58), .A2(
        DP_OP_425J2_127_3477_n61), .Y(DP_OP_425J2_127_3477_n56) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U17 ( .A1(DP_OP_422J2_124_3477_n44), .A2(
        DP_OP_422J2_124_3477_n47), .Y(DP_OP_422J2_124_3477_n42) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U18 ( .A1(DP_OP_423J2_125_3477_n44), .A2(
        DP_OP_423J2_125_3477_n48), .A3(DP_OP_423J2_125_3477_n45), .Y(
        DP_OP_423J2_125_3477_n43) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U18 ( .A1(DP_OP_425J2_127_3477_n44), .A2(
        DP_OP_425J2_127_3477_n48), .A3(DP_OP_425J2_127_3477_n45), .Y(
        DP_OP_425J2_127_3477_n43) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U18 ( .A1(DP_OP_422J2_124_3477_n44), .A2(
        DP_OP_422J2_124_3477_n48), .A3(DP_OP_422J2_124_3477_n45), .Y(
        DP_OP_422J2_124_3477_n43) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U17 ( .A1(DP_OP_423J2_125_3477_n44), .A2(
        DP_OP_423J2_125_3477_n47), .Y(DP_OP_423J2_125_3477_n42) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U17 ( .A1(DP_OP_425J2_127_3477_n44), .A2(
        DP_OP_425J2_127_3477_n47), .Y(DP_OP_425J2_127_3477_n42) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U17 ( .A1(DP_OP_424J2_126_3477_n44), .A2(
        DP_OP_424J2_126_3477_n47), .Y(DP_OP_424J2_126_3477_n42) );
  XNOR2X1_HVT DP_OP_424J2_126_3477_U208 ( .A1(DP_OP_424J2_126_3477_n182), .A2(
        DP_OP_424J2_126_3477_n26), .Y(n_conv2_sum_c[10]) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U18 ( .A1(DP_OP_424J2_126_3477_n44), .A2(
        DP_OP_424J2_126_3477_n48), .A3(DP_OP_424J2_126_3477_n45), .Y(
        DP_OP_424J2_126_3477_n43) );
  XOR2X1_HVT DP_OP_423J2_125_3477_U200 ( .A1(DP_OP_423J2_125_3477_n177), .A2(
        DP_OP_423J2_125_3477_n25), .Y(n_conv2_sum_b[11]) );
  XOR2X1_HVT DP_OP_423J2_125_3477_U147 ( .A1(DP_OP_423J2_125_3477_n141), .A2(
        DP_OP_423J2_125_3477_n20), .Y(n_conv2_sum_b[16]) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U170 ( .A1(DP_OP_422J2_124_3477_n151), .A2(
        DP_OP_422J2_124_3477_n161), .A3(DP_OP_422J2_124_3477_n152), .Y(
        DP_OP_422J2_124_3477_n150) );
  XOR2X1_HVT DP_OP_422J2_124_3477_U169 ( .A1(DP_OP_422J2_124_3477_n161), .A2(
        DP_OP_422J2_124_3477_n22), .Y(n_conv2_sum_a[14]) );
  XOR2X1_HVT DP_OP_425J2_127_3477_U147 ( .A1(DP_OP_425J2_127_3477_n141), .A2(
        DP_OP_425J2_127_3477_n20), .Y(n_conv2_sum_d[16]) );
  XOR2X1_HVT DP_OP_424J2_126_3477_U200 ( .A1(DP_OP_424J2_126_3477_n177), .A2(
        DP_OP_424J2_126_3477_n25), .Y(n_conv2_sum_c[11]) );
  XOR2X1_HVT DP_OP_422J2_124_3477_U200 ( .A1(DP_OP_422J2_124_3477_n177), .A2(
        DP_OP_422J2_124_3477_n25), .Y(n_conv2_sum_a[11]) );
  XOR2X1_HVT DP_OP_424J2_126_3477_U169 ( .A1(DP_OP_424J2_126_3477_n161), .A2(
        DP_OP_424J2_126_3477_n22), .Y(n_conv2_sum_c[14]) );
  XOR2X1_HVT DP_OP_425J2_127_3477_U200 ( .A1(DP_OP_425J2_127_3477_n177), .A2(
        DP_OP_425J2_127_3477_n25), .Y(n_conv2_sum_d[11]) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U170 ( .A1(DP_OP_424J2_126_3477_n151), .A2(
        DP_OP_424J2_126_3477_n161), .A3(DP_OP_424J2_126_3477_n152), .Y(
        DP_OP_424J2_126_3477_n150) );
  XNOR2X1_HVT DP_OP_422J2_124_3477_U157 ( .A1(DP_OP_422J2_124_3477_n150), .A2(
        DP_OP_422J2_124_3477_n21), .Y(n_conv2_sum_a[15]) );
  XNOR2X1_HVT DP_OP_424J2_126_3477_U157 ( .A1(DP_OP_424J2_126_3477_n150), .A2(
        DP_OP_424J2_126_3477_n21), .Y(n_conv2_sum_c[15]) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1528 ( .A1(DP_OP_425J2_127_3477_n2305), 
        .A2(DP_OP_425J2_127_3477_n2314), .Y(DP_OP_425J2_127_3477_n2289) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1968 ( .A1(DP_OP_423J2_125_3477_n2745), 
        .A2(DP_OP_423J2_125_3477_n2754), .Y(DP_OP_423J2_125_3477_n2729) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1968 ( .A1(DP_OP_425J2_127_3477_n2745), 
        .A2(DP_OP_425J2_127_3477_n2754), .Y(DP_OP_425J2_127_3477_n2729) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1529 ( .A1(DP_OP_423J2_125_3477_n2746), 
        .A2(DP_OP_425J2_127_3477_n2314), .Y(DP_OP_425J2_127_3477_n2290) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1528 ( .A1(DP_OP_422J2_124_3477_n2745), 
        .A2(DP_OP_424J2_126_3477_n2314), .Y(DP_OP_424J2_126_3477_n2289) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1440 ( .A1(DP_OP_424J2_126_3477_n2217), 
        .A2(DP_OP_424J2_126_3477_n2226), .Y(DP_OP_424J2_126_3477_n2201) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1115 ( .A1(n334), .A2(n389), .Y(
        DP_OP_425J2_127_3477_n460) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1107 ( .A1(n485), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_424J2_126_3477_n276) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1113 ( .A1(n5001), .A2(n389), .Y(
        DP_OP_424J2_126_3477_n1875) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1113 ( .A1(n365), .A2(n390), .Y(
        DP_OP_425J2_127_3477_n1875) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1115 ( .A1(n486), .A2(
        DP_OP_425J2_127_3477_n2), .Y(DP_OP_424J2_126_3477_n460) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1099 ( .A1(n371), .A2(n386), .Y(
        DP_OP_423J2_125_3477_n260) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1102 ( .A1(n517), .A2(n386), .Y(
        DP_OP_424J2_126_3477_n266) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1113 ( .A1(n495), .A2(
        DP_OP_423J2_125_3477_n2), .Y(DP_OP_422J2_124_3477_n1875) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1114 ( .A1(n539), .A2(n390), .Y(
        DP_OP_422J2_124_3477_n1876) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1564 ( .A1(DP_OP_424J2_126_3477_n2613), 
        .A2(DP_OP_425J2_127_3477_n2357), .Y(DP_OP_425J2_127_3477_n2325) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1168 ( .A1(DP_OP_425J2_127_3477_n2965), 
        .A2(DP_OP_424J2_126_3477_n1961), .Y(DP_OP_424J2_126_3477_n1929) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1364 ( .A1(DP_OP_425J2_127_3477_n2705), 
        .A2(DP_OP_423J2_125_3477_n2139), .Y(DP_OP_423J2_125_3477_n2125) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1363 ( .A1(DP_OP_422J2_124_3477_n2924), 
        .A2(DP_OP_422J2_124_3477_n2139), .Y(DP_OP_424J2_126_3477_n2124) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2136 ( .A1(DP_OP_425J2_127_3477_n2921), 
        .A2(DP_OP_425J2_127_3477_n2929), .Y(DP_OP_425J2_127_3477_n2897) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1388 ( .A1(DP_OP_423J2_125_3477_n2877), 
        .A2(DP_OP_425J2_127_3477_n2181), .Y(DP_OP_425J2_127_3477_n2149) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2180 ( .A1(DP_OP_425J2_127_3477_n2965), 
        .A2(DP_OP_425J2_127_3477_n2973), .Y(DP_OP_425J2_127_3477_n2941) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1300 ( .A1(DP_OP_425J2_127_3477_n2085), 
        .A2(DP_OP_425J2_127_3477_n2093), .Y(DP_OP_425J2_127_3477_n2061) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1264 ( .A1(DP_OP_425J2_127_3477_n2789), 
        .A2(DP_OP_423J2_125_3477_n2050), .Y(DP_OP_423J2_125_3477_n2025) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1608 ( .A1(DP_OP_425J2_127_3477_n2525), 
        .A2(DP_OP_424J2_126_3477_n2401), .Y(DP_OP_424J2_126_3477_n2369) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1396 ( .A1(DP_OP_422J2_124_3477_n2789), 
        .A2(DP_OP_422J2_124_3477_n2182), .Y(DP_OP_423J2_125_3477_n2157) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1362 ( .A1(DP_OP_422J2_124_3477_n2923), 
        .A2(DP_OP_422J2_124_3477_n2139), .Y(DP_OP_424J2_126_3477_n2123) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1790 ( .A1(DP_OP_422J2_124_3477_n2575), 
        .A2(DP_OP_422J2_124_3477_n2577), .Y(DP_OP_422J2_124_3477_n2551) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1366 ( .A1(DP_OP_422J2_124_3477_n2135), 
        .A2(DP_OP_422J2_124_3477_n2139), .Y(DP_OP_422J2_124_3477_n2127) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1365 ( .A1(DP_OP_422J2_124_3477_n2926), 
        .A2(DP_OP_425J2_127_3477_n2139), .Y(DP_OP_424J2_126_3477_n2126) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2096 ( .A1(DP_OP_423J2_125_3477_n2969), 
        .A2(DP_OP_424J2_126_3477_n2885), .Y(DP_OP_424J2_126_3477_n2857) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2093 ( .A1(DP_OP_423J2_125_3477_n2878), 
        .A2(DP_OP_423J2_125_3477_n2885), .Y(DP_OP_423J2_125_3477_n2854) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1696 ( .A1(DP_OP_425J2_127_3477_n2481), 
        .A2(DP_OP_425J2_127_3477_n2489), .Y(DP_OP_425J2_127_3477_n2457) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1652 ( .A1(DP_OP_423J2_125_3477_n2613), 
        .A2(DP_OP_425J2_127_3477_n2445), .Y(DP_OP_425J2_127_3477_n2413) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1784 ( .A1(DP_OP_423J2_125_3477_n2261), 
        .A2(DP_OP_425J2_127_3477_n2577), .Y(DP_OP_425J2_127_3477_n2545) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1362 ( .A1(DP_OP_424J2_126_3477_n2703), 
        .A2(DP_OP_422J2_124_3477_n2139), .Y(DP_OP_422J2_124_3477_n2123) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1652 ( .A1(DP_OP_422J2_124_3477_n2613), 
        .A2(DP_OP_424J2_126_3477_n2445), .Y(DP_OP_424J2_126_3477_n2413) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1363 ( .A1(DP_OP_425J2_127_3477_n2704), 
        .A2(DP_OP_423J2_125_3477_n2139), .Y(DP_OP_423J2_125_3477_n2124) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2096 ( .A1(DP_OP_424J2_126_3477_n2177), 
        .A2(DP_OP_422J2_124_3477_n2885), .Y(DP_OP_422J2_124_3477_n2857) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1788 ( .A1(DP_OP_423J2_125_3477_n2397), 
        .A2(DP_OP_422J2_124_3477_n2577), .Y(DP_OP_422J2_124_3477_n2549) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2020 ( .A1(DP_OP_424J2_126_3477_n2789), 
        .A2(DP_OP_424J2_126_3477_n2799), .Y(DP_OP_424J2_126_3477_n2781) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1256 ( .A1(DP_OP_423J2_125_3477_n3007), 
        .A2(DP_OP_425J2_127_3477_n2049), .Y(DP_OP_425J2_127_3477_n2017) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2097 ( .A1(DP_OP_422J2_124_3477_n1958), 
        .A2(DP_OP_424J2_126_3477_n2885), .Y(DP_OP_424J2_126_3477_n2858) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1788 ( .A1(DP_OP_422J2_124_3477_n2265), 
        .A2(DP_OP_425J2_127_3477_n2577), .Y(DP_OP_424J2_126_3477_n2549) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1476 ( .A1(DP_OP_425J2_127_3477_n2261), 
        .A2(DP_OP_425J2_127_3477_n2269), .Y(DP_OP_425J2_127_3477_n2237) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1784 ( .A1(DP_OP_424J2_126_3477_n2569), 
        .A2(DP_OP_422J2_124_3477_n2577), .Y(DP_OP_424J2_126_3477_n2545) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1960 ( .A1(DP_OP_425J2_127_3477_n2745), 
        .A2(DP_OP_423J2_125_3477_n2753), .Y(DP_OP_425J2_127_3477_n2721) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1828 ( .A1(DP_OP_422J2_124_3477_n2745), 
        .A2(DP_OP_425J2_127_3477_n2621), .Y(DP_OP_425J2_127_3477_n2589) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1872 ( .A1(DP_OP_422J2_124_3477_n2789), 
        .A2(DP_OP_425J2_127_3477_n2665), .Y(DP_OP_425J2_127_3477_n2633) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2224 ( .A1(DP_OP_425J2_127_3477_n3007), 
        .A2(DP_OP_425J2_127_3477_n3015), .Y(DP_OP_425J2_127_3477_n2983) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1365 ( .A1(DP_OP_422J2_124_3477_n2134), 
        .A2(DP_OP_422J2_124_3477_n2139), .Y(DP_OP_422J2_124_3477_n2126) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1789 ( .A1(DP_OP_423J2_125_3477_n2662), 
        .A2(DP_OP_423J2_125_3477_n2577), .Y(DP_OP_424J2_126_3477_n2550) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2188 ( .A1(DP_OP_425J2_127_3477_n2085), 
        .A2(DP_OP_423J2_125_3477_n2974), .Y(DP_OP_423J2_125_3477_n2949) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1363 ( .A1(DP_OP_422J2_124_3477_n2132), 
        .A2(DP_OP_422J2_124_3477_n2139), .Y(DP_OP_422J2_124_3477_n2124) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2180 ( .A1(DP_OP_425J2_127_3477_n1997), 
        .A2(DP_OP_423J2_125_3477_n2973), .Y(DP_OP_424J2_126_3477_n2941) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1789 ( .A1(DP_OP_423J2_125_3477_n2398), 
        .A2(DP_OP_422J2_124_3477_n2577), .Y(DP_OP_422J2_124_3477_n2550) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2097 ( .A1(DP_OP_425J2_127_3477_n2750), 
        .A2(DP_OP_422J2_124_3477_n2885), .Y(DP_OP_422J2_124_3477_n2858) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1787 ( .A1(DP_OP_423J2_125_3477_n2572), 
        .A2(DP_OP_423J2_125_3477_n2577), .Y(DP_OP_423J2_125_3477_n2548) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2136 ( .A1(DP_OP_424J2_126_3477_n2921), 
        .A2(DP_OP_424J2_126_3477_n2929), .Y(DP_OP_424J2_126_3477_n2897) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1388 ( .A1(DP_OP_422J2_124_3477_n2877), 
        .A2(DP_OP_425J2_127_3477_n2181), .Y(DP_OP_424J2_126_3477_n2149) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1361 ( .A1(DP_OP_422J2_124_3477_n2834), 
        .A2(DP_OP_423J2_125_3477_n2139), .Y(DP_OP_423J2_125_3477_n2122) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1520 ( .A1(DP_OP_423J2_125_3477_n2217), 
        .A2(DP_OP_422J2_124_3477_n2313), .Y(DP_OP_424J2_126_3477_n2281) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1366 ( .A1(DP_OP_422J2_124_3477_n2927), 
        .A2(DP_OP_423J2_125_3477_n2139), .Y(DP_OP_424J2_126_3477_n2127) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1366 ( .A1(DP_OP_423J2_125_3477_n2135), 
        .A2(DP_OP_423J2_125_3477_n2139), .Y(DP_OP_423J2_125_3477_n2127) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2098 ( .A1(DP_OP_424J2_126_3477_n2795), 
        .A2(DP_OP_423J2_125_3477_n2885), .Y(DP_OP_423J2_125_3477_n2859) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2098 ( .A1(DP_OP_422J2_124_3477_n2883), 
        .A2(DP_OP_422J2_124_3477_n2885), .Y(DP_OP_422J2_124_3477_n2859) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1785 ( .A1(DP_OP_423J2_125_3477_n2570), 
        .A2(DP_OP_423J2_125_3477_n2577), .Y(DP_OP_423J2_125_3477_n2546) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2095 ( .A1(DP_OP_423J2_125_3477_n2880), 
        .A2(DP_OP_423J2_125_3477_n2885), .Y(DP_OP_423J2_125_3477_n2856) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1364 ( .A1(DP_OP_424J2_126_3477_n2133), 
        .A2(DP_OP_425J2_127_3477_n2139), .Y(DP_OP_424J2_126_3477_n2125) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1924 ( .A1(DP_OP_424J2_126_3477_n2613), 
        .A2(DP_OP_423J2_125_3477_n2710), .Y(DP_OP_423J2_125_3477_n2685) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2056 ( .A1(DP_OP_425J2_127_3477_n2217), 
        .A2(DP_OP_423J2_125_3477_n2842), .Y(DP_OP_423J2_125_3477_n2817) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1828 ( .A1(DP_OP_424J2_126_3477_n2613), 
        .A2(DP_OP_422J2_124_3477_n2621), .Y(DP_OP_424J2_126_3477_n2589) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1790 ( .A1(DP_OP_423J2_125_3477_n2575), 
        .A2(DP_OP_423J2_125_3477_n2577), .Y(DP_OP_423J2_125_3477_n2551) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1484 ( .A1(DP_OP_423J2_125_3477_n2261), 
        .A2(DP_OP_423J2_125_3477_n2270), .Y(DP_OP_423J2_125_3477_n2245) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1300 ( .A1(DP_OP_425J2_127_3477_n2833), 
        .A2(DP_OP_422J2_124_3477_n2093), .Y(DP_OP_424J2_126_3477_n2061) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2100 ( .A1(DP_OP_423J2_125_3477_n2877), 
        .A2(DP_OP_423J2_125_3477_n2886), .Y(DP_OP_423J2_125_3477_n2861) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1220 ( .A1(DP_OP_423J2_125_3477_n1997), 
        .A2(DP_OP_423J2_125_3477_n2006), .Y(DP_OP_423J2_125_3477_n1981) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1790 ( .A1(DP_OP_423J2_125_3477_n2663), 
        .A2(DP_OP_423J2_125_3477_n2577), .Y(DP_OP_424J2_126_3477_n2551) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2224 ( .A1(DP_OP_424J2_126_3477_n3007), 
        .A2(DP_OP_424J2_126_3477_n3015), .Y(DP_OP_424J2_126_3477_n2983) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1364 ( .A1(DP_OP_424J2_126_3477_n2705), 
        .A2(DP_OP_422J2_124_3477_n2139), .Y(DP_OP_422J2_124_3477_n2125) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1365 ( .A1(DP_OP_423J2_125_3477_n2134), 
        .A2(DP_OP_423J2_125_3477_n2139), .Y(DP_OP_423J2_125_3477_n2126) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2098 ( .A1(DP_OP_424J2_126_3477_n2883), 
        .A2(DP_OP_424J2_126_3477_n2885), .Y(DP_OP_424J2_126_3477_n2859) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1704 ( .A1(DP_OP_423J2_125_3477_n2481), 
        .A2(DP_OP_423J2_125_3477_n2490), .Y(DP_OP_423J2_125_3477_n2465) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2144 ( .A1(DP_OP_423J2_125_3477_n2921), 
        .A2(DP_OP_423J2_125_3477_n2930), .Y(DP_OP_423J2_125_3477_n2905) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2097 ( .A1(DP_OP_423J2_125_3477_n1958), 
        .A2(DP_OP_424J2_126_3477_n2885), .Y(DP_OP_425J2_127_3477_n2858) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1520 ( .A1(DP_OP_423J2_125_3477_n2305), 
        .A2(DP_OP_423J2_125_3477_n2313), .Y(DP_OP_423J2_125_3477_n2281) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1789 ( .A1(DP_OP_423J2_125_3477_n2266), 
        .A2(DP_OP_425J2_127_3477_n2577), .Y(DP_OP_425J2_127_3477_n2550) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1432 ( .A1(DP_OP_423J2_125_3477_n2217), 
        .A2(DP_OP_423J2_125_3477_n2225), .Y(DP_OP_423J2_125_3477_n2193) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2136 ( .A1(DP_OP_423J2_125_3477_n2921), 
        .A2(DP_OP_423J2_125_3477_n2929), .Y(DP_OP_423J2_125_3477_n2897) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1388 ( .A1(DP_OP_424J2_126_3477_n2261), 
        .A2(DP_OP_423J2_125_3477_n2181), .Y(DP_OP_423J2_125_3477_n2149) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1344 ( .A1(DP_OP_424J2_126_3477_n2217), 
        .A2(DP_OP_424J2_126_3477_n2137), .Y(DP_OP_423J2_125_3477_n2105) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2180 ( .A1(DP_OP_424J2_126_3477_n2877), 
        .A2(DP_OP_423J2_125_3477_n2973), .Y(DP_OP_423J2_125_3477_n2941) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1756 ( .A1(DP_OP_423J2_125_3477_n2525), 
        .A2(DP_OP_423J2_125_3477_n2535), .Y(DP_OP_423J2_125_3477_n2517) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1300 ( .A1(DP_OP_422J2_124_3477_n2877), 
        .A2(DP_OP_423J2_125_3477_n2093), .Y(DP_OP_423J2_125_3477_n2061) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1256 ( .A1(DP_OP_425J2_127_3477_n2789), 
        .A2(DP_OP_422J2_124_3477_n2049), .Y(DP_OP_423J2_125_3477_n2017) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2224 ( .A1(DP_OP_423J2_125_3477_n3007), 
        .A2(DP_OP_425J2_127_3477_n3015), .Y(DP_OP_423J2_125_3477_n2983) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1872 ( .A1(DP_OP_424J2_126_3477_n2569), 
        .A2(DP_OP_423J2_125_3477_n2665), .Y(DP_OP_423J2_125_3477_n2633) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1828 ( .A1(DP_OP_423J2_125_3477_n2613), 
        .A2(DP_OP_423J2_125_3477_n2621), .Y(DP_OP_423J2_125_3477_n2589) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1960 ( .A1(DP_OP_423J2_125_3477_n2745), 
        .A2(DP_OP_423J2_125_3477_n2753), .Y(DP_OP_423J2_125_3477_n2721) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1786 ( .A1(DP_OP_423J2_125_3477_n2571), 
        .A2(DP_OP_423J2_125_3477_n2577), .Y(DP_OP_423J2_125_3477_n2547) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1476 ( .A1(DP_OP_423J2_125_3477_n2261), 
        .A2(DP_OP_422J2_124_3477_n2269), .Y(DP_OP_423J2_125_3477_n2237) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1256 ( .A1(DP_OP_424J2_126_3477_n2789), 
        .A2(DP_OP_422J2_124_3477_n2049), .Y(DP_OP_422J2_124_3477_n2017) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2224 ( .A1(DP_OP_422J2_124_3477_n3007), 
        .A2(DP_OP_422J2_124_3477_n3015), .Y(DP_OP_422J2_124_3477_n2983) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1872 ( .A1(DP_OP_425J2_127_3477_n2525), 
        .A2(DP_OP_425J2_127_3477_n2665), .Y(DP_OP_422J2_124_3477_n2633) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1476 ( .A1(DP_OP_422J2_124_3477_n2261), 
        .A2(DP_OP_422J2_124_3477_n2269), .Y(DP_OP_422J2_124_3477_n2237) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1787 ( .A1(DP_OP_424J2_126_3477_n2572), 
        .A2(DP_OP_422J2_124_3477_n2577), .Y(DP_OP_424J2_126_3477_n2548) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2096 ( .A1(DP_OP_422J2_124_3477_n2045), 
        .A2(DP_OP_423J2_125_3477_n2885), .Y(DP_OP_423J2_125_3477_n2857) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1696 ( .A1(DP_OP_423J2_125_3477_n2481), 
        .A2(DP_OP_423J2_125_3477_n2489), .Y(DP_OP_423J2_125_3477_n2457) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1652 ( .A1(DP_OP_423J2_125_3477_n2437), 
        .A2(DP_OP_423J2_125_3477_n2445), .Y(DP_OP_423J2_125_3477_n2413) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1608 ( .A1(DP_OP_422J2_124_3477_n2569), 
        .A2(DP_OP_423J2_125_3477_n2401), .Y(DP_OP_423J2_125_3477_n2369) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1363 ( .A1(DP_OP_423J2_125_3477_n2924), 
        .A2(DP_OP_425J2_127_3477_n2139), .Y(DP_OP_425J2_127_3477_n2124) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1564 ( .A1(DP_OP_422J2_124_3477_n2613), 
        .A2(DP_OP_423J2_125_3477_n2357), .Y(DP_OP_423J2_125_3477_n2325) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2096 ( .A1(DP_OP_423J2_125_3477_n1957), 
        .A2(DP_OP_423J2_125_3477_n2885), .Y(DP_OP_425J2_127_3477_n2857) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2197 ( .A1(DP_OP_423J2_125_3477_n1998), 
        .A2(DP_OP_422J2_124_3477_n2975), .Y(DP_OP_422J2_124_3477_n2958) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1581 ( .A1(DP_OP_424J2_126_3477_n2482), 
        .A2(DP_OP_422J2_124_3477_n2359), .Y(DP_OP_422J2_124_3477_n2342) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1624 ( .A1(DP_OP_422J2_124_3477_n2569), 
        .A2(DP_OP_423J2_125_3477_n2403), .Y(DP_OP_423J2_125_3477_n2385) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1449 ( .A1(DP_OP_422J2_124_3477_n2218), 
        .A2(DP_OP_422J2_124_3477_n2227), .Y(DP_OP_422J2_124_3477_n2210) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1362 ( .A1(DP_OP_424J2_126_3477_n2835), 
        .A2(DP_OP_425J2_127_3477_n2139), .Y(DP_OP_425J2_127_3477_n2123) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1788 ( .A1(DP_OP_423J2_125_3477_n2265), 
        .A2(DP_OP_425J2_127_3477_n2577), .Y(DP_OP_425J2_127_3477_n2549) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2095 ( .A1(DP_OP_422J2_124_3477_n2880), 
        .A2(DP_OP_422J2_124_3477_n2885), .Y(DP_OP_422J2_124_3477_n2856) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2020 ( .A1(DP_OP_425J2_127_3477_n2789), 
        .A2(DP_OP_425J2_127_3477_n2799), .Y(DP_OP_425J2_127_3477_n2781) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1844 ( .A1(DP_OP_423J2_125_3477_n2217), 
        .A2(DP_OP_425J2_127_3477_n2623), .Y(DP_OP_425J2_127_3477_n2605) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2240 ( .A1(DP_OP_425J2_127_3477_n3007), 
        .A2(DP_OP_425J2_127_3477_n3017), .Y(DP_OP_425J2_127_3477_n2999) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1668 ( .A1(DP_OP_423J2_125_3477_n2613), 
        .A2(DP_OP_425J2_127_3477_n2447), .Y(DP_OP_425J2_127_3477_n2429) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1786 ( .A1(DP_OP_423J2_125_3477_n2263), 
        .A2(DP_OP_425J2_127_3477_n2577), .Y(DP_OP_425J2_127_3477_n2547) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2108 ( .A1(DP_OP_423J2_125_3477_n2877), 
        .A2(DP_OP_422J2_124_3477_n2887), .Y(DP_OP_423J2_125_3477_n2869) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2095 ( .A1(DP_OP_424J2_126_3477_n2880), 
        .A2(DP_OP_424J2_126_3477_n2885), .Y(DP_OP_424J2_126_3477_n2856) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1580 ( .A1(DP_OP_425J2_127_3477_n2481), 
        .A2(DP_OP_423J2_125_3477_n2359), .Y(DP_OP_423J2_125_3477_n2341) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1365 ( .A1(DP_OP_425J2_127_3477_n2134), 
        .A2(DP_OP_425J2_127_3477_n2139), .Y(DP_OP_425J2_127_3477_n2126) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1264 ( .A1(DP_OP_422J2_124_3477_n3007), 
        .A2(DP_OP_425J2_127_3477_n2050), .Y(DP_OP_424J2_126_3477_n2025) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2093 ( .A1(DP_OP_424J2_126_3477_n2878), 
        .A2(DP_OP_424J2_126_3477_n2885), .Y(DP_OP_424J2_126_3477_n2854) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1366 ( .A1(DP_OP_425J2_127_3477_n2135), 
        .A2(DP_OP_425J2_127_3477_n2139), .Y(DP_OP_425J2_127_3477_n2127) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1788 ( .A1(DP_OP_423J2_125_3477_n2573), 
        .A2(DP_OP_423J2_125_3477_n2577), .Y(DP_OP_423J2_125_3477_n2549) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2144 ( .A1(DP_OP_424J2_126_3477_n2921), 
        .A2(DP_OP_425J2_127_3477_n2930), .Y(DP_OP_424J2_126_3477_n2905) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1785 ( .A1(DP_OP_422J2_124_3477_n2262), 
        .A2(DP_OP_422J2_124_3477_n2577), .Y(DP_OP_424J2_126_3477_n2546) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1748 ( .A1(DP_OP_423J2_125_3477_n2613), 
        .A2(DP_OP_425J2_127_3477_n2534), .Y(DP_OP_424J2_126_3477_n2509) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1844 ( .A1(DP_OP_423J2_125_3477_n2613), 
        .A2(DP_OP_423J2_125_3477_n2623), .Y(DP_OP_423J2_125_3477_n2605) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2241 ( .A1(DP_OP_424J2_126_3477_n3008), 
        .A2(DP_OP_422J2_124_3477_n3017), .Y(DP_OP_424J2_126_3477_n3000) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1176 ( .A1(DP_OP_425J2_127_3477_n2965), 
        .A2(DP_OP_424J2_126_3477_n1962), .Y(DP_OP_424J2_126_3477_n1937) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1361 ( .A1(DP_OP_422J2_124_3477_n2922), 
        .A2(DP_OP_423J2_125_3477_n2139), .Y(DP_OP_424J2_126_3477_n2122) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1564 ( .A1(DP_OP_424J2_126_3477_n2481), 
        .A2(DP_OP_422J2_124_3477_n2357), .Y(DP_OP_422J2_124_3477_n2325) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2180 ( .A1(DP_OP_425J2_127_3477_n2833), 
        .A2(DP_OP_422J2_124_3477_n2973), .Y(DP_OP_422J2_124_3477_n2941) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1362 ( .A1(DP_OP_424J2_126_3477_n2219), 
        .A2(DP_OP_423J2_125_3477_n2139), .Y(DP_OP_423J2_125_3477_n2123) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1364 ( .A1(DP_OP_425J2_127_3477_n2133), 
        .A2(DP_OP_425J2_127_3477_n2139), .Y(DP_OP_425J2_127_3477_n2125) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2098 ( .A1(DP_OP_422J2_124_3477_n3013), 
        .A2(DP_OP_422J2_124_3477_n2885), .Y(DP_OP_425J2_127_3477_n2859) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1790 ( .A1(DP_OP_423J2_125_3477_n2267), 
        .A2(DP_OP_425J2_127_3477_n2577), .Y(DP_OP_425J2_127_3477_n2551) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2232 ( .A1(DP_OP_422J2_124_3477_n3007), 
        .A2(DP_OP_422J2_124_3477_n3016), .Y(DP_OP_422J2_124_3477_n2991) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1484 ( .A1(DP_OP_425J2_127_3477_n2261), 
        .A2(DP_OP_425J2_127_3477_n2270), .Y(DP_OP_425J2_127_3477_n2245) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2108 ( .A1(DP_OP_424J2_126_3477_n2877), 
        .A2(DP_OP_424J2_126_3477_n2887), .Y(DP_OP_424J2_126_3477_n2869) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1748 ( .A1(DP_OP_425J2_127_3477_n2525), 
        .A2(DP_OP_425J2_127_3477_n2534), .Y(DP_OP_425J2_127_3477_n2509) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1785 ( .A1(DP_OP_423J2_125_3477_n2262), 
        .A2(DP_OP_425J2_127_3477_n2577), .Y(DP_OP_425J2_127_3477_n2546) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1617 ( .A1(DP_OP_422J2_124_3477_n2570), 
        .A2(DP_OP_423J2_125_3477_n2402), .Y(DP_OP_423J2_125_3477_n2378) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1880 ( .A1(DP_OP_422J2_124_3477_n2789), 
        .A2(DP_OP_425J2_127_3477_n2666), .Y(DP_OP_425J2_127_3477_n2641) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1660 ( .A1(DP_OP_423J2_125_3477_n2613), 
        .A2(DP_OP_425J2_127_3477_n2446), .Y(DP_OP_425J2_127_3477_n2421) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2233 ( .A1(DP_OP_423J2_125_3477_n3008), 
        .A2(DP_OP_423J2_125_3477_n3016), .Y(DP_OP_423J2_125_3477_n2992) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1360 ( .A1(DP_OP_422J2_124_3477_n2129), 
        .A2(DP_OP_422J2_124_3477_n2139), .Y(DP_OP_422J2_124_3477_n2121) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1616 ( .A1(DP_OP_424J2_126_3477_n2569), 
        .A2(DP_OP_425J2_127_3477_n2402), .Y(DP_OP_425J2_127_3477_n2377) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1617 ( .A1(DP_OP_423J2_125_3477_n2526), 
        .A2(DP_OP_423J2_125_3477_n2402), .Y(DP_OP_422J2_124_3477_n2378) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1352 ( .A1(DP_OP_423J2_125_3477_n2921), 
        .A2(DP_OP_425J2_127_3477_n2138), .Y(DP_OP_425J2_127_3477_n2113) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2012 ( .A1(DP_OP_425J2_127_3477_n2789), 
        .A2(DP_OP_425J2_127_3477_n2798), .Y(DP_OP_425J2_127_3477_n2773) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1396 ( .A1(DP_OP_423J2_125_3477_n2877), 
        .A2(DP_OP_425J2_127_3477_n2182), .Y(DP_OP_425J2_127_3477_n2157) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2094 ( .A1(DP_OP_423J2_125_3477_n2967), 
        .A2(DP_OP_424J2_126_3477_n2885), .Y(DP_OP_424J2_126_3477_n2855) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2093 ( .A1(DP_OP_425J2_127_3477_n2878), 
        .A2(DP_OP_424J2_126_3477_n2885), .Y(DP_OP_425J2_127_3477_n2854) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1264 ( .A1(DP_OP_423J2_125_3477_n3007), 
        .A2(DP_OP_425J2_127_3477_n2050), .Y(DP_OP_425J2_127_3477_n2025) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1573 ( .A1(DP_OP_424J2_126_3477_n2482), 
        .A2(DP_OP_422J2_124_3477_n2358), .Y(DP_OP_422J2_124_3477_n2334) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2196 ( .A1(DP_OP_423J2_125_3477_n1997), 
        .A2(DP_OP_422J2_124_3477_n2975), .Y(DP_OP_422J2_124_3477_n2957) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1924 ( .A1(DP_OP_424J2_126_3477_n2217), 
        .A2(DP_OP_425J2_127_3477_n2710), .Y(DP_OP_425J2_127_3477_n2685) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1932 ( .A1(DP_OP_422J2_124_3477_n2701), 
        .A2(DP_OP_422J2_124_3477_n2711), .Y(DP_OP_422J2_124_3477_n2693) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1704 ( .A1(DP_OP_425J2_127_3477_n2481), 
        .A2(DP_OP_425J2_127_3477_n2490), .Y(DP_OP_425J2_127_3477_n2465) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2144 ( .A1(DP_OP_425J2_127_3477_n2921), 
        .A2(DP_OP_425J2_127_3477_n2930), .Y(DP_OP_425J2_127_3477_n2905) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2108 ( .A1(DP_OP_422J2_124_3477_n2877), 
        .A2(DP_OP_422J2_124_3477_n2887), .Y(DP_OP_422J2_124_3477_n2869) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1228 ( .A1(DP_OP_423J2_125_3477_n1997), 
        .A2(DP_OP_423J2_125_3477_n2007), .Y(DP_OP_423J2_125_3477_n1989) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1616 ( .A1(DP_OP_423J2_125_3477_n2525), 
        .A2(DP_OP_424J2_126_3477_n2402), .Y(DP_OP_422J2_124_3477_n2377) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2101 ( .A1(DP_OP_422J2_124_3477_n2878), 
        .A2(DP_OP_422J2_124_3477_n2886), .Y(DP_OP_422J2_124_3477_n2862) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2094 ( .A1(DP_OP_425J2_127_3477_n2747), 
        .A2(DP_OP_422J2_124_3477_n2885), .Y(DP_OP_422J2_124_3477_n2855) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1785 ( .A1(DP_OP_422J2_124_3477_n2570), 
        .A2(DP_OP_422J2_124_3477_n2577), .Y(DP_OP_422J2_124_3477_n2546) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2013 ( .A1(DP_OP_423J2_125_3477_n2790), 
        .A2(DP_OP_423J2_125_3477_n2798), .Y(DP_OP_423J2_125_3477_n2774) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2232 ( .A1(DP_OP_425J2_127_3477_n3007), 
        .A2(DP_OP_423J2_125_3477_n3016), .Y(DP_OP_425J2_127_3477_n2991) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1176 ( .A1(DP_OP_424J2_126_3477_n3007), 
        .A2(DP_OP_424J2_126_3477_n1962), .Y(DP_OP_425J2_127_3477_n1937) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2064 ( .A1(DP_OP_422J2_124_3477_n2833), 
        .A2(DP_OP_422J2_124_3477_n2843), .Y(DP_OP_422J2_124_3477_n2825) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1916 ( .A1(DP_OP_422J2_124_3477_n2129), 
        .A2(DP_OP_423J2_125_3477_n2709), .Y(DP_OP_424J2_126_3477_n2677) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2188 ( .A1(DP_OP_425J2_127_3477_n2965), 
        .A2(DP_OP_425J2_127_3477_n2974), .Y(DP_OP_425J2_127_3477_n2949) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1360 ( .A1(DP_OP_422J2_124_3477_n2833), 
        .A2(DP_OP_423J2_125_3477_n2139), .Y(DP_OP_423J2_125_3477_n2121) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2188 ( .A1(DP_OP_425J2_127_3477_n2833), 
        .A2(DP_OP_422J2_124_3477_n2974), .Y(DP_OP_422J2_124_3477_n2949) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1792 ( .A1(DP_OP_423J2_125_3477_n2261), 
        .A2(DP_OP_425J2_127_3477_n2578), .Y(DP_OP_425J2_127_3477_n2553) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1228 ( .A1(DP_OP_424J2_126_3477_n2833), 
        .A2(DP_OP_422J2_124_3477_n2007), .Y(DP_OP_422J2_124_3477_n1989) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1176 ( .A1(DP_OP_425J2_127_3477_n2085), 
        .A2(DP_OP_422J2_124_3477_n1962), .Y(DP_OP_422J2_124_3477_n1937) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1228 ( .A1(DP_OP_425J2_127_3477_n2921), 
        .A2(DP_OP_422J2_124_3477_n2007), .Y(DP_OP_424J2_126_3477_n1989) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2095 ( .A1(DP_OP_422J2_124_3477_n3010), 
        .A2(DP_OP_424J2_126_3477_n2885), .Y(DP_OP_425J2_127_3477_n2856) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1361 ( .A1(DP_OP_423J2_125_3477_n2922), 
        .A2(DP_OP_425J2_127_3477_n2139), .Y(DP_OP_425J2_127_3477_n2122) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1932 ( .A1(DP_OP_422J2_124_3477_n2129), 
        .A2(DP_OP_424J2_126_3477_n2711), .Y(DP_OP_424J2_126_3477_n2693) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1787 ( .A1(DP_OP_425J2_127_3477_n2572), 
        .A2(DP_OP_425J2_127_3477_n2577), .Y(DP_OP_425J2_127_3477_n2548) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1177 ( .A1(DP_OP_422J2_124_3477_n3008), 
        .A2(DP_OP_423J2_125_3477_n1962), .Y(DP_OP_423J2_125_3477_n1938) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1353 ( .A1(DP_OP_422J2_124_3477_n2922), 
        .A2(DP_OP_423J2_125_3477_n2138), .Y(DP_OP_424J2_126_3477_n2114) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1360 ( .A1(DP_OP_422J2_124_3477_n2921), 
        .A2(DP_OP_422J2_124_3477_n2139), .Y(DP_OP_424J2_126_3477_n2121) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1536 ( .A1(DP_OP_423J2_125_3477_n2305), 
        .A2(DP_OP_423J2_125_3477_n2315), .Y(DP_OP_423J2_125_3477_n2297) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2152 ( .A1(DP_OP_423J2_125_3477_n2921), 
        .A2(DP_OP_423J2_125_3477_n2931), .Y(DP_OP_423J2_125_3477_n2913) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1617 ( .A1(DP_OP_422J2_124_3477_n2658), 
        .A2(DP_OP_424J2_126_3477_n2402), .Y(DP_OP_424J2_126_3477_n2378) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1220 ( .A1(DP_OP_425J2_127_3477_n1997), 
        .A2(DP_OP_425J2_127_3477_n2006), .Y(DP_OP_425J2_127_3477_n1981) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2196 ( .A1(DP_OP_425J2_127_3477_n2085), 
        .A2(DP_OP_424J2_126_3477_n2975), .Y(DP_OP_423J2_125_3477_n2957) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1888 ( .A1(DP_OP_423J2_125_3477_n2745), 
        .A2(DP_OP_425J2_127_3477_n2667), .Y(DP_OP_424J2_126_3477_n2649) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1536 ( .A1(DP_OP_423J2_125_3477_n2217), 
        .A2(DP_OP_424J2_126_3477_n2315), .Y(DP_OP_424J2_126_3477_n2297) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2152 ( .A1(DP_OP_422J2_124_3477_n2921), 
        .A2(DP_OP_422J2_124_3477_n2931), .Y(DP_OP_422J2_124_3477_n2913) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1177 ( .A1(DP_OP_425J2_127_3477_n2086), 
        .A2(DP_OP_422J2_124_3477_n1962), .Y(DP_OP_422J2_124_3477_n1938) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1448 ( .A1(DP_OP_424J2_126_3477_n2217), 
        .A2(DP_OP_424J2_126_3477_n2227), .Y(DP_OP_424J2_126_3477_n2209) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1360 ( .A1(DP_OP_424J2_126_3477_n2833), 
        .A2(DP_OP_425J2_127_3477_n2139), .Y(DP_OP_425J2_127_3477_n2121) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1793 ( .A1(DP_OP_422J2_124_3477_n2570), 
        .A2(DP_OP_422J2_124_3477_n2578), .Y(DP_OP_422J2_124_3477_n2554) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1668 ( .A1(DP_OP_422J2_124_3477_n2613), 
        .A2(DP_OP_424J2_126_3477_n2447), .Y(DP_OP_424J2_126_3477_n2429) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1228 ( .A1(DP_OP_425J2_127_3477_n1997), 
        .A2(DP_OP_425J2_127_3477_n2007), .Y(DP_OP_425J2_127_3477_n1989) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1668 ( .A1(DP_OP_423J2_125_3477_n2481), 
        .A2(DP_OP_422J2_124_3477_n2447), .Y(DP_OP_422J2_124_3477_n2429) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1932 ( .A1(DP_OP_422J2_124_3477_n2833), 
        .A2(DP_OP_425J2_127_3477_n2711), .Y(DP_OP_425J2_127_3477_n2693) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2094 ( .A1(DP_OP_425J2_127_3477_n2175), 
        .A2(DP_OP_423J2_125_3477_n2885), .Y(DP_OP_423J2_125_3477_n2855) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2196 ( .A1(DP_OP_425J2_127_3477_n2965), 
        .A2(DP_OP_425J2_127_3477_n2975), .Y(DP_OP_425J2_127_3477_n2957) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1448 ( .A1(DP_OP_425J2_127_3477_n2217), 
        .A2(DP_OP_425J2_127_3477_n2227), .Y(DP_OP_425J2_127_3477_n2209) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2240 ( .A1(DP_OP_422J2_124_3477_n3007), 
        .A2(DP_OP_422J2_124_3477_n3017), .Y(DP_OP_422J2_124_3477_n2999) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1844 ( .A1(DP_OP_424J2_126_3477_n2613), 
        .A2(DP_OP_424J2_126_3477_n2623), .Y(DP_OP_424J2_126_3477_n2605) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1786 ( .A1(DP_OP_423J2_125_3477_n2659), 
        .A2(DP_OP_425J2_127_3477_n2577), .Y(DP_OP_424J2_126_3477_n2547) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2100 ( .A1(DP_OP_422J2_124_3477_n2877), 
        .A2(DP_OP_422J2_124_3477_n2886), .Y(DP_OP_422J2_124_3477_n2861) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2094 ( .A1(DP_OP_425J2_127_3477_n2879), 
        .A2(DP_OP_423J2_125_3477_n2885), .Y(DP_OP_425J2_127_3477_n2855) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1787 ( .A1(DP_OP_423J2_125_3477_n2396), 
        .A2(DP_OP_422J2_124_3477_n2577), .Y(DP_OP_422J2_124_3477_n2548) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2144 ( .A1(DP_OP_422J2_124_3477_n2921), 
        .A2(DP_OP_422J2_124_3477_n2930), .Y(DP_OP_422J2_124_3477_n2905) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1704 ( .A1(DP_OP_422J2_124_3477_n2481), 
        .A2(DP_OP_422J2_124_3477_n2490), .Y(DP_OP_422J2_124_3477_n2465) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1572 ( .A1(DP_OP_424J2_126_3477_n2481), 
        .A2(DP_OP_422J2_124_3477_n2358), .Y(DP_OP_422J2_124_3477_n2333) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1924 ( .A1(DP_OP_422J2_124_3477_n2701), 
        .A2(DP_OP_422J2_124_3477_n2710), .Y(DP_OP_422J2_124_3477_n2685) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1404 ( .A1(DP_OP_422J2_124_3477_n2877), 
        .A2(DP_OP_424J2_126_3477_n2183), .Y(DP_OP_424J2_126_3477_n2165) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1264 ( .A1(DP_OP_424J2_126_3477_n2789), 
        .A2(DP_OP_422J2_124_3477_n2050), .Y(DP_OP_422J2_124_3477_n2025) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2108 ( .A1(DP_OP_425J2_127_3477_n2877), 
        .A2(DP_OP_425J2_127_3477_n2887), .Y(DP_OP_425J2_127_3477_n2869) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2093 ( .A1(DP_OP_422J2_124_3477_n2878), 
        .A2(DP_OP_422J2_124_3477_n2885), .Y(DP_OP_422J2_124_3477_n2854) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1789 ( .A1(DP_OP_423J2_125_3477_n2574), 
        .A2(DP_OP_423J2_125_3477_n2577), .Y(DP_OP_423J2_125_3477_n2550) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2241 ( .A1(DP_OP_422J2_124_3477_n3008), 
        .A2(DP_OP_422J2_124_3477_n3017), .Y(DP_OP_422J2_124_3477_n3000) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1756 ( .A1(DP_OP_423J2_125_3477_n2437), 
        .A2(DP_OP_422J2_124_3477_n2535), .Y(DP_OP_422J2_124_3477_n2517) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1361 ( .A1(DP_OP_422J2_124_3477_n2130), 
        .A2(DP_OP_422J2_124_3477_n2139), .Y(DP_OP_422J2_124_3477_n2122) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2097 ( .A1(DP_OP_425J2_127_3477_n2178), 
        .A2(DP_OP_423J2_125_3477_n2885), .Y(DP_OP_423J2_125_3477_n2858) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1786 ( .A1(DP_OP_422J2_124_3477_n2571), 
        .A2(DP_OP_422J2_124_3477_n2577), .Y(DP_OP_422J2_124_3477_n2547) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1404 ( .A1(DP_OP_425J2_127_3477_n2305), 
        .A2(DP_OP_422J2_124_3477_n2183), .Y(DP_OP_422J2_124_3477_n2165) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1756 ( .A1(DP_OP_422J2_124_3477_n2305), 
        .A2(DP_OP_425J2_127_3477_n2535), .Y(DP_OP_424J2_126_3477_n2517) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U95 ( .A1(DP_OP_424J2_126_3477_n101), .A2(
        DP_OP_424J2_126_3477_n104), .Y(DP_OP_424J2_126_3477_n99) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U95 ( .A1(DP_OP_422J2_124_3477_n101), .A2(
        DP_OP_422J2_124_3477_n104), .Y(DP_OP_422J2_124_3477_n99) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U75 ( .A1(DP_OP_422J2_124_3477_n87), .A2(
        DP_OP_422J2_124_3477_n90), .Y(DP_OP_422J2_124_3477_n85) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U75 ( .A1(DP_OP_424J2_126_3477_n87), .A2(
        DP_OP_424J2_126_3477_n90), .Y(DP_OP_424J2_126_3477_n85) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U155 ( .A1(DP_OP_422J2_124_3477_n281), .A2(
        DP_OP_422J2_124_3477_n282), .Y(DP_OP_422J2_124_3477_n137) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U155 ( .A1(DP_OP_423J2_125_3477_n281), .A2(
        DP_OP_423J2_125_3477_n282), .Y(DP_OP_423J2_125_3477_n137) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U155 ( .A1(DP_OP_425J2_127_3477_n281), .A2(
        DP_OP_425J2_127_3477_n282), .Y(DP_OP_425J2_127_3477_n137) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U149 ( .A1(DP_OP_422J2_124_3477_n137), .A2(
        DP_OP_422J2_124_3477_n144), .Y(DP_OP_422J2_124_3477_n135) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U149 ( .A1(DP_OP_423J2_125_3477_n137), .A2(
        DP_OP_423J2_125_3477_n144), .Y(DP_OP_423J2_125_3477_n135) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U149 ( .A1(DP_OP_425J2_127_3477_n137), .A2(
        DP_OP_425J2_127_3477_n144), .Y(DP_OP_425J2_127_3477_n135) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U149 ( .A1(DP_OP_424J2_126_3477_n137), .A2(
        DP_OP_424J2_126_3477_n144), .Y(DP_OP_424J2_126_3477_n135) );
  AO221X1_HVT U3 ( .A1(1'b1), .A2(n567), .A3(n497), .A4(conv2_sum_b[20]), .A5(
        n270), .Y(n601) );
  AO221X1_HVT U4 ( .A1(1'b1), .A2(n698), .A3(tmp_big2[20]), .A4(n171), .A5(
        n172), .Y(n731) );
  AO221X1_HVT U5 ( .A1(1'b1), .A2(n632), .A3(n502), .A4(conv2_sum_d[20]), .A5(
        n141), .Y(n665) );
  AO221X1_HVT U6 ( .A1(1'b1), .A2(n578), .A3(n495), .A4(conv2_sum_b[12]), .A5(
        n139), .Y(n581) );
  AO221X1_HVT U7 ( .A1(1'b1), .A2(n622), .A3(n522), .A4(conv2_sum_d[28]), .A5(
        n119), .Y(n623) );
  AO221X1_HVT U8 ( .A1(1'b1), .A2(n557), .A3(n520), .A4(conv2_sum_b[28]), .A5(
        n117), .Y(n558) );
  AO221X1_HVT U9 ( .A1(1'b1), .A2(n645), .A3(n5001), .A4(conv2_sum_d[12]), 
        .A5(n115), .Y(n648) );
  AO221X1_HVT U10 ( .A1(1'b1), .A2(n685), .A3(tmp_big2[28]), .A4(n81), .A5(n82), .Y(n686) );
  OA221X1_HVT U11 ( .A1(1'b0), .A2(DP_OP_424J2_126_3477_n70), .A3(
        DP_OP_424J2_126_3477_n65), .A4(DP_OP_424J2_126_3477_n149), .A5(n226), 
        .Y(DP_OP_424J2_126_3477_n62) );
  OA221X1_HVT U12 ( .A1(1'b0), .A2(DP_OP_422J2_124_3477_n70), .A3(
        DP_OP_422J2_124_3477_n65), .A4(DP_OP_422J2_124_3477_n149), .A5(n223), 
        .Y(DP_OP_422J2_124_3477_n62) );
  OA221X1_HVT U13 ( .A1(1'b0), .A2(n664), .A3(conv2_sum_c[16]), .A4(n494), 
        .A5(n214), .Y(n491) );
  OA221X1_HVT U14 ( .A1(1'b0), .A2(DP_OP_425J2_127_3477_n70), .A3(
        DP_OP_425J2_127_3477_n65), .A4(DP_OP_425J2_127_3477_n149), .A5(n150), 
        .Y(DP_OP_425J2_127_3477_n62) );
  OA221X1_HVT U15 ( .A1(1'b0), .A2(DP_OP_423J2_125_3477_n70), .A3(
        DP_OP_423J2_125_3477_n65), .A4(DP_OP_423J2_125_3477_n149), .A5(n147), 
        .Y(DP_OP_423J2_125_3477_n62) );
  INVX2_HVT U16 ( .A(n403), .Y(n381) );
  OAI21X1_HVT U17 ( .A1(DP_OP_422J2_124_3477_n163), .A2(
        DP_OP_422J2_124_3477_n183), .A3(DP_OP_422J2_124_3477_n164), .Y(
        DP_OP_422J2_124_3477_n162) );
  OAI21X1_HVT U18 ( .A1(DP_OP_424J2_126_3477_n163), .A2(
        DP_OP_424J2_126_3477_n183), .A3(DP_OP_424J2_126_3477_n164), .Y(
        DP_OP_424J2_126_3477_n162) );
  NOR2X0_HVT U19 ( .A1(DP_OP_423J2_125_3477_n2482), .A2(
        DP_OP_422J2_124_3477_n2445), .Y(DP_OP_422J2_124_3477_n2414) );
  NOR2X0_HVT U20 ( .A1(DP_OP_423J2_125_3477_n2484), .A2(
        DP_OP_422J2_124_3477_n2445), .Y(DP_OP_422J2_124_3477_n2416) );
  NOR2X0_HVT U21 ( .A1(DP_OP_423J2_125_3477_n2481), .A2(
        DP_OP_422J2_124_3477_n2445), .Y(DP_OP_422J2_124_3477_n2413) );
  NOR2X0_HVT U22 ( .A1(DP_OP_422J2_124_3477_n3007), .A2(
        DP_OP_424J2_126_3477_n2051), .Y(DP_OP_424J2_126_3477_n2033) );
  OR2X1_HVT U23 ( .A1(DP_OP_422J2_124_3477_n3006), .A2(
        DP_OP_424J2_126_3477_n2051), .Y(DP_OP_424J2_126_3477_n2032) );
  MUX21X1_HVT U24 ( .A1(conv2_sram_rdata_weight[7]), .A2(
        conv1_sram_rdata_weight[7]), .S0(n392), .Y(conv_weight_box[7]) );
  MUX21X1_HVT U25 ( .A1(conv2_sram_rdata_weight[63]), .A2(
        conv1_sram_rdata_weight[63]), .S0(n397), .Y(conv_weight_box[63]) );
  NOR2X0_HVT U26 ( .A1(DP_OP_425J2_127_3477_n2791), .A2(
        DP_OP_424J2_126_3477_n2051), .Y(DP_OP_423J2_125_3477_n2035) );
  NOR2X0_HVT U27 ( .A1(DP_OP_425J2_127_3477_n2790), .A2(
        DP_OP_424J2_126_3477_n2051), .Y(DP_OP_423J2_125_3477_n2034) );
  NOR2X0_HVT U28 ( .A1(DP_OP_422J2_124_3477_n2441), .A2(
        DP_OP_422J2_124_3477_n2445), .Y(DP_OP_422J2_124_3477_n2417) );
  NOR2X0_HVT U29 ( .A1(DP_OP_422J2_124_3477_n2439), .A2(
        DP_OP_422J2_124_3477_n2445), .Y(DP_OP_422J2_124_3477_n2415) );
  INVX1_HVT U30 ( .A(conv_weight_box[7]), .Y(DP_OP_422J2_124_3477_n1960) );
  OR2X1_HVT U31 ( .A1(DP_OP_422J2_124_3477_n2436), .A2(
        DP_OP_422J2_124_3477_n2445), .Y(DP_OP_422J2_124_3477_n2412) );
  NOR2X0_HVT U32 ( .A1(DP_OP_422J2_124_3477_n3009), .A2(
        DP_OP_424J2_126_3477_n2051), .Y(DP_OP_424J2_126_3477_n2035) );
  OR2X1_HVT U33 ( .A1(DP_OP_423J2_125_3477_n2707), .A2(
        DP_OP_424J2_126_3477_n2620), .Y(DP_OP_424J2_126_3477_n2587) );
  NOR2X0_HVT U34 ( .A1(DP_OP_422J2_124_3477_n3008), .A2(
        DP_OP_424J2_126_3477_n2051), .Y(DP_OP_424J2_126_3477_n2034) );
  MUX21X1_HVT U35 ( .A1(conv2_sram_rdata_weight[78]), .A2(
        conv1_sram_rdata_weight[78]), .S0(n399), .Y(conv_weight_box[78]) );
  INVX1_HVT U36 ( .A(tmp_big1[17]), .Y(n748) );
  INVX1_HVT U37 ( .A(tmp_big1[19]), .Y(n750) );
  INVX1_HVT U38 ( .A(tmp_big1[11]), .Y(n742) );
  MUX21X1_HVT U39 ( .A1(conv2_sum_b[17]), .A2(conv2_sum_a[17]), .S0(n412), .Y(
        tmp_big1[17]) );
  MUX21X1_HVT U40 ( .A1(conv2_sum_b[19]), .A2(conv2_sum_a[19]), .S0(n412), .Y(
        tmp_big1[19]) );
  NOR2X0_HVT U41 ( .A1(DP_OP_425J2_127_3477_n2793), .A2(
        DP_OP_424J2_126_3477_n2051), .Y(DP_OP_423J2_125_3477_n2037) );
  NOR2X0_HVT U42 ( .A1(DP_OP_423J2_125_3477_n2487), .A2(
        DP_OP_422J2_124_3477_n2445), .Y(DP_OP_422J2_124_3477_n2419) );
  NOR2X0_HVT U43 ( .A1(DP_OP_422J2_124_3477_n3011), .A2(
        DP_OP_424J2_126_3477_n2051), .Y(DP_OP_424J2_126_3477_n2037) );
  MUX21X1_HVT U44 ( .A1(tmp_big2[15]), .A2(tmp_big1[15]), .S0(n471), .Y(
        data_out[15]) );
  INVX2_HVT U45 ( .A(n381), .Y(n400) );
  NOR2X0_HVT U46 ( .A1(DP_OP_422J2_124_3477_n3012), .A2(
        DP_OP_424J2_126_3477_n2051), .Y(DP_OP_424J2_126_3477_n2038) );
  MUX21X1_HVT U47 ( .A1(conv2_sum_b[11]), .A2(conv2_sum_a[11]), .S0(n412), .Y(
        tmp_big1[11]) );
  AND2X1_HVT U48 ( .A1(n765), .A2(n381), .Y(DP_OP_425J2_127_3477_n3054) );
  INVX1_HVT U49 ( .A(DP_OP_425J2_127_3477_n3054), .Y(DP_OP_422J2_124_3477_n2)
         );
  INVX1_HVT U50 ( .A(DP_OP_425J2_127_3477_n3054), .Y(DP_OP_423J2_125_3477_n2)
         );
  INVX1_HVT U51 ( .A(DP_OP_425J2_127_3477_n3054), .Y(DP_OP_424J2_126_3477_n2)
         );
  MUX21X1_HVT U52 ( .A1(tmp_big2[5]), .A2(tmp_big1[5]), .S0(n471), .Y(
        data_out[5]) );
  MUX21X1_HVT U53 ( .A1(tmp_big2[6]), .A2(tmp_big1[6]), .S0(n471), .Y(
        data_out[6]) );
  NOR2X0_HVT U54 ( .A1(DP_OP_425J2_127_3477_n2795), .A2(
        DP_OP_424J2_126_3477_n2051), .Y(DP_OP_423J2_125_3477_n2039) );
  OAI21X1_HVT U55 ( .A1(DP_OP_422J2_124_3477_n181), .A2(
        DP_OP_422J2_124_3477_n175), .A3(DP_OP_422J2_124_3477_n176), .Y(
        DP_OP_422J2_124_3477_n174) );
  NOR2X0_HVT U56 ( .A1(DP_OP_424J2_126_3477_n2047), .A2(
        DP_OP_424J2_126_3477_n2051), .Y(DP_OP_424J2_126_3477_n2039) );
  OAI21X1_HVT U57 ( .A1(DP_OP_424J2_126_3477_n181), .A2(
        DP_OP_424J2_126_3477_n175), .A3(DP_OP_424J2_126_3477_n176), .Y(
        DP_OP_424J2_126_3477_n174) );
  AOI21X1_HVT U58 ( .A1(DP_OP_422J2_124_3477_n162), .A2(
        DP_OP_422J2_124_3477_n135), .A3(DP_OP_422J2_124_3477_n136), .Y(
        DP_OP_422J2_124_3477_n3) );
  AOI21X1_HVT U59 ( .A1(DP_OP_424J2_126_3477_n162), .A2(
        DP_OP_424J2_126_3477_n135), .A3(DP_OP_424J2_126_3477_n136), .Y(
        DP_OP_424J2_126_3477_n3) );
  INVX1_HVT U60 ( .A(n465), .Y(tmp_big1[3]) );
  XOR2X1_HVT U61 ( .A1(DP_OP_423J2_125_3477_n3), .A2(DP_OP_423J2_125_3477_n19), 
        .Y(n_conv2_sum_b[17]) );
  INVX1_HVT U62 ( .A(DP_OP_422J2_124_3477_n181), .Y(DP_OP_422J2_124_3477_n179)
         );
  XOR2X1_HVT U63 ( .A1(DP_OP_425J2_127_3477_n3), .A2(DP_OP_425J2_127_3477_n19), 
        .Y(n_conv2_sum_d[17]) );
  INVX0_HVT U64 ( .A(DP_OP_422J2_124_3477_n137), .Y(n1) );
  NAND2X0_HVT U65 ( .A1(n1), .A2(DP_OP_422J2_124_3477_n140), .Y(n2) );
  HADDX1_HVT U66 ( .A0(DP_OP_422J2_124_3477_n141), .B0(n2), .SO(
        n_conv2_sum_a[16]) );
  INVX0_HVT U67 ( .A(DP_OP_424J2_126_3477_n137), .Y(n3) );
  NAND2X0_HVT U68 ( .A1(n3), .A2(DP_OP_424J2_126_3477_n140), .Y(n4) );
  HADDX1_HVT U69 ( .A0(DP_OP_424J2_126_3477_n141), .B0(n4), .SO(
        n_conv2_sum_c[16]) );
  INVX0_HVT U70 ( .A(DP_OP_423J2_125_3477_n162), .Y(n5010) );
  OA21X1_HVT U71 ( .A1(DP_OP_423J2_125_3477_n144), .A2(n5010), .A3(
        DP_OP_423J2_125_3477_n145), .Y(DP_OP_423J2_125_3477_n141) );
  INVX0_HVT U72 ( .A(DP_OP_425J2_127_3477_n162), .Y(n6) );
  OA21X1_HVT U73 ( .A1(DP_OP_425J2_127_3477_n144), .A2(n6), .A3(
        DP_OP_425J2_127_3477_n145), .Y(DP_OP_425J2_127_3477_n141) );
  INVX0_HVT U74 ( .A(DP_OP_422J2_124_3477_n132), .Y(n7010) );
  NAND2X0_HVT U75 ( .A1(n7010), .A2(DP_OP_422J2_124_3477_n133), .Y(n8) );
  HADDX1_HVT U76 ( .A0(DP_OP_422J2_124_3477_n3), .B0(n8), .SO(
        n_conv2_sum_a[17]) );
  INVX0_HVT U77 ( .A(DP_OP_424J2_126_3477_n132), .Y(n9) );
  NAND2X0_HVT U78 ( .A1(n9), .A2(DP_OP_424J2_126_3477_n133), .Y(n10) );
  HADDX1_HVT U79 ( .A0(DP_OP_424J2_126_3477_n3), .B0(n10), .SO(
        n_conv2_sum_c[17]) );
  NAND2X0_HVT U80 ( .A1(conv2_sum_b[27]), .A2(n523), .Y(n11) );
  NAND2X0_HVT U81 ( .A1(conv2_sum_a[26]), .A2(n11), .Y(n12) );
  NAND2X0_HVT U82 ( .A1(n611), .A2(conv2_sum_a[24]), .Y(n13) );
  OA22X1_HVT U83 ( .A1(conv2_sum_b[25]), .A2(n511), .A3(conv2_sum_b[24]), .A4(
        n13), .Y(n14) );
  OA222X1_HVT U84 ( .A1(n12), .A2(conv2_sum_b[26]), .A3(conv2_sum_b[27]), .A4(
        n523), .A5(n14), .A6(n559), .Y(n555) );
  NAND2X0_HVT U85 ( .A1(DP_OP_423J2_125_3477_n237), .A2(
        DP_OP_423J2_125_3477_n152), .Y(n15) );
  HADDX1_HVT U86 ( .A0(DP_OP_423J2_125_3477_n161), .B0(n15), .SO(
        n_conv2_sum_b[14]) );
  OA21X1_HVT U87 ( .A1(DP_OP_422J2_124_3477_n132), .A2(DP_OP_422J2_124_3477_n3), .A3(DP_OP_422J2_124_3477_n133), .Y(n16) );
  NAND2X0_HVT U88 ( .A1(DP_OP_422J2_124_3477_n233), .A2(
        DP_OP_422J2_124_3477_n130), .Y(n17) );
  HADDX1_HVT U89 ( .A0(n16), .B0(n17), .SO(n_conv2_sum_a[18]) );
  NAND2X0_HVT U90 ( .A1(DP_OP_425J2_127_3477_n237), .A2(
        DP_OP_425J2_127_3477_n152), .Y(n18) );
  HADDX1_HVT U91 ( .A0(DP_OP_425J2_127_3477_n161), .B0(n18), .SO(
        n_conv2_sum_d[14]) );
  OA21X1_HVT U92 ( .A1(DP_OP_424J2_126_3477_n132), .A2(DP_OP_424J2_126_3477_n3), .A3(DP_OP_424J2_126_3477_n133), .Y(n19) );
  NAND2X0_HVT U93 ( .A1(DP_OP_424J2_126_3477_n233), .A2(
        DP_OP_424J2_126_3477_n130), .Y(n20) );
  HADDX1_HVT U94 ( .A0(n19), .B0(n20), .SO(n_conv2_sum_c[18]) );
  NAND2X0_HVT U95 ( .A1(conv2_sum_d[27]), .A2(n525), .Y(n21) );
  NAND2X0_HVT U96 ( .A1(conv2_sum_c[26]), .A2(n21), .Y(n22) );
  NAND2X0_HVT U97 ( .A1(n673), .A2(conv2_sum_c[24]), .Y(n23) );
  OA22X1_HVT U98 ( .A1(conv2_sum_d[25]), .A2(n518), .A3(conv2_sum_d[24]), .A4(
        n23), .Y(n24) );
  OA222X1_HVT U99 ( .A1(n22), .A2(conv2_sum_d[26]), .A3(conv2_sum_d[27]), .A4(
        n525), .A5(n24), .A6(n624), .Y(n620) );
  OA21X1_HVT U100 ( .A1(DP_OP_423J2_125_3477_n151), .A2(
        DP_OP_423J2_125_3477_n161), .A3(DP_OP_423J2_125_3477_n152), .Y(n25) );
  NAND2X0_HVT U101 ( .A1(DP_OP_423J2_125_3477_n236), .A2(
        DP_OP_423J2_125_3477_n149), .Y(n26) );
  HADDX1_HVT U102 ( .A0(n25), .B0(n26), .SO(n_conv2_sum_b[15]) );
  OA21X1_HVT U103 ( .A1(DP_OP_422J2_124_3477_n125), .A2(
        DP_OP_422J2_124_3477_n3), .A3(DP_OP_422J2_124_3477_n126), .Y(n27) );
  NAND2X0_HVT U104 ( .A1(n430), .A2(DP_OP_422J2_124_3477_n123), .Y(n28) );
  HADDX1_HVT U105 ( .A0(n27), .B0(n28), .SO(n_conv2_sum_a[19]) );
  OA21X1_HVT U106 ( .A1(DP_OP_425J2_127_3477_n151), .A2(
        DP_OP_425J2_127_3477_n161), .A3(DP_OP_425J2_127_3477_n152), .Y(n29) );
  NAND2X0_HVT U107 ( .A1(DP_OP_425J2_127_3477_n236), .A2(
        DP_OP_425J2_127_3477_n149), .Y(n30) );
  HADDX1_HVT U108 ( .A0(n29), .B0(n30), .SO(n_conv2_sum_d[15]) );
  OA21X1_HVT U109 ( .A1(DP_OP_424J2_126_3477_n125), .A2(
        DP_OP_424J2_126_3477_n3), .A3(DP_OP_424J2_126_3477_n126), .Y(n31) );
  NAND2X0_HVT U110 ( .A1(n452), .A2(DP_OP_424J2_126_3477_n123), .Y(n32) );
  HADDX1_HVT U111 ( .A0(n31), .B0(n32), .SO(n_conv2_sum_c[19]) );
  OA21X1_HVT U112 ( .A1(DP_OP_423J2_125_3477_n90), .A2(DP_OP_423J2_125_3477_n3), .A3(DP_OP_423J2_125_3477_n91), .Y(n33) );
  NAND2X0_HVT U113 ( .A1(DP_OP_423J2_125_3477_n227), .A2(
        DP_OP_423J2_125_3477_n88), .Y(n34) );
  HADDX1_HVT U114 ( .A0(n33), .B0(n34), .SO(n_conv2_sum_b[24]) );
  OA21X1_HVT U115 ( .A1(DP_OP_422J2_124_3477_n118), .A2(
        DP_OP_422J2_124_3477_n3), .A3(DP_OP_422J2_124_3477_n119), .Y(n35) );
  NAND2X0_HVT U116 ( .A1(DP_OP_422J2_124_3477_n231), .A2(
        DP_OP_422J2_124_3477_n116), .Y(n36) );
  HADDX1_HVT U117 ( .A0(n35), .B0(n36), .SO(n_conv2_sum_a[20]) );
  OA21X1_HVT U118 ( .A1(DP_OP_425J2_127_3477_n90), .A2(DP_OP_425J2_127_3477_n3), .A3(DP_OP_425J2_127_3477_n91), .Y(n37) );
  NAND2X0_HVT U119 ( .A1(DP_OP_425J2_127_3477_n227), .A2(
        DP_OP_425J2_127_3477_n88), .Y(n38) );
  HADDX1_HVT U120 ( .A0(n37), .B0(n38), .SO(n_conv2_sum_d[24]) );
  OA21X1_HVT U121 ( .A1(DP_OP_424J2_126_3477_n118), .A2(
        DP_OP_424J2_126_3477_n3), .A3(DP_OP_424J2_126_3477_n119), .Y(n39) );
  NAND2X0_HVT U122 ( .A1(DP_OP_424J2_126_3477_n231), .A2(
        DP_OP_424J2_126_3477_n116), .Y(n40) );
  HADDX1_HVT U123 ( .A0(n39), .B0(n40), .SO(n_conv2_sum_c[20]) );
  OA21X1_HVT U124 ( .A1(DP_OP_423J2_125_3477_n83), .A2(DP_OP_423J2_125_3477_n3), .A3(DP_OP_423J2_125_3477_n84), .Y(n41) );
  NAND2X0_HVT U125 ( .A1(n434), .A2(DP_OP_423J2_125_3477_n81), .Y(n42) );
  HADDX1_HVT U126 ( .A0(n41), .B0(n42), .SO(n_conv2_sum_b[25]) );
  OA21X1_HVT U127 ( .A1(DP_OP_422J2_124_3477_n111), .A2(
        DP_OP_422J2_124_3477_n3), .A3(DP_OP_422J2_124_3477_n112), .Y(n43) );
  NAND2X0_HVT U128 ( .A1(n429), .A2(DP_OP_422J2_124_3477_n109), .Y(n44) );
  HADDX1_HVT U129 ( .A0(n43), .B0(n44), .SO(n_conv2_sum_a[21]) );
  OA21X1_HVT U130 ( .A1(DP_OP_425J2_127_3477_n83), .A2(DP_OP_425J2_127_3477_n3), .A3(DP_OP_425J2_127_3477_n84), .Y(n45) );
  NAND2X0_HVT U131 ( .A1(n456), .A2(DP_OP_425J2_127_3477_n81), .Y(n46) );
  HADDX1_HVT U132 ( .A0(n45), .B0(n46), .SO(n_conv2_sum_d[25]) );
  OA21X1_HVT U133 ( .A1(DP_OP_424J2_126_3477_n111), .A2(
        DP_OP_424J2_126_3477_n3), .A3(DP_OP_424J2_126_3477_n112), .Y(n47) );
  NAND2X0_HVT U134 ( .A1(n451), .A2(DP_OP_424J2_126_3477_n109), .Y(n48) );
  HADDX1_HVT U135 ( .A0(n47), .B0(n48), .SO(n_conv2_sum_c[21]) );
  OA21X1_HVT U136 ( .A1(DP_OP_423J2_125_3477_n72), .A2(
        DP_OP_423J2_125_3477_n141), .A3(DP_OP_423J2_125_3477_n73), .Y(n49) );
  NAND2X0_HVT U137 ( .A1(n433), .A2(DP_OP_423J2_125_3477_n70), .Y(n5000) );
  HADDX1_HVT U138 ( .A0(n49), .B0(n5000), .SO(n_conv2_sum_b[26]) );
  OA21X1_HVT U139 ( .A1(DP_OP_422J2_124_3477_n104), .A2(
        DP_OP_422J2_124_3477_n3), .A3(DP_OP_422J2_124_3477_n105), .Y(n51) );
  NAND2X0_HVT U140 ( .A1(DP_OP_422J2_124_3477_n229), .A2(
        DP_OP_422J2_124_3477_n102), .Y(n52) );
  HADDX1_HVT U141 ( .A0(n51), .B0(n52), .SO(n_conv2_sum_a[22]) );
  OA21X1_HVT U142 ( .A1(DP_OP_425J2_127_3477_n72), .A2(
        DP_OP_425J2_127_3477_n141), .A3(DP_OP_425J2_127_3477_n73), .Y(n53) );
  NAND2X0_HVT U143 ( .A1(n455), .A2(DP_OP_425J2_127_3477_n70), .Y(n54) );
  HADDX1_HVT U144 ( .A0(n53), .B0(n54), .SO(n_conv2_sum_d[26]) );
  OA21X1_HVT U145 ( .A1(DP_OP_424J2_126_3477_n104), .A2(
        DP_OP_424J2_126_3477_n3), .A3(DP_OP_424J2_126_3477_n105), .Y(n55) );
  NAND2X0_HVT U146 ( .A1(DP_OP_424J2_126_3477_n229), .A2(
        DP_OP_424J2_126_3477_n102), .Y(n56) );
  HADDX1_HVT U147 ( .A0(n55), .B0(n56), .SO(n_conv2_sum_c[22]) );
  OA21X1_HVT U148 ( .A1(DP_OP_423J2_125_3477_n61), .A2(
        DP_OP_423J2_125_3477_n161), .A3(DP_OP_423J2_125_3477_n62), .Y(n57) );
  INVX0_HVT U149 ( .A(DP_OP_423J2_125_3477_n58), .Y(n58) );
  NAND2X0_HVT U150 ( .A1(n58), .A2(DP_OP_423J2_125_3477_n59), .Y(n59) );
  HADDX1_HVT U151 ( .A0(n57), .B0(n59), .SO(n_conv2_sum_b[27]) );
  OA21X1_HVT U152 ( .A1(DP_OP_422J2_124_3477_n97), .A2(DP_OP_422J2_124_3477_n3), .A3(DP_OP_422J2_124_3477_n98), .Y(n60) );
  NAND2X0_HVT U153 ( .A1(n425), .A2(DP_OP_422J2_124_3477_n95), .Y(n61) );
  HADDX1_HVT U154 ( .A0(n60), .B0(n61), .SO(n_conv2_sum_a[23]) );
  OA21X1_HVT U155 ( .A1(DP_OP_425J2_127_3477_n61), .A2(
        DP_OP_425J2_127_3477_n161), .A3(DP_OP_425J2_127_3477_n62), .Y(n62) );
  INVX0_HVT U156 ( .A(DP_OP_425J2_127_3477_n58), .Y(n63) );
  NAND2X0_HVT U157 ( .A1(n63), .A2(DP_OP_425J2_127_3477_n59), .Y(n64) );
  HADDX1_HVT U158 ( .A0(n62), .B0(n64), .SO(n_conv2_sum_d[27]) );
  OA21X1_HVT U159 ( .A1(DP_OP_424J2_126_3477_n97), .A2(DP_OP_424J2_126_3477_n3), .A3(DP_OP_424J2_126_3477_n98), .Y(n65) );
  NAND2X0_HVT U160 ( .A1(n447), .A2(DP_OP_424J2_126_3477_n95), .Y(n66) );
  HADDX1_HVT U161 ( .A0(n65), .B0(n66), .SO(n_conv2_sum_c[23]) );
  OA22X1_HVT U162 ( .A1(n763), .A2(tmp_big2[7]), .A3(tmp_big2[6]), .A4(n726), 
        .Y(n67) );
  AO222X1_HVT U163 ( .A1(n763), .A2(tmp_big2[7]), .A3(n762), .A4(tmp_big2[6]), 
        .A5(n727), .A6(n728), .Y(n68) );
  NAND2X0_HVT U164 ( .A1(n67), .A2(n68), .Y(n470) );
  OA21X1_HVT U165 ( .A1(DP_OP_423J2_125_3477_n118), .A2(
        DP_OP_423J2_125_3477_n3), .A3(DP_OP_423J2_125_3477_n119), .Y(n69) );
  NAND2X0_HVT U166 ( .A1(DP_OP_423J2_125_3477_n231), .A2(
        DP_OP_423J2_125_3477_n116), .Y(n7000) );
  HADDX1_HVT U167 ( .A0(n69), .B0(n7000), .SO(n_conv2_sum_b[20]) );
  OA21X1_HVT U168 ( .A1(DP_OP_422J2_124_3477_n90), .A2(DP_OP_422J2_124_3477_n3), .A3(DP_OP_422J2_124_3477_n91), .Y(n71) );
  NAND2X0_HVT U169 ( .A1(DP_OP_422J2_124_3477_n227), .A2(
        DP_OP_422J2_124_3477_n88), .Y(n72) );
  HADDX1_HVT U170 ( .A0(n71), .B0(n72), .SO(n_conv2_sum_a[24]) );
  OA21X1_HVT U171 ( .A1(DP_OP_425J2_127_3477_n118), .A2(
        DP_OP_425J2_127_3477_n3), .A3(DP_OP_425J2_127_3477_n119), .Y(n73) );
  NAND2X0_HVT U172 ( .A1(DP_OP_425J2_127_3477_n231), .A2(
        DP_OP_425J2_127_3477_n116), .Y(n74) );
  HADDX1_HVT U173 ( .A0(n73), .B0(n74), .SO(n_conv2_sum_d[20]) );
  OA21X1_HVT U174 ( .A1(DP_OP_424J2_126_3477_n90), .A2(DP_OP_424J2_126_3477_n3), .A3(DP_OP_424J2_126_3477_n91), .Y(n75) );
  NAND2X0_HVT U175 ( .A1(DP_OP_424J2_126_3477_n227), .A2(
        DP_OP_424J2_126_3477_n88), .Y(n76) );
  HADDX1_HVT U176 ( .A0(n75), .B0(n76), .SO(n_conv2_sum_c[24]) );
  OA22X1_HVT U177 ( .A1(tmp_big2[8]), .A2(n704), .A3(n547), .A4(tmp_big2[9]), 
        .Y(n77) );
  OA222X1_HVT U178 ( .A1(tmp_big2[10]), .A2(n703), .A3(tmp_big2[11]), .A4(n742), .A5(n714), .A6(n77), .Y(n708) );
  OA22X1_HVT U179 ( .A1(n661), .A2(conv2_sum_d[6]), .A3(n475), .A4(
        conv2_sum_d[7]), .Y(n78) );
  AO222X1_HVT U180 ( .A1(conv2_sum_d[6]), .A2(n487), .A3(conv2_sum_d[7]), .A4(
        n475), .A5(n663), .A6(n662), .Y(n79) );
  NAND3X0_HVT U181 ( .A1(n78), .A2(n668), .A3(n79), .Y(n541) );
  INVX0_HVT U183 ( .A(tmp_big1[28]), .Y(n81) );
  INVX0_HVT U184 ( .A(n678), .Y(n82) );
  NAND2X0_HVT U185 ( .A1(n438), .A2(DP_OP_423J2_125_3477_n216), .Y(n83) );
  AND2X1_HVT U186 ( .A1(n83), .A2(DP_OP_423J2_125_3477_n215), .Y(
        DP_OP_423J2_125_3477_n211) );
  OA21X1_HVT U187 ( .A1(DP_OP_423J2_125_3477_n111), .A2(
        DP_OP_423J2_125_3477_n3), .A3(DP_OP_423J2_125_3477_n112), .Y(n84) );
  NAND2X0_HVT U188 ( .A1(n439), .A2(DP_OP_423J2_125_3477_n109), .Y(n85) );
  HADDX1_HVT U189 ( .A0(n84), .B0(n85), .SO(n_conv2_sum_b[21]) );
  OA21X1_HVT U190 ( .A1(DP_OP_422J2_124_3477_n83), .A2(DP_OP_422J2_124_3477_n3), .A3(DP_OP_422J2_124_3477_n84), .Y(n86) );
  NAND2X0_HVT U191 ( .A1(n424), .A2(DP_OP_422J2_124_3477_n81), .Y(n87) );
  HADDX1_HVT U192 ( .A0(n86), .B0(n87), .SO(n_conv2_sum_a[25]) );
  OA21X1_HVT U193 ( .A1(DP_OP_425J2_127_3477_n111), .A2(
        DP_OP_425J2_127_3477_n3), .A3(DP_OP_425J2_127_3477_n112), .Y(n88) );
  NAND2X0_HVT U194 ( .A1(n461), .A2(DP_OP_425J2_127_3477_n109), .Y(n89) );
  HADDX1_HVT U195 ( .A0(n88), .B0(n89), .SO(n_conv2_sum_d[21]) );
  OA21X1_HVT U196 ( .A1(DP_OP_424J2_126_3477_n83), .A2(DP_OP_424J2_126_3477_n3), .A3(DP_OP_424J2_126_3477_n84), .Y(n90) );
  NAND2X0_HVT U197 ( .A1(n446), .A2(DP_OP_424J2_126_3477_n81), .Y(n91) );
  HADDX1_HVT U198 ( .A0(n90), .B0(n91), .SO(n_conv2_sum_c[25]) );
  OA22X1_HVT U199 ( .A1(n572), .A2(conv2_sum_b[8]), .A3(n549), .A4(
        conv2_sum_b[9]), .Y(n92) );
  OA222X1_HVT U200 ( .A1(conv2_sum_b[10]), .A2(n571), .A3(conv2_sum_b[11]), 
        .A4(n539), .A5(n582), .A6(n92), .Y(n576) );
  AO22X1_HVT U201 ( .A1(conv2_sum_c[9]), .A2(n417), .A3(conv2_sum_d[9]), .A4(
        N7), .Y(tmp_big2[9]) );
  OR2X1_HVT U202 ( .A1(DP_OP_423J2_125_3477_n76), .A2(
        DP_OP_423J2_125_3477_n140), .Y(n93) );
  NAND2X0_HVT U203 ( .A1(n434), .A2(DP_OP_423J2_125_3477_n86), .Y(n94) );
  NAND3X0_HVT U204 ( .A1(n93), .A2(DP_OP_423J2_125_3477_n81), .A3(n94), .Y(
        DP_OP_423J2_125_3477_n75) );
  OR2X1_HVT U205 ( .A1(DP_OP_425J2_127_3477_n76), .A2(
        DP_OP_425J2_127_3477_n140), .Y(n95) );
  NAND2X0_HVT U206 ( .A1(n456), .A2(DP_OP_425J2_127_3477_n86), .Y(n96) );
  NAND3X0_HVT U207 ( .A1(n95), .A2(DP_OP_425J2_127_3477_n81), .A3(n96), .Y(
        DP_OP_425J2_127_3477_n75) );
  NAND2X0_HVT U208 ( .A1(n428), .A2(DP_OP_422J2_124_3477_n216), .Y(n97) );
  AND2X1_HVT U209 ( .A1(n97), .A2(DP_OP_422J2_124_3477_n215), .Y(
        DP_OP_422J2_124_3477_n211) );
  NAND2X0_HVT U210 ( .A1(DP_OP_422J2_124_3477_n57), .A2(n422), .Y(n98) );
  AND2X1_HVT U211 ( .A1(n98), .A2(DP_OP_422J2_124_3477_n52), .Y(
        DP_OP_422J2_124_3477_n48) );
  NAND2X0_HVT U212 ( .A1(DP_OP_425J2_127_3477_n200), .A2(n458), .Y(n99) );
  AND2X1_HVT U213 ( .A1(n99), .A2(DP_OP_425J2_127_3477_n199), .Y(
        DP_OP_425J2_127_3477_n195) );
  NAND2X0_HVT U214 ( .A1(n450), .A2(DP_OP_424J2_126_3477_n216), .Y(n100) );
  AND2X1_HVT U215 ( .A1(n100), .A2(DP_OP_424J2_126_3477_n215), .Y(
        DP_OP_424J2_126_3477_n211) );
  NAND2X0_HVT U216 ( .A1(DP_OP_424J2_126_3477_n57), .A2(n444), .Y(n101) );
  AND2X1_HVT U217 ( .A1(n101), .A2(DP_OP_424J2_126_3477_n52), .Y(
        DP_OP_424J2_126_3477_n48) );
  INVX0_HVT U218 ( .A(DP_OP_423J2_125_3477_n209), .Y(n102) );
  NAND2X0_HVT U219 ( .A1(n102), .A2(DP_OP_423J2_125_3477_n210), .Y(n103) );
  HADDX1_HVT U220 ( .A0(DP_OP_423J2_125_3477_n211), .B0(n103), .SO(
        n_conv2_sum_b[3]) );
  OA21X1_HVT U221 ( .A1(DP_OP_423J2_125_3477_n104), .A2(
        DP_OP_423J2_125_3477_n3), .A3(DP_OP_423J2_125_3477_n105), .Y(n104) );
  NAND2X0_HVT U222 ( .A1(DP_OP_423J2_125_3477_n229), .A2(
        DP_OP_423J2_125_3477_n102), .Y(n105) );
  HADDX1_HVT U223 ( .A0(n104), .B0(n105), .SO(n_conv2_sum_b[22]) );
  OA21X1_HVT U224 ( .A1(DP_OP_422J2_124_3477_n72), .A2(
        DP_OP_422J2_124_3477_n141), .A3(DP_OP_422J2_124_3477_n73), .Y(n106) );
  NAND2X0_HVT U225 ( .A1(n423), .A2(DP_OP_422J2_124_3477_n70), .Y(n107) );
  HADDX1_HVT U226 ( .A0(n106), .B0(n107), .SO(n_conv2_sum_a[26]) );
  INVX0_HVT U227 ( .A(DP_OP_425J2_127_3477_n209), .Y(n108) );
  NAND2X0_HVT U228 ( .A1(n108), .A2(DP_OP_425J2_127_3477_n210), .Y(n109) );
  HADDX1_HVT U229 ( .A0(DP_OP_425J2_127_3477_n211), .B0(n109), .SO(
        n_conv2_sum_d[3]) );
  OA21X1_HVT U230 ( .A1(DP_OP_425J2_127_3477_n104), .A2(
        DP_OP_425J2_127_3477_n3), .A3(DP_OP_425J2_127_3477_n105), .Y(n110) );
  NAND2X0_HVT U231 ( .A1(DP_OP_425J2_127_3477_n229), .A2(
        DP_OP_425J2_127_3477_n102), .Y(n111) );
  HADDX1_HVT U232 ( .A0(n110), .B0(n111), .SO(n_conv2_sum_d[22]) );
  OA21X1_HVT U233 ( .A1(DP_OP_424J2_126_3477_n72), .A2(
        DP_OP_424J2_126_3477_n141), .A3(DP_OP_424J2_126_3477_n73), .Y(n112) );
  NAND2X0_HVT U234 ( .A1(n445), .A2(DP_OP_424J2_126_3477_n70), .Y(n113) );
  HADDX1_HVT U235 ( .A0(n112), .B0(n113), .SO(n_conv2_sum_c[26]) );
  INVX0_HVT U237 ( .A(n634), .Y(n115) );
  INVX0_HVT U239 ( .A(n551), .Y(n117) );
  INVX0_HVT U241 ( .A(n616), .Y(n119) );
  AO22X1_HVT U242 ( .A1(n471), .A2(tmp_big1[10]), .A3(n464), .A4(tmp_big2[10]), 
        .Y(data_out[10]) );
  NAND2X0_HVT U243 ( .A1(DP_OP_423J2_125_3477_n57), .A2(n432), .Y(n120) );
  AND2X1_HVT U244 ( .A1(n120), .A2(DP_OP_423J2_125_3477_n52), .Y(
        DP_OP_423J2_125_3477_n48) );
  NAND2X0_HVT U245 ( .A1(n427), .A2(DP_OP_422J2_124_3477_n208), .Y(n121) );
  AND2X1_HVT U246 ( .A1(n121), .A2(DP_OP_422J2_124_3477_n207), .Y(
        DP_OP_422J2_124_3477_n203) );
  NAND2X0_HVT U247 ( .A1(DP_OP_425J2_127_3477_n57), .A2(n454), .Y(n122) );
  AND2X1_HVT U248 ( .A1(n122), .A2(DP_OP_425J2_127_3477_n52), .Y(
        DP_OP_425J2_127_3477_n48) );
  NAND2X0_HVT U249 ( .A1(n449), .A2(DP_OP_424J2_126_3477_n208), .Y(n123) );
  AND2X1_HVT U250 ( .A1(n123), .A2(DP_OP_424J2_126_3477_n207), .Y(
        DP_OP_424J2_126_3477_n203) );
  AND2X1_HVT U251 ( .A1(DP_OP_423J2_125_3477_n207), .A2(n437), .Y(n124) );
  HADDX1_HVT U252 ( .A0(n124), .B0(DP_OP_423J2_125_3477_n208), .SO(
        n_conv2_sum_b[4]) );
  OA21X1_HVT U253 ( .A1(DP_OP_423J2_125_3477_n97), .A2(DP_OP_423J2_125_3477_n3), .A3(DP_OP_423J2_125_3477_n98), .Y(n125) );
  NAND2X0_HVT U254 ( .A1(n435), .A2(DP_OP_423J2_125_3477_n95), .Y(n126) );
  HADDX1_HVT U255 ( .A0(n125), .B0(n126), .SO(n_conv2_sum_b[23]) );
  OA21X1_HVT U256 ( .A1(DP_OP_422J2_124_3477_n61), .A2(
        DP_OP_422J2_124_3477_n161), .A3(DP_OP_422J2_124_3477_n62), .Y(n127) );
  INVX0_HVT U257 ( .A(DP_OP_422J2_124_3477_n58), .Y(n129) );
  NAND2X0_HVT U258 ( .A1(n129), .A2(DP_OP_422J2_124_3477_n59), .Y(n130) );
  HADDX1_HVT U259 ( .A0(n127), .B0(n130), .SO(n_conv2_sum_a[27]) );
  INVX0_HVT U260 ( .A(DP_OP_425J2_127_3477_n201), .Y(n131) );
  NAND2X0_HVT U261 ( .A1(n131), .A2(DP_OP_425J2_127_3477_n202), .Y(n132) );
  HADDX1_HVT U262 ( .A0(DP_OP_425J2_127_3477_n203), .B0(n132), .SO(
        n_conv2_sum_d[5]) );
  OA21X1_HVT U263 ( .A1(DP_OP_425J2_127_3477_n97), .A2(DP_OP_425J2_127_3477_n3), .A3(DP_OP_425J2_127_3477_n98), .Y(n133) );
  NAND2X0_HVT U264 ( .A1(n457), .A2(DP_OP_425J2_127_3477_n95), .Y(n134) );
  HADDX1_HVT U265 ( .A0(n133), .B0(n134), .SO(n_conv2_sum_d[23]) );
  OA21X1_HVT U266 ( .A1(DP_OP_424J2_126_3477_n61), .A2(
        DP_OP_424J2_126_3477_n161), .A3(DP_OP_424J2_126_3477_n62), .Y(n135) );
  INVX0_HVT U267 ( .A(DP_OP_424J2_126_3477_n58), .Y(n136) );
  NAND2X0_HVT U268 ( .A1(n136), .A2(DP_OP_424J2_126_3477_n59), .Y(n137) );
  HADDX1_HVT U269 ( .A0(n135), .B0(n137), .SO(n_conv2_sum_c[27]) );
  INVX0_HVT U271 ( .A(n569), .Y(n139) );
  INVX0_HVT U273 ( .A(n626), .Y(n141) );
  OR2X1_HVT U274 ( .A1(DP_OP_422J2_124_3477_n76), .A2(
        DP_OP_422J2_124_3477_n140), .Y(n142) );
  NAND2X0_HVT U275 ( .A1(n424), .A2(DP_OP_422J2_124_3477_n86), .Y(n143) );
  NAND3X0_HVT U276 ( .A1(n142), .A2(DP_OP_422J2_124_3477_n81), .A3(n143), .Y(
        DP_OP_422J2_124_3477_n75) );
  NAND2X0_HVT U277 ( .A1(n446), .A2(DP_OP_424J2_126_3477_n86), .Y(n144) );
  OR2X1_HVT U278 ( .A1(DP_OP_424J2_126_3477_n76), .A2(
        DP_OP_424J2_126_3477_n140), .Y(n145) );
  NAND3X0_HVT U279 ( .A1(n145), .A2(DP_OP_424J2_126_3477_n81), .A3(n144), .Y(
        DP_OP_424J2_126_3477_n75) );
  AOI22X1_HVT U281 ( .A1(n433), .A2(DP_OP_423J2_125_3477_n75), .A3(
        DP_OP_423J2_125_3477_n158), .A4(DP_OP_423J2_125_3477_n63), .Y(n147) );
  NAND2X0_HVT U282 ( .A1(DP_OP_422J2_124_3477_n200), .A2(n426), .Y(n148) );
  AND2X1_HVT U283 ( .A1(n148), .A2(DP_OP_422J2_124_3477_n199), .Y(
        DP_OP_422J2_124_3477_n195) );
  AOI22X1_HVT U285 ( .A1(n455), .A2(DP_OP_425J2_127_3477_n75), .A3(
        DP_OP_425J2_127_3477_n158), .A4(DP_OP_425J2_127_3477_n63), .Y(n150) );
  NAND2X0_HVT U286 ( .A1(DP_OP_424J2_126_3477_n200), .A2(n448), .Y(n151) );
  AND2X1_HVT U287 ( .A1(n151), .A2(DP_OP_424J2_126_3477_n199), .Y(
        DP_OP_424J2_126_3477_n195) );
  INVX0_HVT U288 ( .A(DP_OP_423J2_125_3477_n201), .Y(n152) );
  NAND2X0_HVT U289 ( .A1(n152), .A2(DP_OP_423J2_125_3477_n202), .Y(n153) );
  HADDX1_HVT U290 ( .A0(DP_OP_423J2_125_3477_n203), .B0(n153), .SO(
        n_conv2_sum_b[5]) );
  INVX0_HVT U291 ( .A(DP_OP_423J2_125_3477_n193), .Y(n154) );
  NAND2X0_HVT U292 ( .A1(n154), .A2(DP_OP_423J2_125_3477_n194), .Y(n155) );
  HADDX1_HVT U293 ( .A0(DP_OP_423J2_125_3477_n195), .B0(n155), .SO(
        n_conv2_sum_b[7]) );
  AND2X1_HVT U294 ( .A1(DP_OP_423J2_125_3477_n241), .A2(
        DP_OP_423J2_125_3477_n181), .Y(n156) );
  HADDX1_HVT U295 ( .A0(n156), .B0(DP_OP_423J2_125_3477_n182), .SO(
        n_conv2_sum_b[10]) );
  INVX0_HVT U296 ( .A(DP_OP_423J2_125_3477_n39), .Y(n157) );
  NAND2X0_HVT U297 ( .A1(n157), .A2(DP_OP_423J2_125_3477_n40), .Y(n158) );
  HADDX1_HVT U298 ( .A0(DP_OP_423J2_125_3477_n41), .B0(n158), .SO(
        n_conv2_sum_b[30]) );
  INVX0_HVT U299 ( .A(DP_OP_422J2_124_3477_n56), .Y(n159) );
  OA21X1_HVT U300 ( .A1(DP_OP_422J2_124_3477_n161), .A2(n159), .A3(
        DP_OP_422J2_124_3477_n55), .Y(n160) );
  NAND2X0_HVT U301 ( .A1(n422), .A2(DP_OP_422J2_124_3477_n52), .Y(n161) );
  HADDX1_HVT U302 ( .A0(n160), .B0(n161), .SO(n_conv2_sum_a[28]) );
  AND2X1_HVT U303 ( .A1(DP_OP_425J2_127_3477_n207), .A2(n459), .Y(n162) );
  HADDX1_HVT U304 ( .A0(n162), .B0(DP_OP_425J2_127_3477_n208), .SO(
        n_conv2_sum_d[4]) );
  AND2X1_HVT U305 ( .A1(DP_OP_425J2_127_3477_n199), .A2(n458), .Y(n163) );
  HADDX1_HVT U306 ( .A0(n163), .B0(DP_OP_425J2_127_3477_n200), .SO(
        n_conv2_sum_d[6]) );
  INVX0_HVT U307 ( .A(DP_OP_425J2_127_3477_n189), .Y(n164) );
  NAND2X0_HVT U308 ( .A1(n164), .A2(DP_OP_425J2_127_3477_n190), .Y(n165) );
  HADDX1_HVT U309 ( .A0(DP_OP_425J2_127_3477_n191), .B0(n165), .SO(
        n_conv2_sum_d[8]) );
  INVX0_HVT U310 ( .A(DP_OP_425J2_127_3477_n39), .Y(n166) );
  NAND2X0_HVT U311 ( .A1(n166), .A2(DP_OP_425J2_127_3477_n40), .Y(n167) );
  HADDX1_HVT U312 ( .A0(DP_OP_425J2_127_3477_n41), .B0(n167), .SO(
        n_conv2_sum_d[30]) );
  INVX0_HVT U313 ( .A(DP_OP_424J2_126_3477_n56), .Y(n168) );
  OA21X1_HVT U314 ( .A1(DP_OP_424J2_126_3477_n161), .A2(n168), .A3(
        DP_OP_424J2_126_3477_n55), .Y(n169) );
  NAND2X0_HVT U315 ( .A1(n444), .A2(DP_OP_424J2_126_3477_n52), .Y(n170) );
  HADDX1_HVT U316 ( .A0(n169), .B0(n170), .SO(n_conv2_sum_c[28]) );
  INVX0_HVT U317 ( .A(tmp_big1[20]), .Y(n171) );
  INVX0_HVT U318 ( .A(n689), .Y(n172) );
  NAND2X0_HVT U320 ( .A1(DP_OP_422J2_124_3477_n158), .A2(
        DP_OP_422J2_124_3477_n236), .Y(n174) );
  AND2X1_HVT U321 ( .A1(n174), .A2(DP_OP_422J2_124_3477_n149), .Y(
        DP_OP_422J2_124_3477_n145) );
  NAND2X0_HVT U322 ( .A1(DP_OP_424J2_126_3477_n158), .A2(
        DP_OP_424J2_126_3477_n236), .Y(n175) );
  AND2X1_HVT U323 ( .A1(n175), .A2(DP_OP_424J2_126_3477_n149), .Y(
        DP_OP_424J2_126_3477_n145) );
  NAND2X0_HVT U324 ( .A1(n437), .A2(DP_OP_423J2_125_3477_n208), .Y(n176) );
  AND2X1_HVT U325 ( .A1(n176), .A2(DP_OP_423J2_125_3477_n207), .Y(
        DP_OP_423J2_125_3477_n203) );
  NAND2X0_HVT U326 ( .A1(DP_OP_423J2_125_3477_n128), .A2(n440), .Y(n177) );
  AND2X1_HVT U327 ( .A1(n177), .A2(DP_OP_423J2_125_3477_n123), .Y(
        DP_OP_423J2_125_3477_n119) );
  NAND2X0_HVT U328 ( .A1(DP_OP_422J2_124_3477_n100), .A2(n425), .Y(n178) );
  AND2X1_HVT U329 ( .A1(n178), .A2(DP_OP_422J2_124_3477_n95), .Y(
        DP_OP_422J2_124_3477_n91) );
  NAND2X0_HVT U330 ( .A1(n460), .A2(DP_OP_425J2_127_3477_n216), .Y(n179) );
  AND2X1_HVT U331 ( .A1(n179), .A2(DP_OP_425J2_127_3477_n215), .Y(
        DP_OP_425J2_127_3477_n211) );
  NAND2X0_HVT U332 ( .A1(DP_OP_425J2_127_3477_n128), .A2(n462), .Y(n180) );
  AND2X1_HVT U333 ( .A1(n180), .A2(DP_OP_425J2_127_3477_n123), .Y(
        DP_OP_425J2_127_3477_n119) );
  NAND2X0_HVT U334 ( .A1(DP_OP_424J2_126_3477_n100), .A2(n447), .Y(n181) );
  AND2X1_HVT U335 ( .A1(n181), .A2(DP_OP_424J2_126_3477_n95), .Y(
        DP_OP_424J2_126_3477_n91) );
  INVX0_HVT U336 ( .A(DP_OP_423J2_125_3477_n189), .Y(n182) );
  NAND2X0_HVT U337 ( .A1(n182), .A2(DP_OP_423J2_125_3477_n190), .Y(n183) );
  HADDX1_HVT U338 ( .A0(DP_OP_423J2_125_3477_n191), .B0(n183), .SO(
        n_conv2_sum_b[8]) );
  INVX0_HVT U339 ( .A(DP_OP_423J2_125_3477_n170), .Y(n184) );
  NAND2X0_HVT U340 ( .A1(n184), .A2(DP_OP_423J2_125_3477_n171), .Y(n185) );
  HADDX1_HVT U341 ( .A0(DP_OP_423J2_125_3477_n172), .B0(n185), .SO(
        n_conv2_sum_b[12]) );
  OA21X1_HVT U342 ( .A1(DP_OP_423J2_125_3477_n39), .A2(
        DP_OP_423J2_125_3477_n41), .A3(DP_OP_423J2_125_3477_n40), .Y(n186) );
  NAND2X0_HVT U343 ( .A1(n431), .A2(DP_OP_423J2_125_3477_n37), .Y(n187) );
  HADDX1_HVT U344 ( .A0(n186), .B0(n187), .SO(n_conv2_sum_b[31]) );
  INVX0_HVT U345 ( .A(DP_OP_422J2_124_3477_n209), .Y(n188) );
  NAND2X0_HVT U346 ( .A1(n188), .A2(DP_OP_422J2_124_3477_n210), .Y(n189) );
  HADDX1_HVT U347 ( .A0(DP_OP_422J2_124_3477_n211), .B0(n189), .SO(
        n_conv2_sum_a[3]) );
  INVX0_HVT U348 ( .A(DP_OP_422J2_124_3477_n193), .Y(n190) );
  NAND2X0_HVT U349 ( .A1(n190), .A2(DP_OP_422J2_124_3477_n194), .Y(n191) );
  HADDX1_HVT U350 ( .A0(DP_OP_422J2_124_3477_n195), .B0(n191), .SO(
        n_conv2_sum_a[7]) );
  AND2X1_HVT U351 ( .A1(DP_OP_422J2_124_3477_n241), .A2(
        DP_OP_422J2_124_3477_n181), .Y(n192) );
  HADDX1_HVT U352 ( .A0(n192), .B0(DP_OP_422J2_124_3477_n182), .SO(
        n_conv2_sum_a[10]) );
  OA21X1_HVT U353 ( .A1(DP_OP_422J2_124_3477_n47), .A2(
        DP_OP_422J2_124_3477_n161), .A3(DP_OP_422J2_124_3477_n48), .Y(n193) );
  INVX0_HVT U354 ( .A(DP_OP_422J2_124_3477_n44), .Y(n194) );
  NAND2X0_HVT U355 ( .A1(n194), .A2(DP_OP_422J2_124_3477_n45), .Y(n195) );
  HADDX1_HVT U356 ( .A0(n193), .B0(n195), .SO(n_conv2_sum_a[29]) );
  OA21X1_HVT U357 ( .A1(DP_OP_425J2_127_3477_n189), .A2(
        DP_OP_425J2_127_3477_n191), .A3(DP_OP_425J2_127_3477_n190), .Y(n196)
         );
  INVX0_HVT U358 ( .A(DP_OP_425J2_127_3477_n186), .Y(n197) );
  NAND2X0_HVT U359 ( .A1(n197), .A2(DP_OP_425J2_127_3477_n187), .Y(n198) );
  HADDX1_HVT U360 ( .A0(n196), .B0(n198), .SO(n_conv2_sum_d[9]) );
  INVX0_HVT U361 ( .A(DP_OP_425J2_127_3477_n170), .Y(n199) );
  NAND2X0_HVT U362 ( .A1(n199), .A2(DP_OP_425J2_127_3477_n171), .Y(n200) );
  HADDX1_HVT U363 ( .A0(DP_OP_425J2_127_3477_n172), .B0(n200), .SO(
        n_conv2_sum_d[12]) );
  OA21X1_HVT U364 ( .A1(DP_OP_425J2_127_3477_n39), .A2(
        DP_OP_425J2_127_3477_n41), .A3(DP_OP_425J2_127_3477_n40), .Y(n201) );
  NAND2X0_HVT U365 ( .A1(n453), .A2(DP_OP_425J2_127_3477_n37), .Y(n202) );
  HADDX1_HVT U366 ( .A0(n201), .B0(n202), .SO(n_conv2_sum_d[31]) );
  INVX0_HVT U367 ( .A(DP_OP_424J2_126_3477_n209), .Y(n203) );
  NAND2X0_HVT U368 ( .A1(n203), .A2(DP_OP_424J2_126_3477_n210), .Y(n204) );
  HADDX1_HVT U369 ( .A0(DP_OP_424J2_126_3477_n211), .B0(n204), .SO(
        n_conv2_sum_c[3]) );
  INVX0_HVT U370 ( .A(DP_OP_424J2_126_3477_n193), .Y(n205) );
  NAND2X0_HVT U371 ( .A1(n205), .A2(DP_OP_424J2_126_3477_n194), .Y(n206) );
  HADDX1_HVT U372 ( .A0(DP_OP_424J2_126_3477_n195), .B0(n206), .SO(
        n_conv2_sum_c[7]) );
  OA21X1_HVT U373 ( .A1(DP_OP_424J2_126_3477_n47), .A2(
        DP_OP_424J2_126_3477_n161), .A3(DP_OP_424J2_126_3477_n48), .Y(n207) );
  INVX0_HVT U374 ( .A(DP_OP_424J2_126_3477_n44), .Y(n208) );
  NAND2X0_HVT U375 ( .A1(n208), .A2(DP_OP_424J2_126_3477_n45), .Y(n209) );
  HADDX1_HVT U376 ( .A0(n207), .B0(n209), .SO(n_conv2_sum_c[29]) );
  NAND2X0_HVT U377 ( .A1(conv2_sum_b[19]), .A2(n508), .Y(n210) );
  NAND2X0_HVT U378 ( .A1(conv2_sum_a[18]), .A2(n210), .Y(n211) );
  NAND2X0_HVT U379 ( .A1(n599), .A2(conv2_sum_a[16]), .Y(n212) );
  OA22X1_HVT U380 ( .A1(conv2_sum_b[17]), .A2(n507), .A3(conv2_sum_b[16]), 
        .A4(n212), .Y(n213) );
  OA222X1_HVT U381 ( .A1(n211), .A2(conv2_sum_b[18]), .A3(conv2_sum_b[19]), 
        .A4(n508), .A5(n213), .A6(n602), .Y(n565) );
  NOR2X0_HVT U382 ( .A1(n666), .A2(n665), .Y(n214) );
  INVX0_HVT U384 ( .A(tmp_big1[24]), .Y(n216) );
  NAND2X0_HVT U385 ( .A1(tmp_big2[24]), .A2(n216), .Y(n217) );
  INVX0_HVT U386 ( .A(n687), .Y(n218) );
  INVX0_HVT U387 ( .A(n686), .Y(n219) );
  AND4X1_HVT U388 ( .A1(n736), .A2(n217), .A3(n218), .A4(n219), .Y(n534) );
  NAND2X0_HVT U389 ( .A1(DP_OP_423J2_125_3477_n114), .A2(n439), .Y(n220) );
  AND2X1_HVT U390 ( .A1(n220), .A2(DP_OP_423J2_125_3477_n109), .Y(
        DP_OP_423J2_125_3477_n105) );
  NAND2X0_HVT U391 ( .A1(DP_OP_422J2_124_3477_n128), .A2(n430), .Y(n221) );
  AND2X1_HVT U392 ( .A1(n221), .A2(DP_OP_422J2_124_3477_n123), .Y(
        DP_OP_422J2_124_3477_n119) );
  AOI22X1_HVT U394 ( .A1(n423), .A2(DP_OP_422J2_124_3477_n75), .A3(
        DP_OP_422J2_124_3477_n158), .A4(DP_OP_422J2_124_3477_n63), .Y(n223) );
  NAND2X0_HVT U395 ( .A1(DP_OP_425J2_127_3477_n114), .A2(n461), .Y(n224) );
  AND2X1_HVT U396 ( .A1(n224), .A2(DP_OP_425J2_127_3477_n109), .Y(
        DP_OP_425J2_127_3477_n105) );
  NAND2X0_HVT U397 ( .A1(DP_OP_424J2_126_3477_n128), .A2(n452), .Y(n225) );
  AND2X1_HVT U398 ( .A1(n225), .A2(DP_OP_424J2_126_3477_n123), .Y(
        DP_OP_424J2_126_3477_n119) );
  AOI22X1_HVT U399 ( .A1(n445), .A2(DP_OP_424J2_126_3477_n75), .A3(
        DP_OP_424J2_126_3477_n158), .A4(DP_OP_424J2_126_3477_n63), .Y(n226) );
  INVX0_HVT U401 ( .A(DP_OP_423J2_125_3477_n217), .Y(n228) );
  AND2X1_HVT U402 ( .A1(n228), .A2(DP_OP_423J2_125_3477_n218), .Y(n229) );
  HADDX1_HVT U403 ( .A0(n229), .B0(DP_OP_423J2_125_3477_n219), .SO(
        n_conv2_sum_b[1]) );
  AND2X1_HVT U404 ( .A1(DP_OP_423J2_125_3477_n199), .A2(n436), .Y(n230) );
  HADDX1_HVT U405 ( .A0(n230), .B0(DP_OP_423J2_125_3477_n200), .SO(
        n_conv2_sum_b[6]) );
  OA21X1_HVT U406 ( .A1(DP_OP_423J2_125_3477_n189), .A2(
        DP_OP_423J2_125_3477_n191), .A3(DP_OP_423J2_125_3477_n190), .Y(n231)
         );
  INVX0_HVT U407 ( .A(DP_OP_423J2_125_3477_n186), .Y(n232) );
  NAND2X0_HVT U408 ( .A1(n232), .A2(DP_OP_423J2_125_3477_n187), .Y(n233) );
  HADDX1_HVT U409 ( .A0(n231), .B0(n233), .SO(n_conv2_sum_b[9]) );
  OA21X1_HVT U410 ( .A1(DP_OP_423J2_125_3477_n170), .A2(
        DP_OP_423J2_125_3477_n172), .A3(DP_OP_423J2_125_3477_n171), .Y(n234)
         );
  INVX0_HVT U411 ( .A(DP_OP_423J2_125_3477_n167), .Y(n235) );
  NAND2X0_HVT U412 ( .A1(n235), .A2(DP_OP_423J2_125_3477_n168), .Y(n236) );
  HADDX1_HVT U413 ( .A0(n234), .B0(n236), .SO(n_conv2_sum_b[13]) );
  INVX0_HVT U414 ( .A(DP_OP_423J2_125_3477_n56), .Y(n237) );
  OA21X1_HVT U415 ( .A1(DP_OP_423J2_125_3477_n161), .A2(n237), .A3(
        DP_OP_423J2_125_3477_n55), .Y(n238) );
  NAND2X0_HVT U416 ( .A1(n432), .A2(DP_OP_423J2_125_3477_n52), .Y(n239) );
  HADDX1_HVT U417 ( .A0(n238), .B0(n239), .SO(n_conv2_sum_b[28]) );
  INVX0_HVT U418 ( .A(DP_OP_422J2_124_3477_n217), .Y(n240) );
  AND2X1_HVT U419 ( .A1(n240), .A2(DP_OP_422J2_124_3477_n218), .Y(n241) );
  HADDX1_HVT U420 ( .A0(n241), .B0(DP_OP_422J2_124_3477_n219), .SO(
        n_conv2_sum_a[1]) );
  INVX0_HVT U421 ( .A(DP_OP_422J2_124_3477_n201), .Y(n242) );
  NAND2X0_HVT U422 ( .A1(n242), .A2(DP_OP_422J2_124_3477_n202), .Y(n243) );
  HADDX1_HVT U423 ( .A0(DP_OP_422J2_124_3477_n203), .B0(n243), .SO(
        n_conv2_sum_a[5]) );
  INVX0_HVT U424 ( .A(DP_OP_422J2_124_3477_n189), .Y(n244) );
  NAND2X0_HVT U425 ( .A1(n244), .A2(DP_OP_422J2_124_3477_n190), .Y(n245) );
  HADDX1_HVT U426 ( .A0(DP_OP_422J2_124_3477_n191), .B0(n245), .SO(
        n_conv2_sum_a[8]) );
  INVX0_HVT U427 ( .A(DP_OP_422J2_124_3477_n170), .Y(n246) );
  NAND2X0_HVT U428 ( .A1(n246), .A2(DP_OP_422J2_124_3477_n171), .Y(n247) );
  HADDX1_HVT U429 ( .A0(DP_OP_422J2_124_3477_n172), .B0(n247), .SO(
        n_conv2_sum_a[12]) );
  INVX0_HVT U430 ( .A(DP_OP_422J2_124_3477_n39), .Y(n248) );
  NAND2X0_HVT U431 ( .A1(n248), .A2(DP_OP_422J2_124_3477_n40), .Y(n249) );
  HADDX1_HVT U432 ( .A0(DP_OP_422J2_124_3477_n41), .B0(n249), .SO(
        n_conv2_sum_a[30]) );
  INVX0_HVT U433 ( .A(DP_OP_425J2_127_3477_n217), .Y(n250) );
  AND2X1_HVT U434 ( .A1(n250), .A2(DP_OP_425J2_127_3477_n218), .Y(n251) );
  HADDX1_HVT U435 ( .A0(n251), .B0(DP_OP_425J2_127_3477_n219), .SO(
        n_conv2_sum_d[1]) );
  INVX0_HVT U436 ( .A(DP_OP_425J2_127_3477_n193), .Y(n252) );
  NAND2X0_HVT U437 ( .A1(n252), .A2(DP_OP_425J2_127_3477_n194), .Y(n253) );
  HADDX1_HVT U438 ( .A0(DP_OP_425J2_127_3477_n195), .B0(n253), .SO(
        n_conv2_sum_d[7]) );
  OA21X1_HVT U439 ( .A1(DP_OP_425J2_127_3477_n170), .A2(
        DP_OP_425J2_127_3477_n172), .A3(DP_OP_425J2_127_3477_n171), .Y(n254)
         );
  INVX0_HVT U440 ( .A(DP_OP_425J2_127_3477_n167), .Y(n255) );
  NAND2X0_HVT U441 ( .A1(n255), .A2(DP_OP_425J2_127_3477_n168), .Y(n256) );
  HADDX1_HVT U442 ( .A0(n254), .B0(n256), .SO(n_conv2_sum_d[13]) );
  INVX0_HVT U443 ( .A(DP_OP_425J2_127_3477_n56), .Y(n257) );
  OA21X1_HVT U444 ( .A1(DP_OP_425J2_127_3477_n161), .A2(n257), .A3(
        DP_OP_425J2_127_3477_n55), .Y(n258) );
  NAND2X0_HVT U445 ( .A1(n454), .A2(DP_OP_425J2_127_3477_n52), .Y(n259) );
  HADDX1_HVT U446 ( .A0(n258), .B0(n259), .SO(n_conv2_sum_d[28]) );
  INVX0_HVT U447 ( .A(DP_OP_424J2_126_3477_n217), .Y(n260) );
  AND2X1_HVT U448 ( .A1(n260), .A2(DP_OP_424J2_126_3477_n218), .Y(n261) );
  HADDX1_HVT U449 ( .A0(n261), .B0(DP_OP_424J2_126_3477_n219), .SO(
        n_conv2_sum_c[1]) );
  INVX0_HVT U450 ( .A(DP_OP_424J2_126_3477_n201), .Y(n262) );
  NAND2X0_HVT U451 ( .A1(n262), .A2(DP_OP_424J2_126_3477_n202), .Y(n263) );
  HADDX1_HVT U452 ( .A0(DP_OP_424J2_126_3477_n203), .B0(n263), .SO(
        n_conv2_sum_c[5]) );
  INVX0_HVT U453 ( .A(DP_OP_424J2_126_3477_n189), .Y(n264) );
  NAND2X0_HVT U454 ( .A1(n264), .A2(DP_OP_424J2_126_3477_n190), .Y(n265) );
  HADDX1_HVT U455 ( .A0(DP_OP_424J2_126_3477_n191), .B0(n265), .SO(
        n_conv2_sum_c[8]) );
  INVX0_HVT U456 ( .A(DP_OP_424J2_126_3477_n170), .Y(n266) );
  NAND2X0_HVT U457 ( .A1(n266), .A2(DP_OP_424J2_126_3477_n171), .Y(n267) );
  HADDX1_HVT U458 ( .A0(DP_OP_424J2_126_3477_n172), .B0(n267), .SO(
        n_conv2_sum_c[12]) );
  INVX0_HVT U459 ( .A(DP_OP_424J2_126_3477_n39), .Y(n268) );
  NAND2X0_HVT U460 ( .A1(n268), .A2(DP_OP_424J2_126_3477_n40), .Y(n269) );
  HADDX1_HVT U461 ( .A0(DP_OP_424J2_126_3477_n41), .B0(n269), .SO(
        n_conv2_sum_c[30]) );
  INVX0_HVT U462 ( .A(n561), .Y(n270) );
  NAND2X0_HVT U464 ( .A1(conv2_sum_d[19]), .A2(n515), .Y(n272) );
  NAND2X0_HVT U465 ( .A1(conv2_sum_c[18]), .A2(n272), .Y(n273) );
  NAND2X0_HVT U466 ( .A1(n664), .A2(conv2_sum_c[16]), .Y(n274) );
  OA22X1_HVT U467 ( .A1(conv2_sum_d[17]), .A2(n514), .A3(conv2_sum_d[16]), 
        .A4(n274), .Y(n275) );
  OA222X1_HVT U468 ( .A1(n273), .A2(conv2_sum_d[18]), .A3(conv2_sum_d[19]), 
        .A4(n515), .A5(n275), .A6(n666), .Y(n630) );
  NAND2X0_HVT U469 ( .A1(n679), .A2(tmp_big1[26]), .Y(n276) );
  NAND2X0_HVT U470 ( .A1(n736), .A2(tmp_big1[24]), .Y(n277) );
  OA22X1_HVT U471 ( .A1(tmp_big2[25]), .A2(n754), .A3(tmp_big2[24]), .A4(n277), 
        .Y(n278) );
  OA222X1_HVT U472 ( .A1(n276), .A2(tmp_big2[26]), .A3(tmp_big2[27]), .A4(n756), .A5(n687), .A6(n278), .Y(n683) );
  NAND2X0_HVT U473 ( .A1(DP_OP_423J2_125_3477_n158), .A2(
        DP_OP_423J2_125_3477_n236), .Y(n279) );
  AND2X1_HVT U474 ( .A1(n279), .A2(DP_OP_423J2_125_3477_n149), .Y(
        DP_OP_423J2_125_3477_n145) );
  NAND2X0_HVT U475 ( .A1(DP_OP_425J2_127_3477_n158), .A2(
        DP_OP_425J2_127_3477_n236), .Y(n280) );
  AND2X1_HVT U476 ( .A1(n280), .A2(DP_OP_425J2_127_3477_n149), .Y(
        DP_OP_425J2_127_3477_n145) );
  NAND2X0_HVT U477 ( .A1(DP_OP_423J2_125_3477_n200), .A2(n436), .Y(n281) );
  AND2X1_HVT U478 ( .A1(n281), .A2(DP_OP_423J2_125_3477_n199), .Y(
        DP_OP_423J2_125_3477_n195) );
  NAND2X0_HVT U479 ( .A1(DP_OP_423J2_125_3477_n100), .A2(n435), .Y(n282) );
  AND2X1_HVT U480 ( .A1(n282), .A2(DP_OP_423J2_125_3477_n95), .Y(
        DP_OP_423J2_125_3477_n91) );
  NAND2X0_HVT U481 ( .A1(DP_OP_422J2_124_3477_n114), .A2(n429), .Y(n283) );
  AND2X1_HVT U482 ( .A1(n283), .A2(DP_OP_422J2_124_3477_n109), .Y(
        DP_OP_422J2_124_3477_n105) );
  NAND2X0_HVT U483 ( .A1(n459), .A2(DP_OP_425J2_127_3477_n208), .Y(n284) );
  AND2X1_HVT U484 ( .A1(n284), .A2(DP_OP_425J2_127_3477_n207), .Y(
        DP_OP_425J2_127_3477_n203) );
  NAND2X0_HVT U485 ( .A1(DP_OP_425J2_127_3477_n100), .A2(n457), .Y(n285) );
  AND2X1_HVT U486 ( .A1(n285), .A2(DP_OP_425J2_127_3477_n95), .Y(
        DP_OP_425J2_127_3477_n91) );
  NAND2X0_HVT U487 ( .A1(DP_OP_424J2_126_3477_n114), .A2(n451), .Y(n286) );
  AND2X1_HVT U488 ( .A1(n286), .A2(DP_OP_424J2_126_3477_n109), .Y(
        DP_OP_424J2_126_3477_n105) );
  AND2X1_HVT U489 ( .A1(DP_OP_423J2_125_3477_n215), .A2(n438), .Y(n287) );
  HADDX1_HVT U490 ( .A0(n287), .B0(DP_OP_423J2_125_3477_n216), .SO(
        n_conv2_sum_b[2]) );
  OA21X1_HVT U491 ( .A1(DP_OP_423J2_125_3477_n47), .A2(
        DP_OP_423J2_125_3477_n161), .A3(DP_OP_423J2_125_3477_n48), .Y(n288) );
  INVX0_HVT U492 ( .A(DP_OP_423J2_125_3477_n44), .Y(n289) );
  NAND2X0_HVT U493 ( .A1(n289), .A2(DP_OP_423J2_125_3477_n45), .Y(n290) );
  HADDX1_HVT U494 ( .A0(n288), .B0(n290), .SO(n_conv2_sum_b[29]) );
  AND2X1_HVT U495 ( .A1(DP_OP_422J2_124_3477_n215), .A2(n428), .Y(n291) );
  HADDX1_HVT U496 ( .A0(n291), .B0(DP_OP_422J2_124_3477_n216), .SO(
        n_conv2_sum_a[2]) );
  AND2X1_HVT U497 ( .A1(DP_OP_422J2_124_3477_n207), .A2(n427), .Y(n292) );
  HADDX1_HVT U498 ( .A0(n292), .B0(DP_OP_422J2_124_3477_n208), .SO(
        n_conv2_sum_a[4]) );
  AND2X1_HVT U499 ( .A1(DP_OP_422J2_124_3477_n199), .A2(n426), .Y(n293) );
  HADDX1_HVT U500 ( .A0(n293), .B0(DP_OP_422J2_124_3477_n200), .SO(
        n_conv2_sum_a[6]) );
  OA21X1_HVT U501 ( .A1(DP_OP_422J2_124_3477_n189), .A2(
        DP_OP_422J2_124_3477_n191), .A3(DP_OP_422J2_124_3477_n190), .Y(n294)
         );
  INVX0_HVT U502 ( .A(DP_OP_422J2_124_3477_n186), .Y(n295) );
  NAND2X0_HVT U503 ( .A1(n295), .A2(DP_OP_422J2_124_3477_n187), .Y(n296) );
  HADDX1_HVT U504 ( .A0(n294), .B0(n296), .SO(n_conv2_sum_a[9]) );
  OA21X1_HVT U505 ( .A1(DP_OP_422J2_124_3477_n170), .A2(
        DP_OP_422J2_124_3477_n172), .A3(DP_OP_422J2_124_3477_n171), .Y(n297)
         );
  INVX0_HVT U506 ( .A(DP_OP_422J2_124_3477_n167), .Y(n298) );
  NAND2X0_HVT U507 ( .A1(n298), .A2(DP_OP_422J2_124_3477_n168), .Y(n299) );
  HADDX1_HVT U508 ( .A0(n297), .B0(n299), .SO(n_conv2_sum_a[13]) );
  OA21X1_HVT U509 ( .A1(DP_OP_422J2_124_3477_n39), .A2(
        DP_OP_422J2_124_3477_n41), .A3(DP_OP_422J2_124_3477_n40), .Y(n300) );
  NAND2X0_HVT U510 ( .A1(n420), .A2(DP_OP_422J2_124_3477_n37), .Y(n301) );
  HADDX1_HVT U511 ( .A0(n300), .B0(n301), .SO(n_conv2_sum_a[31]) );
  AND2X1_HVT U512 ( .A1(DP_OP_425J2_127_3477_n215), .A2(n460), .Y(n302) );
  HADDX1_HVT U513 ( .A0(n302), .B0(DP_OP_425J2_127_3477_n216), .SO(
        n_conv2_sum_d[2]) );
  AND2X1_HVT U514 ( .A1(DP_OP_425J2_127_3477_n241), .A2(
        DP_OP_425J2_127_3477_n181), .Y(n303) );
  HADDX1_HVT U515 ( .A0(n303), .B0(DP_OP_425J2_127_3477_n182), .SO(
        n_conv2_sum_d[10]) );
  OA21X1_HVT U516 ( .A1(DP_OP_425J2_127_3477_n47), .A2(
        DP_OP_425J2_127_3477_n161), .A3(DP_OP_425J2_127_3477_n48), .Y(n304) );
  INVX0_HVT U517 ( .A(DP_OP_425J2_127_3477_n44), .Y(n305) );
  NAND2X0_HVT U518 ( .A1(n305), .A2(DP_OP_425J2_127_3477_n45), .Y(n306) );
  HADDX1_HVT U519 ( .A0(n304), .B0(n306), .SO(n_conv2_sum_d[29]) );
  AND2X1_HVT U520 ( .A1(DP_OP_424J2_126_3477_n215), .A2(n450), .Y(n307) );
  HADDX1_HVT U521 ( .A0(n307), .B0(DP_OP_424J2_126_3477_n216), .SO(
        n_conv2_sum_c[2]) );
  AND2X1_HVT U522 ( .A1(DP_OP_424J2_126_3477_n207), .A2(n449), .Y(n308) );
  HADDX1_HVT U523 ( .A0(n308), .B0(DP_OP_424J2_126_3477_n208), .SO(
        n_conv2_sum_c[4]) );
  AND2X1_HVT U524 ( .A1(DP_OP_424J2_126_3477_n199), .A2(n448), .Y(n309) );
  HADDX1_HVT U525 ( .A0(n309), .B0(DP_OP_424J2_126_3477_n200), .SO(
        n_conv2_sum_c[6]) );
  OA21X1_HVT U526 ( .A1(DP_OP_424J2_126_3477_n189), .A2(
        DP_OP_424J2_126_3477_n191), .A3(DP_OP_424J2_126_3477_n190), .Y(n310)
         );
  INVX0_HVT U527 ( .A(DP_OP_424J2_126_3477_n186), .Y(n311) );
  NAND2X0_HVT U528 ( .A1(n311), .A2(DP_OP_424J2_126_3477_n187), .Y(n312) );
  HADDX1_HVT U529 ( .A0(n310), .B0(n312), .SO(n_conv2_sum_c[9]) );
  OA21X1_HVT U530 ( .A1(DP_OP_424J2_126_3477_n170), .A2(
        DP_OP_424J2_126_3477_n172), .A3(DP_OP_424J2_126_3477_n171), .Y(n313)
         );
  INVX0_HVT U531 ( .A(DP_OP_424J2_126_3477_n167), .Y(n314) );
  NAND2X0_HVT U532 ( .A1(n314), .A2(DP_OP_424J2_126_3477_n168), .Y(n315) );
  HADDX1_HVT U533 ( .A0(n313), .B0(n315), .SO(n_conv2_sum_c[13]) );
  OA21X1_HVT U534 ( .A1(DP_OP_424J2_126_3477_n39), .A2(
        DP_OP_424J2_126_3477_n41), .A3(DP_OP_424J2_126_3477_n40), .Y(n316) );
  NAND2X0_HVT U535 ( .A1(n442), .A2(DP_OP_424J2_126_3477_n37), .Y(n317) );
  HADDX1_HVT U536 ( .A0(n316), .B0(n317), .SO(n_conv2_sum_c[31]) );
  AND2X1_HVT U537 ( .A1(n537), .A2(mode[1]), .Y(n346) );
  INVX1_HVT U538 ( .A(mode[0]), .Y(n537) );
  MUX21X2_HVT U539 ( .A1(conv2_sram_rdata_weight[94]), .A2(
        conv1_sram_rdata_weight[94]), .S0(n398), .Y(conv_weight_box[94]) );
  MUX21X2_HVT U540 ( .A1(conv2_sram_rdata_weight[27]), .A2(
        conv1_sram_rdata_weight[27]), .S0(n399), .Y(conv_weight_box[27]) );
  INVX2_HVT U541 ( .A(n346), .Y(n403) );
  IBUFFX2_HVT U542 ( .A(DP_OP_425J2_127_3477_n181), .Y(
        DP_OP_425J2_127_3477_n179) );
  NOR2X0_HVT U543 ( .A1(DP_OP_422J2_124_3477_n2442), .A2(
        DP_OP_422J2_124_3477_n2445), .Y(DP_OP_422J2_124_3477_n2418) );
  IBUFFX2_HVT U544 ( .A(DP_OP_423J2_125_3477_n181), .Y(
        DP_OP_423J2_125_3477_n179) );
  MUX21X1_HVT U545 ( .A1(conv2_sram_rdata_weight[62]), .A2(
        conv1_sram_rdata_weight[62]), .S0(n404), .Y(conv_weight_box[62]) );
  MUX21X1_HVT U546 ( .A1(conv2_sram_rdata_weight[42]), .A2(
        conv1_sram_rdata_weight[42]), .S0(n403), .Y(conv_weight_box[42]) );
  MUX21X1_HVT U547 ( .A1(conv2_sram_rdata_weight[47]), .A2(
        conv1_sram_rdata_weight[47]), .S0(n401), .Y(conv_weight_box[47]) );
  MUX21X1_HVT U548 ( .A1(conv2_sram_rdata_weight[55]), .A2(
        conv1_sram_rdata_weight[55]), .S0(n404), .Y(conv_weight_box[55]) );
  MUX21X1_HVT U549 ( .A1(conv2_sram_rdata_weight[3]), .A2(
        conv1_sram_rdata_weight[3]), .S0(n403), .Y(conv_weight_box[3]) );
  INVX4_HVT U550 ( .A(n471), .Y(n464) );
  INVX1_HVT U551 ( .A(n394), .Y(n392) );
  INVX2_HVT U552 ( .A(n381), .Y(n402) );
  INVX2_HVT U553 ( .A(n346), .Y(n384) );
  INVX1_HVT U554 ( .A(n394), .Y(n395) );
  INVX0_HVT U555 ( .A(DP_OP_422J2_124_3477_n192), .Y(DP_OP_422J2_124_3477_n191) );
  INVX0_HVT U556 ( .A(DP_OP_425J2_127_3477_n192), .Y(DP_OP_425J2_127_3477_n191) );
  INVX0_HVT U557 ( .A(DP_OP_424J2_126_3477_n192), .Y(DP_OP_424J2_126_3477_n191) );
  INVX0_HVT U558 ( .A(DP_OP_423J2_125_3477_n192), .Y(DP_OP_423J2_125_3477_n191) );
  INVX0_HVT U559 ( .A(DP_OP_424J2_126_3477_n181), .Y(DP_OP_424J2_126_3477_n179) );
  INVX1_HVT U560 ( .A(N7), .Y(n419) );
  INVX1_HVT U561 ( .A(N7), .Y(n416) );
  MUX21X1_HVT U562 ( .A1(conv2_sram_rdata_weight[26]), .A2(
        conv1_sram_rdata_weight[26]), .S0(n399), .Y(conv_weight_box[26]) );
  INVX1_HVT U563 ( .A(n396), .Y(n399) );
  INVX1_HVT U564 ( .A(srstn), .Y(n382) );
  INVX0_HVT U565 ( .A(DP_OP_422J2_124_3477_n57), .Y(DP_OP_422J2_124_3477_n55)
         );
  INVX0_HVT U566 ( .A(DP_OP_425J2_127_3477_n57), .Y(DP_OP_425J2_127_3477_n55)
         );
  INVX0_HVT U567 ( .A(DP_OP_424J2_126_3477_n57), .Y(DP_OP_424J2_126_3477_n55)
         );
  INVX0_HVT U568 ( .A(DP_OP_423J2_125_3477_n57), .Y(DP_OP_423J2_125_3477_n55)
         );
  INVX0_HVT U569 ( .A(DP_OP_424J2_126_3477_n145), .Y(DP_OP_424J2_126_3477_n143) );
  INVX0_HVT U570 ( .A(DP_OP_424J2_126_3477_n144), .Y(DP_OP_424J2_126_3477_n142) );
  INVX0_HVT U571 ( .A(DP_OP_422J2_124_3477_n144), .Y(DP_OP_422J2_124_3477_n142) );
  INVX0_HVT U572 ( .A(DP_OP_422J2_124_3477_n145), .Y(DP_OP_422J2_124_3477_n143) );
  INVX0_HVT U573 ( .A(DP_OP_425J2_127_3477_n180), .Y(DP_OP_425J2_127_3477_n241) );
  INVX0_HVT U574 ( .A(DP_OP_423J2_125_3477_n180), .Y(DP_OP_423J2_125_3477_n241) );
  INVX0_HVT U575 ( .A(DP_OP_422J2_124_3477_n180), .Y(DP_OP_422J2_124_3477_n241) );
  INVX0_HVT U576 ( .A(DP_OP_424J2_126_3477_n180), .Y(DP_OP_424J2_126_3477_n241) );
  INVX1_HVT U577 ( .A(DP_OP_424J2_126_3477_n151), .Y(DP_OP_424J2_126_3477_n237) );
  INVX1_HVT U578 ( .A(DP_OP_422J2_124_3477_n151), .Y(DP_OP_422J2_124_3477_n237) );
  INVX1_HVT U579 ( .A(DP_OP_425J2_127_3477_n151), .Y(DP_OP_425J2_127_3477_n237) );
  INVX1_HVT U580 ( .A(DP_OP_423J2_125_3477_n151), .Y(DP_OP_423J2_125_3477_n237) );
  INVX0_HVT U581 ( .A(DP_OP_422J2_124_3477_n75), .Y(DP_OP_422J2_124_3477_n73)
         );
  INVX0_HVT U582 ( .A(DP_OP_422J2_124_3477_n74), .Y(DP_OP_422J2_124_3477_n72)
         );
  INVX0_HVT U583 ( .A(DP_OP_425J2_127_3477_n74), .Y(DP_OP_425J2_127_3477_n72)
         );
  INVX0_HVT U584 ( .A(DP_OP_425J2_127_3477_n75), .Y(DP_OP_425J2_127_3477_n73)
         );
  INVX0_HVT U585 ( .A(DP_OP_423J2_125_3477_n75), .Y(DP_OP_423J2_125_3477_n73)
         );
  INVX0_HVT U586 ( .A(DP_OP_424J2_126_3477_n75), .Y(DP_OP_424J2_126_3477_n73)
         );
  INVX0_HVT U587 ( .A(DP_OP_423J2_125_3477_n74), .Y(DP_OP_423J2_125_3477_n72)
         );
  INVX0_HVT U588 ( .A(DP_OP_424J2_126_3477_n74), .Y(DP_OP_424J2_126_3477_n72)
         );
  INVX0_HVT U589 ( .A(DP_OP_425J2_127_3477_n137), .Y(DP_OP_425J2_127_3477_n235) );
  INVX0_HVT U590 ( .A(DP_OP_423J2_125_3477_n137), .Y(DP_OP_423J2_125_3477_n235) );
  INVX0_HVT U591 ( .A(DP_OP_425J2_127_3477_n85), .Y(DP_OP_425J2_127_3477_n83)
         );
  INVX0_HVT U592 ( .A(DP_OP_425J2_127_3477_n86), .Y(DP_OP_425J2_127_3477_n84)
         );
  INVX0_HVT U593 ( .A(DP_OP_422J2_124_3477_n86), .Y(DP_OP_422J2_124_3477_n84)
         );
  INVX0_HVT U594 ( .A(DP_OP_422J2_124_3477_n85), .Y(DP_OP_422J2_124_3477_n83)
         );
  INVX0_HVT U595 ( .A(DP_OP_424J2_126_3477_n86), .Y(DP_OP_424J2_126_3477_n84)
         );
  INVX0_HVT U596 ( .A(DP_OP_424J2_126_3477_n85), .Y(DP_OP_424J2_126_3477_n83)
         );
  INVX0_HVT U597 ( .A(DP_OP_423J2_125_3477_n86), .Y(DP_OP_423J2_125_3477_n84)
         );
  INVX0_HVT U598 ( .A(DP_OP_423J2_125_3477_n85), .Y(DP_OP_423J2_125_3477_n83)
         );
  INVX0_HVT U599 ( .A(DP_OP_424J2_126_3477_n99), .Y(DP_OP_424J2_126_3477_n97)
         );
  INVX0_HVT U600 ( .A(DP_OP_424J2_126_3477_n100), .Y(DP_OP_424J2_126_3477_n98)
         );
  INVX0_HVT U601 ( .A(DP_OP_423J2_125_3477_n99), .Y(DP_OP_423J2_125_3477_n97)
         );
  INVX0_HVT U602 ( .A(DP_OP_423J2_125_3477_n100), .Y(DP_OP_423J2_125_3477_n98)
         );
  INVX0_HVT U603 ( .A(n733), .Y(n536) );
  INVX0_HVT U604 ( .A(DP_OP_422J2_124_3477_n99), .Y(DP_OP_422J2_124_3477_n97)
         );
  INVX0_HVT U605 ( .A(DP_OP_422J2_124_3477_n100), .Y(DP_OP_422J2_124_3477_n98)
         );
  INVX0_HVT U606 ( .A(DP_OP_425J2_127_3477_n99), .Y(DP_OP_425J2_127_3477_n97)
         );
  INVX0_HVT U607 ( .A(DP_OP_425J2_127_3477_n100), .Y(DP_OP_425J2_127_3477_n98)
         );
  INVX0_HVT U608 ( .A(DP_OP_425J2_127_3477_n114), .Y(DP_OP_425J2_127_3477_n112) );
  INVX0_HVT U609 ( .A(DP_OP_425J2_127_3477_n113), .Y(DP_OP_425J2_127_3477_n111) );
  INVX0_HVT U610 ( .A(DP_OP_422J2_124_3477_n114), .Y(DP_OP_422J2_124_3477_n112) );
  INVX0_HVT U611 ( .A(DP_OP_422J2_124_3477_n113), .Y(DP_OP_422J2_124_3477_n111) );
  INVX0_HVT U612 ( .A(DP_OP_423J2_125_3477_n113), .Y(DP_OP_423J2_125_3477_n111) );
  INVX0_HVT U613 ( .A(DP_OP_423J2_125_3477_n114), .Y(DP_OP_423J2_125_3477_n112) );
  INVX0_HVT U614 ( .A(DP_OP_424J2_126_3477_n113), .Y(DP_OP_424J2_126_3477_n111) );
  INVX0_HVT U615 ( .A(DP_OP_424J2_126_3477_n114), .Y(DP_OP_424J2_126_3477_n112) );
  INVX0_HVT U616 ( .A(n732), .Y(n467) );
  INVX0_HVT U617 ( .A(n710), .Y(n747) );
  INVX0_HVT U618 ( .A(DP_OP_425J2_127_3477_n219), .Y(DP_OP_425J2_127_3477_n4)
         );
  INVX0_HVT U619 ( .A(DP_OP_422J2_124_3477_n219), .Y(DP_OP_422J2_124_3477_n4)
         );
  INVX0_HVT U620 ( .A(DP_OP_423J2_125_3477_n219), .Y(DP_OP_423J2_125_3477_n4)
         );
  INVX0_HVT U621 ( .A(DP_OP_424J2_126_3477_n219), .Y(DP_OP_424J2_126_3477_n4)
         );
  INVX0_HVT U622 ( .A(DP_OP_424J2_126_3477_n127), .Y(DP_OP_424J2_126_3477_n125) );
  INVX0_HVT U623 ( .A(DP_OP_424J2_126_3477_n128), .Y(DP_OP_424J2_126_3477_n126) );
  INVX0_HVT U624 ( .A(tmp_big2[8]), .Y(n740) );
  INVX0_HVT U625 ( .A(DP_OP_423J2_125_3477_n127), .Y(DP_OP_423J2_125_3477_n125) );
  INVX0_HVT U626 ( .A(DP_OP_423J2_125_3477_n128), .Y(DP_OP_423J2_125_3477_n126) );
  INVX0_HVT U627 ( .A(DP_OP_422J2_124_3477_n128), .Y(DP_OP_422J2_124_3477_n126) );
  INVX0_HVT U628 ( .A(DP_OP_422J2_124_3477_n127), .Y(DP_OP_422J2_124_3477_n125) );
  INVX0_HVT U629 ( .A(DP_OP_425J2_127_3477_n127), .Y(DP_OP_425J2_127_3477_n125) );
  INVX0_HVT U630 ( .A(DP_OP_425J2_127_3477_n128), .Y(DP_OP_425J2_127_3477_n126) );
  INVX0_HVT U631 ( .A(DP_OP_422J2_124_3477_n87), .Y(DP_OP_422J2_124_3477_n227)
         );
  INVX0_HVT U632 ( .A(DP_OP_422J2_124_3477_n101), .Y(DP_OP_422J2_124_3477_n229) );
  INVX0_HVT U633 ( .A(DP_OP_422J2_124_3477_n115), .Y(DP_OP_422J2_124_3477_n231) );
  INVX0_HVT U634 ( .A(DP_OP_425J2_127_3477_n132), .Y(DP_OP_425J2_127_3477_n234) );
  INVX0_HVT U635 ( .A(DP_OP_425J2_127_3477_n129), .Y(DP_OP_425J2_127_3477_n233) );
  INVX0_HVT U636 ( .A(DP_OP_425J2_127_3477_n115), .Y(DP_OP_425J2_127_3477_n231) );
  INVX0_HVT U637 ( .A(DP_OP_425J2_127_3477_n101), .Y(DP_OP_425J2_127_3477_n229) );
  INVX0_HVT U638 ( .A(DP_OP_422J2_124_3477_n129), .Y(DP_OP_422J2_124_3477_n233) );
  INVX0_HVT U639 ( .A(DP_OP_425J2_127_3477_n87), .Y(DP_OP_425J2_127_3477_n227)
         );
  INVX0_HVT U640 ( .A(tmp_big1[30]), .Y(n759) );
  INVX0_HVT U641 ( .A(DP_OP_423J2_125_3477_n87), .Y(DP_OP_423J2_125_3477_n227)
         );
  INVX0_HVT U642 ( .A(DP_OP_423J2_125_3477_n101), .Y(DP_OP_423J2_125_3477_n229) );
  INVX0_HVT U643 ( .A(DP_OP_423J2_125_3477_n115), .Y(DP_OP_423J2_125_3477_n231) );
  INVX0_HVT U644 ( .A(DP_OP_423J2_125_3477_n129), .Y(DP_OP_423J2_125_3477_n233) );
  INVX0_HVT U645 ( .A(tmp_big1[14]), .Y(n745) );
  INVX0_HVT U646 ( .A(DP_OP_423J2_125_3477_n132), .Y(DP_OP_423J2_125_3477_n234) );
  INVX0_HVT U647 ( .A(DP_OP_424J2_126_3477_n101), .Y(DP_OP_424J2_126_3477_n229) );
  INVX0_HVT U648 ( .A(DP_OP_424J2_126_3477_n129), .Y(DP_OP_424J2_126_3477_n233) );
  INVX0_HVT U649 ( .A(tmp_big1[6]), .Y(n762) );
  INVX0_HVT U650 ( .A(DP_OP_424J2_126_3477_n115), .Y(DP_OP_424J2_126_3477_n231) );
  INVX0_HVT U651 ( .A(tmp_big1[10]), .Y(n741) );
  INVX0_HVT U652 ( .A(tmp_big1[4]), .Y(n760) );
  INVX0_HVT U653 ( .A(DP_OP_424J2_126_3477_n87), .Y(DP_OP_424J2_126_3477_n227)
         );
  INVX0_HVT U654 ( .A(tmp_big1[22]), .Y(n752) );
  INVX0_HVT U655 ( .A(tmp_big1[12]), .Y(n743) );
  INVX0_HVT U656 ( .A(tmp_big1[2]), .Y(n758) );
  INVX1_HVT U657 ( .A(N7), .Y(n417) );
  MUX21X1_HVT U658 ( .A1(conv2_sram_rdata_weight[87]), .A2(
        conv1_sram_rdata_weight[87]), .S0(n393), .Y(conv_weight_box[87]) );
  MUX21X1_HVT U659 ( .A1(conv2_sram_rdata_weight[39]), .A2(
        conv1_sram_rdata_weight[39]), .S0(n402), .Y(conv_weight_box[39]) );
  MUX21X1_HVT U660 ( .A1(conv2_sram_rdata_weight[83]), .A2(
        conv1_sram_rdata_weight[83]), .S0(n402), .Y(conv_weight_box[83]) );
  MUX21X1_HVT U661 ( .A1(conv2_sram_rdata_weight[99]), .A2(
        conv1_sram_rdata_weight[99]), .S0(n401), .Y(conv_weight_box[99]) );
  MUX21X1_HVT U662 ( .A1(conv2_sram_rdata_weight[79]), .A2(
        conv1_sram_rdata_weight[79]), .S0(n393), .Y(conv_weight_box[79]) );
  MUX21X1_HVT U663 ( .A1(conv2_sram_rdata_weight[67]), .A2(
        conv1_sram_rdata_weight[67]), .S0(n400), .Y(conv_weight_box[67]) );
  MUX21X1_HVT U664 ( .A1(conv2_sram_rdata_weight[75]), .A2(
        conv1_sram_rdata_weight[75]), .S0(n399), .Y(conv_weight_box[75]) );
  MUX21X1_HVT U665 ( .A1(conv2_sram_rdata_weight[43]), .A2(
        conv1_sram_rdata_weight[43]), .S0(n395), .Y(conv_weight_box[43]) );
  MUX21X1_HVT U666 ( .A1(conv2_sram_rdata_weight[51]), .A2(
        conv1_sram_rdata_weight[51]), .S0(n402), .Y(conv_weight_box[51]) );
  MUX21X1_HVT U667 ( .A1(conv2_sram_rdata_weight[71]), .A2(
        conv1_sram_rdata_weight[71]), .S0(n398), .Y(conv_weight_box[71]) );
  MUX21X1_HVT U668 ( .A1(conv2_sram_rdata_weight[31]), .A2(
        conv1_sram_rdata_weight[31]), .S0(n401), .Y(conv_weight_box[31]) );
  MUX21X1_HVT U669 ( .A1(conv2_sram_rdata_weight[91]), .A2(
        conv1_sram_rdata_weight[91]), .S0(n393), .Y(conv_weight_box[91]) );
  MUX21X1_HVT U670 ( .A1(conv2_sram_rdata_weight[95]), .A2(
        conv1_sram_rdata_weight[95]), .S0(n384), .Y(conv_weight_box[95]) );
  MUX21X1_HVT U671 ( .A1(conv2_sram_rdata_weight[35]), .A2(
        conv1_sram_rdata_weight[35]), .S0(n398), .Y(conv_weight_box[35]) );
  MUX21X1_HVT U672 ( .A1(conv2_sram_rdata_weight[59]), .A2(
        conv1_sram_rdata_weight[59]), .S0(n398), .Y(conv_weight_box[59]) );
  MUX21X1_HVT U673 ( .A1(conv2_sram_rdata_weight[23]), .A2(
        conv1_sram_rdata_weight[23]), .S0(n395), .Y(conv_weight_box[23]) );
  MUX21X1_HVT U674 ( .A1(conv2_sram_rdata_weight[11]), .A2(
        conv1_sram_rdata_weight[11]), .S0(n393), .Y(conv_weight_box[11]) );
  INVX1_HVT U675 ( .A(DP_OP_425J2_127_3477_n3054), .Y(n391) );
  INVX1_HVT U676 ( .A(DP_OP_425J2_127_3477_n3054), .Y(DP_OP_425J2_127_3477_n2)
         );
  INVX1_HVT U677 ( .A(DP_OP_425J2_127_3477_n3054), .Y(n390) );
  INVX1_HVT U678 ( .A(DP_OP_425J2_127_3477_n3054), .Y(n389) );
  MUX21X1_HVT U679 ( .A1(conv2_sram_rdata_weight[15]), .A2(
        conv1_sram_rdata_weight[15]), .S0(n401), .Y(conv_weight_box[15]) );
  MUX21X1_HVT U680 ( .A1(conv2_sram_rdata_weight[19]), .A2(
        conv1_sram_rdata_weight[19]), .S0(n400), .Y(conv_weight_box[19]) );
  INVX1_HVT U681 ( .A(n396), .Y(n397) );
  INVX1_HVT U682 ( .A(srstn), .Y(n383) );
  NOR2X1_HVT U683 ( .A1(n559), .A2(n558), .Y(n610) );
  NOR2X1_HVT U684 ( .A1(n624), .A2(n623), .Y(n672) );
  INVX1_HVT U685 ( .A(DP_OP_425J2_127_3477_n3054), .Y(n385) );
  INVX1_HVT U686 ( .A(DP_OP_425J2_127_3477_n3054), .Y(n386) );
  INVX1_HVT U687 ( .A(DP_OP_425J2_127_3477_n3054), .Y(n387) );
  INVX1_HVT U688 ( .A(DP_OP_425J2_127_3477_n3054), .Y(n388) );
  INVX2_HVT U689 ( .A(n381), .Y(n393) );
  INVX1_HVT U690 ( .A(n384), .Y(n394) );
  INVX1_HVT U691 ( .A(n384), .Y(n396) );
  INVX1_HVT U692 ( .A(n396), .Y(n398) );
  INVX2_HVT U693 ( .A(srstn), .Y(n407) );
  INVX1_HVT U694 ( .A(srstn), .Y(n408) );
  INVX2_HVT U695 ( .A(srstn), .Y(n406) );
  INVX2_HVT U696 ( .A(srstn), .Y(n405) );
  INVX2_HVT U697 ( .A(n346), .Y(n404) );
  INVX2_HVT U698 ( .A(n381), .Y(n401) );
  INVX8_HVT U699 ( .A(n464), .Y(n409) );
  INVX2_HVT U700 ( .A(n464), .Y(n410) );
  INVX2_HVT U701 ( .A(n464), .Y(n411) );
  AND2X1_HVT U702 ( .A1(n614), .A2(n613), .Y(N5) );
  INVX1_HVT U703 ( .A(N5), .Y(n412) );
  INVX0_HVT U704 ( .A(N5), .Y(n413) );
  INVX0_HVT U705 ( .A(N5), .Y(n414) );
  INVX1_HVT U706 ( .A(N5), .Y(n415) );
  AND2X1_HVT U707 ( .A1(n676), .A2(n675), .Y(N7) );
  INVX0_HVT U708 ( .A(N7), .Y(n418) );
  INVX1_HVT U709 ( .A(DP_OP_422J2_124_3477_n148), .Y(DP_OP_422J2_124_3477_n236) );
  INVX1_HVT U710 ( .A(DP_OP_422J2_124_3477_n152), .Y(DP_OP_422J2_124_3477_n158) );
  INVX1_HVT U711 ( .A(DP_OP_422J2_124_3477_n1678), .Y(
        DP_OP_422J2_124_3477_n1679) );
  INVX1_HVT U712 ( .A(DP_OP_422J2_124_3477_n183), .Y(DP_OP_422J2_124_3477_n182) );
  INVX1_HVT U713 ( .A(src_window[66]), .Y(DP_OP_422J2_124_3477_n1957) );
  INVX1_HVT U714 ( .A(src_window[65]), .Y(DP_OP_422J2_124_3477_n1958) );
  INVX1_HVT U715 ( .A(conv_weight_box[6]), .Y(DP_OP_422J2_124_3477_n1961) );
  INVX1_HVT U716 ( .A(conv_weight_box[5]), .Y(DP_OP_422J2_124_3477_n1962) );
  INVX1_HVT U717 ( .A(conv_weight_box[4]), .Y(DP_OP_422J2_124_3477_n1963) );
  INVX1_HVT U718 ( .A(src_window[83]), .Y(DP_OP_422J2_124_3477_n2000) );
  INVX1_HVT U719 ( .A(conv_weight_box[15]), .Y(DP_OP_422J2_124_3477_n2004) );
  INVX1_HVT U720 ( .A(conv_weight_box[14]), .Y(DP_OP_422J2_124_3477_n2005) );
  INVX1_HVT U721 ( .A(conv_weight_box[13]), .Y(DP_OP_422J2_124_3477_n2006) );
  INVX1_HVT U722 ( .A(conv_weight_box[12]), .Y(DP_OP_422J2_124_3477_n2007) );
  INVX1_HVT U723 ( .A(src_window[111]), .Y(DP_OP_422J2_124_3477_n2040) );
  INVX1_HVT U724 ( .A(src_window[107]), .Y(DP_OP_422J2_124_3477_n2044) );
  INVX1_HVT U725 ( .A(src_window[106]), .Y(DP_OP_422J2_124_3477_n2045) );
  INVX1_HVT U726 ( .A(src_window[104]), .Y(DP_OP_422J2_124_3477_n2047) );
  INVX1_HVT U727 ( .A(conv_weight_box[23]), .Y(DP_OP_422J2_124_3477_n2048) );
  INVX1_HVT U728 ( .A(conv_weight_box[22]), .Y(DP_OP_422J2_124_3477_n2049) );
  INVX1_HVT U729 ( .A(conv_weight_box[21]), .Y(DP_OP_422J2_124_3477_n2050) );
  INVX1_HVT U730 ( .A(conv_weight_box[20]), .Y(DP_OP_422J2_124_3477_n2051) );
  INVX1_HVT U731 ( .A(src_window[127]), .Y(DP_OP_422J2_124_3477_n2084) );
  INVX1_HVT U732 ( .A(src_window[123]), .Y(DP_OP_422J2_124_3477_n2088) );
  INVX1_HVT U733 ( .A(src_window[121]), .Y(DP_OP_422J2_124_3477_n2090) );
  INVX1_HVT U734 ( .A(src_window[120]), .Y(DP_OP_422J2_124_3477_n2091) );
  INVX1_HVT U735 ( .A(conv_weight_box[31]), .Y(DP_OP_422J2_124_3477_n2092) );
  INVX1_HVT U736 ( .A(conv_weight_box[30]), .Y(DP_OP_422J2_124_3477_n2093) );
  INVX1_HVT U737 ( .A(conv_weight_box[29]), .Y(DP_OP_422J2_124_3477_n2094) );
  INVX1_HVT U738 ( .A(conv_weight_box[28]), .Y(DP_OP_422J2_124_3477_n2095) );
  INVX1_HVT U739 ( .A(src_window[142]), .Y(DP_OP_422J2_124_3477_n2129) );
  INVX1_HVT U740 ( .A(src_window[141]), .Y(DP_OP_422J2_124_3477_n2130) );
  INVX1_HVT U741 ( .A(src_window[139]), .Y(DP_OP_422J2_124_3477_n2132) );
  INVX1_HVT U742 ( .A(src_window[137]), .Y(DP_OP_422J2_124_3477_n2134) );
  INVX1_HVT U743 ( .A(src_window[136]), .Y(DP_OP_422J2_124_3477_n2135) );
  INVX1_HVT U744 ( .A(conv_weight_box[39]), .Y(DP_OP_422J2_124_3477_n2136) );
  INVX1_HVT U745 ( .A(conv_weight_box[38]), .Y(DP_OP_422J2_124_3477_n2137) );
  INVX1_HVT U746 ( .A(conv_weight_box[37]), .Y(DP_OP_422J2_124_3477_n2138) );
  INVX1_HVT U747 ( .A(conv_weight_box[36]), .Y(DP_OP_422J2_124_3477_n2139) );
  INVX1_HVT U748 ( .A(src_window[167]), .Y(DP_OP_422J2_124_3477_n2172) );
  INVX1_HVT U749 ( .A(src_window[162]), .Y(DP_OP_422J2_124_3477_n2177) );
  INVX1_HVT U750 ( .A(src_window[161]), .Y(DP_OP_422J2_124_3477_n2178) );
  INVX1_HVT U751 ( .A(src_window[160]), .Y(DP_OP_422J2_124_3477_n2179) );
  INVX1_HVT U752 ( .A(conv_weight_box[47]), .Y(DP_OP_422J2_124_3477_n2180) );
  INVX1_HVT U753 ( .A(conv_weight_box[46]), .Y(DP_OP_422J2_124_3477_n2181) );
  INVX1_HVT U754 ( .A(conv_weight_box[45]), .Y(DP_OP_422J2_124_3477_n2182) );
  INVX1_HVT U755 ( .A(conv_weight_box[44]), .Y(DP_OP_422J2_124_3477_n2183) );
  INVX1_HVT U756 ( .A(src_window[182]), .Y(DP_OP_422J2_124_3477_n2217) );
  INVX1_HVT U757 ( .A(src_window[181]), .Y(DP_OP_422J2_124_3477_n2218) );
  INVX1_HVT U758 ( .A(src_window[180]), .Y(DP_OP_422J2_124_3477_n2219) );
  INVX1_HVT U759 ( .A(src_window[179]), .Y(DP_OP_422J2_124_3477_n2220) );
  INVX1_HVT U760 ( .A(conv_weight_box[55]), .Y(DP_OP_422J2_124_3477_n2224) );
  INVX1_HVT U761 ( .A(conv_weight_box[54]), .Y(DP_OP_422J2_124_3477_n2225) );
  INVX1_HVT U762 ( .A(conv_weight_box[52]), .Y(DP_OP_422J2_124_3477_n2227) );
  INVX1_HVT U763 ( .A(src_window[207]), .Y(DP_OP_422J2_124_3477_n2260) );
  INVX1_HVT U764 ( .A(src_window[206]), .Y(DP_OP_422J2_124_3477_n2261) );
  INVX1_HVT U765 ( .A(src_window[205]), .Y(DP_OP_422J2_124_3477_n2262) );
  INVX1_HVT U766 ( .A(src_window[204]), .Y(DP_OP_422J2_124_3477_n2263) );
  INVX1_HVT U767 ( .A(src_window[202]), .Y(DP_OP_422J2_124_3477_n2265) );
  INVX1_HVT U768 ( .A(src_window[200]), .Y(DP_OP_422J2_124_3477_n2267) );
  INVX1_HVT U769 ( .A(conv_weight_box[63]), .Y(DP_OP_422J2_124_3477_n2268) );
  INVX1_HVT U770 ( .A(conv_weight_box[62]), .Y(DP_OP_422J2_124_3477_n2269) );
  INVX1_HVT U771 ( .A(conv_weight_box[61]), .Y(DP_OP_422J2_124_3477_n2270) );
  INVX1_HVT U772 ( .A(conv_weight_box[60]), .Y(DP_OP_422J2_124_3477_n2271) );
  INVX1_HVT U773 ( .A(src_window[223]), .Y(DP_OP_422J2_124_3477_n2304) );
  INVX1_HVT U774 ( .A(src_window[222]), .Y(DP_OP_422J2_124_3477_n2305) );
  INVX1_HVT U775 ( .A(src_window[220]), .Y(DP_OP_422J2_124_3477_n2307) );
  INVX1_HVT U776 ( .A(src_window[219]), .Y(DP_OP_422J2_124_3477_n2308) );
  INVX1_HVT U777 ( .A(src_window[216]), .Y(DP_OP_422J2_124_3477_n2311) );
  INVX1_HVT U778 ( .A(conv_weight_box[71]), .Y(DP_OP_422J2_124_3477_n2312) );
  INVX1_HVT U779 ( .A(conv_weight_box[70]), .Y(DP_OP_422J2_124_3477_n2313) );
  INVX1_HVT U780 ( .A(conv_weight_box[68]), .Y(DP_OP_422J2_124_3477_n2315) );
  INVX1_HVT U781 ( .A(src_window[239]), .Y(DP_OP_422J2_124_3477_n2348) );
  INVX1_HVT U782 ( .A(src_window[236]), .Y(DP_OP_422J2_124_3477_n2351) );
  INVX1_HVT U783 ( .A(src_window[234]), .Y(DP_OP_422J2_124_3477_n2353) );
  INVX1_HVT U784 ( .A(src_window[233]), .Y(DP_OP_422J2_124_3477_n2354) );
  INVX1_HVT U785 ( .A(src_window[232]), .Y(DP_OP_422J2_124_3477_n2355) );
  INVX1_HVT U786 ( .A(conv_weight_box[79]), .Y(DP_OP_422J2_124_3477_n2356) );
  INVX1_HVT U787 ( .A(conv_weight_box[78]), .Y(DP_OP_422J2_124_3477_n2357) );
  INVX1_HVT U788 ( .A(conv_weight_box[77]), .Y(DP_OP_422J2_124_3477_n2358) );
  INVX1_HVT U789 ( .A(conv_weight_box[76]), .Y(DP_OP_422J2_124_3477_n2359) );
  INVX1_HVT U790 ( .A(src_window[263]), .Y(DP_OP_422J2_124_3477_n2392) );
  INVX1_HVT U791 ( .A(DP_OP_422J2_124_3477_n175), .Y(DP_OP_422J2_124_3477_n240) );
  INVX1_HVT U792 ( .A(conv_weight_box[87]), .Y(DP_OP_422J2_124_3477_n2400) );
  INVX1_HVT U793 ( .A(conv_weight_box[86]), .Y(DP_OP_422J2_124_3477_n2401) );
  INVX1_HVT U794 ( .A(conv_weight_box[84]), .Y(DP_OP_422J2_124_3477_n2403) );
  INVX1_HVT U795 ( .A(src_window[279]), .Y(DP_OP_422J2_124_3477_n2436) );
  INVX1_HVT U796 ( .A(src_window[276]), .Y(DP_OP_422J2_124_3477_n2439) );
  INVX1_HVT U797 ( .A(src_window[274]), .Y(DP_OP_422J2_124_3477_n2441) );
  INVX1_HVT U798 ( .A(src_window[273]), .Y(DP_OP_422J2_124_3477_n2442) );
  INVX1_HVT U799 ( .A(conv_weight_box[95]), .Y(DP_OP_422J2_124_3477_n2444) );
  INVX1_HVT U800 ( .A(conv_weight_box[94]), .Y(DP_OP_422J2_124_3477_n2445) );
  INVX1_HVT U801 ( .A(conv_weight_box[93]), .Y(DP_OP_422J2_124_3477_n2446) );
  INVX1_HVT U802 ( .A(conv_weight_box[92]), .Y(DP_OP_422J2_124_3477_n2447) );
  INVX1_HVT U803 ( .A(src_window[287]), .Y(DP_OP_422J2_124_3477_n2480) );
  INVX1_HVT U804 ( .A(src_window[286]), .Y(DP_OP_422J2_124_3477_n2481) );
  INVX1_HVT U805 ( .A(src_window[285]), .Y(DP_OP_422J2_124_3477_n2482) );
  INVX1_HVT U806 ( .A(src_window[284]), .Y(DP_OP_422J2_124_3477_n2483) );
  INVX1_HVT U807 ( .A(src_window[283]), .Y(DP_OP_422J2_124_3477_n2484) );
  INVX1_HVT U808 ( .A(src_window[282]), .Y(DP_OP_422J2_124_3477_n2485) );
  INVX1_HVT U809 ( .A(src_window[281]), .Y(DP_OP_422J2_124_3477_n2486) );
  INVX1_HVT U810 ( .A(src_window[280]), .Y(DP_OP_422J2_124_3477_n2487) );
  INVX1_HVT U811 ( .A(conv_weight_box[99]), .Y(DP_OP_422J2_124_3477_n2488) );
  INVX1_HVT U812 ( .A(conv_weight_box[98]), .Y(DP_OP_422J2_124_3477_n2489) );
  INVX1_HVT U813 ( .A(conv_weight_box[97]), .Y(DP_OP_422J2_124_3477_n2490) );
  INVX1_HVT U814 ( .A(conv_weight_box[96]), .Y(DP_OP_422J2_124_3477_n2491) );
  INVX1_HVT U815 ( .A(src_window[269]), .Y(DP_OP_422J2_124_3477_n2526) );
  INVX1_HVT U816 ( .A(src_window[267]), .Y(DP_OP_422J2_124_3477_n2528) );
  INVX1_HVT U817 ( .A(DP_OP_422J2_124_3477_n252), .Y(DP_OP_422J2_124_3477_n253) );
  INVX1_HVT U818 ( .A(src_window[264]), .Y(DP_OP_422J2_124_3477_n2531) );
  INVX1_HVT U819 ( .A(conv_weight_box[91]), .Y(DP_OP_422J2_124_3477_n2532) );
  INVX1_HVT U820 ( .A(conv_weight_box[90]), .Y(DP_OP_422J2_124_3477_n2533) );
  INVX1_HVT U821 ( .A(conv_weight_box[89]), .Y(DP_OP_422J2_124_3477_n2534) );
  INVX1_HVT U822 ( .A(conv_weight_box[88]), .Y(DP_OP_422J2_124_3477_n2535) );
  INVX1_HVT U823 ( .A(DP_OP_422J2_124_3477_n254), .Y(DP_OP_422J2_124_3477_n255) );
  INVX1_HVT U824 ( .A(src_window[255]), .Y(DP_OP_422J2_124_3477_n2568) );
  INVX1_HVT U825 ( .A(src_window[254]), .Y(DP_OP_422J2_124_3477_n2569) );
  INVX1_HVT U826 ( .A(DP_OP_422J2_124_3477_n256), .Y(DP_OP_422J2_124_3477_n257) );
  INVX1_HVT U827 ( .A(src_window[253]), .Y(DP_OP_422J2_124_3477_n2570) );
  INVX1_HVT U828 ( .A(src_window[252]), .Y(DP_OP_422J2_124_3477_n2571) );
  INVX1_HVT U829 ( .A(src_window[248]), .Y(DP_OP_422J2_124_3477_n2575) );
  INVX1_HVT U830 ( .A(conv_weight_box[83]), .Y(DP_OP_422J2_124_3477_n2576) );
  INVX1_HVT U831 ( .A(conv_weight_box[82]), .Y(DP_OP_422J2_124_3477_n2577) );
  INVX1_HVT U832 ( .A(conv_weight_box[81]), .Y(DP_OP_422J2_124_3477_n2578) );
  INVX1_HVT U833 ( .A(conv_weight_box[80]), .Y(DP_OP_422J2_124_3477_n2579) );
  INVX1_HVT U834 ( .A(DP_OP_422J2_124_3477_n258), .Y(DP_OP_422J2_124_3477_n259) );
  INVX1_HVT U835 ( .A(DP_OP_422J2_124_3477_n260), .Y(DP_OP_422J2_124_3477_n261) );
  INVX1_HVT U836 ( .A(src_window[231]), .Y(DP_OP_422J2_124_3477_n2612) );
  INVX1_HVT U837 ( .A(src_window[230]), .Y(DP_OP_422J2_124_3477_n2613) );
  INVX1_HVT U838 ( .A(src_window[227]), .Y(DP_OP_422J2_124_3477_n2616) );
  INVX1_HVT U839 ( .A(src_window[226]), .Y(DP_OP_422J2_124_3477_n2617) );
  INVX1_HVT U840 ( .A(src_window[224]), .Y(DP_OP_422J2_124_3477_n2619) );
  INVX1_HVT U841 ( .A(conv_weight_box[75]), .Y(DP_OP_422J2_124_3477_n2620) );
  INVX1_HVT U842 ( .A(conv_weight_box[74]), .Y(DP_OP_422J2_124_3477_n2621) );
  INVX1_HVT U843 ( .A(conv_weight_box[73]), .Y(DP_OP_422J2_124_3477_n2622) );
  INVX1_HVT U844 ( .A(conv_weight_box[72]), .Y(DP_OP_422J2_124_3477_n2623) );
  INVX1_HVT U845 ( .A(DP_OP_422J2_124_3477_n262), .Y(DP_OP_422J2_124_3477_n263) );
  INVX1_HVT U846 ( .A(DP_OP_422J2_124_3477_n264), .Y(DP_OP_422J2_124_3477_n265) );
  INVX1_HVT U847 ( .A(src_window[215]), .Y(DP_OP_422J2_124_3477_n2656) );
  INVX1_HVT U848 ( .A(src_window[213]), .Y(DP_OP_422J2_124_3477_n2658) );
  INVX1_HVT U849 ( .A(src_window[212]), .Y(DP_OP_422J2_124_3477_n2659) );
  INVX1_HVT U850 ( .A(src_window[209]), .Y(DP_OP_422J2_124_3477_n2662) );
  INVX1_HVT U851 ( .A(src_window[208]), .Y(DP_OP_422J2_124_3477_n2663) );
  INVX1_HVT U852 ( .A(conv_weight_box[67]), .Y(DP_OP_422J2_124_3477_n2664) );
  INVX1_HVT U853 ( .A(conv_weight_box[65]), .Y(DP_OP_422J2_124_3477_n2666) );
  INVX1_HVT U854 ( .A(conv_weight_box[64]), .Y(DP_OP_422J2_124_3477_n2667) );
  INVX1_HVT U855 ( .A(DP_OP_422J2_124_3477_n266), .Y(DP_OP_422J2_124_3477_n267) );
  INVX1_HVT U856 ( .A(DP_OP_422J2_124_3477_n268), .Y(DP_OP_422J2_124_3477_n269) );
  INVX1_HVT U857 ( .A(src_window[191]), .Y(DP_OP_422J2_124_3477_n2700) );
  INVX1_HVT U858 ( .A(src_window[190]), .Y(DP_OP_422J2_124_3477_n2701) );
  INVX1_HVT U859 ( .A(src_window[189]), .Y(DP_OP_422J2_124_3477_n2702) );
  INVX1_HVT U860 ( .A(src_window[187]), .Y(DP_OP_422J2_124_3477_n2704) );
  INVX1_HVT U861 ( .A(src_window[184]), .Y(DP_OP_422J2_124_3477_n2707) );
  INVX1_HVT U862 ( .A(conv_weight_box[59]), .Y(DP_OP_422J2_124_3477_n2708) );
  INVX1_HVT U863 ( .A(conv_weight_box[58]), .Y(DP_OP_422J2_124_3477_n2709) );
  INVX1_HVT U864 ( .A(DP_OP_422J2_124_3477_n270), .Y(DP_OP_422J2_124_3477_n271) );
  INVX1_HVT U865 ( .A(conv_weight_box[57]), .Y(DP_OP_422J2_124_3477_n2710) );
  INVX1_HVT U866 ( .A(conv_weight_box[56]), .Y(DP_OP_422J2_124_3477_n2711) );
  INVX1_HVT U867 ( .A(DP_OP_422J2_124_3477_n272), .Y(DP_OP_422J2_124_3477_n273) );
  INVX1_HVT U868 ( .A(src_window[174]), .Y(DP_OP_422J2_124_3477_n2745) );
  INVX1_HVT U869 ( .A(src_window[173]), .Y(DP_OP_422J2_124_3477_n2746) );
  INVX1_HVT U870 ( .A(src_window[172]), .Y(DP_OP_422J2_124_3477_n2747) );
  INVX1_HVT U871 ( .A(src_window[170]), .Y(DP_OP_422J2_124_3477_n2749) );
  INVX1_HVT U872 ( .A(DP_OP_422J2_124_3477_n274), .Y(DP_OP_422J2_124_3477_n275) );
  INVX1_HVT U873 ( .A(src_window[169]), .Y(DP_OP_422J2_124_3477_n2750) );
  INVX1_HVT U874 ( .A(src_window[168]), .Y(DP_OP_422J2_124_3477_n2751) );
  INVX1_HVT U875 ( .A(conv_weight_box[51]), .Y(DP_OP_422J2_124_3477_n2752) );
  INVX1_HVT U876 ( .A(conv_weight_box[50]), .Y(DP_OP_422J2_124_3477_n2753) );
  INVX1_HVT U877 ( .A(conv_weight_box[49]), .Y(DP_OP_422J2_124_3477_n2754) );
  INVX1_HVT U878 ( .A(conv_weight_box[48]), .Y(DP_OP_422J2_124_3477_n2755) );
  INVX1_HVT U879 ( .A(DP_OP_422J2_124_3477_n276), .Y(DP_OP_422J2_124_3477_n277) );
  INVX1_HVT U880 ( .A(src_window[158]), .Y(DP_OP_422J2_124_3477_n2789) );
  INVX1_HVT U881 ( .A(DP_OP_422J2_124_3477_n278), .Y(DP_OP_422J2_124_3477_n279) );
  INVX1_HVT U882 ( .A(src_window[157]), .Y(DP_OP_422J2_124_3477_n2790) );
  INVX1_HVT U883 ( .A(src_window[156]), .Y(DP_OP_422J2_124_3477_n2791) );
  INVX1_HVT U884 ( .A(src_window[155]), .Y(DP_OP_422J2_124_3477_n2792) );
  INVX1_HVT U885 ( .A(src_window[154]), .Y(DP_OP_422J2_124_3477_n2793) );
  INVX1_HVT U886 ( .A(src_window[152]), .Y(DP_OP_422J2_124_3477_n2795) );
  INVX1_HVT U887 ( .A(conv_weight_box[43]), .Y(DP_OP_422J2_124_3477_n2796) );
  INVX1_HVT U888 ( .A(conv_weight_box[42]), .Y(DP_OP_422J2_124_3477_n2797) );
  INVX1_HVT U889 ( .A(conv_weight_box[41]), .Y(DP_OP_422J2_124_3477_n2798) );
  INVX1_HVT U890 ( .A(conv_weight_box[40]), .Y(DP_OP_422J2_124_3477_n2799) );
  INVX1_HVT U891 ( .A(DP_OP_422J2_124_3477_n280), .Y(DP_OP_422J2_124_3477_n281) );
  INVX1_HVT U892 ( .A(src_window[134]), .Y(DP_OP_422J2_124_3477_n2833) );
  INVX1_HVT U893 ( .A(src_window[133]), .Y(DP_OP_422J2_124_3477_n2834) );
  INVX1_HVT U894 ( .A(src_window[132]), .Y(DP_OP_422J2_124_3477_n2835) );
  INVX1_HVT U895 ( .A(src_window[130]), .Y(DP_OP_422J2_124_3477_n2837) );
  INVX1_HVT U896 ( .A(src_window[129]), .Y(DP_OP_422J2_124_3477_n2838) );
  INVX1_HVT U897 ( .A(conv_weight_box[35]), .Y(DP_OP_422J2_124_3477_n2840) );
  INVX1_HVT U898 ( .A(conv_weight_box[34]), .Y(DP_OP_422J2_124_3477_n2841) );
  INVX1_HVT U899 ( .A(conv_weight_box[33]), .Y(DP_OP_422J2_124_3477_n2842) );
  INVX1_HVT U900 ( .A(conv_weight_box[32]), .Y(DP_OP_422J2_124_3477_n2843) );
  INVX1_HVT U901 ( .A(src_window[118]), .Y(DP_OP_422J2_124_3477_n2877) );
  INVX1_HVT U902 ( .A(src_window[117]), .Y(DP_OP_422J2_124_3477_n2878) );
  INVX1_HVT U903 ( .A(src_window[115]), .Y(DP_OP_422J2_124_3477_n2880) );
  INVX1_HVT U904 ( .A(src_window[112]), .Y(DP_OP_422J2_124_3477_n2883) );
  INVX1_HVT U905 ( .A(conv_weight_box[27]), .Y(DP_OP_422J2_124_3477_n2884) );
  INVX1_HVT U906 ( .A(conv_weight_box[26]), .Y(DP_OP_422J2_124_3477_n2885) );
  INVX1_HVT U907 ( .A(conv_weight_box[25]), .Y(DP_OP_422J2_124_3477_n2886) );
  INVX1_HVT U908 ( .A(conv_weight_box[24]), .Y(DP_OP_422J2_124_3477_n2887) );
  INVX1_HVT U909 ( .A(src_window[94]), .Y(DP_OP_422J2_124_3477_n2921) );
  INVX1_HVT U910 ( .A(src_window[93]), .Y(DP_OP_422J2_124_3477_n2922) );
  INVX1_HVT U911 ( .A(src_window[92]), .Y(DP_OP_422J2_124_3477_n2923) );
  INVX1_HVT U912 ( .A(src_window[91]), .Y(DP_OP_422J2_124_3477_n2924) );
  INVX1_HVT U913 ( .A(src_window[89]), .Y(DP_OP_422J2_124_3477_n2926) );
  INVX1_HVT U914 ( .A(src_window[88]), .Y(DP_OP_422J2_124_3477_n2927) );
  INVX1_HVT U915 ( .A(conv_weight_box[19]), .Y(DP_OP_422J2_124_3477_n2928) );
  INVX1_HVT U916 ( .A(conv_weight_box[18]), .Y(DP_OP_422J2_124_3477_n2929) );
  INVX1_HVT U917 ( .A(conv_weight_box[17]), .Y(DP_OP_422J2_124_3477_n2930) );
  INVX1_HVT U918 ( .A(conv_weight_box[16]), .Y(DP_OP_422J2_124_3477_n2931) );
  INVX1_HVT U919 ( .A(src_window[79]), .Y(DP_OP_422J2_124_3477_n2964) );
  INVX1_HVT U920 ( .A(src_window[74]), .Y(DP_OP_422J2_124_3477_n2969) );
  INVX1_HVT U921 ( .A(src_window[73]), .Y(DP_OP_422J2_124_3477_n2970) );
  INVX1_HVT U922 ( .A(src_window[72]), .Y(DP_OP_422J2_124_3477_n2971) );
  INVX1_HVT U923 ( .A(conv_weight_box[11]), .Y(DP_OP_422J2_124_3477_n2972) );
  INVX1_HVT U924 ( .A(conv_weight_box[10]), .Y(DP_OP_422J2_124_3477_n2973) );
  INVX1_HVT U925 ( .A(conv_weight_box[9]), .Y(DP_OP_422J2_124_3477_n2974) );
  INVX1_HVT U926 ( .A(conv_weight_box[8]), .Y(DP_OP_422J2_124_3477_n2975) );
  INVX1_HVT U927 ( .A(src_window[63]), .Y(DP_OP_422J2_124_3477_n3006) );
  INVX1_HVT U928 ( .A(src_window[62]), .Y(DP_OP_422J2_124_3477_n3007) );
  INVX1_HVT U929 ( .A(src_window[61]), .Y(DP_OP_422J2_124_3477_n3008) );
  INVX1_HVT U930 ( .A(src_window[60]), .Y(DP_OP_422J2_124_3477_n3009) );
  INVX1_HVT U931 ( .A(src_window[59]), .Y(DP_OP_422J2_124_3477_n3010) );
  INVX1_HVT U932 ( .A(src_window[58]), .Y(DP_OP_422J2_124_3477_n3011) );
  INVX1_HVT U933 ( .A(src_window[57]), .Y(DP_OP_422J2_124_3477_n3012) );
  INVX1_HVT U934 ( .A(src_window[56]), .Y(DP_OP_422J2_124_3477_n3013) );
  INVX1_HVT U935 ( .A(conv_weight_box[2]), .Y(DP_OP_422J2_124_3477_n3015) );
  INVX1_HVT U936 ( .A(conv_weight_box[1]), .Y(DP_OP_422J2_124_3477_n3016) );
  INVX1_HVT U937 ( .A(conv_weight_box[0]), .Y(DP_OP_422J2_124_3477_n3017) );
  INVX1_HVT U938 ( .A(DP_OP_422J2_124_3477_n460), .Y(DP_OP_422J2_124_3477_n461) );
  INVX1_HVT U939 ( .A(DP_OP_422J2_124_3477_n770), .Y(DP_OP_422J2_124_3477_n771) );
  OR2X1_HVT U940 ( .A1(DP_OP_422J2_124_3477_n252), .A2(n421), .Y(n420) );
  OR2X1_HVT U941 ( .A1(n377), .A2(n391), .Y(n421) );
  OR2X1_HVT U942 ( .A1(DP_OP_422J2_124_3477_n258), .A2(
        DP_OP_422J2_124_3477_n257), .Y(n422) );
  OR2X1_HVT U943 ( .A1(DP_OP_422J2_124_3477_n262), .A2(
        DP_OP_422J2_124_3477_n261), .Y(n423) );
  OR2X1_HVT U944 ( .A1(DP_OP_422J2_124_3477_n264), .A2(
        DP_OP_422J2_124_3477_n263), .Y(n424) );
  OR2X1_HVT U945 ( .A1(DP_OP_422J2_124_3477_n268), .A2(
        DP_OP_422J2_124_3477_n267), .Y(n425) );
  OR2X1_HVT U946 ( .A1(DP_OP_422J2_124_3477_n971), .A2(
        DP_OP_422J2_124_3477_n969), .Y(n426) );
  OR2X1_HVT U947 ( .A1(DP_OP_422J2_124_3477_n1353), .A2(
        DP_OP_422J2_124_3477_n1351), .Y(n427) );
  OR2X1_HVT U948 ( .A1(DP_OP_422J2_124_3477_n1683), .A2(
        DP_OP_422J2_124_3477_n1681), .Y(n428) );
  OR2X1_HVT U949 ( .A1(DP_OP_422J2_124_3477_n272), .A2(
        DP_OP_422J2_124_3477_n271), .Y(n429) );
  OR2X1_HVT U950 ( .A1(DP_OP_422J2_124_3477_n276), .A2(
        DP_OP_422J2_124_3477_n275), .Y(n430) );
  INVX1_HVT U951 ( .A(DP_OP_422J2_124_3477_n288), .Y(DP_OP_422J2_124_3477_n289) );
  INVX1_HVT U952 ( .A(DP_OP_422J2_124_3477_n162), .Y(DP_OP_422J2_124_3477_n161) );
  INVX1_HVT U953 ( .A(conv_weight_box[3]), .Y(DP_OP_422J2_124_3477_n3014) );
  INVX1_HVT U954 ( .A(DP_OP_423J2_125_3477_n148), .Y(DP_OP_423J2_125_3477_n236) );
  INVX1_HVT U955 ( .A(DP_OP_423J2_125_3477_n152), .Y(DP_OP_423J2_125_3477_n158) );
  INVX1_HVT U956 ( .A(DP_OP_423J2_125_3477_n1678), .Y(
        DP_OP_423J2_125_3477_n1679) );
  INVX1_HVT U957 ( .A(DP_OP_423J2_125_3477_n183), .Y(DP_OP_423J2_125_3477_n182) );
  INVX1_HVT U958 ( .A(src_window[63]), .Y(DP_OP_423J2_125_3477_n1952) );
  INVX1_HVT U959 ( .A(src_window[58]), .Y(DP_OP_423J2_125_3477_n1957) );
  INVX1_HVT U960 ( .A(src_window[57]), .Y(DP_OP_423J2_125_3477_n1958) );
  INVX1_HVT U961 ( .A(conv_weight_box[5]), .Y(DP_OP_423J2_125_3477_n1962) );
  INVX1_HVT U962 ( .A(conv_weight_box[4]), .Y(DP_OP_423J2_125_3477_n1963) );
  INVX1_HVT U963 ( .A(src_window[78]), .Y(DP_OP_423J2_125_3477_n1997) );
  INVX1_HVT U964 ( .A(src_window[77]), .Y(DP_OP_423J2_125_3477_n1998) );
  INVX1_HVT U965 ( .A(src_window[75]), .Y(DP_OP_423J2_125_3477_n2000) );
  INVX1_HVT U966 ( .A(src_window[72]), .Y(DP_OP_423J2_125_3477_n2003) );
  INVX1_HVT U967 ( .A(conv_weight_box[15]), .Y(DP_OP_423J2_125_3477_n2004) );
  INVX1_HVT U968 ( .A(conv_weight_box[14]), .Y(DP_OP_423J2_125_3477_n2005) );
  INVX1_HVT U969 ( .A(conv_weight_box[13]), .Y(DP_OP_423J2_125_3477_n2006) );
  INVX1_HVT U970 ( .A(conv_weight_box[12]), .Y(DP_OP_423J2_125_3477_n2007) );
  INVX1_HVT U971 ( .A(src_window[103]), .Y(DP_OP_423J2_125_3477_n2040) );
  INVX1_HVT U972 ( .A(src_window[99]), .Y(DP_OP_423J2_125_3477_n2044) );
  INVX1_HVT U973 ( .A(conv_weight_box[23]), .Y(DP_OP_423J2_125_3477_n2048) );
  INVX1_HVT U974 ( .A(conv_weight_box[21]), .Y(DP_OP_423J2_125_3477_n2050) );
  INVX1_HVT U975 ( .A(src_window[119]), .Y(DP_OP_423J2_125_3477_n2084) );
  INVX1_HVT U976 ( .A(src_window[117]), .Y(DP_OP_423J2_125_3477_n2086) );
  INVX1_HVT U977 ( .A(src_window[116]), .Y(DP_OP_423J2_125_3477_n2087) );
  INVX1_HVT U978 ( .A(src_window[115]), .Y(DP_OP_423J2_125_3477_n2088) );
  INVX1_HVT U979 ( .A(conv_weight_box[31]), .Y(DP_OP_423J2_125_3477_n2092) );
  INVX1_HVT U980 ( .A(conv_weight_box[30]), .Y(DP_OP_423J2_125_3477_n2093) );
  INVX1_HVT U981 ( .A(src_window[135]), .Y(DP_OP_423J2_125_3477_n2128) );
  INVX1_HVT U982 ( .A(src_window[129]), .Y(DP_OP_423J2_125_3477_n2134) );
  INVX1_HVT U983 ( .A(src_window[128]), .Y(DP_OP_423J2_125_3477_n2135) );
  INVX1_HVT U984 ( .A(conv_weight_box[39]), .Y(DP_OP_423J2_125_3477_n2136) );
  INVX1_HVT U985 ( .A(conv_weight_box[37]), .Y(DP_OP_423J2_125_3477_n2138) );
  INVX1_HVT U986 ( .A(conv_weight_box[36]), .Y(DP_OP_423J2_125_3477_n2139) );
  INVX1_HVT U987 ( .A(src_window[159]), .Y(DP_OP_423J2_125_3477_n2172) );
  INVX1_HVT U988 ( .A(src_window[156]), .Y(DP_OP_423J2_125_3477_n2175) );
  INVX1_HVT U989 ( .A(src_window[153]), .Y(DP_OP_423J2_125_3477_n2178) );
  INVX1_HVT U990 ( .A(conv_weight_box[47]), .Y(DP_OP_423J2_125_3477_n2180) );
  INVX1_HVT U991 ( .A(conv_weight_box[46]), .Y(DP_OP_423J2_125_3477_n2181) );
  INVX1_HVT U992 ( .A(conv_weight_box[44]), .Y(DP_OP_423J2_125_3477_n2183) );
  INVX1_HVT U993 ( .A(src_window[174]), .Y(DP_OP_423J2_125_3477_n2217) );
  INVX1_HVT U994 ( .A(src_window[173]), .Y(DP_OP_423J2_125_3477_n2218) );
  INVX1_HVT U995 ( .A(src_window[172]), .Y(DP_OP_423J2_125_3477_n2219) );
  INVX1_HVT U996 ( .A(conv_weight_box[55]), .Y(DP_OP_423J2_125_3477_n2224) );
  INVX1_HVT U997 ( .A(conv_weight_box[54]), .Y(DP_OP_423J2_125_3477_n2225) );
  INVX1_HVT U998 ( .A(conv_weight_box[53]), .Y(DP_OP_423J2_125_3477_n2226) );
  INVX1_HVT U999 ( .A(src_window[199]), .Y(DP_OP_423J2_125_3477_n2260) );
  INVX1_HVT U1000 ( .A(src_window[198]), .Y(DP_OP_423J2_125_3477_n2261) );
  INVX1_HVT U1001 ( .A(src_window[197]), .Y(DP_OP_423J2_125_3477_n2262) );
  INVX1_HVT U1002 ( .A(src_window[196]), .Y(DP_OP_423J2_125_3477_n2263) );
  INVX1_HVT U1003 ( .A(src_window[194]), .Y(DP_OP_423J2_125_3477_n2265) );
  INVX1_HVT U1004 ( .A(src_window[193]), .Y(DP_OP_423J2_125_3477_n2266) );
  INVX1_HVT U1005 ( .A(src_window[192]), .Y(DP_OP_423J2_125_3477_n2267) );
  INVX1_HVT U1006 ( .A(conv_weight_box[63]), .Y(DP_OP_423J2_125_3477_n2268) );
  INVX1_HVT U1007 ( .A(conv_weight_box[61]), .Y(DP_OP_423J2_125_3477_n2270) );
  INVX1_HVT U1008 ( .A(src_window[215]), .Y(DP_OP_423J2_125_3477_n2304) );
  INVX1_HVT U1009 ( .A(src_window[214]), .Y(DP_OP_423J2_125_3477_n2305) );
  INVX1_HVT U1010 ( .A(src_window[212]), .Y(DP_OP_423J2_125_3477_n2307) );
  INVX1_HVT U1011 ( .A(src_window[211]), .Y(DP_OP_423J2_125_3477_n2308) );
  INVX1_HVT U1012 ( .A(src_window[208]), .Y(DP_OP_423J2_125_3477_n2311) );
  INVX1_HVT U1013 ( .A(conv_weight_box[71]), .Y(DP_OP_423J2_125_3477_n2312) );
  INVX1_HVT U1014 ( .A(conv_weight_box[70]), .Y(DP_OP_423J2_125_3477_n2313) );
  INVX1_HVT U1015 ( .A(conv_weight_box[69]), .Y(DP_OP_423J2_125_3477_n2314) );
  INVX1_HVT U1016 ( .A(conv_weight_box[68]), .Y(DP_OP_423J2_125_3477_n2315) );
  INVX1_HVT U1017 ( .A(src_window[231]), .Y(DP_OP_423J2_125_3477_n2348) );
  INVX1_HVT U1018 ( .A(src_window[229]), .Y(DP_OP_423J2_125_3477_n2350) );
  INVX1_HVT U1019 ( .A(src_window[228]), .Y(DP_OP_423J2_125_3477_n2351) );
  INVX1_HVT U1020 ( .A(src_window[226]), .Y(DP_OP_423J2_125_3477_n2353) );
  INVX1_HVT U1021 ( .A(src_window[225]), .Y(DP_OP_423J2_125_3477_n2354) );
  INVX1_HVT U1022 ( .A(src_window[224]), .Y(DP_OP_423J2_125_3477_n2355) );
  INVX1_HVT U1023 ( .A(conv_weight_box[79]), .Y(DP_OP_423J2_125_3477_n2356) );
  INVX1_HVT U1024 ( .A(conv_weight_box[78]), .Y(DP_OP_423J2_125_3477_n2357) );
  INVX1_HVT U1025 ( .A(conv_weight_box[77]), .Y(DP_OP_423J2_125_3477_n2358) );
  INVX1_HVT U1026 ( .A(conv_weight_box[76]), .Y(DP_OP_423J2_125_3477_n2359) );
  INVX1_HVT U1027 ( .A(src_window[251]), .Y(DP_OP_423J2_125_3477_n2396) );
  INVX1_HVT U1028 ( .A(src_window[250]), .Y(DP_OP_423J2_125_3477_n2397) );
  INVX1_HVT U1029 ( .A(src_window[249]), .Y(DP_OP_423J2_125_3477_n2398) );
  INVX1_HVT U1030 ( .A(DP_OP_423J2_125_3477_n175), .Y(
        DP_OP_423J2_125_3477_n240) );
  INVX1_HVT U1031 ( .A(conv_weight_box[87]), .Y(DP_OP_423J2_125_3477_n2400) );
  INVX1_HVT U1032 ( .A(conv_weight_box[86]), .Y(DP_OP_423J2_125_3477_n2401) );
  INVX1_HVT U1033 ( .A(conv_weight_box[85]), .Y(DP_OP_423J2_125_3477_n2402) );
  INVX1_HVT U1034 ( .A(conv_weight_box[84]), .Y(DP_OP_423J2_125_3477_n2403) );
  INVX1_HVT U1035 ( .A(src_window[271]), .Y(DP_OP_423J2_125_3477_n2436) );
  INVX1_HVT U1036 ( .A(src_window[270]), .Y(DP_OP_423J2_125_3477_n2437) );
  INVX1_HVT U1037 ( .A(src_window[268]), .Y(DP_OP_423J2_125_3477_n2439) );
  INVX1_HVT U1038 ( .A(src_window[266]), .Y(DP_OP_423J2_125_3477_n2441) );
  INVX1_HVT U1039 ( .A(src_window[265]), .Y(DP_OP_423J2_125_3477_n2442) );
  INVX1_HVT U1040 ( .A(conv_weight_box[95]), .Y(DP_OP_423J2_125_3477_n2444) );
  INVX1_HVT U1041 ( .A(conv_weight_box[94]), .Y(DP_OP_423J2_125_3477_n2445) );
  INVX1_HVT U1042 ( .A(conv_weight_box[93]), .Y(DP_OP_423J2_125_3477_n2446) );
  INVX1_HVT U1043 ( .A(src_window[278]), .Y(DP_OP_423J2_125_3477_n2481) );
  INVX1_HVT U1044 ( .A(src_window[277]), .Y(DP_OP_423J2_125_3477_n2482) );
  INVX1_HVT U1045 ( .A(src_window[275]), .Y(DP_OP_423J2_125_3477_n2484) );
  INVX1_HVT U1046 ( .A(src_window[272]), .Y(DP_OP_423J2_125_3477_n2487) );
  INVX1_HVT U1047 ( .A(conv_weight_box[99]), .Y(DP_OP_423J2_125_3477_n2488) );
  INVX1_HVT U1048 ( .A(conv_weight_box[98]), .Y(DP_OP_423J2_125_3477_n2489) );
  INVX1_HVT U1049 ( .A(conv_weight_box[97]), .Y(DP_OP_423J2_125_3477_n2490) );
  INVX1_HVT U1050 ( .A(conv_weight_box[96]), .Y(DP_OP_423J2_125_3477_n2491) );
  INVX1_HVT U1051 ( .A(src_window[262]), .Y(DP_OP_423J2_125_3477_n2525) );
  INVX1_HVT U1052 ( .A(src_window[261]), .Y(DP_OP_423J2_125_3477_n2526) );
  INVX1_HVT U1053 ( .A(src_window[260]), .Y(DP_OP_423J2_125_3477_n2527) );
  INVX1_HVT U1054 ( .A(src_window[259]), .Y(DP_OP_423J2_125_3477_n2528) );
  INVX1_HVT U1055 ( .A(src_window[258]), .Y(DP_OP_423J2_125_3477_n2529) );
  INVX1_HVT U1056 ( .A(DP_OP_423J2_125_3477_n252), .Y(
        DP_OP_423J2_125_3477_n253) );
  INVX1_HVT U1057 ( .A(src_window[257]), .Y(DP_OP_423J2_125_3477_n2530) );
  INVX1_HVT U1058 ( .A(src_window[256]), .Y(DP_OP_423J2_125_3477_n2531) );
  INVX1_HVT U1059 ( .A(conv_weight_box[91]), .Y(DP_OP_423J2_125_3477_n2532) );
  INVX1_HVT U1060 ( .A(conv_weight_box[90]), .Y(DP_OP_423J2_125_3477_n2533) );
  INVX1_HVT U1061 ( .A(conv_weight_box[89]), .Y(DP_OP_423J2_125_3477_n2534) );
  INVX1_HVT U1062 ( .A(conv_weight_box[88]), .Y(DP_OP_423J2_125_3477_n2535) );
  INVX1_HVT U1063 ( .A(DP_OP_423J2_125_3477_n254), .Y(
        DP_OP_423J2_125_3477_n255) );
  INVX1_HVT U1064 ( .A(src_window[247]), .Y(DP_OP_423J2_125_3477_n2568) );
  INVX1_HVT U1065 ( .A(src_window[246]), .Y(DP_OP_423J2_125_3477_n2569) );
  INVX1_HVT U1066 ( .A(DP_OP_423J2_125_3477_n256), .Y(
        DP_OP_423J2_125_3477_n257) );
  INVX1_HVT U1067 ( .A(src_window[245]), .Y(DP_OP_423J2_125_3477_n2570) );
  INVX1_HVT U1068 ( .A(src_window[244]), .Y(DP_OP_423J2_125_3477_n2571) );
  INVX1_HVT U1069 ( .A(src_window[243]), .Y(DP_OP_423J2_125_3477_n2572) );
  INVX1_HVT U1070 ( .A(src_window[242]), .Y(DP_OP_423J2_125_3477_n2573) );
  INVX1_HVT U1071 ( .A(src_window[241]), .Y(DP_OP_423J2_125_3477_n2574) );
  INVX1_HVT U1072 ( .A(src_window[240]), .Y(DP_OP_423J2_125_3477_n2575) );
  INVX1_HVT U1073 ( .A(conv_weight_box[83]), .Y(DP_OP_423J2_125_3477_n2576) );
  INVX1_HVT U1074 ( .A(conv_weight_box[82]), .Y(DP_OP_423J2_125_3477_n2577) );
  INVX1_HVT U1075 ( .A(conv_weight_box[80]), .Y(DP_OP_423J2_125_3477_n2579) );
  INVX1_HVT U1076 ( .A(DP_OP_423J2_125_3477_n258), .Y(
        DP_OP_423J2_125_3477_n259) );
  INVX1_HVT U1077 ( .A(DP_OP_423J2_125_3477_n260), .Y(
        DP_OP_423J2_125_3477_n261) );
  INVX1_HVT U1078 ( .A(src_window[223]), .Y(DP_OP_423J2_125_3477_n2612) );
  INVX1_HVT U1079 ( .A(src_window[222]), .Y(DP_OP_423J2_125_3477_n2613) );
  INVX1_HVT U1080 ( .A(src_window[218]), .Y(DP_OP_423J2_125_3477_n2617) );
  INVX1_HVT U1081 ( .A(src_window[216]), .Y(DP_OP_423J2_125_3477_n2619) );
  INVX1_HVT U1082 ( .A(conv_weight_box[74]), .Y(DP_OP_423J2_125_3477_n2621) );
  INVX1_HVT U1083 ( .A(conv_weight_box[72]), .Y(DP_OP_423J2_125_3477_n2623) );
  INVX1_HVT U1084 ( .A(DP_OP_423J2_125_3477_n262), .Y(
        DP_OP_423J2_125_3477_n263) );
  INVX1_HVT U1085 ( .A(DP_OP_423J2_125_3477_n264), .Y(
        DP_OP_423J2_125_3477_n265) );
  INVX1_HVT U1086 ( .A(src_window[207]), .Y(DP_OP_423J2_125_3477_n2656) );
  INVX1_HVT U1087 ( .A(src_window[205]), .Y(DP_OP_423J2_125_3477_n2658) );
  INVX1_HVT U1088 ( .A(src_window[204]), .Y(DP_OP_423J2_125_3477_n2659) );
  INVX1_HVT U1089 ( .A(src_window[201]), .Y(DP_OP_423J2_125_3477_n2662) );
  INVX1_HVT U1090 ( .A(src_window[200]), .Y(DP_OP_423J2_125_3477_n2663) );
  INVX1_HVT U1091 ( .A(conv_weight_box[67]), .Y(DP_OP_423J2_125_3477_n2664) );
  INVX1_HVT U1092 ( .A(conv_weight_box[66]), .Y(DP_OP_423J2_125_3477_n2665) );
  INVX1_HVT U1093 ( .A(conv_weight_box[64]), .Y(DP_OP_423J2_125_3477_n2667) );
  INVX1_HVT U1094 ( .A(DP_OP_423J2_125_3477_n266), .Y(
        DP_OP_423J2_125_3477_n267) );
  INVX1_HVT U1095 ( .A(DP_OP_423J2_125_3477_n268), .Y(
        DP_OP_423J2_125_3477_n269) );
  INVX1_HVT U1096 ( .A(src_window[183]), .Y(DP_OP_423J2_125_3477_n2700) );
  INVX1_HVT U1097 ( .A(src_window[181]), .Y(DP_OP_423J2_125_3477_n2702) );
  INVX1_HVT U1098 ( .A(src_window[178]), .Y(DP_OP_423J2_125_3477_n2705) );
  INVX1_HVT U1099 ( .A(src_window[176]), .Y(DP_OP_423J2_125_3477_n2707) );
  INVX1_HVT U1100 ( .A(conv_weight_box[59]), .Y(DP_OP_423J2_125_3477_n2708) );
  INVX1_HVT U1101 ( .A(conv_weight_box[58]), .Y(DP_OP_423J2_125_3477_n2709) );
  INVX1_HVT U1102 ( .A(DP_OP_423J2_125_3477_n270), .Y(
        DP_OP_423J2_125_3477_n271) );
  INVX1_HVT U1103 ( .A(conv_weight_box[57]), .Y(DP_OP_423J2_125_3477_n2710) );
  INVX1_HVT U1104 ( .A(DP_OP_423J2_125_3477_n272), .Y(
        DP_OP_423J2_125_3477_n273) );
  INVX1_HVT U1105 ( .A(src_window[166]), .Y(DP_OP_423J2_125_3477_n2745) );
  INVX1_HVT U1106 ( .A(src_window[165]), .Y(DP_OP_423J2_125_3477_n2746) );
  INVX1_HVT U1107 ( .A(src_window[164]), .Y(DP_OP_423J2_125_3477_n2747) );
  INVX1_HVT U1108 ( .A(src_window[163]), .Y(DP_OP_423J2_125_3477_n2748) );
  INVX1_HVT U1109 ( .A(src_window[162]), .Y(DP_OP_423J2_125_3477_n2749) );
  INVX1_HVT U1110 ( .A(DP_OP_423J2_125_3477_n274), .Y(
        DP_OP_423J2_125_3477_n275) );
  INVX1_HVT U1111 ( .A(src_window[161]), .Y(DP_OP_423J2_125_3477_n2750) );
  INVX1_HVT U1112 ( .A(conv_weight_box[51]), .Y(DP_OP_423J2_125_3477_n2752) );
  INVX1_HVT U1113 ( .A(conv_weight_box[50]), .Y(DP_OP_423J2_125_3477_n2753) );
  INVX1_HVT U1114 ( .A(conv_weight_box[49]), .Y(DP_OP_423J2_125_3477_n2754) );
  INVX1_HVT U1115 ( .A(conv_weight_box[48]), .Y(DP_OP_423J2_125_3477_n2755) );
  INVX1_HVT U1116 ( .A(DP_OP_423J2_125_3477_n276), .Y(
        DP_OP_423J2_125_3477_n277) );
  INVX1_HVT U1117 ( .A(DP_OP_423J2_125_3477_n278), .Y(
        DP_OP_423J2_125_3477_n279) );
  INVX1_HVT U1118 ( .A(src_window[149]), .Y(DP_OP_423J2_125_3477_n2790) );
  INVX1_HVT U1119 ( .A(src_window[148]), .Y(DP_OP_423J2_125_3477_n2791) );
  INVX1_HVT U1120 ( .A(src_window[146]), .Y(DP_OP_423J2_125_3477_n2793) );
  INVX1_HVT U1121 ( .A(src_window[145]), .Y(DP_OP_423J2_125_3477_n2794) );
  INVX1_HVT U1122 ( .A(src_window[144]), .Y(DP_OP_423J2_125_3477_n2795) );
  INVX1_HVT U1123 ( .A(conv_weight_box[43]), .Y(DP_OP_423J2_125_3477_n2796) );
  INVX1_HVT U1124 ( .A(conv_weight_box[41]), .Y(DP_OP_423J2_125_3477_n2798) );
  INVX1_HVT U1125 ( .A(DP_OP_423J2_125_3477_n280), .Y(
        DP_OP_423J2_125_3477_n281) );
  INVX1_HVT U1126 ( .A(src_window[125]), .Y(DP_OP_423J2_125_3477_n2834) );
  INVX1_HVT U1127 ( .A(src_window[122]), .Y(DP_OP_423J2_125_3477_n2837) );
  INVX1_HVT U1128 ( .A(conv_weight_box[35]), .Y(DP_OP_423J2_125_3477_n2840) );
  INVX1_HVT U1129 ( .A(conv_weight_box[34]), .Y(DP_OP_423J2_125_3477_n2841) );
  INVX1_HVT U1130 ( .A(conv_weight_box[33]), .Y(DP_OP_423J2_125_3477_n2842) );
  INVX1_HVT U1131 ( .A(conv_weight_box[32]), .Y(DP_OP_423J2_125_3477_n2843) );
  INVX1_HVT U1132 ( .A(src_window[110]), .Y(DP_OP_423J2_125_3477_n2877) );
  INVX1_HVT U1133 ( .A(src_window[109]), .Y(DP_OP_423J2_125_3477_n2878) );
  INVX1_HVT U1134 ( .A(src_window[107]), .Y(DP_OP_423J2_125_3477_n2880) );
  INVX1_HVT U1135 ( .A(conv_weight_box[27]), .Y(DP_OP_423J2_125_3477_n2884) );
  INVX1_HVT U1136 ( .A(conv_weight_box[26]), .Y(DP_OP_423J2_125_3477_n2885) );
  INVX1_HVT U1137 ( .A(conv_weight_box[25]), .Y(DP_OP_423J2_125_3477_n2886) );
  INVX1_HVT U1138 ( .A(src_window[87]), .Y(DP_OP_423J2_125_3477_n2920) );
  INVX1_HVT U1139 ( .A(src_window[86]), .Y(DP_OP_423J2_125_3477_n2921) );
  INVX1_HVT U1140 ( .A(src_window[85]), .Y(DP_OP_423J2_125_3477_n2922) );
  INVX1_HVT U1141 ( .A(src_window[84]), .Y(DP_OP_423J2_125_3477_n2923) );
  INVX1_HVT U1142 ( .A(src_window[83]), .Y(DP_OP_423J2_125_3477_n2924) );
  INVX1_HVT U1143 ( .A(src_window[81]), .Y(DP_OP_423J2_125_3477_n2926) );
  INVX1_HVT U1144 ( .A(src_window[80]), .Y(DP_OP_423J2_125_3477_n2927) );
  INVX1_HVT U1145 ( .A(conv_weight_box[19]), .Y(DP_OP_423J2_125_3477_n2928) );
  INVX1_HVT U1146 ( .A(conv_weight_box[18]), .Y(DP_OP_423J2_125_3477_n2929) );
  INVX1_HVT U1147 ( .A(conv_weight_box[17]), .Y(DP_OP_423J2_125_3477_n2930) );
  INVX1_HVT U1148 ( .A(conv_weight_box[16]), .Y(DP_OP_423J2_125_3477_n2931) );
  INVX1_HVT U1149 ( .A(src_window[71]), .Y(DP_OP_423J2_125_3477_n2964) );
  INVX1_HVT U1150 ( .A(src_window[68]), .Y(DP_OP_423J2_125_3477_n2967) );
  INVX1_HVT U1151 ( .A(src_window[66]), .Y(DP_OP_423J2_125_3477_n2969) );
  INVX1_HVT U1152 ( .A(src_window[65]), .Y(DP_OP_423J2_125_3477_n2970) );
  INVX1_HVT U1153 ( .A(src_window[64]), .Y(DP_OP_423J2_125_3477_n2971) );
  INVX1_HVT U1154 ( .A(conv_weight_box[11]), .Y(DP_OP_423J2_125_3477_n2972) );
  INVX1_HVT U1155 ( .A(conv_weight_box[10]), .Y(DP_OP_423J2_125_3477_n2973) );
  INVX1_HVT U1156 ( .A(conv_weight_box[9]), .Y(DP_OP_423J2_125_3477_n2974) );
  INVX1_HVT U1157 ( .A(src_window[55]), .Y(DP_OP_423J2_125_3477_n3006) );
  INVX1_HVT U1158 ( .A(src_window[54]), .Y(DP_OP_423J2_125_3477_n3007) );
  INVX1_HVT U1159 ( .A(src_window[53]), .Y(DP_OP_423J2_125_3477_n3008) );
  INVX1_HVT U1160 ( .A(src_window[52]), .Y(DP_OP_423J2_125_3477_n3009) );
  INVX1_HVT U1161 ( .A(src_window[51]), .Y(DP_OP_423J2_125_3477_n3010) );
  INVX1_HVT U1162 ( .A(src_window[50]), .Y(DP_OP_423J2_125_3477_n3011) );
  INVX1_HVT U1163 ( .A(src_window[49]), .Y(DP_OP_423J2_125_3477_n3012) );
  INVX1_HVT U1164 ( .A(conv_weight_box[1]), .Y(DP_OP_423J2_125_3477_n3016) );
  INVX1_HVT U1165 ( .A(conv_weight_box[0]), .Y(DP_OP_423J2_125_3477_n3017) );
  INVX1_HVT U1166 ( .A(DP_OP_423J2_125_3477_n460), .Y(
        DP_OP_423J2_125_3477_n461) );
  INVX1_HVT U1167 ( .A(DP_OP_423J2_125_3477_n770), .Y(
        DP_OP_423J2_125_3477_n771) );
  OR2X1_HVT U1168 ( .A1(DP_OP_423J2_125_3477_n252), .A2(n441), .Y(n431) );
  OR2X1_HVT U1169 ( .A1(DP_OP_423J2_125_3477_n258), .A2(
        DP_OP_423J2_125_3477_n257), .Y(n432) );
  OR2X1_HVT U1170 ( .A1(DP_OP_423J2_125_3477_n262), .A2(
        DP_OP_423J2_125_3477_n261), .Y(n433) );
  OR2X1_HVT U1171 ( .A1(DP_OP_423J2_125_3477_n264), .A2(
        DP_OP_423J2_125_3477_n263), .Y(n434) );
  OR2X1_HVT U1172 ( .A1(DP_OP_423J2_125_3477_n268), .A2(
        DP_OP_423J2_125_3477_n267), .Y(n435) );
  OR2X1_HVT U1173 ( .A1(DP_OP_423J2_125_3477_n971), .A2(
        DP_OP_423J2_125_3477_n969), .Y(n436) );
  OR2X1_HVT U1174 ( .A1(DP_OP_423J2_125_3477_n1353), .A2(
        DP_OP_423J2_125_3477_n1351), .Y(n437) );
  OR2X1_HVT U1175 ( .A1(DP_OP_423J2_125_3477_n1683), .A2(
        DP_OP_423J2_125_3477_n1681), .Y(n438) );
  OR2X1_HVT U1176 ( .A1(DP_OP_423J2_125_3477_n272), .A2(
        DP_OP_423J2_125_3477_n271), .Y(n439) );
  OR2X1_HVT U1177 ( .A1(DP_OP_423J2_125_3477_n276), .A2(
        DP_OP_423J2_125_3477_n275), .Y(n440) );
  OR2X1_HVT U1178 ( .A1(n529), .A2(n386), .Y(n441) );
  AOI21X2_HVT U1179 ( .A1(DP_OP_423J2_125_3477_n162), .A2(
        DP_OP_423J2_125_3477_n135), .A3(DP_OP_423J2_125_3477_n136), .Y(
        DP_OP_423J2_125_3477_n3) );
  INVX1_HVT U1180 ( .A(DP_OP_423J2_125_3477_n288), .Y(
        DP_OP_423J2_125_3477_n289) );
  INVX1_HVT U1181 ( .A(DP_OP_423J2_125_3477_n162), .Y(
        DP_OP_423J2_125_3477_n161) );
  INVX1_HVT U1182 ( .A(conv_weight_box[7]), .Y(DP_OP_423J2_125_3477_n1960) );
  INVX1_HVT U1183 ( .A(conv_weight_box[3]), .Y(DP_OP_423J2_125_3477_n3014) );
  INVX1_HVT U1184 ( .A(DP_OP_424J2_126_3477_n148), .Y(
        DP_OP_424J2_126_3477_n236) );
  INVX1_HVT U1185 ( .A(DP_OP_424J2_126_3477_n152), .Y(
        DP_OP_424J2_126_3477_n158) );
  INVX1_HVT U1186 ( .A(DP_OP_424J2_126_3477_n1678), .Y(
        DP_OP_424J2_126_3477_n1679) );
  INVX1_HVT U1187 ( .A(DP_OP_424J2_126_3477_n183), .Y(
        DP_OP_424J2_126_3477_n182) );
  INVX1_HVT U1188 ( .A(src_window[21]), .Y(DP_OP_424J2_126_3477_n1954) );
  INVX1_HVT U1189 ( .A(src_window[19]), .Y(DP_OP_424J2_126_3477_n1956) );
  INVX1_HVT U1190 ( .A(src_window[18]), .Y(DP_OP_424J2_126_3477_n1957) );
  INVX1_HVT U1191 ( .A(src_window[17]), .Y(DP_OP_424J2_126_3477_n1958) );
  INVX1_HVT U1192 ( .A(conv_weight_box[6]), .Y(DP_OP_424J2_126_3477_n1961) );
  INVX1_HVT U1193 ( .A(conv_weight_box[5]), .Y(DP_OP_424J2_126_3477_n1962) );
  INVX1_HVT U1194 ( .A(src_window[34]), .Y(DP_OP_424J2_126_3477_n2001) );
  INVX1_HVT U1195 ( .A(src_window[59]), .Y(DP_OP_424J2_126_3477_n2044) );
  INVX1_HVT U1196 ( .A(src_window[56]), .Y(DP_OP_424J2_126_3477_n2047) );
  INVX1_HVT U1197 ( .A(conv_weight_box[22]), .Y(DP_OP_424J2_126_3477_n2049) );
  INVX1_HVT U1198 ( .A(conv_weight_box[20]), .Y(DP_OP_424J2_126_3477_n2051) );
  INVX1_HVT U1199 ( .A(src_window[79]), .Y(DP_OP_424J2_126_3477_n2084) );
  INVX1_HVT U1200 ( .A(src_window[76]), .Y(DP_OP_424J2_126_3477_n2087) );
  INVX1_HVT U1201 ( .A(src_window[75]), .Y(DP_OP_424J2_126_3477_n2088) );
  INVX1_HVT U1202 ( .A(src_window[73]), .Y(DP_OP_424J2_126_3477_n2090) );
  INVX1_HVT U1203 ( .A(conv_weight_box[29]), .Y(DP_OP_424J2_126_3477_n2094) );
  INVX1_HVT U1204 ( .A(conv_weight_box[28]), .Y(DP_OP_424J2_126_3477_n2095) );
  INVX1_HVT U1205 ( .A(src_window[95]), .Y(DP_OP_424J2_126_3477_n2128) );
  INVX1_HVT U1206 ( .A(src_window[90]), .Y(DP_OP_424J2_126_3477_n2133) );
  INVX1_HVT U1207 ( .A(conv_weight_box[38]), .Y(DP_OP_424J2_126_3477_n2137) );
  INVX1_HVT U1208 ( .A(src_window[119]), .Y(DP_OP_424J2_126_3477_n2172) );
  INVX1_HVT U1209 ( .A(src_window[114]), .Y(DP_OP_424J2_126_3477_n2177) );
  INVX1_HVT U1210 ( .A(src_window[113]), .Y(DP_OP_424J2_126_3477_n2178) );
  INVX1_HVT U1211 ( .A(src_window[112]), .Y(DP_OP_424J2_126_3477_n2179) );
  INVX1_HVT U1212 ( .A(conv_weight_box[45]), .Y(DP_OP_424J2_126_3477_n2182) );
  INVX1_HVT U1213 ( .A(conv_weight_box[44]), .Y(DP_OP_424J2_126_3477_n2183) );
  INVX1_HVT U1214 ( .A(src_window[134]), .Y(DP_OP_424J2_126_3477_n2217) );
  INVX1_HVT U1215 ( .A(src_window[133]), .Y(DP_OP_424J2_126_3477_n2218) );
  INVX1_HVT U1216 ( .A(src_window[132]), .Y(DP_OP_424J2_126_3477_n2219) );
  INVX1_HVT U1217 ( .A(src_window[131]), .Y(DP_OP_424J2_126_3477_n2220) );
  INVX1_HVT U1218 ( .A(conv_weight_box[54]), .Y(DP_OP_424J2_126_3477_n2225) );
  INVX1_HVT U1219 ( .A(conv_weight_box[53]), .Y(DP_OP_424J2_126_3477_n2226) );
  INVX1_HVT U1220 ( .A(conv_weight_box[52]), .Y(DP_OP_424J2_126_3477_n2227) );
  INVX1_HVT U1221 ( .A(src_window[159]), .Y(DP_OP_424J2_126_3477_n2260) );
  INVX1_HVT U1222 ( .A(src_window[158]), .Y(DP_OP_424J2_126_3477_n2261) );
  INVX1_HVT U1223 ( .A(src_window[155]), .Y(DP_OP_424J2_126_3477_n2264) );
  INVX1_HVT U1224 ( .A(src_window[154]), .Y(DP_OP_424J2_126_3477_n2265) );
  INVX1_HVT U1225 ( .A(conv_weight_box[62]), .Y(DP_OP_424J2_126_3477_n2269) );
  INVX1_HVT U1226 ( .A(conv_weight_box[61]), .Y(DP_OP_424J2_126_3477_n2270) );
  INVX1_HVT U1227 ( .A(conv_weight_box[60]), .Y(DP_OP_424J2_126_3477_n2271) );
  INVX1_HVT U1228 ( .A(src_window[175]), .Y(DP_OP_424J2_126_3477_n2304) );
  INVX1_HVT U1229 ( .A(src_window[171]), .Y(DP_OP_424J2_126_3477_n2308) );
  INVX1_HVT U1230 ( .A(src_window[169]), .Y(DP_OP_424J2_126_3477_n2310) );
  INVX1_HVT U1231 ( .A(conv_weight_box[69]), .Y(DP_OP_424J2_126_3477_n2314) );
  INVX1_HVT U1232 ( .A(conv_weight_box[68]), .Y(DP_OP_424J2_126_3477_n2315) );
  INVX1_HVT U1233 ( .A(src_window[188]), .Y(DP_OP_424J2_126_3477_n2351) );
  INVX1_HVT U1234 ( .A(src_window[186]), .Y(DP_OP_424J2_126_3477_n2353) );
  INVX1_HVT U1235 ( .A(src_window[185]), .Y(DP_OP_424J2_126_3477_n2354) );
  INVX1_HVT U1236 ( .A(conv_weight_box[78]), .Y(DP_OP_424J2_126_3477_n2357) );
  INVX1_HVT U1237 ( .A(conv_weight_box[77]), .Y(DP_OP_424J2_126_3477_n2358) );
  INVX1_HVT U1238 ( .A(src_window[210]), .Y(DP_OP_424J2_126_3477_n2397) );
  INVX1_HVT U1239 ( .A(DP_OP_424J2_126_3477_n175), .Y(
        DP_OP_424J2_126_3477_n240) );
  INVX1_HVT U1240 ( .A(conv_weight_box[86]), .Y(DP_OP_424J2_126_3477_n2401) );
  INVX1_HVT U1241 ( .A(conv_weight_box[85]), .Y(DP_OP_424J2_126_3477_n2402) );
  INVX1_HVT U1242 ( .A(src_window[228]), .Y(DP_OP_424J2_126_3477_n2439) );
  INVX1_HVT U1243 ( .A(src_window[225]), .Y(DP_OP_424J2_126_3477_n2442) );
  INVX1_HVT U1244 ( .A(conv_weight_box[95]), .Y(DP_OP_424J2_126_3477_n2444) );
  INVX1_HVT U1245 ( .A(conv_weight_box[94]), .Y(DP_OP_424J2_126_3477_n2445) );
  INVX1_HVT U1246 ( .A(conv_weight_box[93]), .Y(DP_OP_424J2_126_3477_n2446) );
  INVX1_HVT U1247 ( .A(conv_weight_box[92]), .Y(DP_OP_424J2_126_3477_n2447) );
  INVX1_HVT U1248 ( .A(src_window[238]), .Y(DP_OP_424J2_126_3477_n2481) );
  INVX1_HVT U1249 ( .A(src_window[237]), .Y(DP_OP_424J2_126_3477_n2482) );
  INVX1_HVT U1250 ( .A(src_window[235]), .Y(DP_OP_424J2_126_3477_n2484) );
  INVX1_HVT U1251 ( .A(conv_weight_box[99]), .Y(DP_OP_424J2_126_3477_n2488) );
  INVX1_HVT U1252 ( .A(conv_weight_box[98]), .Y(DP_OP_424J2_126_3477_n2489) );
  INVX1_HVT U1253 ( .A(src_window[221]), .Y(DP_OP_424J2_126_3477_n2526) );
  INVX1_HVT U1254 ( .A(src_window[219]), .Y(DP_OP_424J2_126_3477_n2528) );
  INVX1_HVT U1255 ( .A(DP_OP_424J2_126_3477_n252), .Y(
        DP_OP_424J2_126_3477_n253) );
  INVX1_HVT U1256 ( .A(src_window[217]), .Y(DP_OP_424J2_126_3477_n2530) );
  INVX1_HVT U1257 ( .A(conv_weight_box[91]), .Y(DP_OP_424J2_126_3477_n2532) );
  INVX1_HVT U1258 ( .A(conv_weight_box[90]), .Y(DP_OP_424J2_126_3477_n2533) );
  INVX1_HVT U1259 ( .A(DP_OP_424J2_126_3477_n254), .Y(
        DP_OP_424J2_126_3477_n255) );
  INVX1_HVT U1260 ( .A(src_window[206]), .Y(DP_OP_424J2_126_3477_n2569) );
  INVX1_HVT U1261 ( .A(DP_OP_424J2_126_3477_n256), .Y(
        DP_OP_424J2_126_3477_n257) );
  INVX1_HVT U1262 ( .A(src_window[203]), .Y(DP_OP_424J2_126_3477_n2572) );
  INVX1_HVT U1263 ( .A(conv_weight_box[81]), .Y(DP_OP_424J2_126_3477_n2578) );
  INVX1_HVT U1264 ( .A(DP_OP_424J2_126_3477_n258), .Y(
        DP_OP_424J2_126_3477_n259) );
  INVX1_HVT U1265 ( .A(DP_OP_424J2_126_3477_n260), .Y(
        DP_OP_424J2_126_3477_n261) );
  INVX1_HVT U1266 ( .A(src_window[183]), .Y(DP_OP_424J2_126_3477_n2612) );
  INVX1_HVT U1267 ( .A(src_window[182]), .Y(DP_OP_424J2_126_3477_n2613) );
  INVX1_HVT U1268 ( .A(src_window[179]), .Y(DP_OP_424J2_126_3477_n2616) );
  INVX1_HVT U1269 ( .A(src_window[177]), .Y(DP_OP_424J2_126_3477_n2618) );
  INVX1_HVT U1270 ( .A(conv_weight_box[75]), .Y(DP_OP_424J2_126_3477_n2620) );
  INVX1_HVT U1271 ( .A(conv_weight_box[73]), .Y(DP_OP_424J2_126_3477_n2622) );
  INVX1_HVT U1272 ( .A(conv_weight_box[72]), .Y(DP_OP_424J2_126_3477_n2623) );
  INVX1_HVT U1273 ( .A(DP_OP_424J2_126_3477_n262), .Y(
        DP_OP_424J2_126_3477_n263) );
  INVX1_HVT U1274 ( .A(DP_OP_424J2_126_3477_n264), .Y(
        DP_OP_424J2_126_3477_n265) );
  INVX1_HVT U1275 ( .A(src_window[165]), .Y(DP_OP_424J2_126_3477_n2658) );
  INVX1_HVT U1276 ( .A(src_window[160]), .Y(DP_OP_424J2_126_3477_n2663) );
  INVX1_HVT U1277 ( .A(conv_weight_box[66]), .Y(DP_OP_424J2_126_3477_n2665) );
  INVX1_HVT U1278 ( .A(conv_weight_box[65]), .Y(DP_OP_424J2_126_3477_n2666) );
  INVX1_HVT U1279 ( .A(DP_OP_424J2_126_3477_n266), .Y(
        DP_OP_424J2_126_3477_n267) );
  INVX1_HVT U1280 ( .A(DP_OP_424J2_126_3477_n268), .Y(
        DP_OP_424J2_126_3477_n269) );
  INVX1_HVT U1281 ( .A(src_window[143]), .Y(DP_OP_424J2_126_3477_n2700) );
  INVX1_HVT U1282 ( .A(src_window[140]), .Y(DP_OP_424J2_126_3477_n2703) );
  INVX1_HVT U1283 ( .A(src_window[138]), .Y(DP_OP_424J2_126_3477_n2705) );
  INVX1_HVT U1284 ( .A(DP_OP_424J2_126_3477_n270), .Y(
        DP_OP_424J2_126_3477_n271) );
  INVX1_HVT U1285 ( .A(conv_weight_box[56]), .Y(DP_OP_424J2_126_3477_n2711) );
  INVX1_HVT U1286 ( .A(DP_OP_424J2_126_3477_n272), .Y(
        DP_OP_424J2_126_3477_n273) );
  INVX1_HVT U1287 ( .A(src_window[126]), .Y(DP_OP_424J2_126_3477_n2745) );
  INVX1_HVT U1288 ( .A(src_window[124]), .Y(DP_OP_424J2_126_3477_n2747) );
  INVX1_HVT U1289 ( .A(src_window[122]), .Y(DP_OP_424J2_126_3477_n2749) );
  INVX1_HVT U1290 ( .A(DP_OP_424J2_126_3477_n274), .Y(
        DP_OP_424J2_126_3477_n275) );
  INVX1_HVT U1291 ( .A(src_window[121]), .Y(DP_OP_424J2_126_3477_n2750) );
  INVX1_HVT U1292 ( .A(src_window[120]), .Y(DP_OP_424J2_126_3477_n2751) );
  INVX1_HVT U1293 ( .A(conv_weight_box[50]), .Y(DP_OP_424J2_126_3477_n2753) );
  INVX1_HVT U1294 ( .A(conv_weight_box[48]), .Y(DP_OP_424J2_126_3477_n2755) );
  INVX1_HVT U1295 ( .A(DP_OP_424J2_126_3477_n276), .Y(
        DP_OP_424J2_126_3477_n277) );
  INVX1_HVT U1296 ( .A(src_window[110]), .Y(DP_OP_424J2_126_3477_n2789) );
  INVX1_HVT U1297 ( .A(DP_OP_424J2_126_3477_n278), .Y(
        DP_OP_424J2_126_3477_n279) );
  INVX1_HVT U1298 ( .A(src_window[109]), .Y(DP_OP_424J2_126_3477_n2790) );
  INVX1_HVT U1299 ( .A(src_window[108]), .Y(DP_OP_424J2_126_3477_n2791) );
  INVX1_HVT U1300 ( .A(src_window[106]), .Y(DP_OP_424J2_126_3477_n2793) );
  INVX1_HVT U1301 ( .A(src_window[105]), .Y(DP_OP_424J2_126_3477_n2794) );
  INVX1_HVT U1302 ( .A(src_window[104]), .Y(DP_OP_424J2_126_3477_n2795) );
  INVX1_HVT U1303 ( .A(conv_weight_box[42]), .Y(DP_OP_424J2_126_3477_n2797) );
  INVX1_HVT U1304 ( .A(conv_weight_box[40]), .Y(DP_OP_424J2_126_3477_n2799) );
  INVX1_HVT U1305 ( .A(DP_OP_424J2_126_3477_n280), .Y(
        DP_OP_424J2_126_3477_n281) );
  INVX1_HVT U1306 ( .A(src_window[86]), .Y(DP_OP_424J2_126_3477_n2833) );
  INVX1_HVT U1307 ( .A(src_window[85]), .Y(DP_OP_424J2_126_3477_n2834) );
  INVX1_HVT U1308 ( .A(src_window[84]), .Y(DP_OP_424J2_126_3477_n2835) );
  INVX1_HVT U1309 ( .A(src_window[82]), .Y(DP_OP_424J2_126_3477_n2837) );
  INVX1_HVT U1310 ( .A(conv_weight_box[34]), .Y(DP_OP_424J2_126_3477_n2841) );
  INVX1_HVT U1311 ( .A(src_window[70]), .Y(DP_OP_424J2_126_3477_n2877) );
  INVX1_HVT U1312 ( .A(src_window[69]), .Y(DP_OP_424J2_126_3477_n2878) );
  INVX1_HVT U1313 ( .A(src_window[67]), .Y(DP_OP_424J2_126_3477_n2880) );
  INVX1_HVT U1314 ( .A(src_window[64]), .Y(DP_OP_424J2_126_3477_n2883) );
  INVX1_HVT U1315 ( .A(conv_weight_box[26]), .Y(DP_OP_424J2_126_3477_n2885) );
  INVX1_HVT U1316 ( .A(conv_weight_box[25]), .Y(DP_OP_424J2_126_3477_n2886) );
  INVX1_HVT U1317 ( .A(conv_weight_box[24]), .Y(DP_OP_424J2_126_3477_n2887) );
  INVX1_HVT U1318 ( .A(src_window[47]), .Y(DP_OP_424J2_126_3477_n2920) );
  INVX1_HVT U1319 ( .A(src_window[46]), .Y(DP_OP_424J2_126_3477_n2921) );
  INVX1_HVT U1320 ( .A(src_window[45]), .Y(DP_OP_424J2_126_3477_n2922) );
  INVX1_HVT U1321 ( .A(src_window[44]), .Y(DP_OP_424J2_126_3477_n2923) );
  INVX1_HVT U1322 ( .A(src_window[43]), .Y(DP_OP_424J2_126_3477_n2924) );
  INVX1_HVT U1323 ( .A(src_window[42]), .Y(DP_OP_424J2_126_3477_n2925) );
  INVX1_HVT U1324 ( .A(src_window[41]), .Y(DP_OP_424J2_126_3477_n2926) );
  INVX1_HVT U1325 ( .A(src_window[40]), .Y(DP_OP_424J2_126_3477_n2927) );
  INVX1_HVT U1326 ( .A(conv_weight_box[18]), .Y(DP_OP_424J2_126_3477_n2929) );
  INVX1_HVT U1327 ( .A(src_window[31]), .Y(DP_OP_424J2_126_3477_n2964) );
  INVX1_HVT U1328 ( .A(src_window[28]), .Y(DP_OP_424J2_126_3477_n2967) );
  INVX1_HVT U1329 ( .A(src_window[26]), .Y(DP_OP_424J2_126_3477_n2969) );
  INVX1_HVT U1330 ( .A(src_window[25]), .Y(DP_OP_424J2_126_3477_n2970) );
  INVX1_HVT U1331 ( .A(conv_weight_box[8]), .Y(DP_OP_424J2_126_3477_n2975) );
  INVX1_HVT U1332 ( .A(src_window[15]), .Y(DP_OP_424J2_126_3477_n3006) );
  INVX1_HVT U1333 ( .A(src_window[14]), .Y(DP_OP_424J2_126_3477_n3007) );
  INVX1_HVT U1334 ( .A(src_window[13]), .Y(DP_OP_424J2_126_3477_n3008) );
  INVX1_HVT U1335 ( .A(src_window[12]), .Y(DP_OP_424J2_126_3477_n3009) );
  INVX1_HVT U1336 ( .A(src_window[11]), .Y(DP_OP_424J2_126_3477_n3010) );
  INVX1_HVT U1337 ( .A(src_window[10]), .Y(DP_OP_424J2_126_3477_n3011) );
  INVX1_HVT U1338 ( .A(src_window[9]), .Y(DP_OP_424J2_126_3477_n3012) );
  INVX1_HVT U1339 ( .A(src_window[8]), .Y(DP_OP_424J2_126_3477_n3013) );
  INVX1_HVT U1340 ( .A(conv_weight_box[2]), .Y(DP_OP_424J2_126_3477_n3015) );
  INVX1_HVT U1341 ( .A(conv_weight_box[1]), .Y(DP_OP_424J2_126_3477_n3016) );
  INVX1_HVT U1342 ( .A(DP_OP_424J2_126_3477_n460), .Y(
        DP_OP_424J2_126_3477_n461) );
  INVX1_HVT U1343 ( .A(DP_OP_424J2_126_3477_n770), .Y(
        DP_OP_424J2_126_3477_n771) );
  OR2X1_HVT U1344 ( .A1(DP_OP_424J2_126_3477_n252), .A2(n443), .Y(n442) );
  OR2X1_HVT U1345 ( .A1(n378), .A2(n385), .Y(n443) );
  OR2X1_HVT U1346 ( .A1(DP_OP_424J2_126_3477_n258), .A2(
        DP_OP_424J2_126_3477_n257), .Y(n444) );
  OR2X1_HVT U1347 ( .A1(DP_OP_424J2_126_3477_n262), .A2(
        DP_OP_424J2_126_3477_n261), .Y(n445) );
  OR2X1_HVT U1348 ( .A1(DP_OP_424J2_126_3477_n264), .A2(
        DP_OP_424J2_126_3477_n263), .Y(n446) );
  OR2X1_HVT U1349 ( .A1(DP_OP_424J2_126_3477_n268), .A2(
        DP_OP_424J2_126_3477_n267), .Y(n447) );
  OR2X1_HVT U1350 ( .A1(DP_OP_424J2_126_3477_n971), .A2(
        DP_OP_424J2_126_3477_n969), .Y(n448) );
  OR2X1_HVT U1351 ( .A1(DP_OP_424J2_126_3477_n1353), .A2(
        DP_OP_424J2_126_3477_n1351), .Y(n449) );
  OR2X1_HVT U1352 ( .A1(DP_OP_424J2_126_3477_n1683), .A2(
        DP_OP_424J2_126_3477_n1681), .Y(n450) );
  OR2X1_HVT U1353 ( .A1(DP_OP_424J2_126_3477_n272), .A2(
        DP_OP_424J2_126_3477_n271), .Y(n451) );
  OR2X1_HVT U1354 ( .A1(DP_OP_424J2_126_3477_n276), .A2(
        DP_OP_424J2_126_3477_n275), .Y(n452) );
  INVX1_HVT U1355 ( .A(DP_OP_424J2_126_3477_n288), .Y(
        DP_OP_424J2_126_3477_n289) );
  INVX1_HVT U1356 ( .A(DP_OP_424J2_126_3477_n162), .Y(
        DP_OP_424J2_126_3477_n161) );
  INVX1_HVT U1357 ( .A(DP_OP_425J2_127_3477_n148), .Y(
        DP_OP_425J2_127_3477_n236) );
  INVX1_HVT U1358 ( .A(DP_OP_425J2_127_3477_n152), .Y(
        DP_OP_425J2_127_3477_n158) );
  INVX1_HVT U1359 ( .A(DP_OP_425J2_127_3477_n1678), .Y(
        DP_OP_425J2_127_3477_n1679) );
  INVX1_HVT U1360 ( .A(DP_OP_425J2_127_3477_n183), .Y(
        DP_OP_425J2_127_3477_n182) );
  INVX1_HVT U1361 ( .A(conv_weight_box[6]), .Y(DP_OP_425J2_127_3477_n1961) );
  INVX1_HVT U1362 ( .A(conv_weight_box[4]), .Y(DP_OP_425J2_127_3477_n1963) );
  INVX1_HVT U1363 ( .A(src_window[30]), .Y(DP_OP_425J2_127_3477_n1997) );
  INVX1_HVT U1364 ( .A(src_window[29]), .Y(DP_OP_425J2_127_3477_n1998) );
  INVX1_HVT U1365 ( .A(src_window[27]), .Y(DP_OP_425J2_127_3477_n2000) );
  INVX1_HVT U1366 ( .A(src_window[24]), .Y(DP_OP_425J2_127_3477_n2003) );
  INVX1_HVT U1367 ( .A(conv_weight_box[15]), .Y(DP_OP_425J2_127_3477_n2004) );
  INVX1_HVT U1368 ( .A(conv_weight_box[14]), .Y(DP_OP_425J2_127_3477_n2005) );
  INVX1_HVT U1369 ( .A(conv_weight_box[13]), .Y(DP_OP_425J2_127_3477_n2006) );
  INVX1_HVT U1370 ( .A(conv_weight_box[12]), .Y(DP_OP_425J2_127_3477_n2007) );
  INVX1_HVT U1371 ( .A(src_window[48]), .Y(DP_OP_425J2_127_3477_n2047) );
  INVX1_HVT U1372 ( .A(conv_weight_box[23]), .Y(DP_OP_425J2_127_3477_n2048) );
  INVX1_HVT U1373 ( .A(conv_weight_box[22]), .Y(DP_OP_425J2_127_3477_n2049) );
  INVX1_HVT U1374 ( .A(conv_weight_box[21]), .Y(DP_OP_425J2_127_3477_n2050) );
  INVX1_HVT U1375 ( .A(conv_weight_box[20]), .Y(DP_OP_425J2_127_3477_n2051) );
  INVX1_HVT U1376 ( .A(src_window[71]), .Y(DP_OP_425J2_127_3477_n2084) );
  INVX1_HVT U1377 ( .A(src_window[70]), .Y(DP_OP_425J2_127_3477_n2085) );
  INVX1_HVT U1378 ( .A(src_window[69]), .Y(DP_OP_425J2_127_3477_n2086) );
  INVX1_HVT U1379 ( .A(src_window[68]), .Y(DP_OP_425J2_127_3477_n2087) );
  INVX1_HVT U1380 ( .A(src_window[67]), .Y(DP_OP_425J2_127_3477_n2088) );
  INVX1_HVT U1381 ( .A(conv_weight_box[31]), .Y(DP_OP_425J2_127_3477_n2092) );
  INVX1_HVT U1382 ( .A(conv_weight_box[30]), .Y(DP_OP_425J2_127_3477_n2093) );
  INVX1_HVT U1383 ( .A(conv_weight_box[29]), .Y(DP_OP_425J2_127_3477_n2094) );
  INVX1_HVT U1384 ( .A(conv_weight_box[28]), .Y(DP_OP_425J2_127_3477_n2095) );
  INVX1_HVT U1385 ( .A(src_window[87]), .Y(DP_OP_425J2_127_3477_n2128) );
  INVX1_HVT U1386 ( .A(src_window[82]), .Y(DP_OP_425J2_127_3477_n2133) );
  INVX1_HVT U1387 ( .A(src_window[81]), .Y(DP_OP_425J2_127_3477_n2134) );
  INVX1_HVT U1388 ( .A(src_window[80]), .Y(DP_OP_425J2_127_3477_n2135) );
  INVX1_HVT U1389 ( .A(conv_weight_box[39]), .Y(DP_OP_425J2_127_3477_n2136) );
  INVX1_HVT U1390 ( .A(conv_weight_box[38]), .Y(DP_OP_425J2_127_3477_n2137) );
  INVX1_HVT U1391 ( .A(conv_weight_box[37]), .Y(DP_OP_425J2_127_3477_n2138) );
  INVX1_HVT U1392 ( .A(conv_weight_box[36]), .Y(DP_OP_425J2_127_3477_n2139) );
  INVX1_HVT U1393 ( .A(src_window[111]), .Y(DP_OP_425J2_127_3477_n2172) );
  INVX1_HVT U1394 ( .A(src_window[108]), .Y(DP_OP_425J2_127_3477_n2175) );
  INVX1_HVT U1395 ( .A(src_window[105]), .Y(DP_OP_425J2_127_3477_n2178) );
  INVX1_HVT U1396 ( .A(conv_weight_box[47]), .Y(DP_OP_425J2_127_3477_n2180) );
  INVX1_HVT U1397 ( .A(conv_weight_box[46]), .Y(DP_OP_425J2_127_3477_n2181) );
  INVX1_HVT U1398 ( .A(conv_weight_box[45]), .Y(DP_OP_425J2_127_3477_n2182) );
  INVX1_HVT U1399 ( .A(src_window[127]), .Y(DP_OP_425J2_127_3477_n2216) );
  INVX1_HVT U1400 ( .A(src_window[126]), .Y(DP_OP_425J2_127_3477_n2217) );
  INVX1_HVT U1401 ( .A(src_window[125]), .Y(DP_OP_425J2_127_3477_n2218) );
  INVX1_HVT U1402 ( .A(src_window[124]), .Y(DP_OP_425J2_127_3477_n2219) );
  INVX1_HVT U1403 ( .A(src_window[123]), .Y(DP_OP_425J2_127_3477_n2220) );
  INVX1_HVT U1404 ( .A(conv_weight_box[55]), .Y(DP_OP_425J2_127_3477_n2224) );
  INVX1_HVT U1405 ( .A(conv_weight_box[53]), .Y(DP_OP_425J2_127_3477_n2226) );
  INVX1_HVT U1406 ( .A(conv_weight_box[52]), .Y(DP_OP_425J2_127_3477_n2227) );
  INVX1_HVT U1407 ( .A(src_window[151]), .Y(DP_OP_425J2_127_3477_n2260) );
  INVX1_HVT U1408 ( .A(src_window[150]), .Y(DP_OP_425J2_127_3477_n2261) );
  INVX1_HVT U1409 ( .A(src_window[147]), .Y(DP_OP_425J2_127_3477_n2264) );
  INVX1_HVT U1410 ( .A(conv_weight_box[63]), .Y(DP_OP_425J2_127_3477_n2268) );
  INVX1_HVT U1411 ( .A(conv_weight_box[62]), .Y(DP_OP_425J2_127_3477_n2269) );
  INVX1_HVT U1412 ( .A(conv_weight_box[61]), .Y(DP_OP_425J2_127_3477_n2270) );
  INVX1_HVT U1413 ( .A(conv_weight_box[60]), .Y(DP_OP_425J2_127_3477_n2271) );
  INVX1_HVT U1414 ( .A(src_window[167]), .Y(DP_OP_425J2_127_3477_n2304) );
  INVX1_HVT U1415 ( .A(src_window[166]), .Y(DP_OP_425J2_127_3477_n2305) );
  INVX1_HVT U1416 ( .A(src_window[164]), .Y(DP_OP_425J2_127_3477_n2307) );
  INVX1_HVT U1417 ( .A(src_window[163]), .Y(DP_OP_425J2_127_3477_n2308) );
  INVX1_HVT U1418 ( .A(conv_weight_box[71]), .Y(DP_OP_425J2_127_3477_n2312) );
  INVX1_HVT U1419 ( .A(conv_weight_box[70]), .Y(DP_OP_425J2_127_3477_n2313) );
  INVX1_HVT U1420 ( .A(conv_weight_box[69]), .Y(DP_OP_425J2_127_3477_n2314) );
  INVX1_HVT U1421 ( .A(conv_weight_box[68]), .Y(DP_OP_425J2_127_3477_n2315) );
  INVX1_HVT U1422 ( .A(src_window[180]), .Y(DP_OP_425J2_127_3477_n2351) );
  INVX1_HVT U1423 ( .A(src_window[178]), .Y(DP_OP_425J2_127_3477_n2353) );
  INVX1_HVT U1424 ( .A(src_window[177]), .Y(DP_OP_425J2_127_3477_n2354) );
  INVX1_HVT U1425 ( .A(src_window[176]), .Y(DP_OP_425J2_127_3477_n2355) );
  INVX1_HVT U1426 ( .A(conv_weight_box[79]), .Y(DP_OP_425J2_127_3477_n2356) );
  INVX1_HVT U1427 ( .A(conv_weight_box[78]), .Y(DP_OP_425J2_127_3477_n2357) );
  INVX1_HVT U1428 ( .A(conv_weight_box[77]), .Y(DP_OP_425J2_127_3477_n2358) );
  INVX1_HVT U1429 ( .A(conv_weight_box[76]), .Y(DP_OP_425J2_127_3477_n2359) );
  INVX1_HVT U1430 ( .A(src_window[203]), .Y(DP_OP_425J2_127_3477_n2396) );
  INVX1_HVT U1431 ( .A(src_window[202]), .Y(DP_OP_425J2_127_3477_n2397) );
  INVX1_HVT U1432 ( .A(src_window[201]), .Y(DP_OP_425J2_127_3477_n2398) );
  INVX1_HVT U1433 ( .A(DP_OP_425J2_127_3477_n175), .Y(
        DP_OP_425J2_127_3477_n240) );
  INVX1_HVT U1434 ( .A(conv_weight_box[87]), .Y(DP_OP_425J2_127_3477_n2400) );
  INVX1_HVT U1435 ( .A(conv_weight_box[86]), .Y(DP_OP_425J2_127_3477_n2401) );
  INVX1_HVT U1436 ( .A(conv_weight_box[85]), .Y(DP_OP_425J2_127_3477_n2402) );
  INVX1_HVT U1437 ( .A(conv_weight_box[84]), .Y(DP_OP_425J2_127_3477_n2403) );
  INVX1_HVT U1438 ( .A(src_window[221]), .Y(DP_OP_425J2_127_3477_n2438) );
  INVX1_HVT U1439 ( .A(src_window[220]), .Y(DP_OP_425J2_127_3477_n2439) );
  INVX1_HVT U1440 ( .A(src_window[218]), .Y(DP_OP_425J2_127_3477_n2441) );
  INVX1_HVT U1441 ( .A(src_window[217]), .Y(DP_OP_425J2_127_3477_n2442) );
  INVX1_HVT U1442 ( .A(conv_weight_box[94]), .Y(DP_OP_425J2_127_3477_n2445) );
  INVX1_HVT U1443 ( .A(conv_weight_box[93]), .Y(DP_OP_425J2_127_3477_n2446) );
  INVX1_HVT U1444 ( .A(conv_weight_box[92]), .Y(DP_OP_425J2_127_3477_n2447) );
  INVX1_HVT U1445 ( .A(src_window[230]), .Y(DP_OP_425J2_127_3477_n2481) );
  INVX1_HVT U1446 ( .A(src_window[229]), .Y(DP_OP_425J2_127_3477_n2482) );
  INVX1_HVT U1447 ( .A(src_window[227]), .Y(DP_OP_425J2_127_3477_n2484) );
  INVX1_HVT U1448 ( .A(conv_weight_box[99]), .Y(DP_OP_425J2_127_3477_n2488) );
  INVX1_HVT U1449 ( .A(conv_weight_box[98]), .Y(DP_OP_425J2_127_3477_n2489) );
  INVX1_HVT U1450 ( .A(conv_weight_box[97]), .Y(DP_OP_425J2_127_3477_n2490) );
  INVX1_HVT U1451 ( .A(conv_weight_box[96]), .Y(DP_OP_425J2_127_3477_n2491) );
  INVX1_HVT U1452 ( .A(src_window[214]), .Y(DP_OP_425J2_127_3477_n2525) );
  INVX1_HVT U1453 ( .A(src_window[213]), .Y(DP_OP_425J2_127_3477_n2526) );
  INVX1_HVT U1454 ( .A(src_window[211]), .Y(DP_OP_425J2_127_3477_n2528) );
  INVX1_HVT U1455 ( .A(src_window[210]), .Y(DP_OP_425J2_127_3477_n2529) );
  INVX1_HVT U1456 ( .A(DP_OP_425J2_127_3477_n252), .Y(
        DP_OP_425J2_127_3477_n253) );
  INVX1_HVT U1457 ( .A(src_window[209]), .Y(DP_OP_425J2_127_3477_n2530) );
  INVX1_HVT U1458 ( .A(conv_weight_box[89]), .Y(DP_OP_425J2_127_3477_n2534) );
  INVX1_HVT U1459 ( .A(conv_weight_box[88]), .Y(DP_OP_425J2_127_3477_n2535) );
  INVX1_HVT U1460 ( .A(DP_OP_425J2_127_3477_n254), .Y(
        DP_OP_425J2_127_3477_n255) );
  INVX1_HVT U1461 ( .A(DP_OP_425J2_127_3477_n256), .Y(
        DP_OP_425J2_127_3477_n257) );
  INVX1_HVT U1462 ( .A(src_window[195]), .Y(DP_OP_425J2_127_3477_n2572) );
  INVX1_HVT U1463 ( .A(conv_weight_box[83]), .Y(DP_OP_425J2_127_3477_n2576) );
  INVX1_HVT U1464 ( .A(conv_weight_box[82]), .Y(DP_OP_425J2_127_3477_n2577) );
  INVX1_HVT U1465 ( .A(conv_weight_box[81]), .Y(DP_OP_425J2_127_3477_n2578) );
  INVX1_HVT U1466 ( .A(conv_weight_box[80]), .Y(DP_OP_425J2_127_3477_n2579) );
  INVX1_HVT U1467 ( .A(DP_OP_425J2_127_3477_n258), .Y(
        DP_OP_425J2_127_3477_n259) );
  INVX1_HVT U1468 ( .A(DP_OP_425J2_127_3477_n260), .Y(
        DP_OP_425J2_127_3477_n261) );
  INVX1_HVT U1469 ( .A(src_window[175]), .Y(DP_OP_425J2_127_3477_n2612) );
  INVX1_HVT U1470 ( .A(src_window[171]), .Y(DP_OP_425J2_127_3477_n2616) );
  INVX1_HVT U1471 ( .A(src_window[170]), .Y(DP_OP_425J2_127_3477_n2617) );
  INVX1_HVT U1472 ( .A(src_window[168]), .Y(DP_OP_425J2_127_3477_n2619) );
  INVX1_HVT U1473 ( .A(conv_weight_box[75]), .Y(DP_OP_425J2_127_3477_n2620) );
  INVX1_HVT U1474 ( .A(conv_weight_box[74]), .Y(DP_OP_425J2_127_3477_n2621) );
  INVX1_HVT U1475 ( .A(conv_weight_box[73]), .Y(DP_OP_425J2_127_3477_n2622) );
  INVX1_HVT U1476 ( .A(conv_weight_box[72]), .Y(DP_OP_425J2_127_3477_n2623) );
  INVX1_HVT U1477 ( .A(DP_OP_425J2_127_3477_n262), .Y(
        DP_OP_425J2_127_3477_n263) );
  INVX1_HVT U1478 ( .A(DP_OP_425J2_127_3477_n264), .Y(
        DP_OP_425J2_127_3477_n265) );
  INVX1_HVT U1479 ( .A(src_window[157]), .Y(DP_OP_425J2_127_3477_n2658) );
  INVX1_HVT U1480 ( .A(src_window[153]), .Y(DP_OP_425J2_127_3477_n2662) );
  INVX1_HVT U1481 ( .A(src_window[152]), .Y(DP_OP_425J2_127_3477_n2663) );
  INVX1_HVT U1482 ( .A(conv_weight_box[67]), .Y(DP_OP_425J2_127_3477_n2664) );
  INVX1_HVT U1483 ( .A(conv_weight_box[66]), .Y(DP_OP_425J2_127_3477_n2665) );
  INVX1_HVT U1484 ( .A(conv_weight_box[65]), .Y(DP_OP_425J2_127_3477_n2666) );
  INVX1_HVT U1485 ( .A(conv_weight_box[64]), .Y(DP_OP_425J2_127_3477_n2667) );
  INVX1_HVT U1486 ( .A(DP_OP_425J2_127_3477_n266), .Y(
        DP_OP_425J2_127_3477_n267) );
  INVX1_HVT U1487 ( .A(DP_OP_425J2_127_3477_n268), .Y(
        DP_OP_425J2_127_3477_n269) );
  INVX1_HVT U1488 ( .A(src_window[135]), .Y(DP_OP_425J2_127_3477_n2700) );
  INVX1_HVT U1489 ( .A(src_window[131]), .Y(DP_OP_425J2_127_3477_n2704) );
  INVX1_HVT U1490 ( .A(src_window[130]), .Y(DP_OP_425J2_127_3477_n2705) );
  INVX1_HVT U1491 ( .A(src_window[128]), .Y(DP_OP_425J2_127_3477_n2707) );
  INVX1_HVT U1492 ( .A(conv_weight_box[59]), .Y(DP_OP_425J2_127_3477_n2708) );
  INVX1_HVT U1493 ( .A(conv_weight_box[58]), .Y(DP_OP_425J2_127_3477_n2709) );
  INVX1_HVT U1494 ( .A(DP_OP_425J2_127_3477_n270), .Y(
        DP_OP_425J2_127_3477_n271) );
  INVX1_HVT U1495 ( .A(conv_weight_box[57]), .Y(DP_OP_425J2_127_3477_n2710) );
  INVX1_HVT U1496 ( .A(conv_weight_box[56]), .Y(DP_OP_425J2_127_3477_n2711) );
  INVX1_HVT U1497 ( .A(DP_OP_425J2_127_3477_n272), .Y(
        DP_OP_425J2_127_3477_n273) );
  INVX1_HVT U1498 ( .A(src_window[118]), .Y(DP_OP_425J2_127_3477_n2745) );
  INVX1_HVT U1499 ( .A(src_window[116]), .Y(DP_OP_425J2_127_3477_n2747) );
  INVX1_HVT U1500 ( .A(src_window[114]), .Y(DP_OP_425J2_127_3477_n2749) );
  INVX1_HVT U1501 ( .A(DP_OP_425J2_127_3477_n274), .Y(
        DP_OP_425J2_127_3477_n275) );
  INVX1_HVT U1502 ( .A(src_window[113]), .Y(DP_OP_425J2_127_3477_n2750) );
  INVX1_HVT U1503 ( .A(conv_weight_box[51]), .Y(DP_OP_425J2_127_3477_n2752) );
  INVX1_HVT U1504 ( .A(conv_weight_box[49]), .Y(DP_OP_425J2_127_3477_n2754) );
  INVX1_HVT U1505 ( .A(conv_weight_box[48]), .Y(DP_OP_425J2_127_3477_n2755) );
  INVX1_HVT U1506 ( .A(DP_OP_425J2_127_3477_n276), .Y(
        DP_OP_425J2_127_3477_n277) );
  INVX1_HVT U1507 ( .A(src_window[102]), .Y(DP_OP_425J2_127_3477_n2789) );
  INVX1_HVT U1508 ( .A(DP_OP_425J2_127_3477_n278), .Y(
        DP_OP_425J2_127_3477_n279) );
  INVX1_HVT U1509 ( .A(src_window[101]), .Y(DP_OP_425J2_127_3477_n2790) );
  INVX1_HVT U1510 ( .A(src_window[100]), .Y(DP_OP_425J2_127_3477_n2791) );
  INVX1_HVT U1511 ( .A(src_window[98]), .Y(DP_OP_425J2_127_3477_n2793) );
  INVX1_HVT U1512 ( .A(src_window[97]), .Y(DP_OP_425J2_127_3477_n2794) );
  INVX1_HVT U1513 ( .A(src_window[96]), .Y(DP_OP_425J2_127_3477_n2795) );
  INVX1_HVT U1514 ( .A(conv_weight_box[43]), .Y(DP_OP_425J2_127_3477_n2796) );
  INVX1_HVT U1515 ( .A(conv_weight_box[42]), .Y(DP_OP_425J2_127_3477_n2797) );
  INVX1_HVT U1516 ( .A(conv_weight_box[41]), .Y(DP_OP_425J2_127_3477_n2798) );
  INVX1_HVT U1517 ( .A(conv_weight_box[40]), .Y(DP_OP_425J2_127_3477_n2799) );
  INVX1_HVT U1518 ( .A(DP_OP_425J2_127_3477_n280), .Y(
        DP_OP_425J2_127_3477_n281) );
  INVX1_HVT U1519 ( .A(src_window[78]), .Y(DP_OP_425J2_127_3477_n2833) );
  INVX1_HVT U1520 ( .A(src_window[77]), .Y(DP_OP_425J2_127_3477_n2834) );
  INVX1_HVT U1521 ( .A(src_window[76]), .Y(DP_OP_425J2_127_3477_n2835) );
  INVX1_HVT U1522 ( .A(src_window[74]), .Y(DP_OP_425J2_127_3477_n2837) );
  INVX1_HVT U1523 ( .A(conv_weight_box[35]), .Y(DP_OP_425J2_127_3477_n2840) );
  INVX1_HVT U1524 ( .A(conv_weight_box[34]), .Y(DP_OP_425J2_127_3477_n2841) );
  INVX1_HVT U1525 ( .A(conv_weight_box[33]), .Y(DP_OP_425J2_127_3477_n2842) );
  INVX1_HVT U1526 ( .A(conv_weight_box[32]), .Y(DP_OP_425J2_127_3477_n2843) );
  INVX1_HVT U1527 ( .A(src_window[62]), .Y(DP_OP_425J2_127_3477_n2877) );
  INVX1_HVT U1528 ( .A(src_window[61]), .Y(DP_OP_425J2_127_3477_n2878) );
  INVX1_HVT U1529 ( .A(src_window[60]), .Y(DP_OP_425J2_127_3477_n2879) );
  INVX1_HVT U1530 ( .A(conv_weight_box[27]), .Y(DP_OP_425J2_127_3477_n2884) );
  INVX1_HVT U1531 ( .A(conv_weight_box[24]), .Y(DP_OP_425J2_127_3477_n2887) );
  INVX1_HVT U1532 ( .A(src_window[39]), .Y(DP_OP_425J2_127_3477_n2920) );
  INVX1_HVT U1533 ( .A(src_window[38]), .Y(DP_OP_425J2_127_3477_n2921) );
  INVX1_HVT U1534 ( .A(src_window[37]), .Y(DP_OP_425J2_127_3477_n2922) );
  INVX1_HVT U1535 ( .A(src_window[36]), .Y(DP_OP_425J2_127_3477_n2923) );
  INVX1_HVT U1536 ( .A(src_window[35]), .Y(DP_OP_425J2_127_3477_n2924) );
  INVX1_HVT U1537 ( .A(src_window[33]), .Y(DP_OP_425J2_127_3477_n2926) );
  INVX1_HVT U1538 ( .A(src_window[32]), .Y(DP_OP_425J2_127_3477_n2927) );
  INVX1_HVT U1539 ( .A(conv_weight_box[19]), .Y(DP_OP_425J2_127_3477_n2928) );
  INVX1_HVT U1540 ( .A(conv_weight_box[18]), .Y(DP_OP_425J2_127_3477_n2929) );
  INVX1_HVT U1541 ( .A(conv_weight_box[17]), .Y(DP_OP_425J2_127_3477_n2930) );
  INVX1_HVT U1542 ( .A(conv_weight_box[16]), .Y(DP_OP_425J2_127_3477_n2931) );
  INVX1_HVT U1543 ( .A(src_window[23]), .Y(DP_OP_425J2_127_3477_n2964) );
  INVX1_HVT U1544 ( .A(src_window[22]), .Y(DP_OP_425J2_127_3477_n2965) );
  INVX1_HVT U1545 ( .A(src_window[20]), .Y(DP_OP_425J2_127_3477_n2967) );
  INVX1_HVT U1546 ( .A(src_window[16]), .Y(DP_OP_425J2_127_3477_n2971) );
  INVX1_HVT U1547 ( .A(conv_weight_box[11]), .Y(DP_OP_425J2_127_3477_n2972) );
  INVX1_HVT U1548 ( .A(conv_weight_box[10]), .Y(DP_OP_425J2_127_3477_n2973) );
  INVX1_HVT U1549 ( .A(conv_weight_box[9]), .Y(DP_OP_425J2_127_3477_n2974) );
  INVX1_HVT U1550 ( .A(conv_weight_box[8]), .Y(DP_OP_425J2_127_3477_n2975) );
  INVX1_HVT U1551 ( .A(src_window[7]), .Y(DP_OP_425J2_127_3477_n3006) );
  INVX1_HVT U1552 ( .A(src_window[6]), .Y(DP_OP_425J2_127_3477_n3007) );
  INVX1_HVT U1553 ( .A(src_window[5]), .Y(DP_OP_425J2_127_3477_n3008) );
  INVX1_HVT U1554 ( .A(src_window[4]), .Y(DP_OP_425J2_127_3477_n3009) );
  INVX1_HVT U1555 ( .A(src_window[3]), .Y(DP_OP_425J2_127_3477_n3010) );
  INVX1_HVT U1556 ( .A(src_window[2]), .Y(DP_OP_425J2_127_3477_n3011) );
  INVX1_HVT U1557 ( .A(src_window[1]), .Y(DP_OP_425J2_127_3477_n3012) );
  INVX1_HVT U1558 ( .A(src_window[0]), .Y(DP_OP_425J2_127_3477_n3013) );
  INVX1_HVT U1559 ( .A(conv_weight_box[2]), .Y(DP_OP_425J2_127_3477_n3015) );
  INVX1_HVT U1560 ( .A(conv_weight_box[0]), .Y(DP_OP_425J2_127_3477_n3017) );
  INVX1_HVT U1561 ( .A(DP_OP_425J2_127_3477_n460), .Y(
        DP_OP_425J2_127_3477_n461) );
  INVX1_HVT U1562 ( .A(DP_OP_425J2_127_3477_n770), .Y(
        DP_OP_425J2_127_3477_n771) );
  OR2X1_HVT U1563 ( .A1(DP_OP_425J2_127_3477_n252), .A2(n463), .Y(n453) );
  OR2X1_HVT U1564 ( .A1(DP_OP_425J2_127_3477_n258), .A2(
        DP_OP_425J2_127_3477_n257), .Y(n454) );
  OR2X1_HVT U1565 ( .A1(DP_OP_425J2_127_3477_n262), .A2(
        DP_OP_425J2_127_3477_n261), .Y(n455) );
  OR2X1_HVT U1566 ( .A1(DP_OP_425J2_127_3477_n264), .A2(
        DP_OP_425J2_127_3477_n263), .Y(n456) );
  OR2X1_HVT U1567 ( .A1(DP_OP_425J2_127_3477_n268), .A2(
        DP_OP_425J2_127_3477_n267), .Y(n457) );
  OR2X1_HVT U1568 ( .A1(DP_OP_425J2_127_3477_n971), .A2(
        DP_OP_425J2_127_3477_n969), .Y(n458) );
  OR2X1_HVT U1569 ( .A1(DP_OP_425J2_127_3477_n1353), .A2(
        DP_OP_425J2_127_3477_n1351), .Y(n459) );
  OR2X1_HVT U1570 ( .A1(DP_OP_425J2_127_3477_n1683), .A2(
        DP_OP_425J2_127_3477_n1681), .Y(n460) );
  OR2X1_HVT U1571 ( .A1(DP_OP_425J2_127_3477_n272), .A2(
        DP_OP_425J2_127_3477_n271), .Y(n461) );
  OR2X1_HVT U1572 ( .A1(DP_OP_425J2_127_3477_n276), .A2(
        DP_OP_425J2_127_3477_n275), .Y(n462) );
  OR2X1_HVT U1573 ( .A1(n530), .A2(n388), .Y(n463) );
  AOI21X2_HVT U1574 ( .A1(DP_OP_425J2_127_3477_n162), .A2(
        DP_OP_425J2_127_3477_n135), .A3(DP_OP_425J2_127_3477_n136), .Y(
        DP_OP_425J2_127_3477_n3) );
  INVX1_HVT U1575 ( .A(DP_OP_425J2_127_3477_n288), .Y(
        DP_OP_425J2_127_3477_n289) );
  INVX1_HVT U1576 ( .A(DP_OP_425J2_127_3477_n162), .Y(
        DP_OP_425J2_127_3477_n161) );
  INVX1_HVT U1577 ( .A(conv_weight_box[7]), .Y(DP_OP_425J2_127_3477_n1960) );
  INVX1_HVT U1578 ( .A(conv_weight_box[3]), .Y(DP_OP_425J2_127_3477_n3014) );
  MUX21X1_HVT U1579 ( .A1(tmp_big2[11]), .A2(tmp_big1[11]), .S0(n471), .Y(
        data_out[11]) );
  MUX21X1_HVT U1580 ( .A1(n466), .A2(n545), .S0(n412), .Y(n465) );
  OAI22X1_HVT U1581 ( .A1(n469), .A2(n468), .A3(n469), .A4(n467), .Y(n696) );
  OAI22X1_HVT U1582 ( .A1(n748), .A2(tmp_big2[17]), .A3(n692), .A4(
        tmp_big2[16]), .Y(n468) );
  OAI22X1_HVT U1583 ( .A1(tmp_big2[19]), .A2(n750), .A3(tmp_big2[18]), .A4(
        n691), .Y(n469) );
  MUX21X1_HVT U1584 ( .A1(conv2_sram_rdata_weight[6]), .A2(
        conv1_sram_rdata_weight[6]), .S0(n393), .Y(conv_weight_box[6]) );
  MUX21X1_HVT U1585 ( .A1(conv2_sram_rdata_weight[50]), .A2(
        conv1_sram_rdata_weight[50]), .S0(n395), .Y(conv_weight_box[50]) );
  MUX21X1_HVT U1586 ( .A1(conv2_sram_rdata_weight[58]), .A2(
        conv1_sram_rdata_weight[58]), .S0(n392), .Y(conv_weight_box[58]) );
  MUX21X1_HVT U1587 ( .A1(conv2_sram_rdata_weight[46]), .A2(
        conv1_sram_rdata_weight[46]), .S0(n400), .Y(conv_weight_box[46]) );
  MUX21X1_HVT U1588 ( .A1(conv2_sram_rdata_weight[82]), .A2(
        conv1_sram_rdata_weight[82]), .S0(n399), .Y(conv_weight_box[82]) );
  MUX21X1_HVT U1589 ( .A1(conv2_sram_rdata_weight[38]), .A2(
        conv1_sram_rdata_weight[38]), .S0(n393), .Y(conv_weight_box[38]) );
  MUX21X1_HVT U1590 ( .A1(conv2_sram_rdata_weight[30]), .A2(
        conv1_sram_rdata_weight[30]), .S0(n401), .Y(conv_weight_box[30]) );
  MUX21X1_HVT U1591 ( .A1(conv2_sram_rdata_weight[2]), .A2(
        conv1_sram_rdata_weight[2]), .S0(n400), .Y(conv_weight_box[2]) );
  MUX21X1_HVT U1592 ( .A1(conv2_sram_rdata_weight[18]), .A2(
        conv1_sram_rdata_weight[18]), .S0(n393), .Y(conv_weight_box[18]) );
  MUX21X1_HVT U1593 ( .A1(conv2_sram_rdata_weight[90]), .A2(
        conv1_sram_rdata_weight[90]), .S0(n395), .Y(conv_weight_box[90]) );
  MUX21X1_HVT U1594 ( .A1(conv2_sram_rdata_weight[70]), .A2(
        conv1_sram_rdata_weight[70]), .S0(n384), .Y(conv_weight_box[70]) );
  MUX21X1_HVT U1595 ( .A1(conv2_sram_rdata_weight[54]), .A2(
        conv1_sram_rdata_weight[54]), .S0(n397), .Y(conv_weight_box[54]) );
  MUX21X1_HVT U1596 ( .A1(conv2_sram_rdata_weight[66]), .A2(
        conv1_sram_rdata_weight[66]), .S0(n402), .Y(conv_weight_box[66]) );
  MUX21X1_HVT U1597 ( .A1(conv2_sram_rdata_weight[34]), .A2(
        conv1_sram_rdata_weight[34]), .S0(n399), .Y(conv_weight_box[34]) );
  MUX21X1_HVT U1598 ( .A1(conv2_sram_rdata_weight[14]), .A2(
        conv1_sram_rdata_weight[14]), .S0(n392), .Y(conv_weight_box[14]) );
  MUX21X1_HVT U1599 ( .A1(conv2_sram_rdata_weight[22]), .A2(
        conv1_sram_rdata_weight[22]), .S0(n400), .Y(conv_weight_box[22]) );
  MUX21X1_HVT U1600 ( .A1(conv2_sram_rdata_weight[74]), .A2(
        conv1_sram_rdata_weight[74]), .S0(n404), .Y(conv_weight_box[74]) );
  MUX21X1_HVT U1601 ( .A1(conv2_sram_rdata_weight[10]), .A2(
        conv1_sram_rdata_weight[10]), .S0(n400), .Y(conv_weight_box[10]) );
  MUX21X1_HVT U1602 ( .A1(conv2_sram_rdata_weight[98]), .A2(
        conv1_sram_rdata_weight[98]), .S0(n398), .Y(conv_weight_box[98]) );
  MUX21X1_HVT U1603 ( .A1(conv2_sram_rdata_weight[86]), .A2(
        conv1_sram_rdata_weight[86]), .S0(n392), .Y(conv_weight_box[86]) );
  MUX21X1_HVT U1604 ( .A1(conv2_sram_rdata_weight[81]), .A2(
        conv1_sram_rdata_weight[81]), .S0(n404), .Y(conv_weight_box[81]) );
  MUX21X1_HVT U1605 ( .A1(conv2_sram_rdata_weight[73]), .A2(
        conv1_sram_rdata_weight[73]), .S0(n403), .Y(conv_weight_box[73]) );
  MUX21X1_HVT U1606 ( .A1(conv2_sram_rdata_weight[85]), .A2(
        conv1_sram_rdata_weight[85]), .S0(n402), .Y(conv_weight_box[85]) );
  MUX21X1_HVT U1607 ( .A1(conv2_sram_rdata_weight[61]), .A2(
        conv1_sram_rdata_weight[61]), .S0(n392), .Y(conv_weight_box[61]) );
  MUX21X1_HVT U1608 ( .A1(conv2_sram_rdata_weight[93]), .A2(
        conv1_sram_rdata_weight[93]), .S0(n397), .Y(conv_weight_box[93]) );
  MUX21X1_HVT U1609 ( .A1(conv2_sram_rdata_weight[21]), .A2(
        conv1_sram_rdata_weight[21]), .S0(n402), .Y(conv_weight_box[21]) );
  MUX21X1_HVT U1610 ( .A1(conv2_sram_rdata_weight[33]), .A2(
        conv1_sram_rdata_weight[33]), .S0(n395), .Y(conv_weight_box[33]) );
  MUX21X1_HVT U1611 ( .A1(conv2_sram_rdata_weight[97]), .A2(
        conv1_sram_rdata_weight[97]), .S0(n401), .Y(conv_weight_box[97]) );
  MUX21X1_HVT U1612 ( .A1(conv2_sram_rdata_weight[89]), .A2(
        conv1_sram_rdata_weight[89]), .S0(n399), .Y(conv_weight_box[89]) );
  MUX21X1_HVT U1613 ( .A1(conv2_sram_rdata_weight[37]), .A2(
        conv1_sram_rdata_weight[37]), .S0(n384), .Y(conv_weight_box[37]) );
  MUX21X1_HVT U1614 ( .A1(conv2_sram_rdata_weight[41]), .A2(
        conv1_sram_rdata_weight[41]), .S0(n400), .Y(conv_weight_box[41]) );
  MUX21X1_HVT U1615 ( .A1(conv2_sram_rdata_weight[77]), .A2(
        conv1_sram_rdata_weight[77]), .S0(n402), .Y(conv_weight_box[77]) );
  MUX21X1_HVT U1616 ( .A1(conv2_sram_rdata_weight[49]), .A2(
        conv1_sram_rdata_weight[49]), .S0(n403), .Y(conv_weight_box[49]) );
  MUX21X1_HVT U1617 ( .A1(conv2_sram_rdata_weight[13]), .A2(
        conv1_sram_rdata_weight[13]), .S0(n395), .Y(conv_weight_box[13]) );
  MUX21X1_HVT U1618 ( .A1(conv2_sram_rdata_weight[69]), .A2(
        conv1_sram_rdata_weight[69]), .S0(n403), .Y(conv_weight_box[69]) );
  MUX21X1_HVT U1619 ( .A1(conv2_sram_rdata_weight[57]), .A2(
        conv1_sram_rdata_weight[57]), .S0(n404), .Y(conv_weight_box[57]) );
  MUX21X1_HVT U1620 ( .A1(conv2_sram_rdata_weight[25]), .A2(
        conv1_sram_rdata_weight[25]), .S0(n397), .Y(conv_weight_box[25]) );
  MUX21X1_HVT U1621 ( .A1(conv2_sram_rdata_weight[53]), .A2(
        conv1_sram_rdata_weight[53]), .S0(n403), .Y(conv_weight_box[53]) );
  MUX21X1_HVT U1622 ( .A1(conv2_sram_rdata_weight[1]), .A2(
        conv1_sram_rdata_weight[1]), .S0(n398), .Y(conv_weight_box[1]) );
  MUX21X1_HVT U1623 ( .A1(conv2_sram_rdata_weight[65]), .A2(
        conv1_sram_rdata_weight[65]), .S0(n401), .Y(conv_weight_box[65]) );
  MUX21X1_HVT U1624 ( .A1(tmp_big2[30]), .A2(tmp_big1[30]), .S0(n410), .Y(
        data_out[30]) );
  MUX21X1_HVT U1625 ( .A1(conv2_sram_rdata_weight[5]), .A2(
        conv1_sram_rdata_weight[5]), .S0(n398), .Y(conv_weight_box[5]) );
  MUX21X1_HVT U1626 ( .A1(conv2_sram_rdata_weight[80]), .A2(
        conv1_sram_rdata_weight[80]), .S0(n403), .Y(conv_weight_box[80]) );
  MUX21X1_HVT U1627 ( .A1(conv2_sram_rdata_weight[72]), .A2(
        conv1_sram_rdata_weight[72]), .S0(n393), .Y(conv_weight_box[72]) );
  MUX21X1_HVT U1628 ( .A1(conv2_sram_rdata_weight[0]), .A2(
        conv1_sram_rdata_weight[0]), .S0(n395), .Y(conv_weight_box[0]) );
  MUX21X1_HVT U1629 ( .A1(conv2_sram_rdata_weight[92]), .A2(
        conv1_sram_rdata_weight[92]), .S0(n397), .Y(conv_weight_box[92]) );
  MUX21X1_HVT U1630 ( .A1(conv2_sram_rdata_weight[56]), .A2(
        conv1_sram_rdata_weight[56]), .S0(n393), .Y(conv_weight_box[56]) );
  MUX21X1_HVT U1631 ( .A1(conv2_sram_rdata_weight[4]), .A2(
        conv1_sram_rdata_weight[4]), .S0(n403), .Y(conv_weight_box[4]) );
  MUX21X1_HVT U1632 ( .A1(conv2_sram_rdata_weight[40]), .A2(
        conv1_sram_rdata_weight[40]), .S0(n404), .Y(conv_weight_box[40]) );
  MUX21X1_HVT U1633 ( .A1(conv2_sram_rdata_weight[36]), .A2(
        conv1_sram_rdata_weight[36]), .S0(n399), .Y(conv_weight_box[36]) );
  MUX21X1_HVT U1634 ( .A1(conv2_sram_rdata_weight[29]), .A2(
        conv1_sram_rdata_weight[29]), .S0(n403), .Y(conv_weight_box[29]) );
  MUX21X1_HVT U1635 ( .A1(conv2_sram_rdata_weight[9]), .A2(
        conv1_sram_rdata_weight[9]), .S0(n400), .Y(conv_weight_box[9]) );
  MUX21X1_HVT U1636 ( .A1(conv2_sram_rdata_weight[8]), .A2(
        conv1_sram_rdata_weight[8]), .S0(n398), .Y(conv_weight_box[8]) );
  MUX21X1_HVT U1637 ( .A1(conv2_sram_rdata_weight[76]), .A2(
        conv1_sram_rdata_weight[76]), .S0(n384), .Y(conv_weight_box[76]) );
  MUX21X1_HVT U1638 ( .A1(conv2_sram_rdata_weight[17]), .A2(
        conv1_sram_rdata_weight[17]), .S0(n400), .Y(conv_weight_box[17]) );
  MUX21X1_HVT U1639 ( .A1(conv2_sram_rdata_weight[68]), .A2(
        conv1_sram_rdata_weight[68]), .S0(n392), .Y(conv_weight_box[68]) );
  MUX21X1_HVT U1640 ( .A1(conv2_sram_rdata_weight[60]), .A2(
        conv1_sram_rdata_weight[60]), .S0(n397), .Y(conv_weight_box[60]) );
  MUX21X1_HVT U1641 ( .A1(conv2_sram_rdata_weight[48]), .A2(
        conv1_sram_rdata_weight[48]), .S0(n401), .Y(conv_weight_box[48]) );
  MUX21X1_HVT U1642 ( .A1(conv2_sram_rdata_weight[84]), .A2(
        conv1_sram_rdata_weight[84]), .S0(n392), .Y(conv_weight_box[84]) );
  MUX21X1_HVT U1643 ( .A1(conv2_sram_rdata_weight[45]), .A2(
        conv1_sram_rdata_weight[45]), .S0(n402), .Y(conv_weight_box[45]) );
  MUX21X1_HVT U1644 ( .A1(conv2_sram_rdata_weight[88]), .A2(
        conv1_sram_rdata_weight[88]), .S0(n384), .Y(conv_weight_box[88]) );
  MUX21X1_HVT U1645 ( .A1(conv2_sram_rdata_weight[32]), .A2(
        conv1_sram_rdata_weight[32]), .S0(n384), .Y(conv_weight_box[32]) );
  MUX21X1_HVT U1646 ( .A1(conv2_sram_rdata_weight[20]), .A2(
        conv1_sram_rdata_weight[20]), .S0(n401), .Y(conv_weight_box[20]) );
  MUX21X1_HVT U1647 ( .A1(conv2_sram_rdata_weight[28]), .A2(
        conv1_sram_rdata_weight[28]), .S0(n404), .Y(conv_weight_box[28]) );
  MUX21X1_HVT U1648 ( .A1(conv2_sram_rdata_weight[52]), .A2(
        conv1_sram_rdata_weight[52]), .S0(n397), .Y(conv_weight_box[52]) );
  MUX21X1_HVT U1649 ( .A1(conv2_sram_rdata_weight[16]), .A2(
        conv1_sram_rdata_weight[16]), .S0(n402), .Y(conv_weight_box[16]) );
  MUX21X1_HVT U1650 ( .A1(conv2_sram_rdata_weight[96]), .A2(
        conv1_sram_rdata_weight[96]), .S0(n404), .Y(conv_weight_box[96]) );
  MUX21X1_HVT U1651 ( .A1(conv2_sram_rdata_weight[12]), .A2(
        conv1_sram_rdata_weight[12]), .S0(n400), .Y(conv_weight_box[12]) );
  MUX21X1_HVT U1652 ( .A1(conv2_sram_rdata_weight[24]), .A2(
        conv1_sram_rdata_weight[24]), .S0(n402), .Y(conv_weight_box[24]) );
  MUX21X1_HVT U1653 ( .A1(conv2_sram_rdata_weight[64]), .A2(
        conv1_sram_rdata_weight[64]), .S0(n393), .Y(conv_weight_box[64]) );
  MUX21X1_HVT U1654 ( .A1(conv2_sram_rdata_weight[44]), .A2(
        conv1_sram_rdata_weight[44]), .S0(n404), .Y(conv_weight_box[44]) );
  MUX21X1_HVT U1655 ( .A1(tmp_big2[31]), .A2(tmp_big1[31]), .S0(n411), .Y(
        data_out[31]) );
  OAI21X1_HVT U1656 ( .A1(tmp_big1[16]), .A2(n738), .A3(n729), .Y(n730) );
  MUX21X1_HVT U1657 ( .A1(conv2_sum_b[31]), .A2(conv2_sum_a[31]), .S0(n413), 
        .Y(tmp_big1[31]) );
  MUX21X1_HVT U1658 ( .A1(tmp_big2[7]), .A2(tmp_big1[7]), .S0(n409), .Y(
        data_out[7]) );
  MUX21X1_HVT U1659 ( .A1(tmp_big2[8]), .A2(tmp_big1[8]), .S0(n471), .Y(
        data_out[8]) );
  MUX21X1_HVT U1660 ( .A1(tmp_big2[9]), .A2(tmp_big1[9]), .S0(n471), .Y(
        data_out[9]) );
  MUX21X1_HVT U1661 ( .A1(tmp_big2[12]), .A2(tmp_big1[12]), .S0(n409), .Y(
        data_out[12]) );
  MUX21X1_HVT U1662 ( .A1(tmp_big2[13]), .A2(tmp_big1[13]), .S0(n471), .Y(
        data_out[13]) );
  MUX21X1_HVT U1663 ( .A1(tmp_big2[29]), .A2(tmp_big1[29]), .S0(n411), .Y(
        data_out[29]) );
  MUX21X1_HVT U1664 ( .A1(tmp_big2[23]), .A2(tmp_big1[23]), .S0(n410), .Y(
        data_out[23]) );
  MUX21X1_HVT U1665 ( .A1(tmp_big2[22]), .A2(tmp_big1[22]), .S0(n409), .Y(
        data_out[22]) );
  MUX21X1_HVT U1666 ( .A1(conv2_sum_d[31]), .A2(conv2_sum_c[31]), .S0(n417), 
        .Y(tmp_big2[31]) );
  MUX21X1_HVT U1667 ( .A1(conv2_sum_b[30]), .A2(conv2_sum_a[30]), .S0(n413), 
        .Y(tmp_big1[30]) );
  MUX21X1_HVT U1668 ( .A1(conv2_sum_d[30]), .A2(conv2_sum_c[30]), .S0(n419), 
        .Y(tmp_big2[30]) );
  MUX21X1_HVT U1669 ( .A1(conv2_sum_b[7]), .A2(conv2_sum_a[7]), .S0(n414), .Y(
        tmp_big1[7]) );
  MUX21X1_HVT U1670 ( .A1(conv2_sum_d[7]), .A2(conv2_sum_c[7]), .S0(n419), .Y(
        tmp_big2[7]) );
  MUX21X1_HVT U1671 ( .A1(conv2_sum_b[6]), .A2(conv2_sum_a[6]), .S0(n415), .Y(
        tmp_big1[6]) );
  MUX21X1_HVT U1672 ( .A1(conv2_sum_d[6]), .A2(conv2_sum_c[6]), .S0(n418), .Y(
        tmp_big2[6]) );
  MUX21X1_HVT U1673 ( .A1(conv2_sum_b[4]), .A2(conv2_sum_a[4]), .S0(n413), .Y(
        tmp_big1[4]) );
  MUX21X1_HVT U1674 ( .A1(conv2_sum_d[4]), .A2(conv2_sum_c[4]), .S0(n417), .Y(
        tmp_big2[4]) );
  MUX21X1_HVT U1675 ( .A1(conv2_sum_b[5]), .A2(conv2_sum_a[5]), .S0(n413), .Y(
        tmp_big1[5]) );
  MUX21X1_HVT U1676 ( .A1(conv2_sum_d[5]), .A2(conv2_sum_c[5]), .S0(n418), .Y(
        tmp_big2[5]) );
  MUX21X1_HVT U1677 ( .A1(conv2_sum_b[1]), .A2(conv2_sum_a[1]), .S0(n412), .Y(
        tmp_big1[1]) );
  MUX21X1_HVT U1678 ( .A1(n543), .A2(n544), .S0(n416), .Y(n542) );
  MUX21X1_HVT U1679 ( .A1(conv2_sum_d[0]), .A2(conv2_sum_c[0]), .S0(n416), .Y(
        tmp_big2[0]) );
  MUX21X1_HVT U1680 ( .A1(conv2_sum_b[0]), .A2(conv2_sum_a[0]), .S0(n415), .Y(
        tmp_big1[0]) );
  MUX21X1_HVT U1681 ( .A1(conv2_sum_b[2]), .A2(conv2_sum_a[2]), .S0(n412), .Y(
        tmp_big1[2]) );
  MUX21X1_HVT U1682 ( .A1(conv2_sum_d[2]), .A2(conv2_sum_c[2]), .S0(n419), .Y(
        tmp_big2[2]) );
  MUX21X1_HVT U1683 ( .A1(conv2_sum_d[3]), .A2(conv2_sum_c[3]), .S0(n416), .Y(
        tmp_big2[3]) );
  MUX21X1_HVT U1684 ( .A1(conv2_sum_d[8]), .A2(conv2_sum_c[8]), .S0(n417), .Y(
        tmp_big2[8]) );
  NAND2X4_HVT U1685 ( .A1(n533), .A2(n737), .Y(n471) );
  INVX1_HVT U1686 ( .A(n542), .Y(tmp_big2[1]) );
  INVX1_HVT U1687 ( .A(n547), .Y(tmp_big1[9]) );
  INVX1_HVT U1688 ( .A(tmp_big1[25]), .Y(n754) );
  INVX1_HVT U1689 ( .A(tmp_big1[29]), .Y(n757) );
  INVX1_HVT U1690 ( .A(tmp_big2[31]), .Y(n739) );
  INVX1_HVT U1691 ( .A(tmp_big1[27]), .Y(n756) );
  INVX1_HVT U1692 ( .A(tmp_big1[26]), .Y(n755) );
  INVX1_HVT U1693 ( .A(tmp_big1[7]), .Y(n763) );
  INVX1_HVT U1694 ( .A(tmp_big1[5]), .Y(n761) );
  AO22X1_HVT U1695 ( .A1(tmp_big2[2]), .A2(n758), .A3(tmp_big2[3]), .A4(n465), 
        .Y(n721) );
  INVX1_HVT U1696 ( .A(tmp_big2[16]), .Y(n738) );
  INVX1_HVT U1697 ( .A(tmp_big1[21]), .Y(n751) );
  INVX1_HVT U1698 ( .A(tmp_big1[23]), .Y(n753) );
  INVX1_HVT U1699 ( .A(tmp_big1[18]), .Y(n749) );
  INVX1_HVT U1700 ( .A(tmp_big1[13]), .Y(n744) );
  INVX1_HVT U1701 ( .A(tmp_big1[15]), .Y(n746) );
  AO22X1_HVT U1702 ( .A1(conv2_sum_d[2]), .A2(n481), .A3(conv2_sum_d[3]), .A4(
        n490), .Y(n656) );
  NOR3X0_HVT U1703 ( .A1(n714), .A2(n713), .A3(n712), .Y(n492) );
  NAND2X0_HVT U1704 ( .A1(n532), .A2(n531), .Y(n535) );
  NAND3X0_HVT U1705 ( .A1(n470), .A2(n536), .A3(n492), .Y(n531) );
  OA21X1_HVT U1706 ( .A1(n734), .A2(n733), .A3(n735), .Y(n532) );
  NAND2X0_HVT U1707 ( .A1(n535), .A2(n534), .Y(n533) );
  OR2X1_HVT U1708 ( .A1(n538), .A2(conv2_sum_c[3]), .Y(n650) );
  NAND2X0_HVT U1709 ( .A1(n668), .A2(n667), .Y(n540) );
  NAND3X0_HVT U1710 ( .A1(n541), .A2(n540), .A3(n491), .Y(n669) );
  OR2X1_HVT U1711 ( .A1(n548), .A2(conv2_sum_a[9]), .Y(n579) );
  MUX21X1_HVT U1712 ( .A1(n548), .A2(n549), .S0(n412), .Y(n547) );
  AO22X1_HVT U1713 ( .A1(conv2_sum_b[30]), .A2(n527), .A3(conv2_sum_a[31]), 
        .A4(n529), .Y(n557) );
  NAND2X0_HVT U1714 ( .A1(conv2_sum_b[29]), .A2(n524), .Y(n551) );
  NAND2X0_HVT U1715 ( .A1(conv2_sum_a[28]), .A2(n551), .Y(n550) );
  OA22X1_HVT U1716 ( .A1(n524), .A2(conv2_sum_b[29]), .A3(n550), .A4(
        conv2_sum_b[28]), .Y(n556) );
  NAND2X0_HVT U1717 ( .A1(conv2_sum_b[25]), .A2(n511), .Y(n611) );
  AO22X1_HVT U1718 ( .A1(conv2_sum_b[26]), .A2(n519), .A3(conv2_sum_b[27]), 
        .A4(n523), .Y(n559) );
  NAND2X0_HVT U1719 ( .A1(conv2_sum_a[31]), .A2(n529), .Y(n552) );
  NAND2X0_HVT U1720 ( .A1(conv2_sum_a[30]), .A2(n552), .Y(n553) );
  OA22X1_HVT U1721 ( .A1(n529), .A2(conv2_sum_a[31]), .A3(n553), .A4(
        conv2_sum_b[30]), .Y(n554) );
  NAND2X0_HVT U1722 ( .A1(conv2_sum_b[24]), .A2(n499), .Y(n612) );
  AO22X1_HVT U1723 ( .A1(conv2_sum_b[22]), .A2(n498), .A3(conv2_sum_b[23]), 
        .A4(n510), .Y(n567) );
  NAND2X0_HVT U1724 ( .A1(conv2_sum_b[21]), .A2(n509), .Y(n561) );
  NAND2X0_HVT U1725 ( .A1(conv2_sum_a[20]), .A2(n561), .Y(n560) );
  OA22X1_HVT U1726 ( .A1(n509), .A2(conv2_sum_b[21]), .A3(n560), .A4(
        conv2_sum_b[20]), .Y(n566) );
  NAND2X0_HVT U1727 ( .A1(conv2_sum_b[17]), .A2(n507), .Y(n599) );
  AO22X1_HVT U1728 ( .A1(conv2_sum_b[18]), .A2(n482), .A3(conv2_sum_b[19]), 
        .A4(n508), .Y(n602) );
  NAND2X0_HVT U1729 ( .A1(conv2_sum_b[23]), .A2(n510), .Y(n562) );
  NAND2X0_HVT U1730 ( .A1(conv2_sum_a[22]), .A2(n562), .Y(n563) );
  OA22X1_HVT U1731 ( .A1(n510), .A2(conv2_sum_b[23]), .A3(n563), .A4(
        conv2_sum_b[22]), .Y(n564) );
  AO22X1_HVT U1732 ( .A1(conv2_sum_b[14]), .A2(n496), .A3(conv2_sum_b[15]), 
        .A4(n506), .Y(n578) );
  NAND2X0_HVT U1733 ( .A1(conv2_sum_b[13]), .A2(n505), .Y(n569) );
  NAND2X0_HVT U1734 ( .A1(conv2_sum_a[12]), .A2(n569), .Y(n568) );
  OA22X1_HVT U1735 ( .A1(n505), .A2(conv2_sum_b[13]), .A3(n568), .A4(
        conv2_sum_b[12]), .Y(n577) );
  NAND2X0_HVT U1736 ( .A1(conv2_sum_b[11]), .A2(n539), .Y(n570) );
  NAND2X0_HVT U1737 ( .A1(conv2_sum_a[10]), .A2(n570), .Y(n571) );
  NAND2X0_HVT U1738 ( .A1(conv2_sum_a[8]), .A2(n579), .Y(n572) );
  AO22X1_HVT U1739 ( .A1(conv2_sum_b[10]), .A2(n483), .A3(conv2_sum_b[11]), 
        .A4(n539), .Y(n582) );
  NAND2X0_HVT U1740 ( .A1(conv2_sum_b[15]), .A2(n506), .Y(n573) );
  NAND2X0_HVT U1741 ( .A1(conv2_sum_a[14]), .A2(n573), .Y(n574) );
  OA22X1_HVT U1742 ( .A1(n506), .A2(conv2_sum_b[15]), .A3(n574), .A4(
        conv2_sum_b[14]), .Y(n575) );
  OAI21X1_HVT U1743 ( .A1(conv2_sum_a[8]), .A2(n477), .A3(n579), .Y(n580) );
  OR3X1_HVT U1744 ( .A1(n582), .A2(n581), .A3(n580), .Y(n605) );
  NAND2X0_HVT U1745 ( .A1(conv2_sum_b[3]), .A2(n545), .Y(n583) );
  NAND2X0_HVT U1746 ( .A1(n583), .A2(conv2_sum_a[2]), .Y(n584) );
  OA22X1_HVT U1747 ( .A1(conv2_sum_b[3]), .A2(n545), .A3(conv2_sum_b[2]), .A4(
        n584), .Y(n590) );
  AO22X1_HVT U1748 ( .A1(conv2_sum_b[2]), .A2(n488), .A3(conv2_sum_b[3]), .A4(
        n545), .Y(n589) );
  NAND2X0_HVT U1749 ( .A1(conv2_sum_a[1]), .A2(n546), .Y(n585) );
  NAND2X0_HVT U1750 ( .A1(n585), .A2(conv2_sum_b[0]), .Y(n586) );
  OAI22X1_HVT U1751 ( .A1(conv2_sum_a[0]), .A2(n586), .A3(n546), .A4(
        conv2_sum_a[1]), .Y(n588) );
  AO22X1_HVT U1752 ( .A1(conv2_sum_b[5]), .A2(n472), .A3(conv2_sum_b[4]), .A4(
        n479), .Y(n587) );
  AO221X1_HVT U1753 ( .A1(n590), .A2(n589), .A3(n588), .A4(n590), .A5(n587), 
        .Y(n598) );
  AO22X1_HVT U1754 ( .A1(conv2_sum_b[6]), .A2(n484), .A3(conv2_sum_b[7]), .A4(
        n473), .Y(n597) );
  NAND2X0_HVT U1755 ( .A1(conv2_sum_b[5]), .A2(n472), .Y(n591) );
  NAND2X0_HVT U1756 ( .A1(conv2_sum_a[4]), .A2(n591), .Y(n592) );
  OA22X1_HVT U1757 ( .A1(n592), .A2(conv2_sum_b[4]), .A3(n472), .A4(
        conv2_sum_b[5]), .Y(n596) );
  NAND2X0_HVT U1758 ( .A1(conv2_sum_b[7]), .A2(n473), .Y(n593) );
  NAND2X0_HVT U1759 ( .A1(conv2_sum_a[6]), .A2(n593), .Y(n594) );
  OA22X1_HVT U1760 ( .A1(n473), .A2(conv2_sum_b[7]), .A3(n594), .A4(
        conv2_sum_b[6]), .Y(n595) );
  OA221X1_HVT U1761 ( .A1(n598), .A2(n597), .A3(n596), .A4(n597), .A5(n595), 
        .Y(n604) );
  OAI21X1_HVT U1762 ( .A1(conv2_sum_a[16]), .A2(n493), .A3(n599), .Y(n600) );
  OR3X1_HVT U1763 ( .A1(n602), .A2(n601), .A3(n600), .Y(n603) );
  AO221X1_HVT U1764 ( .A1(n606), .A2(n605), .A3(n606), .A4(n604), .A5(n603), 
        .Y(n607) );
  NAND2X0_HVT U1765 ( .A1(n608), .A2(n607), .Y(n609) );
  NAND4X0_HVT U1766 ( .A1(n612), .A2(n611), .A3(n610), .A4(n609), .Y(n613) );
  OA221X1_HVT U1767 ( .A1(n555), .A2(n558), .A3(n556), .A4(n557), .A5(n554), 
        .Y(n614) );
  OA221X1_HVT U1768 ( .A1(n565), .A2(n601), .A3(n566), .A4(n567), .A5(n564), 
        .Y(n608) );
  OA221X1_HVT U1769 ( .A1(n581), .A2(n576), .A3(n577), .A4(n578), .A5(n575), 
        .Y(n606) );
  AO22X1_HVT U1770 ( .A1(conv2_sum_d[30]), .A2(n528), .A3(conv2_sum_c[31]), 
        .A4(n530), .Y(n622) );
  NAND2X0_HVT U1771 ( .A1(conv2_sum_d[29]), .A2(n526), .Y(n616) );
  NAND2X0_HVT U1772 ( .A1(conv2_sum_c[28]), .A2(n616), .Y(n615) );
  OA22X1_HVT U1773 ( .A1(n526), .A2(conv2_sum_d[29]), .A3(n615), .A4(
        conv2_sum_d[28]), .Y(n621) );
  NAND2X0_HVT U1774 ( .A1(conv2_sum_d[25]), .A2(n518), .Y(n673) );
  AO22X1_HVT U1775 ( .A1(conv2_sum_d[26]), .A2(n521), .A3(conv2_sum_d[27]), 
        .A4(n525), .Y(n624) );
  NAND2X0_HVT U1776 ( .A1(conv2_sum_c[31]), .A2(n530), .Y(n617) );
  NAND2X0_HVT U1777 ( .A1(conv2_sum_c[30]), .A2(n617), .Y(n618) );
  OA22X1_HVT U1778 ( .A1(n530), .A2(conv2_sum_c[31]), .A3(n618), .A4(
        conv2_sum_d[30]), .Y(n619) );
  NAND2X0_HVT U1779 ( .A1(conv2_sum_d[24]), .A2(n504), .Y(n674) );
  AO22X1_HVT U1780 ( .A1(conv2_sum_d[22]), .A2(n503), .A3(conv2_sum_d[23]), 
        .A4(n517), .Y(n632) );
  NAND2X0_HVT U1781 ( .A1(conv2_sum_d[21]), .A2(n516), .Y(n626) );
  NAND2X0_HVT U1782 ( .A1(conv2_sum_c[20]), .A2(n626), .Y(n625) );
  OA22X1_HVT U1783 ( .A1(n516), .A2(conv2_sum_d[21]), .A3(n625), .A4(
        conv2_sum_d[20]), .Y(n631) );
  NAND2X0_HVT U1784 ( .A1(conv2_sum_d[17]), .A2(n514), .Y(n664) );
  AO22X1_HVT U1785 ( .A1(conv2_sum_d[18]), .A2(n485), .A3(conv2_sum_d[19]), 
        .A4(n515), .Y(n666) );
  NAND2X0_HVT U1786 ( .A1(conv2_sum_d[23]), .A2(n517), .Y(n627) );
  NAND2X0_HVT U1787 ( .A1(conv2_sum_c[22]), .A2(n627), .Y(n628) );
  OA22X1_HVT U1788 ( .A1(n517), .A2(conv2_sum_d[23]), .A3(n628), .A4(
        conv2_sum_d[22]), .Y(n629) );
  AO22X1_HVT U1789 ( .A1(conv2_sum_d[14]), .A2(n501), .A3(conv2_sum_d[15]), 
        .A4(n513), .Y(n645) );
  NAND2X0_HVT U1790 ( .A1(conv2_sum_d[13]), .A2(n512), .Y(n634) );
  NAND2X0_HVT U1791 ( .A1(conv2_sum_c[12]), .A2(n634), .Y(n633) );
  OA22X1_HVT U1792 ( .A1(n512), .A2(conv2_sum_d[13]), .A3(n633), .A4(
        conv2_sum_d[12]), .Y(n644) );
  NAND2X0_HVT U1793 ( .A1(conv2_sum_d[11]), .A2(n476), .Y(n635) );
  NAND2X0_HVT U1794 ( .A1(conv2_sum_c[10]), .A2(n635), .Y(n636) );
  OA22X1_HVT U1795 ( .A1(conv2_sum_d[11]), .A2(n476), .A3(conv2_sum_d[10]), 
        .A4(n636), .Y(n639) );
  NAND2X0_HVT U1796 ( .A1(conv2_sum_d[9]), .A2(n489), .Y(n646) );
  NAND2X0_HVT U1797 ( .A1(conv2_sum_c[8]), .A2(n646), .Y(n637) );
  OA22X1_HVT U1798 ( .A1(n489), .A2(conv2_sum_d[9]), .A3(n637), .A4(
        conv2_sum_d[8]), .Y(n638) );
  AO22X1_HVT U1799 ( .A1(conv2_sum_d[10]), .A2(n486), .A3(conv2_sum_d[11]), 
        .A4(n476), .Y(n649) );
  AO22X1_HVT U1800 ( .A1(n639), .A2(n638), .A3(n639), .A4(n649), .Y(n643) );
  NAND2X0_HVT U1801 ( .A1(conv2_sum_d[15]), .A2(n513), .Y(n640) );
  NAND2X0_HVT U1802 ( .A1(conv2_sum_c[14]), .A2(n640), .Y(n641) );
  OA22X1_HVT U1803 ( .A1(n513), .A2(conv2_sum_d[15]), .A3(n641), .A4(
        conv2_sum_d[14]), .Y(n642) );
  OAI21X1_HVT U1804 ( .A1(conv2_sum_c[8]), .A2(n478), .A3(n646), .Y(n647) );
  OR3X1_HVT U1805 ( .A1(n649), .A2(n648), .A3(n647), .Y(n667) );
  NAND2X0_HVT U1806 ( .A1(conv2_sum_c[2]), .A2(n650), .Y(n651) );
  OA22X1_HVT U1807 ( .A1(conv2_sum_d[3]), .A2(n490), .A3(conv2_sum_d[2]), .A4(
        n651), .Y(n657) );
  NAND2X0_HVT U1808 ( .A1(n543), .A2(conv2_sum_c[1]), .Y(n652) );
  NAND2X0_HVT U1809 ( .A1(conv2_sum_d[0]), .A2(n652), .Y(n653) );
  OAI22X1_HVT U1810 ( .A1(conv2_sum_c[0]), .A2(n653), .A3(n543), .A4(
        conv2_sum_c[1]), .Y(n655) );
  AO22X1_HVT U1811 ( .A1(conv2_sum_d[5]), .A2(n474), .A3(conv2_sum_d[4]), .A4(
        n480), .Y(n654) );
  AO221X1_HVT U1812 ( .A1(n657), .A2(n656), .A3(n657), .A4(n655), .A5(n654), 
        .Y(n663) );
  NAND2X0_HVT U1813 ( .A1(conv2_sum_d[5]), .A2(n474), .Y(n658) );
  NAND2X0_HVT U1814 ( .A1(conv2_sum_c[4]), .A2(n658), .Y(n659) );
  OA22X1_HVT U1815 ( .A1(n659), .A2(conv2_sum_d[4]), .A3(n474), .A4(
        conv2_sum_d[5]), .Y(n662) );
  NAND2X0_HVT U1816 ( .A1(conv2_sum_d[7]), .A2(n475), .Y(n660) );
  NAND2X0_HVT U1817 ( .A1(conv2_sum_c[6]), .A2(n660), .Y(n661) );
  NAND2X0_HVT U1818 ( .A1(n669), .A2(n670), .Y(n671) );
  NAND4X0_HVT U1819 ( .A1(n671), .A2(n673), .A3(n672), .A4(n674), .Y(n675) );
  OA221X1_HVT U1820 ( .A1(n620), .A2(n623), .A3(n621), .A4(n622), .A5(n619), 
        .Y(n676) );
  OA221X1_HVT U1821 ( .A1(n630), .A2(n665), .A3(n631), .A4(n632), .A5(n629), 
        .Y(n670) );
  OA221X1_HVT U1822 ( .A1(n643), .A2(n648), .A3(n644), .A4(n645), .A5(n642), 
        .Y(n668) );
  AO22X1_HVT U1823 ( .A1(tmp_big2[30]), .A2(n759), .A3(tmp_big1[31]), .A4(n739), .Y(n685) );
  NAND2X0_HVT U1824 ( .A1(tmp_big2[29]), .A2(n757), .Y(n678) );
  NAND2X0_HVT U1825 ( .A1(tmp_big1[28]), .A2(n678), .Y(n677) );
  OA22X1_HVT U1826 ( .A1(n757), .A2(tmp_big2[29]), .A3(n677), .A4(tmp_big2[28]), .Y(n684) );
  NAND2X0_HVT U1827 ( .A1(tmp_big2[27]), .A2(n756), .Y(n679) );
  NAND2X0_HVT U1828 ( .A1(tmp_big2[25]), .A2(n754), .Y(n736) );
  AO22X1_HVT U1829 ( .A1(tmp_big2[26]), .A2(n755), .A3(tmp_big2[27]), .A4(n756), .Y(n687) );
  NAND2X0_HVT U1830 ( .A1(tmp_big1[31]), .A2(n739), .Y(n680) );
  NAND2X0_HVT U1831 ( .A1(tmp_big1[30]), .A2(n680), .Y(n681) );
  OA22X1_HVT U1832 ( .A1(n739), .A2(tmp_big1[31]), .A3(n681), .A4(tmp_big2[30]), .Y(n682) );
  AO22X1_HVT U1833 ( .A1(tmp_big2[22]), .A2(n752), .A3(tmp_big2[23]), .A4(n753), .Y(n698) );
  NAND2X0_HVT U1834 ( .A1(tmp_big2[21]), .A2(n751), .Y(n689) );
  NAND2X0_HVT U1835 ( .A1(tmp_big1[20]), .A2(n689), .Y(n688) );
  OA22X1_HVT U1836 ( .A1(n751), .A2(tmp_big2[21]), .A3(n688), .A4(tmp_big2[20]), .Y(n697) );
  NAND2X0_HVT U1837 ( .A1(tmp_big2[19]), .A2(n750), .Y(n690) );
  NAND2X0_HVT U1838 ( .A1(tmp_big1[18]), .A2(n690), .Y(n691) );
  NAND2X0_HVT U1839 ( .A1(tmp_big2[17]), .A2(n748), .Y(n729) );
  NAND2X0_HVT U1840 ( .A1(tmp_big1[16]), .A2(n729), .Y(n692) );
  AO22X1_HVT U1841 ( .A1(tmp_big2[18]), .A2(n749), .A3(tmp_big2[19]), .A4(n750), .Y(n732) );
  NAND2X0_HVT U1842 ( .A1(tmp_big2[23]), .A2(n753), .Y(n693) );
  NAND2X0_HVT U1843 ( .A1(tmp_big1[22]), .A2(n693), .Y(n694) );
  OA22X1_HVT U1844 ( .A1(n753), .A2(tmp_big2[23]), .A3(n694), .A4(tmp_big2[22]), .Y(n695) );
  AO22X1_HVT U1845 ( .A1(tmp_big2[14]), .A2(n745), .A3(tmp_big2[15]), .A4(n746), .Y(n710) );
  NAND2X0_HVT U1846 ( .A1(tmp_big2[13]), .A2(n744), .Y(n7001) );
  NAND2X0_HVT U1847 ( .A1(tmp_big1[12]), .A2(n7001), .Y(n699) );
  OA22X1_HVT U1848 ( .A1(n744), .A2(tmp_big2[13]), .A3(n699), .A4(tmp_big2[12]), .Y(n709) );
  NAND2X0_HVT U1849 ( .A1(tmp_big2[12]), .A2(n743), .Y(n701) );
  NAND3X0_HVT U1850 ( .A1(n701), .A2(n747), .A3(n7001), .Y(n713) );
  NAND2X0_HVT U1851 ( .A1(tmp_big2[11]), .A2(n742), .Y(n702) );
  NAND2X0_HVT U1852 ( .A1(tmp_big1[10]), .A2(n702), .Y(n703) );
  NAND2X0_HVT U1853 ( .A1(n547), .A2(tmp_big2[9]), .Y(n711) );
  NAND2X0_HVT U1854 ( .A1(tmp_big1[8]), .A2(n711), .Y(n704) );
  AO22X1_HVT U1855 ( .A1(tmp_big2[10]), .A2(n741), .A3(tmp_big2[11]), .A4(n742), .Y(n714) );
  NAND2X0_HVT U1856 ( .A1(tmp_big2[15]), .A2(n746), .Y(n705) );
  NAND2X0_HVT U1857 ( .A1(tmp_big1[14]), .A2(n705), .Y(n706) );
  OA22X1_HVT U1858 ( .A1(n746), .A2(tmp_big2[15]), .A3(n706), .A4(tmp_big2[14]), .Y(n707) );
  OAI21X1_HVT U1859 ( .A1(tmp_big1[8]), .A2(n740), .A3(n711), .Y(n712) );
  NAND2X0_HVT U1860 ( .A1(tmp_big2[3]), .A2(n465), .Y(n715) );
  NAND2X0_HVT U1861 ( .A1(tmp_big1[2]), .A2(n715), .Y(n716) );
  OA22X1_HVT U1862 ( .A1(tmp_big2[3]), .A2(n465), .A3(tmp_big2[2]), .A4(n716), 
        .Y(n722) );
  NAND2X0_HVT U1863 ( .A1(n542), .A2(tmp_big1[1]), .Y(n717) );
  NAND2X0_HVT U1864 ( .A1(tmp_big2[0]), .A2(n717), .Y(n718) );
  OAI22X1_HVT U1865 ( .A1(tmp_big1[0]), .A2(n718), .A3(n542), .A4(tmp_big1[1]), 
        .Y(n720) );
  AO22X1_HVT U1866 ( .A1(tmp_big2[5]), .A2(n761), .A3(tmp_big2[4]), .A4(n760), 
        .Y(n719) );
  AO221X1_HVT U1867 ( .A1(n722), .A2(n721), .A3(n722), .A4(n720), .A5(n719), 
        .Y(n728) );
  NAND2X0_HVT U1868 ( .A1(tmp_big2[5]), .A2(n761), .Y(n723) );
  NAND2X0_HVT U1869 ( .A1(tmp_big1[4]), .A2(n723), .Y(n724) );
  OA22X1_HVT U1870 ( .A1(n724), .A2(tmp_big2[4]), .A3(n761), .A4(tmp_big2[5]), 
        .Y(n727) );
  NAND2X0_HVT U1871 ( .A1(tmp_big2[7]), .A2(n763), .Y(n725) );
  NAND2X0_HVT U1872 ( .A1(tmp_big1[6]), .A2(n725), .Y(n726) );
  OR3X1_HVT U1873 ( .A1(n732), .A2(n731), .A3(n730), .Y(n733) );
  OA221X1_HVT U1874 ( .A1(n683), .A2(n686), .A3(n684), .A4(n685), .A5(n682), 
        .Y(n737) );
  OA221X1_HVT U1875 ( .A1(n696), .A2(n731), .A3(n697), .A4(n698), .A5(n695), 
        .Y(n735) );
  OA221X1_HVT U1876 ( .A1(n713), .A2(n708), .A3(n709), .A4(n710), .A5(n707), 
        .Y(n734) );
  OR3X1_HVT U1877 ( .A1(channel[4]), .A2(channel[0]), .A3(channel[1]), .Y(n764) );
  OR3X1_HVT U1878 ( .A1(channel[2]), .A2(channel[3]), .A3(n764), .Y(n765) );
  MUX21X1_HVT U1879 ( .A1(conv2_sum_b[29]), .A2(conv2_sum_a[29]), .S0(n414), 
        .Y(tmp_big1[29]) );
  MUX21X1_HVT U1880 ( .A1(conv2_sum_b[28]), .A2(conv2_sum_a[28]), .S0(n413), 
        .Y(tmp_big1[28]) );
  MUX21X1_HVT U1881 ( .A1(conv2_sum_b[27]), .A2(conv2_sum_a[27]), .S0(n413), 
        .Y(tmp_big1[27]) );
  MUX21X1_HVT U1882 ( .A1(conv2_sum_b[26]), .A2(conv2_sum_a[26]), .S0(n415), 
        .Y(tmp_big1[26]) );
  MUX21X1_HVT U1883 ( .A1(conv2_sum_b[25]), .A2(conv2_sum_a[25]), .S0(n415), 
        .Y(tmp_big1[25]) );
  MUX21X1_HVT U1884 ( .A1(conv2_sum_b[24]), .A2(conv2_sum_a[24]), .S0(n414), 
        .Y(tmp_big1[24]) );
  MUX21X1_HVT U1885 ( .A1(conv2_sum_b[23]), .A2(conv2_sum_a[23]), .S0(n414), 
        .Y(tmp_big1[23]) );
  MUX21X1_HVT U1886 ( .A1(conv2_sum_b[22]), .A2(conv2_sum_a[22]), .S0(n414), 
        .Y(tmp_big1[22]) );
  MUX21X1_HVT U1887 ( .A1(conv2_sum_b[21]), .A2(conv2_sum_a[21]), .S0(n413), 
        .Y(tmp_big1[21]) );
  MUX21X1_HVT U1888 ( .A1(conv2_sum_b[20]), .A2(conv2_sum_a[20]), .S0(n414), 
        .Y(tmp_big1[20]) );
  MUX21X1_HVT U1889 ( .A1(conv2_sum_b[18]), .A2(conv2_sum_a[18]), .S0(n412), 
        .Y(tmp_big1[18]) );
  MUX21X1_HVT U1890 ( .A1(conv2_sum_b[16]), .A2(conv2_sum_a[16]), .S0(n413), 
        .Y(tmp_big1[16]) );
  MUX21X1_HVT U1891 ( .A1(conv2_sum_b[15]), .A2(conv2_sum_a[15]), .S0(n415), 
        .Y(tmp_big1[15]) );
  MUX21X1_HVT U1892 ( .A1(conv2_sum_b[14]), .A2(conv2_sum_a[14]), .S0(n414), 
        .Y(tmp_big1[14]) );
  MUX21X1_HVT U1893 ( .A1(conv2_sum_b[13]), .A2(conv2_sum_a[13]), .S0(n415), 
        .Y(tmp_big1[13]) );
  MUX21X1_HVT U1894 ( .A1(conv2_sum_b[12]), .A2(conv2_sum_a[12]), .S0(n415), 
        .Y(tmp_big1[12]) );
  MUX21X1_HVT U1895 ( .A1(conv2_sum_b[10]), .A2(conv2_sum_a[10]), .S0(n415), 
        .Y(tmp_big1[10]) );
  MUX21X1_HVT U1896 ( .A1(conv2_sum_b[8]), .A2(conv2_sum_a[8]), .S0(n414), .Y(
        tmp_big1[8]) );
  MUX21X1_HVT U1897 ( .A1(conv2_sum_d[29]), .A2(conv2_sum_c[29]), .S0(n417), 
        .Y(tmp_big2[29]) );
  MUX21X1_HVT U1898 ( .A1(conv2_sum_d[28]), .A2(conv2_sum_c[28]), .S0(n418), 
        .Y(tmp_big2[28]) );
  MUX21X1_HVT U1899 ( .A1(conv2_sum_d[27]), .A2(conv2_sum_c[27]), .S0(n418), 
        .Y(tmp_big2[27]) );
  MUX21X1_HVT U1900 ( .A1(conv2_sum_d[26]), .A2(conv2_sum_c[26]), .S0(n419), 
        .Y(tmp_big2[26]) );
  MUX21X1_HVT U1901 ( .A1(conv2_sum_d[25]), .A2(conv2_sum_c[25]), .S0(n418), 
        .Y(tmp_big2[25]) );
  MUX21X1_HVT U1902 ( .A1(conv2_sum_d[24]), .A2(conv2_sum_c[24]), .S0(n417), 
        .Y(tmp_big2[24]) );
  MUX21X1_HVT U1903 ( .A1(conv2_sum_d[23]), .A2(conv2_sum_c[23]), .S0(n419), 
        .Y(tmp_big2[23]) );
  MUX21X1_HVT U1904 ( .A1(conv2_sum_d[22]), .A2(conv2_sum_c[22]), .S0(n417), 
        .Y(tmp_big2[22]) );
  MUX21X1_HVT U1905 ( .A1(conv2_sum_d[21]), .A2(conv2_sum_c[21]), .S0(n418), 
        .Y(tmp_big2[21]) );
  MUX21X1_HVT U1906 ( .A1(conv2_sum_d[20]), .A2(conv2_sum_c[20]), .S0(n419), 
        .Y(tmp_big2[20]) );
  MUX21X1_HVT U1907 ( .A1(conv2_sum_d[19]), .A2(conv2_sum_c[19]), .S0(n416), 
        .Y(tmp_big2[19]) );
  MUX21X1_HVT U1908 ( .A1(conv2_sum_d[18]), .A2(conv2_sum_c[18]), .S0(n416), 
        .Y(tmp_big2[18]) );
  MUX21X1_HVT U1909 ( .A1(conv2_sum_d[17]), .A2(conv2_sum_c[17]), .S0(n416), 
        .Y(tmp_big2[17]) );
  MUX21X1_HVT U1910 ( .A1(conv2_sum_d[16]), .A2(conv2_sum_c[16]), .S0(n417), 
        .Y(tmp_big2[16]) );
  MUX21X1_HVT U1911 ( .A1(conv2_sum_d[15]), .A2(conv2_sum_c[15]), .S0(n419), 
        .Y(tmp_big2[15]) );
  MUX21X1_HVT U1912 ( .A1(conv2_sum_d[14]), .A2(conv2_sum_c[14]), .S0(n418), 
        .Y(tmp_big2[14]) );
  MUX21X1_HVT U1913 ( .A1(conv2_sum_d[13]), .A2(conv2_sum_c[13]), .S0(n418), 
        .Y(tmp_big2[13]) );
  MUX21X1_HVT U1914 ( .A1(conv2_sum_d[12]), .A2(conv2_sum_c[12]), .S0(n417), 
        .Y(tmp_big2[12]) );
  MUX21X1_HVT U1915 ( .A1(conv2_sum_d[11]), .A2(conv2_sum_c[11]), .S0(n416), 
        .Y(tmp_big2[11]) );
  MUX21X1_HVT U1916 ( .A1(conv2_sum_d[10]), .A2(conv2_sum_c[10]), .S0(n419), 
        .Y(tmp_big2[10]) );
  MUX21X1_HVT U1917 ( .A1(tmp_big2[0]), .A2(tmp_big1[0]), .S0(n410), .Y(
        data_out[0]) );
  MUX21X1_HVT U1918 ( .A1(tmp_big2[1]), .A2(tmp_big1[1]), .S0(n411), .Y(
        data_out[1]) );
  MUX21X1_HVT U1919 ( .A1(tmp_big2[2]), .A2(tmp_big1[2]), .S0(n411), .Y(
        data_out[2]) );
  MUX21X1_HVT U1920 ( .A1(tmp_big2[3]), .A2(tmp_big1[3]), .S0(n410), .Y(
        data_out[3]) );
  MUX21X1_HVT U1921 ( .A1(tmp_big2[4]), .A2(tmp_big1[4]), .S0(n410), .Y(
        data_out[4]) );
  MUX21X1_HVT U1922 ( .A1(tmp_big2[14]), .A2(tmp_big1[14]), .S0(n471), .Y(
        data_out[14]) );
  MUX21X1_HVT U1923 ( .A1(tmp_big2[16]), .A2(tmp_big1[16]), .S0(n409), .Y(
        data_out[16]) );
  MUX21X1_HVT U1924 ( .A1(tmp_big2[17]), .A2(tmp_big1[17]), .S0(n409), .Y(
        data_out[17]) );
  MUX21X1_HVT U1925 ( .A1(tmp_big2[18]), .A2(tmp_big1[18]), .S0(n409), .Y(
        data_out[18]) );
  MUX21X1_HVT U1926 ( .A1(tmp_big2[19]), .A2(tmp_big1[19]), .S0(n409), .Y(
        data_out[19]) );
  MUX21X1_HVT U1927 ( .A1(tmp_big2[20]), .A2(tmp_big1[20]), .S0(n410), .Y(
        data_out[20]) );
  MUX21X1_HVT U1928 ( .A1(tmp_big2[21]), .A2(tmp_big1[21]), .S0(n411), .Y(
        data_out[21]) );
  MUX21X1_HVT U1929 ( .A1(tmp_big2[24]), .A2(tmp_big1[24]), .S0(n411), .Y(
        data_out[24]) );
  MUX21X1_HVT U1930 ( .A1(tmp_big2[25]), .A2(tmp_big1[25]), .S0(n411), .Y(
        data_out[25]) );
  MUX21X1_HVT U1931 ( .A1(tmp_big2[26]), .A2(tmp_big1[26]), .S0(n410), .Y(
        data_out[26]) );
  MUX21X1_HVT U1932 ( .A1(tmp_big2[27]), .A2(tmp_big1[27]), .S0(n410), .Y(
        data_out[27]) );
  MUX21X1_HVT U1933 ( .A1(tmp_big2[28]), .A2(tmp_big1[28]), .S0(n411), .Y(
        data_out[28]) );
endmodule


module quantize ( clk, srstn, bias_data, mode, quantized_data, ori_data_31_, 
        ori_data_30_, ori_data_29_, ori_data_28_, ori_data_27_, ori_data_26_, 
        ori_data_25_, ori_data_24_, ori_data_23_, ori_data_22_, ori_data_21_, 
        ori_data_20_, ori_data_19_, ori_data_18_, ori_data_17_, ori_data_16_, 
        ori_data_15_, ori_data_14_, ori_data_13_, ori_data_12_, ori_data_11_, 
        ori_data_10_, ori_data_9_, ori_data_8_, ori_data_7_, ori_data_6_, 
        ori_data_5_ );
  input [3:0] bias_data;
  input [1:0] mode;
  output [7:0] quantized_data;
  input clk, srstn, ori_data_31_, ori_data_30_, ori_data_29_, ori_data_28_,
         ori_data_27_, ori_data_26_, ori_data_25_, ori_data_24_, ori_data_23_,
         ori_data_22_, ori_data_21_, ori_data_20_, ori_data_19_, ori_data_18_,
         ori_data_17_, ori_data_16_, ori_data_15_, ori_data_14_, ori_data_13_,
         ori_data_12_, ori_data_11_, ori_data_10_, ori_data_9_, ori_data_8_,
         ori_data_7_, ori_data_6_, ori_data_5_;
  wire   N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, n13, DP_OP_26J6_124_4249_n586,
         DP_OP_26J6_124_4249_n584, DP_OP_26J6_124_4249_n582,
         DP_OP_26J6_124_4249_n580, DP_OP_26J6_124_4249_n576,
         DP_OP_26J6_124_4249_n574, DP_OP_26J6_124_4249_n570,
         DP_OP_26J6_124_4249_n563, DP_OP_26J6_124_4249_n562,
         DP_OP_26J6_124_4249_n561, DP_OP_26J6_124_4249_n560,
         DP_OP_26J6_124_4249_n559, DP_OP_26J6_124_4249_n558,
         DP_OP_26J6_124_4249_n557, DP_OP_26J6_124_4249_n551,
         DP_OP_26J6_124_4249_n550, DP_OP_26J6_124_4249_n549,
         DP_OP_26J6_124_4249_n548, DP_OP_26J6_124_4249_n547,
         DP_OP_26J6_124_4249_n546, DP_OP_26J6_124_4249_n545,
         DP_OP_26J6_124_4249_n544, DP_OP_26J6_124_4249_n536,
         DP_OP_26J6_124_4249_n535, DP_OP_26J6_124_4249_n534,
         DP_OP_26J6_124_4249_n533, DP_OP_26J6_124_4249_n528,
         DP_OP_26J6_124_4249_n527, DP_OP_26J6_124_4249_n526,
         DP_OP_26J6_124_4249_n516, DP_OP_26J6_124_4249_n515,
         DP_OP_26J6_124_4249_n514, DP_OP_26J6_124_4249_n513,
         DP_OP_26J6_124_4249_n512, DP_OP_26J6_124_4249_n511,
         DP_OP_26J6_124_4249_n510, DP_OP_26J6_124_4249_n509,
         DP_OP_26J6_124_4249_n508, DP_OP_26J6_124_4249_n507,
         DP_OP_26J6_124_4249_n497, DP_OP_26J6_124_4249_n496,
         DP_OP_26J6_124_4249_n491, DP_OP_26J6_124_4249_n490,
         DP_OP_26J6_124_4249_n489, DP_OP_26J6_124_4249_n488,
         DP_OP_26J6_124_4249_n486, DP_OP_26J6_124_4249_n485,
         DP_OP_26J6_124_4249_n478, DP_OP_26J6_124_4249_n477,
         DP_OP_26J6_124_4249_n476, DP_OP_26J6_124_4249_n475,
         DP_OP_26J6_124_4249_n474, DP_OP_26J6_124_4249_n473,
         DP_OP_26J6_124_4249_n472, DP_OP_26J6_124_4249_n469,
         DP_OP_26J6_124_4249_n468, DP_OP_26J6_124_4249_n467,
         DP_OP_26J6_124_4249_n466, DP_OP_26J6_124_4249_n464,
         DP_OP_26J6_124_4249_n456, DP_OP_26J6_124_4249_n455,
         DP_OP_26J6_124_4249_n454, DP_OP_26J6_124_4249_n453,
         DP_OP_26J6_124_4249_n452, DP_OP_26J6_124_4249_n447,
         DP_OP_26J6_124_4249_n446, DP_OP_26J6_124_4249_n445,
         DP_OP_26J6_124_4249_n442, DP_OP_26J6_124_4249_n437,
         DP_OP_26J6_124_4249_n435, DP_OP_26J6_124_4249_n434,
         DP_OP_26J6_124_4249_n433, DP_OP_26J6_124_4249_n432,
         DP_OP_26J6_124_4249_n431, DP_OP_26J6_124_4249_n430,
         DP_OP_26J6_124_4249_n429, DP_OP_26J6_124_4249_n428,
         DP_OP_26J6_124_4249_n427, DP_OP_26J6_124_4249_n426,
         DP_OP_26J6_124_4249_n425, DP_OP_26J6_124_4249_n424,
         DP_OP_26J6_124_4249_n422, DP_OP_26J6_124_4249_n421,
         DP_OP_26J6_124_4249_n411, DP_OP_26J6_124_4249_n410,
         DP_OP_26J6_124_4249_n405, DP_OP_26J6_124_4249_n404,
         DP_OP_26J6_124_4249_n403, DP_OP_26J6_124_4249_n402,
         DP_OP_26J6_124_4249_n400, DP_OP_26J6_124_4249_n394,
         DP_OP_26J6_124_4249_n392, DP_OP_26J6_124_4249_n391,
         DP_OP_26J6_124_4249_n389, DP_OP_26J6_124_4249_n388,
         DP_OP_26J6_124_4249_n387, DP_OP_26J6_124_4249_n386,
         DP_OP_26J6_124_4249_n383, DP_OP_26J6_124_4249_n382,
         DP_OP_26J6_124_4249_n381, DP_OP_26J6_124_4249_n380,
         DP_OP_26J6_124_4249_n378, DP_OP_26J6_124_4249_n377,
         DP_OP_26J6_124_4249_n370, DP_OP_26J6_124_4249_n369,
         DP_OP_26J6_124_4249_n367, DP_OP_26J6_124_4249_n366,
         DP_OP_26J6_124_4249_n361, DP_OP_26J6_124_4249_n360,
         DP_OP_26J6_124_4249_n359, DP_OP_26J6_124_4249_n358,
         DP_OP_26J6_124_4249_n356, DP_OP_26J6_124_4249_n351,
         DP_OP_26J6_124_4249_n349, DP_OP_26J6_124_4249_n348,
         DP_OP_26J6_124_4249_n347, DP_OP_26J6_124_4249_n345,
         DP_OP_26J6_124_4249_n344, DP_OP_26J6_124_4249_n343,
         DP_OP_26J6_124_4249_n342, DP_OP_26J6_124_4249_n341,
         DP_OP_26J6_124_4249_n340, DP_OP_26J6_124_4249_n339,
         DP_OP_26J6_124_4249_n338, DP_OP_26J6_124_4249_n337,
         DP_OP_26J6_124_4249_n336, DP_OP_26J6_124_4249_n334,
         DP_OP_26J6_124_4249_n332, DP_OP_26J6_124_4249_n330,
         DP_OP_26J6_124_4249_n329, DP_OP_26J6_124_4249_n328,
         DP_OP_26J6_124_4249_n310, DP_OP_26J6_124_4249_n309,
         DP_OP_26J6_124_4249_n306, DP_OP_26J6_124_4249_n294,
         DP_OP_26J6_124_4249_n289, DP_OP_26J6_124_4249_n287,
         DP_OP_26J6_124_4249_n285, DP_OP_26J6_124_4249_n283,
         DP_OP_26J6_124_4249_n282, DP_OP_26J6_124_4249_n281,
         DP_OP_26J6_124_4249_n279, DP_OP_26J6_124_4249_n277,
         DP_OP_26J6_124_4249_n272, DP_OP_26J6_124_4249_n271,
         DP_OP_26J6_124_4249_n263, DP_OP_26J6_124_4249_n262,
         DP_OP_26J6_124_4249_n261, DP_OP_26J6_124_4249_n260,
         DP_OP_26J6_124_4249_n259, DP_OP_26J6_124_4249_n258,
         DP_OP_26J6_124_4249_n252, DP_OP_26J6_124_4249_n251,
         DP_OP_26J6_124_4249_n250, DP_OP_26J6_124_4249_n249,
         DP_OP_26J6_124_4249_n248, DP_OP_26J6_124_4249_n247,
         DP_OP_26J6_124_4249_n246, DP_OP_26J6_124_4249_n245,
         DP_OP_26J6_124_4249_n240, DP_OP_26J6_124_4249_n238,
         DP_OP_26J6_124_4249_n237, DP_OP_26J6_124_4249_n236,
         DP_OP_26J6_124_4249_n233, DP_OP_26J6_124_4249_n231,
         DP_OP_26J6_124_4249_n230, DP_OP_26J6_124_4249_n228,
         DP_OP_26J6_124_4249_n223, DP_OP_26J6_124_4249_n219,
         DP_OP_26J6_124_4249_n218, DP_OP_26J6_124_4249_n217,
         DP_OP_26J6_124_4249_n216, DP_OP_26J6_124_4249_n215,
         DP_OP_26J6_124_4249_n214, DP_OP_26J6_124_4249_n213,
         DP_OP_26J6_124_4249_n212, DP_OP_26J6_124_4249_n211,
         DP_OP_26J6_124_4249_n210, DP_OP_26J6_124_4249_n200,
         DP_OP_26J6_124_4249_n199, DP_OP_26J6_124_4249_n194,
         DP_OP_26J6_124_4249_n193, DP_OP_26J6_124_4249_n192,
         DP_OP_26J6_124_4249_n191, DP_OP_26J6_124_4249_n189,
         DP_OP_26J6_124_4249_n188, DP_OP_26J6_124_4249_n181,
         DP_OP_26J6_124_4249_n180, DP_OP_26J6_124_4249_n178,
         DP_OP_26J6_124_4249_n177, DP_OP_26J6_124_4249_n176,
         DP_OP_26J6_124_4249_n175, DP_OP_26J6_124_4249_n172,
         DP_OP_26J6_124_4249_n171, DP_OP_26J6_124_4249_n170,
         DP_OP_26J6_124_4249_n169, DP_OP_26J6_124_4249_n167,
         DP_OP_26J6_124_4249_n166, DP_OP_26J6_124_4249_n161,
         DP_OP_26J6_124_4249_n156, DP_OP_26J6_124_4249_n155,
         DP_OP_26J6_124_4249_n152, DP_OP_26J6_124_4249_n150,
         DP_OP_26J6_124_4249_n149, DP_OP_26J6_124_4249_n148,
         DP_OP_26J6_124_4249_n147, DP_OP_26J6_124_4249_n145,
         DP_OP_26J6_124_4249_n140, DP_OP_26J6_124_4249_n139,
         DP_OP_26J6_124_4249_n138, DP_OP_26J6_124_4249_n134,
         DP_OP_26J6_124_4249_n133, DP_OP_26J6_124_4249_n132,
         DP_OP_26J6_124_4249_n131, DP_OP_26J6_124_4249_n130,
         DP_OP_26J6_124_4249_n129, DP_OP_26J6_124_4249_n128,
         DP_OP_26J6_124_4249_n127, DP_OP_26J6_124_4249_n123,
         DP_OP_26J6_124_4249_n117, DP_OP_26J6_124_4249_n116,
         DP_OP_26J6_124_4249_n107, DP_OP_26J6_124_4249_n106,
         DP_OP_26J6_124_4249_n105, DP_OP_26J6_124_4249_n103,
         DP_OP_26J6_124_4249_n102, DP_OP_26J6_124_4249_n96,
         DP_OP_26J6_124_4249_n95, DP_OP_26J6_124_4249_n92,
         DP_OP_26J6_124_4249_n91, DP_OP_26J6_124_4249_n84,
         DP_OP_26J6_124_4249_n83, DP_OP_26J6_124_4249_n81,
         DP_OP_26J6_124_4249_n80, DP_OP_26J6_124_4249_n74,
         DP_OP_26J6_124_4249_n73, DP_OP_26J6_124_4249_n72,
         DP_OP_26J6_124_4249_n71, DP_OP_26J6_124_4249_n70,
         DP_OP_26J6_124_4249_n69, DP_OP_26J6_124_4249_n64,
         DP_OP_26J6_124_4249_n63, DP_OP_26J6_124_4249_n62,
         DP_OP_26J6_124_4249_n61, DP_OP_26J6_124_4249_n60,
         DP_OP_26J6_124_4249_n59, DP_OP_26J6_124_4249_n54,
         DP_OP_26J6_124_4249_n52, DP_OP_26J6_124_4249_n51,
         DP_OP_26J6_124_4249_n48, DP_OP_26J6_124_4249_n47,
         DP_OP_26J6_124_4249_n45, DP_OP_26J6_124_4249_n40,
         DP_OP_26J6_124_4249_n39, DP_OP_26J6_124_4249_n38,
         DP_OP_26J6_124_4249_n37, DP_OP_26J6_124_4249_n35,
         DP_OP_26J6_124_4249_n33, DP_OP_26J6_124_4249_n32,
         DP_OP_26J6_124_4249_n24, DP_OP_26J6_124_4249_n8,
         DP_OP_26J6_124_4249_n7, DP_OP_26J6_124_4249_n4,
         DP_OP_26J6_124_4249_n3, DP_OP_26J6_124_4249_n2,
         DP_OP_26J6_124_4249_n1, n1, n2, n3, n4, n5, n6, n7, n9, n10, n11, n12,
         n14, n15, n16, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n33, n34, n35, n360, n370, n380, n390, n410, n420,
         n430, n440, n450, n460, n470, n490, n500, n510, n520, n530, n540,
         n550, n560, n570, n580, n590, n600, n610, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n1070, n1080,
         n1090, n1100, n1110, n1120, n1130, n1140, n1150, n1160, n1170, n1180,
         n1190, n1200, n1210, n1220, n1230, n1240, n1250, n1260, n1270, n1280,
         n1290, n1300, n1310, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202;
  wire   [7:0] n_quantized_data;

  DFFSSRX1_HVT quantized_data_reg_7_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[7]), .CLK(clk), .Q(quantized_data[7]) );
  DFFSSRX1_HVT quantized_data_reg_6_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[6]), .CLK(clk), .Q(quantized_data[6]) );
  DFFSSRX1_HVT quantized_data_reg_5_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[5]), .CLK(clk), .Q(quantized_data[5]) );
  DFFSSRX1_HVT quantized_data_reg_4_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[4]), .CLK(clk), .Q(quantized_data[4]) );
  DFFSSRX1_HVT quantized_data_reg_3_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[3]), .CLK(clk), .Q(quantized_data[3]) );
  DFFSSRX1_HVT quantized_data_reg_2_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[2]), .CLK(clk), .Q(quantized_data[2]) );
  DFFSSRX1_HVT quantized_data_reg_1_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[1]), .CLK(clk), .Q(quantized_data[1]) );
  DFFSSRX1_HVT quantized_data_reg_0_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[0]), .CLK(clk), .Q(quantized_data[0]) );
  XOR2X1_HVT DP_OP_26J6_124_4249_U262 ( .A1(DP_OP_26J6_124_4249_n238), .A2(
        DP_OP_26J6_124_4249_n24), .Y(N111) );
  XOR2X1_HVT DP_OP_26J6_124_4249_U305 ( .A1(DP_OP_26J6_124_4249_n263), .A2(
        DP_OP_26J6_124_4249_n262), .Y(N107) );
  OAI21X2_HVT DP_OP_26J6_124_4249_U350 ( .A1(DP_OP_26J6_124_4249_n340), .A2(
        DP_OP_26J6_124_4249_n381), .A3(DP_OP_26J6_124_4249_n341), .Y(
        DP_OP_26J6_124_4249_n339) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U620 ( .A1(DP_OP_26J6_124_4249_n558), .A2(
        DP_OP_26J6_124_4249_n550), .A3(DP_OP_26J6_124_4249_n551), .Y(
        DP_OP_26J6_124_4249_n549) );
  OAI21X2_HVT DP_OP_26J6_124_4249_U132 ( .A1(DP_OP_26J6_124_4249_n129), .A2(
        DP_OP_26J6_124_4249_n170), .A3(DP_OP_26J6_124_4249_n130), .Y(
        DP_OP_26J6_124_4249_n128) );
  OAI21X2_HVT DP_OP_26J6_124_4249_U569 ( .A1(DP_OP_26J6_124_4249_n511), .A2(
        DP_OP_26J6_124_4249_n547), .A3(DP_OP_26J6_124_4249_n512), .Y(
        DP_OP_26J6_124_4249_n510) );
  XNOR2X2_HVT DP_OP_26J6_124_4249_U31 ( .A1(DP_OP_26J6_124_4249_n60), .A2(
        DP_OP_26J6_124_4249_n7), .Y(N128) );
  OAI21X2_HVT DP_OP_26J6_124_4249_U241 ( .A1(DP_OP_26J6_124_4249_n214), .A2(
        DP_OP_26J6_124_4249_n248), .A3(DP_OP_26J6_124_4249_n215), .Y(
        DP_OP_26J6_124_4249_n213) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U470 ( .A1(DP_OP_26J6_124_4249_n433), .A2(
        DP_OP_26J6_124_4249_n509), .A3(DP_OP_26J6_124_4249_n434), .Y(
        DP_OP_26J6_124_4249_n432) );
  XNOR2X1_HVT DP_OP_26J6_124_4249_U511 ( .A1(DP_OP_26J6_124_4249_n476), .A2(
        DP_OP_26J6_124_4249_n310), .Y(N46) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U354 ( .A1(DP_OP_26J6_124_4249_n356), .A2(
        DP_OP_26J6_124_4249_n344), .A3(DP_OP_26J6_124_4249_n345), .Y(
        DP_OP_26J6_124_4249_n343) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U382 ( .A1(DP_OP_26J6_124_4249_n378), .A2(
        DP_OP_26J6_124_4249_n366), .A3(DP_OP_26J6_124_4249_n367), .Y(
        DP_OP_26J6_124_4249_n361) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U410 ( .A1(DP_OP_26J6_124_4249_n400), .A2(
        DP_OP_26J6_124_4249_n388), .A3(DP_OP_26J6_124_4249_n389), .Y(
        DP_OP_26J6_124_4249_n387) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U438 ( .A1(DP_OP_26J6_124_4249_n422), .A2(
        DP_OP_26J6_124_4249_n410), .A3(DP_OP_26J6_124_4249_n411), .Y(
        DP_OP_26J6_124_4249_n405) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U464 ( .A1(DP_OP_26J6_124_4249_n442), .A2(
        DP_OP_26J6_124_4249_n430), .A3(DP_OP_26J6_124_4249_n431), .Y(
        DP_OP_26J6_124_4249_n429) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U492 ( .A1(DP_OP_26J6_124_4249_n464), .A2(
        DP_OP_26J6_124_4249_n452), .A3(DP_OP_26J6_124_4249_n453), .Y(
        DP_OP_26J6_124_4249_n447) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U520 ( .A1(DP_OP_26J6_124_4249_n486), .A2(
        DP_OP_26J6_124_4249_n474), .A3(DP_OP_26J6_124_4249_n475), .Y(
        DP_OP_26J6_124_4249_n473) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U548 ( .A1(DP_OP_26J6_124_4249_n508), .A2(
        DP_OP_26J6_124_4249_n496), .A3(DP_OP_26J6_124_4249_n497), .Y(
        DP_OP_26J6_124_4249_n491) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U573 ( .A1(DP_OP_26J6_124_4249_n527), .A2(
        DP_OP_26J6_124_4249_n515), .A3(DP_OP_26J6_124_4249_n516), .Y(
        DP_OP_26J6_124_4249_n514) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U146 ( .A1(DP_OP_26J6_124_4249_n140), .A2(
        DP_OP_26J6_124_4249_n152), .A3(DP_OP_26J6_124_4249_n145), .Y(
        DP_OP_26J6_124_4249_n139) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U54 ( .A1(DP_OP_26J6_124_4249_n81), .A2(
        DP_OP_26J6_124_4249_n69), .A3(DP_OP_26J6_124_4249_n70), .Y(
        DP_OP_26J6_124_4249_n64) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U136 ( .A1(DP_OP_26J6_124_4249_n145), .A2(
        DP_OP_26J6_124_4249_n133), .A3(DP_OP_26J6_124_4249_n134), .Y(
        DP_OP_26J6_124_4249_n132) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U164 ( .A1(DP_OP_26J6_124_4249_n167), .A2(
        DP_OP_26J6_124_4249_n155), .A3(DP_OP_26J6_124_4249_n156), .Y(
        DP_OP_26J6_124_4249_n150) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U192 ( .A1(DP_OP_26J6_124_4249_n189), .A2(
        DP_OP_26J6_124_4249_n177), .A3(DP_OP_26J6_124_4249_n178), .Y(
        DP_OP_26J6_124_4249_n176) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U220 ( .A1(DP_OP_26J6_124_4249_n211), .A2(
        DP_OP_26J6_124_4249_n199), .A3(DP_OP_26J6_124_4249_n200), .Y(
        DP_OP_26J6_124_4249_n194) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U245 ( .A1(DP_OP_26J6_124_4249_n228), .A2(
        DP_OP_26J6_124_4249_n218), .A3(DP_OP_26J6_124_4249_n219), .Y(
        DP_OP_26J6_124_4249_n217) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U290 ( .A1(DP_OP_26J6_124_4249_n259), .A2(
        DP_OP_26J6_124_4249_n251), .A3(DP_OP_26J6_124_4249_n252), .Y(
        DP_OP_26J6_124_4249_n250) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U641 ( .A1(ori_data_6_), .A2(bias_data[1]), 
        .Y(DP_OP_26J6_124_4249_n562) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U640 ( .A1(bias_data[1]), .A2(ori_data_6_), 
        .Y(DP_OP_26J6_124_4249_n561) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U634 ( .A1(ori_data_7_), .A2(bias_data[2]), 
        .Y(DP_OP_26J6_124_4249_n558) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U633 ( .A1(bias_data[2]), .A2(ori_data_7_), 
        .Y(DP_OP_26J6_124_4249_n557) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U624 ( .A1(ori_data_8_), .A2(n1290), .Y(
        DP_OP_26J6_124_4249_n551) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U619 ( .A1(DP_OP_26J6_124_4249_n557), .A2(
        DP_OP_26J6_124_4249_n550), .Y(DP_OP_26J6_124_4249_n548) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U618 ( .A1(DP_OP_26J6_124_4249_n560), .A2(
        DP_OP_26J6_124_4249_n548), .A3(DP_OP_26J6_124_4249_n549), .Y(
        DP_OP_26J6_124_4249_n547) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U615 ( .A1(ori_data_9_), .A2(n1290), .Y(
        DP_OP_26J6_124_4249_n545) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U603 ( .A1(ori_data_10_), .A2(n1260), .Y(
        DP_OP_26J6_124_4249_n536) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U602 ( .A1(n1260), .A2(ori_data_10_), .Y(
        DP_OP_26J6_124_4249_n535) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U598 ( .A1(DP_OP_26J6_124_4249_n544), .A2(
        DP_OP_26J6_124_4249_n535), .Y(DP_OP_26J6_124_4249_n533) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U591 ( .A1(ori_data_11_), .A2(n1280), .Y(
        DP_OP_26J6_124_4249_n527) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U577 ( .A1(ori_data_12_), .A2(n1280), .Y(
        DP_OP_26J6_124_4249_n516) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U576 ( .A1(n1260), .A2(ori_data_12_), .Y(
        DP_OP_26J6_124_4249_n515) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U572 ( .A1(DP_OP_26J6_124_4249_n515), .A2(
        DP_OP_26J6_124_4249_n526), .Y(DP_OP_26J6_124_4249_n513) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U571 ( .A1(DP_OP_26J6_124_4249_n534), .A2(
        DP_OP_26J6_124_4249_n513), .A3(DP_OP_26J6_124_4249_n514), .Y(
        DP_OP_26J6_124_4249_n512) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U570 ( .A1(DP_OP_26J6_124_4249_n533), .A2(
        DP_OP_26J6_124_4249_n513), .Y(DP_OP_26J6_124_4249_n511) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U566 ( .A1(ori_data_13_), .A2(n1270), .Y(
        DP_OP_26J6_124_4249_n508) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U552 ( .A1(ori_data_14_), .A2(n1280), .Y(
        DP_OP_26J6_124_4249_n497) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U551 ( .A1(n1270), .A2(ori_data_14_), .Y(
        DP_OP_26J6_124_4249_n496) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U547 ( .A1(DP_OP_26J6_124_4249_n496), .A2(
        DP_OP_26J6_124_4249_n507), .Y(DP_OP_26J6_124_4249_n490) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U538 ( .A1(ori_data_15_), .A2(n1260), .Y(
        DP_OP_26J6_124_4249_n486) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U537 ( .A1(n1280), .A2(ori_data_15_), .Y(
        DP_OP_26J6_124_4249_n485) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U527 ( .A1(DP_OP_26J6_124_4249_n490), .A2(
        DP_OP_26J6_124_4249_n580), .Y(DP_OP_26J6_124_4249_n477) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U524 ( .A1(ori_data_16_), .A2(n1270), .Y(
        DP_OP_26J6_124_4249_n475) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U523 ( .A1(n1290), .A2(ori_data_16_), .Y(
        DP_OP_26J6_124_4249_n474) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U521 ( .A1(DP_OP_26J6_124_4249_n283), .A2(
        DP_OP_26J6_124_4249_n475), .Y(DP_OP_26J6_124_4249_n310) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U519 ( .A1(DP_OP_26J6_124_4249_n474), .A2(
        DP_OP_26J6_124_4249_n485), .Y(DP_OP_26J6_124_4249_n472) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U518 ( .A1(DP_OP_26J6_124_4249_n491), .A2(
        DP_OP_26J6_124_4249_n472), .A3(DP_OP_26J6_124_4249_n473), .Y(
        DP_OP_26J6_124_4249_n467) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U517 ( .A1(DP_OP_26J6_124_4249_n490), .A2(
        DP_OP_26J6_124_4249_n472), .Y(DP_OP_26J6_124_4249_n466) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U510 ( .A1(ori_data_17_), .A2(n1260), .Y(
        DP_OP_26J6_124_4249_n464) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U507 ( .A1(DP_OP_26J6_124_4249_n282), .A2(
        DP_OP_26J6_124_4249_n464), .Y(DP_OP_26J6_124_4249_n309) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U499 ( .A1(DP_OP_26J6_124_4249_n468), .A2(
        DP_OP_26J6_124_4249_n282), .Y(DP_OP_26J6_124_4249_n455) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U496 ( .A1(ori_data_18_), .A2(n1270), .Y(
        DP_OP_26J6_124_4249_n453) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U495 ( .A1(n1280), .A2(ori_data_18_), .Y(
        DP_OP_26J6_124_4249_n452) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U486 ( .A1(DP_OP_26J6_124_4249_n469), .A2(
        DP_OP_26J6_124_4249_n446), .A3(DP_OP_26J6_124_4249_n447), .Y(
        DP_OP_26J6_124_4249_n445) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U482 ( .A1(ori_data_19_), .A2(n1290), .Y(
        DP_OP_26J6_124_4249_n442) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U481 ( .A1(n1290), .A2(ori_data_19_), .Y(
        DP_OP_26J6_124_4249_n437) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U471 ( .A1(DP_OP_26J6_124_4249_n435), .A2(
        DP_OP_26J6_124_4249_n468), .Y(DP_OP_26J6_124_4249_n433) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U468 ( .A1(ori_data_20_), .A2(n1260), .Y(
        DP_OP_26J6_124_4249_n431) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U467 ( .A1(n1290), .A2(ori_data_20_), .Y(
        DP_OP_26J6_124_4249_n430) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U465 ( .A1(DP_OP_26J6_124_4249_n279), .A2(
        DP_OP_26J6_124_4249_n431), .Y(DP_OP_26J6_124_4249_n306) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U463 ( .A1(DP_OP_26J6_124_4249_n430), .A2(
        DP_OP_26J6_124_4249_n437), .Y(DP_OP_26J6_124_4249_n428) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U462 ( .A1(DP_OP_26J6_124_4249_n447), .A2(
        DP_OP_26J6_124_4249_n428), .A3(DP_OP_26J6_124_4249_n429), .Y(
        DP_OP_26J6_124_4249_n427) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U461 ( .A1(DP_OP_26J6_124_4249_n446), .A2(
        DP_OP_26J6_124_4249_n428), .Y(DP_OP_26J6_124_4249_n426) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U456 ( .A1(ori_data_21_), .A2(n1270), .Y(
        DP_OP_26J6_124_4249_n422) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U455 ( .A1(n1270), .A2(ori_data_21_), .Y(
        DP_OP_26J6_124_4249_n421) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U442 ( .A1(ori_data_22_), .A2(n1260), .Y(
        DP_OP_26J6_124_4249_n411) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U437 ( .A1(DP_OP_26J6_124_4249_n410), .A2(
        DP_OP_26J6_124_4249_n421), .Y(DP_OP_26J6_124_4249_n404) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U428 ( .A1(ori_data_23_), .A2(n1280), .Y(
        DP_OP_26J6_124_4249_n400) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U418 ( .A1(DP_OP_26J6_124_4249_n405), .A2(
        n140), .A3(DP_OP_26J6_124_4249_n394), .Y(DP_OP_26J6_124_4249_n392) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U417 ( .A1(DP_OP_26J6_124_4249_n404), .A2(
        n140), .Y(DP_OP_26J6_124_4249_n391) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U414 ( .A1(ori_data_24_), .A2(n1280), .Y(
        DP_OP_26J6_124_4249_n389) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U413 ( .A1(n1260), .A2(ori_data_24_), .Y(
        DP_OP_26J6_124_4249_n388) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U408 ( .A1(DP_OP_26J6_124_4249_n405), .A2(
        DP_OP_26J6_124_4249_n386), .A3(DP_OP_26J6_124_4249_n387), .Y(
        DP_OP_26J6_124_4249_n381) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U407 ( .A1(DP_OP_26J6_124_4249_n404), .A2(
        DP_OP_26J6_124_4249_n386), .Y(DP_OP_26J6_124_4249_n380) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U400 ( .A1(ori_data_25_), .A2(n1260), .Y(
        DP_OP_26J6_124_4249_n378) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U399 ( .A1(n1290), .A2(ori_data_25_), .Y(
        DP_OP_26J6_124_4249_n377) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U389 ( .A1(DP_OP_26J6_124_4249_n382), .A2(
        DP_OP_26J6_124_4249_n570), .Y(DP_OP_26J6_124_4249_n369) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U386 ( .A1(ori_data_26_), .A2(n1270), .Y(
        DP_OP_26J6_124_4249_n367) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U385 ( .A1(n1270), .A2(ori_data_26_), .Y(
        DP_OP_26J6_124_4249_n366) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U381 ( .A1(DP_OP_26J6_124_4249_n366), .A2(
        DP_OP_26J6_124_4249_n377), .Y(DP_OP_26J6_124_4249_n360) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U376 ( .A1(DP_OP_26J6_124_4249_n383), .A2(
        DP_OP_26J6_124_4249_n360), .A3(DP_OP_26J6_124_4249_n361), .Y(
        DP_OP_26J6_124_4249_n359) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U375 ( .A1(DP_OP_26J6_124_4249_n382), .A2(
        DP_OP_26J6_124_4249_n360), .Y(DP_OP_26J6_124_4249_n358) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U372 ( .A1(ori_data_27_), .A2(n1270), .Y(
        DP_OP_26J6_124_4249_n356) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U361 ( .A1(DP_OP_26J6_124_4249_n349), .A2(
        DP_OP_26J6_124_4249_n382), .Y(DP_OP_26J6_124_4249_n347) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U358 ( .A1(ori_data_28_), .A2(n1260), .Y(
        DP_OP_26J6_124_4249_n345) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U353 ( .A1(DP_OP_26J6_124_4249_n344), .A2(
        DP_OP_26J6_124_4249_n351), .Y(DP_OP_26J6_124_4249_n342) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U352 ( .A1(DP_OP_26J6_124_4249_n361), .A2(
        DP_OP_26J6_124_4249_n342), .A3(DP_OP_26J6_124_4249_n343), .Y(
        DP_OP_26J6_124_4249_n341) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U351 ( .A1(DP_OP_26J6_124_4249_n360), .A2(
        DP_OP_26J6_124_4249_n342), .Y(DP_OP_26J6_124_4249_n340) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U349 ( .A1(DP_OP_26J6_124_4249_n340), .A2(
        DP_OP_26J6_124_4249_n380), .Y(DP_OP_26J6_124_4249_n338) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U344 ( .A1(ori_data_29_), .A2(n1290), .Y(
        DP_OP_26J6_124_4249_n334) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U338 ( .A1(DP_OP_26J6_124_4249_n339), .A2(
        n139), .A3(DP_OP_26J6_124_4249_n332), .Y(DP_OP_26J6_124_4249_n330) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U337 ( .A1(DP_OP_26J6_124_4249_n338), .A2(
        n139), .Y(DP_OP_26J6_124_4249_n329) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U312 ( .A1(ori_data_6_), .A2(ori_data_5_), 
        .Y(DP_OP_26J6_124_4249_n263) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U307 ( .A1(DP_OP_26J6_124_4249_n262), .A2(
        DP_OP_26J6_124_4249_n263), .Y(DP_OP_26J6_124_4249_n261) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U304 ( .A1(ori_data_8_), .A2(bias_data[0]), 
        .Y(DP_OP_26J6_124_4249_n259) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U294 ( .A1(ori_data_9_), .A2(bias_data[1]), 
        .Y(DP_OP_26J6_124_4249_n252) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U289 ( .A1(DP_OP_26J6_124_4249_n251), .A2(
        DP_OP_26J6_124_4249_n258), .Y(DP_OP_26J6_124_4249_n249) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U288 ( .A1(DP_OP_26J6_124_4249_n249), .A2(
        DP_OP_26J6_124_4249_n261), .A3(DP_OP_26J6_124_4249_n250), .Y(
        DP_OP_26J6_124_4249_n248) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U285 ( .A1(ori_data_10_), .A2(bias_data[2]), 
        .Y(DP_OP_26J6_124_4249_n246) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U275 ( .A1(DP_OP_26J6_124_4249_n247), .A2(
        DP_OP_26J6_124_4249_n289), .A3(DP_OP_26J6_124_4249_n240), .Y(
        DP_OP_26J6_124_4249_n238) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U273 ( .A1(ori_data_11_), .A2(n1250), .Y(
        DP_OP_26J6_124_4249_n237) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U272 ( .A1(n1240), .A2(ori_data_11_), .Y(
        DP_OP_26J6_124_4249_n236) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U270 ( .A1(DP_OP_26J6_124_4249_n584), .A2(
        DP_OP_26J6_124_4249_n237), .Y(DP_OP_26J6_124_4249_n24) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U268 ( .A1(DP_OP_26J6_124_4249_n236), .A2(
        DP_OP_26J6_124_4249_n245), .Y(DP_OP_26J6_124_4249_n230) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U261 ( .A1(ori_data_12_), .A2(n1240), .Y(
        DP_OP_26J6_124_4249_n228) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U260 ( .A1(n1280), .A2(ori_data_12_), .Y(
        DP_OP_26J6_124_4249_n223) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U249 ( .A1(ori_data_13_), .A2(n1240), .Y(
        DP_OP_26J6_124_4249_n219) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U244 ( .A1(DP_OP_26J6_124_4249_n218), .A2(
        DP_OP_26J6_124_4249_n223), .Y(DP_OP_26J6_124_4249_n216) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U243 ( .A1(DP_OP_26J6_124_4249_n231), .A2(
        DP_OP_26J6_124_4249_n216), .A3(DP_OP_26J6_124_4249_n217), .Y(
        DP_OP_26J6_124_4249_n215) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U242 ( .A1(DP_OP_26J6_124_4249_n230), .A2(
        DP_OP_26J6_124_4249_n216), .Y(DP_OP_26J6_124_4249_n214) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U238 ( .A1(ori_data_14_), .A2(n1240), .Y(
        DP_OP_26J6_124_4249_n211) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U224 ( .A1(ori_data_15_), .A2(bias_data[3]), 
        .Y(DP_OP_26J6_124_4249_n200) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U223 ( .A1(n1250), .A2(ori_data_15_), .Y(
        DP_OP_26J6_124_4249_n199) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U219 ( .A1(DP_OP_26J6_124_4249_n199), .A2(
        DP_OP_26J6_124_4249_n210), .Y(DP_OP_26J6_124_4249_n193) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U210 ( .A1(ori_data_16_), .A2(bias_data[3]), 
        .Y(DP_OP_26J6_124_4249_n189) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U209 ( .A1(n1240), .A2(ori_data_16_), .Y(
        DP_OP_26J6_124_4249_n188) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U199 ( .A1(DP_OP_26J6_124_4249_n193), .A2(
        DP_OP_26J6_124_4249_n283), .Y(DP_OP_26J6_124_4249_n180) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U196 ( .A1(ori_data_17_), .A2(n1250), .Y(
        DP_OP_26J6_124_4249_n178) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U195 ( .A1(n1260), .A2(ori_data_17_), .Y(
        DP_OP_26J6_124_4249_n177) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U191 ( .A1(DP_OP_26J6_124_4249_n177), .A2(
        DP_OP_26J6_124_4249_n188), .Y(DP_OP_26J6_124_4249_n175) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U190 ( .A1(DP_OP_26J6_124_4249_n194), .A2(
        DP_OP_26J6_124_4249_n175), .A3(DP_OP_26J6_124_4249_n176), .Y(
        DP_OP_26J6_124_4249_n170) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U189 ( .A1(DP_OP_26J6_124_4249_n193), .A2(
        DP_OP_26J6_124_4249_n175), .Y(DP_OP_26J6_124_4249_n169) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U182 ( .A1(ori_data_18_), .A2(n1250), .Y(
        DP_OP_26J6_124_4249_n167) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U181 ( .A1(bias_data[3]), .A2(ori_data_18_), 
        .Y(DP_OP_26J6_124_4249_n166) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U168 ( .A1(ori_data_19_), .A2(bias_data[3]), 
        .Y(DP_OP_26J6_124_4249_n156) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U167 ( .A1(n1240), .A2(ori_data_19_), .Y(
        DP_OP_26J6_124_4249_n155) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U163 ( .A1(DP_OP_26J6_124_4249_n155), .A2(
        DP_OP_26J6_124_4249_n166), .Y(DP_OP_26J6_124_4249_n149) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U158 ( .A1(DP_OP_26J6_124_4249_n172), .A2(
        DP_OP_26J6_124_4249_n149), .A3(DP_OP_26J6_124_4249_n150), .Y(
        DP_OP_26J6_124_4249_n148) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U157 ( .A1(DP_OP_26J6_124_4249_n171), .A2(
        DP_OP_26J6_124_4249_n149), .Y(DP_OP_26J6_124_4249_n147) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U154 ( .A1(ori_data_20_), .A2(n1250), .Y(
        DP_OP_26J6_124_4249_n145) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U153 ( .A1(bias_data[3]), .A2(ori_data_20_), 
        .Y(DP_OP_26J6_124_4249_n140) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U140 ( .A1(ori_data_21_), .A2(n1250), .Y(
        DP_OP_26J6_124_4249_n134) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U139 ( .A1(n1250), .A2(ori_data_21_), .Y(
        DP_OP_26J6_124_4249_n133) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U135 ( .A1(DP_OP_26J6_124_4249_n133), .A2(
        DP_OP_26J6_124_4249_n140), .Y(DP_OP_26J6_124_4249_n131) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U134 ( .A1(DP_OP_26J6_124_4249_n150), .A2(
        DP_OP_26J6_124_4249_n131), .A3(DP_OP_26J6_124_4249_n132), .Y(
        DP_OP_26J6_124_4249_n130) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U133 ( .A1(DP_OP_26J6_124_4249_n149), .A2(
        DP_OP_26J6_124_4249_n131), .Y(DP_OP_26J6_124_4249_n129) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U131 ( .A1(DP_OP_26J6_124_4249_n129), .A2(
        DP_OP_26J6_124_4249_n169), .Y(DP_OP_26J6_124_4249_n127) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U128 ( .A1(ori_data_22_), .A2(n1250), .Y(
        DP_OP_26J6_124_4249_n117) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U108 ( .A1(n140), .A2(
        DP_OP_26J6_124_4249_n123), .A3(DP_OP_26J6_124_4249_n394), .Y(
        DP_OP_26J6_124_4249_n106) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U100 ( .A1(ori_data_24_), .A2(n1250), .Y(
        DP_OP_26J6_124_4249_n103) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U99 ( .A1(n1240), .A2(ori_data_24_), .Y(
        DP_OP_26J6_124_4249_n102) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U86 ( .A1(ori_data_25_), .A2(bias_data[3]), 
        .Y(DP_OP_26J6_124_4249_n92) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U85 ( .A1(n1290), .A2(ori_data_25_), .Y(
        DP_OP_26J6_124_4249_n91) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U77 ( .A1(DP_OP_26J6_124_4249_n105), .A2(n141), .Y(DP_OP_26J6_124_4249_n3) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U72 ( .A1(ori_data_26_), .A2(n1240), .Y(
        DP_OP_26J6_124_4249_n81) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U71 ( .A1(bias_data[3]), .A2(ori_data_26_), 
        .Y(DP_OP_26J6_124_4249_n80) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U61 ( .A1(DP_OP_26J6_124_4249_n3), .A2(
        DP_OP_26J6_124_4249_n74), .Y(DP_OP_26J6_124_4249_n72) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U58 ( .A1(ori_data_27_), .A2(n1240), .Y(
        DP_OP_26J6_124_4249_n70) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U57 ( .A1(bias_data[3]), .A2(ori_data_27_), 
        .Y(DP_OP_26J6_124_4249_n69) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U55 ( .A1(DP_OP_26J6_124_4249_n272), .A2(
        DP_OP_26J6_124_4249_n70), .Y(DP_OP_26J6_124_4249_n8) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U53 ( .A1(DP_OP_26J6_124_4249_n69), .A2(
        DP_OP_26J6_124_4249_n80), .Y(DP_OP_26J6_124_4249_n63) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U48 ( .A1(DP_OP_26J6_124_4249_n2), .A2(
        DP_OP_26J6_124_4249_n63), .A3(DP_OP_26J6_124_4249_n64), .Y(
        DP_OP_26J6_124_4249_n62) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U47 ( .A1(DP_OP_26J6_124_4249_n3), .A2(
        DP_OP_26J6_124_4249_n63), .Y(DP_OP_26J6_124_4249_n61) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U44 ( .A1(ori_data_28_), .A2(n1240), .Y(
        DP_OP_26J6_124_4249_n59) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U43 ( .A1(n1290), .A2(ori_data_28_), .Y(
        DP_OP_26J6_124_4249_n54) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U41 ( .A1(DP_OP_26J6_124_4249_n271), .A2(
        DP_OP_26J6_124_4249_n59), .Y(DP_OP_26J6_124_4249_n7) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U30 ( .A1(ori_data_29_), .A2(n1250), .Y(
        DP_OP_26J6_124_4249_n48) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U25 ( .A1(DP_OP_26J6_124_4249_n47), .A2(
        DP_OP_26J6_124_4249_n54), .Y(DP_OP_26J6_124_4249_n45) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U20 ( .A1(DP_OP_26J6_124_4249_n2), .A2(n142), 
        .A3(n134), .Y(DP_OP_26J6_124_4249_n40) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U19 ( .A1(DP_OP_26J6_124_4249_n3), .A2(n142), 
        .Y(DP_OP_26J6_124_4249_n39) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U16 ( .A1(ori_data_30_), .A2(n1270), .Y(
        DP_OP_26J6_124_4249_n37) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U10 ( .A1(DP_OP_26J6_124_4249_n38), .A2(n135), .A3(DP_OP_26J6_124_4249_n35), .Y(DP_OP_26J6_124_4249_n33) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U8 ( .A1(ori_data_31_), .A2(n1250), .Y(
        DP_OP_26J6_124_4249_n32) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U5 ( .A1(n132), .A2(DP_OP_26J6_124_4249_n32), 
        .Y(DP_OP_26J6_124_4249_n4) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U614 ( .A1(n1270), .A2(ori_data_9_), .Y(
        DP_OP_26J6_124_4249_n544) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U293 ( .A1(bias_data[1]), .A2(ori_data_9_), 
        .Y(DP_OP_26J6_124_4249_n251) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U565 ( .A1(n1280), .A2(ori_data_13_), .Y(
        DP_OP_26J6_124_4249_n507) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U303 ( .A1(bias_data[0]), .A2(ori_data_8_), 
        .Y(DP_OP_26J6_124_4249_n258) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U29 ( .A1(n1250), .A2(ori_data_29_), .Y(
        DP_OP_26J6_124_4249_n47) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U78 ( .A1(n141), .A2(
        DP_OP_26J6_124_4249_n106), .A3(n137), .Y(DP_OP_26J6_124_4249_n2) );
  XNOR2X1_HVT DP_OP_26J6_124_4249_U45 ( .A1(DP_OP_26J6_124_4249_n71), .A2(
        DP_OP_26J6_124_4249_n8), .Y(N127) );
  XOR2X1_HVT DP_OP_26J6_124_4249_U4 ( .A1(DP_OP_26J6_124_4249_n33), .A2(
        DP_OP_26J6_124_4249_n4), .Y(N131) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U623 ( .A1(n1280), .A2(ori_data_8_), .Y(
        DP_OP_26J6_124_4249_n550) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U248 ( .A1(n1240), .A2(ori_data_13_), .Y(
        DP_OP_26J6_124_4249_n218) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U237 ( .A1(n1240), .A2(ori_data_14_), .Y(
        DP_OP_26J6_124_4249_n210) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U441 ( .A1(n1290), .A2(ori_data_22_), .Y(
        DP_OP_26J6_124_4249_n410) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U127 ( .A1(n1240), .A2(ori_data_22_), .Y(
        DP_OP_26J6_124_4249_n116) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U357 ( .A1(n1290), .A2(ori_data_28_), .Y(
        DP_OP_26J6_124_4249_n344) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U371 ( .A1(n1290), .A2(ori_data_27_), .Y(
        DP_OP_26J6_124_4249_n351) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U459 ( .A1(DP_OP_26J6_124_4249_n426), .A2(
        DP_OP_26J6_124_4249_n466), .Y(DP_OP_26J6_124_4249_n424) );
  AO221X1_HVT U3 ( .A1(1'b1), .A2(n470), .A3(DP_OP_26J6_124_4249_n281), .A4(
        DP_OP_26J6_124_4249_n172), .A5(DP_OP_26J6_124_4249_n161), .Y(n490) );
  AO221X1_HVT U4 ( .A1(1'b1), .A2(n390), .A3(DP_OP_26J6_124_4249_n138), .A4(
        DP_OP_26J6_124_4249_n172), .A5(DP_OP_26J6_124_4249_n139), .Y(n410) );
  OA221X1_HVT U5 ( .A1(1'b0), .A2(DP_OP_26J6_124_4249_n228), .A3(
        DP_OP_26J6_124_4249_n223), .A4(DP_OP_26J6_124_4249_n233), .A5(n105), 
        .Y(n1070) );
  OA221X1_HVT U6 ( .A1(1'b0), .A2(DP_OP_26J6_124_4249_n442), .A3(
        DP_OP_26J6_124_4249_n437), .A4(n85), .A5(n86), .Y(
        DP_OP_26J6_124_4249_n434) );
  OA221X1_HVT U7 ( .A1(1'b0), .A2(DP_OP_26J6_124_4249_n356), .A3(
        DP_OP_26J6_124_4249_n351), .A4(n33), .A5(n34), .Y(
        DP_OP_26J6_124_4249_n348) );
  OA221X1_HVT U8 ( .A1(1'b0), .A2(DP_OP_26J6_124_4249_n59), .A3(
        DP_OP_26J6_124_4249_n54), .A4(n18), .A5(n19), .Y(
        DP_OP_26J6_124_4249_n51) );
  NOR2X0_HVT U9 ( .A1(bias_data[2]), .A2(ori_data_10_), .Y(
        DP_OP_26J6_124_4249_n245) );
  AOI21X1_HVT U10 ( .A1(DP_OP_26J6_124_4249_n510), .A2(
        DP_OP_26J6_124_4249_n424), .A3(DP_OP_26J6_124_4249_n425), .Y(
        DP_OP_26J6_124_4249_n294) );
  OAI21X1_HVT U11 ( .A1(DP_OP_26J6_124_4249_n426), .A2(
        DP_OP_26J6_124_4249_n467), .A3(DP_OP_26J6_124_4249_n427), .Y(
        DP_OP_26J6_124_4249_n425) );
  INVX1_HVT U12 ( .A(DP_OP_26J6_124_4249_n213), .Y(DP_OP_26J6_124_4249_n212)
         );
  OAI21X1_HVT U13 ( .A1(DP_OP_26J6_124_4249_n545), .A2(
        DP_OP_26J6_124_4249_n535), .A3(DP_OP_26J6_124_4249_n536), .Y(
        DP_OP_26J6_124_4249_n534) );
  XOR2X1_HVT U14 ( .A1(DP_OP_26J6_124_4249_n454), .A2(n138), .Y(N48) );
  OAI21X1_HVT U15 ( .A1(DP_OP_26J6_124_4249_n455), .A2(
        DP_OP_26J6_124_4249_n509), .A3(DP_OP_26J6_124_4249_n456), .Y(
        DP_OP_26J6_124_4249_n454) );
  OAI21X1_HVT U16 ( .A1(DP_OP_26J6_124_4249_n39), .A2(DP_OP_26J6_124_4249_n1), 
        .A3(DP_OP_26J6_124_4249_n40), .Y(DP_OP_26J6_124_4249_n38) );
  OAI21X1_HVT U17 ( .A1(DP_OP_26J6_124_4249_n246), .A2(
        DP_OP_26J6_124_4249_n236), .A3(DP_OP_26J6_124_4249_n237), .Y(
        DP_OP_26J6_124_4249_n231) );
  INVX1_HVT U18 ( .A(DP_OP_26J6_124_4249_n246), .Y(DP_OP_26J6_124_4249_n240)
         );
  OA21X1_HVT U19 ( .A1(DP_OP_26J6_124_4249_n509), .A2(DP_OP_26J6_124_4249_n488), .A3(DP_OP_26J6_124_4249_n489), .Y(n1) );
  NAND2X0_HVT U20 ( .A1(DP_OP_26J6_124_4249_n580), .A2(
        DP_OP_26J6_124_4249_n486), .Y(n2) );
  HADDX1_HVT U21 ( .A0(n1), .B0(n2), .SO(N45) );
  OA21X1_HVT U22 ( .A1(DP_OP_26J6_124_4249_n147), .A2(DP_OP_26J6_124_4249_n212), .A3(DP_OP_26J6_124_4249_n148), .Y(n3) );
  NAND2X0_HVT U23 ( .A1(DP_OP_26J6_124_4249_n279), .A2(
        DP_OP_26J6_124_4249_n145), .Y(n4) );
  HADDX1_HVT U24 ( .A0(n3), .B0(n4), .SO(N120) );
  INVX0_HVT U25 ( .A(DP_OP_26J6_124_4249_n509), .Y(n5) );
  NAND3X0_HVT U26 ( .A1(DP_OP_26J6_124_4249_n446), .A2(
        DP_OP_26J6_124_4249_n468), .A3(n5), .Y(n6) );
  AO22X1_HVT U27 ( .A1(DP_OP_26J6_124_4249_n442), .A2(DP_OP_26J6_124_4249_n576), .A3(DP_OP_26J6_124_4249_n445), .A4(n6), .Y(n7) );
  NAND4X0_HVT U28 ( .A1(DP_OP_26J6_124_4249_n442), .A2(
        DP_OP_26J6_124_4249_n576), .A3(DP_OP_26J6_124_4249_n445), .A4(n6), .Y(
        n9) );
  NAND2X0_HVT U29 ( .A1(n7), .A2(n9), .Y(N49) );
  OA21X1_HVT U30 ( .A1(DP_OP_26J6_124_4249_n210), .A2(DP_OP_26J6_124_4249_n212), .A3(DP_OP_26J6_124_4249_n211), .Y(n10) );
  NAND2X0_HVT U31 ( .A1(DP_OP_26J6_124_4249_n580), .A2(
        DP_OP_26J6_124_4249_n200), .Y(n11) );
  HADDX1_HVT U32 ( .A0(n10), .B0(n11), .SO(N115) );
  INVX0_HVT U33 ( .A(DP_OP_26J6_124_4249_n388), .Y(n12) );
  OA21X1_HVT U34 ( .A1(ori_data_23_), .A2(n1280), .A3(n12), .Y(
        DP_OP_26J6_124_4249_n386) );
  NAND2X0_HVT U35 ( .A1(DP_OP_26J6_124_4249_n574), .A2(
        DP_OP_26J6_124_4249_n422), .Y(n14) );
  HADDX1_HVT U36 ( .A0(DP_OP_26J6_124_4249_n294), .B0(n14), .SO(N51) );
  OA21X1_HVT U37 ( .A1(DP_OP_26J6_124_4249_n191), .A2(DP_OP_26J6_124_4249_n212), .A3(DP_OP_26J6_124_4249_n192), .Y(n15) );
  NAND2X0_HVT U38 ( .A1(DP_OP_26J6_124_4249_n283), .A2(
        DP_OP_26J6_124_4249_n189), .Y(n16) );
  HADDX1_HVT U39 ( .A0(n15), .B0(n16), .SO(N116) );
  INVX0_HVT U41 ( .A(DP_OP_26J6_124_4249_n64), .Y(n18) );
  NAND2X0_HVT U42 ( .A1(DP_OP_26J6_124_4249_n2), .A2(DP_OP_26J6_124_4249_n52), 
        .Y(n19) );
  OA21X1_HVT U43 ( .A1(DP_OP_26J6_124_4249_n507), .A2(DP_OP_26J6_124_4249_n509), .A3(DP_OP_26J6_124_4249_n508), .Y(n20) );
  NAND2X0_HVT U44 ( .A1(DP_OP_26J6_124_4249_n285), .A2(
        DP_OP_26J6_124_4249_n497), .Y(n21) );
  HADDX1_HVT U45 ( .A0(n20), .B0(n21), .SO(N44) );
  NAND2X0_HVT U46 ( .A1(DP_OP_26J6_124_4249_n277), .A2(
        DP_OP_26J6_124_4249_n117), .Y(n22) );
  HADDX1_HVT U47 ( .A0(DP_OP_26J6_124_4249_n1), .B0(n22), .SO(N122) );
  OA21X1_HVT U48 ( .A1(DP_OP_26J6_124_4249_n402), .A2(DP_OP_26J6_124_4249_n294), .A3(DP_OP_26J6_124_4249_n403), .Y(n23) );
  NAND2X0_HVT U49 ( .A1(n140), .A2(DP_OP_26J6_124_4249_n400), .Y(n24) );
  HADDX1_HVT U50 ( .A0(n23), .B0(n24), .SO(N53) );
  NAND2X0_HVT U51 ( .A1(DP_OP_26J6_124_4249_n285), .A2(
        DP_OP_26J6_124_4249_n211), .Y(n25) );
  HADDX1_HVT U52 ( .A0(DP_OP_26J6_124_4249_n212), .B0(n25), .SO(N114) );
  OA21X1_HVT U53 ( .A1(DP_OP_26J6_124_4249_n294), .A2(DP_OP_26J6_124_4249_n336), .A3(DP_OP_26J6_124_4249_n337), .Y(n26) );
  NAND2X0_HVT U54 ( .A1(n139), .A2(DP_OP_26J6_124_4249_n334), .Y(n27) );
  HADDX1_HVT U55 ( .A0(n26), .B0(n27), .SO(N59) );
  OA21X1_HVT U56 ( .A1(DP_OP_26J6_124_4249_n180), .A2(DP_OP_26J6_124_4249_n212), .A3(DP_OP_26J6_124_4249_n181), .Y(n28) );
  NAND2X0_HVT U57 ( .A1(DP_OP_26J6_124_4249_n282), .A2(
        DP_OP_26J6_124_4249_n178), .Y(n29) );
  HADDX1_HVT U58 ( .A0(n28), .B0(n29), .SO(N117) );
  AND2X1_HVT U59 ( .A1(n135), .A2(DP_OP_26J6_124_4249_n37), .Y(n30) );
  HADDX1_HVT U60 ( .A0(n30), .B0(DP_OP_26J6_124_4249_n38), .SO(N130) );
  NAND2X0_HVT U61 ( .A1(DP_OP_26J6_124_4249_n469), .A2(
        DP_OP_26J6_124_4249_n282), .Y(n31) );
  AND2X1_HVT U62 ( .A1(n31), .A2(DP_OP_26J6_124_4249_n464), .Y(
        DP_OP_26J6_124_4249_n456) );
  INVX0_HVT U64 ( .A(DP_OP_26J6_124_4249_n361), .Y(n33) );
  NAND2X0_HVT U65 ( .A1(DP_OP_26J6_124_4249_n383), .A2(
        DP_OP_26J6_124_4249_n349), .Y(n34) );
  NAND2X0_HVT U66 ( .A1(DP_OP_26J6_124_4249_n2), .A2(DP_OP_26J6_124_4249_n74), 
        .Y(n35) );
  AND2X1_HVT U67 ( .A1(n35), .A2(DP_OP_26J6_124_4249_n81), .Y(
        DP_OP_26J6_124_4249_n73) );
  OA21X1_HVT U68 ( .A1(DP_OP_26J6_124_4249_n391), .A2(DP_OP_26J6_124_4249_n294), .A3(DP_OP_26J6_124_4249_n392), .Y(n360) );
  NAND2X0_HVT U69 ( .A1(DP_OP_26J6_124_4249_n96), .A2(DP_OP_26J6_124_4249_n389), .Y(n370) );
  HADDX1_HVT U70 ( .A0(n360), .B0(n370), .SO(N54) );
  INVX0_HVT U71 ( .A(DP_OP_26J6_124_4249_n212), .Y(n380) );
  AND3X1_HVT U72 ( .A1(DP_OP_26J6_124_4249_n171), .A2(DP_OP_26J6_124_4249_n138), .A3(n380), .Y(n390) );
  AND2X1_HVT U74 ( .A1(DP_OP_26J6_124_4249_n574), .A2(DP_OP_26J6_124_4249_n134), .Y(n420) );
  HADDX1_HVT U75 ( .A0(n420), .B0(n410), .SO(N121) );
  OA21X1_HVT U76 ( .A1(DP_OP_26J6_124_4249_n294), .A2(DP_OP_26J6_124_4249_n347), .A3(DP_OP_26J6_124_4249_n348), .Y(n430) );
  NAND2X0_HVT U77 ( .A1(DP_OP_26J6_124_4249_n271), .A2(
        DP_OP_26J6_124_4249_n345), .Y(n440) );
  HADDX1_HVT U78 ( .A0(n430), .B0(n440), .SO(N58) );
  INVX0_HVT U79 ( .A(DP_OP_26J6_124_4249_n96), .Y(n450) );
  OA21X1_HVT U80 ( .A1(DP_OP_26J6_124_4249_n106), .A2(n450), .A3(
        DP_OP_26J6_124_4249_n103), .Y(DP_OP_26J6_124_4249_n95) );
  INVX0_HVT U81 ( .A(DP_OP_26J6_124_4249_n212), .Y(n460) );
  AND3X1_HVT U82 ( .A1(DP_OP_26J6_124_4249_n171), .A2(DP_OP_26J6_124_4249_n281), .A3(n460), .Y(n470) );
  AND2X1_HVT U84 ( .A1(DP_OP_26J6_124_4249_n576), .A2(DP_OP_26J6_124_4249_n156), .Y(n500) );
  HADDX1_HVT U85 ( .A0(n500), .B0(n490), .SO(N119) );
  INVX0_HVT U86 ( .A(DP_OP_26J6_124_4249_n437), .Y(n510) );
  AND2X1_HVT U87 ( .A1(DP_OP_26J6_124_4249_n446), .A2(n510), .Y(
        DP_OP_26J6_124_4249_n435) );
  OA21X1_HVT U88 ( .A1(DP_OP_26J6_124_4249_n294), .A2(DP_OP_26J6_124_4249_n369), .A3(DP_OP_26J6_124_4249_n370), .Y(n520) );
  NAND2X0_HVT U89 ( .A1(DP_OP_26J6_124_4249_n74), .A2(DP_OP_26J6_124_4249_n367), .Y(n530) );
  HADDX1_HVT U90 ( .A0(n520), .B0(n530), .SO(N56) );
  NAND2X0_HVT U91 ( .A1(DP_OP_26J6_124_4249_n52), .A2(DP_OP_26J6_124_4249_n3), 
        .Y(n540) );
  OA21X1_HVT U92 ( .A1(DP_OP_26J6_124_4249_n1), .A2(n540), .A3(
        DP_OP_26J6_124_4249_n51), .Y(n550) );
  NAND2X0_HVT U93 ( .A1(n139), .A2(DP_OP_26J6_124_4249_n48), .Y(n560) );
  HADDX1_HVT U94 ( .A0(n550), .B0(n560), .SO(N129) );
  INVX0_HVT U95 ( .A(DP_OP_26J6_124_4249_n351), .Y(n570) );
  AND2X1_HVT U96 ( .A1(DP_OP_26J6_124_4249_n360), .A2(n570), .Y(
        DP_OP_26J6_124_4249_n349) );
  OA21X1_HVT U97 ( .A1(DP_OP_26J6_124_4249_n421), .A2(DP_OP_26J6_124_4249_n294), .A3(DP_OP_26J6_124_4249_n422), .Y(n580) );
  NAND2X0_HVT U98 ( .A1(DP_OP_26J6_124_4249_n277), .A2(
        DP_OP_26J6_124_4249_n411), .Y(n590) );
  HADDX1_HVT U99 ( .A0(n580), .B0(n590), .SO(N52) );
  NAND2X0_HVT U100 ( .A1(DP_OP_26J6_124_4249_n491), .A2(
        DP_OP_26J6_124_4249_n580), .Y(n600) );
  AND2X1_HVT U101 ( .A1(n600), .A2(DP_OP_26J6_124_4249_n486), .Y(
        DP_OP_26J6_124_4249_n478) );
  NAND2X0_HVT U102 ( .A1(DP_OP_26J6_124_4249_n194), .A2(
        DP_OP_26J6_124_4249_n283), .Y(n610) );
  AND2X1_HVT U103 ( .A1(n610), .A2(DP_OP_26J6_124_4249_n189), .Y(
        DP_OP_26J6_124_4249_n181) );
  NAND2X0_HVT U104 ( .A1(n1290), .A2(ori_data_31_), .Y(n62) );
  AND2X1_HVT U105 ( .A1(n62), .A2(n133), .Y(n63) );
  AO21X1_HVT U106 ( .A1(n136), .A2(DP_OP_26J6_124_4249_n328), .A3(
        DP_OP_26J6_124_4249_n35), .Y(n64) );
  HADDX1_HVT U107 ( .A0(n63), .B0(n64), .SO(N61) );
  OA21X1_HVT U108 ( .A1(DP_OP_26J6_124_4249_n1), .A2(DP_OP_26J6_124_4249_n105), 
        .A3(DP_OP_26J6_124_4249_n106), .Y(n65) );
  NAND2X0_HVT U109 ( .A1(DP_OP_26J6_124_4249_n96), .A2(
        DP_OP_26J6_124_4249_n103), .Y(n66) );
  HADDX1_HVT U110 ( .A0(n65), .B0(n66), .SO(N124) );
  NAND2X0_HVT U111 ( .A1(DP_OP_26J6_124_4249_n64), .A2(DP_OP_26J6_124_4249_n45), .Y(n67) );
  OR2X1_HVT U112 ( .A1(DP_OP_26J6_124_4249_n47), .A2(DP_OP_26J6_124_4249_n59), 
        .Y(n68) );
  NAND3X0_HVT U113 ( .A1(n68), .A2(DP_OP_26J6_124_4249_n48), .A3(n67), .Y(n134) );
  NAND2X0_HVT U114 ( .A1(n1260), .A2(ori_data_30_), .Y(n69) );
  AND2X1_HVT U115 ( .A1(n136), .A2(n69), .Y(n70) );
  HADDX1_HVT U116 ( .A0(n70), .B0(DP_OP_26J6_124_4249_n328), .SO(N60) );
  NAND2X0_HVT U117 ( .A1(DP_OP_26J6_124_4249_n96), .A2(
        DP_OP_26J6_124_4249_n107), .Y(n71) );
  OA21X1_HVT U118 ( .A1(DP_OP_26J6_124_4249_n1), .A2(n71), .A3(
        DP_OP_26J6_124_4249_n95), .Y(n72) );
  NAND2X0_HVT U119 ( .A1(DP_OP_26J6_124_4249_n92), .A2(
        DP_OP_26J6_124_4249_n570), .Y(n73) );
  HADDX1_HVT U120 ( .A0(n72), .B0(n73), .SO(N125) );
  OA21X1_HVT U121 ( .A1(DP_OP_26J6_124_4249_n557), .A2(
        DP_OP_26J6_124_4249_n559), .A3(DP_OP_26J6_124_4249_n558), .Y(n74) );
  INVX0_HVT U122 ( .A(DP_OP_26J6_124_4249_n550), .Y(n75) );
  NAND2X0_HVT U123 ( .A1(n75), .A2(DP_OP_26J6_124_4249_n551), .Y(n76) );
  HADDX1_HVT U124 ( .A0(n74), .B0(n76), .SO(N38) );
  INVX0_HVT U125 ( .A(DP_OP_26J6_124_4249_n452), .Y(n77) );
  OA21X1_HVT U126 ( .A1(ori_data_17_), .A2(n1260), .A3(n77), .Y(
        DP_OP_26J6_124_4249_n446) );
  NAND2X0_HVT U127 ( .A1(DP_OP_26J6_124_4249_n582), .A2(
        DP_OP_26J6_124_4249_n508), .Y(n78) );
  HADDX1_HVT U128 ( .A0(DP_OP_26J6_124_4249_n509), .B0(n78), .SO(N43) );
  OA21X1_HVT U129 ( .A1(DP_OP_26J6_124_4249_n1), .A2(DP_OP_26J6_124_4249_n116), 
        .A3(DP_OP_26J6_124_4249_n117), .Y(n79) );
  NAND2X0_HVT U130 ( .A1(ori_data_23_), .A2(bias_data[3]), .Y(n80) );
  NAND2X0_HVT U131 ( .A1(n80), .A2(n140), .Y(n81) );
  HADDX1_HVT U132 ( .A0(n79), .B0(n81), .SO(N123) );
  INVX0_HVT U133 ( .A(DP_OP_26J6_124_4249_n561), .Y(n82) );
  NAND2X0_HVT U134 ( .A1(n82), .A2(DP_OP_26J6_124_4249_n562), .Y(n83) );
  HADDX1_HVT U135 ( .A0(DP_OP_26J6_124_4249_n563), .B0(n83), .SO(N36) );
  AND2X1_HVT U136 ( .A1(DP_OP_26J6_124_4249_n586), .A2(
        DP_OP_26J6_124_4249_n545), .Y(n84) );
  HADDX1_HVT U137 ( .A0(n84), .B0(DP_OP_26J6_124_4249_n546), .SO(N39) );
  INVX0_HVT U138 ( .A(DP_OP_26J6_124_4249_n447), .Y(n85) );
  NAND2X0_HVT U139 ( .A1(DP_OP_26J6_124_4249_n469), .A2(
        DP_OP_26J6_124_4249_n435), .Y(n86) );
  INVX0_HVT U141 ( .A(DP_OP_26J6_124_4249_n140), .Y(n88) );
  AND2X1_HVT U142 ( .A1(DP_OP_26J6_124_4249_n149), .A2(n88), .Y(
        DP_OP_26J6_124_4249_n138) );
  OA21X1_HVT U143 ( .A1(DP_OP_26J6_124_4249_n380), .A2(
        DP_OP_26J6_124_4249_n294), .A3(DP_OP_26J6_124_4249_n381), .Y(n89) );
  NAND2X0_HVT U144 ( .A1(DP_OP_26J6_124_4249_n570), .A2(
        DP_OP_26J6_124_4249_n378), .Y(n90) );
  HADDX1_HVT U145 ( .A0(n89), .B0(n90), .SO(N55) );
  OA21X1_HVT U146 ( .A1(DP_OP_26J6_124_4249_n83), .A2(DP_OP_26J6_124_4249_n1), 
        .A3(DP_OP_26J6_124_4249_n84), .Y(n91) );
  NAND2X0_HVT U147 ( .A1(DP_OP_26J6_124_4249_n74), .A2(DP_OP_26J6_124_4249_n81), .Y(n92) );
  HADDX1_HVT U148 ( .A0(n91), .B0(n92), .SO(N126) );
  OR4X1_HVT U149 ( .A1(N128), .A2(N124), .A3(N125), .A4(N123), .Y(n162) );
  HADDX1_HVT U150 ( .A0(ori_data_5_), .B0(ori_data_6_), .SO(N106) );
  AND2X1_HVT U151 ( .A1(DP_OP_26J6_124_4249_n289), .A2(
        DP_OP_26J6_124_4249_n246), .Y(n93) );
  HADDX1_HVT U152 ( .A0(n93), .B0(DP_OP_26J6_124_4249_n247), .SO(N110) );
  OA21X1_HVT U153 ( .A1(DP_OP_26J6_124_4249_n526), .A2(
        DP_OP_26J6_124_4249_n528), .A3(DP_OP_26J6_124_4249_n527), .Y(n94) );
  NAND2X0_HVT U154 ( .A1(DP_OP_26J6_124_4249_n287), .A2(
        DP_OP_26J6_124_4249_n516), .Y(n95) );
  HADDX1_HVT U155 ( .A0(n94), .B0(n95), .SO(N42) );
  OA21X1_HVT U156 ( .A1(DP_OP_26J6_124_4249_n358), .A2(
        DP_OP_26J6_124_4249_n294), .A3(DP_OP_26J6_124_4249_n359), .Y(n96) );
  NAND2X0_HVT U157 ( .A1(DP_OP_26J6_124_4249_n272), .A2(
        DP_OP_26J6_124_4249_n356), .Y(n97) );
  HADDX1_HVT U158 ( .A0(n96), .B0(n97), .SO(N57) );
  INVX0_HVT U159 ( .A(DP_OP_26J6_124_4249_n258), .Y(n98) );
  NAND2X0_HVT U160 ( .A1(n98), .A2(DP_OP_26J6_124_4249_n259), .Y(n99) );
  HADDX1_HVT U161 ( .A0(DP_OP_26J6_124_4249_n260), .B0(n99), .SO(N108) );
  INVX0_HVT U162 ( .A(DP_OP_26J6_124_4249_n535), .Y(n100) );
  NAND2X0_HVT U163 ( .A1(DP_OP_26J6_124_4249_n546), .A2(
        DP_OP_26J6_124_4249_n586), .Y(n101) );
  AO22X1_HVT U164 ( .A1(n100), .A2(DP_OP_26J6_124_4249_n536), .A3(
        DP_OP_26J6_124_4249_n545), .A4(n101), .Y(n102) );
  NAND4X0_HVT U165 ( .A1(n100), .A2(DP_OP_26J6_124_4249_n536), .A3(
        DP_OP_26J6_124_4249_n545), .A4(n101), .Y(n103) );
  NAND2X0_HVT U166 ( .A1(n102), .A2(n103), .Y(N40) );
  INVX0_HVT U167 ( .A(DP_OP_26J6_124_4249_n223), .Y(n104) );
  NAND3X0_HVT U168 ( .A1(DP_OP_26J6_124_4249_n230), .A2(
        DP_OP_26J6_124_4249_n247), .A3(n104), .Y(n105) );
  NAND2X0_HVT U170 ( .A1(DP_OP_26J6_124_4249_n582), .A2(
        DP_OP_26J6_124_4249_n219), .Y(n1080) );
  HADDX1_HVT U171 ( .A0(n1070), .B0(n1080), .SO(N113) );
  NAND2X0_HVT U172 ( .A1(DP_OP_26J6_124_4249_n383), .A2(
        DP_OP_26J6_124_4249_n570), .Y(n1090) );
  AND2X1_HVT U173 ( .A1(n1090), .A2(DP_OP_26J6_124_4249_n378), .Y(
        DP_OP_26J6_124_4249_n370) );
  INVX0_HVT U174 ( .A(DP_OP_26J6_124_4249_n54), .Y(n1100) );
  AND2X1_HVT U175 ( .A1(DP_OP_26J6_124_4249_n63), .A2(n1100), .Y(
        DP_OP_26J6_124_4249_n52) );
  OA21X1_HVT U176 ( .A1(DP_OP_26J6_124_4249_n169), .A2(
        DP_OP_26J6_124_4249_n212), .A3(DP_OP_26J6_124_4249_n170), .Y(n1110) );
  NAND2X0_HVT U177 ( .A1(DP_OP_26J6_124_4249_n281), .A2(
        DP_OP_26J6_124_4249_n167), .Y(n1120) );
  HADDX1_HVT U178 ( .A0(n1110), .B0(n1120), .SO(N118) );
  INVX0_HVT U179 ( .A(DP_OP_26J6_124_4249_n557), .Y(n1130) );
  NAND2X0_HVT U180 ( .A1(n1130), .A2(DP_OP_26J6_124_4249_n558), .Y(n1140) );
  HADDX1_HVT U181 ( .A0(DP_OP_26J6_124_4249_n559), .B0(n1140), .SO(N37) );
  OA21X1_HVT U182 ( .A1(DP_OP_26J6_124_4249_n258), .A2(
        DP_OP_26J6_124_4249_n260), .A3(DP_OP_26J6_124_4249_n259), .Y(n1150) );
  INVX0_HVT U183 ( .A(DP_OP_26J6_124_4249_n251), .Y(n1160) );
  NAND2X0_HVT U184 ( .A1(n1160), .A2(DP_OP_26J6_124_4249_n252), .Y(n1170) );
  HADDX1_HVT U185 ( .A0(n1150), .B0(n1170), .SO(N109) );
  NAND2X0_HVT U186 ( .A1(DP_OP_26J6_124_4249_n584), .A2(
        DP_OP_26J6_124_4249_n527), .Y(n1180) );
  HADDX1_HVT U187 ( .A0(DP_OP_26J6_124_4249_n528), .B0(n1180), .SO(N41) );
  AOI21X1_HVT U188 ( .A1(DP_OP_26J6_124_4249_n230), .A2(
        DP_OP_26J6_124_4249_n247), .A3(DP_OP_26J6_124_4249_n231), .Y(n1190) );
  NAND2X0_HVT U189 ( .A1(DP_OP_26J6_124_4249_n287), .A2(
        DP_OP_26J6_124_4249_n228), .Y(n1200) );
  HADDX1_HVT U190 ( .A0(n1190), .B0(n1200), .SO(N112) );
  INVX0_HVT U191 ( .A(N113), .Y(n1210) );
  AO21X1_HVT U192 ( .A1(n202), .A2(n1210), .A3(n201), .Y(n1220) );
  AO21X1_HVT U193 ( .A1(n200), .A2(n199), .A3(n198), .Y(n1230) );
  NAND2X0_HVT U194 ( .A1(n1230), .A2(n1220), .Y(n_quantized_data[7]) );
  NAND2X2_HVT U195 ( .A1(n198), .A2(n201), .Y(n195) );
  INVX0_HVT U196 ( .A(DP_OP_26J6_124_4249_n485), .Y(DP_OP_26J6_124_4249_n580)
         );
  INVX0_HVT U197 ( .A(N131), .Y(n165) );
  INVX0_HVT U198 ( .A(N119), .Y(n155) );
  INVX0_HVT U199 ( .A(N121), .Y(n154) );
  AND3X1_HVT U200 ( .A1(N44), .A2(N43), .A3(N51), .Y(n167) );
  XNOR2X1_HVT U201 ( .A1(DP_OP_26J6_124_4249_n432), .A2(
        DP_OP_26J6_124_4249_n306), .Y(N50) );
  INVX0_HVT U202 ( .A(DP_OP_26J6_124_4249_n3), .Y(DP_OP_26J6_124_4249_n83) );
  INVX0_HVT U203 ( .A(DP_OP_26J6_124_4249_n338), .Y(DP_OP_26J6_124_4249_n336)
         );
  AOI21X1_HVT U204 ( .A1(DP_OP_26J6_124_4249_n546), .A2(
        DP_OP_26J6_124_4249_n533), .A3(DP_OP_26J6_124_4249_n534), .Y(
        DP_OP_26J6_124_4249_n528) );
  INVX0_HVT U205 ( .A(DP_OP_26J6_124_4249_n2), .Y(DP_OP_26J6_124_4249_n84) );
  INVX0_HVT U206 ( .A(DP_OP_26J6_124_4249_n169), .Y(DP_OP_26J6_124_4249_n171)
         );
  INVX0_HVT U207 ( .A(DP_OP_26J6_124_4249_n466), .Y(DP_OP_26J6_124_4249_n468)
         );
  INVX0_HVT U208 ( .A(DP_OP_26J6_124_4249_n105), .Y(DP_OP_26J6_124_4249_n107)
         );
  INVX0_HVT U209 ( .A(DP_OP_26J6_124_4249_n380), .Y(DP_OP_26J6_124_4249_n382)
         );
  INVX0_HVT U210 ( .A(DP_OP_26J6_124_4249_n404), .Y(DP_OP_26J6_124_4249_n402)
         );
  INVX0_HVT U211 ( .A(DP_OP_26J6_124_4249_n177), .Y(DP_OP_26J6_124_4249_n282)
         );
  INVX0_HVT U212 ( .A(DP_OP_26J6_124_4249_n188), .Y(DP_OP_26J6_124_4249_n283)
         );
  INVX0_HVT U213 ( .A(DP_OP_26J6_124_4249_n37), .Y(DP_OP_26J6_124_4249_n35) );
  INVX0_HVT U214 ( .A(DP_OP_26J6_124_4249_n69), .Y(DP_OP_26J6_124_4249_n272)
         );
  INVX0_HVT U215 ( .A(DP_OP_26J6_124_4249_n140), .Y(DP_OP_26J6_124_4249_n279)
         );
  INVX0_HVT U216 ( .A(DP_OP_26J6_124_4249_n334), .Y(DP_OP_26J6_124_4249_n332)
         );
  INVX0_HVT U217 ( .A(DP_OP_26J6_124_4249_n437), .Y(DP_OP_26J6_124_4249_n576)
         );
  INVX0_HVT U218 ( .A(DP_OP_26J6_124_4249_n167), .Y(DP_OP_26J6_124_4249_n161)
         );
  INVX0_HVT U219 ( .A(DP_OP_26J6_124_4249_n421), .Y(DP_OP_26J6_124_4249_n574)
         );
  INVX0_HVT U220 ( .A(DP_OP_26J6_124_4249_n223), .Y(DP_OP_26J6_124_4249_n287)
         );
  INVX0_HVT U221 ( .A(DP_OP_26J6_124_4249_n117), .Y(DP_OP_26J6_124_4249_n123)
         );
  INVX0_HVT U222 ( .A(DP_OP_26J6_124_4249_n54), .Y(DP_OP_26J6_124_4249_n271)
         );
  INVX0_HVT U223 ( .A(DP_OP_26J6_124_4249_n400), .Y(DP_OP_26J6_124_4249_n394)
         );
  INVX0_HVT U224 ( .A(DP_OP_26J6_124_4249_n193), .Y(DP_OP_26J6_124_4249_n191)
         );
  INVX0_HVT U225 ( .A(DP_OP_26J6_124_4249_n194), .Y(DP_OP_26J6_124_4249_n192)
         );
  INVX0_HVT U226 ( .A(DP_OP_26J6_124_4249_n491), .Y(DP_OP_26J6_124_4249_n489)
         );
  INVX0_HVT U227 ( .A(DP_OP_26J6_124_4249_n490), .Y(DP_OP_26J6_124_4249_n488)
         );
  INVX0_HVT U228 ( .A(DP_OP_26J6_124_4249_n507), .Y(DP_OP_26J6_124_4249_n582)
         );
  INVX0_HVT U229 ( .A(DP_OP_26J6_124_4249_n210), .Y(DP_OP_26J6_124_4249_n285)
         );
  INVX0_HVT U230 ( .A(DP_OP_26J6_124_4249_n526), .Y(DP_OP_26J6_124_4249_n584)
         );
  INVX1_HVT U231 ( .A(n1300), .Y(n1290) );
  INVX1_HVT U232 ( .A(n1300), .Y(n1240) );
  INVX1_HVT U233 ( .A(n1300), .Y(n1250) );
  INVX1_HVT U234 ( .A(n1300), .Y(n1260) );
  INVX1_HVT U235 ( .A(n1300), .Y(n1280) );
  INVX1_HVT U236 ( .A(n1300), .Y(n1270) );
  INVX0_HVT U237 ( .A(n180), .Y(n173) );
  INVX1_HVT U238 ( .A(bias_data[3]), .Y(n1300) );
  INVX0_HVT U239 ( .A(srstn), .Y(n13) );
  INVX1_HVT U240 ( .A(DP_OP_26J6_124_4249_n116), .Y(DP_OP_26J6_124_4249_n277)
         );
  INVX1_HVT U241 ( .A(DP_OP_26J6_124_4249_n150), .Y(DP_OP_26J6_124_4249_n152)
         );
  INVX1_HVT U242 ( .A(DP_OP_26J6_124_4249_n166), .Y(DP_OP_26J6_124_4249_n281)
         );
  INVX1_HVT U243 ( .A(DP_OP_26J6_124_4249_n170), .Y(DP_OP_26J6_124_4249_n172)
         );
  INVX1_HVT U244 ( .A(DP_OP_26J6_124_4249_n245), .Y(DP_OP_26J6_124_4249_n289)
         );
  INVX1_HVT U245 ( .A(DP_OP_26J6_124_4249_n261), .Y(DP_OP_26J6_124_4249_n260)
         );
  INVX1_HVT U246 ( .A(ori_data_7_), .Y(DP_OP_26J6_124_4249_n262) );
  INVX1_HVT U247 ( .A(DP_OP_26J6_124_4249_n80), .Y(DP_OP_26J6_124_4249_n74) );
  INVX1_HVT U248 ( .A(DP_OP_26J6_124_4249_n102), .Y(DP_OP_26J6_124_4249_n96)
         );
  INVX1_HVT U249 ( .A(DP_OP_26J6_124_4249_n339), .Y(DP_OP_26J6_124_4249_n337)
         );
  INVX1_HVT U250 ( .A(DP_OP_26J6_124_4249_n377), .Y(DP_OP_26J6_124_4249_n570)
         );
  INVX1_HVT U251 ( .A(DP_OP_26J6_124_4249_n381), .Y(DP_OP_26J6_124_4249_n383)
         );
  INVX1_HVT U252 ( .A(DP_OP_26J6_124_4249_n405), .Y(DP_OP_26J6_124_4249_n403)
         );
  INVX1_HVT U253 ( .A(DP_OP_26J6_124_4249_n467), .Y(DP_OP_26J6_124_4249_n469)
         );
  INVX1_HVT U254 ( .A(DP_OP_26J6_124_4249_n544), .Y(DP_OP_26J6_124_4249_n586)
         );
  OAI21X1_HVT U255 ( .A1(DP_OP_26J6_124_4249_n61), .A2(DP_OP_26J6_124_4249_n1), 
        .A3(DP_OP_26J6_124_4249_n62), .Y(DP_OP_26J6_124_4249_n60) );
  OAI21X1_HVT U256 ( .A1(DP_OP_26J6_124_4249_n72), .A2(DP_OP_26J6_124_4249_n1), 
        .A3(DP_OP_26J6_124_4249_n73), .Y(DP_OP_26J6_124_4249_n71) );
  OAI21X1_HVT U257 ( .A1(DP_OP_26J6_124_4249_n477), .A2(
        DP_OP_26J6_124_4249_n509), .A3(DP_OP_26J6_124_4249_n478), .Y(
        DP_OP_26J6_124_4249_n476) );
  OR2X1_HVT U258 ( .A1(n1240), .A2(ori_data_31_), .Y(n132) );
  OR2X1_HVT U259 ( .A1(n1280), .A2(ori_data_31_), .Y(n133) );
  OR2X1_HVT U260 ( .A1(bias_data[3]), .A2(ori_data_30_), .Y(n135) );
  OR2X1_HVT U261 ( .A1(n1270), .A2(ori_data_30_), .Y(n136) );
  OA21X1_HVT U262 ( .A1(DP_OP_26J6_124_4249_n103), .A2(DP_OP_26J6_124_4249_n91), .A3(DP_OP_26J6_124_4249_n92), .Y(n137) );
  AND2X1_HVT U263 ( .A1(DP_OP_26J6_124_4249_n281), .A2(
        DP_OP_26J6_124_4249_n453), .Y(n138) );
  OR2X1_HVT U264 ( .A1(n1280), .A2(ori_data_29_), .Y(n139) );
  OR2X1_HVT U265 ( .A1(n1250), .A2(ori_data_23_), .Y(n140) );
  OR2X1_HVT U266 ( .A1(DP_OP_26J6_124_4249_n91), .A2(DP_OP_26J6_124_4249_n102), 
        .Y(n141) );
  AND2X1_HVT U267 ( .A1(DP_OP_26J6_124_4249_n63), .A2(DP_OP_26J6_124_4249_n45), 
        .Y(n142) );
  NAND2X0_HVT U268 ( .A1(DP_OP_26J6_124_4249_n277), .A2(n140), .Y(
        DP_OP_26J6_124_4249_n105) );
  INVX1_HVT U269 ( .A(DP_OP_26J6_124_4249_n231), .Y(DP_OP_26J6_124_4249_n233)
         );
  NOR2X0_HVT U270 ( .A1(n1270), .A2(ori_data_11_), .Y(DP_OP_26J6_124_4249_n526) );
  OA21X1_HVT U271 ( .A1(DP_OP_26J6_124_4249_n466), .A2(
        DP_OP_26J6_124_4249_n509), .A3(DP_OP_26J6_124_4249_n467), .Y(n1310) );
  XOR2X1_HVT U272 ( .A1(n1310), .A2(DP_OP_26J6_124_4249_n309), .Y(N47) );
  INVX1_HVT U273 ( .A(DP_OP_26J6_124_4249_n547), .Y(DP_OP_26J6_124_4249_n546)
         );
  INVX1_HVT U274 ( .A(DP_OP_26J6_124_4249_n560), .Y(DP_OP_26J6_124_4249_n559)
         );
  AOI21X2_HVT U275 ( .A1(DP_OP_26J6_124_4249_n213), .A2(
        DP_OP_26J6_124_4249_n127), .A3(DP_OP_26J6_124_4249_n128), .Y(
        DP_OP_26J6_124_4249_n1) );
  INVX1_HVT U276 ( .A(DP_OP_26J6_124_4249_n248), .Y(DP_OP_26J6_124_4249_n247)
         );
  INVX4_HVT U277 ( .A(DP_OP_26J6_124_4249_n510), .Y(DP_OP_26J6_124_4249_n509)
         );
  OAI21X2_HVT U278 ( .A1(DP_OP_26J6_124_4249_n563), .A2(
        DP_OP_26J6_124_4249_n561), .A3(DP_OP_26J6_124_4249_n562), .Y(
        DP_OP_26J6_124_4249_n560) );
  NOR2X0_HVT U279 ( .A1(bias_data[0]), .A2(ori_data_5_), .Y(
        DP_OP_26J6_124_4249_n563) );
  OAI21X2_HVT U280 ( .A1(DP_OP_26J6_124_4249_n329), .A2(
        DP_OP_26J6_124_4249_n294), .A3(DP_OP_26J6_124_4249_n330), .Y(
        DP_OP_26J6_124_4249_n328) );
  AND2X1_HVT U281 ( .A1(N49), .A2(N50), .Y(n143) );
  AND3X1_HVT U282 ( .A1(n143), .A2(n168), .A3(n167), .Y(n169) );
  INVX1_HVT U283 ( .A(mode[0]), .Y(n151) );
  INVX1_HVT U284 ( .A(N43), .Y(n200) );
  INVX1_HVT U285 ( .A(N129), .Y(n158) );
  INVX1_HVT U286 ( .A(N126), .Y(n159) );
  INVX1_HVT U287 ( .A(N127), .Y(n160) );
  INVX1_HVT U288 ( .A(N130), .Y(n157) );
  OR3X1_HVT U289 ( .A1(N45), .A2(N46), .A3(n144), .Y(n145) );
  OR2X1_HVT U290 ( .A1(N47), .A2(N48), .Y(n144) );
  INVX1_HVT U291 ( .A(N61), .Y(n153) );
  INVX1_HVT U292 ( .A(n195), .Y(n196) );
  NOR4X1_HVT U293 ( .A1(N52), .A2(N53), .A3(N54), .A4(N55), .Y(n150) );
  NOR4X1_HVT U294 ( .A1(N58), .A2(N56), .A3(N59), .A4(N57), .Y(n149) );
  OR2X1_HVT U295 ( .A1(N49), .A2(N50), .Y(n147) );
  OR3X1_HVT U296 ( .A1(N43), .A2(N51), .A3(N44), .Y(n146) );
  NOR4X1_HVT U297 ( .A1(n147), .A2(N60), .A3(n146), .A4(n145), .Y(n148) );
  NAND3X0_HVT U298 ( .A1(n150), .A2(n149), .A3(n148), .Y(n152) );
  NAND2X0_HVT U299 ( .A1(n151), .A2(mode[1]), .Y(n180) );
  AO21X1_HVT U300 ( .A1(n153), .A2(n152), .A3(n180), .Y(n198) );
  NOR4X1_HVT U301 ( .A1(N114), .A2(N122), .A3(N113), .A4(N116), .Y(n156) );
  NAND4X0_HVT U302 ( .A1(n157), .A2(n156), .A3(n155), .A4(n154), .Y(n164) );
  NOR4X1_HVT U303 ( .A1(N115), .A2(N118), .A3(N117), .A4(N120), .Y(n161) );
  NAND4X0_HVT U304 ( .A1(n161), .A2(n160), .A3(n159), .A4(n158), .Y(n163) );
  OR3X1_HVT U305 ( .A1(n164), .A2(n163), .A3(n162), .Y(n166) );
  AO21X1_HVT U306 ( .A1(n166), .A2(n165), .A3(n173), .Y(n201) );
  AND4X1_HVT U307 ( .A1(N52), .A2(N53), .A3(N54), .A4(N55), .Y(n171) );
  AND4X1_HVT U308 ( .A1(N57), .A2(N56), .A3(N58), .A4(N59), .Y(n170) );
  AND4X1_HVT U309 ( .A1(N46), .A2(N45), .A3(N48), .A4(N47), .Y(n168) );
  NAND4X0_HVT U310 ( .A1(n171), .A2(n170), .A3(N60), .A4(n169), .Y(n172) );
  NAND2X0_HVT U311 ( .A1(N61), .A2(n172), .Y(n199) );
  AND2X1_HVT U312 ( .A1(n199), .A2(n173), .Y(n193) );
  NAND2X0_HVT U313 ( .A1(n193), .A2(N36), .Y(n182) );
  AND4X1_HVT U314 ( .A1(N116), .A2(N114), .A3(N122), .A4(N113), .Y(n174) );
  NAND4X0_HVT U315 ( .A1(N130), .A2(n174), .A3(N119), .A4(N121), .Y(n178) );
  NAND4X0_HVT U316 ( .A1(N128), .A2(N123), .A3(N125), .A4(N124), .Y(n177) );
  AND4X1_HVT U317 ( .A1(N115), .A2(N118), .A3(N117), .A4(N120), .Y(n175) );
  NAND4X0_HVT U318 ( .A1(N127), .A2(n175), .A3(N126), .A4(N129), .Y(n176) );
  OR3X1_HVT U319 ( .A1(n178), .A2(n177), .A3(n176), .Y(n179) );
  NAND2X0_HVT U320 ( .A1(n179), .A2(N131), .Y(n202) );
  AND2X1_HVT U321 ( .A1(n202), .A2(n180), .Y(n194) );
  NAND2X0_HVT U322 ( .A1(n194), .A2(N106), .Y(n181) );
  NAND3X0_HVT U323 ( .A1(n195), .A2(n182), .A3(n181), .Y(n_quantized_data[0])
         );
  NAND2X0_HVT U324 ( .A1(n193), .A2(N37), .Y(n184) );
  NAND2X0_HVT U325 ( .A1(n194), .A2(N107), .Y(n183) );
  NAND3X0_HVT U326 ( .A1(n195), .A2(n184), .A3(n183), .Y(n_quantized_data[1])
         );
  NAND2X0_HVT U327 ( .A1(n193), .A2(N38), .Y(n186) );
  NAND2X0_HVT U328 ( .A1(n194), .A2(N108), .Y(n185) );
  NAND3X0_HVT U329 ( .A1(n195), .A2(n186), .A3(n185), .Y(n_quantized_data[2])
         );
  NAND2X0_HVT U330 ( .A1(n193), .A2(N39), .Y(n188) );
  NAND2X0_HVT U331 ( .A1(n194), .A2(N109), .Y(n187) );
  NAND3X0_HVT U332 ( .A1(n195), .A2(n188), .A3(n187), .Y(n_quantized_data[3])
         );
  NAND2X0_HVT U333 ( .A1(n193), .A2(N40), .Y(n190) );
  NAND2X0_HVT U334 ( .A1(n194), .A2(N110), .Y(n189) );
  NAND3X0_HVT U335 ( .A1(n195), .A2(n190), .A3(n189), .Y(n_quantized_data[4])
         );
  NAND2X0_HVT U336 ( .A1(n193), .A2(N41), .Y(n192) );
  NAND2X0_HVT U337 ( .A1(n194), .A2(N111), .Y(n191) );
  NAND3X0_HVT U338 ( .A1(n195), .A2(n192), .A3(n191), .Y(n_quantized_data[5])
         );
  AO22X1_HVT U339 ( .A1(n194), .A2(N112), .A3(n193), .A4(N42), .Y(n197) );
  OR2X1_HVT U340 ( .A1(n197), .A2(n196), .Y(n_quantized_data[6]) );
endmodule


module conv_top ( clk, srstn, conv_start, fc_done, sram_rdata_a0, 
        sram_rdata_a1, sram_rdata_a2, sram_rdata_a3, sram_rdata_a4, 
        sram_rdata_a5, sram_rdata_a6, sram_rdata_a7, sram_rdata_a8, 
        sram_rdata_b0, sram_rdata_b1, sram_rdata_b2, sram_rdata_b3, 
        sram_rdata_b4, sram_rdata_b5, sram_rdata_b6, sram_rdata_b7, 
        sram_rdata_b8, sram_rdata_weight, sram_raddr_weight, sram_raddr_a0, 
        sram_raddr_a1, sram_raddr_a2, sram_raddr_a3, sram_raddr_a4, 
        sram_raddr_a5, sram_raddr_a6, sram_raddr_a7, sram_raddr_a8, 
        sram_write_enable_b0, sram_write_enable_b1, sram_write_enable_b2, 
        sram_write_enable_b3, sram_write_enable_b4, sram_write_enable_b5, 
        sram_write_enable_b6, sram_write_enable_b7, sram_write_enable_b8, 
        sram_bytemask_b, sram_waddr_b, sram_wdata_b, sram_raddr_b0, 
        sram_raddr_b1, sram_raddr_b2, sram_raddr_b3, sram_raddr_b4, 
        sram_raddr_b5, sram_raddr_b6, sram_raddr_b7, sram_raddr_b8, 
        sram_write_enable_c0, sram_write_enable_c1, sram_write_enable_c2, 
        sram_write_enable_c3, sram_write_enable_c4, sram_bytemask_c, 
        sram_waddr_c, sram_wdata_c, sram_write_enable_d0, sram_write_enable_d1, 
        sram_write_enable_d2, sram_write_enable_d3, sram_write_enable_d4, 
        sram_bytemask_d, sram_waddr_d, sram_wdata_d, conv1_done, conv_done, 
        mem_sel );
  input [31:0] sram_rdata_a0;
  input [31:0] sram_rdata_a1;
  input [31:0] sram_rdata_a2;
  input [31:0] sram_rdata_a3;
  input [31:0] sram_rdata_a4;
  input [31:0] sram_rdata_a5;
  input [31:0] sram_rdata_a6;
  input [31:0] sram_rdata_a7;
  input [31:0] sram_rdata_a8;
  input [31:0] sram_rdata_b0;
  input [31:0] sram_rdata_b1;
  input [31:0] sram_rdata_b2;
  input [31:0] sram_rdata_b3;
  input [31:0] sram_rdata_b4;
  input [31:0] sram_rdata_b5;
  input [31:0] sram_rdata_b6;
  input [31:0] sram_rdata_b7;
  input [31:0] sram_rdata_b8;
  input [99:0] sram_rdata_weight;
  output [16:0] sram_raddr_weight;
  output [9:0] sram_raddr_a0;
  output [9:0] sram_raddr_a1;
  output [9:0] sram_raddr_a2;
  output [9:0] sram_raddr_a3;
  output [9:0] sram_raddr_a4;
  output [9:0] sram_raddr_a5;
  output [9:0] sram_raddr_a6;
  output [9:0] sram_raddr_a7;
  output [9:0] sram_raddr_a8;
  output [3:0] sram_bytemask_b;
  output [9:0] sram_waddr_b;
  output [7:0] sram_wdata_b;
  output [9:0] sram_raddr_b0;
  output [9:0] sram_raddr_b1;
  output [9:0] sram_raddr_b2;
  output [9:0] sram_raddr_b3;
  output [9:0] sram_raddr_b4;
  output [9:0] sram_raddr_b5;
  output [9:0] sram_raddr_b6;
  output [9:0] sram_raddr_b7;
  output [9:0] sram_raddr_b8;
  output [3:0] sram_bytemask_c;
  output [9:0] sram_waddr_c;
  output [7:0] sram_wdata_c;
  output [3:0] sram_bytemask_d;
  output [9:0] sram_waddr_d;
  output [7:0] sram_wdata_d;
  input clk, srstn, conv_start, fc_done;
  output sram_write_enable_b0, sram_write_enable_b1, sram_write_enable_b2,
         sram_write_enable_b3, sram_write_enable_b4, sram_write_enable_b5,
         sram_write_enable_b6, sram_write_enable_b7, sram_write_enable_b8,
         sram_write_enable_c0, sram_write_enable_c1, sram_write_enable_c2,
         sram_write_enable_c3, sram_write_enable_c4, sram_write_enable_d0,
         sram_write_enable_d1, sram_write_enable_d2, sram_write_enable_d3,
         sram_write_enable_d4, conv1_done, conv_done, mem_sel;
  wire   load_conv1_bias_enable, conv1_bias_set_16_, conv1_bias_set_15_,
         conv1_bias_set_14_, conv1_bias_set_13_, conv1_bias_set_12_,
         conv1_bias_set_11_, conv1_bias_set_10_, conv1_bias_set_9_,
         conv1_bias_set_8_, conv1_bias_set_7_, conv1_bias_set_6_,
         conv1_bias_set_5_, conv1_bias_set_4_, conv1_bias_set_3_,
         conv1_bias_set_2_, conv1_bias_set_1_, conv1_bias_set_0_, set_7_,
         set_6_, set_5_, set_4_, set_3_, set_2_, set_1_, set_0_,
         load_conv2_bias0_enable, load_conv2_bias1_enable, data_out_31_,
         data_out_30_, data_out_29_, data_out_28_, data_out_27_, data_out_26_,
         data_out_25_, data_out_24_, data_out_23_, data_out_22_, data_out_21_,
         data_out_20_, data_out_19_, data_out_18_, data_out_17_, data_out_16_,
         data_out_15_, data_out_14_, data_out_13_, data_out_12_, data_out_11_,
         data_out_10_, data_out_9_, data_out_8_, data_out_7_, data_out_6_,
         data_out_5_, data_out_4_, data_out_3_, data_out_2_, data_out_1_,
         data_out_0_, n1, n2, n3;
  wire   [1:0] mode;
  wire   [3:0] box_sel;
  wire   [4:0] channel;
  wire   [99:0] conv1_weight;
  wire   [99:0] weight;
  wire   [287:0] src_window;
  wire   [3:0] bias_data;

  fsm fsm ( .clk(clk), .srstn(n3), .conv_start(conv_start), .conv1_done(
        conv1_done), .conv_done(conv_done), .fc_done(fc_done), .mode(mode), 
        .mem_sel(mem_sel) );
  conv_control conv_control ( .clk(clk), .srstn(srstn), .mode(mode), .mem_sel(
        mem_sel), .conv1_done(conv1_done), .sram_raddr_weight(
        sram_raddr_weight), .box_sel(box_sel), .load_conv1_bias_enable(
        load_conv1_bias_enable), .conv1_bias_set({conv1_bias_set_16_, 
        conv1_bias_set_15_, conv1_bias_set_14_, conv1_bias_set_13_, 
        conv1_bias_set_12_, conv1_bias_set_11_, conv1_bias_set_10_, 
        conv1_bias_set_9_, conv1_bias_set_8_, conv1_bias_set_7_, 
        conv1_bias_set_6_, conv1_bias_set_5_, conv1_bias_set_4_, 
        conv1_bias_set_3_, conv1_bias_set_2_, conv1_bias_set_1_, 
        conv1_bias_set_0_}), .sram_raddr_a0(sram_raddr_a0), .sram_raddr_a1(
        sram_raddr_a1), .sram_raddr_a2(sram_raddr_a2), .sram_raddr_a3(
        sram_raddr_a3), .sram_raddr_a4(sram_raddr_a4), .sram_raddr_a5(
        sram_raddr_a5), .sram_raddr_a6(sram_raddr_a6), .sram_raddr_a7(
        sram_raddr_a7), .sram_raddr_a8(sram_raddr_a8), .sram_write_enable_b0(
        sram_write_enable_b0), .sram_write_enable_b1(sram_write_enable_b1), 
        .sram_write_enable_b2(sram_write_enable_b2), .sram_write_enable_b3(
        sram_write_enable_b3), .sram_write_enable_b4(sram_write_enable_b4), 
        .sram_write_enable_b5(sram_write_enable_b5), .sram_write_enable_b6(
        sram_write_enable_b6), .sram_write_enable_b7(sram_write_enable_b7), 
        .sram_write_enable_b8(sram_write_enable_b8), .sram_bytemask_b(
        sram_bytemask_b), .sram_waddr_b(sram_waddr_b), .conv_done(conv_done), 
        .channel(channel), .set({set_7_, set_6_, set_5_, set_4_, set_3_, 
        set_2_, set_1_, set_0_}), .load_conv2_bias0_enable(
        load_conv2_bias0_enable), .load_conv2_bias1_enable(
        load_conv2_bias1_enable), .sram_raddr_b0(sram_raddr_b0), 
        .sram_raddr_b1(sram_raddr_b1), .sram_raddr_b2(sram_raddr_b2), 
        .sram_raddr_b3(sram_raddr_b3), .sram_raddr_b4(sram_raddr_b4), 
        .sram_raddr_b5(sram_raddr_b5), .sram_raddr_b6(sram_raddr_b6), 
        .sram_raddr_b7(sram_raddr_b7), .sram_raddr_b8(sram_raddr_b8), 
        .sram_write_enable_c0(sram_write_enable_c0), .sram_write_enable_c1(
        sram_write_enable_c1), .sram_write_enable_c2(sram_write_enable_c2), 
        .sram_write_enable_c3(sram_write_enable_c3), .sram_write_enable_c4(
        sram_write_enable_c4), .sram_bytemask_c(sram_bytemask_c), 
        .sram_waddr_c(sram_waddr_c), .sram_write_enable_d0(
        sram_write_enable_d0), .sram_write_enable_d1(sram_write_enable_d1), 
        .sram_write_enable_d2(sram_write_enable_d2), .sram_write_enable_d3(
        sram_write_enable_d3), .sram_write_enable_d4(sram_write_enable_d4), 
        .sram_bytemask_d(sram_bytemask_d), .sram_waddr_d(sram_waddr_d) );
  data_reg data_reg ( .clk(clk), .srstn(n2), .mode(mode), .box_sel(box_sel), 
        .sram_rdata_a0(sram_rdata_a0), .sram_rdata_a1(sram_rdata_a1), 
        .sram_rdata_a2(sram_rdata_a2), .sram_rdata_a3(sram_rdata_a3), 
        .sram_rdata_a4(sram_rdata_a4), .sram_rdata_a5(sram_rdata_a5), 
        .sram_rdata_a6(sram_rdata_a6), .sram_rdata_a7(sram_rdata_a7), 
        .sram_rdata_a8(sram_rdata_a8), .sram_rdata_b0(sram_rdata_b0), 
        .sram_rdata_b1(sram_rdata_b1), .sram_rdata_b2(sram_rdata_b2), 
        .sram_rdata_b3(sram_rdata_b3), .sram_rdata_b4(sram_rdata_b4), 
        .sram_rdata_b5(sram_rdata_b5), .sram_rdata_b6(sram_rdata_b6), 
        .sram_rdata_b7(sram_rdata_b7), .sram_rdata_b8(sram_rdata_b8), 
        .sram_rdata_weight(sram_rdata_weight), .conv1_weight(conv1_weight), 
        .weight(weight), .src_window(src_window) );
  bias_sel bias_sel ( .clk(clk), .srstn(srstn), .mode(mode), 
        .load_conv1_bias_enable(load_conv1_bias_enable), 
        .load_conv2_bias0_enable(load_conv2_bias0_enable), 
        .load_conv2_bias1_enable(load_conv2_bias1_enable), .sram_rdata_weight(
        sram_rdata_weight), .bias_data(bias_data), .conv1_bias_set_5_(
        conv1_bias_set_5_), .conv1_bias_set_4_(conv1_bias_set_4_), 
        .conv1_bias_set_3_(conv1_bias_set_3_), .conv1_bias_set_2_(
        conv1_bias_set_2_), .conv1_bias_set_1_(conv1_bias_set_1_), 
        .conv1_bias_set_0_(conv1_bias_set_0_), .set_5_(set_5_), .set_4_(set_4_), .set_3_(set_3_), .set_2_(set_2_), .set_1_(set_1_), .set_0_(set_0_) );
  multiply_compare multiply_compare ( .clk(clk), .srstn(n3), .mode(mode), 
        .channel(channel), .conv1_sram_rdata_weight(conv1_weight), 
        .conv2_sram_rdata_weight(weight), .src_window(src_window), .data_out({
        data_out_31_, data_out_30_, data_out_29_, data_out_28_, data_out_27_, 
        data_out_26_, data_out_25_, data_out_24_, data_out_23_, data_out_22_, 
        data_out_21_, data_out_20_, data_out_19_, data_out_18_, data_out_17_, 
        data_out_16_, data_out_15_, data_out_14_, data_out_13_, data_out_12_, 
        data_out_11_, data_out_10_, data_out_9_, data_out_8_, data_out_7_, 
        data_out_6_, data_out_5_, data_out_4_, data_out_3_, data_out_2_, 
        data_out_1_, data_out_0_}) );
  quantize quantize ( .clk(clk), .srstn(n2), .bias_data(bias_data), .mode(mode), .quantized_data(sram_wdata_c), .ori_data_31_(data_out_31_), .ori_data_30_(
        data_out_30_), .ori_data_29_(data_out_29_), .ori_data_28_(data_out_28_), .ori_data_27_(data_out_27_), .ori_data_26_(data_out_26_), .ori_data_25_(
        data_out_25_), .ori_data_24_(data_out_24_), .ori_data_23_(data_out_23_), .ori_data_22_(data_out_22_), .ori_data_21_(data_out_21_), .ori_data_20_(
        data_out_20_), .ori_data_19_(data_out_19_), .ori_data_18_(data_out_18_), .ori_data_17_(data_out_17_), .ori_data_16_(data_out_16_), .ori_data_15_(
        data_out_15_), .ori_data_14_(data_out_14_), .ori_data_13_(data_out_13_), .ori_data_12_(data_out_12_), .ori_data_11_(data_out_11_), .ori_data_10_(
        data_out_10_), .ori_data_9_(data_out_9_), .ori_data_8_(data_out_8_), 
        .ori_data_7_(data_out_7_), .ori_data_6_(data_out_6_), .ori_data_5_(
        data_out_5_) );
  INVX1_HVT U1 ( .A(srstn), .Y(n1) );
  INVX1_HVT U2 ( .A(n1), .Y(n3) );
  INVX0_HVT U3 ( .A(n1), .Y(n2) );
  DELLN1X2_HVT U4 ( .A(sram_wdata_c[0]), .Y(sram_wdata_b[0]) );
  DELLN1X2_HVT U5 ( .A(sram_wdata_c[1]), .Y(sram_wdata_b[1]) );
  DELLN1X2_HVT U6 ( .A(sram_wdata_c[2]), .Y(sram_wdata_d[2]) );
  DELLN1X2_HVT U7 ( .A(sram_wdata_c[3]), .Y(sram_wdata_b[3]) );
  DELLN1X2_HVT U8 ( .A(sram_wdata_c[4]), .Y(sram_wdata_d[4]) );
  DELLN1X2_HVT U9 ( .A(sram_wdata_c[5]), .Y(sram_wdata_d[5]) );
  DELLN1X2_HVT U10 ( .A(sram_wdata_c[6]), .Y(sram_wdata_b[6]) );
  DELLN1X2_HVT U11 ( .A(sram_wdata_c[7]), .Y(sram_wdata_b[7]) );
  NBUFFX2_HVT U12 ( .A(sram_wdata_c[3]), .Y(sram_wdata_d[3]) );
  NBUFFX2_HVT U13 ( .A(sram_wdata_c[5]), .Y(sram_wdata_b[5]) );
  NBUFFX2_HVT U14 ( .A(sram_wdata_c[6]), .Y(sram_wdata_d[6]) );
  NBUFFX2_HVT U15 ( .A(sram_wdata_c[0]), .Y(sram_wdata_d[0]) );
  NBUFFX2_HVT U16 ( .A(sram_wdata_c[7]), .Y(sram_wdata_d[7]) );
  NBUFFX2_HVT U17 ( .A(sram_wdata_c[1]), .Y(sram_wdata_d[1]) );
  NBUFFX2_HVT U18 ( .A(sram_wdata_c[2]), .Y(sram_wdata_b[2]) );
  NBUFFX2_HVT U19 ( .A(sram_wdata_c[4]), .Y(sram_wdata_b[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fc_controller_mydesign_0 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net21977, n1;

  AND2X1_HVT main_gate ( .A1(net21977), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n1), .D(EN), .Q(net21977) );
  INVX0_HVT U1 ( .A(CLK), .Y(n1) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fc_controller_mydesign_1 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net21977, n2;

  AND2X1_HVT main_gate ( .A1(net21977), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net21977) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module fc_controller ( clk, srstn, conv_done, mem_sel, accumulate_reset, 
        fc_state, sram_sel, sram_raddr_c0, sram_raddr_c1, sram_raddr_c2, 
        sram_raddr_c3, sram_raddr_c4, sram_raddr_d0, sram_raddr_d1, 
        sram_raddr_d2, sram_raddr_d3, sram_raddr_d4, sram_raddr_e0, 
        sram_raddr_e1, sram_raddr_e2, sram_raddr_e3, sram_raddr_e4, 
        sram_write_enable_e0, sram_write_enable_e1, sram_write_enable_e2, 
        sram_write_enable_e3, sram_write_enable_e4, sram_write_enable_f, 
        sram_waddr, sram_bytemask, sram_raddr_weight, fc1_done, fc2_done );
  output [1:0] sram_sel;
  output [5:0] sram_raddr_c0;
  output [5:0] sram_raddr_c1;
  output [5:0] sram_raddr_c2;
  output [5:0] sram_raddr_c3;
  output [5:0] sram_raddr_c4;
  output [5:0] sram_raddr_d0;
  output [5:0] sram_raddr_d1;
  output [5:0] sram_raddr_d2;
  output [5:0] sram_raddr_d3;
  output [5:0] sram_raddr_d4;
  output [4:0] sram_raddr_e0;
  output [4:0] sram_raddr_e1;
  output [4:0] sram_raddr_e2;
  output [4:0] sram_raddr_e3;
  output [4:0] sram_raddr_e4;
  output [5:0] sram_waddr;
  output [3:0] sram_bytemask;
  output [14:0] sram_raddr_weight;
  input clk, srstn, conv_done, mem_sel;
  output accumulate_reset, fc_state, sram_write_enable_e0,
         sram_write_enable_e1, sram_write_enable_e2, sram_write_enable_e3,
         sram_write_enable_e4, sram_write_enable_f, fc1_done, fc2_done;
  wire   n_sram_sel_0_, n_write_enable, write_enable, write_e_sram_cnt_2_,
         n_write_enable_delay3, n_write_enable_delay1, n_write_enable_delay2,
         fetch_done, n_data_addr_complete, data_addr_complete, busy,
         n_conv_done_record, conv_done_record, N414, net21994, net22000,
         net22005, net22008, net22011, net22014, net22017, net22020, net22025,
         net22027, net22028, net22029, net22032, n17, n54, n55, n58, n60, n69,
         n99, n127, n128, n129, n1, n2, n5, n6, n7, n8, n10, n11, n12, n13,
         n18, n19, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n48, n49, n50, n51, n52, n53, n56, n57, n59, n61, n62, n63, n64, n65,
         n66, n67, n68, n70, n71, n72, n73, n148, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260;
  wire   [2:0] n_state;
  wire   [1:0] state;
  wire   [1:0] bytemask_sel;
  wire   [13:0] n_weight_cnt;
  wire   [5:1] n_row_cnt;

  SNPS_CLOCK_GATE_HIGH_fc_controller_mydesign_0 clk_gate_sram_waddr_reg ( 
        .CLK(clk), .EN(net21994), .ENCLK(net22020) );
  SNPS_CLOCK_GATE_HIGH_fc_controller_mydesign_1 clk_gate_write_e_sram_cnt_reg ( 
        .CLK(clk), .EN(net22025), .ENCLK(net22032) );
  DFFSSRX1_HVT state_reg_0_ ( .D(1'b0), .SETB(n36), .RSTB(n_state[0]), .CLK(
        clk), .Q(state[0]), .QN(n52) );
  DFFSSRX1_HVT n_write_enable_delay2_reg ( .D(1'b0), .SETB(n37), .RSTB(
        n_write_enable_delay3), .CLK(clk), .Q(n_write_enable_delay2) );
  DFFSSRX1_HVT n_write_enable_delay1_reg ( .D(1'b0), .SETB(n36), .RSTB(
        n_write_enable_delay2), .CLK(clk), .Q(n_write_enable_delay1) );
  DFFSSRX1_HVT n_write_enable_reg ( .D(1'b0), .SETB(n36), .RSTB(
        n_write_enable_delay1), .CLK(clk), .Q(n_write_enable), .QN(n43) );
  DFFSSRX1_HVT write_enable_reg ( .D(1'b0), .SETB(n37), .RSTB(n_write_enable), 
        .CLK(clk), .Q(write_enable), .QN(n57) );
  DFFSSRX1_HVT state_reg_2_ ( .D(1'b0), .SETB(n36), .RSTB(n_state[2]), .CLK(
        clk), .Q(n56), .QN(n69) );
  DFFSSRX1_HVT state_reg_1_ ( .D(1'b0), .SETB(n36), .RSTB(n_state[1]), .CLK(
        clk), .Q(state[1]) );
  DFFSSRX1_HVT data_addr_complete_reg ( .D(1'b0), .SETB(n36), .RSTB(
        n_data_addr_complete), .CLK(clk), .Q(data_addr_complete), .QN(n63) );
  DFFSSRX1_HVT row_cnt_reg_5_ ( .D(1'b0), .SETB(n36), .RSTB(n_row_cnt[5]), 
        .CLK(clk), .Q(sram_raddr_d3[5]), .QN(n51) );
  DFFSSRX1_HVT row_cnt_reg_4_ ( .D(1'b0), .SETB(n36), .RSTB(n_row_cnt[4]), 
        .CLK(clk), .Q(sram_raddr_e3[4]), .QN(n49) );
  DFFSSRX1_HVT row_cnt_reg_3_ ( .D(1'b0), .SETB(n37), .RSTB(n_row_cnt[3]), 
        .CLK(clk), .Q(sram_raddr_e3[3]), .QN(n44) );
  DFFSSRX1_HVT row_cnt_reg_2_ ( .D(1'b0), .SETB(n36), .RSTB(n_row_cnt[2]), 
        .CLK(clk), .Q(sram_raddr_e3[2]), .QN(n45) );
  DFFSSRX1_HVT row_cnt_reg_1_ ( .D(1'b0), .SETB(n36), .RSTB(n_row_cnt[1]), 
        .CLK(clk), .Q(sram_raddr_e3[1]), .QN(n53) );
  DFFSSRX1_HVT row_cnt_reg_0_ ( .D(1'b0), .SETB(n37), .RSTB(n209), .CLK(clk), 
        .Q(sram_raddr_e3[0]), .QN(n50) );
  DFFSSRX1_HVT weight_cnt_reg_12_ ( .D(1'b0), .SETB(n36), .RSTB(n60), .CLK(clk), .Q(sram_raddr_weight[12]) );
  DFFSSRX1_HVT weight_cnt_reg_0_ ( .D(1'b0), .SETB(n36), .RSTB(n_weight_cnt[0]), .CLK(clk), .Q(sram_raddr_weight[0]), .QN(n64) );
  DFFSSRX1_HVT weight_cnt_reg_10_ ( .D(1'b0), .SETB(n37), .RSTB(n199), .CLK(
        clk), .Q(sram_raddr_weight[10]), .QN(n68) );
  DFFSSRX1_HVT weight_cnt_reg_11_ ( .D(1'b0), .SETB(n36), .RSTB(n200), .CLK(
        clk), .Q(sram_raddr_weight[11]), .QN(n70) );
  DFFSSRX1_HVT weight_cnt_reg_3_ ( .D(1'b0), .SETB(n36), .RSTB(n201), .CLK(clk), .Q(sram_raddr_weight[3]), .QN(n72) );
  DFFSSRX1_HVT weight_cnt_reg_4_ ( .D(1'b0), .SETB(n36), .RSTB(n204), .CLK(clk), .Q(sram_raddr_weight[4]), .QN(n59) );
  DFFSSRX1_HVT weight_cnt_reg_6_ ( .D(1'b0), .SETB(n37), .RSTB(n205), .CLK(clk), .Q(sram_raddr_weight[6]), .QN(n73) );
  DFFSSRX1_HVT weight_cnt_reg_5_ ( .D(1'b0), .SETB(n37), .RSTB(n_weight_cnt[5]), .CLK(clk), .Q(sram_raddr_weight[5]) );
  DFFSSRX1_HVT weight_cnt_reg_8_ ( .D(1'b0), .SETB(n37), .RSTB(n202), .CLK(clk), .Q(sram_raddr_weight[8]) );
  DFFSSRX1_HVT weight_cnt_reg_9_ ( .D(1'b0), .SETB(n36), .RSTB(n198), .CLK(clk), .Q(sram_raddr_weight[9]), .QN(n67) );
  DFFSSRX1_HVT weight_cnt_reg_7_ ( .D(1'b0), .SETB(n36), .RSTB(n206), .CLK(clk), .Q(sram_raddr_weight[7]), .QN(n66) );
  DFFSSRX1_HVT weight_cnt_reg_14_ ( .D(1'b0), .SETB(n37), .RSTB(n208), .CLK(
        clk), .Q(sram_raddr_weight[14]), .QN(n65) );
  DFFSSRX1_HVT weight_cnt_reg_13_ ( .D(1'b0), .SETB(n36), .RSTB(
        n_weight_cnt[13]), .CLK(clk), .Q(sram_raddr_weight[13]) );
  DFFSSRX1_HVT weight_cnt_reg_1_ ( .D(1'b0), .SETB(n37), .RSTB(n_weight_cnt[1]), .CLK(clk), .Q(sram_raddr_weight[1]) );
  DFFSSRX1_HVT weight_cnt_reg_2_ ( .D(1'b0), .SETB(n36), .RSTB(n203), .CLK(clk), .Q(sram_raddr_weight[2]), .QN(n61) );
  DFFSSRX1_HVT sram_sel_reg_0_ ( .D(1'b0), .SETB(n37), .RSTB(n_sram_sel_0_), 
        .CLK(clk), .Q(sram_sel[0]) );
  DFFSSRX1_HVT sram_sel_reg_1_ ( .D(n17), .SETB(n99), .RSTB(srstn), .CLK(clk), 
        .Q(sram_sel[1]) );
  DFFSSRX1_HVT fetch_done_reg ( .D(1'b0), .SETB(n37), .RSTB(n129), .CLK(clk), 
        .Q(fetch_done), .QN(n62) );
  DFFSSRX1_HVT fc2_done_reg ( .D(1'b0), .SETB(n37), .RSTB(n207), .CLK(clk), 
        .Q(fc2_done), .QN(n58) );
  DFFSSRX1_HVT fc1_done_reg ( .D(1'b0), .SETB(n37), .RSTB(n210), .CLK(clk), 
        .Q(fc1_done) );
  DFFSSRX1_HVT bytemask_sel_reg_0_ ( .D(1'b0), .SETB(n36), .RSTB(n128), .CLK(
        clk), .Q(bytemask_sel[0]), .QN(n48) );
  DFFSSRX1_HVT bytemask_sel_reg_1_ ( .D(1'b0), .SETB(n37), .RSTB(n127), .CLK(
        clk), .Q(bytemask_sel[1]), .QN(n42) );
  DFFSSRX1_HVT write_e_sram_cnt_reg_0_ ( .D(1'b0), .SETB(n36), .RSTB(net22029), 
        .CLK(net22032), .Q(n41), .QN(n55) );
  DFFSSRX1_HVT write_e_sram_cnt_reg_1_ ( .D(1'b0), .SETB(n37), .RSTB(net22028), 
        .CLK(net22032), .Q(n46), .QN(n54) );
  DFFSSRX1_HVT write_e_sram_cnt_reg_2_ ( .D(1'b0), .SETB(n37), .RSTB(net22027), 
        .CLK(net22032), .Q(write_e_sram_cnt_2_) );
  DFFSSRX1_HVT sram_waddr_reg_0_ ( .D(1'b0), .SETB(n37), .RSTB(net22017), 
        .CLK(net22020), .Q(sram_waddr[0]) );
  DFFSSRX1_HVT sram_waddr_reg_1_ ( .D(1'b0), .SETB(n37), .RSTB(net22014), 
        .CLK(net22020), .Q(sram_waddr[1]) );
  DFFSSRX1_HVT sram_waddr_reg_2_ ( .D(1'b0), .SETB(n37), .RSTB(net22011), 
        .CLK(net22020), .Q(sram_waddr[2]) );
  DFFSSRX1_HVT sram_waddr_reg_3_ ( .D(1'b0), .SETB(n36), .RSTB(net22008), 
        .CLK(net22020), .Q(sram_waddr[3]) );
  DFFSSRX1_HVT sram_waddr_reg_4_ ( .D(1'b0), .SETB(n36), .RSTB(net22005), 
        .CLK(net22020), .Q(sram_waddr[4]) );
  DFFSSRX1_HVT sram_waddr_reg_5_ ( .D(1'b0), .SETB(n37), .RSTB(net22000), 
        .CLK(net22020), .Q(sram_waddr[5]), .QN(n71) );
  DFFSSRX1_HVT busy_reg ( .D(1'b0), .SETB(n37), .RSTB(N414), .CLK(clk), .Q(
        busy) );
  DFFSSRX1_HVT conv_done_record_reg ( .D(1'b0), .SETB(n36), .RSTB(
        n_conv_done_record), .CLK(clk), .Q(conv_done_record) );
  OA221X1_HVT U3 ( .A1(1'b0), .A2(n174), .A3(n171), .A4(sram_raddr_e3[2]), 
        .A5(n19), .Y(n_row_cnt[2]) );
  OA221X1_HVT U4 ( .A1(1'b0), .A2(n248), .A3(sram_waddr[3]), .A4(n18), .A5(
        n251), .Y(net22008) );
  OA221X1_HVT U5 ( .A1(1'b0), .A2(n237), .A3(sram_raddr_weight[12]), .A4(n238), 
        .A5(n195), .Y(n60) );
  OA221X1_HVT U6 ( .A1(1'b0), .A2(n247), .A3(sram_waddr[4]), .A4(n246), .A5(
        n251), .Y(net22005) );
  OA221X1_HVT U7 ( .A1(1'b0), .A2(n195), .A3(sram_raddr_weight[8]), .A4(n224), 
        .A5(n223), .Y(n202) );
  OA221X1_HVT U8 ( .A1(1'b0), .A2(n236), .A3(sram_raddr_weight[13]), .A4(n219), 
        .A5(n195), .Y(n_weight_cnt[13]) );
  OA221X1_HVT U9 ( .A1(1'b0), .A2(n195), .A3(sram_raddr_weight[1]), .A4(
        sram_raddr_weight[0]), .A5(n218), .Y(n_weight_cnt[1]) );
  INVX0_HVT U10 ( .A(state[1]), .Y(n1) );
  NAND2X0_HVT U11 ( .A1(n161), .A2(n1), .Y(n168) );
  NOR4X0_HVT U12 ( .A1(state[0]), .A2(state[1]), .A3(n56), .A4(busy), .Y(n2)
         );
  AO222X1_HVT U13 ( .A1(n193), .A2(n62), .A3(n210), .A4(n197), .A5(n217), .A6(
        n2), .Y(n162) );
  INVX0_HVT U16 ( .A(n65), .Y(n5) );
  INVX0_HVT U17 ( .A(n236), .Y(n6) );
  OA221X1_HVT U18 ( .A1(n65), .A2(n236), .A3(n5), .A4(n6), .A5(n195), .Y(n208)
         );
  INVX0_HVT U19 ( .A(n66), .Y(n7) );
  INVX0_HVT U20 ( .A(n227), .Y(n8) );
  OA221X1_HVT U21 ( .A1(n66), .A2(n227), .A3(n7), .A4(n8), .A5(n195), .Y(n206)
         );
  NAND3X0_HVT U23 ( .A1(sram_waddr[3]), .A2(sram_waddr[4]), .A3(n250), .Y(n10)
         );
  OR3X1_HVT U24 ( .A1(sram_waddr[0]), .A2(sram_waddr[5]), .A3(n10), .Y(n11) );
  AO221X1_HVT U25 ( .A1(n197), .A2(sram_waddr[2]), .A3(n197), .A4(n11), .A5(
        n188), .Y(n251) );
  INVX0_HVT U26 ( .A(n231), .Y(n12) );
  INVX0_HVT U27 ( .A(n59), .Y(n13) );
  OA221X1_HVT U28 ( .A1(n231), .A2(n59), .A3(n12), .A4(n13), .A5(n195), .Y(
        n204) );
  INVX0_HVT U32 ( .A(n249), .Y(n18) );
  INVX0_HVT U33 ( .A(n172), .Y(n19) );
  AO21X1_HVT U35 ( .A1(sram_waddr[1]), .A2(sram_waddr[0]), .A3(sram_waddr[2]), 
        .Y(n21) );
  AND3X1_HVT U36 ( .A1(n249), .A2(n251), .A3(n21), .Y(net22011) );
  INVX0_HVT U37 ( .A(n172), .Y(n22) );
  INVX0_HVT U38 ( .A(sram_raddr_e3[3]), .Y(n23) );
  OA221X1_HVT U39 ( .A1(n172), .A2(sram_raddr_e3[3]), .A3(n22), .A4(n23), .A5(
        n174), .Y(n_row_cnt[3]) );
  AO21X1_HVT U40 ( .A1(n57), .A2(bytemask_sel[1]), .A3(sram_bytemask[1]), .Y(
        n24) );
  OA221X1_HVT U41 ( .A1(n24), .A2(sram_bytemask[2]), .A3(n24), .A4(
        write_enable), .A5(n58), .Y(n127) );
  INVX0_HVT U42 ( .A(n173), .Y(n25) );
  INVX0_HVT U43 ( .A(sram_raddr_e3[4]), .Y(n26) );
  OA221X1_HVT U44 ( .A1(n173), .A2(sram_raddr_e3[4]), .A3(n25), .A4(n26), .A5(
        n174), .Y(n_row_cnt[4]) );
  NOR4X0_HVT U45 ( .A1(sram_raddr_weight[0]), .A2(sram_raddr_weight[1]), .A3(
        n239), .A4(n203), .Y(n27) );
  NAND4X0_HVT U46 ( .A1(n202), .A2(n201), .A3(n204), .A4(n27), .Y(n28) );
  OR3X1_HVT U47 ( .A1(n205), .A2(n206), .A3(n28), .Y(n29) );
  NAND3X0_HVT U48 ( .A1(n199), .A2(n198), .A3(n200), .Y(n30) );
  NOR4X0_HVT U49 ( .A1(n60), .A2(n_weight_cnt[13]), .A3(n29), .A4(n30), .Y(n31) );
  OA221X1_HVT U50 ( .A1(data_addr_complete), .A2(n208), .A3(data_addr_complete), .A4(n31), .A5(n188), .Y(n_data_addr_complete) );
  INVX0_HVT U51 ( .A(bytemask_sel[0]), .Y(n32) );
  INVX0_HVT U52 ( .A(write_enable), .Y(n33) );
  OA221X1_HVT U53 ( .A1(bytemask_sel[0]), .A2(write_enable), .A3(n32), .A4(n33), .A5(n58), .Y(n128) );
  NAND2X0_HVT U54 ( .A1(n173), .A2(sram_raddr_e3[4]), .Y(n34) );
  HADDX1_HVT U55 ( .A0(n51), .B0(n34), .SO(n35) );
  AND2X1_HVT U56 ( .A1(n174), .A2(n35), .Y(n_row_cnt[5]) );
  INVX1_HVT U57 ( .A(n232), .Y(n238) );
  INVX2_HVT U58 ( .A(srstn), .Y(n36) );
  INVX0_HVT U59 ( .A(n237), .Y(n219) );
  INVX0_HVT U60 ( .A(n234), .Y(n233) );
  INVX0_HVT U61 ( .A(n221), .Y(n235) );
  INVX0_HVT U62 ( .A(n223), .Y(n222) );
  INVX0_HVT U63 ( .A(n227), .Y(n220) );
  INVX0_HVT U64 ( .A(n225), .Y(n228) );
  INVX0_HVT U65 ( .A(n247), .Y(n245) );
  INVX0_HVT U66 ( .A(n50), .Y(sram_raddr_e4[0]) );
  INVX0_HVT U67 ( .A(n38), .Y(sram_raddr_e4[1]) );
  INVX0_HVT U68 ( .A(n214), .Y(n215) );
  INVX0_HVT U69 ( .A(n50), .Y(sram_raddr_c1[0]) );
  INVX0_HVT U70 ( .A(n38), .Y(sram_raddr_c0[1]) );
  INVX0_HVT U71 ( .A(n50), .Y(sram_raddr_d2[0]) );
  INVX0_HVT U72 ( .A(n40), .Y(sram_raddr_c1[4]) );
  INVX0_HVT U73 ( .A(n49), .Y(sram_raddr_d3[4]) );
  INVX0_HVT U74 ( .A(n39), .Y(sram_raddr_c4[0]) );
  INVX0_HVT U75 ( .A(n53), .Y(sram_raddr_d3[1]) );
  INVX0_HVT U76 ( .A(n40), .Y(sram_raddr_d0[4]) );
  INVX0_HVT U77 ( .A(n39), .Y(sram_raddr_d1[0]) );
  INVX0_HVT U78 ( .A(n40), .Y(sram_raddr_c2[4]) );
  INVX0_HVT U79 ( .A(n39), .Y(sram_raddr_d3[0]) );
  INVX0_HVT U80 ( .A(n163), .Y(n165) );
  INVX0_HVT U81 ( .A(n39), .Y(sram_raddr_c3[0]) );
  INVX0_HVT U82 ( .A(n53), .Y(sram_raddr_d1[1]) );
  INVX0_HVT U83 ( .A(n49), .Y(sram_raddr_d4[4]) );
  INVX0_HVT U84 ( .A(n38), .Y(sram_raddr_c4[1]) );
  INVX0_HVT U85 ( .A(n49), .Y(sram_raddr_d2[4]) );
  INVX0_HVT U86 ( .A(n40), .Y(sram_raddr_c4[4]) );
  INVX0_HVT U87 ( .A(n53), .Y(sram_raddr_d2[1]) );
  INVX0_HVT U88 ( .A(n40), .Y(sram_raddr_e1[4]) );
  INVX0_HVT U89 ( .A(n38), .Y(sram_raddr_c2[1]) );
  INVX0_HVT U90 ( .A(n39), .Y(sram_raddr_d0[0]) );
  INVX0_HVT U91 ( .A(n53), .Y(sram_raddr_e1[1]) );
  INVX0_HVT U92 ( .A(n39), .Y(sram_raddr_e1[0]) );
  INVX0_HVT U93 ( .A(n40), .Y(sram_raddr_e2[4]) );
  INVX0_HVT U94 ( .A(n38), .Y(sram_raddr_d0[1]) );
  INVX0_HVT U95 ( .A(n53), .Y(sram_raddr_e2[1]) );
  INVX0_HVT U96 ( .A(n39), .Y(sram_raddr_e2[0]) );
  INVX0_HVT U97 ( .A(n39), .Y(sram_raddr_c0[0]) );
  INVX0_HVT U98 ( .A(n40), .Y(sram_raddr_e4[4]) );
  INVX0_HVT U99 ( .A(n38), .Y(sram_raddr_c3[1]) );
  INVX0_HVT U100 ( .A(n40), .Y(sram_raddr_e0[4]) );
  INVX0_HVT U101 ( .A(n53), .Y(sram_raddr_e0[1]) );
  INVX0_HVT U102 ( .A(n40), .Y(sram_raddr_c3[4]) );
  INVX0_HVT U103 ( .A(n39), .Y(sram_raddr_d4[0]) );
  INVX0_HVT U104 ( .A(n53), .Y(sram_raddr_d4[1]) );
  INVX0_HVT U105 ( .A(n38), .Y(sram_raddr_c1[1]) );
  INVX0_HVT U106 ( .A(n39), .Y(sram_raddr_e0[0]) );
  INVX0_HVT U107 ( .A(n40), .Y(sram_raddr_d1[4]) );
  INVX0_HVT U108 ( .A(n39), .Y(sram_raddr_c2[0]) );
  INVX0_HVT U109 ( .A(n40), .Y(sram_raddr_c0[4]) );
  INVX0_HVT U110 ( .A(n188), .Y(n184) );
  INVX0_HVT U111 ( .A(n148), .Y(sram_raddr_d1[5]) );
  INVX0_HVT U112 ( .A(n148), .Y(sram_raddr_d2[5]) );
  INVX0_HVT U113 ( .A(n148), .Y(sram_raddr_c4[5]) );
  INVX0_HVT U114 ( .A(n148), .Y(sram_raddr_c3[5]) );
  INVX0_HVT U115 ( .A(n148), .Y(sram_raddr_d0[5]) );
  INVX0_HVT U116 ( .A(n190), .Y(sram_raddr_e4[2]) );
  INVX0_HVT U117 ( .A(n166), .Y(sram_raddr_e4[3]) );
  INVX0_HVT U118 ( .A(n231), .Y(n229) );
  INVX0_HVT U119 ( .A(n148), .Y(sram_raddr_d4[5]) );
  INVX0_HVT U120 ( .A(n148), .Y(sram_raddr_c1[5]) );
  INVX0_HVT U121 ( .A(sram_waddr[0]), .Y(n252) );
  INVX0_HVT U122 ( .A(n166), .Y(sram_raddr_c0[3]) );
  INVX0_HVT U123 ( .A(n190), .Y(sram_raddr_c0[2]) );
  INVX0_HVT U124 ( .A(n148), .Y(sram_raddr_c0[5]) );
  INVX0_HVT U125 ( .A(sram_waddr[1]), .Y(n250) );
  INVX0_HVT U126 ( .A(n190), .Y(sram_raddr_c1[2]) );
  INVX0_HVT U127 ( .A(n166), .Y(sram_raddr_c1[3]) );
  INVX0_HVT U128 ( .A(n148), .Y(sram_raddr_c2[5]) );
  INVX0_HVT U129 ( .A(n44), .Y(sram_raddr_d0[3]) );
  INVX0_HVT U130 ( .A(n44), .Y(sram_raddr_c2[3]) );
  INVX0_HVT U131 ( .A(n45), .Y(sram_raddr_d0[2]) );
  INVX0_HVT U132 ( .A(n45), .Y(sram_raddr_c4[2]) );
  INVX0_HVT U133 ( .A(n44), .Y(sram_raddr_e0[3]) );
  INVX0_HVT U134 ( .A(n45), .Y(sram_raddr_e0[2]) );
  INVX0_HVT U135 ( .A(n44), .Y(sram_raddr_e1[3]) );
  INVX0_HVT U136 ( .A(n45), .Y(sram_raddr_e1[2]) );
  INVX0_HVT U137 ( .A(n44), .Y(sram_raddr_c4[3]) );
  INVX0_HVT U138 ( .A(n44), .Y(sram_raddr_d2[3]) );
  INVX0_HVT U139 ( .A(n45), .Y(sram_raddr_d4[2]) );
  INVX0_HVT U140 ( .A(n44), .Y(sram_raddr_d4[3]) );
  INVX0_HVT U141 ( .A(n44), .Y(sram_raddr_e2[3]) );
  INVX0_HVT U142 ( .A(n45), .Y(sram_raddr_e2[2]) );
  INVX0_HVT U143 ( .A(n45), .Y(sram_raddr_d1[2]) );
  INVX0_HVT U144 ( .A(n44), .Y(sram_raddr_d3[3]) );
  INVX0_HVT U145 ( .A(n45), .Y(sram_raddr_d2[2]) );
  INVX0_HVT U146 ( .A(n45), .Y(sram_raddr_c2[2]) );
  INVX0_HVT U147 ( .A(n45), .Y(sram_raddr_c3[2]) );
  INVX0_HVT U148 ( .A(n44), .Y(sram_raddr_c3[3]) );
  INVX0_HVT U149 ( .A(n45), .Y(sram_raddr_d3[2]) );
  INVX0_HVT U150 ( .A(n44), .Y(sram_raddr_d1[3]) );
  INVX2_HVT U151 ( .A(srstn), .Y(n37) );
  INVX1_HVT U152 ( .A(sram_raddr_e3[1]), .Y(n38) );
  INVX1_HVT U153 ( .A(sram_raddr_e3[0]), .Y(n39) );
  INVX1_HVT U154 ( .A(sram_raddr_e3[4]), .Y(n40) );
  INVX1_HVT U155 ( .A(n168), .Y(n193) );
  NAND3X0_HVT U156 ( .A1(n163), .A2(n186), .A3(n168), .Y(n195) );
  INVX1_HVT U157 ( .A(n197), .Y(n186) );
  AND2X1_HVT U158 ( .A1(n158), .A2(n52), .Y(n197) );
  INVX1_HVT U159 ( .A(sram_raddr_d3[5]), .Y(n148) );
  INVX1_HVT U160 ( .A(sram_raddr_e3[2]), .Y(n190) );
  INVX1_HVT U161 ( .A(sram_raddr_e3[3]), .Y(n166) );
  AO21X1_HVT U162 ( .A1(n188), .A2(n177), .A3(n162), .Y(n_state[0]) );
  AND2X1_HVT U163 ( .A1(n48), .A2(n42), .Y(sram_bytemask[3]) );
  AND2X1_HVT U164 ( .A1(bytemask_sel[0]), .A2(n42), .Y(sram_bytemask[2]) );
  AND2X1_HVT U165 ( .A1(bytemask_sel[0]), .A2(bytemask_sel[1]), .Y(
        sram_bytemask[0]) );
  INVX1_HVT U166 ( .A(n248), .Y(n246) );
  INVX1_HVT U167 ( .A(n177), .Y(n207) );
  NOR4X1_HVT U168 ( .A1(sram_raddr_weight[11]), .A2(sram_raddr_weight[10]), 
        .A3(sram_raddr_weight[9]), .A4(n213), .Y(n258) );
  OR2X1_HVT U169 ( .A1(n57), .A2(n243), .Y(n177) );
  AND2X1_HVT U170 ( .A1(state[1]), .A2(n69), .Y(n158) );
  NAND2X0_HVT U171 ( .A1(n177), .A2(n158), .Y(n160) );
  AND2X1_HVT U172 ( .A1(state[0]), .A2(n69), .Y(n161) );
  NAND2X0_HVT U173 ( .A1(n193), .A2(fetch_done), .Y(n159) );
  NAND3X0_HVT U174 ( .A1(n160), .A2(n186), .A3(n159), .Y(n_state[1]) );
  AND2X1_HVT U175 ( .A1(n161), .A2(state[1]), .Y(n188) );
  AND4X1_HVT U176 ( .A1(n257), .A2(write_enable), .A3(n240), .A4(
        sram_raddr_weight[0]), .Y(n210) );
  OR3X1_HVT U177 ( .A1(n188), .A2(n162), .A3(n_state[1]), .Y(N414) );
  NAND2X0_HVT U178 ( .A1(n188), .A2(n63), .Y(n163) );
  AND2X1_HVT U179 ( .A1(n195), .A2(n64), .Y(n_weight_cnt[0]) );
  AND4X1_HVT U180 ( .A1(n53), .A2(n51), .A3(n50), .A4(sram_raddr_e3[4]), .Y(
        n164) );
  NAND3X0_HVT U181 ( .A1(n164), .A2(sram_raddr_e3[3]), .A3(n190), .Y(n175) );
  NAND2X0_HVT U182 ( .A1(n165), .A2(n175), .Y(n169) );
  AND2X1_HVT U183 ( .A1(sram_raddr_e3[1]), .A2(sram_raddr_e3[0]), .Y(n171) );
  AND2X1_HVT U184 ( .A1(n171), .A2(sram_raddr_e3[2]), .Y(n172) );
  AND2X1_HVT U185 ( .A1(n166), .A2(n49), .Y(n192) );
  NAND3X0_HVT U186 ( .A1(n172), .A2(sram_raddr_d3[5]), .A3(n192), .Y(n176) );
  NAND2X0_HVT U187 ( .A1(n176), .A2(n197), .Y(n167) );
  NAND3X0_HVT U188 ( .A1(n169), .A2(n168), .A3(n167), .Y(n174) );
  AND2X1_HVT U189 ( .A1(n174), .A2(n50), .Y(n209) );
  AND2X1_HVT U190 ( .A1(n53), .A2(sram_raddr_e3[0]), .Y(n170) );
  AO22X1_HVT U191 ( .A1(n170), .A2(n174), .A3(n209), .A4(sram_raddr_e3[1]), 
        .Y(n_row_cnt[1]) );
  AND2X1_HVT U192 ( .A1(n172), .A2(sram_raddr_e3[3]), .Y(n173) );
  OAI22X1_HVT U193 ( .A1(n186), .A2(n176), .A3(n184), .A4(n175), .Y(
        n_write_enable_delay3) );
  AND2X1_HVT U194 ( .A1(n207), .A2(n188), .Y(n_state[2]) );
  NAND2X0_HVT U195 ( .A1(n225), .A2(n73), .Y(n178) );
  AND3X1_HVT U196 ( .A1(n178), .A2(n227), .A3(n195), .Y(n205) );
  NAND2X0_HVT U197 ( .A1(n218), .A2(n61), .Y(n179) );
  AND3X1_HVT U198 ( .A1(n195), .A2(n230), .A3(n179), .Y(n203) );
  NAND2X0_HVT U199 ( .A1(n230), .A2(n72), .Y(n180) );
  AND3X1_HVT U200 ( .A1(n195), .A2(n231), .A3(n180), .Y(n201) );
  NAND2X0_HVT U201 ( .A1(n70), .A2(n234), .Y(n181) );
  AND3X1_HVT U202 ( .A1(n195), .A2(n232), .A3(n181), .Y(n200) );
  NAND2X0_HVT U203 ( .A1(n68), .A2(n221), .Y(n182) );
  AND3X1_HVT U204 ( .A1(n195), .A2(n234), .A3(n182), .Y(n199) );
  NAND2X0_HVT U205 ( .A1(n67), .A2(n223), .Y(n183) );
  AND3X1_HVT U206 ( .A1(n195), .A2(n221), .A3(n183), .Y(n198) );
  AND3X1_HVT U207 ( .A1(n197), .A2(n260), .A3(n55), .Y(net22029) );
  NAND2X0_HVT U208 ( .A1(n186), .A2(n184), .Y(n185) );
  NAND2X0_HVT U209 ( .A1(write_enable), .A2(sram_bytemask[0]), .Y(n196) );
  AND2X1_HVT U210 ( .A1(n197), .A2(n260), .Y(n187) );
  AO21X1_HVT U211 ( .A1(n185), .A2(n196), .A3(n187), .Y(n244) );
  OR3X1_HVT U212 ( .A1(write_e_sram_cnt_2_), .A2(n255), .A3(n186), .Y(n254) );
  NAND3X0_HVT U213 ( .A1(n187), .A2(write_e_sram_cnt_2_), .A3(n255), .Y(n253)
         );
  NAND2X0_HVT U214 ( .A1(n197), .A2(write_enable), .Y(n189) );
  NOR2X0_HVT U215 ( .A1(write_e_sram_cnt_2_), .A2(n189), .Y(n259) );
  NAND2X0_HVT U216 ( .A1(n188), .A2(write_enable), .Y(sram_write_enable_f) );
  OR2X1_HVT U217 ( .A1(n260), .A2(n189), .Y(sram_write_enable_e4) );
  AND4X1_HVT U218 ( .A1(n190), .A2(n51), .A3(n50), .A4(sram_raddr_e3[1]), .Y(
        n191) );
  NAND3X0_HVT U219 ( .A1(n193), .A2(n192), .A3(n191), .Y(n194) );
  NAND2X0_HVT U220 ( .A1(n194), .A2(n43), .Y(accumulate_reset) );
  AND3X1_HVT U221 ( .A1(n197), .A2(n255), .A3(n256), .Y(net22028) );
  AND2X1_HVT U222 ( .A1(n239), .A2(n195), .Y(n_weight_cnt[5]) );
  NAND3X0_HVT U223 ( .A1(srstn), .A2(n197), .A3(n196), .Y(net22025) );
  OR4X1_HVT U224 ( .A1(sram_raddr_weight[7]), .A2(sram_raddr_weight[6]), .A3(
        sram_raddr_weight[4]), .A4(sram_raddr_weight[2]), .Y(n211) );
  OR3X1_HVT U225 ( .A1(sram_raddr_weight[8]), .A2(sram_raddr_weight[3]), .A3(
        n211), .Y(n212) );
  OR3X1_HVT U226 ( .A1(sram_raddr_weight[13]), .A2(sram_raddr_weight[12]), 
        .A3(n212), .Y(n214) );
  NOR3X0_HVT U227 ( .A1(sram_raddr_weight[0]), .A2(sram_raddr_weight[1]), .A3(
        n214), .Y(n241) );
  OR2X1_HVT U228 ( .A1(sram_raddr_weight[14]), .A2(sram_raddr_weight[5]), .Y(
        n213) );
  NAND2X0_HVT U229 ( .A1(n241), .A2(n258), .Y(n243) );
  AND2X1_HVT U230 ( .A1(sram_raddr_weight[1]), .A2(n215), .Y(n257) );
  AND3X1_HVT U231 ( .A1(sram_raddr_weight[14]), .A2(sram_raddr_weight[11]), 
        .A3(sram_raddr_weight[5]), .Y(n216) );
  AND3X1_HVT U232 ( .A1(sram_raddr_weight[10]), .A2(sram_raddr_weight[9]), 
        .A3(n216), .Y(n240) );
  OR2X1_HVT U233 ( .A1(conv_done_record), .A2(conv_done), .Y(n217) );
  AND2X1_HVT U234 ( .A1(n_state[1]), .A2(n_state[0]), .Y(fc_state) );
  AND2X1_HVT U235 ( .A1(busy), .A2(n217), .Y(n_conv_done_record) );
  NAND2X0_HVT U237 ( .A1(sram_raddr_weight[0]), .A2(sram_raddr_weight[1]), .Y(
        n218) );
  NAND3X0_HVT U238 ( .A1(sram_raddr_weight[2]), .A2(sram_raddr_weight[0]), 
        .A3(sram_raddr_weight[1]), .Y(n230) );
  NAND4X0_HVT U239 ( .A1(sram_raddr_weight[3]), .A2(sram_raddr_weight[2]), 
        .A3(sram_raddr_weight[0]), .A4(sram_raddr_weight[1]), .Y(n231) );
  AND2X1_HVT U240 ( .A1(sram_raddr_weight[4]), .A2(n229), .Y(n226) );
  NAND2X0_HVT U241 ( .A1(sram_raddr_weight[5]), .A2(n226), .Y(n225) );
  NAND2X0_HVT U242 ( .A1(sram_raddr_weight[6]), .A2(n228), .Y(n227) );
  AND2X1_HVT U243 ( .A1(sram_raddr_weight[7]), .A2(n220), .Y(n224) );
  NAND2X0_HVT U244 ( .A1(sram_raddr_weight[8]), .A2(n224), .Y(n223) );
  NAND2X0_HVT U245 ( .A1(sram_raddr_weight[9]), .A2(n222), .Y(n221) );
  NAND2X0_HVT U246 ( .A1(sram_raddr_weight[10]), .A2(n235), .Y(n234) );
  NAND2X0_HVT U247 ( .A1(sram_raddr_weight[11]), .A2(n233), .Y(n232) );
  NAND2X0_HVT U248 ( .A1(sram_raddr_weight[12]), .A2(n238), .Y(n237) );
  NAND2X0_HVT U249 ( .A1(sram_raddr_weight[13]), .A2(n219), .Y(n236) );
  OA21X1_HVT U250 ( .A1(sram_raddr_weight[5]), .A2(n226), .A3(n225), .Y(n239)
         );
  AND2X1_HVT U251 ( .A1(n241), .A2(n240), .Y(n17) );
  NAND2X0_HVT U252 ( .A1(sram_sel[0]), .A2(n243), .Y(n242) );
  OAI22X1_HVT U253 ( .A1(n17), .A2(n242), .A3(mem_sel), .A4(n243), .Y(
        n_sram_sel_0_) );
  NAND2X0_HVT U254 ( .A1(sram_sel[1]), .A2(n243), .Y(n99) );
  NAND3X0_HVT U255 ( .A1(n55), .A2(n54), .A3(write_e_sram_cnt_2_), .Y(n260) );
  NAND2X0_HVT U256 ( .A1(srstn), .A2(n244), .Y(net21994) );
  NAND4X0_HVT U257 ( .A1(sram_waddr[2]), .A2(sram_waddr[0]), .A3(sram_waddr[1]), .A4(sram_waddr[3]), .Y(n248) );
  NAND2X0_HVT U258 ( .A1(sram_waddr[4]), .A2(n246), .Y(n247) );
  OA221X1_HVT U259 ( .A1(sram_waddr[5]), .A2(n245), .A3(n71), .A4(n247), .A5(
        n251), .Y(net22000) );
  NAND3X0_HVT U260 ( .A1(sram_waddr[2]), .A2(sram_waddr[0]), .A3(sram_waddr[1]), .Y(n249) );
  OA221X1_HVT U261 ( .A1(sram_waddr[1]), .A2(sram_waddr[0]), .A3(n250), .A4(
        n252), .A5(n251), .Y(net22014) );
  AND2X1_HVT U262 ( .A1(n252), .A2(n251), .Y(net22017) );
  NAND2X0_HVT U263 ( .A1(n41), .A2(n46), .Y(n255) );
  NAND2X0_HVT U264 ( .A1(n254), .A2(n253), .Y(net22027) );
  NAND2X0_HVT U265 ( .A1(n55), .A2(n54), .Y(n256) );
  AND3X1_HVT U266 ( .A1(n258), .A2(n257), .A3(n64), .Y(n129) );
  AND2X1_HVT U267 ( .A1(bytemask_sel[1]), .A2(n48), .Y(sram_bytemask[1]) );
  NAND3X0_HVT U268 ( .A1(n55), .A2(n54), .A3(n259), .Y(sram_write_enable_e0)
         );
  NAND3X0_HVT U269 ( .A1(n54), .A2(n259), .A3(n41), .Y(sram_write_enable_e1)
         );
  NAND3X0_HVT U270 ( .A1(n55), .A2(n259), .A3(n46), .Y(sram_write_enable_e2)
         );
  NAND3X0_HVT U271 ( .A1(n259), .A2(n41), .A3(n46), .Y(sram_write_enable_e3)
         );
endmodule


module fc_data_reg ( clk, srstn, sram_rdata_c0, sram_rdata_c1, sram_rdata_c2, 
        sram_rdata_c3, sram_rdata_c4, sram_rdata_d0, sram_rdata_d1, 
        sram_rdata_d2, sram_rdata_d3, sram_rdata_d4, sram_rdata_e0, 
        sram_rdata_e1, sram_rdata_e2, sram_rdata_e3, sram_rdata_e4, sram_sel, 
        src_window );
  input [31:0] sram_rdata_c0;
  input [31:0] sram_rdata_c1;
  input [31:0] sram_rdata_c2;
  input [31:0] sram_rdata_c3;
  input [31:0] sram_rdata_c4;
  input [31:0] sram_rdata_d0;
  input [31:0] sram_rdata_d1;
  input [31:0] sram_rdata_d2;
  input [31:0] sram_rdata_d3;
  input [31:0] sram_rdata_d4;
  input [31:0] sram_rdata_e0;
  input [31:0] sram_rdata_e1;
  input [31:0] sram_rdata_e2;
  input [31:0] sram_rdata_e3;
  input [31:0] sram_rdata_e4;
  input [1:0] sram_sel;
  output [159:0] src_window;
  input clk, srstn;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45;
  wire   [159:0] n_src_box;

  DFFSSRX1_HVT src_box_reg_159_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[159]), 
        .CLK(clk), .Q(src_window[159]) );
  DFFSSRX1_HVT src_box_reg_158_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[158]), 
        .CLK(clk), .Q(src_window[158]) );
  DFFSSRX1_HVT src_box_reg_157_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[157]), 
        .CLK(clk), .Q(src_window[157]) );
  DFFSSRX1_HVT src_box_reg_156_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[156]), 
        .CLK(clk), .Q(src_window[156]) );
  DFFSSRX1_HVT src_box_reg_155_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[155]), 
        .CLK(clk), .Q(src_window[155]) );
  DFFSSRX1_HVT src_box_reg_154_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[154]), 
        .CLK(clk), .Q(src_window[154]) );
  DFFSSRX1_HVT src_box_reg_153_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[153]), 
        .CLK(clk), .Q(src_window[153]) );
  DFFSSRX1_HVT src_box_reg_152_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[152]), 
        .CLK(clk), .Q(src_window[152]) );
  DFFSSRX1_HVT src_box_reg_151_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[151]), 
        .CLK(clk), .Q(src_window[151]) );
  DFFSSRX1_HVT src_box_reg_150_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[150]), 
        .CLK(clk), .Q(src_window[150]) );
  DFFSSRX1_HVT src_box_reg_149_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[149]), 
        .CLK(clk), .Q(src_window[149]) );
  DFFSSRX1_HVT src_box_reg_148_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[148]), 
        .CLK(clk), .Q(src_window[148]) );
  DFFSSRX1_HVT src_box_reg_147_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[147]), 
        .CLK(clk), .Q(src_window[147]) );
  DFFSSRX1_HVT src_box_reg_146_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[146]), 
        .CLK(clk), .Q(src_window[146]) );
  DFFSSRX1_HVT src_box_reg_145_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[145]), 
        .CLK(clk), .Q(src_window[145]) );
  DFFSSRX1_HVT src_box_reg_144_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[144]), 
        .CLK(clk), .Q(src_window[144]) );
  DFFSSRX1_HVT src_box_reg_143_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[143]), 
        .CLK(clk), .Q(src_window[143]) );
  DFFSSRX1_HVT src_box_reg_142_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[142]), 
        .CLK(clk), .Q(src_window[142]) );
  DFFSSRX1_HVT src_box_reg_141_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[141]), 
        .CLK(clk), .Q(src_window[141]) );
  DFFSSRX1_HVT src_box_reg_140_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[140]), 
        .CLK(clk), .Q(src_window[140]) );
  DFFSSRX1_HVT src_box_reg_139_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[139]), 
        .CLK(clk), .Q(src_window[139]) );
  DFFSSRX1_HVT src_box_reg_138_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[138]), 
        .CLK(clk), .Q(src_window[138]) );
  DFFSSRX1_HVT src_box_reg_137_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[137]), 
        .CLK(clk), .Q(src_window[137]) );
  DFFSSRX1_HVT src_box_reg_136_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[136]), 
        .CLK(clk), .Q(src_window[136]) );
  DFFSSRX1_HVT src_box_reg_135_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[135]), 
        .CLK(clk), .Q(src_window[135]) );
  DFFSSRX1_HVT src_box_reg_134_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[134]), 
        .CLK(clk), .Q(src_window[134]) );
  DFFSSRX1_HVT src_box_reg_133_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[133]), 
        .CLK(clk), .Q(src_window[133]) );
  DFFSSRX1_HVT src_box_reg_132_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[132]), 
        .CLK(clk), .Q(src_window[132]) );
  DFFSSRX1_HVT src_box_reg_131_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[131]), 
        .CLK(clk), .Q(src_window[131]) );
  DFFSSRX1_HVT src_box_reg_130_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[130]), 
        .CLK(clk), .Q(src_window[130]) );
  DFFSSRX1_HVT src_box_reg_129_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[129]), 
        .CLK(clk), .Q(src_window[129]) );
  DFFSSRX1_HVT src_box_reg_128_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[128]), 
        .CLK(clk), .Q(src_window[128]) );
  DFFSSRX1_HVT src_box_reg_127_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[127]), 
        .CLK(clk), .Q(src_window[127]) );
  DFFSSRX1_HVT src_box_reg_126_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[126]), 
        .CLK(clk), .Q(src_window[126]) );
  DFFSSRX1_HVT src_box_reg_125_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[125]), 
        .CLK(clk), .Q(src_window[125]) );
  DFFSSRX1_HVT src_box_reg_124_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[124]), 
        .CLK(clk), .Q(src_window[124]) );
  DFFSSRX1_HVT src_box_reg_123_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[123]), 
        .CLK(clk), .Q(src_window[123]) );
  DFFSSRX1_HVT src_box_reg_122_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[122]), 
        .CLK(clk), .Q(src_window[122]) );
  DFFSSRX1_HVT src_box_reg_121_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[121]), 
        .CLK(clk), .Q(src_window[121]) );
  DFFSSRX1_HVT src_box_reg_120_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[120]), 
        .CLK(clk), .Q(src_window[120]) );
  DFFSSRX1_HVT src_box_reg_119_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[119]), 
        .CLK(clk), .Q(src_window[119]) );
  DFFSSRX1_HVT src_box_reg_118_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[118]), 
        .CLK(clk), .Q(src_window[118]) );
  DFFSSRX1_HVT src_box_reg_117_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[117]), 
        .CLK(clk), .Q(src_window[117]) );
  DFFSSRX1_HVT src_box_reg_116_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[116]), 
        .CLK(clk), .Q(src_window[116]) );
  DFFSSRX1_HVT src_box_reg_115_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[115]), 
        .CLK(clk), .Q(src_window[115]) );
  DFFSSRX1_HVT src_box_reg_114_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[114]), 
        .CLK(clk), .Q(src_window[114]) );
  DFFSSRX1_HVT src_box_reg_113_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[113]), 
        .CLK(clk), .Q(src_window[113]) );
  DFFSSRX1_HVT src_box_reg_112_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[112]), 
        .CLK(clk), .Q(src_window[112]) );
  DFFSSRX1_HVT src_box_reg_111_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[111]), 
        .CLK(clk), .Q(src_window[111]) );
  DFFSSRX1_HVT src_box_reg_110_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[110]), 
        .CLK(clk), .Q(src_window[110]) );
  DFFSSRX1_HVT src_box_reg_109_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[109]), 
        .CLK(clk), .Q(src_window[109]) );
  DFFSSRX1_HVT src_box_reg_108_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[108]), 
        .CLK(clk), .Q(src_window[108]) );
  DFFSSRX1_HVT src_box_reg_107_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[107]), 
        .CLK(clk), .Q(src_window[107]) );
  DFFSSRX1_HVT src_box_reg_106_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[106]), 
        .CLK(clk), .Q(src_window[106]) );
  DFFSSRX1_HVT src_box_reg_105_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[105]), 
        .CLK(clk), .Q(src_window[105]) );
  DFFSSRX1_HVT src_box_reg_104_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[104]), 
        .CLK(clk), .Q(src_window[104]) );
  DFFSSRX1_HVT src_box_reg_103_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[103]), 
        .CLK(clk), .Q(src_window[103]) );
  DFFSSRX1_HVT src_box_reg_102_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[102]), 
        .CLK(clk), .Q(src_window[102]) );
  DFFSSRX1_HVT src_box_reg_101_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[101]), 
        .CLK(clk), .Q(src_window[101]) );
  DFFSSRX1_HVT src_box_reg_100_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[100]), 
        .CLK(clk), .Q(src_window[100]) );
  DFFSSRX1_HVT src_box_reg_99_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[99]), 
        .CLK(clk), .Q(src_window[99]) );
  DFFSSRX1_HVT src_box_reg_98_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[98]), 
        .CLK(clk), .Q(src_window[98]) );
  DFFSSRX1_HVT src_box_reg_97_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[97]), 
        .CLK(clk), .Q(src_window[97]) );
  DFFSSRX1_HVT src_box_reg_96_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[96]), 
        .CLK(clk), .Q(src_window[96]) );
  DFFSSRX1_HVT src_box_reg_95_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[95]), 
        .CLK(clk), .Q(src_window[95]) );
  DFFSSRX1_HVT src_box_reg_94_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[94]), 
        .CLK(clk), .Q(src_window[94]) );
  DFFSSRX1_HVT src_box_reg_93_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[93]), 
        .CLK(clk), .Q(src_window[93]) );
  DFFSSRX1_HVT src_box_reg_92_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[92]), 
        .CLK(clk), .Q(src_window[92]) );
  DFFSSRX1_HVT src_box_reg_91_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[91]), 
        .CLK(clk), .Q(src_window[91]) );
  DFFSSRX1_HVT src_box_reg_90_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[90]), 
        .CLK(clk), .Q(src_window[90]) );
  DFFSSRX1_HVT src_box_reg_89_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[89]), 
        .CLK(clk), .Q(src_window[89]) );
  DFFSSRX1_HVT src_box_reg_88_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[88]), 
        .CLK(clk), .Q(src_window[88]) );
  DFFSSRX1_HVT src_box_reg_87_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[87]), 
        .CLK(clk), .Q(src_window[87]) );
  DFFSSRX1_HVT src_box_reg_86_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[86]), 
        .CLK(clk), .Q(src_window[86]) );
  DFFSSRX1_HVT src_box_reg_85_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[85]), 
        .CLK(clk), .Q(src_window[85]) );
  DFFSSRX1_HVT src_box_reg_84_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[84]), 
        .CLK(clk), .Q(src_window[84]) );
  DFFSSRX1_HVT src_box_reg_83_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[83]), 
        .CLK(clk), .Q(src_window[83]) );
  DFFSSRX1_HVT src_box_reg_82_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[82]), 
        .CLK(clk), .Q(src_window[82]) );
  DFFSSRX1_HVT src_box_reg_81_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[81]), 
        .CLK(clk), .Q(src_window[81]) );
  DFFSSRX1_HVT src_box_reg_80_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[80]), 
        .CLK(clk), .Q(src_window[80]) );
  DFFSSRX1_HVT src_box_reg_79_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[79]), 
        .CLK(clk), .Q(src_window[79]) );
  DFFSSRX1_HVT src_box_reg_78_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[78]), 
        .CLK(clk), .Q(src_window[78]) );
  DFFSSRX1_HVT src_box_reg_77_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[77]), 
        .CLK(clk), .Q(src_window[77]) );
  DFFSSRX1_HVT src_box_reg_76_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[76]), 
        .CLK(clk), .Q(src_window[76]) );
  DFFSSRX1_HVT src_box_reg_75_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[75]), 
        .CLK(clk), .Q(src_window[75]) );
  DFFSSRX1_HVT src_box_reg_74_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[74]), 
        .CLK(clk), .Q(src_window[74]) );
  DFFSSRX1_HVT src_box_reg_73_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[73]), 
        .CLK(clk), .Q(src_window[73]) );
  DFFSSRX1_HVT src_box_reg_72_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[72]), 
        .CLK(clk), .Q(src_window[72]) );
  DFFSSRX1_HVT src_box_reg_71_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[71]), 
        .CLK(clk), .Q(src_window[71]) );
  DFFSSRX1_HVT src_box_reg_70_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[70]), 
        .CLK(clk), .Q(src_window[70]) );
  DFFSSRX1_HVT src_box_reg_69_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[69]), 
        .CLK(clk), .Q(src_window[69]) );
  DFFSSRX1_HVT src_box_reg_68_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[68]), 
        .CLK(clk), .Q(src_window[68]) );
  DFFSSRX1_HVT src_box_reg_67_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[67]), 
        .CLK(clk), .Q(src_window[67]) );
  DFFSSRX1_HVT src_box_reg_66_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[66]), 
        .CLK(clk), .Q(src_window[66]) );
  DFFSSRX1_HVT src_box_reg_65_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[65]), 
        .CLK(clk), .Q(src_window[65]) );
  DFFSSRX1_HVT src_box_reg_64_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[64]), 
        .CLK(clk), .Q(src_window[64]) );
  DFFSSRX1_HVT src_box_reg_63_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[63]), 
        .CLK(clk), .Q(src_window[63]) );
  DFFSSRX1_HVT src_box_reg_62_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[62]), 
        .CLK(clk), .Q(src_window[62]) );
  DFFSSRX1_HVT src_box_reg_61_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[61]), 
        .CLK(clk), .Q(src_window[61]) );
  DFFSSRX1_HVT src_box_reg_60_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[60]), 
        .CLK(clk), .Q(src_window[60]) );
  DFFSSRX1_HVT src_box_reg_59_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[59]), 
        .CLK(clk), .Q(src_window[59]) );
  DFFSSRX1_HVT src_box_reg_58_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[58]), 
        .CLK(clk), .Q(src_window[58]) );
  DFFSSRX1_HVT src_box_reg_57_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[57]), 
        .CLK(clk), .Q(src_window[57]) );
  DFFSSRX1_HVT src_box_reg_56_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[56]), 
        .CLK(clk), .Q(src_window[56]) );
  DFFSSRX1_HVT src_box_reg_55_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[55]), 
        .CLK(clk), .Q(src_window[55]) );
  DFFSSRX1_HVT src_box_reg_54_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[54]), 
        .CLK(clk), .Q(src_window[54]) );
  DFFSSRX1_HVT src_box_reg_53_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[53]), 
        .CLK(clk), .Q(src_window[53]) );
  DFFSSRX1_HVT src_box_reg_52_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[52]), 
        .CLK(clk), .Q(src_window[52]) );
  DFFSSRX1_HVT src_box_reg_51_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[51]), 
        .CLK(clk), .Q(src_window[51]) );
  DFFSSRX1_HVT src_box_reg_50_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[50]), 
        .CLK(clk), .Q(src_window[50]) );
  DFFSSRX1_HVT src_box_reg_49_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[49]), 
        .CLK(clk), .Q(src_window[49]) );
  DFFSSRX1_HVT src_box_reg_48_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[48]), 
        .CLK(clk), .Q(src_window[48]) );
  DFFSSRX1_HVT src_box_reg_47_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[47]), 
        .CLK(clk), .Q(src_window[47]) );
  DFFSSRX1_HVT src_box_reg_46_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[46]), 
        .CLK(clk), .Q(src_window[46]) );
  DFFSSRX1_HVT src_box_reg_45_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[45]), 
        .CLK(clk), .Q(src_window[45]) );
  DFFSSRX1_HVT src_box_reg_44_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[44]), 
        .CLK(clk), .Q(src_window[44]) );
  DFFSSRX1_HVT src_box_reg_43_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[43]), 
        .CLK(clk), .Q(src_window[43]) );
  DFFSSRX1_HVT src_box_reg_42_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[42]), 
        .CLK(clk), .Q(src_window[42]) );
  DFFSSRX1_HVT src_box_reg_41_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[41]), 
        .CLK(clk), .Q(src_window[41]) );
  DFFSSRX1_HVT src_box_reg_40_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[40]), 
        .CLK(clk), .Q(src_window[40]) );
  DFFSSRX1_HVT src_box_reg_39_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[39]), 
        .CLK(clk), .Q(src_window[39]) );
  DFFSSRX1_HVT src_box_reg_38_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[38]), 
        .CLK(clk), .Q(src_window[38]) );
  DFFSSRX1_HVT src_box_reg_37_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[37]), 
        .CLK(clk), .Q(src_window[37]) );
  DFFSSRX1_HVT src_box_reg_36_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[36]), 
        .CLK(clk), .Q(src_window[36]) );
  DFFSSRX1_HVT src_box_reg_35_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[35]), 
        .CLK(clk), .Q(src_window[35]) );
  DFFSSRX1_HVT src_box_reg_34_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[34]), 
        .CLK(clk), .Q(src_window[34]) );
  DFFSSRX1_HVT src_box_reg_33_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[33]), 
        .CLK(clk), .Q(src_window[33]) );
  DFFSSRX1_HVT src_box_reg_32_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[32]), 
        .CLK(clk), .Q(src_window[32]) );
  DFFSSRX1_HVT src_box_reg_31_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[31]), 
        .CLK(clk), .Q(src_window[31]) );
  DFFSSRX1_HVT src_box_reg_30_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[30]), 
        .CLK(clk), .Q(src_window[30]) );
  DFFSSRX1_HVT src_box_reg_29_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[29]), 
        .CLK(clk), .Q(src_window[29]) );
  DFFSSRX1_HVT src_box_reg_28_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[28]), 
        .CLK(clk), .Q(src_window[28]) );
  DFFSSRX1_HVT src_box_reg_27_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[27]), 
        .CLK(clk), .Q(src_window[27]) );
  DFFSSRX1_HVT src_box_reg_26_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[26]), 
        .CLK(clk), .Q(src_window[26]) );
  DFFSSRX1_HVT src_box_reg_25_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[25]), 
        .CLK(clk), .Q(src_window[25]) );
  DFFSSRX1_HVT src_box_reg_24_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[24]), 
        .CLK(clk), .Q(src_window[24]) );
  DFFSSRX1_HVT src_box_reg_23_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[23]), 
        .CLK(clk), .Q(src_window[23]) );
  DFFSSRX1_HVT src_box_reg_22_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[22]), 
        .CLK(clk), .Q(src_window[22]) );
  DFFSSRX1_HVT src_box_reg_21_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[21]), 
        .CLK(clk), .Q(src_window[21]) );
  DFFSSRX1_HVT src_box_reg_20_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[20]), 
        .CLK(clk), .Q(src_window[20]) );
  DFFSSRX1_HVT src_box_reg_19_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[19]), 
        .CLK(clk), .Q(src_window[19]) );
  DFFSSRX1_HVT src_box_reg_18_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[18]), 
        .CLK(clk), .Q(src_window[18]) );
  DFFSSRX1_HVT src_box_reg_17_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[17]), 
        .CLK(clk), .Q(src_window[17]) );
  DFFSSRX1_HVT src_box_reg_16_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[16]), 
        .CLK(clk), .Q(src_window[16]) );
  DFFSSRX1_HVT src_box_reg_15_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[15]), 
        .CLK(clk), .Q(src_window[15]) );
  DFFSSRX1_HVT src_box_reg_14_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[14]), 
        .CLK(clk), .Q(src_window[14]) );
  DFFSSRX1_HVT src_box_reg_13_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[13]), 
        .CLK(clk), .Q(src_window[13]) );
  DFFSSRX1_HVT src_box_reg_12_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[12]), 
        .CLK(clk), .Q(src_window[12]) );
  DFFSSRX1_HVT src_box_reg_11_ ( .D(1'b0), .SETB(n26), .RSTB(n_src_box[11]), 
        .CLK(clk), .Q(src_window[11]) );
  DFFSSRX1_HVT src_box_reg_10_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[10]), 
        .CLK(clk), .Q(src_window[10]) );
  DFFSSRX1_HVT src_box_reg_9_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[9]), 
        .CLK(clk), .Q(src_window[9]) );
  DFFSSRX1_HVT src_box_reg_8_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[8]), 
        .CLK(clk), .Q(src_window[8]) );
  DFFSSRX1_HVT src_box_reg_7_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[7]), 
        .CLK(clk), .Q(src_window[7]) );
  DFFSSRX1_HVT src_box_reg_6_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[6]), 
        .CLK(clk), .Q(src_window[6]) );
  DFFSSRX1_HVT src_box_reg_5_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[5]), 
        .CLK(clk), .Q(src_window[5]) );
  DFFSSRX1_HVT src_box_reg_4_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[4]), 
        .CLK(clk), .Q(src_window[4]) );
  DFFSSRX1_HVT src_box_reg_3_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[3]), 
        .CLK(clk), .Q(src_window[3]) );
  DFFSSRX1_HVT src_box_reg_2_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[2]), 
        .CLK(clk), .Q(src_window[2]) );
  DFFSSRX1_HVT src_box_reg_1_ ( .D(1'b0), .SETB(n45), .RSTB(n_src_box[1]), 
        .CLK(clk), .Q(src_window[1]) );
  DFFSSRX1_HVT src_box_reg_0_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[0]), 
        .CLK(clk), .Q(src_window[0]) );
  NAND2X0_HVT U3 ( .A1(n40), .A2(sram_sel[1]), .Y(n43) );
  INVX1_HVT U4 ( .A(n43), .Y(n30) );
  INVX2_HVT U5 ( .A(n25), .Y(n1) );
  INVX2_HVT U6 ( .A(srstn), .Y(n45) );
  INVX1_HVT U7 ( .A(n4), .Y(n8) );
  INVX1_HVT U8 ( .A(n4), .Y(n7) );
  INVX2_HVT U9 ( .A(n4), .Y(n2) );
  INVX1_HVT U10 ( .A(n43), .Y(n16) );
  INVX1_HVT U11 ( .A(n43), .Y(n18) );
  INVX1_HVT U12 ( .A(n20), .Y(n21) );
  INVX1_HVT U13 ( .A(n43), .Y(n17) );
  INVX1_HVT U14 ( .A(n43), .Y(n19) );
  INVX1_HVT U15 ( .A(n33), .Y(n13) );
  INVX1_HVT U16 ( .A(n33), .Y(n11) );
  INVX1_HVT U17 ( .A(n20), .Y(n23) );
  INVX1_HVT U18 ( .A(n33), .Y(n9) );
  INVX1_HVT U19 ( .A(n20), .Y(n24) );
  INVX1_HVT U20 ( .A(n33), .Y(n12) );
  INVX1_HVT U21 ( .A(n20), .Y(n22) );
  INVX1_HVT U22 ( .A(n33), .Y(n15) );
  INVX1_HVT U23 ( .A(n33), .Y(n14) );
  INVX1_HVT U24 ( .A(n33), .Y(n10) );
  INVX2_HVT U25 ( .A(n4), .Y(n3) );
  INVX1_HVT U26 ( .A(n31), .Y(n20) );
  INVX1_HVT U27 ( .A(n4), .Y(n6) );
  INVX1_HVT U28 ( .A(n4), .Y(n5) );
  INVX1_HVT U29 ( .A(n42), .Y(n4) );
  INVX2_HVT U30 ( .A(n25), .Y(n26) );
  INVX2_HVT U31 ( .A(n25), .Y(n28) );
  DELLN1X2_HVT U32 ( .A(n42), .Y(n37) );
  DELLN1X2_HVT U33 ( .A(n42), .Y(n39) );
  DELLN1X2_HVT U34 ( .A(n42), .Y(n38) );
  INVX2_HVT U35 ( .A(n25), .Y(n29) );
  INVX2_HVT U36 ( .A(n25), .Y(n27) );
  INVX1_HVT U37 ( .A(n33), .Y(n36) );
  INVX1_HVT U38 ( .A(n33), .Y(n35) );
  INVX1_HVT U39 ( .A(n33), .Y(n34) );
  AND2X1_HVT U40 ( .A1(n41), .A2(n40), .Y(n44) );
  INVX1_HVT U41 ( .A(n43), .Y(n32) );
  INVX1_HVT U42 ( .A(n43), .Y(n31) );
  INVX1_HVT U43 ( .A(n45), .Y(n25) );
  INVX1_HVT U44 ( .A(n44), .Y(n33) );
  INVX1_HVT U45 ( .A(sram_sel[1]), .Y(n41) );
  INVX1_HVT U46 ( .A(sram_sel[0]), .Y(n40) );
  AND2X1_HVT U47 ( .A1(n41), .A2(sram_sel[0]), .Y(n42) );
  AO222X1_HVT U48 ( .A1(n18), .A2(sram_rdata_e4[0]), .A3(n8), .A4(
        sram_rdata_d4[0]), .A5(n12), .A6(sram_rdata_c4[0]), .Y(n_src_box[0])
         );
  AO222X1_HVT U49 ( .A1(n16), .A2(sram_rdata_e4[1]), .A3(n14), .A4(
        sram_rdata_c4[1]), .A5(sram_rdata_d4[1]), .A6(n6), .Y(n_src_box[1]) );
  AO222X1_HVT U50 ( .A1(n16), .A2(sram_rdata_e4[8]), .A3(n36), .A4(
        sram_rdata_c4[8]), .A5(sram_rdata_d4[8]), .A6(n5), .Y(n_src_box[8]) );
  AO222X1_HVT U51 ( .A1(n16), .A2(sram_rdata_e4[9]), .A3(n36), .A4(
        sram_rdata_c4[9]), .A5(sram_rdata_d4[9]), .A6(n2), .Y(n_src_box[9]) );
  AO222X1_HVT U52 ( .A1(n21), .A2(sram_rdata_e4[16]), .A3(n36), .A4(
        sram_rdata_c4[16]), .A5(sram_rdata_d4[16]), .A6(n5), .Y(n_src_box[16])
         );
  AO222X1_HVT U53 ( .A1(n21), .A2(sram_rdata_e4[17]), .A3(n12), .A4(
        sram_rdata_c4[17]), .A5(sram_rdata_d4[17]), .A6(n6), .Y(n_src_box[17])
         );
  AO222X1_HVT U54 ( .A1(n23), .A2(sram_rdata_e4[18]), .A3(n9), .A4(
        sram_rdata_c4[18]), .A5(sram_rdata_d4[18]), .A6(n6), .Y(n_src_box[18])
         );
  AO222X1_HVT U55 ( .A1(n18), .A2(sram_rdata_e4[25]), .A3(n14), .A4(
        sram_rdata_c4[25]), .A5(sram_rdata_d4[25]), .A6(n8), .Y(n_src_box[25])
         );
  AO222X1_HVT U56 ( .A1(n16), .A2(sram_rdata_e4[26]), .A3(n12), .A4(
        sram_rdata_c4[26]), .A5(sram_rdata_d4[26]), .A6(n39), .Y(n_src_box[26]) );
  AO222X1_HVT U57 ( .A1(n21), .A2(sram_rdata_e3[0]), .A3(n12), .A4(
        sram_rdata_c3[0]), .A5(sram_rdata_d3[0]), .A6(n37), .Y(n_src_box[32])
         );
  AO222X1_HVT U58 ( .A1(n30), .A2(sram_rdata_e3[1]), .A3(n10), .A4(
        sram_rdata_c3[1]), .A5(sram_rdata_d3[1]), .A6(n2), .Y(n_src_box[33])
         );
  AO222X1_HVT U59 ( .A1(n19), .A2(sram_rdata_e3[2]), .A3(n10), .A4(
        sram_rdata_c3[2]), .A5(sram_rdata_d3[2]), .A6(n3), .Y(n_src_box[34])
         );
  AO222X1_HVT U60 ( .A1(n22), .A2(sram_rdata_e3[8]), .A3(n14), .A4(
        sram_rdata_c3[8]), .A5(sram_rdata_d3[8]), .A6(n37), .Y(n_src_box[40])
         );
  AO222X1_HVT U61 ( .A1(n17), .A2(sram_rdata_e3[9]), .A3(n13), .A4(
        sram_rdata_c3[9]), .A5(sram_rdata_d3[9]), .A6(n6), .Y(n_src_box[41])
         );
  AO222X1_HVT U62 ( .A1(n17), .A2(sram_rdata_e3[16]), .A3(n12), .A4(
        sram_rdata_c3[16]), .A5(sram_rdata_d3[16]), .A6(n5), .Y(n_src_box[48])
         );
  AO222X1_HVT U63 ( .A1(n17), .A2(sram_rdata_e3[17]), .A3(n10), .A4(
        sram_rdata_c3[17]), .A5(sram_rdata_d3[17]), .A6(n2), .Y(n_src_box[49])
         );
  AO222X1_HVT U64 ( .A1(n22), .A2(sram_rdata_e3[24]), .A3(n14), .A4(
        sram_rdata_c3[24]), .A5(sram_rdata_d3[24]), .A6(n7), .Y(n_src_box[56])
         );
  AO222X1_HVT U65 ( .A1(n22), .A2(sram_rdata_e3[25]), .A3(n14), .A4(
        sram_rdata_c3[25]), .A5(sram_rdata_d3[25]), .A6(n39), .Y(n_src_box[57]) );
  AO222X1_HVT U66 ( .A1(n30), .A2(sram_rdata_e2[0]), .A3(n9), .A4(
        sram_rdata_c2[0]), .A5(sram_rdata_d2[0]), .A6(n8), .Y(n_src_box[64])
         );
  AO222X1_HVT U67 ( .A1(n16), .A2(sram_rdata_e2[1]), .A3(n12), .A4(
        sram_rdata_c2[1]), .A5(sram_rdata_d2[1]), .A6(n3), .Y(n_src_box[65])
         );
  AO222X1_HVT U68 ( .A1(n18), .A2(sram_rdata_e2[2]), .A3(n10), .A4(
        sram_rdata_c2[2]), .A5(sram_rdata_d2[2]), .A6(n6), .Y(n_src_box[66])
         );
  AO222X1_HVT U69 ( .A1(n30), .A2(sram_rdata_e2[8]), .A3(n13), .A4(
        sram_rdata_c2[8]), .A5(sram_rdata_d2[8]), .A6(n38), .Y(n_src_box[72])
         );
  AO222X1_HVT U70 ( .A1(n30), .A2(sram_rdata_e2[9]), .A3(n12), .A4(
        sram_rdata_c2[9]), .A5(sram_rdata_d2[9]), .A6(n5), .Y(n_src_box[73])
         );
  AO222X1_HVT U71 ( .A1(n19), .A2(sram_rdata_e2[16]), .A3(n14), .A4(
        sram_rdata_c2[16]), .A5(sram_rdata_d2[16]), .A6(n5), .Y(n_src_box[80])
         );
  AO222X1_HVT U72 ( .A1(n19), .A2(sram_rdata_e2[17]), .A3(n13), .A4(
        sram_rdata_c2[17]), .A5(sram_rdata_d2[17]), .A6(n6), .Y(n_src_box[81])
         );
  AO222X1_HVT U73 ( .A1(n18), .A2(sram_rdata_e2[24]), .A3(n15), .A4(
        sram_rdata_c2[24]), .A5(sram_rdata_d2[24]), .A6(n5), .Y(n_src_box[88])
         );
  AO222X1_HVT U74 ( .A1(n18), .A2(sram_rdata_e2[25]), .A3(n35), .A4(
        sram_rdata_c2[25]), .A5(sram_rdata_d2[25]), .A6(n6), .Y(n_src_box[89])
         );
  AO222X1_HVT U75 ( .A1(n17), .A2(sram_rdata_e1[0]), .A3(n35), .A4(
        sram_rdata_c1[0]), .A5(sram_rdata_d1[0]), .A6(n2), .Y(n_src_box[96])
         );
  AO222X1_HVT U76 ( .A1(n23), .A2(sram_rdata_e1[1]), .A3(n35), .A4(
        sram_rdata_c1[1]), .A5(sram_rdata_d1[1]), .A6(n2), .Y(n_src_box[97])
         );
  AO222X1_HVT U77 ( .A1(n23), .A2(sram_rdata_e1[2]), .A3(n11), .A4(
        sram_rdata_c1[2]), .A5(sram_rdata_d1[2]), .A6(n3), .Y(n_src_box[98])
         );
  AO222X1_HVT U78 ( .A1(n24), .A2(sram_rdata_e1[8]), .A3(n10), .A4(
        sram_rdata_c1[8]), .A5(sram_rdata_d1[8]), .A6(n7), .Y(n_src_box[104])
         );
  AO222X1_HVT U79 ( .A1(n23), .A2(sram_rdata_e1[9]), .A3(n13), .A4(
        sram_rdata_c1[9]), .A5(sram_rdata_d1[9]), .A6(n8), .Y(n_src_box[105])
         );
  AO222X1_HVT U80 ( .A1(n24), .A2(sram_rdata_e1[10]), .A3(n9), .A4(
        sram_rdata_c1[10]), .A5(sram_rdata_d1[10]), .A6(n8), .Y(n_src_box[106]) );
  AO222X1_HVT U81 ( .A1(n22), .A2(sram_rdata_e1[16]), .A3(n14), .A4(
        sram_rdata_c1[16]), .A5(sram_rdata_d1[16]), .A6(n38), .Y(
        n_src_box[112]) );
  AO222X1_HVT U82 ( .A1(n30), .A2(sram_rdata_e1[17]), .A3(n11), .A4(
        sram_rdata_c1[17]), .A5(sram_rdata_d1[17]), .A6(n8), .Y(n_src_box[113]) );
  AO222X1_HVT U83 ( .A1(n16), .A2(sram_rdata_e1[24]), .A3(n11), .A4(
        sram_rdata_c1[24]), .A5(sram_rdata_d1[24]), .A6(n38), .Y(
        n_src_box[120]) );
  AO222X1_HVT U84 ( .A1(n18), .A2(sram_rdata_e1[25]), .A3(n13), .A4(
        sram_rdata_c1[25]), .A5(sram_rdata_d1[25]), .A6(n3), .Y(n_src_box[121]) );
  AO222X1_HVT U85 ( .A1(n19), .A2(sram_rdata_e1[26]), .A3(n9), .A4(
        sram_rdata_c1[26]), .A5(sram_rdata_d1[26]), .A6(n6), .Y(n_src_box[122]) );
  AO222X1_HVT U86 ( .A1(n19), .A2(sram_rdata_e0[0]), .A3(n13), .A4(
        sram_rdata_c0[0]), .A5(sram_rdata_d0[0]), .A6(n5), .Y(n_src_box[128])
         );
  AO222X1_HVT U87 ( .A1(n17), .A2(sram_rdata_e0[1]), .A3(n9), .A4(
        sram_rdata_c0[1]), .A5(sram_rdata_d0[1]), .A6(n7), .Y(n_src_box[129])
         );
  AO222X1_HVT U88 ( .A1(n24), .A2(sram_rdata_e0[2]), .A3(n15), .A4(
        sram_rdata_c0[2]), .A5(sram_rdata_d0[2]), .A6(n5), .Y(n_src_box[130])
         );
  AO222X1_HVT U89 ( .A1(n24), .A2(sram_rdata_e0[8]), .A3(n15), .A4(
        sram_rdata_c0[8]), .A5(sram_rdata_d0[8]), .A6(n6), .Y(n_src_box[136])
         );
  AO222X1_HVT U90 ( .A1(n30), .A2(sram_rdata_e0[9]), .A3(n11), .A4(
        sram_rdata_c0[9]), .A5(sram_rdata_d0[9]), .A6(n5), .Y(n_src_box[137])
         );
  AO222X1_HVT U91 ( .A1(n17), .A2(sram_rdata_e0[16]), .A3(n13), .A4(
        sram_rdata_c0[16]), .A5(sram_rdata_d0[16]), .A6(n3), .Y(n_src_box[144]) );
  AO222X1_HVT U92 ( .A1(n16), .A2(sram_rdata_e0[17]), .A3(n9), .A4(
        sram_rdata_c0[17]), .A5(sram_rdata_d0[17]), .A6(n37), .Y(
        n_src_box[145]) );
  AO222X1_HVT U93 ( .A1(n30), .A2(sram_rdata_e0[24]), .A3(n15), .A4(
        sram_rdata_c0[24]), .A5(sram_rdata_d0[24]), .A6(n39), .Y(
        n_src_box[152]) );
  AO222X1_HVT U94 ( .A1(n30), .A2(sram_rdata_e0[25]), .A3(n11), .A4(
        sram_rdata_c0[25]), .A5(sram_rdata_d0[25]), .A6(n7), .Y(n_src_box[153]) );
  AO222X1_HVT U95 ( .A1(n19), .A2(sram_rdata_e0[26]), .A3(n15), .A4(
        sram_rdata_c0[26]), .A5(sram_rdata_d0[26]), .A6(n3), .Y(n_src_box[154]) );
  AO222X1_HVT U96 ( .A1(n35), .A2(sram_rdata_c1[4]), .A3(n23), .A4(
        sram_rdata_e1[4]), .A5(sram_rdata_d1[4]), .A6(n7), .Y(n_src_box[100])
         );
  AO222X1_HVT U97 ( .A1(n35), .A2(sram_rdata_c1[5]), .A3(n31), .A4(
        sram_rdata_e1[5]), .A5(sram_rdata_d1[5]), .A6(n7), .Y(n_src_box[101])
         );
  AO222X1_HVT U98 ( .A1(n44), .A2(sram_rdata_c1[6]), .A3(n22), .A4(
        sram_rdata_e1[6]), .A5(sram_rdata_d1[6]), .A6(n39), .Y(n_src_box[102])
         );
  AO222X1_HVT U99 ( .A1(n15), .A2(sram_rdata_c1[7]), .A3(n21), .A4(
        sram_rdata_e1[7]), .A5(sram_rdata_d1[7]), .A6(n8), .Y(n_src_box[103])
         );
  AO222X1_HVT U100 ( .A1(n10), .A2(sram_rdata_c1[11]), .A3(n17), .A4(
        sram_rdata_e1[11]), .A5(sram_rdata_d1[11]), .A6(n3), .Y(n_src_box[107]) );
  AO222X1_HVT U101 ( .A1(n11), .A2(sram_rdata_c1[12]), .A3(n17), .A4(
        sram_rdata_e1[12]), .A5(sram_rdata_d1[12]), .A6(n2), .Y(n_src_box[108]) );
  AO222X1_HVT U102 ( .A1(n11), .A2(sram_rdata_c1[13]), .A3(n31), .A4(
        sram_rdata_e1[13]), .A5(sram_rdata_d1[13]), .A6(n6), .Y(n_src_box[109]) );
  AO222X1_HVT U103 ( .A1(n13), .A2(sram_rdata_c4[10]), .A3(n31), .A4(
        sram_rdata_e4[10]), .A5(sram_rdata_d4[10]), .A6(n39), .Y(n_src_box[10]) );
  AO222X1_HVT U104 ( .A1(n36), .A2(sram_rdata_c1[14]), .A3(n30), .A4(
        sram_rdata_e1[14]), .A5(sram_rdata_d1[14]), .A6(n3), .Y(n_src_box[110]) );
  AO222X1_HVT U105 ( .A1(n34), .A2(sram_rdata_c1[15]), .A3(n22), .A4(
        sram_rdata_e1[15]), .A5(sram_rdata_d1[15]), .A6(n5), .Y(n_src_box[111]) );
  AO222X1_HVT U106 ( .A1(n34), .A2(sram_rdata_c1[18]), .A3(n24), .A4(
        sram_rdata_e1[18]), .A5(sram_rdata_d1[18]), .A6(n7), .Y(n_src_box[114]) );
  AO222X1_HVT U107 ( .A1(n44), .A2(sram_rdata_c1[19]), .A3(n31), .A4(
        sram_rdata_e1[19]), .A5(sram_rdata_d1[19]), .A6(n38), .Y(
        n_src_box[115]) );
  AO222X1_HVT U108 ( .A1(n36), .A2(sram_rdata_c1[20]), .A3(n18), .A4(
        sram_rdata_e1[20]), .A5(sram_rdata_d1[20]), .A6(n2), .Y(n_src_box[116]) );
  AO222X1_HVT U109 ( .A1(n9), .A2(sram_rdata_c1[21]), .A3(n19), .A4(
        sram_rdata_e1[21]), .A5(sram_rdata_d1[21]), .A6(n37), .Y(
        n_src_box[117]) );
  AO222X1_HVT U110 ( .A1(n12), .A2(sram_rdata_c1[22]), .A3(n17), .A4(
        sram_rdata_e1[22]), .A5(sram_rdata_d1[22]), .A6(n39), .Y(
        n_src_box[118]) );
  AO222X1_HVT U111 ( .A1(n14), .A2(sram_rdata_c1[23]), .A3(n17), .A4(
        sram_rdata_e1[23]), .A5(sram_rdata_d1[23]), .A6(n3), .Y(n_src_box[119]) );
  AO222X1_HVT U112 ( .A1(n35), .A2(sram_rdata_c4[11]), .A3(n30), .A4(
        sram_rdata_e4[11]), .A5(sram_rdata_d4[11]), .A6(n42), .Y(n_src_box[11]) );
  AO222X1_HVT U113 ( .A1(n34), .A2(sram_rdata_c1[27]), .A3(n30), .A4(
        sram_rdata_e1[27]), .A5(sram_rdata_d1[27]), .A6(n37), .Y(
        n_src_box[123]) );
  AO222X1_HVT U114 ( .A1(n10), .A2(sram_rdata_c1[28]), .A3(n16), .A4(
        sram_rdata_e1[28]), .A5(sram_rdata_d1[28]), .A6(n39), .Y(
        n_src_box[124]) );
  AO222X1_HVT U115 ( .A1(n44), .A2(sram_rdata_c1[29]), .A3(n19), .A4(
        sram_rdata_e1[29]), .A5(sram_rdata_d1[29]), .A6(n39), .Y(
        n_src_box[125]) );
  AO222X1_HVT U116 ( .A1(n10), .A2(sram_rdata_c1[30]), .A3(n19), .A4(
        sram_rdata_e1[30]), .A5(sram_rdata_d1[30]), .A6(n3), .Y(n_src_box[126]) );
  AO222X1_HVT U117 ( .A1(n34), .A2(sram_rdata_c1[31]), .A3(n32), .A4(
        sram_rdata_e1[31]), .A5(sram_rdata_d1[31]), .A6(n7), .Y(n_src_box[127]) );
  AO222X1_HVT U118 ( .A1(n13), .A2(sram_rdata_c4[12]), .A3(n31), .A4(
        sram_rdata_e4[12]), .A5(sram_rdata_d4[12]), .A6(n3), .Y(n_src_box[12])
         );
  AO222X1_HVT U119 ( .A1(n15), .A2(sram_rdata_c0[3]), .A3(n21), .A4(
        sram_rdata_e0[3]), .A5(sram_rdata_d0[3]), .A6(n2), .Y(n_src_box[131])
         );
  AO222X1_HVT U120 ( .A1(n35), .A2(sram_rdata_c0[4]), .A3(n32), .A4(
        sram_rdata_e0[4]), .A5(sram_rdata_d0[4]), .A6(n2), .Y(n_src_box[132])
         );
  AO222X1_HVT U121 ( .A1(n36), .A2(sram_rdata_c0[5]), .A3(n23), .A4(
        sram_rdata_e0[5]), .A5(sram_rdata_d0[5]), .A6(n39), .Y(n_src_box[133])
         );
  AO222X1_HVT U122 ( .A1(n44), .A2(sram_rdata_c0[6]), .A3(n32), .A4(
        sram_rdata_e0[6]), .A5(sram_rdata_d0[6]), .A6(n37), .Y(n_src_box[134])
         );
  AO222X1_HVT U123 ( .A1(n13), .A2(sram_rdata_c0[7]), .A3(n21), .A4(
        sram_rdata_e0[7]), .A5(sram_rdata_d0[7]), .A6(n5), .Y(n_src_box[135])
         );
  AO222X1_HVT U124 ( .A1(n9), .A2(sram_rdata_c0[10]), .A3(n23), .A4(
        sram_rdata_e0[10]), .A5(sram_rdata_d0[10]), .A6(n42), .Y(
        n_src_box[138]) );
  AO222X1_HVT U125 ( .A1(n11), .A2(sram_rdata_c0[11]), .A3(n16), .A4(
        sram_rdata_e0[11]), .A5(sram_rdata_d0[11]), .A6(n6), .Y(n_src_box[139]) );
  AO222X1_HVT U126 ( .A1(n9), .A2(sram_rdata_c4[13]), .A3(n16), .A4(
        sram_rdata_e4[13]), .A5(sram_rdata_d4[13]), .A6(n38), .Y(n_src_box[13]) );
  AO222X1_HVT U127 ( .A1(n12), .A2(sram_rdata_c0[12]), .A3(n18), .A4(
        sram_rdata_e0[12]), .A5(sram_rdata_d0[12]), .A6(n37), .Y(
        n_src_box[140]) );
  AO222X1_HVT U128 ( .A1(n35), .A2(sram_rdata_c0[13]), .A3(n24), .A4(
        sram_rdata_e0[13]), .A5(sram_rdata_d0[13]), .A6(n3), .Y(n_src_box[141]) );
  AO222X1_HVT U129 ( .A1(n34), .A2(sram_rdata_c0[14]), .A3(n19), .A4(
        sram_rdata_e0[14]), .A5(sram_rdata_d0[14]), .A6(n38), .Y(
        n_src_box[142]) );
  AO222X1_HVT U130 ( .A1(n34), .A2(sram_rdata_c0[15]), .A3(n22), .A4(
        sram_rdata_e0[15]), .A5(sram_rdata_d0[15]), .A6(n37), .Y(
        n_src_box[143]) );
  AO222X1_HVT U131 ( .A1(n44), .A2(sram_rdata_c0[18]), .A3(n21), .A4(
        sram_rdata_e0[18]), .A5(sram_rdata_d0[18]), .A6(n38), .Y(
        n_src_box[146]) );
  AO222X1_HVT U132 ( .A1(n36), .A2(sram_rdata_c0[19]), .A3(n30), .A4(
        sram_rdata_e0[19]), .A5(sram_rdata_d0[19]), .A6(n7), .Y(n_src_box[147]) );
  AO222X1_HVT U133 ( .A1(n15), .A2(sram_rdata_c0[20]), .A3(n31), .A4(
        sram_rdata_e0[20]), .A5(sram_rdata_d0[20]), .A6(n6), .Y(n_src_box[148]) );
  AO222X1_HVT U134 ( .A1(n15), .A2(sram_rdata_c0[21]), .A3(n21), .A4(
        sram_rdata_e0[21]), .A5(sram_rdata_d0[21]), .A6(n42), .Y(
        n_src_box[149]) );
  AO222X1_HVT U135 ( .A1(n12), .A2(sram_rdata_c4[14]), .A3(n32), .A4(
        sram_rdata_e4[14]), .A5(sram_rdata_d4[14]), .A6(n6), .Y(n_src_box[14])
         );
  AO222X1_HVT U136 ( .A1(n36), .A2(sram_rdata_c0[22]), .A3(n18), .A4(
        sram_rdata_e0[22]), .A5(sram_rdata_d0[22]), .A6(n8), .Y(n_src_box[150]) );
  AO222X1_HVT U137 ( .A1(n34), .A2(sram_rdata_c0[23]), .A3(n21), .A4(
        sram_rdata_e0[23]), .A5(sram_rdata_d0[23]), .A6(n2), .Y(n_src_box[151]) );
  AO222X1_HVT U138 ( .A1(n10), .A2(sram_rdata_c0[27]), .A3(n24), .A4(
        sram_rdata_e0[27]), .A5(sram_rdata_d0[27]), .A6(n37), .Y(
        n_src_box[155]) );
  AO222X1_HVT U139 ( .A1(n44), .A2(sram_rdata_c0[28]), .A3(n22), .A4(
        sram_rdata_e0[28]), .A5(sram_rdata_d0[28]), .A6(n37), .Y(
        n_src_box[156]) );
  AO222X1_HVT U140 ( .A1(n11), .A2(sram_rdata_c0[29]), .A3(n16), .A4(
        sram_rdata_e0[29]), .A5(sram_rdata_d0[29]), .A6(n8), .Y(n_src_box[157]) );
  AO222X1_HVT U141 ( .A1(n34), .A2(sram_rdata_c0[30]), .A3(n19), .A4(
        sram_rdata_e0[30]), .A5(sram_rdata_d0[30]), .A6(n39), .Y(
        n_src_box[158]) );
  AO222X1_HVT U142 ( .A1(n12), .A2(sram_rdata_c0[31]), .A3(n17), .A4(
        sram_rdata_e0[31]), .A5(sram_rdata_d0[31]), .A6(n5), .Y(n_src_box[159]) );
  AO222X1_HVT U143 ( .A1(n14), .A2(sram_rdata_c4[15]), .A3(n32), .A4(
        sram_rdata_e4[15]), .A5(sram_rdata_d4[15]), .A6(n38), .Y(n_src_box[15]) );
  AO222X1_HVT U144 ( .A1(n35), .A2(sram_rdata_c4[19]), .A3(n22), .A4(
        sram_rdata_e4[19]), .A5(sram_rdata_d4[19]), .A6(n2), .Y(n_src_box[19])
         );
  AO222X1_HVT U145 ( .A1(n35), .A2(sram_rdata_c4[20]), .A3(n32), .A4(
        sram_rdata_e4[20]), .A5(sram_rdata_d4[20]), .A6(n38), .Y(n_src_box[20]) );
  AO222X1_HVT U146 ( .A1(n44), .A2(sram_rdata_c4[21]), .A3(n18), .A4(
        sram_rdata_e4[21]), .A5(sram_rdata_d4[21]), .A6(n42), .Y(n_src_box[21]) );
  AO222X1_HVT U147 ( .A1(n15), .A2(sram_rdata_c4[22]), .A3(n21), .A4(
        sram_rdata_e4[22]), .A5(sram_rdata_d4[22]), .A6(n3), .Y(n_src_box[22])
         );
  AO222X1_HVT U148 ( .A1(n9), .A2(sram_rdata_c4[23]), .A3(n18), .A4(
        sram_rdata_e4[23]), .A5(sram_rdata_d4[23]), .A6(n42), .Y(n_src_box[23]) );
  AO222X1_HVT U149 ( .A1(n10), .A2(sram_rdata_c4[24]), .A3(n24), .A4(
        sram_rdata_e4[24]), .A5(sram_rdata_d4[24]), .A6(n37), .Y(n_src_box[24]) );
  AO222X1_HVT U150 ( .A1(n11), .A2(sram_rdata_c4[27]), .A3(n31), .A4(
        sram_rdata_e4[27]), .A5(sram_rdata_d4[27]), .A6(n42), .Y(n_src_box[27]) );
  AO222X1_HVT U151 ( .A1(n15), .A2(sram_rdata_c4[28]), .A3(n31), .A4(
        sram_rdata_e4[28]), .A5(sram_rdata_d4[28]), .A6(n38), .Y(n_src_box[28]) );
  AO222X1_HVT U152 ( .A1(n36), .A2(sram_rdata_c4[29]), .A3(n19), .A4(
        sram_rdata_e4[29]), .A5(sram_rdata_d4[29]), .A6(n3), .Y(n_src_box[29])
         );
  AO222X1_HVT U153 ( .A1(n34), .A2(sram_rdata_c4[2]), .A3(n23), .A4(
        sram_rdata_e4[2]), .A5(sram_rdata_d4[2]), .A6(n2), .Y(n_src_box[2]) );
  AO222X1_HVT U154 ( .A1(n34), .A2(sram_rdata_c4[30]), .A3(n21), .A4(
        sram_rdata_e4[30]), .A5(sram_rdata_d4[30]), .A6(n8), .Y(n_src_box[30])
         );
  AO222X1_HVT U155 ( .A1(n44), .A2(sram_rdata_c4[31]), .A3(n19), .A4(
        sram_rdata_e4[31]), .A5(sram_rdata_d4[31]), .A6(n2), .Y(n_src_box[31])
         );
  AO222X1_HVT U156 ( .A1(n36), .A2(sram_rdata_c3[3]), .A3(n17), .A4(
        sram_rdata_e3[3]), .A5(sram_rdata_d3[3]), .A6(n2), .Y(n_src_box[35])
         );
  AO222X1_HVT U157 ( .A1(n11), .A2(sram_rdata_c3[4]), .A3(n16), .A4(
        sram_rdata_e3[4]), .A5(sram_rdata_d3[4]), .A6(n39), .Y(n_src_box[36])
         );
  AO222X1_HVT U158 ( .A1(n14), .A2(sram_rdata_c3[5]), .A3(n31), .A4(
        sram_rdata_e3[5]), .A5(sram_rdata_d3[5]), .A6(n37), .Y(n_src_box[37])
         );
  AO222X1_HVT U159 ( .A1(n14), .A2(sram_rdata_c3[6]), .A3(n18), .A4(
        sram_rdata_e3[6]), .A5(sram_rdata_d3[6]), .A6(n39), .Y(n_src_box[38])
         );
  AO222X1_HVT U160 ( .A1(n35), .A2(sram_rdata_c3[7]), .A3(n30), .A4(
        sram_rdata_e3[7]), .A5(sram_rdata_d3[7]), .A6(n37), .Y(n_src_box[39])
         );
  AO222X1_HVT U161 ( .A1(n34), .A2(sram_rdata_c4[3]), .A3(n16), .A4(
        sram_rdata_e4[3]), .A5(sram_rdata_d4[3]), .A6(n39), .Y(n_src_box[3])
         );
  AO222X1_HVT U162 ( .A1(n10), .A2(sram_rdata_c3[10]), .A3(n24), .A4(
        sram_rdata_e3[10]), .A5(sram_rdata_d3[10]), .A6(n6), .Y(n_src_box[42])
         );
  AO222X1_HVT U163 ( .A1(n44), .A2(sram_rdata_c3[11]), .A3(n16), .A4(
        sram_rdata_e3[11]), .A5(sram_rdata_d3[11]), .A6(n42), .Y(n_src_box[43]) );
  AO222X1_HVT U164 ( .A1(n10), .A2(sram_rdata_c3[12]), .A3(n24), .A4(
        sram_rdata_e3[12]), .A5(sram_rdata_d3[12]), .A6(n3), .Y(n_src_box[44])
         );
  AO222X1_HVT U165 ( .A1(n34), .A2(sram_rdata_c3[13]), .A3(n32), .A4(
        sram_rdata_e3[13]), .A5(sram_rdata_d3[13]), .A6(n37), .Y(n_src_box[45]) );
  AO222X1_HVT U166 ( .A1(n15), .A2(sram_rdata_c3[14]), .A3(n31), .A4(
        sram_rdata_e3[14]), .A5(sram_rdata_d3[14]), .A6(n42), .Y(n_src_box[46]) );
  AO222X1_HVT U167 ( .A1(n13), .A2(sram_rdata_c3[15]), .A3(n21), .A4(
        sram_rdata_e3[15]), .A5(sram_rdata_d3[15]), .A6(n37), .Y(n_src_box[47]) );
  AO222X1_HVT U168 ( .A1(n35), .A2(sram_rdata_c4[4]), .A3(n30), .A4(
        sram_rdata_e4[4]), .A5(sram_rdata_d4[4]), .A6(n7), .Y(n_src_box[4]) );
  AO222X1_HVT U169 ( .A1(n36), .A2(sram_rdata_c3[18]), .A3(n22), .A4(
        sram_rdata_e3[18]), .A5(sram_rdata_d3[18]), .A6(n42), .Y(n_src_box[50]) );
  AO222X1_HVT U170 ( .A1(n44), .A2(sram_rdata_c3[19]), .A3(n19), .A4(
        sram_rdata_e3[19]), .A5(sram_rdata_d3[19]), .A6(n7), .Y(n_src_box[51])
         );
  AO222X1_HVT U171 ( .A1(n13), .A2(sram_rdata_c3[20]), .A3(n22), .A4(
        sram_rdata_e3[20]), .A5(sram_rdata_d3[20]), .A6(n5), .Y(n_src_box[52])
         );
  AO222X1_HVT U172 ( .A1(n11), .A2(sram_rdata_c3[21]), .A3(n24), .A4(
        sram_rdata_e3[21]), .A5(sram_rdata_d3[21]), .A6(n3), .Y(n_src_box[53])
         );
  AO222X1_HVT U173 ( .A1(n9), .A2(sram_rdata_c3[22]), .A3(n32), .A4(
        sram_rdata_e3[22]), .A5(sram_rdata_d3[22]), .A6(n7), .Y(n_src_box[54])
         );
  AO222X1_HVT U174 ( .A1(n9), .A2(sram_rdata_c3[23]), .A3(n17), .A4(
        sram_rdata_e3[23]), .A5(sram_rdata_d3[23]), .A6(n39), .Y(n_src_box[55]) );
  AO222X1_HVT U175 ( .A1(n14), .A2(sram_rdata_c3[26]), .A3(n19), .A4(
        sram_rdata_e3[26]), .A5(sram_rdata_d3[26]), .A6(n38), .Y(n_src_box[58]) );
  AO222X1_HVT U176 ( .A1(n35), .A2(sram_rdata_c3[27]), .A3(n32), .A4(
        sram_rdata_e3[27]), .A5(sram_rdata_d3[27]), .A6(n3), .Y(n_src_box[59])
         );
  AO222X1_HVT U177 ( .A1(n34), .A2(sram_rdata_c4[5]), .A3(n17), .A4(
        sram_rdata_e4[5]), .A5(sram_rdata_d4[5]), .A6(n38), .Y(n_src_box[5])
         );
  AO222X1_HVT U178 ( .A1(n15), .A2(sram_rdata_c3[28]), .A3(n32), .A4(
        sram_rdata_e3[28]), .A5(sram_rdata_d3[28]), .A6(n38), .Y(n_src_box[60]) );
  AO222X1_HVT U179 ( .A1(n44), .A2(sram_rdata_c3[29]), .A3(n23), .A4(
        sram_rdata_e3[29]), .A5(sram_rdata_d3[29]), .A6(n39), .Y(n_src_box[61]) );
  AO222X1_HVT U180 ( .A1(n36), .A2(sram_rdata_c3[30]), .A3(n30), .A4(
        sram_rdata_e3[30]), .A5(sram_rdata_d3[30]), .A6(n2), .Y(n_src_box[62])
         );
  AO222X1_HVT U181 ( .A1(n10), .A2(sram_rdata_c3[31]), .A3(n31), .A4(
        sram_rdata_e3[31]), .A5(sram_rdata_d3[31]), .A6(n38), .Y(n_src_box[63]) );
  AO222X1_HVT U182 ( .A1(n13), .A2(sram_rdata_c2[3]), .A3(n18), .A4(
        sram_rdata_e2[3]), .A5(sram_rdata_d2[3]), .A6(n7), .Y(n_src_box[67])
         );
  AO222X1_HVT U183 ( .A1(n12), .A2(sram_rdata_c2[4]), .A3(n31), .A4(
        sram_rdata_e2[4]), .A5(sram_rdata_d2[4]), .A6(n3), .Y(n_src_box[68])
         );
  AO222X1_HVT U184 ( .A1(n36), .A2(sram_rdata_c2[5]), .A3(n17), .A4(
        sram_rdata_e2[5]), .A5(sram_rdata_d2[5]), .A6(n7), .Y(n_src_box[69])
         );
  AO222X1_HVT U185 ( .A1(n34), .A2(sram_rdata_c4[6]), .A3(n32), .A4(
        sram_rdata_e4[6]), .A5(sram_rdata_d4[6]), .A6(n8), .Y(n_src_box[6]) );
  AO222X1_HVT U186 ( .A1(n11), .A2(sram_rdata_c2[6]), .A3(n21), .A4(
        sram_rdata_e2[6]), .A5(sram_rdata_d2[6]), .A6(n38), .Y(n_src_box[70])
         );
  AO222X1_HVT U187 ( .A1(n44), .A2(sram_rdata_c2[7]), .A3(n23), .A4(
        sram_rdata_e2[7]), .A5(sram_rdata_d2[7]), .A6(n7), .Y(n_src_box[71])
         );
  AO222X1_HVT U188 ( .A1(n9), .A2(sram_rdata_c2[10]), .A3(n32), .A4(
        sram_rdata_e2[10]), .A5(sram_rdata_d2[10]), .A6(n8), .Y(n_src_box[74])
         );
  AO222X1_HVT U189 ( .A1(n34), .A2(sram_rdata_c2[11]), .A3(n16), .A4(
        sram_rdata_e2[11]), .A5(sram_rdata_d2[11]), .A6(n2), .Y(n_src_box[75])
         );
  AO222X1_HVT U190 ( .A1(n14), .A2(sram_rdata_c2[12]), .A3(n18), .A4(
        sram_rdata_e2[12]), .A5(sram_rdata_d2[12]), .A6(n8), .Y(n_src_box[76])
         );
  AO222X1_HVT U191 ( .A1(n12), .A2(sram_rdata_c2[13]), .A3(n18), .A4(
        sram_rdata_e2[13]), .A5(sram_rdata_d2[13]), .A6(n2), .Y(n_src_box[77])
         );
  AO222X1_HVT U192 ( .A1(n35), .A2(sram_rdata_c2[14]), .A3(n21), .A4(
        sram_rdata_e2[14]), .A5(sram_rdata_d2[14]), .A6(n2), .Y(n_src_box[78])
         );
  AO222X1_HVT U193 ( .A1(n35), .A2(sram_rdata_c2[15]), .A3(n32), .A4(
        sram_rdata_e2[15]), .A5(sram_rdata_d2[15]), .A6(n5), .Y(n_src_box[79])
         );
  AO222X1_HVT U194 ( .A1(n44), .A2(sram_rdata_c4[7]), .A3(n23), .A4(
        sram_rdata_e4[7]), .A5(sram_rdata_d4[7]), .A6(n38), .Y(n_src_box[7])
         );
  AO222X1_HVT U195 ( .A1(n15), .A2(sram_rdata_c2[18]), .A3(n31), .A4(
        sram_rdata_e2[18]), .A5(sram_rdata_d2[18]), .A6(n37), .Y(n_src_box[82]) );
  AO222X1_HVT U196 ( .A1(n10), .A2(sram_rdata_c2[19]), .A3(n21), .A4(
        sram_rdata_e2[19]), .A5(sram_rdata_d2[19]), .A6(n37), .Y(n_src_box[83]) );
  AO222X1_HVT U197 ( .A1(n9), .A2(sram_rdata_c2[20]), .A3(n21), .A4(
        sram_rdata_e2[20]), .A5(sram_rdata_d2[20]), .A6(n39), .Y(n_src_box[84]) );
  AO222X1_HVT U198 ( .A1(n11), .A2(sram_rdata_c2[21]), .A3(n32), .A4(
        sram_rdata_e2[21]), .A5(sram_rdata_d2[21]), .A6(n37), .Y(n_src_box[85]) );
  AO222X1_HVT U199 ( .A1(n13), .A2(sram_rdata_c2[22]), .A3(n32), .A4(
        sram_rdata_e2[22]), .A5(sram_rdata_d2[22]), .A6(n8), .Y(n_src_box[86])
         );
  AO222X1_HVT U200 ( .A1(n36), .A2(sram_rdata_c2[23]), .A3(n30), .A4(
        sram_rdata_e2[23]), .A5(sram_rdata_d2[23]), .A6(n8), .Y(n_src_box[87])
         );
  AO222X1_HVT U201 ( .A1(n34), .A2(sram_rdata_c2[26]), .A3(n24), .A4(
        sram_rdata_e2[26]), .A5(sram_rdata_d2[26]), .A6(n8), .Y(n_src_box[90])
         );
  AO222X1_HVT U202 ( .A1(n44), .A2(sram_rdata_c2[27]), .A3(n22), .A4(
        sram_rdata_e2[27]), .A5(sram_rdata_d2[27]), .A6(n38), .Y(n_src_box[91]) );
  AO222X1_HVT U203 ( .A1(n44), .A2(sram_rdata_c2[28]), .A3(n31), .A4(
        sram_rdata_e2[28]), .A5(sram_rdata_d2[28]), .A6(n39), .Y(n_src_box[92]) );
  AO222X1_HVT U204 ( .A1(n36), .A2(sram_rdata_c2[29]), .A3(n16), .A4(
        sram_rdata_e2[29]), .A5(sram_rdata_d2[29]), .A6(n7), .Y(n_src_box[93])
         );
  AO222X1_HVT U205 ( .A1(n9), .A2(sram_rdata_c2[30]), .A3(n17), .A4(
        sram_rdata_e2[30]), .A5(sram_rdata_d2[30]), .A6(n42), .Y(n_src_box[94]) );
  AO222X1_HVT U206 ( .A1(n12), .A2(sram_rdata_c2[31]), .A3(n18), .A4(
        sram_rdata_e2[31]), .A5(sram_rdata_d2[31]), .A6(n38), .Y(n_src_box[95]) );
  AO222X1_HVT U207 ( .A1(n14), .A2(sram_rdata_c1[3]), .A3(n19), .A4(
        sram_rdata_e1[3]), .A5(sram_rdata_d1[3]), .A6(n39), .Y(n_src_box[99])
         );
endmodule


module fc_multiplier_accumulator ( clk, srstn, src_window, sram_rdata_weight, 
        accumulate_reset, data_out );
  input [159:0] src_window;
  input [79:0] sram_rdata_weight;
  output [22:0] data_out;
  input clk, srstn, accumulate_reset;
  wire   DP_OP_102J5_124_3590_n2362, DP_OP_102J5_124_3590_n2330,
         DP_OP_102J5_124_3590_n2329, DP_OP_102J5_124_3590_n2328,
         DP_OP_102J5_124_3590_n2327, DP_OP_102J5_124_3590_n2326,
         DP_OP_102J5_124_3590_n2325, DP_OP_102J5_124_3590_n2324,
         DP_OP_102J5_124_3590_n2323, DP_OP_102J5_124_3590_n2322,
         DP_OP_102J5_124_3590_n2321, DP_OP_102J5_124_3590_n2320,
         DP_OP_102J5_124_3590_n2319, DP_OP_102J5_124_3590_n2318,
         DP_OP_102J5_124_3590_n2317, DP_OP_102J5_124_3590_n2316,
         DP_OP_102J5_124_3590_n2315, DP_OP_102J5_124_3590_n2314,
         DP_OP_102J5_124_3590_n2313, DP_OP_102J5_124_3590_n2312,
         DP_OP_102J5_124_3590_n2311, DP_OP_102J5_124_3590_n2310,
         DP_OP_102J5_124_3590_n2309, DP_OP_102J5_124_3590_n2308,
         DP_OP_102J5_124_3590_n2307, DP_OP_102J5_124_3590_n2306,
         DP_OP_102J5_124_3590_n2305, DP_OP_102J5_124_3590_n2304,
         DP_OP_102J5_124_3590_n2303, DP_OP_102J5_124_3590_n2302,
         DP_OP_102J5_124_3590_n2301, DP_OP_102J5_124_3590_n2300,
         DP_OP_102J5_124_3590_n2299, DP_OP_102J5_124_3590_n2298,
         DP_OP_102J5_124_3590_n2297, DP_OP_102J5_124_3590_n2296,
         DP_OP_102J5_124_3590_n2295, DP_OP_102J5_124_3590_n2294,
         DP_OP_102J5_124_3590_n2293, DP_OP_102J5_124_3590_n2292,
         DP_OP_102J5_124_3590_n2287, DP_OP_102J5_124_3590_n2286,
         DP_OP_102J5_124_3590_n2285, DP_OP_102J5_124_3590_n2284,
         DP_OP_102J5_124_3590_n2283, DP_OP_102J5_124_3590_n2282,
         DP_OP_102J5_124_3590_n2281, DP_OP_102J5_124_3590_n2280,
         DP_OP_102J5_124_3590_n2279, DP_OP_102J5_124_3590_n2278,
         DP_OP_102J5_124_3590_n2277, DP_OP_102J5_124_3590_n2276,
         DP_OP_102J5_124_3590_n2275, DP_OP_102J5_124_3590_n2274,
         DP_OP_102J5_124_3590_n2273, DP_OP_102J5_124_3590_n2272,
         DP_OP_102J5_124_3590_n2271, DP_OP_102J5_124_3590_n2270,
         DP_OP_102J5_124_3590_n2269, DP_OP_102J5_124_3590_n2268,
         DP_OP_102J5_124_3590_n2267, DP_OP_102J5_124_3590_n2266,
         DP_OP_102J5_124_3590_n2265, DP_OP_102J5_124_3590_n2264,
         DP_OP_102J5_124_3590_n2263, DP_OP_102J5_124_3590_n2262,
         DP_OP_102J5_124_3590_n2261, DP_OP_102J5_124_3590_n2260,
         DP_OP_102J5_124_3590_n2259, DP_OP_102J5_124_3590_n2258,
         DP_OP_102J5_124_3590_n2257, DP_OP_102J5_124_3590_n2256,
         DP_OP_102J5_124_3590_n2255, DP_OP_102J5_124_3590_n2254,
         DP_OP_102J5_124_3590_n2253, DP_OP_102J5_124_3590_n2252,
         DP_OP_102J5_124_3590_n2251, DP_OP_102J5_124_3590_n2250,
         DP_OP_102J5_124_3590_n2249, DP_OP_102J5_124_3590_n2248,
         DP_OP_102J5_124_3590_n2243, DP_OP_102J5_124_3590_n2242,
         DP_OP_102J5_124_3590_n2241, DP_OP_102J5_124_3590_n2240,
         DP_OP_102J5_124_3590_n2239, DP_OP_102J5_124_3590_n2238,
         DP_OP_102J5_124_3590_n2237, DP_OP_102J5_124_3590_n2236,
         DP_OP_102J5_124_3590_n2235, DP_OP_102J5_124_3590_n2234,
         DP_OP_102J5_124_3590_n2233, DP_OP_102J5_124_3590_n2232,
         DP_OP_102J5_124_3590_n2231, DP_OP_102J5_124_3590_n2230,
         DP_OP_102J5_124_3590_n2229, DP_OP_102J5_124_3590_n2228,
         DP_OP_102J5_124_3590_n2227, DP_OP_102J5_124_3590_n2226,
         DP_OP_102J5_124_3590_n2225, DP_OP_102J5_124_3590_n2224,
         DP_OP_102J5_124_3590_n2223, DP_OP_102J5_124_3590_n2222,
         DP_OP_102J5_124_3590_n2221, DP_OP_102J5_124_3590_n2220,
         DP_OP_102J5_124_3590_n2219, DP_OP_102J5_124_3590_n2218,
         DP_OP_102J5_124_3590_n2217, DP_OP_102J5_124_3590_n2216,
         DP_OP_102J5_124_3590_n2215, DP_OP_102J5_124_3590_n2214,
         DP_OP_102J5_124_3590_n2213, DP_OP_102J5_124_3590_n2212,
         DP_OP_102J5_124_3590_n2211, DP_OP_102J5_124_3590_n2210,
         DP_OP_102J5_124_3590_n2209, DP_OP_102J5_124_3590_n2208,
         DP_OP_102J5_124_3590_n2207, DP_OP_102J5_124_3590_n2206,
         DP_OP_102J5_124_3590_n2205, DP_OP_102J5_124_3590_n2204,
         DP_OP_102J5_124_3590_n2199, DP_OP_102J5_124_3590_n2198,
         DP_OP_102J5_124_3590_n2197, DP_OP_102J5_124_3590_n2196,
         DP_OP_102J5_124_3590_n2195, DP_OP_102J5_124_3590_n2194,
         DP_OP_102J5_124_3590_n2193, DP_OP_102J5_124_3590_n2192,
         DP_OP_102J5_124_3590_n2191, DP_OP_102J5_124_3590_n2190,
         DP_OP_102J5_124_3590_n2189, DP_OP_102J5_124_3590_n2188,
         DP_OP_102J5_124_3590_n2187, DP_OP_102J5_124_3590_n2186,
         DP_OP_102J5_124_3590_n2185, DP_OP_102J5_124_3590_n2184,
         DP_OP_102J5_124_3590_n2183, DP_OP_102J5_124_3590_n2182,
         DP_OP_102J5_124_3590_n2181, DP_OP_102J5_124_3590_n2180,
         DP_OP_102J5_124_3590_n2179, DP_OP_102J5_124_3590_n2178,
         DP_OP_102J5_124_3590_n2177, DP_OP_102J5_124_3590_n2176,
         DP_OP_102J5_124_3590_n2175, DP_OP_102J5_124_3590_n2174,
         DP_OP_102J5_124_3590_n2173, DP_OP_102J5_124_3590_n2172,
         DP_OP_102J5_124_3590_n2171, DP_OP_102J5_124_3590_n2170,
         DP_OP_102J5_124_3590_n2169, DP_OP_102J5_124_3590_n2168,
         DP_OP_102J5_124_3590_n2167, DP_OP_102J5_124_3590_n2166,
         DP_OP_102J5_124_3590_n2165, DP_OP_102J5_124_3590_n2164,
         DP_OP_102J5_124_3590_n2163, DP_OP_102J5_124_3590_n2162,
         DP_OP_102J5_124_3590_n2161, DP_OP_102J5_124_3590_n2160,
         DP_OP_102J5_124_3590_n2155, DP_OP_102J5_124_3590_n2154,
         DP_OP_102J5_124_3590_n2153, DP_OP_102J5_124_3590_n2152,
         DP_OP_102J5_124_3590_n2151, DP_OP_102J5_124_3590_n2150,
         DP_OP_102J5_124_3590_n2149, DP_OP_102J5_124_3590_n2148,
         DP_OP_102J5_124_3590_n2147, DP_OP_102J5_124_3590_n2146,
         DP_OP_102J5_124_3590_n2145, DP_OP_102J5_124_3590_n2144,
         DP_OP_102J5_124_3590_n2143, DP_OP_102J5_124_3590_n2142,
         DP_OP_102J5_124_3590_n2141, DP_OP_102J5_124_3590_n2140,
         DP_OP_102J5_124_3590_n2139, DP_OP_102J5_124_3590_n2138,
         DP_OP_102J5_124_3590_n2137, DP_OP_102J5_124_3590_n2136,
         DP_OP_102J5_124_3590_n2135, DP_OP_102J5_124_3590_n2134,
         DP_OP_102J5_124_3590_n2133, DP_OP_102J5_124_3590_n2132,
         DP_OP_102J5_124_3590_n2131, DP_OP_102J5_124_3590_n2130,
         DP_OP_102J5_124_3590_n2129, DP_OP_102J5_124_3590_n2128,
         DP_OP_102J5_124_3590_n2127, DP_OP_102J5_124_3590_n2126,
         DP_OP_102J5_124_3590_n2125, DP_OP_102J5_124_3590_n2124,
         DP_OP_102J5_124_3590_n2123, DP_OP_102J5_124_3590_n2122,
         DP_OP_102J5_124_3590_n2121, DP_OP_102J5_124_3590_n2120,
         DP_OP_102J5_124_3590_n2119, DP_OP_102J5_124_3590_n2118,
         DP_OP_102J5_124_3590_n2117, DP_OP_102J5_124_3590_n2116,
         DP_OP_102J5_124_3590_n2111, DP_OP_102J5_124_3590_n2110,
         DP_OP_102J5_124_3590_n2109, DP_OP_102J5_124_3590_n2108,
         DP_OP_102J5_124_3590_n2107, DP_OP_102J5_124_3590_n2106,
         DP_OP_102J5_124_3590_n2105, DP_OP_102J5_124_3590_n2104,
         DP_OP_102J5_124_3590_n2103, DP_OP_102J5_124_3590_n2102,
         DP_OP_102J5_124_3590_n2101, DP_OP_102J5_124_3590_n2100,
         DP_OP_102J5_124_3590_n2099, DP_OP_102J5_124_3590_n2098,
         DP_OP_102J5_124_3590_n2097, DP_OP_102J5_124_3590_n2096,
         DP_OP_102J5_124_3590_n2095, DP_OP_102J5_124_3590_n2094,
         DP_OP_102J5_124_3590_n2093, DP_OP_102J5_124_3590_n2092,
         DP_OP_102J5_124_3590_n2091, DP_OP_102J5_124_3590_n2090,
         DP_OP_102J5_124_3590_n2089, DP_OP_102J5_124_3590_n2088,
         DP_OP_102J5_124_3590_n2087, DP_OP_102J5_124_3590_n2086,
         DP_OP_102J5_124_3590_n2085, DP_OP_102J5_124_3590_n2084,
         DP_OP_102J5_124_3590_n2083, DP_OP_102J5_124_3590_n2082,
         DP_OP_102J5_124_3590_n2081, DP_OP_102J5_124_3590_n2080,
         DP_OP_102J5_124_3590_n2079, DP_OP_102J5_124_3590_n2078,
         DP_OP_102J5_124_3590_n2077, DP_OP_102J5_124_3590_n2076,
         DP_OP_102J5_124_3590_n2075, DP_OP_102J5_124_3590_n2074,
         DP_OP_102J5_124_3590_n2073, DP_OP_102J5_124_3590_n2072,
         DP_OP_102J5_124_3590_n2067, DP_OP_102J5_124_3590_n2066,
         DP_OP_102J5_124_3590_n2065, DP_OP_102J5_124_3590_n2064,
         DP_OP_102J5_124_3590_n2063, DP_OP_102J5_124_3590_n2062,
         DP_OP_102J5_124_3590_n2061, DP_OP_102J5_124_3590_n2060,
         DP_OP_102J5_124_3590_n2059, DP_OP_102J5_124_3590_n2058,
         DP_OP_102J5_124_3590_n2057, DP_OP_102J5_124_3590_n2056,
         DP_OP_102J5_124_3590_n2055, DP_OP_102J5_124_3590_n2054,
         DP_OP_102J5_124_3590_n2053, DP_OP_102J5_124_3590_n2052,
         DP_OP_102J5_124_3590_n2051, DP_OP_102J5_124_3590_n2050,
         DP_OP_102J5_124_3590_n2049, DP_OP_102J5_124_3590_n2048,
         DP_OP_102J5_124_3590_n2047, DP_OP_102J5_124_3590_n2046,
         DP_OP_102J5_124_3590_n2045, DP_OP_102J5_124_3590_n2044,
         DP_OP_102J5_124_3590_n2043, DP_OP_102J5_124_3590_n2042,
         DP_OP_102J5_124_3590_n2041, DP_OP_102J5_124_3590_n2040,
         DP_OP_102J5_124_3590_n2039, DP_OP_102J5_124_3590_n2038,
         DP_OP_102J5_124_3590_n2037, DP_OP_102J5_124_3590_n2036,
         DP_OP_102J5_124_3590_n2035, DP_OP_102J5_124_3590_n2034,
         DP_OP_102J5_124_3590_n2033, DP_OP_102J5_124_3590_n2032,
         DP_OP_102J5_124_3590_n2031, DP_OP_102J5_124_3590_n2030,
         DP_OP_102J5_124_3590_n2029, DP_OP_102J5_124_3590_n2028,
         DP_OP_102J5_124_3590_n2023, DP_OP_102J5_124_3590_n2022,
         DP_OP_102J5_124_3590_n2021, DP_OP_102J5_124_3590_n2020,
         DP_OP_102J5_124_3590_n2019, DP_OP_102J5_124_3590_n2018,
         DP_OP_102J5_124_3590_n2017, DP_OP_102J5_124_3590_n2016,
         DP_OP_102J5_124_3590_n2015, DP_OP_102J5_124_3590_n2014,
         DP_OP_102J5_124_3590_n2013, DP_OP_102J5_124_3590_n2012,
         DP_OP_102J5_124_3590_n2011, DP_OP_102J5_124_3590_n2010,
         DP_OP_102J5_124_3590_n2009, DP_OP_102J5_124_3590_n2008,
         DP_OP_102J5_124_3590_n2007, DP_OP_102J5_124_3590_n2006,
         DP_OP_102J5_124_3590_n2005, DP_OP_102J5_124_3590_n2004,
         DP_OP_102J5_124_3590_n2003, DP_OP_102J5_124_3590_n2002,
         DP_OP_102J5_124_3590_n2001, DP_OP_102J5_124_3590_n2000,
         DP_OP_102J5_124_3590_n1999, DP_OP_102J5_124_3590_n1998,
         DP_OP_102J5_124_3590_n1997, DP_OP_102J5_124_3590_n1996,
         DP_OP_102J5_124_3590_n1995, DP_OP_102J5_124_3590_n1994,
         DP_OP_102J5_124_3590_n1993, DP_OP_102J5_124_3590_n1992,
         DP_OP_102J5_124_3590_n1991, DP_OP_102J5_124_3590_n1990,
         DP_OP_102J5_124_3590_n1989, DP_OP_102J5_124_3590_n1988,
         DP_OP_102J5_124_3590_n1987, DP_OP_102J5_124_3590_n1986,
         DP_OP_102J5_124_3590_n1985, DP_OP_102J5_124_3590_n1984,
         DP_OP_102J5_124_3590_n1979, DP_OP_102J5_124_3590_n1978,
         DP_OP_102J5_124_3590_n1977, DP_OP_102J5_124_3590_n1976,
         DP_OP_102J5_124_3590_n1975, DP_OP_102J5_124_3590_n1974,
         DP_OP_102J5_124_3590_n1973, DP_OP_102J5_124_3590_n1972,
         DP_OP_102J5_124_3590_n1971, DP_OP_102J5_124_3590_n1970,
         DP_OP_102J5_124_3590_n1969, DP_OP_102J5_124_3590_n1968,
         DP_OP_102J5_124_3590_n1967, DP_OP_102J5_124_3590_n1966,
         DP_OP_102J5_124_3590_n1965, DP_OP_102J5_124_3590_n1964,
         DP_OP_102J5_124_3590_n1963, DP_OP_102J5_124_3590_n1962,
         DP_OP_102J5_124_3590_n1961, DP_OP_102J5_124_3590_n1960,
         DP_OP_102J5_124_3590_n1959, DP_OP_102J5_124_3590_n1958,
         DP_OP_102J5_124_3590_n1957, DP_OP_102J5_124_3590_n1956,
         DP_OP_102J5_124_3590_n1955, DP_OP_102J5_124_3590_n1954,
         DP_OP_102J5_124_3590_n1953, DP_OP_102J5_124_3590_n1952,
         DP_OP_102J5_124_3590_n1951, DP_OP_102J5_124_3590_n1950,
         DP_OP_102J5_124_3590_n1949, DP_OP_102J5_124_3590_n1948,
         DP_OP_102J5_124_3590_n1947, DP_OP_102J5_124_3590_n1946,
         DP_OP_102J5_124_3590_n1945, DP_OP_102J5_124_3590_n1944,
         DP_OP_102J5_124_3590_n1943, DP_OP_102J5_124_3590_n1942,
         DP_OP_102J5_124_3590_n1941, DP_OP_102J5_124_3590_n1940,
         DP_OP_102J5_124_3590_n1935, DP_OP_102J5_124_3590_n1934,
         DP_OP_102J5_124_3590_n1933, DP_OP_102J5_124_3590_n1932,
         DP_OP_102J5_124_3590_n1931, DP_OP_102J5_124_3590_n1930,
         DP_OP_102J5_124_3590_n1929, DP_OP_102J5_124_3590_n1928,
         DP_OP_102J5_124_3590_n1927, DP_OP_102J5_124_3590_n1926,
         DP_OP_102J5_124_3590_n1925, DP_OP_102J5_124_3590_n1924,
         DP_OP_102J5_124_3590_n1923, DP_OP_102J5_124_3590_n1922,
         DP_OP_102J5_124_3590_n1921, DP_OP_102J5_124_3590_n1920,
         DP_OP_102J5_124_3590_n1919, DP_OP_102J5_124_3590_n1918,
         DP_OP_102J5_124_3590_n1917, DP_OP_102J5_124_3590_n1916,
         DP_OP_102J5_124_3590_n1915, DP_OP_102J5_124_3590_n1914,
         DP_OP_102J5_124_3590_n1913, DP_OP_102J5_124_3590_n1912,
         DP_OP_102J5_124_3590_n1911, DP_OP_102J5_124_3590_n1910,
         DP_OP_102J5_124_3590_n1909, DP_OP_102J5_124_3590_n1908,
         DP_OP_102J5_124_3590_n1907, DP_OP_102J5_124_3590_n1906,
         DP_OP_102J5_124_3590_n1905, DP_OP_102J5_124_3590_n1904,
         DP_OP_102J5_124_3590_n1903, DP_OP_102J5_124_3590_n1902,
         DP_OP_102J5_124_3590_n1901, DP_OP_102J5_124_3590_n1900,
         DP_OP_102J5_124_3590_n1899, DP_OP_102J5_124_3590_n1898,
         DP_OP_102J5_124_3590_n1897, DP_OP_102J5_124_3590_n1896,
         DP_OP_102J5_124_3590_n1891, DP_OP_102J5_124_3590_n1890,
         DP_OP_102J5_124_3590_n1889, DP_OP_102J5_124_3590_n1888,
         DP_OP_102J5_124_3590_n1887, DP_OP_102J5_124_3590_n1886,
         DP_OP_102J5_124_3590_n1885, DP_OP_102J5_124_3590_n1884,
         DP_OP_102J5_124_3590_n1883, DP_OP_102J5_124_3590_n1882,
         DP_OP_102J5_124_3590_n1881, DP_OP_102J5_124_3590_n1880,
         DP_OP_102J5_124_3590_n1879, DP_OP_102J5_124_3590_n1878,
         DP_OP_102J5_124_3590_n1877, DP_OP_102J5_124_3590_n1876,
         DP_OP_102J5_124_3590_n1875, DP_OP_102J5_124_3590_n1874,
         DP_OP_102J5_124_3590_n1873, DP_OP_102J5_124_3590_n1872,
         DP_OP_102J5_124_3590_n1871, DP_OP_102J5_124_3590_n1870,
         DP_OP_102J5_124_3590_n1869, DP_OP_102J5_124_3590_n1868,
         DP_OP_102J5_124_3590_n1867, DP_OP_102J5_124_3590_n1866,
         DP_OP_102J5_124_3590_n1865, DP_OP_102J5_124_3590_n1864,
         DP_OP_102J5_124_3590_n1863, DP_OP_102J5_124_3590_n1862,
         DP_OP_102J5_124_3590_n1861, DP_OP_102J5_124_3590_n1860,
         DP_OP_102J5_124_3590_n1859, DP_OP_102J5_124_3590_n1858,
         DP_OP_102J5_124_3590_n1857, DP_OP_102J5_124_3590_n1856,
         DP_OP_102J5_124_3590_n1855, DP_OP_102J5_124_3590_n1854,
         DP_OP_102J5_124_3590_n1853, DP_OP_102J5_124_3590_n1852,
         DP_OP_102J5_124_3590_n1847, DP_OP_102J5_124_3590_n1846,
         DP_OP_102J5_124_3590_n1845, DP_OP_102J5_124_3590_n1844,
         DP_OP_102J5_124_3590_n1843, DP_OP_102J5_124_3590_n1842,
         DP_OP_102J5_124_3590_n1841, DP_OP_102J5_124_3590_n1840,
         DP_OP_102J5_124_3590_n1839, DP_OP_102J5_124_3590_n1838,
         DP_OP_102J5_124_3590_n1837, DP_OP_102J5_124_3590_n1836,
         DP_OP_102J5_124_3590_n1835, DP_OP_102J5_124_3590_n1834,
         DP_OP_102J5_124_3590_n1833, DP_OP_102J5_124_3590_n1832,
         DP_OP_102J5_124_3590_n1831, DP_OP_102J5_124_3590_n1830,
         DP_OP_102J5_124_3590_n1829, DP_OP_102J5_124_3590_n1828,
         DP_OP_102J5_124_3590_n1827, DP_OP_102J5_124_3590_n1826,
         DP_OP_102J5_124_3590_n1825, DP_OP_102J5_124_3590_n1824,
         DP_OP_102J5_124_3590_n1823, DP_OP_102J5_124_3590_n1822,
         DP_OP_102J5_124_3590_n1821, DP_OP_102J5_124_3590_n1820,
         DP_OP_102J5_124_3590_n1819, DP_OP_102J5_124_3590_n1818,
         DP_OP_102J5_124_3590_n1817, DP_OP_102J5_124_3590_n1816,
         DP_OP_102J5_124_3590_n1815, DP_OP_102J5_124_3590_n1814,
         DP_OP_102J5_124_3590_n1813, DP_OP_102J5_124_3590_n1812,
         DP_OP_102J5_124_3590_n1811, DP_OP_102J5_124_3590_n1810,
         DP_OP_102J5_124_3590_n1809, DP_OP_102J5_124_3590_n1808,
         DP_OP_102J5_124_3590_n1803, DP_OP_102J5_124_3590_n1802,
         DP_OP_102J5_124_3590_n1801, DP_OP_102J5_124_3590_n1800,
         DP_OP_102J5_124_3590_n1799, DP_OP_102J5_124_3590_n1798,
         DP_OP_102J5_124_3590_n1797, DP_OP_102J5_124_3590_n1796,
         DP_OP_102J5_124_3590_n1795, DP_OP_102J5_124_3590_n1794,
         DP_OP_102J5_124_3590_n1793, DP_OP_102J5_124_3590_n1792,
         DP_OP_102J5_124_3590_n1791, DP_OP_102J5_124_3590_n1790,
         DP_OP_102J5_124_3590_n1789, DP_OP_102J5_124_3590_n1788,
         DP_OP_102J5_124_3590_n1787, DP_OP_102J5_124_3590_n1786,
         DP_OP_102J5_124_3590_n1785, DP_OP_102J5_124_3590_n1784,
         DP_OP_102J5_124_3590_n1783, DP_OP_102J5_124_3590_n1782,
         DP_OP_102J5_124_3590_n1781, DP_OP_102J5_124_3590_n1780,
         DP_OP_102J5_124_3590_n1779, DP_OP_102J5_124_3590_n1778,
         DP_OP_102J5_124_3590_n1777, DP_OP_102J5_124_3590_n1776,
         DP_OP_102J5_124_3590_n1775, DP_OP_102J5_124_3590_n1774,
         DP_OP_102J5_124_3590_n1773, DP_OP_102J5_124_3590_n1772,
         DP_OP_102J5_124_3590_n1771, DP_OP_102J5_124_3590_n1770,
         DP_OP_102J5_124_3590_n1769, DP_OP_102J5_124_3590_n1768,
         DP_OP_102J5_124_3590_n1767, DP_OP_102J5_124_3590_n1766,
         DP_OP_102J5_124_3590_n1765, DP_OP_102J5_124_3590_n1760,
         DP_OP_102J5_124_3590_n1759, DP_OP_102J5_124_3590_n1758,
         DP_OP_102J5_124_3590_n1757, DP_OP_102J5_124_3590_n1756,
         DP_OP_102J5_124_3590_n1755, DP_OP_102J5_124_3590_n1754,
         DP_OP_102J5_124_3590_n1753, DP_OP_102J5_124_3590_n1752,
         DP_OP_102J5_124_3590_n1751, DP_OP_102J5_124_3590_n1750,
         DP_OP_102J5_124_3590_n1749, DP_OP_102J5_124_3590_n1748,
         DP_OP_102J5_124_3590_n1747, DP_OP_102J5_124_3590_n1746,
         DP_OP_102J5_124_3590_n1745, DP_OP_102J5_124_3590_n1744,
         DP_OP_102J5_124_3590_n1743, DP_OP_102J5_124_3590_n1742,
         DP_OP_102J5_124_3590_n1741, DP_OP_102J5_124_3590_n1740,
         DP_OP_102J5_124_3590_n1739, DP_OP_102J5_124_3590_n1738,
         DP_OP_102J5_124_3590_n1737, DP_OP_102J5_124_3590_n1736,
         DP_OP_102J5_124_3590_n1735, DP_OP_102J5_124_3590_n1734,
         DP_OP_102J5_124_3590_n1733, DP_OP_102J5_124_3590_n1732,
         DP_OP_102J5_124_3590_n1731, DP_OP_102J5_124_3590_n1730,
         DP_OP_102J5_124_3590_n1729, DP_OP_102J5_124_3590_n1728,
         DP_OP_102J5_124_3590_n1727, DP_OP_102J5_124_3590_n1726,
         DP_OP_102J5_124_3590_n1725, DP_OP_102J5_124_3590_n1724,
         DP_OP_102J5_124_3590_n1723, DP_OP_102J5_124_3590_n1722,
         DP_OP_102J5_124_3590_n1721, DP_OP_102J5_124_3590_n1716,
         DP_OP_102J5_124_3590_n1715, DP_OP_102J5_124_3590_n1714,
         DP_OP_102J5_124_3590_n1713, DP_OP_102J5_124_3590_n1712,
         DP_OP_102J5_124_3590_n1711, DP_OP_102J5_124_3590_n1710,
         DP_OP_102J5_124_3590_n1709, DP_OP_102J5_124_3590_n1708,
         DP_OP_102J5_124_3590_n1707, DP_OP_102J5_124_3590_n1706,
         DP_OP_102J5_124_3590_n1705, DP_OP_102J5_124_3590_n1704,
         DP_OP_102J5_124_3590_n1703, DP_OP_102J5_124_3590_n1702,
         DP_OP_102J5_124_3590_n1701, DP_OP_102J5_124_3590_n1700,
         DP_OP_102J5_124_3590_n1699, DP_OP_102J5_124_3590_n1698,
         DP_OP_102J5_124_3590_n1697, DP_OP_102J5_124_3590_n1696,
         DP_OP_102J5_124_3590_n1695, DP_OP_102J5_124_3590_n1694,
         DP_OP_102J5_124_3590_n1693, DP_OP_102J5_124_3590_n1692,
         DP_OP_102J5_124_3590_n1691, DP_OP_102J5_124_3590_n1690,
         DP_OP_102J5_124_3590_n1689, DP_OP_102J5_124_3590_n1688,
         DP_OP_102J5_124_3590_n1687, DP_OP_102J5_124_3590_n1686,
         DP_OP_102J5_124_3590_n1685, DP_OP_102J5_124_3590_n1684,
         DP_OP_102J5_124_3590_n1683, DP_OP_102J5_124_3590_n1682,
         DP_OP_102J5_124_3590_n1681, DP_OP_102J5_124_3590_n1680,
         DP_OP_102J5_124_3590_n1679, DP_OP_102J5_124_3590_n1678,
         DP_OP_102J5_124_3590_n1677, DP_OP_102J5_124_3590_n1672,
         DP_OP_102J5_124_3590_n1671, DP_OP_102J5_124_3590_n1670,
         DP_OP_102J5_124_3590_n1669, DP_OP_102J5_124_3590_n1668,
         DP_OP_102J5_124_3590_n1667, DP_OP_102J5_124_3590_n1666,
         DP_OP_102J5_124_3590_n1665, DP_OP_102J5_124_3590_n1664,
         DP_OP_102J5_124_3590_n1663, DP_OP_102J5_124_3590_n1662,
         DP_OP_102J5_124_3590_n1661, DP_OP_102J5_124_3590_n1660,
         DP_OP_102J5_124_3590_n1659, DP_OP_102J5_124_3590_n1658,
         DP_OP_102J5_124_3590_n1657, DP_OP_102J5_124_3590_n1656,
         DP_OP_102J5_124_3590_n1655, DP_OP_102J5_124_3590_n1654,
         DP_OP_102J5_124_3590_n1653, DP_OP_102J5_124_3590_n1652,
         DP_OP_102J5_124_3590_n1651, DP_OP_102J5_124_3590_n1650,
         DP_OP_102J5_124_3590_n1649, DP_OP_102J5_124_3590_n1648,
         DP_OP_102J5_124_3590_n1647, DP_OP_102J5_124_3590_n1646,
         DP_OP_102J5_124_3590_n1645, DP_OP_102J5_124_3590_n1644,
         DP_OP_102J5_124_3590_n1643, DP_OP_102J5_124_3590_n1642,
         DP_OP_102J5_124_3590_n1641, DP_OP_102J5_124_3590_n1640,
         DP_OP_102J5_124_3590_n1639, DP_OP_102J5_124_3590_n1638,
         DP_OP_102J5_124_3590_n1637, DP_OP_102J5_124_3590_n1636,
         DP_OP_102J5_124_3590_n1635, DP_OP_102J5_124_3590_n1634,
         DP_OP_102J5_124_3590_n1633, DP_OP_102J5_124_3590_n1628,
         DP_OP_102J5_124_3590_n1627, DP_OP_102J5_124_3590_n1626,
         DP_OP_102J5_124_3590_n1625, DP_OP_102J5_124_3590_n1624,
         DP_OP_102J5_124_3590_n1623, DP_OP_102J5_124_3590_n1622,
         DP_OP_102J5_124_3590_n1621, DP_OP_102J5_124_3590_n1620,
         DP_OP_102J5_124_3590_n1619, DP_OP_102J5_124_3590_n1618,
         DP_OP_102J5_124_3590_n1617, DP_OP_102J5_124_3590_n1616,
         DP_OP_102J5_124_3590_n1615, DP_OP_102J5_124_3590_n1614,
         DP_OP_102J5_124_3590_n1613, DP_OP_102J5_124_3590_n1612,
         DP_OP_102J5_124_3590_n1611, DP_OP_102J5_124_3590_n1610,
         DP_OP_102J5_124_3590_n1609, DP_OP_102J5_124_3590_n1608,
         DP_OP_102J5_124_3590_n1607, DP_OP_102J5_124_3590_n1606,
         DP_OP_102J5_124_3590_n1605, DP_OP_102J5_124_3590_n1604,
         DP_OP_102J5_124_3590_n1603, DP_OP_102J5_124_3590_n1602,
         DP_OP_102J5_124_3590_n1601, DP_OP_102J5_124_3590_n1600,
         DP_OP_102J5_124_3590_n1599, DP_OP_102J5_124_3590_n1598,
         DP_OP_102J5_124_3590_n1597, DP_OP_102J5_124_3590_n1596,
         DP_OP_102J5_124_3590_n1595, DP_OP_102J5_124_3590_n1594,
         DP_OP_102J5_124_3590_n1593, DP_OP_102J5_124_3590_n1592,
         DP_OP_102J5_124_3590_n1591, DP_OP_102J5_124_3590_n1590,
         DP_OP_102J5_124_3590_n1589, DP_OP_102J5_124_3590_n1584,
         DP_OP_102J5_124_3590_n1583, DP_OP_102J5_124_3590_n1582,
         DP_OP_102J5_124_3590_n1581, DP_OP_102J5_124_3590_n1580,
         DP_OP_102J5_124_3590_n1579, DP_OP_102J5_124_3590_n1578,
         DP_OP_102J5_124_3590_n1577, DP_OP_102J5_124_3590_n1576,
         DP_OP_102J5_124_3590_n1575, DP_OP_102J5_124_3590_n1574,
         DP_OP_102J5_124_3590_n1573, DP_OP_102J5_124_3590_n1572,
         DP_OP_102J5_124_3590_n1571, DP_OP_102J5_124_3590_n1570,
         DP_OP_102J5_124_3590_n1569, DP_OP_102J5_124_3590_n1568,
         DP_OP_102J5_124_3590_n1567, DP_OP_102J5_124_3590_n1566,
         DP_OP_102J5_124_3590_n1565, DP_OP_102J5_124_3590_n1564,
         DP_OP_102J5_124_3590_n1563, DP_OP_102J5_124_3590_n1562,
         DP_OP_102J5_124_3590_n1561, DP_OP_102J5_124_3590_n1560,
         DP_OP_102J5_124_3590_n1559, DP_OP_102J5_124_3590_n1558,
         DP_OP_102J5_124_3590_n1557, DP_OP_102J5_124_3590_n1556,
         DP_OP_102J5_124_3590_n1555, DP_OP_102J5_124_3590_n1554,
         DP_OP_102J5_124_3590_n1553, DP_OP_102J5_124_3590_n1552,
         DP_OP_102J5_124_3590_n1551, DP_OP_102J5_124_3590_n1550,
         DP_OP_102J5_124_3590_n1549, DP_OP_102J5_124_3590_n1548,
         DP_OP_102J5_124_3590_n1547, DP_OP_102J5_124_3590_n1546,
         DP_OP_102J5_124_3590_n1545, DP_OP_102J5_124_3590_n1540,
         DP_OP_102J5_124_3590_n1539, DP_OP_102J5_124_3590_n1538,
         DP_OP_102J5_124_3590_n1537, DP_OP_102J5_124_3590_n1536,
         DP_OP_102J5_124_3590_n1535, DP_OP_102J5_124_3590_n1534,
         DP_OP_102J5_124_3590_n1533, DP_OP_102J5_124_3590_n1532,
         DP_OP_102J5_124_3590_n1531, DP_OP_102J5_124_3590_n1530,
         DP_OP_102J5_124_3590_n1529, DP_OP_102J5_124_3590_n1528,
         DP_OP_102J5_124_3590_n1527, DP_OP_102J5_124_3590_n1526,
         DP_OP_102J5_124_3590_n1525, DP_OP_102J5_124_3590_n1524,
         DP_OP_102J5_124_3590_n1523, DP_OP_102J5_124_3590_n1522,
         DP_OP_102J5_124_3590_n1521, DP_OP_102J5_124_3590_n1520,
         DP_OP_102J5_124_3590_n1519, DP_OP_102J5_124_3590_n1518,
         DP_OP_102J5_124_3590_n1517, DP_OP_102J5_124_3590_n1516,
         DP_OP_102J5_124_3590_n1515, DP_OP_102J5_124_3590_n1514,
         DP_OP_102J5_124_3590_n1513, DP_OP_102J5_124_3590_n1512,
         DP_OP_102J5_124_3590_n1511, DP_OP_102J5_124_3590_n1510,
         DP_OP_102J5_124_3590_n1509, DP_OP_102J5_124_3590_n1508,
         DP_OP_102J5_124_3590_n1507, DP_OP_102J5_124_3590_n1506,
         DP_OP_102J5_124_3590_n1505, DP_OP_102J5_124_3590_n1504,
         DP_OP_102J5_124_3590_n1503, DP_OP_102J5_124_3590_n1502,
         DP_OP_102J5_124_3590_n1501, DP_OP_102J5_124_3590_n1496,
         DP_OP_102J5_124_3590_n1495, DP_OP_102J5_124_3590_n1494,
         DP_OP_102J5_124_3590_n1493, DP_OP_102J5_124_3590_n1492,
         DP_OP_102J5_124_3590_n1491, DP_OP_102J5_124_3590_n1490,
         DP_OP_102J5_124_3590_n1489, DP_OP_102J5_124_3590_n1488,
         DP_OP_102J5_124_3590_n1487, DP_OP_102J5_124_3590_n1486,
         DP_OP_102J5_124_3590_n1485, DP_OP_102J5_124_3590_n1484,
         DP_OP_102J5_124_3590_n1483, DP_OP_102J5_124_3590_n1482,
         DP_OP_102J5_124_3590_n1481, DP_OP_102J5_124_3590_n1480,
         DP_OP_102J5_124_3590_n1479, DP_OP_102J5_124_3590_n1478,
         DP_OP_102J5_124_3590_n1477, DP_OP_102J5_124_3590_n1476,
         DP_OP_102J5_124_3590_n1475, DP_OP_102J5_124_3590_n1474,
         DP_OP_102J5_124_3590_n1473, DP_OP_102J5_124_3590_n1472,
         DP_OP_102J5_124_3590_n1471, DP_OP_102J5_124_3590_n1470,
         DP_OP_102J5_124_3590_n1469, DP_OP_102J5_124_3590_n1468,
         DP_OP_102J5_124_3590_n1467, DP_OP_102J5_124_3590_n1466,
         DP_OP_102J5_124_3590_n1465, DP_OP_102J5_124_3590_n1464,
         DP_OP_102J5_124_3590_n1463, DP_OP_102J5_124_3590_n1462,
         DP_OP_102J5_124_3590_n1461, DP_OP_102J5_124_3590_n1460,
         DP_OP_102J5_124_3590_n1459, DP_OP_102J5_124_3590_n1458,
         DP_OP_102J5_124_3590_n1457, DP_OP_102J5_124_3590_n1432,
         DP_OP_102J5_124_3590_n1431, DP_OP_102J5_124_3590_n1430,
         DP_OP_102J5_124_3590_n1429, DP_OP_102J5_124_3590_n1428,
         DP_OP_102J5_124_3590_n1427, DP_OP_102J5_124_3590_n1426,
         DP_OP_102J5_124_3590_n1425, DP_OP_102J5_124_3590_n1424,
         DP_OP_102J5_124_3590_n1423, DP_OP_102J5_124_3590_n1422,
         DP_OP_102J5_124_3590_n1421, DP_OP_102J5_124_3590_n1420,
         DP_OP_102J5_124_3590_n1419, DP_OP_102J5_124_3590_n1417,
         DP_OP_102J5_124_3590_n1416, DP_OP_102J5_124_3590_n1415,
         DP_OP_102J5_124_3590_n1414, DP_OP_102J5_124_3590_n1413,
         DP_OP_102J5_124_3590_n1412, DP_OP_102J5_124_3590_n1411,
         DP_OP_102J5_124_3590_n1410, DP_OP_102J5_124_3590_n1409,
         DP_OP_102J5_124_3590_n1408, DP_OP_102J5_124_3590_n1407,
         DP_OP_102J5_124_3590_n1406, DP_OP_102J5_124_3590_n1405,
         DP_OP_102J5_124_3590_n1404, DP_OP_102J5_124_3590_n1403,
         DP_OP_102J5_124_3590_n1402, DP_OP_102J5_124_3590_n1401,
         DP_OP_102J5_124_3590_n1400, DP_OP_102J5_124_3590_n1399,
         DP_OP_102J5_124_3590_n1398, DP_OP_102J5_124_3590_n1397,
         DP_OP_102J5_124_3590_n1396, DP_OP_102J5_124_3590_n1395,
         DP_OP_102J5_124_3590_n1394, DP_OP_102J5_124_3590_n1393,
         DP_OP_102J5_124_3590_n1392, DP_OP_102J5_124_3590_n1391,
         DP_OP_102J5_124_3590_n1390, DP_OP_102J5_124_3590_n1389,
         DP_OP_102J5_124_3590_n1388, DP_OP_102J5_124_3590_n1387,
         DP_OP_102J5_124_3590_n1386, DP_OP_102J5_124_3590_n1385,
         DP_OP_102J5_124_3590_n1384, DP_OP_102J5_124_3590_n1383,
         DP_OP_102J5_124_3590_n1382, DP_OP_102J5_124_3590_n1381,
         DP_OP_102J5_124_3590_n1380, DP_OP_102J5_124_3590_n1379,
         DP_OP_102J5_124_3590_n1378, DP_OP_102J5_124_3590_n1377,
         DP_OP_102J5_124_3590_n1376, DP_OP_102J5_124_3590_n1375,
         DP_OP_102J5_124_3590_n1374, DP_OP_102J5_124_3590_n1373,
         DP_OP_102J5_124_3590_n1372, DP_OP_102J5_124_3590_n1371,
         DP_OP_102J5_124_3590_n1370, DP_OP_102J5_124_3590_n1369,
         DP_OP_102J5_124_3590_n1368, DP_OP_102J5_124_3590_n1367,
         DP_OP_102J5_124_3590_n1366, DP_OP_102J5_124_3590_n1365,
         DP_OP_102J5_124_3590_n1364, DP_OP_102J5_124_3590_n1363,
         DP_OP_102J5_124_3590_n1362, DP_OP_102J5_124_3590_n1361,
         DP_OP_102J5_124_3590_n1360, DP_OP_102J5_124_3590_n1359,
         DP_OP_102J5_124_3590_n1358, DP_OP_102J5_124_3590_n1357,
         DP_OP_102J5_124_3590_n1356, DP_OP_102J5_124_3590_n1355,
         DP_OP_102J5_124_3590_n1354, DP_OP_102J5_124_3590_n1353,
         DP_OP_102J5_124_3590_n1352, DP_OP_102J5_124_3590_n1351,
         DP_OP_102J5_124_3590_n1350, DP_OP_102J5_124_3590_n1349,
         DP_OP_102J5_124_3590_n1348, DP_OP_102J5_124_3590_n1347,
         DP_OP_102J5_124_3590_n1346, DP_OP_102J5_124_3590_n1345,
         DP_OP_102J5_124_3590_n1344, DP_OP_102J5_124_3590_n1343,
         DP_OP_102J5_124_3590_n1342, DP_OP_102J5_124_3590_n1341,
         DP_OP_102J5_124_3590_n1340, DP_OP_102J5_124_3590_n1339,
         DP_OP_102J5_124_3590_n1338, DP_OP_102J5_124_3590_n1337,
         DP_OP_102J5_124_3590_n1336, DP_OP_102J5_124_3590_n1335,
         DP_OP_102J5_124_3590_n1334, DP_OP_102J5_124_3590_n1333,
         DP_OP_102J5_124_3590_n1332, DP_OP_102J5_124_3590_n1331,
         DP_OP_102J5_124_3590_n1330, DP_OP_102J5_124_3590_n1329,
         DP_OP_102J5_124_3590_n1328, DP_OP_102J5_124_3590_n1327,
         DP_OP_102J5_124_3590_n1326, DP_OP_102J5_124_3590_n1325,
         DP_OP_102J5_124_3590_n1324, DP_OP_102J5_124_3590_n1323,
         DP_OP_102J5_124_3590_n1322, DP_OP_102J5_124_3590_n1321,
         DP_OP_102J5_124_3590_n1320, DP_OP_102J5_124_3590_n1319,
         DP_OP_102J5_124_3590_n1318, DP_OP_102J5_124_3590_n1317,
         DP_OP_102J5_124_3590_n1316, DP_OP_102J5_124_3590_n1315,
         DP_OP_102J5_124_3590_n1314, DP_OP_102J5_124_3590_n1313,
         DP_OP_102J5_124_3590_n1312, DP_OP_102J5_124_3590_n1311,
         DP_OP_102J5_124_3590_n1310, DP_OP_102J5_124_3590_n1309,
         DP_OP_102J5_124_3590_n1308, DP_OP_102J5_124_3590_n1307,
         DP_OP_102J5_124_3590_n1306, DP_OP_102J5_124_3590_n1305,
         DP_OP_102J5_124_3590_n1304, DP_OP_102J5_124_3590_n1303,
         DP_OP_102J5_124_3590_n1302, DP_OP_102J5_124_3590_n1301,
         DP_OP_102J5_124_3590_n1300, DP_OP_102J5_124_3590_n1299,
         DP_OP_102J5_124_3590_n1298, DP_OP_102J5_124_3590_n1297,
         DP_OP_102J5_124_3590_n1296, DP_OP_102J5_124_3590_n1295,
         DP_OP_102J5_124_3590_n1294, DP_OP_102J5_124_3590_n1293,
         DP_OP_102J5_124_3590_n1292, DP_OP_102J5_124_3590_n1291,
         DP_OP_102J5_124_3590_n1290, DP_OP_102J5_124_3590_n1289,
         DP_OP_102J5_124_3590_n1288, DP_OP_102J5_124_3590_n1287,
         DP_OP_102J5_124_3590_n1286, DP_OP_102J5_124_3590_n1285,
         DP_OP_102J5_124_3590_n1284, DP_OP_102J5_124_3590_n1283,
         DP_OP_102J5_124_3590_n1282, DP_OP_102J5_124_3590_n1281,
         DP_OP_102J5_124_3590_n1280, DP_OP_102J5_124_3590_n1279,
         DP_OP_102J5_124_3590_n1278, DP_OP_102J5_124_3590_n1277,
         DP_OP_102J5_124_3590_n1276, DP_OP_102J5_124_3590_n1275,
         DP_OP_102J5_124_3590_n1274, DP_OP_102J5_124_3590_n1273,
         DP_OP_102J5_124_3590_n1272, DP_OP_102J5_124_3590_n1271,
         DP_OP_102J5_124_3590_n1270, DP_OP_102J5_124_3590_n1269,
         DP_OP_102J5_124_3590_n1268, DP_OP_102J5_124_3590_n1267,
         DP_OP_102J5_124_3590_n1266, DP_OP_102J5_124_3590_n1265,
         DP_OP_102J5_124_3590_n1264, DP_OP_102J5_124_3590_n1263,
         DP_OP_102J5_124_3590_n1262, DP_OP_102J5_124_3590_n1261,
         DP_OP_102J5_124_3590_n1260, DP_OP_102J5_124_3590_n1259,
         DP_OP_102J5_124_3590_n1258, DP_OP_102J5_124_3590_n1257,
         DP_OP_102J5_124_3590_n1256, DP_OP_102J5_124_3590_n1255,
         DP_OP_102J5_124_3590_n1254, DP_OP_102J5_124_3590_n1253,
         DP_OP_102J5_124_3590_n1252, DP_OP_102J5_124_3590_n1251,
         DP_OP_102J5_124_3590_n1250, DP_OP_102J5_124_3590_n1249,
         DP_OP_102J5_124_3590_n1248, DP_OP_102J5_124_3590_n1247,
         DP_OP_102J5_124_3590_n1246, DP_OP_102J5_124_3590_n1245,
         DP_OP_102J5_124_3590_n1244, DP_OP_102J5_124_3590_n1243,
         DP_OP_102J5_124_3590_n1242, DP_OP_102J5_124_3590_n1241,
         DP_OP_102J5_124_3590_n1240, DP_OP_102J5_124_3590_n1239,
         DP_OP_102J5_124_3590_n1238, DP_OP_102J5_124_3590_n1237,
         DP_OP_102J5_124_3590_n1236, DP_OP_102J5_124_3590_n1235,
         DP_OP_102J5_124_3590_n1234, DP_OP_102J5_124_3590_n1233,
         DP_OP_102J5_124_3590_n1232, DP_OP_102J5_124_3590_n1231,
         DP_OP_102J5_124_3590_n1230, DP_OP_102J5_124_3590_n1229,
         DP_OP_102J5_124_3590_n1228, DP_OP_102J5_124_3590_n1227,
         DP_OP_102J5_124_3590_n1226, DP_OP_102J5_124_3590_n1225,
         DP_OP_102J5_124_3590_n1224, DP_OP_102J5_124_3590_n1223,
         DP_OP_102J5_124_3590_n1222, DP_OP_102J5_124_3590_n1221,
         DP_OP_102J5_124_3590_n1220, DP_OP_102J5_124_3590_n1219,
         DP_OP_102J5_124_3590_n1218, DP_OP_102J5_124_3590_n1217,
         DP_OP_102J5_124_3590_n1216, DP_OP_102J5_124_3590_n1215,
         DP_OP_102J5_124_3590_n1214, DP_OP_102J5_124_3590_n1213,
         DP_OP_102J5_124_3590_n1212, DP_OP_102J5_124_3590_n1211,
         DP_OP_102J5_124_3590_n1210, DP_OP_102J5_124_3590_n1209,
         DP_OP_102J5_124_3590_n1208, DP_OP_102J5_124_3590_n1207,
         DP_OP_102J5_124_3590_n1206, DP_OP_102J5_124_3590_n1205,
         DP_OP_102J5_124_3590_n1204, DP_OP_102J5_124_3590_n1203,
         DP_OP_102J5_124_3590_n1202, DP_OP_102J5_124_3590_n1201,
         DP_OP_102J5_124_3590_n1200, DP_OP_102J5_124_3590_n1199,
         DP_OP_102J5_124_3590_n1198, DP_OP_102J5_124_3590_n1197,
         DP_OP_102J5_124_3590_n1196, DP_OP_102J5_124_3590_n1195,
         DP_OP_102J5_124_3590_n1194, DP_OP_102J5_124_3590_n1193,
         DP_OP_102J5_124_3590_n1192, DP_OP_102J5_124_3590_n1191,
         DP_OP_102J5_124_3590_n1190, DP_OP_102J5_124_3590_n1189,
         DP_OP_102J5_124_3590_n1188, DP_OP_102J5_124_3590_n1187,
         DP_OP_102J5_124_3590_n1186, DP_OP_102J5_124_3590_n1185,
         DP_OP_102J5_124_3590_n1184, DP_OP_102J5_124_3590_n1183,
         DP_OP_102J5_124_3590_n1182, DP_OP_102J5_124_3590_n1181,
         DP_OP_102J5_124_3590_n1180, DP_OP_102J5_124_3590_n1179,
         DP_OP_102J5_124_3590_n1178, DP_OP_102J5_124_3590_n1177,
         DP_OP_102J5_124_3590_n1176, DP_OP_102J5_124_3590_n1175,
         DP_OP_102J5_124_3590_n1174, DP_OP_102J5_124_3590_n1173,
         DP_OP_102J5_124_3590_n1172, DP_OP_102J5_124_3590_n1171,
         DP_OP_102J5_124_3590_n1170, DP_OP_102J5_124_3590_n1169,
         DP_OP_102J5_124_3590_n1168, DP_OP_102J5_124_3590_n1167,
         DP_OP_102J5_124_3590_n1166, DP_OP_102J5_124_3590_n1165,
         DP_OP_102J5_124_3590_n1164, DP_OP_102J5_124_3590_n1163,
         DP_OP_102J5_124_3590_n1162, DP_OP_102J5_124_3590_n1161,
         DP_OP_102J5_124_3590_n1160, DP_OP_102J5_124_3590_n1159,
         DP_OP_102J5_124_3590_n1158, DP_OP_102J5_124_3590_n1157,
         DP_OP_102J5_124_3590_n1156, DP_OP_102J5_124_3590_n1155,
         DP_OP_102J5_124_3590_n1154, DP_OP_102J5_124_3590_n1153,
         DP_OP_102J5_124_3590_n1152, DP_OP_102J5_124_3590_n1151,
         DP_OP_102J5_124_3590_n1150, DP_OP_102J5_124_3590_n1149,
         DP_OP_102J5_124_3590_n1148, DP_OP_102J5_124_3590_n1147,
         DP_OP_102J5_124_3590_n1146, DP_OP_102J5_124_3590_n1145,
         DP_OP_102J5_124_3590_n1144, DP_OP_102J5_124_3590_n1143,
         DP_OP_102J5_124_3590_n1142, DP_OP_102J5_124_3590_n1141,
         DP_OP_102J5_124_3590_n1140, DP_OP_102J5_124_3590_n1139,
         DP_OP_102J5_124_3590_n1138, DP_OP_102J5_124_3590_n1137,
         DP_OP_102J5_124_3590_n1136, DP_OP_102J5_124_3590_n1135,
         DP_OP_102J5_124_3590_n1134, DP_OP_102J5_124_3590_n1133,
         DP_OP_102J5_124_3590_n1132, DP_OP_102J5_124_3590_n1131,
         DP_OP_102J5_124_3590_n1130, DP_OP_102J5_124_3590_n1129,
         DP_OP_102J5_124_3590_n1128, DP_OP_102J5_124_3590_n1127,
         DP_OP_102J5_124_3590_n1126, DP_OP_102J5_124_3590_n1125,
         DP_OP_102J5_124_3590_n1124, DP_OP_102J5_124_3590_n1123,
         DP_OP_102J5_124_3590_n1122, DP_OP_102J5_124_3590_n1121,
         DP_OP_102J5_124_3590_n1120, DP_OP_102J5_124_3590_n1119,
         DP_OP_102J5_124_3590_n1118, DP_OP_102J5_124_3590_n1117,
         DP_OP_102J5_124_3590_n1116, DP_OP_102J5_124_3590_n1115,
         DP_OP_102J5_124_3590_n1114, DP_OP_102J5_124_3590_n1113,
         DP_OP_102J5_124_3590_n1112, DP_OP_102J5_124_3590_n1111,
         DP_OP_102J5_124_3590_n1110, DP_OP_102J5_124_3590_n1109,
         DP_OP_102J5_124_3590_n1108, DP_OP_102J5_124_3590_n1107,
         DP_OP_102J5_124_3590_n1106, DP_OP_102J5_124_3590_n1105,
         DP_OP_102J5_124_3590_n1104, DP_OP_102J5_124_3590_n1103,
         DP_OP_102J5_124_3590_n1102, DP_OP_102J5_124_3590_n1101,
         DP_OP_102J5_124_3590_n1100, DP_OP_102J5_124_3590_n1099,
         DP_OP_102J5_124_3590_n1098, DP_OP_102J5_124_3590_n1097,
         DP_OP_102J5_124_3590_n1096, DP_OP_102J5_124_3590_n1095,
         DP_OP_102J5_124_3590_n1094, DP_OP_102J5_124_3590_n1093,
         DP_OP_102J5_124_3590_n1092, DP_OP_102J5_124_3590_n1091,
         DP_OP_102J5_124_3590_n1090, DP_OP_102J5_124_3590_n1089,
         DP_OP_102J5_124_3590_n1088, DP_OP_102J5_124_3590_n1087,
         DP_OP_102J5_124_3590_n1086, DP_OP_102J5_124_3590_n1085,
         DP_OP_102J5_124_3590_n1084, DP_OP_102J5_124_3590_n1083,
         DP_OP_102J5_124_3590_n1082, DP_OP_102J5_124_3590_n1081,
         DP_OP_102J5_124_3590_n1080, DP_OP_102J5_124_3590_n1079,
         DP_OP_102J5_124_3590_n1078, DP_OP_102J5_124_3590_n1077,
         DP_OP_102J5_124_3590_n1076, DP_OP_102J5_124_3590_n1075,
         DP_OP_102J5_124_3590_n1074, DP_OP_102J5_124_3590_n1073,
         DP_OP_102J5_124_3590_n1072, DP_OP_102J5_124_3590_n1071,
         DP_OP_102J5_124_3590_n1070, DP_OP_102J5_124_3590_n1069,
         DP_OP_102J5_124_3590_n1068, DP_OP_102J5_124_3590_n1067,
         DP_OP_102J5_124_3590_n1066, DP_OP_102J5_124_3590_n1065,
         DP_OP_102J5_124_3590_n1064, DP_OP_102J5_124_3590_n1063,
         DP_OP_102J5_124_3590_n1062, DP_OP_102J5_124_3590_n1061,
         DP_OP_102J5_124_3590_n1060, DP_OP_102J5_124_3590_n1059,
         DP_OP_102J5_124_3590_n1058, DP_OP_102J5_124_3590_n1057,
         DP_OP_102J5_124_3590_n1056, DP_OP_102J5_124_3590_n1055,
         DP_OP_102J5_124_3590_n1054, DP_OP_102J5_124_3590_n1053,
         DP_OP_102J5_124_3590_n1052, DP_OP_102J5_124_3590_n1051,
         DP_OP_102J5_124_3590_n1050, DP_OP_102J5_124_3590_n1049,
         DP_OP_102J5_124_3590_n1048, DP_OP_102J5_124_3590_n1047,
         DP_OP_102J5_124_3590_n1046, DP_OP_102J5_124_3590_n1045,
         DP_OP_102J5_124_3590_n1044, DP_OP_102J5_124_3590_n1043,
         DP_OP_102J5_124_3590_n1042, DP_OP_102J5_124_3590_n1041,
         DP_OP_102J5_124_3590_n1040, DP_OP_102J5_124_3590_n1039,
         DP_OP_102J5_124_3590_n1038, DP_OP_102J5_124_3590_n1037,
         DP_OP_102J5_124_3590_n1036, DP_OP_102J5_124_3590_n1035,
         DP_OP_102J5_124_3590_n1034, DP_OP_102J5_124_3590_n1033,
         DP_OP_102J5_124_3590_n1032, DP_OP_102J5_124_3590_n1031,
         DP_OP_102J5_124_3590_n1030, DP_OP_102J5_124_3590_n1029,
         DP_OP_102J5_124_3590_n1028, DP_OP_102J5_124_3590_n1027,
         DP_OP_102J5_124_3590_n1026, DP_OP_102J5_124_3590_n1025,
         DP_OP_102J5_124_3590_n1024, DP_OP_102J5_124_3590_n1023,
         DP_OP_102J5_124_3590_n1022, DP_OP_102J5_124_3590_n1021,
         DP_OP_102J5_124_3590_n1020, DP_OP_102J5_124_3590_n1019,
         DP_OP_102J5_124_3590_n1018, DP_OP_102J5_124_3590_n1017,
         DP_OP_102J5_124_3590_n1016, DP_OP_102J5_124_3590_n1015,
         DP_OP_102J5_124_3590_n1014, DP_OP_102J5_124_3590_n1013,
         DP_OP_102J5_124_3590_n1012, DP_OP_102J5_124_3590_n1011,
         DP_OP_102J5_124_3590_n1010, DP_OP_102J5_124_3590_n1009,
         DP_OP_102J5_124_3590_n1008, DP_OP_102J5_124_3590_n1007,
         DP_OP_102J5_124_3590_n1006, DP_OP_102J5_124_3590_n1005,
         DP_OP_102J5_124_3590_n1004, DP_OP_102J5_124_3590_n1003,
         DP_OP_102J5_124_3590_n1002, DP_OP_102J5_124_3590_n1001,
         DP_OP_102J5_124_3590_n1000, DP_OP_102J5_124_3590_n999,
         DP_OP_102J5_124_3590_n998, DP_OP_102J5_124_3590_n997,
         DP_OP_102J5_124_3590_n996, DP_OP_102J5_124_3590_n995,
         DP_OP_102J5_124_3590_n994, DP_OP_102J5_124_3590_n993,
         DP_OP_102J5_124_3590_n992, DP_OP_102J5_124_3590_n991,
         DP_OP_102J5_124_3590_n990, DP_OP_102J5_124_3590_n989,
         DP_OP_102J5_124_3590_n988, DP_OP_102J5_124_3590_n987,
         DP_OP_102J5_124_3590_n986, DP_OP_102J5_124_3590_n985,
         DP_OP_102J5_124_3590_n984, DP_OP_102J5_124_3590_n983,
         DP_OP_102J5_124_3590_n982, DP_OP_102J5_124_3590_n981,
         DP_OP_102J5_124_3590_n980, DP_OP_102J5_124_3590_n979,
         DP_OP_102J5_124_3590_n978, DP_OP_102J5_124_3590_n977,
         DP_OP_102J5_124_3590_n976, DP_OP_102J5_124_3590_n975,
         DP_OP_102J5_124_3590_n974, DP_OP_102J5_124_3590_n973,
         DP_OP_102J5_124_3590_n972, DP_OP_102J5_124_3590_n971,
         DP_OP_102J5_124_3590_n970, DP_OP_102J5_124_3590_n969,
         DP_OP_102J5_124_3590_n968, DP_OP_102J5_124_3590_n967,
         DP_OP_102J5_124_3590_n966, DP_OP_102J5_124_3590_n965,
         DP_OP_102J5_124_3590_n964, DP_OP_102J5_124_3590_n963,
         DP_OP_102J5_124_3590_n962, DP_OP_102J5_124_3590_n961,
         DP_OP_102J5_124_3590_n960, DP_OP_102J5_124_3590_n959,
         DP_OP_102J5_124_3590_n958, DP_OP_102J5_124_3590_n957,
         DP_OP_102J5_124_3590_n956, DP_OP_102J5_124_3590_n955,
         DP_OP_102J5_124_3590_n954, DP_OP_102J5_124_3590_n953,
         DP_OP_102J5_124_3590_n952, DP_OP_102J5_124_3590_n951,
         DP_OP_102J5_124_3590_n950, DP_OP_102J5_124_3590_n949,
         DP_OP_102J5_124_3590_n948, DP_OP_102J5_124_3590_n947,
         DP_OP_102J5_124_3590_n946, DP_OP_102J5_124_3590_n945,
         DP_OP_102J5_124_3590_n944, DP_OP_102J5_124_3590_n943,
         DP_OP_102J5_124_3590_n942, DP_OP_102J5_124_3590_n941,
         DP_OP_102J5_124_3590_n940, DP_OP_102J5_124_3590_n939,
         DP_OP_102J5_124_3590_n938, DP_OP_102J5_124_3590_n937,
         DP_OP_102J5_124_3590_n936, DP_OP_102J5_124_3590_n935,
         DP_OP_102J5_124_3590_n934, DP_OP_102J5_124_3590_n933,
         DP_OP_102J5_124_3590_n932, DP_OP_102J5_124_3590_n931,
         DP_OP_102J5_124_3590_n930, DP_OP_102J5_124_3590_n929,
         DP_OP_102J5_124_3590_n928, DP_OP_102J5_124_3590_n927,
         DP_OP_102J5_124_3590_n926, DP_OP_102J5_124_3590_n925,
         DP_OP_102J5_124_3590_n924, DP_OP_102J5_124_3590_n923,
         DP_OP_102J5_124_3590_n922, DP_OP_102J5_124_3590_n921,
         DP_OP_102J5_124_3590_n920, DP_OP_102J5_124_3590_n919,
         DP_OP_102J5_124_3590_n918, DP_OP_102J5_124_3590_n917,
         DP_OP_102J5_124_3590_n916, DP_OP_102J5_124_3590_n915,
         DP_OP_102J5_124_3590_n914, DP_OP_102J5_124_3590_n913,
         DP_OP_102J5_124_3590_n912, DP_OP_102J5_124_3590_n911,
         DP_OP_102J5_124_3590_n910, DP_OP_102J5_124_3590_n909,
         DP_OP_102J5_124_3590_n908, DP_OP_102J5_124_3590_n907,
         DP_OP_102J5_124_3590_n906, DP_OP_102J5_124_3590_n905,
         DP_OP_102J5_124_3590_n904, DP_OP_102J5_124_3590_n903,
         DP_OP_102J5_124_3590_n902, DP_OP_102J5_124_3590_n901,
         DP_OP_102J5_124_3590_n900, DP_OP_102J5_124_3590_n899,
         DP_OP_102J5_124_3590_n898, DP_OP_102J5_124_3590_n897,
         DP_OP_102J5_124_3590_n896, DP_OP_102J5_124_3590_n895,
         DP_OP_102J5_124_3590_n894, DP_OP_102J5_124_3590_n893,
         DP_OP_102J5_124_3590_n892, DP_OP_102J5_124_3590_n891,
         DP_OP_102J5_124_3590_n890, DP_OP_102J5_124_3590_n889,
         DP_OP_102J5_124_3590_n888, DP_OP_102J5_124_3590_n887,
         DP_OP_102J5_124_3590_n886, DP_OP_102J5_124_3590_n885,
         DP_OP_102J5_124_3590_n884, DP_OP_102J5_124_3590_n883,
         DP_OP_102J5_124_3590_n882, DP_OP_102J5_124_3590_n881,
         DP_OP_102J5_124_3590_n880, DP_OP_102J5_124_3590_n879,
         DP_OP_102J5_124_3590_n878, DP_OP_102J5_124_3590_n877,
         DP_OP_102J5_124_3590_n876, DP_OP_102J5_124_3590_n875,
         DP_OP_102J5_124_3590_n874, DP_OP_102J5_124_3590_n873,
         DP_OP_102J5_124_3590_n872, DP_OP_102J5_124_3590_n871,
         DP_OP_102J5_124_3590_n870, DP_OP_102J5_124_3590_n869,
         DP_OP_102J5_124_3590_n868, DP_OP_102J5_124_3590_n867,
         DP_OP_102J5_124_3590_n866, DP_OP_102J5_124_3590_n865,
         DP_OP_102J5_124_3590_n864, DP_OP_102J5_124_3590_n863,
         DP_OP_102J5_124_3590_n862, DP_OP_102J5_124_3590_n861,
         DP_OP_102J5_124_3590_n860, DP_OP_102J5_124_3590_n859,
         DP_OP_102J5_124_3590_n858, DP_OP_102J5_124_3590_n857,
         DP_OP_102J5_124_3590_n856, DP_OP_102J5_124_3590_n855,
         DP_OP_102J5_124_3590_n854, DP_OP_102J5_124_3590_n853,
         DP_OP_102J5_124_3590_n852, DP_OP_102J5_124_3590_n851,
         DP_OP_102J5_124_3590_n850, DP_OP_102J5_124_3590_n849,
         DP_OP_102J5_124_3590_n848, DP_OP_102J5_124_3590_n847,
         DP_OP_102J5_124_3590_n846, DP_OP_102J5_124_3590_n845,
         DP_OP_102J5_124_3590_n844, DP_OP_102J5_124_3590_n843,
         DP_OP_102J5_124_3590_n842, DP_OP_102J5_124_3590_n841,
         DP_OP_102J5_124_3590_n840, DP_OP_102J5_124_3590_n839,
         DP_OP_102J5_124_3590_n838, DP_OP_102J5_124_3590_n837,
         DP_OP_102J5_124_3590_n836, DP_OP_102J5_124_3590_n835,
         DP_OP_102J5_124_3590_n834, DP_OP_102J5_124_3590_n833,
         DP_OP_102J5_124_3590_n832, DP_OP_102J5_124_3590_n831,
         DP_OP_102J5_124_3590_n830, DP_OP_102J5_124_3590_n829,
         DP_OP_102J5_124_3590_n828, DP_OP_102J5_124_3590_n827,
         DP_OP_102J5_124_3590_n826, DP_OP_102J5_124_3590_n825,
         DP_OP_102J5_124_3590_n824, DP_OP_102J5_124_3590_n823,
         DP_OP_102J5_124_3590_n822, DP_OP_102J5_124_3590_n821,
         DP_OP_102J5_124_3590_n820, DP_OP_102J5_124_3590_n819,
         DP_OP_102J5_124_3590_n818, DP_OP_102J5_124_3590_n817,
         DP_OP_102J5_124_3590_n816, DP_OP_102J5_124_3590_n815,
         DP_OP_102J5_124_3590_n814, DP_OP_102J5_124_3590_n813,
         DP_OP_102J5_124_3590_n812, DP_OP_102J5_124_3590_n811,
         DP_OP_102J5_124_3590_n810, DP_OP_102J5_124_3590_n809,
         DP_OP_102J5_124_3590_n808, DP_OP_102J5_124_3590_n807,
         DP_OP_102J5_124_3590_n806, DP_OP_102J5_124_3590_n805,
         DP_OP_102J5_124_3590_n804, DP_OP_102J5_124_3590_n803,
         DP_OP_102J5_124_3590_n802, DP_OP_102J5_124_3590_n801,
         DP_OP_102J5_124_3590_n800, DP_OP_102J5_124_3590_n799,
         DP_OP_102J5_124_3590_n798, DP_OP_102J5_124_3590_n797,
         DP_OP_102J5_124_3590_n796, DP_OP_102J5_124_3590_n795,
         DP_OP_102J5_124_3590_n794, DP_OP_102J5_124_3590_n793,
         DP_OP_102J5_124_3590_n792, DP_OP_102J5_124_3590_n791,
         DP_OP_102J5_124_3590_n790, DP_OP_102J5_124_3590_n789,
         DP_OP_102J5_124_3590_n788, DP_OP_102J5_124_3590_n787,
         DP_OP_102J5_124_3590_n786, DP_OP_102J5_124_3590_n785,
         DP_OP_102J5_124_3590_n784, DP_OP_102J5_124_3590_n783,
         DP_OP_102J5_124_3590_n782, DP_OP_102J5_124_3590_n781,
         DP_OP_102J5_124_3590_n780, DP_OP_102J5_124_3590_n779,
         DP_OP_102J5_124_3590_n778, DP_OP_102J5_124_3590_n777,
         DP_OP_102J5_124_3590_n776, DP_OP_102J5_124_3590_n775,
         DP_OP_102J5_124_3590_n774, DP_OP_102J5_124_3590_n773,
         DP_OP_102J5_124_3590_n772, DP_OP_102J5_124_3590_n771,
         DP_OP_102J5_124_3590_n770, DP_OP_102J5_124_3590_n769,
         DP_OP_102J5_124_3590_n768, DP_OP_102J5_124_3590_n767,
         DP_OP_102J5_124_3590_n766, DP_OP_102J5_124_3590_n765,
         DP_OP_102J5_124_3590_n764, DP_OP_102J5_124_3590_n763,
         DP_OP_102J5_124_3590_n762, DP_OP_102J5_124_3590_n761,
         DP_OP_102J5_124_3590_n760, DP_OP_102J5_124_3590_n759,
         DP_OP_102J5_124_3590_n758, DP_OP_102J5_124_3590_n757,
         DP_OP_102J5_124_3590_n756, DP_OP_102J5_124_3590_n755,
         DP_OP_102J5_124_3590_n754, DP_OP_102J5_124_3590_n753,
         DP_OP_102J5_124_3590_n752, DP_OP_102J5_124_3590_n751,
         DP_OP_102J5_124_3590_n750, DP_OP_102J5_124_3590_n749,
         DP_OP_102J5_124_3590_n748, DP_OP_102J5_124_3590_n747,
         DP_OP_102J5_124_3590_n746, DP_OP_102J5_124_3590_n745,
         DP_OP_102J5_124_3590_n744, DP_OP_102J5_124_3590_n743,
         DP_OP_102J5_124_3590_n742, DP_OP_102J5_124_3590_n741,
         DP_OP_102J5_124_3590_n740, DP_OP_102J5_124_3590_n739,
         DP_OP_102J5_124_3590_n738, DP_OP_102J5_124_3590_n737,
         DP_OP_102J5_124_3590_n736, DP_OP_102J5_124_3590_n735,
         DP_OP_102J5_124_3590_n734, DP_OP_102J5_124_3590_n733,
         DP_OP_102J5_124_3590_n732, DP_OP_102J5_124_3590_n731,
         DP_OP_102J5_124_3590_n730, DP_OP_102J5_124_3590_n729,
         DP_OP_102J5_124_3590_n728, DP_OP_102J5_124_3590_n727,
         DP_OP_102J5_124_3590_n726, DP_OP_102J5_124_3590_n725,
         DP_OP_102J5_124_3590_n724, DP_OP_102J5_124_3590_n723,
         DP_OP_102J5_124_3590_n722, DP_OP_102J5_124_3590_n721,
         DP_OP_102J5_124_3590_n720, DP_OP_102J5_124_3590_n719,
         DP_OP_102J5_124_3590_n718, DP_OP_102J5_124_3590_n717,
         DP_OP_102J5_124_3590_n716, DP_OP_102J5_124_3590_n715,
         DP_OP_102J5_124_3590_n714, DP_OP_102J5_124_3590_n713,
         DP_OP_102J5_124_3590_n712, DP_OP_102J5_124_3590_n711,
         DP_OP_102J5_124_3590_n710, DP_OP_102J5_124_3590_n709,
         DP_OP_102J5_124_3590_n708, DP_OP_102J5_124_3590_n707,
         DP_OP_102J5_124_3590_n706, DP_OP_102J5_124_3590_n705,
         DP_OP_102J5_124_3590_n704, DP_OP_102J5_124_3590_n703,
         DP_OP_102J5_124_3590_n702, DP_OP_102J5_124_3590_n701,
         DP_OP_102J5_124_3590_n700, DP_OP_102J5_124_3590_n699,
         DP_OP_102J5_124_3590_n698, DP_OP_102J5_124_3590_n697,
         DP_OP_102J5_124_3590_n696, DP_OP_102J5_124_3590_n695,
         DP_OP_102J5_124_3590_n694, DP_OP_102J5_124_3590_n693,
         DP_OP_102J5_124_3590_n692, DP_OP_102J5_124_3590_n691,
         DP_OP_102J5_124_3590_n690, DP_OP_102J5_124_3590_n689,
         DP_OP_102J5_124_3590_n688, DP_OP_102J5_124_3590_n687,
         DP_OP_102J5_124_3590_n686, DP_OP_102J5_124_3590_n685,
         DP_OP_102J5_124_3590_n684, DP_OP_102J5_124_3590_n683,
         DP_OP_102J5_124_3590_n682, DP_OP_102J5_124_3590_n681,
         DP_OP_102J5_124_3590_n680, DP_OP_102J5_124_3590_n679,
         DP_OP_102J5_124_3590_n678, DP_OP_102J5_124_3590_n677,
         DP_OP_102J5_124_3590_n676, DP_OP_102J5_124_3590_n675,
         DP_OP_102J5_124_3590_n674, DP_OP_102J5_124_3590_n673,
         DP_OP_102J5_124_3590_n672, DP_OP_102J5_124_3590_n671,
         DP_OP_102J5_124_3590_n670, DP_OP_102J5_124_3590_n669,
         DP_OP_102J5_124_3590_n668, DP_OP_102J5_124_3590_n667,
         DP_OP_102J5_124_3590_n666, DP_OP_102J5_124_3590_n665,
         DP_OP_102J5_124_3590_n664, DP_OP_102J5_124_3590_n663,
         DP_OP_102J5_124_3590_n662, DP_OP_102J5_124_3590_n661,
         DP_OP_102J5_124_3590_n660, DP_OP_102J5_124_3590_n659,
         DP_OP_102J5_124_3590_n658, DP_OP_102J5_124_3590_n657,
         DP_OP_102J5_124_3590_n656, DP_OP_102J5_124_3590_n655,
         DP_OP_102J5_124_3590_n654, DP_OP_102J5_124_3590_n653,
         DP_OP_102J5_124_3590_n652, DP_OP_102J5_124_3590_n651,
         DP_OP_102J5_124_3590_n650, DP_OP_102J5_124_3590_n649,
         DP_OP_102J5_124_3590_n648, DP_OP_102J5_124_3590_n647,
         DP_OP_102J5_124_3590_n646, DP_OP_102J5_124_3590_n645,
         DP_OP_102J5_124_3590_n644, DP_OP_102J5_124_3590_n643,
         DP_OP_102J5_124_3590_n642, DP_OP_102J5_124_3590_n641,
         DP_OP_102J5_124_3590_n640, DP_OP_102J5_124_3590_n639,
         DP_OP_102J5_124_3590_n638, DP_OP_102J5_124_3590_n637,
         DP_OP_102J5_124_3590_n636, DP_OP_102J5_124_3590_n635,
         DP_OP_102J5_124_3590_n634, DP_OP_102J5_124_3590_n633,
         DP_OP_102J5_124_3590_n632, DP_OP_102J5_124_3590_n631,
         DP_OP_102J5_124_3590_n630, DP_OP_102J5_124_3590_n629,
         DP_OP_102J5_124_3590_n628, DP_OP_102J5_124_3590_n627,
         DP_OP_102J5_124_3590_n626, DP_OP_102J5_124_3590_n625,
         DP_OP_102J5_124_3590_n624, DP_OP_102J5_124_3590_n623,
         DP_OP_102J5_124_3590_n622, DP_OP_102J5_124_3590_n621,
         DP_OP_102J5_124_3590_n620, DP_OP_102J5_124_3590_n619,
         DP_OP_102J5_124_3590_n618, DP_OP_102J5_124_3590_n617,
         DP_OP_102J5_124_3590_n616, DP_OP_102J5_124_3590_n615,
         DP_OP_102J5_124_3590_n614, DP_OP_102J5_124_3590_n613,
         DP_OP_102J5_124_3590_n612, DP_OP_102J5_124_3590_n611,
         DP_OP_102J5_124_3590_n610, DP_OP_102J5_124_3590_n609,
         DP_OP_102J5_124_3590_n608, DP_OP_102J5_124_3590_n607,
         DP_OP_102J5_124_3590_n606, DP_OP_102J5_124_3590_n605,
         DP_OP_102J5_124_3590_n604, DP_OP_102J5_124_3590_n603,
         DP_OP_102J5_124_3590_n602, DP_OP_102J5_124_3590_n601,
         DP_OP_102J5_124_3590_n600, DP_OP_102J5_124_3590_n599,
         DP_OP_102J5_124_3590_n598, DP_OP_102J5_124_3590_n597,
         DP_OP_102J5_124_3590_n596, DP_OP_102J5_124_3590_n595,
         DP_OP_102J5_124_3590_n594, DP_OP_102J5_124_3590_n593,
         DP_OP_102J5_124_3590_n592, DP_OP_102J5_124_3590_n591,
         DP_OP_102J5_124_3590_n590, DP_OP_102J5_124_3590_n589,
         DP_OP_102J5_124_3590_n588, DP_OP_102J5_124_3590_n587,
         DP_OP_102J5_124_3590_n586, DP_OP_102J5_124_3590_n585,
         DP_OP_102J5_124_3590_n584, DP_OP_102J5_124_3590_n583,
         DP_OP_102J5_124_3590_n582, DP_OP_102J5_124_3590_n581,
         DP_OP_102J5_124_3590_n580, DP_OP_102J5_124_3590_n579,
         DP_OP_102J5_124_3590_n578, DP_OP_102J5_124_3590_n577,
         DP_OP_102J5_124_3590_n576, DP_OP_102J5_124_3590_n575,
         DP_OP_102J5_124_3590_n574, DP_OP_102J5_124_3590_n573,
         DP_OP_102J5_124_3590_n572, DP_OP_102J5_124_3590_n571,
         DP_OP_102J5_124_3590_n570, DP_OP_102J5_124_3590_n569,
         DP_OP_102J5_124_3590_n568, DP_OP_102J5_124_3590_n567,
         DP_OP_102J5_124_3590_n566, DP_OP_102J5_124_3590_n565,
         DP_OP_102J5_124_3590_n564, DP_OP_102J5_124_3590_n563,
         DP_OP_102J5_124_3590_n562, DP_OP_102J5_124_3590_n561,
         DP_OP_102J5_124_3590_n560, DP_OP_102J5_124_3590_n559,
         DP_OP_102J5_124_3590_n558, DP_OP_102J5_124_3590_n557,
         DP_OP_102J5_124_3590_n556, DP_OP_102J5_124_3590_n555,
         DP_OP_102J5_124_3590_n554, DP_OP_102J5_124_3590_n553,
         DP_OP_102J5_124_3590_n552, DP_OP_102J5_124_3590_n551,
         DP_OP_102J5_124_3590_n550, DP_OP_102J5_124_3590_n549,
         DP_OP_102J5_124_3590_n548, DP_OP_102J5_124_3590_n547,
         DP_OP_102J5_124_3590_n546, DP_OP_102J5_124_3590_n545,
         DP_OP_102J5_124_3590_n544, DP_OP_102J5_124_3590_n543,
         DP_OP_102J5_124_3590_n542, DP_OP_102J5_124_3590_n541,
         DP_OP_102J5_124_3590_n540, DP_OP_102J5_124_3590_n539,
         DP_OP_102J5_124_3590_n538, DP_OP_102J5_124_3590_n537,
         DP_OP_102J5_124_3590_n536, DP_OP_102J5_124_3590_n535,
         DP_OP_102J5_124_3590_n534, DP_OP_102J5_124_3590_n533,
         DP_OP_102J5_124_3590_n532, DP_OP_102J5_124_3590_n531,
         DP_OP_102J5_124_3590_n530, DP_OP_102J5_124_3590_n529,
         DP_OP_102J5_124_3590_n528, DP_OP_102J5_124_3590_n527,
         DP_OP_102J5_124_3590_n526, DP_OP_102J5_124_3590_n525,
         DP_OP_102J5_124_3590_n524, DP_OP_102J5_124_3590_n523,
         DP_OP_102J5_124_3590_n522, DP_OP_102J5_124_3590_n521,
         DP_OP_102J5_124_3590_n520, DP_OP_102J5_124_3590_n519,
         DP_OP_102J5_124_3590_n518, DP_OP_102J5_124_3590_n517,
         DP_OP_102J5_124_3590_n516, DP_OP_102J5_124_3590_n515,
         DP_OP_102J5_124_3590_n514, DP_OP_102J5_124_3590_n513,
         DP_OP_102J5_124_3590_n512, DP_OP_102J5_124_3590_n511,
         DP_OP_102J5_124_3590_n510, DP_OP_102J5_124_3590_n509,
         DP_OP_102J5_124_3590_n508, DP_OP_102J5_124_3590_n507,
         DP_OP_102J5_124_3590_n506, DP_OP_102J5_124_3590_n505,
         DP_OP_102J5_124_3590_n504, DP_OP_102J5_124_3590_n503,
         DP_OP_102J5_124_3590_n502, DP_OP_102J5_124_3590_n501,
         DP_OP_102J5_124_3590_n500, DP_OP_102J5_124_3590_n499,
         DP_OP_102J5_124_3590_n498, DP_OP_102J5_124_3590_n497,
         DP_OP_102J5_124_3590_n496, DP_OP_102J5_124_3590_n495,
         DP_OP_102J5_124_3590_n494, DP_OP_102J5_124_3590_n493,
         DP_OP_102J5_124_3590_n492, DP_OP_102J5_124_3590_n491,
         DP_OP_102J5_124_3590_n490, DP_OP_102J5_124_3590_n489,
         DP_OP_102J5_124_3590_n488, DP_OP_102J5_124_3590_n487,
         DP_OP_102J5_124_3590_n486, DP_OP_102J5_124_3590_n485,
         DP_OP_102J5_124_3590_n484, DP_OP_102J5_124_3590_n483,
         DP_OP_102J5_124_3590_n482, DP_OP_102J5_124_3590_n481,
         DP_OP_102J5_124_3590_n480, DP_OP_102J5_124_3590_n479,
         DP_OP_102J5_124_3590_n478, DP_OP_102J5_124_3590_n477,
         DP_OP_102J5_124_3590_n476, DP_OP_102J5_124_3590_n475,
         DP_OP_102J5_124_3590_n474, DP_OP_102J5_124_3590_n473,
         DP_OP_102J5_124_3590_n472, DP_OP_102J5_124_3590_n471,
         DP_OP_102J5_124_3590_n470, DP_OP_102J5_124_3590_n469,
         DP_OP_102J5_124_3590_n468, DP_OP_102J5_124_3590_n467,
         DP_OP_102J5_124_3590_n466, DP_OP_102J5_124_3590_n465,
         DP_OP_102J5_124_3590_n464, DP_OP_102J5_124_3590_n463,
         DP_OP_102J5_124_3590_n462, DP_OP_102J5_124_3590_n461,
         DP_OP_102J5_124_3590_n460, DP_OP_102J5_124_3590_n459,
         DP_OP_102J5_124_3590_n458, DP_OP_102J5_124_3590_n457,
         DP_OP_102J5_124_3590_n456, DP_OP_102J5_124_3590_n455,
         DP_OP_102J5_124_3590_n454, DP_OP_102J5_124_3590_n453,
         DP_OP_102J5_124_3590_n452, DP_OP_102J5_124_3590_n451,
         DP_OP_102J5_124_3590_n450, DP_OP_102J5_124_3590_n449,
         DP_OP_102J5_124_3590_n448, DP_OP_102J5_124_3590_n447,
         DP_OP_102J5_124_3590_n446, DP_OP_102J5_124_3590_n445,
         DP_OP_102J5_124_3590_n444, DP_OP_102J5_124_3590_n443,
         DP_OP_102J5_124_3590_n442, DP_OP_102J5_124_3590_n441,
         DP_OP_102J5_124_3590_n440, DP_OP_102J5_124_3590_n439,
         DP_OP_102J5_124_3590_n438, DP_OP_102J5_124_3590_n437,
         DP_OP_102J5_124_3590_n436, DP_OP_102J5_124_3590_n435,
         DP_OP_102J5_124_3590_n434, DP_OP_102J5_124_3590_n433,
         DP_OP_102J5_124_3590_n432, DP_OP_102J5_124_3590_n431,
         DP_OP_102J5_124_3590_n430, DP_OP_102J5_124_3590_n429,
         DP_OP_102J5_124_3590_n428, DP_OP_102J5_124_3590_n427,
         DP_OP_102J5_124_3590_n426, DP_OP_102J5_124_3590_n425,
         DP_OP_102J5_124_3590_n424, DP_OP_102J5_124_3590_n423,
         DP_OP_102J5_124_3590_n422, DP_OP_102J5_124_3590_n421,
         DP_OP_102J5_124_3590_n420, DP_OP_102J5_124_3590_n419,
         DP_OP_102J5_124_3590_n418, DP_OP_102J5_124_3590_n417,
         DP_OP_102J5_124_3590_n416, DP_OP_102J5_124_3590_n415,
         DP_OP_102J5_124_3590_n414, DP_OP_102J5_124_3590_n413,
         DP_OP_102J5_124_3590_n412, DP_OP_102J5_124_3590_n411,
         DP_OP_102J5_124_3590_n410, DP_OP_102J5_124_3590_n409,
         DP_OP_102J5_124_3590_n408, DP_OP_102J5_124_3590_n407,
         DP_OP_102J5_124_3590_n406, DP_OP_102J5_124_3590_n405,
         DP_OP_102J5_124_3590_n404, DP_OP_102J5_124_3590_n403,
         DP_OP_102J5_124_3590_n402, DP_OP_102J5_124_3590_n401,
         DP_OP_102J5_124_3590_n400, DP_OP_102J5_124_3590_n399,
         DP_OP_102J5_124_3590_n398, DP_OP_102J5_124_3590_n397,
         DP_OP_102J5_124_3590_n396, DP_OP_102J5_124_3590_n395,
         DP_OP_102J5_124_3590_n394, DP_OP_102J5_124_3590_n393,
         DP_OP_102J5_124_3590_n392, DP_OP_102J5_124_3590_n391,
         DP_OP_102J5_124_3590_n390, DP_OP_102J5_124_3590_n389,
         DP_OP_102J5_124_3590_n388, DP_OP_102J5_124_3590_n387,
         DP_OP_102J5_124_3590_n386, DP_OP_102J5_124_3590_n385,
         DP_OP_102J5_124_3590_n384, DP_OP_102J5_124_3590_n383,
         DP_OP_102J5_124_3590_n382, DP_OP_102J5_124_3590_n381,
         DP_OP_102J5_124_3590_n380, DP_OP_102J5_124_3590_n379,
         DP_OP_102J5_124_3590_n378, DP_OP_102J5_124_3590_n377,
         DP_OP_102J5_124_3590_n376, DP_OP_102J5_124_3590_n375,
         DP_OP_102J5_124_3590_n374, DP_OP_102J5_124_3590_n373,
         DP_OP_102J5_124_3590_n372, DP_OP_102J5_124_3590_n371,
         DP_OP_102J5_124_3590_n370, DP_OP_102J5_124_3590_n369,
         DP_OP_102J5_124_3590_n368, DP_OP_102J5_124_3590_n367,
         DP_OP_102J5_124_3590_n366, DP_OP_102J5_124_3590_n365,
         DP_OP_102J5_124_3590_n364, DP_OP_102J5_124_3590_n363,
         DP_OP_102J5_124_3590_n362, DP_OP_102J5_124_3590_n361,
         DP_OP_102J5_124_3590_n360, DP_OP_102J5_124_3590_n359,
         DP_OP_102J5_124_3590_n358, DP_OP_102J5_124_3590_n357,
         DP_OP_102J5_124_3590_n356, DP_OP_102J5_124_3590_n355,
         DP_OP_102J5_124_3590_n354, DP_OP_102J5_124_3590_n353,
         DP_OP_102J5_124_3590_n352, DP_OP_102J5_124_3590_n351,
         DP_OP_102J5_124_3590_n350, DP_OP_102J5_124_3590_n349,
         DP_OP_102J5_124_3590_n348, DP_OP_102J5_124_3590_n347,
         DP_OP_102J5_124_3590_n346, DP_OP_102J5_124_3590_n345,
         DP_OP_102J5_124_3590_n344, DP_OP_102J5_124_3590_n343,
         DP_OP_102J5_124_3590_n342, DP_OP_102J5_124_3590_n341,
         DP_OP_102J5_124_3590_n340, DP_OP_102J5_124_3590_n339,
         DP_OP_102J5_124_3590_n338, DP_OP_102J5_124_3590_n337,
         DP_OP_102J5_124_3590_n336, DP_OP_102J5_124_3590_n335,
         DP_OP_102J5_124_3590_n334, DP_OP_102J5_124_3590_n333,
         DP_OP_102J5_124_3590_n332, DP_OP_102J5_124_3590_n331,
         DP_OP_102J5_124_3590_n330, DP_OP_102J5_124_3590_n329,
         DP_OP_102J5_124_3590_n328, DP_OP_102J5_124_3590_n327,
         DP_OP_102J5_124_3590_n326, DP_OP_102J5_124_3590_n325,
         DP_OP_102J5_124_3590_n324, DP_OP_102J5_124_3590_n323,
         DP_OP_102J5_124_3590_n322, DP_OP_102J5_124_3590_n321,
         DP_OP_102J5_124_3590_n320, DP_OP_102J5_124_3590_n319,
         DP_OP_102J5_124_3590_n318, DP_OP_102J5_124_3590_n317,
         DP_OP_102J5_124_3590_n316, DP_OP_102J5_124_3590_n315,
         DP_OP_102J5_124_3590_n314, DP_OP_102J5_124_3590_n313,
         DP_OP_102J5_124_3590_n312, DP_OP_102J5_124_3590_n311,
         DP_OP_102J5_124_3590_n310, DP_OP_102J5_124_3590_n309,
         DP_OP_102J5_124_3590_n308, DP_OP_102J5_124_3590_n307,
         DP_OP_102J5_124_3590_n306, DP_OP_102J5_124_3590_n305,
         DP_OP_102J5_124_3590_n304, DP_OP_102J5_124_3590_n303,
         DP_OP_102J5_124_3590_n302, DP_OP_102J5_124_3590_n301,
         DP_OP_102J5_124_3590_n300, DP_OP_102J5_124_3590_n299,
         DP_OP_102J5_124_3590_n298, DP_OP_102J5_124_3590_n297,
         DP_OP_102J5_124_3590_n296, DP_OP_102J5_124_3590_n295,
         DP_OP_102J5_124_3590_n294, DP_OP_102J5_124_3590_n293,
         DP_OP_102J5_124_3590_n292, DP_OP_102J5_124_3590_n291,
         DP_OP_102J5_124_3590_n290, DP_OP_102J5_124_3590_n289,
         DP_OP_102J5_124_3590_n288, DP_OP_102J5_124_3590_n287,
         DP_OP_102J5_124_3590_n286, DP_OP_102J5_124_3590_n285,
         DP_OP_102J5_124_3590_n284, DP_OP_102J5_124_3590_n283,
         DP_OP_102J5_124_3590_n282, DP_OP_102J5_124_3590_n281,
         DP_OP_102J5_124_3590_n280, DP_OP_102J5_124_3590_n279,
         DP_OP_102J5_124_3590_n278, DP_OP_102J5_124_3590_n277,
         DP_OP_102J5_124_3590_n276, DP_OP_102J5_124_3590_n275,
         DP_OP_102J5_124_3590_n274, DP_OP_102J5_124_3590_n273,
         DP_OP_102J5_124_3590_n272, DP_OP_102J5_124_3590_n271,
         DP_OP_102J5_124_3590_n270, DP_OP_102J5_124_3590_n269,
         DP_OP_102J5_124_3590_n268, DP_OP_102J5_124_3590_n267,
         DP_OP_102J5_124_3590_n266, DP_OP_102J5_124_3590_n265,
         DP_OP_102J5_124_3590_n264, DP_OP_102J5_124_3590_n263,
         DP_OP_102J5_124_3590_n262, DP_OP_102J5_124_3590_n261,
         DP_OP_102J5_124_3590_n260, DP_OP_102J5_124_3590_n259,
         DP_OP_102J5_124_3590_n258, DP_OP_102J5_124_3590_n257,
         DP_OP_102J5_124_3590_n256, DP_OP_102J5_124_3590_n255,
         DP_OP_102J5_124_3590_n254, DP_OP_102J5_124_3590_n253,
         DP_OP_102J5_124_3590_n252, DP_OP_102J5_124_3590_n251,
         DP_OP_102J5_124_3590_n250, DP_OP_102J5_124_3590_n249,
         DP_OP_102J5_124_3590_n248, DP_OP_102J5_124_3590_n247,
         DP_OP_102J5_124_3590_n246, DP_OP_102J5_124_3590_n245,
         DP_OP_102J5_124_3590_n244, DP_OP_102J5_124_3590_n243,
         DP_OP_102J5_124_3590_n242, DP_OP_102J5_124_3590_n241,
         DP_OP_102J5_124_3590_n240, DP_OP_102J5_124_3590_n239,
         DP_OP_102J5_124_3590_n238, DP_OP_102J5_124_3590_n237,
         DP_OP_102J5_124_3590_n236, DP_OP_102J5_124_3590_n235,
         DP_OP_102J5_124_3590_n234, DP_OP_102J5_124_3590_n233,
         DP_OP_102J5_124_3590_n232, DP_OP_102J5_124_3590_n231,
         DP_OP_102J5_124_3590_n230, DP_OP_102J5_124_3590_n229,
         DP_OP_102J5_124_3590_n228, DP_OP_102J5_124_3590_n227,
         DP_OP_102J5_124_3590_n226, DP_OP_102J5_124_3590_n225,
         DP_OP_102J5_124_3590_n224, DP_OP_102J5_124_3590_n223,
         DP_OP_102J5_124_3590_n222, DP_OP_102J5_124_3590_n221,
         DP_OP_102J5_124_3590_n220, DP_OP_102J5_124_3590_n219,
         DP_OP_102J5_124_3590_n218, DP_OP_102J5_124_3590_n217,
         DP_OP_102J5_124_3590_n216, DP_OP_102J5_124_3590_n215,
         DP_OP_102J5_124_3590_n214, DP_OP_102J5_124_3590_n213,
         DP_OP_102J5_124_3590_n212, DP_OP_102J5_124_3590_n211,
         DP_OP_102J5_124_3590_n210, DP_OP_102J5_124_3590_n209,
         DP_OP_102J5_124_3590_n208, DP_OP_102J5_124_3590_n207,
         DP_OP_102J5_124_3590_n206, DP_OP_102J5_124_3590_n205,
         DP_OP_102J5_124_3590_n204, DP_OP_102J5_124_3590_n203,
         DP_OP_102J5_124_3590_n202, DP_OP_102J5_124_3590_n201,
         DP_OP_102J5_124_3590_n200, DP_OP_102J5_124_3590_n199,
         DP_OP_102J5_124_3590_n198, DP_OP_102J5_124_3590_n197,
         DP_OP_102J5_124_3590_n196, DP_OP_102J5_124_3590_n195,
         DP_OP_102J5_124_3590_n194, DP_OP_102J5_124_3590_n193,
         DP_OP_102J5_124_3590_n192, DP_OP_102J5_124_3590_n191,
         DP_OP_102J5_124_3590_n190, DP_OP_102J5_124_3590_n189,
         DP_OP_102J5_124_3590_n188, DP_OP_102J5_124_3590_n187,
         DP_OP_102J5_124_3590_n186, DP_OP_102J5_124_3590_n185,
         DP_OP_102J5_124_3590_n184, DP_OP_102J5_124_3590_n183,
         DP_OP_102J5_124_3590_n182, DP_OP_102J5_124_3590_n181,
         DP_OP_102J5_124_3590_n180, DP_OP_102J5_124_3590_n179,
         DP_OP_102J5_124_3590_n178, DP_OP_102J5_124_3590_n177,
         DP_OP_102J5_124_3590_n176, DP_OP_102J5_124_3590_n175,
         DP_OP_102J5_124_3590_n174, DP_OP_102J5_124_3590_n173,
         DP_OP_102J5_124_3590_n172, DP_OP_102J5_124_3590_n171,
         DP_OP_102J5_124_3590_n170, DP_OP_102J5_124_3590_n169,
         DP_OP_102J5_124_3590_n168, DP_OP_102J5_124_3590_n167,
         DP_OP_102J5_124_3590_n166, DP_OP_102J5_124_3590_n165,
         DP_OP_102J5_124_3590_n164, DP_OP_102J5_124_3590_n163,
         DP_OP_102J5_124_3590_n162, DP_OP_102J5_124_3590_n161,
         DP_OP_102J5_124_3590_n160, DP_OP_102J5_124_3590_n159,
         DP_OP_102J5_124_3590_n158, DP_OP_102J5_124_3590_n157,
         DP_OP_102J5_124_3590_n156, DP_OP_102J5_124_3590_n155,
         DP_OP_102J5_124_3590_n154, DP_OP_102J5_124_3590_n153,
         DP_OP_102J5_124_3590_n152, DP_OP_102J5_124_3590_n151,
         DP_OP_102J5_124_3590_n150, DP_OP_102J5_124_3590_n149,
         DP_OP_102J5_124_3590_n148, DP_OP_102J5_124_3590_n147,
         DP_OP_102J5_124_3590_n146, DP_OP_102J5_124_3590_n145,
         DP_OP_102J5_124_3590_n144, DP_OP_102J5_124_3590_n143,
         DP_OP_102J5_124_3590_n142, DP_OP_102J5_124_3590_n141,
         DP_OP_102J5_124_3590_n140, DP_OP_102J5_124_3590_n139,
         DP_OP_102J5_124_3590_n138, DP_OP_102J5_124_3590_n137,
         DP_OP_102J5_124_3590_n116, DP_OP_102J5_124_3590_n115,
         DP_OP_102J5_124_3590_n114, DP_OP_102J5_124_3590_n113,
         DP_OP_102J5_124_3590_n112, DP_OP_102J5_124_3590_n106,
         DP_OP_102J5_124_3590_n102, DP_OP_102J5_124_3590_n101,
         DP_OP_102J5_124_3590_n100, DP_OP_102J5_124_3590_n99,
         DP_OP_102J5_124_3590_n98, DP_OP_102J5_124_3590_n94,
         DP_OP_102J5_124_3590_n93, DP_OP_102J5_124_3590_n92,
         DP_OP_102J5_124_3590_n91, DP_OP_102J5_124_3590_n90,
         DP_OP_102J5_124_3590_n89, DP_OP_102J5_124_3590_n88,
         DP_OP_102J5_124_3590_n86, DP_OP_102J5_124_3590_n85,
         DP_OP_102J5_124_3590_n82, DP_OP_102J5_124_3590_n81,
         DP_OP_102J5_124_3590_n80, DP_OP_102J5_124_3590_n79,
         DP_OP_102J5_124_3590_n77, DP_OP_102J5_124_3590_n75,
         DP_OP_102J5_124_3590_n74, DP_OP_102J5_124_3590_n73,
         DP_OP_102J5_124_3590_n72, DP_OP_102J5_124_3590_n71,
         DP_OP_102J5_124_3590_n70, DP_OP_102J5_124_3590_n69,
         DP_OP_102J5_124_3590_n67, DP_OP_102J5_124_3590_n66,
         DP_OP_102J5_124_3590_n61, DP_OP_102J5_124_3590_n60,
         DP_OP_102J5_124_3590_n59, DP_OP_102J5_124_3590_n58,
         DP_OP_102J5_124_3590_n57, DP_OP_102J5_124_3590_n56,
         DP_OP_102J5_124_3590_n54, DP_OP_102J5_124_3590_n52,
         DP_OP_102J5_124_3590_n51, DP_OP_102J5_124_3590_n50,
         DP_OP_102J5_124_3590_n48, DP_OP_102J5_124_3590_n47,
         DP_OP_102J5_124_3590_n45, DP_OP_102J5_124_3590_n43,
         DP_OP_102J5_124_3590_n42, DP_OP_102J5_124_3590_n41,
         DP_OP_102J5_124_3590_n37, DP_OP_102J5_124_3590_n33,
         DP_OP_102J5_124_3590_n32, DP_OP_102J5_124_3590_n30,
         DP_OP_102J5_124_3590_n29, DP_OP_102J5_124_3590_n28,
         DP_OP_102J5_124_3590_n27, DP_OP_102J5_124_3590_n25,
         DP_OP_102J5_124_3590_n24, DP_OP_102J5_124_3590_n23,
         DP_OP_102J5_124_3590_n4, DP_OP_102J5_124_3590_n2, n104, n105, n107,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272;
  wire   [22:0] n_accumulator_sum;

  DFFSSRX1_HVT fc_weight_box_reg_0__3_ ( .D(1'b0), .SETB(n160), .RSTB(
        sram_rdata_weight[79]), .CLK(clk), .QN(n177) );
  DFFSSRX1_HVT fc_weight_box_reg_0__2_ ( .D(1'b0), .SETB(n272), .RSTB(
        sram_rdata_weight[78]), .CLK(clk), .QN(n215) );
  DFFSSRX1_HVT fc_weight_box_reg_0__1_ ( .D(1'b0), .SETB(n159), .RSTB(
        sram_rdata_weight[77]), .CLK(clk), .QN(n216) );
  DFFSSRX1_HVT fc_weight_box_reg_0__0_ ( .D(1'b0), .SETB(n161), .RSTB(
        sram_rdata_weight[76]), .CLK(clk), .QN(n217) );
  DFFSSRX1_HVT fc_weight_box_reg_1__3_ ( .D(1'b0), .SETB(n160), .RSTB(
        sram_rdata_weight[75]), .CLK(clk), .QN(n178) );
  DFFSSRX1_HVT fc_weight_box_reg_1__2_ ( .D(1'b0), .SETB(n272), .RSTB(
        sram_rdata_weight[74]), .CLK(clk), .QN(n218) );
  DFFSSRX1_HVT fc_weight_box_reg_1__1_ ( .D(1'b0), .SETB(n159), .RSTB(
        sram_rdata_weight[73]), .CLK(clk), .QN(n219) );
  DFFSSRX1_HVT fc_weight_box_reg_1__0_ ( .D(1'b0), .SETB(n161), .RSTB(
        sram_rdata_weight[72]), .CLK(clk), .QN(n220) );
  DFFSSRX1_HVT fc_weight_box_reg_2__3_ ( .D(1'b0), .SETB(n160), .RSTB(
        sram_rdata_weight[71]), .CLK(clk), .QN(n176) );
  DFFSSRX1_HVT fc_weight_box_reg_2__2_ ( .D(1'b0), .SETB(n272), .RSTB(
        sram_rdata_weight[70]), .CLK(clk), .QN(n212) );
  DFFSSRX1_HVT fc_weight_box_reg_2__1_ ( .D(1'b0), .SETB(n159), .RSTB(
        sram_rdata_weight[69]), .CLK(clk), .QN(n213) );
  DFFSSRX1_HVT fc_weight_box_reg_2__0_ ( .D(1'b0), .SETB(n161), .RSTB(
        sram_rdata_weight[68]), .CLK(clk), .QN(n214) );
  DFFSSRX1_HVT fc_weight_box_reg_3__3_ ( .D(1'b0), .SETB(n160), .RSTB(
        sram_rdata_weight[67]), .CLK(clk), .QN(n179) );
  DFFSSRX1_HVT fc_weight_box_reg_3__2_ ( .D(1'b0), .SETB(n272), .RSTB(
        sram_rdata_weight[66]), .CLK(clk), .QN(n221) );
  DFFSSRX1_HVT fc_weight_box_reg_3__1_ ( .D(1'b0), .SETB(n159), .RSTB(
        sram_rdata_weight[65]), .CLK(clk), .QN(n222) );
  DFFSSRX1_HVT fc_weight_box_reg_3__0_ ( .D(1'b0), .SETB(n161), .RSTB(
        sram_rdata_weight[64]), .CLK(clk), .QN(n223) );
  DFFSSRX1_HVT fc_weight_box_reg_4__3_ ( .D(1'b0), .SETB(n160), .RSTB(
        sram_rdata_weight[63]), .CLK(clk), .QN(n175) );
  DFFSSRX1_HVT fc_weight_box_reg_4__2_ ( .D(1'b0), .SETB(n272), .RSTB(
        sram_rdata_weight[62]), .CLK(clk), .QN(n209) );
  DFFSSRX1_HVT fc_weight_box_reg_4__1_ ( .D(1'b0), .SETB(n159), .RSTB(
        sram_rdata_weight[61]), .CLK(clk), .QN(n210) );
  DFFSSRX1_HVT fc_weight_box_reg_4__0_ ( .D(1'b0), .SETB(n161), .RSTB(
        sram_rdata_weight[60]), .CLK(clk), .QN(n211) );
  DFFSSRX1_HVT fc_weight_box_reg_5__3_ ( .D(1'b0), .SETB(n160), .RSTB(
        sram_rdata_weight[59]), .CLK(clk), .QN(n180) );
  DFFSSRX1_HVT fc_weight_box_reg_5__2_ ( .D(1'b0), .SETB(n272), .RSTB(
        sram_rdata_weight[58]), .CLK(clk), .QN(n224) );
  DFFSSRX1_HVT fc_weight_box_reg_5__1_ ( .D(1'b0), .SETB(n159), .RSTB(
        sram_rdata_weight[57]), .CLK(clk), .QN(n225) );
  DFFSSRX1_HVT fc_weight_box_reg_5__0_ ( .D(1'b0), .SETB(n161), .RSTB(
        sram_rdata_weight[56]), .CLK(clk), .QN(n226) );
  DFFSSRX1_HVT fc_weight_box_reg_6__3_ ( .D(1'b0), .SETB(n160), .RSTB(
        sram_rdata_weight[55]), .CLK(clk), .QN(n174) );
  DFFSSRX1_HVT fc_weight_box_reg_6__2_ ( .D(1'b0), .SETB(n272), .RSTB(
        sram_rdata_weight[54]), .CLK(clk), .QN(n206) );
  DFFSSRX1_HVT fc_weight_box_reg_6__1_ ( .D(1'b0), .SETB(n159), .RSTB(
        sram_rdata_weight[53]), .CLK(clk), .QN(n207) );
  DFFSSRX1_HVT fc_weight_box_reg_6__0_ ( .D(1'b0), .SETB(n161), .RSTB(
        sram_rdata_weight[52]), .CLK(clk), .QN(n208) );
  DFFSSRX1_HVT fc_weight_box_reg_7__3_ ( .D(1'b0), .SETB(n160), .RSTB(
        sram_rdata_weight[51]), .CLK(clk), .QN(n181) );
  DFFSSRX1_HVT fc_weight_box_reg_7__2_ ( .D(1'b0), .SETB(n272), .RSTB(
        sram_rdata_weight[50]), .CLK(clk), .QN(n227) );
  DFFSSRX1_HVT fc_weight_box_reg_7__1_ ( .D(1'b0), .SETB(n159), .RSTB(
        sram_rdata_weight[49]), .CLK(clk), .QN(n228) );
  DFFSSRX1_HVT fc_weight_box_reg_7__0_ ( .D(1'b0), .SETB(n161), .RSTB(
        sram_rdata_weight[48]), .CLK(clk), .QN(n229) );
  DFFSSRX1_HVT fc_weight_box_reg_8__3_ ( .D(1'b0), .SETB(n160), .RSTB(
        sram_rdata_weight[47]), .CLK(clk), .QN(n173) );
  DFFSSRX1_HVT fc_weight_box_reg_8__2_ ( .D(1'b0), .SETB(n272), .RSTB(
        sram_rdata_weight[46]), .CLK(clk), .QN(n203) );
  DFFSSRX1_HVT fc_weight_box_reg_8__1_ ( .D(1'b0), .SETB(n159), .RSTB(
        sram_rdata_weight[45]), .CLK(clk), .QN(n204) );
  DFFSSRX1_HVT fc_weight_box_reg_8__0_ ( .D(1'b0), .SETB(n161), .RSTB(
        sram_rdata_weight[44]), .CLK(clk), .QN(n205) );
  DFFSSRX1_HVT fc_weight_box_reg_9__3_ ( .D(1'b0), .SETB(n160), .RSTB(
        sram_rdata_weight[43]), .CLK(clk), .QN(n182) );
  DFFSSRX1_HVT fc_weight_box_reg_9__2_ ( .D(1'b0), .SETB(n272), .RSTB(
        sram_rdata_weight[42]), .CLK(clk), .QN(n230) );
  DFFSSRX1_HVT fc_weight_box_reg_9__1_ ( .D(1'b0), .SETB(n159), .RSTB(
        sram_rdata_weight[41]), .CLK(clk), .QN(n231) );
  DFFSSRX1_HVT fc_weight_box_reg_9__0_ ( .D(1'b0), .SETB(n161), .RSTB(
        sram_rdata_weight[40]), .CLK(clk), .QN(n232) );
  DFFSSRX1_HVT fc_weight_box_reg_10__3_ ( .D(1'b0), .SETB(n160), .RSTB(
        sram_rdata_weight[39]), .CLK(clk), .QN(n172) );
  DFFSSRX1_HVT fc_weight_box_reg_10__2_ ( .D(1'b0), .SETB(n272), .RSTB(
        sram_rdata_weight[38]), .CLK(clk), .QN(n200) );
  DFFSSRX1_HVT fc_weight_box_reg_10__1_ ( .D(1'b0), .SETB(n159), .RSTB(
        sram_rdata_weight[37]), .CLK(clk), .QN(n201) );
  DFFSSRX1_HVT fc_weight_box_reg_10__0_ ( .D(1'b0), .SETB(n161), .RSTB(
        sram_rdata_weight[36]), .CLK(clk), .QN(n202) );
  DFFSSRX1_HVT fc_weight_box_reg_11__3_ ( .D(1'b0), .SETB(n160), .RSTB(
        sram_rdata_weight[35]), .CLK(clk), .QN(n183) );
  DFFSSRX1_HVT fc_weight_box_reg_11__2_ ( .D(1'b0), .SETB(n272), .RSTB(
        sram_rdata_weight[34]), .CLK(clk), .QN(n233) );
  DFFSSRX1_HVT fc_weight_box_reg_11__1_ ( .D(1'b0), .SETB(n159), .RSTB(
        sram_rdata_weight[33]), .CLK(clk), .QN(n234) );
  DFFSSRX1_HVT fc_weight_box_reg_11__0_ ( .D(1'b0), .SETB(n161), .RSTB(
        sram_rdata_weight[32]), .CLK(clk), .QN(n235) );
  DFFSSRX1_HVT fc_weight_box_reg_12__3_ ( .D(1'b0), .SETB(n160), .RSTB(
        sram_rdata_weight[31]), .CLK(clk), .QN(n171) );
  DFFSSRX1_HVT fc_weight_box_reg_12__2_ ( .D(1'b0), .SETB(n272), .RSTB(
        sram_rdata_weight[30]), .CLK(clk), .QN(n197) );
  DFFSSRX1_HVT fc_weight_box_reg_12__1_ ( .D(1'b0), .SETB(n159), .RSTB(
        sram_rdata_weight[29]), .CLK(clk), .QN(n198) );
  DFFSSRX1_HVT fc_weight_box_reg_12__0_ ( .D(1'b0), .SETB(n161), .RSTB(
        sram_rdata_weight[28]), .CLK(clk), .QN(n199) );
  DFFSSRX1_HVT fc_weight_box_reg_13__3_ ( .D(1'b0), .SETB(n160), .RSTB(
        sram_rdata_weight[27]), .CLK(clk), .QN(n184) );
  DFFSSRX1_HVT fc_weight_box_reg_13__2_ ( .D(1'b0), .SETB(n272), .RSTB(
        sram_rdata_weight[26]), .CLK(clk), .QN(n236) );
  DFFSSRX1_HVT fc_weight_box_reg_13__1_ ( .D(1'b0), .SETB(n159), .RSTB(
        sram_rdata_weight[25]), .CLK(clk), .QN(n237) );
  DFFSSRX1_HVT fc_weight_box_reg_13__0_ ( .D(1'b0), .SETB(n161), .RSTB(
        sram_rdata_weight[24]), .CLK(clk), .QN(n238) );
  DFFSSRX1_HVT fc_weight_box_reg_14__3_ ( .D(1'b0), .SETB(n160), .RSTB(
        sram_rdata_weight[23]), .CLK(clk), .QN(n170) );
  DFFSSRX1_HVT fc_weight_box_reg_14__2_ ( .D(1'b0), .SETB(n272), .RSTB(
        sram_rdata_weight[22]), .CLK(clk), .QN(n194) );
  DFFSSRX1_HVT fc_weight_box_reg_14__1_ ( .D(1'b0), .SETB(n159), .RSTB(
        sram_rdata_weight[21]), .CLK(clk), .QN(n195) );
  DFFSSRX1_HVT fc_weight_box_reg_14__0_ ( .D(1'b0), .SETB(n161), .RSTB(
        sram_rdata_weight[20]), .CLK(clk), .QN(n196) );
  DFFSSRX1_HVT fc_weight_box_reg_15__3_ ( .D(1'b0), .SETB(n160), .RSTB(
        sram_rdata_weight[19]), .CLK(clk), .QN(n185) );
  DFFSSRX1_HVT fc_weight_box_reg_15__2_ ( .D(1'b0), .SETB(n272), .RSTB(
        sram_rdata_weight[18]), .CLK(clk), .QN(n239) );
  DFFSSRX1_HVT fc_weight_box_reg_15__1_ ( .D(1'b0), .SETB(n159), .RSTB(
        sram_rdata_weight[17]), .CLK(clk), .QN(n240) );
  DFFSSRX1_HVT fc_weight_box_reg_15__0_ ( .D(1'b0), .SETB(n161), .RSTB(
        sram_rdata_weight[16]), .CLK(clk), .QN(n241) );
  DFFSSRX1_HVT fc_weight_box_reg_16__3_ ( .D(1'b0), .SETB(n160), .RSTB(
        sram_rdata_weight[15]), .CLK(clk), .QN(n169) );
  DFFSSRX1_HVT fc_weight_box_reg_16__2_ ( .D(1'b0), .SETB(n272), .RSTB(
        sram_rdata_weight[14]), .CLK(clk), .QN(n191) );
  DFFSSRX1_HVT fc_weight_box_reg_16__1_ ( .D(1'b0), .SETB(n159), .RSTB(
        sram_rdata_weight[13]), .CLK(clk), .QN(n192) );
  DFFSSRX1_HVT fc_weight_box_reg_16__0_ ( .D(1'b0), .SETB(n161), .RSTB(
        sram_rdata_weight[12]), .CLK(clk), .QN(n193) );
  DFFSSRX1_HVT fc_weight_box_reg_17__3_ ( .D(1'b0), .SETB(n160), .RSTB(
        sram_rdata_weight[11]), .CLK(clk), .QN(n186) );
  DFFSSRX1_HVT fc_weight_box_reg_17__2_ ( .D(1'b0), .SETB(n272), .RSTB(
        sram_rdata_weight[10]), .CLK(clk), .QN(n242) );
  DFFSSRX1_HVT fc_weight_box_reg_17__1_ ( .D(1'b0), .SETB(n159), .RSTB(
        sram_rdata_weight[9]), .CLK(clk), .QN(n243) );
  DFFSSRX1_HVT fc_weight_box_reg_17__0_ ( .D(1'b0), .SETB(n161), .RSTB(
        sram_rdata_weight[8]), .CLK(clk), .QN(n244) );
  DFFSSRX1_HVT fc_weight_box_reg_18__3_ ( .D(1'b0), .SETB(n160), .RSTB(
        sram_rdata_weight[7]), .CLK(clk), .QN(n168) );
  DFFSSRX1_HVT fc_weight_box_reg_18__2_ ( .D(1'b0), .SETB(n272), .RSTB(
        sram_rdata_weight[6]), .CLK(clk), .QN(n188) );
  DFFSSRX1_HVT fc_weight_box_reg_18__1_ ( .D(1'b0), .SETB(n159), .RSTB(
        sram_rdata_weight[5]), .CLK(clk), .QN(n189) );
  DFFSSRX1_HVT fc_weight_box_reg_18__0_ ( .D(1'b0), .SETB(n161), .RSTB(
        sram_rdata_weight[4]), .CLK(clk), .QN(n190) );
  DFFSSRX1_HVT fc_weight_box_reg_19__3_ ( .D(1'b0), .SETB(n160), .RSTB(
        sram_rdata_weight[3]), .CLK(clk), .QN(n187) );
  DFFSSRX1_HVT fc_weight_box_reg_19__2_ ( .D(1'b0), .SETB(n272), .RSTB(
        sram_rdata_weight[2]), .CLK(clk), .QN(n245) );
  DFFSSRX1_HVT fc_weight_box_reg_19__1_ ( .D(1'b0), .SETB(n159), .RSTB(
        sram_rdata_weight[1]), .CLK(clk), .QN(n246) );
  DFFSSRX1_HVT fc_weight_box_reg_19__0_ ( .D(1'b0), .SETB(n160), .RSTB(
        sram_rdata_weight[0]), .CLK(clk), .QN(n247) );
  DFFSSRX1_HVT accumulator_sum_reg_22_ ( .D(1'b0), .SETB(n161), .RSTB(
        n_accumulator_sum[22]), .CLK(clk), .Q(data_out[22]), .QN(n271) );
  DFFSSRX1_HVT accumulator_sum_reg_21_ ( .D(1'b0), .SETB(n160), .RSTB(
        n_accumulator_sum[21]), .CLK(clk), .Q(data_out[21]), .QN(n270) );
  DFFSSRX1_HVT accumulator_sum_reg_20_ ( .D(1'b0), .SETB(n272), .RSTB(
        n_accumulator_sum[20]), .CLK(clk), .Q(data_out[20]), .QN(n167) );
  DFFSSRX1_HVT accumulator_sum_reg_19_ ( .D(1'b0), .SETB(n159), .RSTB(
        n_accumulator_sum[19]), .CLK(clk), .Q(data_out[19]), .QN(n269) );
  DFFSSRX1_HVT accumulator_sum_reg_18_ ( .D(1'b0), .SETB(n161), .RSTB(
        n_accumulator_sum[18]), .CLK(clk), .Q(data_out[18]), .QN(n261) );
  DFFSSRX1_HVT accumulator_sum_reg_17_ ( .D(1'b0), .SETB(n160), .RSTB(
        n_accumulator_sum[17]), .CLK(clk), .Q(data_out[17]), .QN(n262) );
  DFFSSRX1_HVT accumulator_sum_reg_16_ ( .D(1'b0), .SETB(n272), .RSTB(
        n_accumulator_sum[16]), .CLK(clk), .Q(data_out[16]), .QN(n260) );
  DFFSSRX1_HVT accumulator_sum_reg_15_ ( .D(1'b0), .SETB(n159), .RSTB(
        n_accumulator_sum[15]), .CLK(clk), .Q(data_out[15]), .QN(n165) );
  DFFSSRX1_HVT accumulator_sum_reg_14_ ( .D(1'b0), .SETB(n161), .RSTB(
        n_accumulator_sum[14]), .CLK(clk), .Q(data_out[14]), .QN(n258) );
  DFFSSRX1_HVT accumulator_sum_reg_13_ ( .D(1'b0), .SETB(n160), .RSTB(
        n_accumulator_sum[13]), .CLK(clk), .Q(data_out[13]), .QN(n268) );
  DFFSSRX1_HVT accumulator_sum_reg_12_ ( .D(1'b0), .SETB(n272), .RSTB(
        n_accumulator_sum[12]), .CLK(clk), .Q(data_out[12]), .QN(n163) );
  DFFSSRX1_HVT accumulator_sum_reg_11_ ( .D(1'b0), .SETB(n159), .RSTB(
        n_accumulator_sum[11]), .CLK(clk), .Q(data_out[11]), .QN(n164) );
  DFFSSRX1_HVT accumulator_sum_reg_10_ ( .D(1'b0), .SETB(n161), .RSTB(
        n_accumulator_sum[10]), .CLK(clk), .Q(data_out[10]), .QN(n263) );
  DFFSSRX1_HVT accumulator_sum_reg_9_ ( .D(1'b0), .SETB(n160), .RSTB(
        n_accumulator_sum[9]), .CLK(clk), .Q(data_out[9]), .QN(n266) );
  DFFSSRX1_HVT accumulator_sum_reg_8_ ( .D(1'b0), .SETB(n159), .RSTB(
        n_accumulator_sum[8]), .CLK(clk), .Q(data_out[8]), .QN(n166) );
  DFFSSRX1_HVT accumulator_sum_reg_7_ ( .D(1'b0), .SETB(n159), .RSTB(
        n_accumulator_sum[7]), .CLK(clk), .Q(data_out[7]), .QN(n267) );
  DFFSSRX1_HVT accumulator_sum_reg_6_ ( .D(1'b0), .SETB(n161), .RSTB(
        n_accumulator_sum[6]), .CLK(clk), .Q(data_out[6]), .QN(n264) );
  DFFSSRX1_HVT accumulator_sum_reg_5_ ( .D(1'b0), .SETB(n160), .RSTB(
        n_accumulator_sum[5]), .CLK(clk), .Q(data_out[5]), .QN(n265) );
  DFFSSRX1_HVT accumulator_sum_reg_4_ ( .D(1'b0), .SETB(n159), .RSTB(
        n_accumulator_sum[4]), .CLK(clk), .Q(data_out[4]), .QN(n248) );
  DFFSSRX1_HVT accumulator_sum_reg_3_ ( .D(1'b0), .SETB(n159), .RSTB(
        n_accumulator_sum[3]), .CLK(clk), .Q(data_out[3]), .QN(n251) );
  DFFSSRX1_HVT accumulator_sum_reg_2_ ( .D(1'b0), .SETB(n161), .RSTB(
        n_accumulator_sum[2]), .CLK(clk), .Q(data_out[2]), .QN(n252) );
  DFFSSRX1_HVT accumulator_sum_reg_1_ ( .D(1'b0), .SETB(n160), .RSTB(
        n_accumulator_sum[1]), .CLK(clk), .Q(data_out[1]), .QN(n253) );
  DFFSSRX1_HVT accumulator_sum_reg_0_ ( .D(1'b0), .SETB(n161), .RSTB(
        n_accumulator_sum[0]), .CLK(clk), .Q(data_out[0]), .QN(n254) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1712 ( .A1(n247), .A2(
        DP_OP_102J5_124_3590_n2330), .Y(DP_OP_102J5_124_3590_n2322) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1711 ( .A1(n247), .A2(
        DP_OP_102J5_124_3590_n2329), .Y(DP_OP_102J5_124_3590_n2321) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1710 ( .A1(n247), .A2(
        DP_OP_102J5_124_3590_n2328), .Y(DP_OP_102J5_124_3590_n2320) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1709 ( .A1(n247), .A2(
        DP_OP_102J5_124_3590_n2327), .Y(DP_OP_102J5_124_3590_n2319) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1708 ( .A1(n247), .A2(
        DP_OP_102J5_124_3590_n2326), .Y(DP_OP_102J5_124_3590_n2318) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1707 ( .A1(n247), .A2(
        DP_OP_102J5_124_3590_n2325), .Y(DP_OP_102J5_124_3590_n2317) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1706 ( .A1(n247), .A2(
        DP_OP_102J5_124_3590_n2324), .Y(DP_OP_102J5_124_3590_n2316) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1705 ( .A1(n247), .A2(
        DP_OP_102J5_124_3590_n2323), .Y(DP_OP_102J5_124_3590_n700) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1704 ( .A1(n246), .A2(
        DP_OP_102J5_124_3590_n2330), .Y(DP_OP_102J5_124_3590_n2315) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1703 ( .A1(n246), .A2(
        DP_OP_102J5_124_3590_n2329), .Y(DP_OP_102J5_124_3590_n2314) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1702 ( .A1(n246), .A2(
        DP_OP_102J5_124_3590_n2328), .Y(DP_OP_102J5_124_3590_n2313) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1701 ( .A1(n246), .A2(
        DP_OP_102J5_124_3590_n2327), .Y(DP_OP_102J5_124_3590_n2312) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1700 ( .A1(n246), .A2(
        DP_OP_102J5_124_3590_n2326), .Y(DP_OP_102J5_124_3590_n2311) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1699 ( .A1(n246), .A2(
        DP_OP_102J5_124_3590_n2325), .Y(DP_OP_102J5_124_3590_n2310) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1698 ( .A1(n246), .A2(
        DP_OP_102J5_124_3590_n2324), .Y(DP_OP_102J5_124_3590_n2309) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1697 ( .A1(n246), .A2(
        DP_OP_102J5_124_3590_n2323), .Y(DP_OP_102J5_124_3590_n2308) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1696 ( .A1(n245), .A2(
        DP_OP_102J5_124_3590_n2330), .Y(DP_OP_102J5_124_3590_n2307) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1695 ( .A1(n245), .A2(
        DP_OP_102J5_124_3590_n2329), .Y(DP_OP_102J5_124_3590_n2306) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1694 ( .A1(n245), .A2(
        DP_OP_102J5_124_3590_n2328), .Y(DP_OP_102J5_124_3590_n2305) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1693 ( .A1(n245), .A2(
        DP_OP_102J5_124_3590_n2327), .Y(DP_OP_102J5_124_3590_n2304) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1692 ( .A1(n245), .A2(
        DP_OP_102J5_124_3590_n2326), .Y(DP_OP_102J5_124_3590_n2303) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1691 ( .A1(n245), .A2(
        DP_OP_102J5_124_3590_n2325), .Y(DP_OP_102J5_124_3590_n2302) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1690 ( .A1(n245), .A2(
        DP_OP_102J5_124_3590_n2324), .Y(DP_OP_102J5_124_3590_n2301) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1689 ( .A1(n245), .A2(
        DP_OP_102J5_124_3590_n2323), .Y(DP_OP_102J5_124_3590_n2300) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1688 ( .A1(n187), .A2(
        DP_OP_102J5_124_3590_n2330), .Y(DP_OP_102J5_124_3590_n2299) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1687 ( .A1(n187), .A2(
        DP_OP_102J5_124_3590_n2329), .Y(DP_OP_102J5_124_3590_n2298) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1686 ( .A1(n187), .A2(
        DP_OP_102J5_124_3590_n2328), .Y(DP_OP_102J5_124_3590_n2297) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1685 ( .A1(n187), .A2(
        DP_OP_102J5_124_3590_n2327), .Y(DP_OP_102J5_124_3590_n2296) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1684 ( .A1(n187), .A2(
        DP_OP_102J5_124_3590_n2326), .Y(DP_OP_102J5_124_3590_n2295) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1683 ( .A1(n187), .A2(
        DP_OP_102J5_124_3590_n2325), .Y(DP_OP_102J5_124_3590_n2294) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1682 ( .A1(n187), .A2(
        DP_OP_102J5_124_3590_n2324), .Y(DP_OP_102J5_124_3590_n2293) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1681 ( .A1(n187), .A2(
        DP_OP_102J5_124_3590_n2323), .Y(DP_OP_102J5_124_3590_n2292) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1668 ( .A1(n244), .A2(
        DP_OP_102J5_124_3590_n2287), .Y(DP_OP_102J5_124_3590_n2279) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1667 ( .A1(n244), .A2(
        DP_OP_102J5_124_3590_n2286), .Y(DP_OP_102J5_124_3590_n2278) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1666 ( .A1(n244), .A2(
        DP_OP_102J5_124_3590_n2285), .Y(DP_OP_102J5_124_3590_n2277) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1665 ( .A1(n244), .A2(
        DP_OP_102J5_124_3590_n2284), .Y(DP_OP_102J5_124_3590_n2276) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1664 ( .A1(n244), .A2(
        DP_OP_102J5_124_3590_n2283), .Y(DP_OP_102J5_124_3590_n2275) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1663 ( .A1(n244), .A2(
        DP_OP_102J5_124_3590_n2282), .Y(DP_OP_102J5_124_3590_n2274) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1662 ( .A1(n244), .A2(
        DP_OP_102J5_124_3590_n2281), .Y(DP_OP_102J5_124_3590_n2273) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1661 ( .A1(n244), .A2(
        DP_OP_102J5_124_3590_n2280), .Y(DP_OP_102J5_124_3590_n2272) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1660 ( .A1(n243), .A2(
        DP_OP_102J5_124_3590_n2287), .Y(DP_OP_102J5_124_3590_n2271) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1659 ( .A1(n243), .A2(
        DP_OP_102J5_124_3590_n2286), .Y(DP_OP_102J5_124_3590_n2270) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1658 ( .A1(n243), .A2(
        DP_OP_102J5_124_3590_n2285), .Y(DP_OP_102J5_124_3590_n2269) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1657 ( .A1(n243), .A2(
        DP_OP_102J5_124_3590_n2284), .Y(DP_OP_102J5_124_3590_n2268) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1656 ( .A1(n243), .A2(
        DP_OP_102J5_124_3590_n2283), .Y(DP_OP_102J5_124_3590_n2267) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1655 ( .A1(n243), .A2(
        DP_OP_102J5_124_3590_n2282), .Y(DP_OP_102J5_124_3590_n2266) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1654 ( .A1(n243), .A2(
        DP_OP_102J5_124_3590_n2281), .Y(DP_OP_102J5_124_3590_n2265) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1653 ( .A1(n243), .A2(
        DP_OP_102J5_124_3590_n2280), .Y(DP_OP_102J5_124_3590_n2264) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1652 ( .A1(n242), .A2(
        DP_OP_102J5_124_3590_n2287), .Y(DP_OP_102J5_124_3590_n2263) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1651 ( .A1(n242), .A2(
        DP_OP_102J5_124_3590_n2286), .Y(DP_OP_102J5_124_3590_n2262) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1650 ( .A1(n242), .A2(
        DP_OP_102J5_124_3590_n2285), .Y(DP_OP_102J5_124_3590_n2261) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1649 ( .A1(n242), .A2(
        DP_OP_102J5_124_3590_n2284), .Y(DP_OP_102J5_124_3590_n2260) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1648 ( .A1(n242), .A2(
        DP_OP_102J5_124_3590_n2283), .Y(DP_OP_102J5_124_3590_n2259) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1647 ( .A1(n242), .A2(
        DP_OP_102J5_124_3590_n2282), .Y(DP_OP_102J5_124_3590_n2258) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1646 ( .A1(n242), .A2(
        DP_OP_102J5_124_3590_n2281), .Y(DP_OP_102J5_124_3590_n2257) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1645 ( .A1(n242), .A2(
        DP_OP_102J5_124_3590_n2280), .Y(DP_OP_102J5_124_3590_n2256) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1644 ( .A1(n186), .A2(
        DP_OP_102J5_124_3590_n2287), .Y(DP_OP_102J5_124_3590_n2255) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1643 ( .A1(n186), .A2(
        DP_OP_102J5_124_3590_n2286), .Y(DP_OP_102J5_124_3590_n2254) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1642 ( .A1(n186), .A2(
        DP_OP_102J5_124_3590_n2285), .Y(DP_OP_102J5_124_3590_n2253) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1641 ( .A1(n186), .A2(
        DP_OP_102J5_124_3590_n2284), .Y(DP_OP_102J5_124_3590_n2252) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1640 ( .A1(n186), .A2(
        DP_OP_102J5_124_3590_n2283), .Y(DP_OP_102J5_124_3590_n2251) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1639 ( .A1(n186), .A2(
        DP_OP_102J5_124_3590_n2282), .Y(DP_OP_102J5_124_3590_n2250) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1638 ( .A1(n186), .A2(
        DP_OP_102J5_124_3590_n2281), .Y(DP_OP_102J5_124_3590_n2249) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1637 ( .A1(n186), .A2(
        DP_OP_102J5_124_3590_n2280), .Y(DP_OP_102J5_124_3590_n2248) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1624 ( .A1(n241), .A2(
        DP_OP_102J5_124_3590_n2243), .Y(DP_OP_102J5_124_3590_n2235) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1623 ( .A1(n241), .A2(
        DP_OP_102J5_124_3590_n2242), .Y(DP_OP_102J5_124_3590_n2234) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1622 ( .A1(n241), .A2(
        DP_OP_102J5_124_3590_n2241), .Y(DP_OP_102J5_124_3590_n2233) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1621 ( .A1(n241), .A2(
        DP_OP_102J5_124_3590_n2240), .Y(DP_OP_102J5_124_3590_n2232) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1620 ( .A1(n241), .A2(
        DP_OP_102J5_124_3590_n2239), .Y(DP_OP_102J5_124_3590_n2231) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1619 ( .A1(n241), .A2(
        DP_OP_102J5_124_3590_n2238), .Y(DP_OP_102J5_124_3590_n2230) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1618 ( .A1(n241), .A2(
        DP_OP_102J5_124_3590_n2237), .Y(DP_OP_102J5_124_3590_n2229) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1617 ( .A1(n241), .A2(
        DP_OP_102J5_124_3590_n2236), .Y(DP_OP_102J5_124_3590_n2228) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1616 ( .A1(n240), .A2(
        DP_OP_102J5_124_3590_n2243), .Y(DP_OP_102J5_124_3590_n2227) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1615 ( .A1(n240), .A2(
        DP_OP_102J5_124_3590_n2242), .Y(DP_OP_102J5_124_3590_n2226) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1614 ( .A1(n240), .A2(
        DP_OP_102J5_124_3590_n2241), .Y(DP_OP_102J5_124_3590_n2225) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1613 ( .A1(n240), .A2(
        DP_OP_102J5_124_3590_n2240), .Y(DP_OP_102J5_124_3590_n2224) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1612 ( .A1(n240), .A2(
        DP_OP_102J5_124_3590_n2239), .Y(DP_OP_102J5_124_3590_n2223) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1611 ( .A1(n240), .A2(
        DP_OP_102J5_124_3590_n2238), .Y(DP_OP_102J5_124_3590_n2222) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1610 ( .A1(n240), .A2(
        DP_OP_102J5_124_3590_n2237), .Y(DP_OP_102J5_124_3590_n2221) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1609 ( .A1(n240), .A2(
        DP_OP_102J5_124_3590_n2236), .Y(DP_OP_102J5_124_3590_n2220) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1608 ( .A1(n239), .A2(
        DP_OP_102J5_124_3590_n2243), .Y(DP_OP_102J5_124_3590_n2219) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1607 ( .A1(n239), .A2(
        DP_OP_102J5_124_3590_n2242), .Y(DP_OP_102J5_124_3590_n2218) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1606 ( .A1(n239), .A2(
        DP_OP_102J5_124_3590_n2241), .Y(DP_OP_102J5_124_3590_n2217) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1605 ( .A1(n239), .A2(
        DP_OP_102J5_124_3590_n2240), .Y(DP_OP_102J5_124_3590_n2216) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1604 ( .A1(n239), .A2(
        DP_OP_102J5_124_3590_n2239), .Y(DP_OP_102J5_124_3590_n2215) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1603 ( .A1(n239), .A2(
        DP_OP_102J5_124_3590_n2238), .Y(DP_OP_102J5_124_3590_n2214) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1602 ( .A1(n239), .A2(
        DP_OP_102J5_124_3590_n2237), .Y(DP_OP_102J5_124_3590_n2213) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1601 ( .A1(n239), .A2(
        DP_OP_102J5_124_3590_n2236), .Y(DP_OP_102J5_124_3590_n2212) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1600 ( .A1(n185), .A2(
        DP_OP_102J5_124_3590_n2243), .Y(DP_OP_102J5_124_3590_n2211) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1599 ( .A1(n185), .A2(
        DP_OP_102J5_124_3590_n2242), .Y(DP_OP_102J5_124_3590_n2210) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1598 ( .A1(n185), .A2(
        DP_OP_102J5_124_3590_n2241), .Y(DP_OP_102J5_124_3590_n2209) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1597 ( .A1(n185), .A2(
        DP_OP_102J5_124_3590_n2240), .Y(DP_OP_102J5_124_3590_n2208) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1596 ( .A1(n185), .A2(
        DP_OP_102J5_124_3590_n2239), .Y(DP_OP_102J5_124_3590_n2207) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1595 ( .A1(n185), .A2(
        DP_OP_102J5_124_3590_n2238), .Y(DP_OP_102J5_124_3590_n2206) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1594 ( .A1(n185), .A2(
        DP_OP_102J5_124_3590_n2237), .Y(DP_OP_102J5_124_3590_n2205) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1593 ( .A1(n185), .A2(
        DP_OP_102J5_124_3590_n2236), .Y(DP_OP_102J5_124_3590_n2204) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1580 ( .A1(n238), .A2(
        DP_OP_102J5_124_3590_n2199), .Y(DP_OP_102J5_124_3590_n2191) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1579 ( .A1(n238), .A2(
        DP_OP_102J5_124_3590_n2198), .Y(DP_OP_102J5_124_3590_n2190) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1578 ( .A1(n238), .A2(
        DP_OP_102J5_124_3590_n2197), .Y(DP_OP_102J5_124_3590_n2189) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1577 ( .A1(n238), .A2(
        DP_OP_102J5_124_3590_n2196), .Y(DP_OP_102J5_124_3590_n2188) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1576 ( .A1(n238), .A2(
        DP_OP_102J5_124_3590_n2195), .Y(DP_OP_102J5_124_3590_n2187) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1575 ( .A1(n238), .A2(
        DP_OP_102J5_124_3590_n2194), .Y(DP_OP_102J5_124_3590_n2186) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1574 ( .A1(n238), .A2(
        DP_OP_102J5_124_3590_n2193), .Y(DP_OP_102J5_124_3590_n2185) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1573 ( .A1(n238), .A2(
        DP_OP_102J5_124_3590_n2192), .Y(DP_OP_102J5_124_3590_n2184) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1572 ( .A1(n237), .A2(
        DP_OP_102J5_124_3590_n2199), .Y(DP_OP_102J5_124_3590_n2183) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1571 ( .A1(n237), .A2(
        DP_OP_102J5_124_3590_n2198), .Y(DP_OP_102J5_124_3590_n2182) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1570 ( .A1(n237), .A2(
        DP_OP_102J5_124_3590_n2197), .Y(DP_OP_102J5_124_3590_n2181) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1569 ( .A1(n237), .A2(
        DP_OP_102J5_124_3590_n2196), .Y(DP_OP_102J5_124_3590_n2180) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1568 ( .A1(n237), .A2(
        DP_OP_102J5_124_3590_n2195), .Y(DP_OP_102J5_124_3590_n2179) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1567 ( .A1(n237), .A2(
        DP_OP_102J5_124_3590_n2194), .Y(DP_OP_102J5_124_3590_n2178) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1566 ( .A1(n237), .A2(
        DP_OP_102J5_124_3590_n2193), .Y(DP_OP_102J5_124_3590_n2177) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1565 ( .A1(n237), .A2(
        DP_OP_102J5_124_3590_n2192), .Y(DP_OP_102J5_124_3590_n2176) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1564 ( .A1(n236), .A2(
        DP_OP_102J5_124_3590_n2199), .Y(DP_OP_102J5_124_3590_n2175) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1563 ( .A1(n236), .A2(
        DP_OP_102J5_124_3590_n2198), .Y(DP_OP_102J5_124_3590_n2174) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1562 ( .A1(n236), .A2(
        DP_OP_102J5_124_3590_n2197), .Y(DP_OP_102J5_124_3590_n2173) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1561 ( .A1(n236), .A2(
        DP_OP_102J5_124_3590_n2196), .Y(DP_OP_102J5_124_3590_n2172) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1560 ( .A1(n236), .A2(
        DP_OP_102J5_124_3590_n2195), .Y(DP_OP_102J5_124_3590_n2171) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1559 ( .A1(n236), .A2(
        DP_OP_102J5_124_3590_n2194), .Y(DP_OP_102J5_124_3590_n2170) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1558 ( .A1(n236), .A2(
        DP_OP_102J5_124_3590_n2193), .Y(DP_OP_102J5_124_3590_n2169) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1557 ( .A1(n236), .A2(
        DP_OP_102J5_124_3590_n2192), .Y(DP_OP_102J5_124_3590_n2168) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1556 ( .A1(n184), .A2(
        DP_OP_102J5_124_3590_n2199), .Y(DP_OP_102J5_124_3590_n2167) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1555 ( .A1(n184), .A2(
        DP_OP_102J5_124_3590_n2198), .Y(DP_OP_102J5_124_3590_n2166) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1554 ( .A1(n184), .A2(
        DP_OP_102J5_124_3590_n2197), .Y(DP_OP_102J5_124_3590_n2165) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1553 ( .A1(n184), .A2(
        DP_OP_102J5_124_3590_n2196), .Y(DP_OP_102J5_124_3590_n2164) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1552 ( .A1(n184), .A2(
        DP_OP_102J5_124_3590_n2195), .Y(DP_OP_102J5_124_3590_n2163) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1551 ( .A1(n184), .A2(
        DP_OP_102J5_124_3590_n2194), .Y(DP_OP_102J5_124_3590_n2162) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1550 ( .A1(n184), .A2(
        DP_OP_102J5_124_3590_n2193), .Y(DP_OP_102J5_124_3590_n2161) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1549 ( .A1(n184), .A2(
        DP_OP_102J5_124_3590_n2192), .Y(DP_OP_102J5_124_3590_n2160) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1536 ( .A1(n235), .A2(
        DP_OP_102J5_124_3590_n2155), .Y(DP_OP_102J5_124_3590_n2147) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1535 ( .A1(n235), .A2(
        DP_OP_102J5_124_3590_n2154), .Y(DP_OP_102J5_124_3590_n2146) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1534 ( .A1(n235), .A2(
        DP_OP_102J5_124_3590_n2153), .Y(DP_OP_102J5_124_3590_n2145) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1533 ( .A1(n235), .A2(
        DP_OP_102J5_124_3590_n2152), .Y(DP_OP_102J5_124_3590_n2144) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1532 ( .A1(n235), .A2(
        DP_OP_102J5_124_3590_n2151), .Y(DP_OP_102J5_124_3590_n2143) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1531 ( .A1(n235), .A2(
        DP_OP_102J5_124_3590_n2150), .Y(DP_OP_102J5_124_3590_n2142) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1530 ( .A1(n235), .A2(
        DP_OP_102J5_124_3590_n2149), .Y(DP_OP_102J5_124_3590_n2141) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1529 ( .A1(n235), .A2(
        DP_OP_102J5_124_3590_n2148), .Y(DP_OP_102J5_124_3590_n2140) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1528 ( .A1(n234), .A2(
        DP_OP_102J5_124_3590_n2155), .Y(DP_OP_102J5_124_3590_n2139) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1527 ( .A1(n234), .A2(
        DP_OP_102J5_124_3590_n2154), .Y(DP_OP_102J5_124_3590_n2138) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1526 ( .A1(n234), .A2(
        DP_OP_102J5_124_3590_n2153), .Y(DP_OP_102J5_124_3590_n2137) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1525 ( .A1(n234), .A2(
        DP_OP_102J5_124_3590_n2152), .Y(DP_OP_102J5_124_3590_n2136) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1524 ( .A1(n234), .A2(
        DP_OP_102J5_124_3590_n2151), .Y(DP_OP_102J5_124_3590_n2135) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1523 ( .A1(n234), .A2(
        DP_OP_102J5_124_3590_n2150), .Y(DP_OP_102J5_124_3590_n2134) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1522 ( .A1(n234), .A2(
        DP_OP_102J5_124_3590_n2149), .Y(DP_OP_102J5_124_3590_n2133) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1521 ( .A1(n234), .A2(
        DP_OP_102J5_124_3590_n2148), .Y(DP_OP_102J5_124_3590_n2132) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1520 ( .A1(n233), .A2(
        DP_OP_102J5_124_3590_n2155), .Y(DP_OP_102J5_124_3590_n2131) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1519 ( .A1(n233), .A2(
        DP_OP_102J5_124_3590_n2154), .Y(DP_OP_102J5_124_3590_n2130) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1518 ( .A1(n233), .A2(
        DP_OP_102J5_124_3590_n2153), .Y(DP_OP_102J5_124_3590_n2129) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1517 ( .A1(n233), .A2(
        DP_OP_102J5_124_3590_n2152), .Y(DP_OP_102J5_124_3590_n2128) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1516 ( .A1(n233), .A2(
        DP_OP_102J5_124_3590_n2151), .Y(DP_OP_102J5_124_3590_n2127) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1515 ( .A1(n233), .A2(
        DP_OP_102J5_124_3590_n2150), .Y(DP_OP_102J5_124_3590_n2126) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1514 ( .A1(n233), .A2(
        DP_OP_102J5_124_3590_n2149), .Y(DP_OP_102J5_124_3590_n2125) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1513 ( .A1(n233), .A2(
        DP_OP_102J5_124_3590_n2148), .Y(DP_OP_102J5_124_3590_n2124) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1512 ( .A1(n183), .A2(
        DP_OP_102J5_124_3590_n2155), .Y(DP_OP_102J5_124_3590_n2123) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1511 ( .A1(n183), .A2(
        DP_OP_102J5_124_3590_n2154), .Y(DP_OP_102J5_124_3590_n2122) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1510 ( .A1(n183), .A2(
        DP_OP_102J5_124_3590_n2153), .Y(DP_OP_102J5_124_3590_n2121) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1509 ( .A1(n183), .A2(
        DP_OP_102J5_124_3590_n2152), .Y(DP_OP_102J5_124_3590_n2120) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1508 ( .A1(n183), .A2(
        DP_OP_102J5_124_3590_n2151), .Y(DP_OP_102J5_124_3590_n2119) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1507 ( .A1(n183), .A2(
        DP_OP_102J5_124_3590_n2150), .Y(DP_OP_102J5_124_3590_n2118) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1506 ( .A1(n183), .A2(
        DP_OP_102J5_124_3590_n2149), .Y(DP_OP_102J5_124_3590_n2117) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1505 ( .A1(n183), .A2(
        DP_OP_102J5_124_3590_n2148), .Y(DP_OP_102J5_124_3590_n2116) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1492 ( .A1(n232), .A2(
        DP_OP_102J5_124_3590_n2111), .Y(DP_OP_102J5_124_3590_n2103) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1491 ( .A1(n232), .A2(
        DP_OP_102J5_124_3590_n2110), .Y(DP_OP_102J5_124_3590_n2102) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1490 ( .A1(n232), .A2(
        DP_OP_102J5_124_3590_n2109), .Y(DP_OP_102J5_124_3590_n2101) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1489 ( .A1(n232), .A2(
        DP_OP_102J5_124_3590_n2108), .Y(DP_OP_102J5_124_3590_n2100) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1488 ( .A1(n232), .A2(
        DP_OP_102J5_124_3590_n2107), .Y(DP_OP_102J5_124_3590_n2099) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1487 ( .A1(n232), .A2(
        DP_OP_102J5_124_3590_n2106), .Y(DP_OP_102J5_124_3590_n2098) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1486 ( .A1(n232), .A2(
        DP_OP_102J5_124_3590_n2105), .Y(DP_OP_102J5_124_3590_n2097) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1485 ( .A1(n232), .A2(
        DP_OP_102J5_124_3590_n2104), .Y(DP_OP_102J5_124_3590_n2096) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1484 ( .A1(n231), .A2(
        DP_OP_102J5_124_3590_n2111), .Y(DP_OP_102J5_124_3590_n2095) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1483 ( .A1(n231), .A2(
        DP_OP_102J5_124_3590_n2110), .Y(DP_OP_102J5_124_3590_n2094) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1482 ( .A1(n231), .A2(
        DP_OP_102J5_124_3590_n2109), .Y(DP_OP_102J5_124_3590_n2093) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1481 ( .A1(n231), .A2(
        DP_OP_102J5_124_3590_n2108), .Y(DP_OP_102J5_124_3590_n2092) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1480 ( .A1(n231), .A2(
        DP_OP_102J5_124_3590_n2107), .Y(DP_OP_102J5_124_3590_n2091) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1479 ( .A1(n231), .A2(
        DP_OP_102J5_124_3590_n2106), .Y(DP_OP_102J5_124_3590_n2090) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1478 ( .A1(n231), .A2(
        DP_OP_102J5_124_3590_n2105), .Y(DP_OP_102J5_124_3590_n2089) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1477 ( .A1(n231), .A2(
        DP_OP_102J5_124_3590_n2104), .Y(DP_OP_102J5_124_3590_n2088) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1476 ( .A1(n230), .A2(
        DP_OP_102J5_124_3590_n2111), .Y(DP_OP_102J5_124_3590_n2087) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1475 ( .A1(n230), .A2(
        DP_OP_102J5_124_3590_n2110), .Y(DP_OP_102J5_124_3590_n2086) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1474 ( .A1(n230), .A2(
        DP_OP_102J5_124_3590_n2109), .Y(DP_OP_102J5_124_3590_n2085) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1473 ( .A1(n230), .A2(
        DP_OP_102J5_124_3590_n2108), .Y(DP_OP_102J5_124_3590_n2084) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1472 ( .A1(n230), .A2(
        DP_OP_102J5_124_3590_n2107), .Y(DP_OP_102J5_124_3590_n2083) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1471 ( .A1(n230), .A2(
        DP_OP_102J5_124_3590_n2106), .Y(DP_OP_102J5_124_3590_n2082) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1470 ( .A1(n230), .A2(
        DP_OP_102J5_124_3590_n2105), .Y(DP_OP_102J5_124_3590_n2081) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1469 ( .A1(n230), .A2(
        DP_OP_102J5_124_3590_n2104), .Y(DP_OP_102J5_124_3590_n2080) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1468 ( .A1(n182), .A2(
        DP_OP_102J5_124_3590_n2111), .Y(DP_OP_102J5_124_3590_n2079) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1467 ( .A1(n182), .A2(
        DP_OP_102J5_124_3590_n2110), .Y(DP_OP_102J5_124_3590_n2078) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1466 ( .A1(n182), .A2(
        DP_OP_102J5_124_3590_n2109), .Y(DP_OP_102J5_124_3590_n2077) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1465 ( .A1(n182), .A2(
        DP_OP_102J5_124_3590_n2108), .Y(DP_OP_102J5_124_3590_n2076) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1464 ( .A1(n182), .A2(
        DP_OP_102J5_124_3590_n2107), .Y(DP_OP_102J5_124_3590_n2075) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1463 ( .A1(n182), .A2(
        DP_OP_102J5_124_3590_n2106), .Y(DP_OP_102J5_124_3590_n2074) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1462 ( .A1(n182), .A2(
        DP_OP_102J5_124_3590_n2105), .Y(DP_OP_102J5_124_3590_n2073) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1461 ( .A1(n182), .A2(
        DP_OP_102J5_124_3590_n2104), .Y(DP_OP_102J5_124_3590_n2072) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1448 ( .A1(n229), .A2(
        DP_OP_102J5_124_3590_n2067), .Y(DP_OP_102J5_124_3590_n2059) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1447 ( .A1(n229), .A2(
        DP_OP_102J5_124_3590_n2066), .Y(DP_OP_102J5_124_3590_n2058) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1446 ( .A1(n229), .A2(
        DP_OP_102J5_124_3590_n2065), .Y(DP_OP_102J5_124_3590_n2057) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1445 ( .A1(n229), .A2(
        DP_OP_102J5_124_3590_n2064), .Y(DP_OP_102J5_124_3590_n2056) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1444 ( .A1(n229), .A2(
        DP_OP_102J5_124_3590_n2063), .Y(DP_OP_102J5_124_3590_n2055) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1443 ( .A1(n229), .A2(
        DP_OP_102J5_124_3590_n2062), .Y(DP_OP_102J5_124_3590_n2054) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1442 ( .A1(n229), .A2(
        DP_OP_102J5_124_3590_n2061), .Y(DP_OP_102J5_124_3590_n2053) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1441 ( .A1(n229), .A2(
        DP_OP_102J5_124_3590_n2060), .Y(DP_OP_102J5_124_3590_n2052) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1440 ( .A1(n228), .A2(
        DP_OP_102J5_124_3590_n2067), .Y(DP_OP_102J5_124_3590_n2051) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1439 ( .A1(n228), .A2(
        DP_OP_102J5_124_3590_n2066), .Y(DP_OP_102J5_124_3590_n2050) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1438 ( .A1(n228), .A2(
        DP_OP_102J5_124_3590_n2065), .Y(DP_OP_102J5_124_3590_n2049) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1437 ( .A1(n228), .A2(
        DP_OP_102J5_124_3590_n2064), .Y(DP_OP_102J5_124_3590_n2048) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1436 ( .A1(n228), .A2(
        DP_OP_102J5_124_3590_n2063), .Y(DP_OP_102J5_124_3590_n2047) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1435 ( .A1(n228), .A2(
        DP_OP_102J5_124_3590_n2062), .Y(DP_OP_102J5_124_3590_n2046) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1434 ( .A1(n228), .A2(
        DP_OP_102J5_124_3590_n2061), .Y(DP_OP_102J5_124_3590_n2045) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1433 ( .A1(n228), .A2(
        DP_OP_102J5_124_3590_n2060), .Y(DP_OP_102J5_124_3590_n2044) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1432 ( .A1(n227), .A2(
        DP_OP_102J5_124_3590_n2067), .Y(DP_OP_102J5_124_3590_n2043) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1431 ( .A1(n227), .A2(
        DP_OP_102J5_124_3590_n2066), .Y(DP_OP_102J5_124_3590_n2042) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1430 ( .A1(n227), .A2(
        DP_OP_102J5_124_3590_n2065), .Y(DP_OP_102J5_124_3590_n2041) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1429 ( .A1(n227), .A2(
        DP_OP_102J5_124_3590_n2064), .Y(DP_OP_102J5_124_3590_n2040) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1428 ( .A1(n227), .A2(
        DP_OP_102J5_124_3590_n2063), .Y(DP_OP_102J5_124_3590_n2039) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1427 ( .A1(n227), .A2(
        DP_OP_102J5_124_3590_n2062), .Y(DP_OP_102J5_124_3590_n2038) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1426 ( .A1(n227), .A2(
        DP_OP_102J5_124_3590_n2061), .Y(DP_OP_102J5_124_3590_n2037) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1425 ( .A1(n227), .A2(
        DP_OP_102J5_124_3590_n2060), .Y(DP_OP_102J5_124_3590_n2036) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1424 ( .A1(n181), .A2(
        DP_OP_102J5_124_3590_n2067), .Y(DP_OP_102J5_124_3590_n2035) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1423 ( .A1(n181), .A2(
        DP_OP_102J5_124_3590_n2066), .Y(DP_OP_102J5_124_3590_n2034) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1422 ( .A1(n181), .A2(
        DP_OP_102J5_124_3590_n2065), .Y(DP_OP_102J5_124_3590_n2033) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1421 ( .A1(n181), .A2(
        DP_OP_102J5_124_3590_n2064), .Y(DP_OP_102J5_124_3590_n2032) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1420 ( .A1(n181), .A2(
        DP_OP_102J5_124_3590_n2063), .Y(DP_OP_102J5_124_3590_n2031) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1419 ( .A1(n181), .A2(
        DP_OP_102J5_124_3590_n2062), .Y(DP_OP_102J5_124_3590_n2030) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1418 ( .A1(n181), .A2(
        DP_OP_102J5_124_3590_n2061), .Y(DP_OP_102J5_124_3590_n2029) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1417 ( .A1(n181), .A2(
        DP_OP_102J5_124_3590_n2060), .Y(DP_OP_102J5_124_3590_n2028) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1404 ( .A1(n226), .A2(
        DP_OP_102J5_124_3590_n2023), .Y(DP_OP_102J5_124_3590_n2015) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1403 ( .A1(n226), .A2(
        DP_OP_102J5_124_3590_n2022), .Y(DP_OP_102J5_124_3590_n2014) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1402 ( .A1(n226), .A2(
        DP_OP_102J5_124_3590_n2021), .Y(DP_OP_102J5_124_3590_n2013) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1401 ( .A1(n226), .A2(
        DP_OP_102J5_124_3590_n2020), .Y(DP_OP_102J5_124_3590_n2012) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1400 ( .A1(n226), .A2(
        DP_OP_102J5_124_3590_n2019), .Y(DP_OP_102J5_124_3590_n2011) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1399 ( .A1(n226), .A2(
        DP_OP_102J5_124_3590_n2018), .Y(DP_OP_102J5_124_3590_n2010) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1398 ( .A1(n226), .A2(
        DP_OP_102J5_124_3590_n2017), .Y(DP_OP_102J5_124_3590_n2009) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1397 ( .A1(n226), .A2(
        DP_OP_102J5_124_3590_n2016), .Y(DP_OP_102J5_124_3590_n2008) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1396 ( .A1(n225), .A2(
        DP_OP_102J5_124_3590_n2023), .Y(DP_OP_102J5_124_3590_n2007) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1395 ( .A1(n225), .A2(
        DP_OP_102J5_124_3590_n2022), .Y(DP_OP_102J5_124_3590_n2006) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1394 ( .A1(n225), .A2(
        DP_OP_102J5_124_3590_n2021), .Y(DP_OP_102J5_124_3590_n2005) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1393 ( .A1(n225), .A2(
        DP_OP_102J5_124_3590_n2020), .Y(DP_OP_102J5_124_3590_n2004) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1392 ( .A1(n225), .A2(
        DP_OP_102J5_124_3590_n2019), .Y(DP_OP_102J5_124_3590_n2003) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1391 ( .A1(n225), .A2(
        DP_OP_102J5_124_3590_n2018), .Y(DP_OP_102J5_124_3590_n2002) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1390 ( .A1(n225), .A2(
        DP_OP_102J5_124_3590_n2017), .Y(DP_OP_102J5_124_3590_n2001) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1389 ( .A1(n225), .A2(
        DP_OP_102J5_124_3590_n2016), .Y(DP_OP_102J5_124_3590_n2000) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1388 ( .A1(n224), .A2(
        DP_OP_102J5_124_3590_n2023), .Y(DP_OP_102J5_124_3590_n1999) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1387 ( .A1(n224), .A2(
        DP_OP_102J5_124_3590_n2022), .Y(DP_OP_102J5_124_3590_n1998) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1386 ( .A1(n224), .A2(
        DP_OP_102J5_124_3590_n2021), .Y(DP_OP_102J5_124_3590_n1997) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1385 ( .A1(n224), .A2(
        DP_OP_102J5_124_3590_n2020), .Y(DP_OP_102J5_124_3590_n1996) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1384 ( .A1(n224), .A2(
        DP_OP_102J5_124_3590_n2019), .Y(DP_OP_102J5_124_3590_n1995) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1383 ( .A1(n224), .A2(
        DP_OP_102J5_124_3590_n2018), .Y(DP_OP_102J5_124_3590_n1994) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1382 ( .A1(n224), .A2(
        DP_OP_102J5_124_3590_n2017), .Y(DP_OP_102J5_124_3590_n1993) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1381 ( .A1(n224), .A2(
        DP_OP_102J5_124_3590_n2016), .Y(DP_OP_102J5_124_3590_n1992) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1380 ( .A1(n180), .A2(
        DP_OP_102J5_124_3590_n2023), .Y(DP_OP_102J5_124_3590_n1991) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1379 ( .A1(n180), .A2(
        DP_OP_102J5_124_3590_n2022), .Y(DP_OP_102J5_124_3590_n1990) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1378 ( .A1(n180), .A2(
        DP_OP_102J5_124_3590_n2021), .Y(DP_OP_102J5_124_3590_n1989) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1377 ( .A1(n180), .A2(
        DP_OP_102J5_124_3590_n2020), .Y(DP_OP_102J5_124_3590_n1988) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1376 ( .A1(n180), .A2(
        DP_OP_102J5_124_3590_n2019), .Y(DP_OP_102J5_124_3590_n1987) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1375 ( .A1(n180), .A2(
        DP_OP_102J5_124_3590_n2018), .Y(DP_OP_102J5_124_3590_n1986) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1374 ( .A1(n180), .A2(
        DP_OP_102J5_124_3590_n2017), .Y(DP_OP_102J5_124_3590_n1985) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1373 ( .A1(n180), .A2(
        DP_OP_102J5_124_3590_n2016), .Y(DP_OP_102J5_124_3590_n1984) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1360 ( .A1(n223), .A2(
        DP_OP_102J5_124_3590_n1979), .Y(DP_OP_102J5_124_3590_n1971) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1359 ( .A1(n223), .A2(
        DP_OP_102J5_124_3590_n1978), .Y(DP_OP_102J5_124_3590_n1970) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1358 ( .A1(n223), .A2(
        DP_OP_102J5_124_3590_n1977), .Y(DP_OP_102J5_124_3590_n1969) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1357 ( .A1(n223), .A2(
        DP_OP_102J5_124_3590_n1976), .Y(DP_OP_102J5_124_3590_n1968) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1356 ( .A1(n223), .A2(
        DP_OP_102J5_124_3590_n1975), .Y(DP_OP_102J5_124_3590_n1967) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1355 ( .A1(n223), .A2(
        DP_OP_102J5_124_3590_n1974), .Y(DP_OP_102J5_124_3590_n1966) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1354 ( .A1(n223), .A2(
        DP_OP_102J5_124_3590_n1973), .Y(DP_OP_102J5_124_3590_n1965) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1353 ( .A1(n223), .A2(
        DP_OP_102J5_124_3590_n1972), .Y(DP_OP_102J5_124_3590_n1964) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1352 ( .A1(n222), .A2(
        DP_OP_102J5_124_3590_n1979), .Y(DP_OP_102J5_124_3590_n1963) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1351 ( .A1(n222), .A2(
        DP_OP_102J5_124_3590_n1978), .Y(DP_OP_102J5_124_3590_n1962) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1350 ( .A1(n222), .A2(
        DP_OP_102J5_124_3590_n1977), .Y(DP_OP_102J5_124_3590_n1961) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1349 ( .A1(n222), .A2(
        DP_OP_102J5_124_3590_n1976), .Y(DP_OP_102J5_124_3590_n1960) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1348 ( .A1(n222), .A2(
        DP_OP_102J5_124_3590_n1975), .Y(DP_OP_102J5_124_3590_n1959) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1347 ( .A1(n222), .A2(
        DP_OP_102J5_124_3590_n1974), .Y(DP_OP_102J5_124_3590_n1958) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1346 ( .A1(n222), .A2(
        DP_OP_102J5_124_3590_n1973), .Y(DP_OP_102J5_124_3590_n1957) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1345 ( .A1(n222), .A2(
        DP_OP_102J5_124_3590_n1972), .Y(DP_OP_102J5_124_3590_n1956) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1344 ( .A1(n221), .A2(
        DP_OP_102J5_124_3590_n1979), .Y(DP_OP_102J5_124_3590_n1955) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1343 ( .A1(n221), .A2(
        DP_OP_102J5_124_3590_n1978), .Y(DP_OP_102J5_124_3590_n1954) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1342 ( .A1(n221), .A2(
        DP_OP_102J5_124_3590_n1977), .Y(DP_OP_102J5_124_3590_n1953) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1341 ( .A1(n221), .A2(
        DP_OP_102J5_124_3590_n1976), .Y(DP_OP_102J5_124_3590_n1952) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1340 ( .A1(n221), .A2(
        DP_OP_102J5_124_3590_n1975), .Y(DP_OP_102J5_124_3590_n1951) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1339 ( .A1(n221), .A2(
        DP_OP_102J5_124_3590_n1974), .Y(DP_OP_102J5_124_3590_n1950) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1338 ( .A1(n221), .A2(
        DP_OP_102J5_124_3590_n1973), .Y(DP_OP_102J5_124_3590_n1949) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1337 ( .A1(n221), .A2(
        DP_OP_102J5_124_3590_n1972), .Y(DP_OP_102J5_124_3590_n1948) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1336 ( .A1(n179), .A2(
        DP_OP_102J5_124_3590_n1979), .Y(DP_OP_102J5_124_3590_n1947) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1335 ( .A1(n179), .A2(
        DP_OP_102J5_124_3590_n1978), .Y(DP_OP_102J5_124_3590_n1946) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1334 ( .A1(n179), .A2(
        DP_OP_102J5_124_3590_n1977), .Y(DP_OP_102J5_124_3590_n1945) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1333 ( .A1(n179), .A2(
        DP_OP_102J5_124_3590_n1976), .Y(DP_OP_102J5_124_3590_n1944) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1332 ( .A1(n179), .A2(
        DP_OP_102J5_124_3590_n1975), .Y(DP_OP_102J5_124_3590_n1943) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1331 ( .A1(n179), .A2(
        DP_OP_102J5_124_3590_n1974), .Y(DP_OP_102J5_124_3590_n1942) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1330 ( .A1(n179), .A2(
        DP_OP_102J5_124_3590_n1973), .Y(DP_OP_102J5_124_3590_n1941) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1329 ( .A1(n179), .A2(
        DP_OP_102J5_124_3590_n1972), .Y(DP_OP_102J5_124_3590_n1940) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1316 ( .A1(n220), .A2(
        DP_OP_102J5_124_3590_n1935), .Y(DP_OP_102J5_124_3590_n1927) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1315 ( .A1(n220), .A2(
        DP_OP_102J5_124_3590_n1934), .Y(DP_OP_102J5_124_3590_n1926) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1314 ( .A1(n220), .A2(
        DP_OP_102J5_124_3590_n1933), .Y(DP_OP_102J5_124_3590_n1925) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1313 ( .A1(n220), .A2(
        DP_OP_102J5_124_3590_n1932), .Y(DP_OP_102J5_124_3590_n1924) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1312 ( .A1(n220), .A2(
        DP_OP_102J5_124_3590_n1931), .Y(DP_OP_102J5_124_3590_n1923) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1311 ( .A1(n220), .A2(
        DP_OP_102J5_124_3590_n1930), .Y(DP_OP_102J5_124_3590_n1922) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1310 ( .A1(n220), .A2(
        DP_OP_102J5_124_3590_n1929), .Y(DP_OP_102J5_124_3590_n1921) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1309 ( .A1(n220), .A2(
        DP_OP_102J5_124_3590_n1928), .Y(DP_OP_102J5_124_3590_n1920) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1308 ( .A1(n219), .A2(
        DP_OP_102J5_124_3590_n1935), .Y(DP_OP_102J5_124_3590_n1919) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1307 ( .A1(n219), .A2(
        DP_OP_102J5_124_3590_n1934), .Y(DP_OP_102J5_124_3590_n1918) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1306 ( .A1(n219), .A2(
        DP_OP_102J5_124_3590_n1933), .Y(DP_OP_102J5_124_3590_n1917) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1305 ( .A1(n219), .A2(
        DP_OP_102J5_124_3590_n1932), .Y(DP_OP_102J5_124_3590_n1916) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1304 ( .A1(n219), .A2(
        DP_OP_102J5_124_3590_n1931), .Y(DP_OP_102J5_124_3590_n1915) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1303 ( .A1(n219), .A2(
        DP_OP_102J5_124_3590_n1930), .Y(DP_OP_102J5_124_3590_n1914) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1302 ( .A1(n219), .A2(
        DP_OP_102J5_124_3590_n1929), .Y(DP_OP_102J5_124_3590_n1913) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1301 ( .A1(n219), .A2(
        DP_OP_102J5_124_3590_n1928), .Y(DP_OP_102J5_124_3590_n1912) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1300 ( .A1(n218), .A2(
        DP_OP_102J5_124_3590_n1935), .Y(DP_OP_102J5_124_3590_n1911) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1299 ( .A1(n218), .A2(
        DP_OP_102J5_124_3590_n1934), .Y(DP_OP_102J5_124_3590_n1910) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1298 ( .A1(n218), .A2(
        DP_OP_102J5_124_3590_n1933), .Y(DP_OP_102J5_124_3590_n1909) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1297 ( .A1(n218), .A2(
        DP_OP_102J5_124_3590_n1932), .Y(DP_OP_102J5_124_3590_n1908) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1296 ( .A1(n218), .A2(
        DP_OP_102J5_124_3590_n1931), .Y(DP_OP_102J5_124_3590_n1907) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1295 ( .A1(n218), .A2(
        DP_OP_102J5_124_3590_n1930), .Y(DP_OP_102J5_124_3590_n1906) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1294 ( .A1(n218), .A2(
        DP_OP_102J5_124_3590_n1929), .Y(DP_OP_102J5_124_3590_n1905) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1293 ( .A1(n218), .A2(
        DP_OP_102J5_124_3590_n1928), .Y(DP_OP_102J5_124_3590_n1904) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1292 ( .A1(n178), .A2(
        DP_OP_102J5_124_3590_n1935), .Y(DP_OP_102J5_124_3590_n1903) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1291 ( .A1(n178), .A2(
        DP_OP_102J5_124_3590_n1934), .Y(DP_OP_102J5_124_3590_n1902) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1290 ( .A1(n178), .A2(
        DP_OP_102J5_124_3590_n1933), .Y(DP_OP_102J5_124_3590_n1901) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1289 ( .A1(n178), .A2(
        DP_OP_102J5_124_3590_n1932), .Y(DP_OP_102J5_124_3590_n1900) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1288 ( .A1(n178), .A2(
        DP_OP_102J5_124_3590_n1931), .Y(DP_OP_102J5_124_3590_n1899) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1287 ( .A1(n178), .A2(
        DP_OP_102J5_124_3590_n1930), .Y(DP_OP_102J5_124_3590_n1898) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1286 ( .A1(n178), .A2(
        DP_OP_102J5_124_3590_n1929), .Y(DP_OP_102J5_124_3590_n1897) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1285 ( .A1(n178), .A2(
        DP_OP_102J5_124_3590_n1928), .Y(DP_OP_102J5_124_3590_n1896) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1272 ( .A1(n217), .A2(
        DP_OP_102J5_124_3590_n1891), .Y(DP_OP_102J5_124_3590_n1883) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1271 ( .A1(n217), .A2(
        DP_OP_102J5_124_3590_n1890), .Y(DP_OP_102J5_124_3590_n1882) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1270 ( .A1(n217), .A2(
        DP_OP_102J5_124_3590_n1889), .Y(DP_OP_102J5_124_3590_n1881) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1269 ( .A1(n217), .A2(
        DP_OP_102J5_124_3590_n1888), .Y(DP_OP_102J5_124_3590_n1880) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1268 ( .A1(n217), .A2(
        DP_OP_102J5_124_3590_n1887), .Y(DP_OP_102J5_124_3590_n1879) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1267 ( .A1(n217), .A2(
        DP_OP_102J5_124_3590_n1886), .Y(DP_OP_102J5_124_3590_n1878) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1266 ( .A1(n217), .A2(
        DP_OP_102J5_124_3590_n1885), .Y(DP_OP_102J5_124_3590_n1877) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1265 ( .A1(n217), .A2(
        DP_OP_102J5_124_3590_n1884), .Y(DP_OP_102J5_124_3590_n1876) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1264 ( .A1(n216), .A2(
        DP_OP_102J5_124_3590_n1891), .Y(DP_OP_102J5_124_3590_n1875) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1263 ( .A1(n216), .A2(
        DP_OP_102J5_124_3590_n1890), .Y(DP_OP_102J5_124_3590_n1874) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1262 ( .A1(n216), .A2(
        DP_OP_102J5_124_3590_n1889), .Y(DP_OP_102J5_124_3590_n1873) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1261 ( .A1(n216), .A2(
        DP_OP_102J5_124_3590_n1888), .Y(DP_OP_102J5_124_3590_n1872) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1260 ( .A1(n216), .A2(
        DP_OP_102J5_124_3590_n1887), .Y(DP_OP_102J5_124_3590_n1871) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1259 ( .A1(n216), .A2(
        DP_OP_102J5_124_3590_n1886), .Y(DP_OP_102J5_124_3590_n1870) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1258 ( .A1(n216), .A2(
        DP_OP_102J5_124_3590_n1885), .Y(DP_OP_102J5_124_3590_n1869) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1257 ( .A1(n216), .A2(
        DP_OP_102J5_124_3590_n1884), .Y(DP_OP_102J5_124_3590_n1868) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1256 ( .A1(n215), .A2(
        DP_OP_102J5_124_3590_n1891), .Y(DP_OP_102J5_124_3590_n1867) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1255 ( .A1(n215), .A2(
        DP_OP_102J5_124_3590_n1890), .Y(DP_OP_102J5_124_3590_n1866) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1254 ( .A1(n215), .A2(
        DP_OP_102J5_124_3590_n1889), .Y(DP_OP_102J5_124_3590_n1865) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1253 ( .A1(n215), .A2(
        DP_OP_102J5_124_3590_n1888), .Y(DP_OP_102J5_124_3590_n1864) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1252 ( .A1(n215), .A2(
        DP_OP_102J5_124_3590_n1887), .Y(DP_OP_102J5_124_3590_n1863) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1251 ( .A1(n215), .A2(
        DP_OP_102J5_124_3590_n1886), .Y(DP_OP_102J5_124_3590_n1862) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1250 ( .A1(n215), .A2(
        DP_OP_102J5_124_3590_n1885), .Y(DP_OP_102J5_124_3590_n1861) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1249 ( .A1(n215), .A2(
        DP_OP_102J5_124_3590_n1884), .Y(DP_OP_102J5_124_3590_n1860) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1248 ( .A1(n177), .A2(
        DP_OP_102J5_124_3590_n1891), .Y(DP_OP_102J5_124_3590_n1859) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1247 ( .A1(n177), .A2(
        DP_OP_102J5_124_3590_n1890), .Y(DP_OP_102J5_124_3590_n1858) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1246 ( .A1(n177), .A2(
        DP_OP_102J5_124_3590_n1889), .Y(DP_OP_102J5_124_3590_n1857) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1245 ( .A1(n177), .A2(
        DP_OP_102J5_124_3590_n1888), .Y(DP_OP_102J5_124_3590_n1856) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1244 ( .A1(n177), .A2(
        DP_OP_102J5_124_3590_n1887), .Y(DP_OP_102J5_124_3590_n1855) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1243 ( .A1(n177), .A2(
        DP_OP_102J5_124_3590_n1886), .Y(DP_OP_102J5_124_3590_n1854) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1242 ( .A1(n177), .A2(
        DP_OP_102J5_124_3590_n1885), .Y(DP_OP_102J5_124_3590_n1853) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1241 ( .A1(n177), .A2(
        DP_OP_102J5_124_3590_n1884), .Y(DP_OP_102J5_124_3590_n1852) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1228 ( .A1(n214), .A2(
        DP_OP_102J5_124_3590_n1847), .Y(DP_OP_102J5_124_3590_n1839) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1227 ( .A1(n214), .A2(
        DP_OP_102J5_124_3590_n1846), .Y(DP_OP_102J5_124_3590_n1838) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1226 ( .A1(n214), .A2(
        DP_OP_102J5_124_3590_n1845), .Y(DP_OP_102J5_124_3590_n1837) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1225 ( .A1(n214), .A2(
        DP_OP_102J5_124_3590_n1844), .Y(DP_OP_102J5_124_3590_n1836) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1224 ( .A1(n214), .A2(
        DP_OP_102J5_124_3590_n1843), .Y(DP_OP_102J5_124_3590_n1835) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1223 ( .A1(n214), .A2(
        DP_OP_102J5_124_3590_n1842), .Y(DP_OP_102J5_124_3590_n1834) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1222 ( .A1(n214), .A2(
        DP_OP_102J5_124_3590_n1841), .Y(DP_OP_102J5_124_3590_n1833) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1221 ( .A1(n214), .A2(
        DP_OP_102J5_124_3590_n1840), .Y(DP_OP_102J5_124_3590_n1832) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1220 ( .A1(n213), .A2(
        DP_OP_102J5_124_3590_n1847), .Y(DP_OP_102J5_124_3590_n1831) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1219 ( .A1(n213), .A2(
        DP_OP_102J5_124_3590_n1846), .Y(DP_OP_102J5_124_3590_n1830) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1218 ( .A1(n213), .A2(
        DP_OP_102J5_124_3590_n1845), .Y(DP_OP_102J5_124_3590_n1829) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1217 ( .A1(n213), .A2(
        DP_OP_102J5_124_3590_n1844), .Y(DP_OP_102J5_124_3590_n1828) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1216 ( .A1(n213), .A2(
        DP_OP_102J5_124_3590_n1843), .Y(DP_OP_102J5_124_3590_n1827) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1215 ( .A1(n213), .A2(
        DP_OP_102J5_124_3590_n1842), .Y(DP_OP_102J5_124_3590_n1826) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1214 ( .A1(n213), .A2(
        DP_OP_102J5_124_3590_n1841), .Y(DP_OP_102J5_124_3590_n1825) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1213 ( .A1(n213), .A2(
        DP_OP_102J5_124_3590_n1840), .Y(DP_OP_102J5_124_3590_n1824) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1212 ( .A1(n212), .A2(
        DP_OP_102J5_124_3590_n1847), .Y(DP_OP_102J5_124_3590_n1823) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1211 ( .A1(n212), .A2(
        DP_OP_102J5_124_3590_n1846), .Y(DP_OP_102J5_124_3590_n1822) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1210 ( .A1(n212), .A2(
        DP_OP_102J5_124_3590_n1845), .Y(DP_OP_102J5_124_3590_n1821) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1209 ( .A1(n212), .A2(
        DP_OP_102J5_124_3590_n1844), .Y(DP_OP_102J5_124_3590_n1820) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1208 ( .A1(n212), .A2(
        DP_OP_102J5_124_3590_n1843), .Y(DP_OP_102J5_124_3590_n1819) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1207 ( .A1(n212), .A2(
        DP_OP_102J5_124_3590_n1842), .Y(DP_OP_102J5_124_3590_n1818) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1206 ( .A1(n212), .A2(
        DP_OP_102J5_124_3590_n1841), .Y(DP_OP_102J5_124_3590_n1817) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1205 ( .A1(n212), .A2(
        DP_OP_102J5_124_3590_n1840), .Y(DP_OP_102J5_124_3590_n1816) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1204 ( .A1(n176), .A2(
        DP_OP_102J5_124_3590_n1847), .Y(DP_OP_102J5_124_3590_n1815) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1203 ( .A1(n176), .A2(
        DP_OP_102J5_124_3590_n1846), .Y(DP_OP_102J5_124_3590_n1814) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1202 ( .A1(n176), .A2(
        DP_OP_102J5_124_3590_n1845), .Y(DP_OP_102J5_124_3590_n1813) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1201 ( .A1(n176), .A2(
        DP_OP_102J5_124_3590_n1844), .Y(DP_OP_102J5_124_3590_n1812) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1200 ( .A1(n176), .A2(
        DP_OP_102J5_124_3590_n1843), .Y(DP_OP_102J5_124_3590_n1811) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1199 ( .A1(n176), .A2(
        DP_OP_102J5_124_3590_n1842), .Y(DP_OP_102J5_124_3590_n1810) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1198 ( .A1(n176), .A2(
        DP_OP_102J5_124_3590_n1841), .Y(DP_OP_102J5_124_3590_n1809) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1197 ( .A1(n176), .A2(
        DP_OP_102J5_124_3590_n1840), .Y(DP_OP_102J5_124_3590_n1808) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1184 ( .A1(n211), .A2(
        DP_OP_102J5_124_3590_n1803), .Y(DP_OP_102J5_124_3590_n1795) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1183 ( .A1(n211), .A2(
        DP_OP_102J5_124_3590_n1802), .Y(DP_OP_102J5_124_3590_n1794) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1182 ( .A1(n211), .A2(
        DP_OP_102J5_124_3590_n1801), .Y(DP_OP_102J5_124_3590_n1793) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1181 ( .A1(n211), .A2(
        DP_OP_102J5_124_3590_n1800), .Y(DP_OP_102J5_124_3590_n1792) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1180 ( .A1(n211), .A2(
        DP_OP_102J5_124_3590_n1799), .Y(DP_OP_102J5_124_3590_n1791) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1179 ( .A1(n211), .A2(
        DP_OP_102J5_124_3590_n1798), .Y(DP_OP_102J5_124_3590_n1790) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1177 ( .A1(n211), .A2(
        DP_OP_102J5_124_3590_n1796), .Y(DP_OP_102J5_124_3590_n1788) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1176 ( .A1(n210), .A2(
        DP_OP_102J5_124_3590_n1803), .Y(DP_OP_102J5_124_3590_n1787) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1175 ( .A1(n210), .A2(
        DP_OP_102J5_124_3590_n1802), .Y(DP_OP_102J5_124_3590_n1786) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1174 ( .A1(n210), .A2(
        DP_OP_102J5_124_3590_n1801), .Y(DP_OP_102J5_124_3590_n1785) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1173 ( .A1(n210), .A2(
        DP_OP_102J5_124_3590_n1800), .Y(DP_OP_102J5_124_3590_n1784) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1172 ( .A1(n210), .A2(
        DP_OP_102J5_124_3590_n1799), .Y(DP_OP_102J5_124_3590_n1783) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1171 ( .A1(n210), .A2(
        DP_OP_102J5_124_3590_n1798), .Y(DP_OP_102J5_124_3590_n1782) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1170 ( .A1(n210), .A2(
        DP_OP_102J5_124_3590_n1797), .Y(DP_OP_102J5_124_3590_n1781) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1169 ( .A1(n210), .A2(
        DP_OP_102J5_124_3590_n1796), .Y(DP_OP_102J5_124_3590_n1780) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1168 ( .A1(n209), .A2(
        DP_OP_102J5_124_3590_n1803), .Y(DP_OP_102J5_124_3590_n1779) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1167 ( .A1(n209), .A2(
        DP_OP_102J5_124_3590_n1802), .Y(DP_OP_102J5_124_3590_n1778) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1166 ( .A1(n209), .A2(
        DP_OP_102J5_124_3590_n1801), .Y(DP_OP_102J5_124_3590_n1777) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1165 ( .A1(n209), .A2(
        DP_OP_102J5_124_3590_n1800), .Y(DP_OP_102J5_124_3590_n1776) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1164 ( .A1(n209), .A2(
        DP_OP_102J5_124_3590_n1799), .Y(DP_OP_102J5_124_3590_n1775) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1163 ( .A1(n209), .A2(
        DP_OP_102J5_124_3590_n1798), .Y(DP_OP_102J5_124_3590_n1774) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1162 ( .A1(n209), .A2(
        DP_OP_102J5_124_3590_n1797), .Y(DP_OP_102J5_124_3590_n1773) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1161 ( .A1(n209), .A2(
        DP_OP_102J5_124_3590_n1796), .Y(DP_OP_102J5_124_3590_n1772) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1160 ( .A1(n175), .A2(
        DP_OP_102J5_124_3590_n1803), .Y(DP_OP_102J5_124_3590_n1771) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1159 ( .A1(n175), .A2(
        DP_OP_102J5_124_3590_n1802), .Y(DP_OP_102J5_124_3590_n1770) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1158 ( .A1(n175), .A2(
        DP_OP_102J5_124_3590_n1801), .Y(DP_OP_102J5_124_3590_n1769) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1157 ( .A1(n175), .A2(
        DP_OP_102J5_124_3590_n1800), .Y(DP_OP_102J5_124_3590_n1768) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1156 ( .A1(n175), .A2(
        DP_OP_102J5_124_3590_n1799), .Y(DP_OP_102J5_124_3590_n1767) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1155 ( .A1(n175), .A2(
        DP_OP_102J5_124_3590_n1798), .Y(DP_OP_102J5_124_3590_n1766) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1154 ( .A1(n175), .A2(
        DP_OP_102J5_124_3590_n1797), .Y(DP_OP_102J5_124_3590_n404) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1153 ( .A1(n175), .A2(
        DP_OP_102J5_124_3590_n1796), .Y(DP_OP_102J5_124_3590_n1765) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1140 ( .A1(n208), .A2(
        DP_OP_102J5_124_3590_n1760), .Y(DP_OP_102J5_124_3590_n1752) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1139 ( .A1(n208), .A2(
        DP_OP_102J5_124_3590_n1759), .Y(DP_OP_102J5_124_3590_n1751) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1138 ( .A1(n208), .A2(
        DP_OP_102J5_124_3590_n1758), .Y(DP_OP_102J5_124_3590_n1750) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1137 ( .A1(n208), .A2(
        DP_OP_102J5_124_3590_n1757), .Y(DP_OP_102J5_124_3590_n1749) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1136 ( .A1(n208), .A2(
        DP_OP_102J5_124_3590_n1756), .Y(DP_OP_102J5_124_3590_n1748) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1135 ( .A1(n208), .A2(
        DP_OP_102J5_124_3590_n1755), .Y(DP_OP_102J5_124_3590_n1747) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1134 ( .A1(n208), .A2(
        DP_OP_102J5_124_3590_n1754), .Y(DP_OP_102J5_124_3590_n1746) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1133 ( .A1(n208), .A2(
        DP_OP_102J5_124_3590_n1753), .Y(DP_OP_102J5_124_3590_n1745) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1132 ( .A1(n207), .A2(
        DP_OP_102J5_124_3590_n1760), .Y(DP_OP_102J5_124_3590_n1744) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1131 ( .A1(n207), .A2(
        DP_OP_102J5_124_3590_n1759), .Y(DP_OP_102J5_124_3590_n1743) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1130 ( .A1(n207), .A2(
        DP_OP_102J5_124_3590_n1758), .Y(DP_OP_102J5_124_3590_n1742) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1129 ( .A1(n207), .A2(
        DP_OP_102J5_124_3590_n1757), .Y(DP_OP_102J5_124_3590_n1741) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1128 ( .A1(n207), .A2(
        DP_OP_102J5_124_3590_n1756), .Y(DP_OP_102J5_124_3590_n1740) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1127 ( .A1(n207), .A2(
        DP_OP_102J5_124_3590_n1755), .Y(DP_OP_102J5_124_3590_n1739) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1126 ( .A1(n207), .A2(
        DP_OP_102J5_124_3590_n1754), .Y(DP_OP_102J5_124_3590_n1738) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1125 ( .A1(n207), .A2(
        DP_OP_102J5_124_3590_n1753), .Y(DP_OP_102J5_124_3590_n1737) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1124 ( .A1(n206), .A2(
        DP_OP_102J5_124_3590_n1760), .Y(DP_OP_102J5_124_3590_n1736) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1123 ( .A1(n206), .A2(
        DP_OP_102J5_124_3590_n1759), .Y(DP_OP_102J5_124_3590_n1735) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1122 ( .A1(n206), .A2(
        DP_OP_102J5_124_3590_n1758), .Y(DP_OP_102J5_124_3590_n1734) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1121 ( .A1(n206), .A2(
        DP_OP_102J5_124_3590_n1757), .Y(DP_OP_102J5_124_3590_n1733) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1120 ( .A1(n206), .A2(
        DP_OP_102J5_124_3590_n1756), .Y(DP_OP_102J5_124_3590_n1732) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1119 ( .A1(n206), .A2(
        DP_OP_102J5_124_3590_n1755), .Y(DP_OP_102J5_124_3590_n1731) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1118 ( .A1(n206), .A2(
        DP_OP_102J5_124_3590_n1754), .Y(DP_OP_102J5_124_3590_n1730) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1117 ( .A1(n206), .A2(
        DP_OP_102J5_124_3590_n1753), .Y(DP_OP_102J5_124_3590_n1729) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1116 ( .A1(n174), .A2(
        DP_OP_102J5_124_3590_n1760), .Y(DP_OP_102J5_124_3590_n1728) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1115 ( .A1(n174), .A2(
        DP_OP_102J5_124_3590_n1759), .Y(DP_OP_102J5_124_3590_n1727) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1114 ( .A1(n174), .A2(
        DP_OP_102J5_124_3590_n1758), .Y(DP_OP_102J5_124_3590_n1726) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1113 ( .A1(n174), .A2(
        DP_OP_102J5_124_3590_n1757), .Y(DP_OP_102J5_124_3590_n1725) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1112 ( .A1(n174), .A2(
        DP_OP_102J5_124_3590_n1756), .Y(DP_OP_102J5_124_3590_n1724) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1111 ( .A1(n174), .A2(
        DP_OP_102J5_124_3590_n1755), .Y(DP_OP_102J5_124_3590_n1723) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1110 ( .A1(n174), .A2(
        DP_OP_102J5_124_3590_n1754), .Y(DP_OP_102J5_124_3590_n1722) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1109 ( .A1(n174), .A2(
        DP_OP_102J5_124_3590_n1753), .Y(DP_OP_102J5_124_3590_n1721) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1096 ( .A1(n205), .A2(
        DP_OP_102J5_124_3590_n1716), .Y(DP_OP_102J5_124_3590_n1708) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1095 ( .A1(n205), .A2(
        DP_OP_102J5_124_3590_n1715), .Y(DP_OP_102J5_124_3590_n1707) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1094 ( .A1(n205), .A2(
        DP_OP_102J5_124_3590_n1714), .Y(DP_OP_102J5_124_3590_n1706) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1093 ( .A1(n205), .A2(
        DP_OP_102J5_124_3590_n1713), .Y(DP_OP_102J5_124_3590_n1705) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1092 ( .A1(n205), .A2(
        DP_OP_102J5_124_3590_n1712), .Y(DP_OP_102J5_124_3590_n1704) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1091 ( .A1(n205), .A2(
        DP_OP_102J5_124_3590_n1711), .Y(DP_OP_102J5_124_3590_n1703) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1090 ( .A1(n205), .A2(
        DP_OP_102J5_124_3590_n1710), .Y(DP_OP_102J5_124_3590_n1702) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1089 ( .A1(n205), .A2(
        DP_OP_102J5_124_3590_n1709), .Y(DP_OP_102J5_124_3590_n1701) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1088 ( .A1(n204), .A2(
        DP_OP_102J5_124_3590_n1716), .Y(DP_OP_102J5_124_3590_n1700) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1087 ( .A1(n204), .A2(
        DP_OP_102J5_124_3590_n1715), .Y(DP_OP_102J5_124_3590_n1699) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1086 ( .A1(n204), .A2(
        DP_OP_102J5_124_3590_n1714), .Y(DP_OP_102J5_124_3590_n1698) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1085 ( .A1(n204), .A2(
        DP_OP_102J5_124_3590_n1713), .Y(DP_OP_102J5_124_3590_n1697) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1084 ( .A1(n204), .A2(
        DP_OP_102J5_124_3590_n1712), .Y(DP_OP_102J5_124_3590_n1696) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1083 ( .A1(n204), .A2(
        DP_OP_102J5_124_3590_n1711), .Y(DP_OP_102J5_124_3590_n1695) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1082 ( .A1(n204), .A2(
        DP_OP_102J5_124_3590_n1710), .Y(DP_OP_102J5_124_3590_n1694) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1081 ( .A1(n204), .A2(
        DP_OP_102J5_124_3590_n1709), .Y(DP_OP_102J5_124_3590_n1693) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1080 ( .A1(n203), .A2(
        DP_OP_102J5_124_3590_n1716), .Y(DP_OP_102J5_124_3590_n1692) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1079 ( .A1(n203), .A2(
        DP_OP_102J5_124_3590_n1715), .Y(DP_OP_102J5_124_3590_n1691) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1078 ( .A1(n203), .A2(
        DP_OP_102J5_124_3590_n1714), .Y(DP_OP_102J5_124_3590_n1690) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1077 ( .A1(n203), .A2(
        DP_OP_102J5_124_3590_n1713), .Y(DP_OP_102J5_124_3590_n1689) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1076 ( .A1(n203), .A2(
        DP_OP_102J5_124_3590_n1712), .Y(DP_OP_102J5_124_3590_n1688) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1075 ( .A1(n203), .A2(
        DP_OP_102J5_124_3590_n1711), .Y(DP_OP_102J5_124_3590_n1687) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1074 ( .A1(n203), .A2(
        DP_OP_102J5_124_3590_n1710), .Y(DP_OP_102J5_124_3590_n1686) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1073 ( .A1(n203), .A2(
        DP_OP_102J5_124_3590_n1709), .Y(DP_OP_102J5_124_3590_n1685) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1072 ( .A1(n173), .A2(
        DP_OP_102J5_124_3590_n1716), .Y(DP_OP_102J5_124_3590_n1684) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1071 ( .A1(n173), .A2(
        DP_OP_102J5_124_3590_n1715), .Y(DP_OP_102J5_124_3590_n1683) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1070 ( .A1(n173), .A2(
        DP_OP_102J5_124_3590_n1714), .Y(DP_OP_102J5_124_3590_n1682) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1069 ( .A1(n173), .A2(
        DP_OP_102J5_124_3590_n1713), .Y(DP_OP_102J5_124_3590_n1681) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1068 ( .A1(n173), .A2(
        DP_OP_102J5_124_3590_n1712), .Y(DP_OP_102J5_124_3590_n1680) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1067 ( .A1(n173), .A2(
        DP_OP_102J5_124_3590_n1711), .Y(DP_OP_102J5_124_3590_n1679) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1066 ( .A1(n173), .A2(
        DP_OP_102J5_124_3590_n1710), .Y(DP_OP_102J5_124_3590_n1678) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1065 ( .A1(n173), .A2(
        DP_OP_102J5_124_3590_n1709), .Y(DP_OP_102J5_124_3590_n1677) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1052 ( .A1(n202), .A2(
        DP_OP_102J5_124_3590_n1672), .Y(DP_OP_102J5_124_3590_n1664) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1051 ( .A1(n202), .A2(
        DP_OP_102J5_124_3590_n1671), .Y(DP_OP_102J5_124_3590_n1663) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1050 ( .A1(n202), .A2(
        DP_OP_102J5_124_3590_n1670), .Y(DP_OP_102J5_124_3590_n1662) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1049 ( .A1(n202), .A2(
        DP_OP_102J5_124_3590_n1669), .Y(DP_OP_102J5_124_3590_n1661) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1048 ( .A1(n202), .A2(
        DP_OP_102J5_124_3590_n1668), .Y(DP_OP_102J5_124_3590_n1660) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1047 ( .A1(n202), .A2(
        DP_OP_102J5_124_3590_n1667), .Y(DP_OP_102J5_124_3590_n1659) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1046 ( .A1(n202), .A2(
        DP_OP_102J5_124_3590_n1666), .Y(DP_OP_102J5_124_3590_n1658) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1045 ( .A1(n202), .A2(
        DP_OP_102J5_124_3590_n1665), .Y(DP_OP_102J5_124_3590_n1657) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1044 ( .A1(n201), .A2(
        DP_OP_102J5_124_3590_n1672), .Y(DP_OP_102J5_124_3590_n1656) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1043 ( .A1(n201), .A2(
        DP_OP_102J5_124_3590_n1671), .Y(DP_OP_102J5_124_3590_n1655) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1042 ( .A1(n201), .A2(
        DP_OP_102J5_124_3590_n1670), .Y(DP_OP_102J5_124_3590_n1654) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1041 ( .A1(n201), .A2(
        DP_OP_102J5_124_3590_n1669), .Y(DP_OP_102J5_124_3590_n1653) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1040 ( .A1(n201), .A2(
        DP_OP_102J5_124_3590_n1668), .Y(DP_OP_102J5_124_3590_n1652) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1039 ( .A1(n201), .A2(
        DP_OP_102J5_124_3590_n1667), .Y(DP_OP_102J5_124_3590_n1651) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1038 ( .A1(n201), .A2(
        DP_OP_102J5_124_3590_n1666), .Y(DP_OP_102J5_124_3590_n1650) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1037 ( .A1(n201), .A2(
        DP_OP_102J5_124_3590_n1665), .Y(DP_OP_102J5_124_3590_n1649) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1036 ( .A1(n200), .A2(
        DP_OP_102J5_124_3590_n1672), .Y(DP_OP_102J5_124_3590_n1648) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1035 ( .A1(n200), .A2(
        DP_OP_102J5_124_3590_n1671), .Y(DP_OP_102J5_124_3590_n1647) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1034 ( .A1(n200), .A2(
        DP_OP_102J5_124_3590_n1670), .Y(DP_OP_102J5_124_3590_n1646) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1033 ( .A1(n200), .A2(
        DP_OP_102J5_124_3590_n1669), .Y(DP_OP_102J5_124_3590_n1645) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1032 ( .A1(n200), .A2(
        DP_OP_102J5_124_3590_n1668), .Y(DP_OP_102J5_124_3590_n1644) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1031 ( .A1(n200), .A2(
        DP_OP_102J5_124_3590_n1667), .Y(DP_OP_102J5_124_3590_n1643) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1030 ( .A1(n200), .A2(
        DP_OP_102J5_124_3590_n1666), .Y(DP_OP_102J5_124_3590_n1642) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1029 ( .A1(n200), .A2(
        DP_OP_102J5_124_3590_n1665), .Y(DP_OP_102J5_124_3590_n1641) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1028 ( .A1(n172), .A2(
        DP_OP_102J5_124_3590_n1672), .Y(DP_OP_102J5_124_3590_n1640) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1027 ( .A1(n172), .A2(
        DP_OP_102J5_124_3590_n1671), .Y(DP_OP_102J5_124_3590_n1639) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1026 ( .A1(n172), .A2(
        DP_OP_102J5_124_3590_n1670), .Y(DP_OP_102J5_124_3590_n1638) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1025 ( .A1(n172), .A2(
        DP_OP_102J5_124_3590_n1669), .Y(DP_OP_102J5_124_3590_n1637) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1024 ( .A1(n172), .A2(
        DP_OP_102J5_124_3590_n1668), .Y(DP_OP_102J5_124_3590_n1636) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1023 ( .A1(n172), .A2(
        DP_OP_102J5_124_3590_n1667), .Y(DP_OP_102J5_124_3590_n1635) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1022 ( .A1(n172), .A2(
        DP_OP_102J5_124_3590_n1666), .Y(DP_OP_102J5_124_3590_n1634) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1021 ( .A1(n172), .A2(
        DP_OP_102J5_124_3590_n1665), .Y(DP_OP_102J5_124_3590_n1633) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1008 ( .A1(n199), .A2(
        DP_OP_102J5_124_3590_n1628), .Y(DP_OP_102J5_124_3590_n1620) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1007 ( .A1(n199), .A2(
        DP_OP_102J5_124_3590_n1627), .Y(DP_OP_102J5_124_3590_n1619) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1006 ( .A1(n199), .A2(
        DP_OP_102J5_124_3590_n1626), .Y(DP_OP_102J5_124_3590_n1618) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1005 ( .A1(n199), .A2(
        DP_OP_102J5_124_3590_n1625), .Y(DP_OP_102J5_124_3590_n1617) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1004 ( .A1(n199), .A2(
        DP_OP_102J5_124_3590_n1624), .Y(DP_OP_102J5_124_3590_n1616) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1003 ( .A1(n199), .A2(
        DP_OP_102J5_124_3590_n1623), .Y(DP_OP_102J5_124_3590_n1615) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1002 ( .A1(n199), .A2(
        DP_OP_102J5_124_3590_n1622), .Y(DP_OP_102J5_124_3590_n1614) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1001 ( .A1(n199), .A2(
        DP_OP_102J5_124_3590_n1621), .Y(DP_OP_102J5_124_3590_n1613) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1000 ( .A1(n198), .A2(
        DP_OP_102J5_124_3590_n1628), .Y(DP_OP_102J5_124_3590_n1612) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U999 ( .A1(n198), .A2(
        DP_OP_102J5_124_3590_n1627), .Y(DP_OP_102J5_124_3590_n1611) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U998 ( .A1(n198), .A2(
        DP_OP_102J5_124_3590_n1626), .Y(DP_OP_102J5_124_3590_n1610) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U997 ( .A1(n198), .A2(
        DP_OP_102J5_124_3590_n1625), .Y(DP_OP_102J5_124_3590_n1609) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U996 ( .A1(n198), .A2(
        DP_OP_102J5_124_3590_n1624), .Y(DP_OP_102J5_124_3590_n1608) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U995 ( .A1(n198), .A2(
        DP_OP_102J5_124_3590_n1623), .Y(DP_OP_102J5_124_3590_n1607) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U994 ( .A1(n198), .A2(
        DP_OP_102J5_124_3590_n1622), .Y(DP_OP_102J5_124_3590_n1606) );
  OR2X1_HVT DP_OP_102J5_124_3590_U993 ( .A1(n198), .A2(
        DP_OP_102J5_124_3590_n1621), .Y(DP_OP_102J5_124_3590_n1605) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U992 ( .A1(n197), .A2(
        DP_OP_102J5_124_3590_n1628), .Y(DP_OP_102J5_124_3590_n1604) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U991 ( .A1(n197), .A2(
        DP_OP_102J5_124_3590_n1627), .Y(DP_OP_102J5_124_3590_n1603) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U990 ( .A1(n197), .A2(
        DP_OP_102J5_124_3590_n1626), .Y(DP_OP_102J5_124_3590_n1602) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U989 ( .A1(n197), .A2(
        DP_OP_102J5_124_3590_n1625), .Y(DP_OP_102J5_124_3590_n1601) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U988 ( .A1(n197), .A2(
        DP_OP_102J5_124_3590_n1624), .Y(DP_OP_102J5_124_3590_n1600) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U987 ( .A1(n197), .A2(
        DP_OP_102J5_124_3590_n1623), .Y(DP_OP_102J5_124_3590_n1599) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U986 ( .A1(n197), .A2(
        DP_OP_102J5_124_3590_n1622), .Y(DP_OP_102J5_124_3590_n1598) );
  OR2X1_HVT DP_OP_102J5_124_3590_U985 ( .A1(n197), .A2(
        DP_OP_102J5_124_3590_n1621), .Y(DP_OP_102J5_124_3590_n1597) );
  OR2X1_HVT DP_OP_102J5_124_3590_U984 ( .A1(n171), .A2(
        DP_OP_102J5_124_3590_n1628), .Y(DP_OP_102J5_124_3590_n1596) );
  OR2X1_HVT DP_OP_102J5_124_3590_U983 ( .A1(n171), .A2(
        DP_OP_102J5_124_3590_n1627), .Y(DP_OP_102J5_124_3590_n1595) );
  OR2X1_HVT DP_OP_102J5_124_3590_U982 ( .A1(n171), .A2(
        DP_OP_102J5_124_3590_n1626), .Y(DP_OP_102J5_124_3590_n1594) );
  OR2X1_HVT DP_OP_102J5_124_3590_U981 ( .A1(n171), .A2(
        DP_OP_102J5_124_3590_n1625), .Y(DP_OP_102J5_124_3590_n1593) );
  OR2X1_HVT DP_OP_102J5_124_3590_U980 ( .A1(n171), .A2(
        DP_OP_102J5_124_3590_n1624), .Y(DP_OP_102J5_124_3590_n1592) );
  OR2X1_HVT DP_OP_102J5_124_3590_U979 ( .A1(n171), .A2(
        DP_OP_102J5_124_3590_n1623), .Y(DP_OP_102J5_124_3590_n1591) );
  OR2X1_HVT DP_OP_102J5_124_3590_U978 ( .A1(n171), .A2(
        DP_OP_102J5_124_3590_n1622), .Y(DP_OP_102J5_124_3590_n1590) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U977 ( .A1(n171), .A2(
        DP_OP_102J5_124_3590_n1621), .Y(DP_OP_102J5_124_3590_n1589) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U964 ( .A1(n196), .A2(
        DP_OP_102J5_124_3590_n1584), .Y(DP_OP_102J5_124_3590_n1576) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U963 ( .A1(n196), .A2(
        DP_OP_102J5_124_3590_n1583), .Y(DP_OP_102J5_124_3590_n1575) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U962 ( .A1(n196), .A2(
        DP_OP_102J5_124_3590_n1582), .Y(DP_OP_102J5_124_3590_n1574) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U961 ( .A1(n196), .A2(
        DP_OP_102J5_124_3590_n1581), .Y(DP_OP_102J5_124_3590_n1573) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U960 ( .A1(n196), .A2(
        DP_OP_102J5_124_3590_n1580), .Y(DP_OP_102J5_124_3590_n1572) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U959 ( .A1(n196), .A2(
        DP_OP_102J5_124_3590_n1579), .Y(DP_OP_102J5_124_3590_n1571) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U958 ( .A1(n196), .A2(
        DP_OP_102J5_124_3590_n1578), .Y(DP_OP_102J5_124_3590_n1570) );
  OR2X1_HVT DP_OP_102J5_124_3590_U957 ( .A1(n196), .A2(
        DP_OP_102J5_124_3590_n1577), .Y(DP_OP_102J5_124_3590_n1569) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U956 ( .A1(n195), .A2(
        DP_OP_102J5_124_3590_n1584), .Y(DP_OP_102J5_124_3590_n1568) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U955 ( .A1(n195), .A2(
        DP_OP_102J5_124_3590_n1583), .Y(DP_OP_102J5_124_3590_n1567) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U954 ( .A1(n195), .A2(
        DP_OP_102J5_124_3590_n1582), .Y(DP_OP_102J5_124_3590_n1566) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U953 ( .A1(n195), .A2(
        DP_OP_102J5_124_3590_n1581), .Y(DP_OP_102J5_124_3590_n1565) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U952 ( .A1(n195), .A2(
        DP_OP_102J5_124_3590_n1580), .Y(DP_OP_102J5_124_3590_n1564) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U951 ( .A1(n195), .A2(
        DP_OP_102J5_124_3590_n1579), .Y(DP_OP_102J5_124_3590_n1563) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U950 ( .A1(n195), .A2(
        DP_OP_102J5_124_3590_n1578), .Y(DP_OP_102J5_124_3590_n1562) );
  OR2X1_HVT DP_OP_102J5_124_3590_U949 ( .A1(n195), .A2(
        DP_OP_102J5_124_3590_n1577), .Y(DP_OP_102J5_124_3590_n1561) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U948 ( .A1(n194), .A2(
        DP_OP_102J5_124_3590_n1584), .Y(DP_OP_102J5_124_3590_n1560) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U947 ( .A1(n194), .A2(
        DP_OP_102J5_124_3590_n1583), .Y(DP_OP_102J5_124_3590_n1559) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U946 ( .A1(n194), .A2(
        DP_OP_102J5_124_3590_n1582), .Y(DP_OP_102J5_124_3590_n1558) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U945 ( .A1(n194), .A2(
        DP_OP_102J5_124_3590_n1581), .Y(DP_OP_102J5_124_3590_n1557) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U944 ( .A1(n194), .A2(
        DP_OP_102J5_124_3590_n1580), .Y(DP_OP_102J5_124_3590_n1556) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U943 ( .A1(n194), .A2(
        DP_OP_102J5_124_3590_n1579), .Y(DP_OP_102J5_124_3590_n1555) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U942 ( .A1(n194), .A2(
        DP_OP_102J5_124_3590_n1578), .Y(DP_OP_102J5_124_3590_n1554) );
  OR2X1_HVT DP_OP_102J5_124_3590_U941 ( .A1(n194), .A2(
        DP_OP_102J5_124_3590_n1577), .Y(DP_OP_102J5_124_3590_n1553) );
  OR2X1_HVT DP_OP_102J5_124_3590_U940 ( .A1(n170), .A2(
        DP_OP_102J5_124_3590_n1584), .Y(DP_OP_102J5_124_3590_n1552) );
  OR2X1_HVT DP_OP_102J5_124_3590_U939 ( .A1(n170), .A2(
        DP_OP_102J5_124_3590_n1583), .Y(DP_OP_102J5_124_3590_n1551) );
  OR2X1_HVT DP_OP_102J5_124_3590_U938 ( .A1(n170), .A2(
        DP_OP_102J5_124_3590_n1582), .Y(DP_OP_102J5_124_3590_n1550) );
  OR2X1_HVT DP_OP_102J5_124_3590_U937 ( .A1(n170), .A2(
        DP_OP_102J5_124_3590_n1581), .Y(DP_OP_102J5_124_3590_n1549) );
  OR2X1_HVT DP_OP_102J5_124_3590_U936 ( .A1(n170), .A2(
        DP_OP_102J5_124_3590_n1580), .Y(DP_OP_102J5_124_3590_n1548) );
  OR2X1_HVT DP_OP_102J5_124_3590_U935 ( .A1(n170), .A2(
        DP_OP_102J5_124_3590_n1579), .Y(DP_OP_102J5_124_3590_n1547) );
  OR2X1_HVT DP_OP_102J5_124_3590_U934 ( .A1(n170), .A2(
        DP_OP_102J5_124_3590_n1578), .Y(DP_OP_102J5_124_3590_n1546) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U933 ( .A1(n170), .A2(
        DP_OP_102J5_124_3590_n1577), .Y(DP_OP_102J5_124_3590_n1545) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U920 ( .A1(n193), .A2(
        DP_OP_102J5_124_3590_n1540), .Y(DP_OP_102J5_124_3590_n1532) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U919 ( .A1(n193), .A2(
        DP_OP_102J5_124_3590_n1539), .Y(DP_OP_102J5_124_3590_n1531) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U918 ( .A1(n193), .A2(
        DP_OP_102J5_124_3590_n1538), .Y(DP_OP_102J5_124_3590_n1530) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U917 ( .A1(n193), .A2(
        DP_OP_102J5_124_3590_n1537), .Y(DP_OP_102J5_124_3590_n1529) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U916 ( .A1(n193), .A2(
        DP_OP_102J5_124_3590_n1536), .Y(DP_OP_102J5_124_3590_n1528) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U915 ( .A1(n193), .A2(
        DP_OP_102J5_124_3590_n1535), .Y(DP_OP_102J5_124_3590_n1527) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U914 ( .A1(n193), .A2(
        DP_OP_102J5_124_3590_n1534), .Y(DP_OP_102J5_124_3590_n1526) );
  OR2X1_HVT DP_OP_102J5_124_3590_U913 ( .A1(n193), .A2(
        DP_OP_102J5_124_3590_n1533), .Y(DP_OP_102J5_124_3590_n1525) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U912 ( .A1(n192), .A2(
        DP_OP_102J5_124_3590_n1540), .Y(DP_OP_102J5_124_3590_n1524) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U911 ( .A1(n192), .A2(
        DP_OP_102J5_124_3590_n1539), .Y(DP_OP_102J5_124_3590_n1523) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U910 ( .A1(n192), .A2(
        DP_OP_102J5_124_3590_n1538), .Y(DP_OP_102J5_124_3590_n1522) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U909 ( .A1(n192), .A2(
        DP_OP_102J5_124_3590_n1537), .Y(DP_OP_102J5_124_3590_n1521) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U908 ( .A1(n192), .A2(
        DP_OP_102J5_124_3590_n1536), .Y(DP_OP_102J5_124_3590_n1520) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U907 ( .A1(n192), .A2(
        DP_OP_102J5_124_3590_n1535), .Y(DP_OP_102J5_124_3590_n1519) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U906 ( .A1(n192), .A2(
        DP_OP_102J5_124_3590_n1534), .Y(DP_OP_102J5_124_3590_n1518) );
  OR2X1_HVT DP_OP_102J5_124_3590_U905 ( .A1(n192), .A2(
        DP_OP_102J5_124_3590_n1533), .Y(DP_OP_102J5_124_3590_n1517) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U904 ( .A1(n191), .A2(
        DP_OP_102J5_124_3590_n1540), .Y(DP_OP_102J5_124_3590_n1516) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U903 ( .A1(n191), .A2(
        DP_OP_102J5_124_3590_n1539), .Y(DP_OP_102J5_124_3590_n1515) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U902 ( .A1(n191), .A2(
        DP_OP_102J5_124_3590_n1538), .Y(DP_OP_102J5_124_3590_n1514) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U901 ( .A1(n191), .A2(
        DP_OP_102J5_124_3590_n1537), .Y(DP_OP_102J5_124_3590_n1513) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U900 ( .A1(n191), .A2(
        DP_OP_102J5_124_3590_n1536), .Y(DP_OP_102J5_124_3590_n1512) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U899 ( .A1(n191), .A2(
        DP_OP_102J5_124_3590_n1535), .Y(DP_OP_102J5_124_3590_n1511) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U898 ( .A1(n191), .A2(
        DP_OP_102J5_124_3590_n1534), .Y(DP_OP_102J5_124_3590_n1510) );
  OR2X1_HVT DP_OP_102J5_124_3590_U897 ( .A1(n191), .A2(
        DP_OP_102J5_124_3590_n1533), .Y(DP_OP_102J5_124_3590_n1509) );
  OR2X1_HVT DP_OP_102J5_124_3590_U896 ( .A1(n169), .A2(
        DP_OP_102J5_124_3590_n1540), .Y(DP_OP_102J5_124_3590_n1508) );
  OR2X1_HVT DP_OP_102J5_124_3590_U895 ( .A1(n169), .A2(
        DP_OP_102J5_124_3590_n1539), .Y(DP_OP_102J5_124_3590_n1507) );
  OR2X1_HVT DP_OP_102J5_124_3590_U894 ( .A1(n169), .A2(
        DP_OP_102J5_124_3590_n1538), .Y(DP_OP_102J5_124_3590_n1506) );
  OR2X1_HVT DP_OP_102J5_124_3590_U893 ( .A1(n169), .A2(
        DP_OP_102J5_124_3590_n1537), .Y(DP_OP_102J5_124_3590_n1505) );
  OR2X1_HVT DP_OP_102J5_124_3590_U892 ( .A1(n169), .A2(
        DP_OP_102J5_124_3590_n1536), .Y(DP_OP_102J5_124_3590_n1504) );
  OR2X1_HVT DP_OP_102J5_124_3590_U891 ( .A1(n169), .A2(
        DP_OP_102J5_124_3590_n1535), .Y(DP_OP_102J5_124_3590_n1503) );
  OR2X1_HVT DP_OP_102J5_124_3590_U890 ( .A1(n169), .A2(
        DP_OP_102J5_124_3590_n1534), .Y(DP_OP_102J5_124_3590_n1502) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U889 ( .A1(n169), .A2(
        DP_OP_102J5_124_3590_n1533), .Y(DP_OP_102J5_124_3590_n1501) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U876 ( .A1(n190), .A2(
        DP_OP_102J5_124_3590_n1496), .Y(DP_OP_102J5_124_3590_n1488) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U875 ( .A1(n190), .A2(
        DP_OP_102J5_124_3590_n1495), .Y(DP_OP_102J5_124_3590_n1487) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U874 ( .A1(n190), .A2(
        DP_OP_102J5_124_3590_n1494), .Y(DP_OP_102J5_124_3590_n1486) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U873 ( .A1(n190), .A2(
        DP_OP_102J5_124_3590_n1493), .Y(DP_OP_102J5_124_3590_n1485) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U872 ( .A1(n190), .A2(
        DP_OP_102J5_124_3590_n1492), .Y(DP_OP_102J5_124_3590_n1484) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U871 ( .A1(n190), .A2(
        DP_OP_102J5_124_3590_n1491), .Y(DP_OP_102J5_124_3590_n1483) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U870 ( .A1(n190), .A2(
        DP_OP_102J5_124_3590_n1490), .Y(DP_OP_102J5_124_3590_n1482) );
  OR2X1_HVT DP_OP_102J5_124_3590_U869 ( .A1(n190), .A2(
        DP_OP_102J5_124_3590_n1489), .Y(DP_OP_102J5_124_3590_n1481) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U868 ( .A1(n189), .A2(
        DP_OP_102J5_124_3590_n1496), .Y(DP_OP_102J5_124_3590_n1480) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U867 ( .A1(n189), .A2(
        DP_OP_102J5_124_3590_n1495), .Y(DP_OP_102J5_124_3590_n1479) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U866 ( .A1(n189), .A2(
        DP_OP_102J5_124_3590_n1494), .Y(DP_OP_102J5_124_3590_n1478) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U865 ( .A1(n189), .A2(
        DP_OP_102J5_124_3590_n1493), .Y(DP_OP_102J5_124_3590_n1477) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U864 ( .A1(n189), .A2(
        DP_OP_102J5_124_3590_n1492), .Y(DP_OP_102J5_124_3590_n1476) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U863 ( .A1(n189), .A2(
        DP_OP_102J5_124_3590_n1491), .Y(DP_OP_102J5_124_3590_n1475) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U862 ( .A1(n189), .A2(
        DP_OP_102J5_124_3590_n1490), .Y(DP_OP_102J5_124_3590_n1474) );
  OR2X1_HVT DP_OP_102J5_124_3590_U861 ( .A1(n189), .A2(
        DP_OP_102J5_124_3590_n1489), .Y(DP_OP_102J5_124_3590_n1473) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U860 ( .A1(n188), .A2(
        DP_OP_102J5_124_3590_n1496), .Y(DP_OP_102J5_124_3590_n1472) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U859 ( .A1(n188), .A2(
        DP_OP_102J5_124_3590_n1495), .Y(DP_OP_102J5_124_3590_n1471) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U858 ( .A1(n188), .A2(
        DP_OP_102J5_124_3590_n1494), .Y(DP_OP_102J5_124_3590_n1470) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U857 ( .A1(n188), .A2(
        DP_OP_102J5_124_3590_n1493), .Y(DP_OP_102J5_124_3590_n1469) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U856 ( .A1(n188), .A2(
        DP_OP_102J5_124_3590_n1492), .Y(DP_OP_102J5_124_3590_n1468) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U855 ( .A1(n188), .A2(
        DP_OP_102J5_124_3590_n1491), .Y(DP_OP_102J5_124_3590_n1467) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U854 ( .A1(n188), .A2(
        DP_OP_102J5_124_3590_n1490), .Y(DP_OP_102J5_124_3590_n1466) );
  OR2X1_HVT DP_OP_102J5_124_3590_U853 ( .A1(n188), .A2(
        DP_OP_102J5_124_3590_n1489), .Y(DP_OP_102J5_124_3590_n1465) );
  OR2X1_HVT DP_OP_102J5_124_3590_U852 ( .A1(n168), .A2(
        DP_OP_102J5_124_3590_n1496), .Y(DP_OP_102J5_124_3590_n1464) );
  OR2X1_HVT DP_OP_102J5_124_3590_U851 ( .A1(n168), .A2(
        DP_OP_102J5_124_3590_n1495), .Y(DP_OP_102J5_124_3590_n1463) );
  OR2X1_HVT DP_OP_102J5_124_3590_U850 ( .A1(n168), .A2(
        DP_OP_102J5_124_3590_n1494), .Y(DP_OP_102J5_124_3590_n1462) );
  OR2X1_HVT DP_OP_102J5_124_3590_U849 ( .A1(n168), .A2(
        DP_OP_102J5_124_3590_n1493), .Y(DP_OP_102J5_124_3590_n1461) );
  OR2X1_HVT DP_OP_102J5_124_3590_U848 ( .A1(n168), .A2(
        DP_OP_102J5_124_3590_n1492), .Y(DP_OP_102J5_124_3590_n1460) );
  OR2X1_HVT DP_OP_102J5_124_3590_U847 ( .A1(n168), .A2(
        DP_OP_102J5_124_3590_n1491), .Y(DP_OP_102J5_124_3590_n1459) );
  OR2X1_HVT DP_OP_102J5_124_3590_U846 ( .A1(n168), .A2(
        DP_OP_102J5_124_3590_n1490), .Y(DP_OP_102J5_124_3590_n1458) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U845 ( .A1(n168), .A2(
        DP_OP_102J5_124_3590_n1489), .Y(DP_OP_102J5_124_3590_n1457) );
  FADDX1_HVT DP_OP_102J5_124_3590_U797 ( .A(DP_OP_102J5_124_3590_n1532), .B(
        DP_OP_102J5_124_3590_n1488), .CI(DP_OP_102J5_124_3590_n1576), .CO(
        DP_OP_102J5_124_3590_n1416), .S(DP_OP_102J5_124_3590_n1417) );
  FADDX1_HVT DP_OP_102J5_124_3590_U796 ( .A(DP_OP_102J5_124_3590_n1664), .B(
        DP_OP_102J5_124_3590_n1620), .CI(DP_OP_102J5_124_3590_n1708), .CO(
        DP_OP_102J5_124_3590_n1414), .S(DP_OP_102J5_124_3590_n1415) );
  FADDX1_HVT DP_OP_102J5_124_3590_U795 ( .A(DP_OP_102J5_124_3590_n1795), .B(
        DP_OP_102J5_124_3590_n1752), .CI(DP_OP_102J5_124_3590_n1839), .CO(
        DP_OP_102J5_124_3590_n1412), .S(DP_OP_102J5_124_3590_n1413) );
  FADDX1_HVT DP_OP_102J5_124_3590_U794 ( .A(DP_OP_102J5_124_3590_n1927), .B(
        DP_OP_102J5_124_3590_n1883), .CI(DP_OP_102J5_124_3590_n1971), .CO(
        DP_OP_102J5_124_3590_n1410), .S(DP_OP_102J5_124_3590_n1411) );
  FADDX1_HVT DP_OP_102J5_124_3590_U793 ( .A(DP_OP_102J5_124_3590_n2059), .B(
        DP_OP_102J5_124_3590_n2015), .CI(DP_OP_102J5_124_3590_n2103), .CO(
        DP_OP_102J5_124_3590_n1408), .S(DP_OP_102J5_124_3590_n1409) );
  FADDX1_HVT DP_OP_102J5_124_3590_U792 ( .A(DP_OP_102J5_124_3590_n2322), .B(
        DP_OP_102J5_124_3590_n2147), .CI(DP_OP_102J5_124_3590_n2191), .CO(
        DP_OP_102J5_124_3590_n1406), .S(DP_OP_102J5_124_3590_n1407) );
  FADDX1_HVT DP_OP_102J5_124_3590_U791 ( .A(DP_OP_102J5_124_3590_n2279), .B(
        DP_OP_102J5_124_3590_n2235), .CI(DP_OP_102J5_124_3590_n1411), .CO(
        DP_OP_102J5_124_3590_n1404), .S(DP_OP_102J5_124_3590_n1405) );
  FADDX1_HVT DP_OP_102J5_124_3590_U790 ( .A(DP_OP_102J5_124_3590_n1407), .B(
        DP_OP_102J5_124_3590_n1413), .CI(DP_OP_102J5_124_3590_n1415), .CO(
        DP_OP_102J5_124_3590_n1402), .S(DP_OP_102J5_124_3590_n1403) );
  FADDX1_HVT DP_OP_102J5_124_3590_U789 ( .A(DP_OP_102J5_124_3590_n1409), .B(
        DP_OP_102J5_124_3590_n1417), .CI(DP_OP_102J5_124_3590_n1432), .CO(
        DP_OP_102J5_124_3590_n1400), .S(DP_OP_102J5_124_3590_n1401) );
  FADDX1_HVT DP_OP_102J5_124_3590_U788 ( .A(DP_OP_102J5_124_3590_n1487), .B(
        DP_OP_102J5_124_3590_n1480), .CI(DP_OP_102J5_124_3590_n1524), .CO(
        DP_OP_102J5_124_3590_n1398), .S(DP_OP_102J5_124_3590_n1399) );
  FADDX1_HVT DP_OP_102J5_124_3590_U787 ( .A(DP_OP_102J5_124_3590_n1568), .B(
        DP_OP_102J5_124_3590_n1531), .CI(DP_OP_102J5_124_3590_n1575), .CO(
        DP_OP_102J5_124_3590_n1396), .S(DP_OP_102J5_124_3590_n1397) );
  FADDX1_HVT DP_OP_102J5_124_3590_U786 ( .A(DP_OP_102J5_124_3590_n1619), .B(
        DP_OP_102J5_124_3590_n1612), .CI(DP_OP_102J5_124_3590_n1656), .CO(
        DP_OP_102J5_124_3590_n1394), .S(DP_OP_102J5_124_3590_n1395) );
  FADDX1_HVT DP_OP_102J5_124_3590_U785 ( .A(DP_OP_102J5_124_3590_n1700), .B(
        DP_OP_102J5_124_3590_n1663), .CI(DP_OP_102J5_124_3590_n1707), .CO(
        DP_OP_102J5_124_3590_n1392), .S(DP_OP_102J5_124_3590_n1393) );
  FADDX1_HVT DP_OP_102J5_124_3590_U784 ( .A(DP_OP_102J5_124_3590_n1751), .B(
        DP_OP_102J5_124_3590_n1744), .CI(DP_OP_102J5_124_3590_n1787), .CO(
        DP_OP_102J5_124_3590_n1390), .S(DP_OP_102J5_124_3590_n1391) );
  FADDX1_HVT DP_OP_102J5_124_3590_U783 ( .A(DP_OP_102J5_124_3590_n1831), .B(
        DP_OP_102J5_124_3590_n1794), .CI(DP_OP_102J5_124_3590_n1838), .CO(
        DP_OP_102J5_124_3590_n1388), .S(DP_OP_102J5_124_3590_n1389) );
  FADDX1_HVT DP_OP_102J5_124_3590_U782 ( .A(DP_OP_102J5_124_3590_n1882), .B(
        DP_OP_102J5_124_3590_n1875), .CI(DP_OP_102J5_124_3590_n1919), .CO(
        DP_OP_102J5_124_3590_n1386), .S(DP_OP_102J5_124_3590_n1387) );
  FADDX1_HVT DP_OP_102J5_124_3590_U781 ( .A(DP_OP_102J5_124_3590_n1963), .B(
        DP_OP_102J5_124_3590_n1926), .CI(DP_OP_102J5_124_3590_n2321), .CO(
        DP_OP_102J5_124_3590_n1384), .S(DP_OP_102J5_124_3590_n1385) );
  FADDX1_HVT DP_OP_102J5_124_3590_U780 ( .A(DP_OP_102J5_124_3590_n2315), .B(
        DP_OP_102J5_124_3590_n1970), .CI(DP_OP_102J5_124_3590_n2007), .CO(
        DP_OP_102J5_124_3590_n1382), .S(DP_OP_102J5_124_3590_n1383) );
  FADDX1_HVT DP_OP_102J5_124_3590_U779 ( .A(DP_OP_102J5_124_3590_n2146), .B(
        DP_OP_102J5_124_3590_n2278), .CI(DP_OP_102J5_124_3590_n2271), .CO(
        DP_OP_102J5_124_3590_n1380), .S(DP_OP_102J5_124_3590_n1381) );
  FADDX1_HVT DP_OP_102J5_124_3590_U778 ( .A(DP_OP_102J5_124_3590_n2234), .B(
        DP_OP_102J5_124_3590_n2014), .CI(DP_OP_102J5_124_3590_n2051), .CO(
        DP_OP_102J5_124_3590_n1378), .S(DP_OP_102J5_124_3590_n1379) );
  FADDX1_HVT DP_OP_102J5_124_3590_U777 ( .A(DP_OP_102J5_124_3590_n2227), .B(
        DP_OP_102J5_124_3590_n2058), .CI(DP_OP_102J5_124_3590_n2095), .CO(
        DP_OP_102J5_124_3590_n1376), .S(DP_OP_102J5_124_3590_n1377) );
  FADDX1_HVT DP_OP_102J5_124_3590_U776 ( .A(DP_OP_102J5_124_3590_n2190), .B(
        DP_OP_102J5_124_3590_n2102), .CI(DP_OP_102J5_124_3590_n2139), .CO(
        DP_OP_102J5_124_3590_n1374), .S(DP_OP_102J5_124_3590_n1375) );
  FADDX1_HVT DP_OP_102J5_124_3590_U775 ( .A(DP_OP_102J5_124_3590_n2183), .B(
        DP_OP_102J5_124_3590_n1408), .CI(DP_OP_102J5_124_3590_n1406), .CO(
        DP_OP_102J5_124_3590_n1372), .S(DP_OP_102J5_124_3590_n1373) );
  FADDX1_HVT DP_OP_102J5_124_3590_U774 ( .A(DP_OP_102J5_124_3590_n1414), .B(
        DP_OP_102J5_124_3590_n1410), .CI(DP_OP_102J5_124_3590_n1412), .CO(
        DP_OP_102J5_124_3590_n1370), .S(DP_OP_102J5_124_3590_n1371) );
  FADDX1_HVT DP_OP_102J5_124_3590_U773 ( .A(DP_OP_102J5_124_3590_n1416), .B(
        DP_OP_102J5_124_3590_n1377), .CI(DP_OP_102J5_124_3590_n1379), .CO(
        DP_OP_102J5_124_3590_n1368), .S(DP_OP_102J5_124_3590_n1369) );
  FADDX1_HVT DP_OP_102J5_124_3590_U772 ( .A(DP_OP_102J5_124_3590_n1375), .B(
        DP_OP_102J5_124_3590_n1389), .CI(DP_OP_102J5_124_3590_n1391), .CO(
        DP_OP_102J5_124_3590_n1366), .S(DP_OP_102J5_124_3590_n1367) );
  FADDX1_HVT DP_OP_102J5_124_3590_U771 ( .A(DP_OP_102J5_124_3590_n1381), .B(
        DP_OP_102J5_124_3590_n1395), .CI(DP_OP_102J5_124_3590_n1393), .CO(
        DP_OP_102J5_124_3590_n1364), .S(DP_OP_102J5_124_3590_n1365) );
  FADDX1_HVT DP_OP_102J5_124_3590_U770 ( .A(DP_OP_102J5_124_3590_n1383), .B(
        DP_OP_102J5_124_3590_n1399), .CI(DP_OP_102J5_124_3590_n1397), .CO(
        DP_OP_102J5_124_3590_n1362), .S(DP_OP_102J5_124_3590_n1363) );
  FADDX1_HVT DP_OP_102J5_124_3590_U769 ( .A(DP_OP_102J5_124_3590_n1385), .B(
        DP_OP_102J5_124_3590_n1387), .CI(DP_OP_102J5_124_3590_n1431), .CO(
        DP_OP_102J5_124_3590_n1360), .S(DP_OP_102J5_124_3590_n1361) );
  FADDX1_HVT DP_OP_102J5_124_3590_U768 ( .A(DP_OP_102J5_124_3590_n1404), .B(
        DP_OP_102J5_124_3590_n1373), .CI(DP_OP_102J5_124_3590_n1402), .CO(
        DP_OP_102J5_124_3590_n1358), .S(DP_OP_102J5_124_3590_n1359) );
  FADDX1_HVT DP_OP_102J5_124_3590_U767 ( .A(DP_OP_102J5_124_3590_n1371), .B(
        DP_OP_102J5_124_3590_n1369), .CI(DP_OP_102J5_124_3590_n1363), .CO(
        DP_OP_102J5_124_3590_n1356), .S(DP_OP_102J5_124_3590_n1357) );
  FADDX1_HVT DP_OP_102J5_124_3590_U766 ( .A(DP_OP_102J5_124_3590_n1367), .B(
        DP_OP_102J5_124_3590_n1365), .CI(DP_OP_102J5_124_3590_n1400), .CO(
        DP_OP_102J5_124_3590_n1354), .S(DP_OP_102J5_124_3590_n1355) );
  FADDX1_HVT DP_OP_102J5_124_3590_U765 ( .A(DP_OP_102J5_124_3590_n1361), .B(
        DP_OP_102J5_124_3590_n1359), .CI(DP_OP_102J5_124_3590_n1357), .CO(
        DP_OP_102J5_124_3590_n1352), .S(DP_OP_102J5_124_3590_n1353) );
  HADDX1_HVT DP_OP_102J5_124_3590_U764 ( .A0(DP_OP_102J5_124_3590_n1479), .B0(
        DP_OP_102J5_124_3590_n1486), .C1(DP_OP_102J5_124_3590_n1350), .SO(
        DP_OP_102J5_124_3590_n1351) );
  FADDX1_HVT DP_OP_102J5_124_3590_U763 ( .A(DP_OP_102J5_124_3590_n1516), .B(
        DP_OP_102J5_124_3590_n1472), .CI(DP_OP_102J5_124_3590_n1523), .CO(
        DP_OP_102J5_124_3590_n1348), .S(DP_OP_102J5_124_3590_n1349) );
  FADDX1_HVT DP_OP_102J5_124_3590_U762 ( .A(DP_OP_102J5_124_3590_n1560), .B(
        DP_OP_102J5_124_3590_n1530), .CI(DP_OP_102J5_124_3590_n1567), .CO(
        DP_OP_102J5_124_3590_n1346), .S(DP_OP_102J5_124_3590_n1347) );
  FADDX1_HVT DP_OP_102J5_124_3590_U761 ( .A(DP_OP_102J5_124_3590_n1604), .B(
        DP_OP_102J5_124_3590_n1574), .CI(DP_OP_102J5_124_3590_n1611), .CO(
        DP_OP_102J5_124_3590_n1344), .S(DP_OP_102J5_124_3590_n1345) );
  FADDX1_HVT DP_OP_102J5_124_3590_U760 ( .A(DP_OP_102J5_124_3590_n1648), .B(
        DP_OP_102J5_124_3590_n1618), .CI(DP_OP_102J5_124_3590_n1655), .CO(
        DP_OP_102J5_124_3590_n1342), .S(DP_OP_102J5_124_3590_n1343) );
  FADDX1_HVT DP_OP_102J5_124_3590_U759 ( .A(DP_OP_102J5_124_3590_n1692), .B(
        DP_OP_102J5_124_3590_n1662), .CI(DP_OP_102J5_124_3590_n1699), .CO(
        DP_OP_102J5_124_3590_n1340), .S(DP_OP_102J5_124_3590_n1341) );
  FADDX1_HVT DP_OP_102J5_124_3590_U758 ( .A(DP_OP_102J5_124_3590_n1736), .B(
        DP_OP_102J5_124_3590_n1706), .CI(DP_OP_102J5_124_3590_n1743), .CO(
        DP_OP_102J5_124_3590_n1338), .S(DP_OP_102J5_124_3590_n1339) );
  FADDX1_HVT DP_OP_102J5_124_3590_U757 ( .A(DP_OP_102J5_124_3590_n1779), .B(
        DP_OP_102J5_124_3590_n1750), .CI(DP_OP_102J5_124_3590_n1786), .CO(
        DP_OP_102J5_124_3590_n1336), .S(DP_OP_102J5_124_3590_n1337) );
  FADDX1_HVT DP_OP_102J5_124_3590_U756 ( .A(DP_OP_102J5_124_3590_n1823), .B(
        DP_OP_102J5_124_3590_n1793), .CI(DP_OP_102J5_124_3590_n1830), .CO(
        DP_OP_102J5_124_3590_n1334), .S(DP_OP_102J5_124_3590_n1335) );
  FADDX1_HVT DP_OP_102J5_124_3590_U755 ( .A(DP_OP_102J5_124_3590_n2057), .B(
        DP_OP_102J5_124_3590_n2320), .CI(DP_OP_102J5_124_3590_n2314), .CO(
        DP_OP_102J5_124_3590_n1332), .S(DP_OP_102J5_124_3590_n1333) );
  FADDX1_HVT DP_OP_102J5_124_3590_U754 ( .A(DP_OP_102J5_124_3590_n2043), .B(
        DP_OP_102J5_124_3590_n2307), .CI(DP_OP_102J5_124_3590_n2277), .CO(
        DP_OP_102J5_124_3590_n1330), .S(DP_OP_102J5_124_3590_n1331) );
  FADDX1_HVT DP_OP_102J5_124_3590_U753 ( .A(DP_OP_102J5_124_3590_n2013), .B(
        DP_OP_102J5_124_3590_n1837), .CI(DP_OP_102J5_124_3590_n1867), .CO(
        DP_OP_102J5_124_3590_n1328), .S(DP_OP_102J5_124_3590_n1329) );
  FADDX1_HVT DP_OP_102J5_124_3590_U752 ( .A(DP_OP_102J5_124_3590_n2050), .B(
        DP_OP_102J5_124_3590_n1874), .CI(DP_OP_102J5_124_3590_n1881), .CO(
        DP_OP_102J5_124_3590_n1326), .S(DP_OP_102J5_124_3590_n1327) );
  FADDX1_HVT DP_OP_102J5_124_3590_U751 ( .A(DP_OP_102J5_124_3590_n2087), .B(
        DP_OP_102J5_124_3590_n1911), .CI(DP_OP_102J5_124_3590_n1918), .CO(
        DP_OP_102J5_124_3590_n1324), .S(DP_OP_102J5_124_3590_n1325) );
  FADDX1_HVT DP_OP_102J5_124_3590_U750 ( .A(DP_OP_102J5_124_3590_n2101), .B(
        DP_OP_102J5_124_3590_n1925), .CI(DP_OP_102J5_124_3590_n2270), .CO(
        DP_OP_102J5_124_3590_n1322), .S(DP_OP_102J5_124_3590_n1323) );
  FADDX1_HVT DP_OP_102J5_124_3590_U749 ( .A(DP_OP_102J5_124_3590_n2094), .B(
        DP_OP_102J5_124_3590_n2263), .CI(DP_OP_102J5_124_3590_n2233), .CO(
        DP_OP_102J5_124_3590_n1320), .S(DP_OP_102J5_124_3590_n1321) );
  FADDX1_HVT DP_OP_102J5_124_3590_U748 ( .A(DP_OP_102J5_124_3590_n2226), .B(
        DP_OP_102J5_124_3590_n1955), .CI(DP_OP_102J5_124_3590_n1962), .CO(
        DP_OP_102J5_124_3590_n1318), .S(DP_OP_102J5_124_3590_n1319) );
  FADDX1_HVT DP_OP_102J5_124_3590_U747 ( .A(DP_OP_102J5_124_3590_n2219), .B(
        DP_OP_102J5_124_3590_n1969), .CI(DP_OP_102J5_124_3590_n1999), .CO(
        DP_OP_102J5_124_3590_n1316), .S(DP_OP_102J5_124_3590_n1317) );
  FADDX1_HVT DP_OP_102J5_124_3590_U746 ( .A(DP_OP_102J5_124_3590_n2189), .B(
        DP_OP_102J5_124_3590_n2006), .CI(DP_OP_102J5_124_3590_n2182), .CO(
        DP_OP_102J5_124_3590_n1314), .S(DP_OP_102J5_124_3590_n1315) );
  FADDX1_HVT DP_OP_102J5_124_3590_U745 ( .A(DP_OP_102J5_124_3590_n2175), .B(
        DP_OP_102J5_124_3590_n2131), .CI(DP_OP_102J5_124_3590_n2138), .CO(
        DP_OP_102J5_124_3590_n1312), .S(DP_OP_102J5_124_3590_n1313) );
  FADDX1_HVT DP_OP_102J5_124_3590_U744 ( .A(DP_OP_102J5_124_3590_n2145), .B(
        DP_OP_102J5_124_3590_n1351), .CI(DP_OP_102J5_124_3590_n1376), .CO(
        DP_OP_102J5_124_3590_n1310), .S(DP_OP_102J5_124_3590_n1311) );
  FADDX1_HVT DP_OP_102J5_124_3590_U743 ( .A(DP_OP_102J5_124_3590_n1378), .B(
        DP_OP_102J5_124_3590_n1380), .CI(DP_OP_102J5_124_3590_n1382), .CO(
        DP_OP_102J5_124_3590_n1308), .S(DP_OP_102J5_124_3590_n1309) );
  FADDX1_HVT DP_OP_102J5_124_3590_U742 ( .A(DP_OP_102J5_124_3590_n1392), .B(
        DP_OP_102J5_124_3590_n1384), .CI(DP_OP_102J5_124_3590_n1374), .CO(
        DP_OP_102J5_124_3590_n1306), .S(DP_OP_102J5_124_3590_n1307) );
  FADDX1_HVT DP_OP_102J5_124_3590_U741 ( .A(DP_OP_102J5_124_3590_n1390), .B(
        DP_OP_102J5_124_3590_n1386), .CI(DP_OP_102J5_124_3590_n1388), .CO(
        DP_OP_102J5_124_3590_n1304), .S(DP_OP_102J5_124_3590_n1305) );
  FADDX1_HVT DP_OP_102J5_124_3590_U740 ( .A(DP_OP_102J5_124_3590_n1394), .B(
        DP_OP_102J5_124_3590_n1396), .CI(DP_OP_102J5_124_3590_n1398), .CO(
        DP_OP_102J5_124_3590_n1302), .S(DP_OP_102J5_124_3590_n1303) );
  FADDX1_HVT DP_OP_102J5_124_3590_U739 ( .A(DP_OP_102J5_124_3590_n1327), .B(
        DP_OP_102J5_124_3590_n1339), .CI(DP_OP_102J5_124_3590_n1337), .CO(
        DP_OP_102J5_124_3590_n1300), .S(DP_OP_102J5_124_3590_n1301) );
  FADDX1_HVT DP_OP_102J5_124_3590_U738 ( .A(DP_OP_102J5_124_3590_n1317), .B(
        DP_OP_102J5_124_3590_n1331), .CI(DP_OP_102J5_124_3590_n1329), .CO(
        DP_OP_102J5_124_3590_n1298), .S(DP_OP_102J5_124_3590_n1299) );
  FADDX1_HVT DP_OP_102J5_124_3590_U737 ( .A(DP_OP_102J5_124_3590_n1315), .B(
        DP_OP_102J5_124_3590_n1341), .CI(DP_OP_102J5_124_3590_n1335), .CO(
        DP_OP_102J5_124_3590_n1296), .S(DP_OP_102J5_124_3590_n1297) );
  FADDX1_HVT DP_OP_102J5_124_3590_U736 ( .A(DP_OP_102J5_124_3590_n1321), .B(
        DP_OP_102J5_124_3590_n1343), .CI(DP_OP_102J5_124_3590_n1345), .CO(
        DP_OP_102J5_124_3590_n1294), .S(DP_OP_102J5_124_3590_n1295) );
  FADDX1_HVT DP_OP_102J5_124_3590_U735 ( .A(DP_OP_102J5_124_3590_n1319), .B(
        DP_OP_102J5_124_3590_n1349), .CI(DP_OP_102J5_124_3590_n1347), .CO(
        DP_OP_102J5_124_3590_n1292), .S(DP_OP_102J5_124_3590_n1293) );
  FADDX1_HVT DP_OP_102J5_124_3590_U734 ( .A(DP_OP_102J5_124_3590_n1325), .B(
        DP_OP_102J5_124_3590_n1323), .CI(DP_OP_102J5_124_3590_n1313), .CO(
        DP_OP_102J5_124_3590_n1290), .S(DP_OP_102J5_124_3590_n1291) );
  FADDX1_HVT DP_OP_102J5_124_3590_U733 ( .A(DP_OP_102J5_124_3590_n1333), .B(
        DP_OP_102J5_124_3590_n1372), .CI(DP_OP_102J5_124_3590_n1370), .CO(
        DP_OP_102J5_124_3590_n1288), .S(DP_OP_102J5_124_3590_n1289) );
  FADDX1_HVT DP_OP_102J5_124_3590_U732 ( .A(DP_OP_102J5_124_3590_n1430), .B(
        DP_OP_102J5_124_3590_n1311), .CI(DP_OP_102J5_124_3590_n1368), .CO(
        DP_OP_102J5_124_3590_n1286), .S(DP_OP_102J5_124_3590_n1287) );
  FADDX1_HVT DP_OP_102J5_124_3590_U731 ( .A(DP_OP_102J5_124_3590_n1305), .B(
        DP_OP_102J5_124_3590_n1303), .CI(DP_OP_102J5_124_3590_n1307), .CO(
        DP_OP_102J5_124_3590_n1284), .S(DP_OP_102J5_124_3590_n1285) );
  FADDX1_HVT DP_OP_102J5_124_3590_U730 ( .A(DP_OP_102J5_124_3590_n1366), .B(
        DP_OP_102J5_124_3590_n1309), .CI(DP_OP_102J5_124_3590_n1364), .CO(
        DP_OP_102J5_124_3590_n1282), .S(DP_OP_102J5_124_3590_n1283) );
  FADDX1_HVT DP_OP_102J5_124_3590_U729 ( .A(DP_OP_102J5_124_3590_n1362), .B(
        DP_OP_102J5_124_3590_n1291), .CI(DP_OP_102J5_124_3590_n1293), .CO(
        DP_OP_102J5_124_3590_n1280), .S(DP_OP_102J5_124_3590_n1281) );
  FADDX1_HVT DP_OP_102J5_124_3590_U728 ( .A(DP_OP_102J5_124_3590_n1295), .B(
        DP_OP_102J5_124_3590_n1301), .CI(DP_OP_102J5_124_3590_n1360), .CO(
        DP_OP_102J5_124_3590_n1278), .S(DP_OP_102J5_124_3590_n1279) );
  FADDX1_HVT DP_OP_102J5_124_3590_U727 ( .A(DP_OP_102J5_124_3590_n1299), .B(
        DP_OP_102J5_124_3590_n1297), .CI(DP_OP_102J5_124_3590_n1358), .CO(
        DP_OP_102J5_124_3590_n1276), .S(DP_OP_102J5_124_3590_n1277) );
  FADDX1_HVT DP_OP_102J5_124_3590_U726 ( .A(DP_OP_102J5_124_3590_n1289), .B(
        DP_OP_102J5_124_3590_n1287), .CI(DP_OP_102J5_124_3590_n1356), .CO(
        DP_OP_102J5_124_3590_n1274), .S(DP_OP_102J5_124_3590_n1275) );
  FADDX1_HVT DP_OP_102J5_124_3590_U725 ( .A(DP_OP_102J5_124_3590_n1354), .B(
        DP_OP_102J5_124_3590_n1285), .CI(DP_OP_102J5_124_3590_n1283), .CO(
        DP_OP_102J5_124_3590_n1272), .S(DP_OP_102J5_124_3590_n1273) );
  FADDX1_HVT DP_OP_102J5_124_3590_U724 ( .A(DP_OP_102J5_124_3590_n1281), .B(
        DP_OP_102J5_124_3590_n1279), .CI(DP_OP_102J5_124_3590_n1277), .CO(
        DP_OP_102J5_124_3590_n1270), .S(DP_OP_102J5_124_3590_n1271) );
  FADDX1_HVT DP_OP_102J5_124_3590_U723 ( .A(DP_OP_102J5_124_3590_n1352), .B(
        DP_OP_102J5_124_3590_n1275), .CI(DP_OP_102J5_124_3590_n1273), .CO(
        DP_OP_102J5_124_3590_n1268), .S(DP_OP_102J5_124_3590_n1269) );
  HADDX1_HVT DP_OP_102J5_124_3590_U722 ( .A0(DP_OP_102J5_124_3590_n1640), .B0(
        DP_OP_102J5_124_3590_n1464), .C1(DP_OP_102J5_124_3590_n1266), .SO(
        DP_OP_102J5_124_3590_n1267) );
  FADDX1_HVT DP_OP_102J5_124_3590_U721 ( .A(DP_OP_102J5_124_3590_n2123), .B(
        DP_OP_102J5_124_3590_n1771), .CI(DP_OP_102J5_124_3590_n1903), .CO(
        DP_OP_102J5_124_3590_n1264), .S(DP_OP_102J5_124_3590_n1265) );
  FADDX1_HVT DP_OP_102J5_124_3590_U720 ( .A(DP_OP_102J5_124_3590_n2035), .B(
        DP_OP_102J5_124_3590_n1991), .CI(DP_OP_102J5_124_3590_n2167), .CO(
        DP_OP_102J5_124_3590_n1262), .S(DP_OP_102J5_124_3590_n1263) );
  FADDX1_HVT DP_OP_102J5_124_3590_U719 ( .A(DP_OP_102J5_124_3590_n1815), .B(
        DP_OP_102J5_124_3590_n1947), .CI(DP_OP_102J5_124_3590_n1596), .CO(
        DP_OP_102J5_124_3590_n1260), .S(DP_OP_102J5_124_3590_n1261) );
  FADDX1_HVT DP_OP_102J5_124_3590_U718 ( .A(DP_OP_102J5_124_3590_n1552), .B(
        DP_OP_102J5_124_3590_n1859), .CI(DP_OP_102J5_124_3590_n2255), .CO(
        DP_OP_102J5_124_3590_n1258), .S(DP_OP_102J5_124_3590_n1259) );
  FADDX1_HVT DP_OP_102J5_124_3590_U717 ( .A(DP_OP_102J5_124_3590_n1728), .B(
        DP_OP_102J5_124_3590_n2079), .CI(DP_OP_102J5_124_3590_n2299), .CO(
        DP_OP_102J5_124_3590_n1256), .S(DP_OP_102J5_124_3590_n1257) );
  FADDX1_HVT DP_OP_102J5_124_3590_U716 ( .A(DP_OP_102J5_124_3590_n1508), .B(
        DP_OP_102J5_124_3590_n1684), .CI(DP_OP_102J5_124_3590_n2211), .CO(
        DP_OP_102J5_124_3590_n1254), .S(DP_OP_102J5_124_3590_n1255) );
  FADDX1_HVT DP_OP_102J5_124_3590_U715 ( .A(DP_OP_102J5_124_3590_n1485), .B(
        DP_OP_102J5_124_3590_n1471), .CI(DP_OP_102J5_124_3590_n1478), .CO(
        DP_OP_102J5_124_3590_n1252), .S(DP_OP_102J5_124_3590_n1253) );
  FADDX1_HVT DP_OP_102J5_124_3590_U714 ( .A(DP_OP_102J5_124_3590_n1522), .B(
        DP_OP_102J5_124_3590_n1515), .CI(DP_OP_102J5_124_3590_n1529), .CO(
        DP_OP_102J5_124_3590_n1250), .S(DP_OP_102J5_124_3590_n1251) );
  FADDX1_HVT DP_OP_102J5_124_3590_U713 ( .A(DP_OP_102J5_124_3590_n1566), .B(
        DP_OP_102J5_124_3590_n1559), .CI(DP_OP_102J5_124_3590_n1573), .CO(
        DP_OP_102J5_124_3590_n1248), .S(DP_OP_102J5_124_3590_n1249) );
  FADDX1_HVT DP_OP_102J5_124_3590_U712 ( .A(DP_OP_102J5_124_3590_n2319), .B(
        DP_OP_102J5_124_3590_n1603), .CI(DP_OP_102J5_124_3590_n2313), .CO(
        DP_OP_102J5_124_3590_n1246), .S(DP_OP_102J5_124_3590_n1247) );
  FADDX1_HVT DP_OP_102J5_124_3590_U711 ( .A(DP_OP_102J5_124_3590_n1917), .B(
        DP_OP_102J5_124_3590_n2306), .CI(DP_OP_102J5_124_3590_n1610), .CO(
        DP_OP_102J5_124_3590_n1244), .S(DP_OP_102J5_124_3590_n1245) );
  FADDX1_HVT DP_OP_102J5_124_3590_U710 ( .A(DP_OP_102J5_124_3590_n1910), .B(
        DP_OP_102J5_124_3590_n2276), .CI(DP_OP_102J5_124_3590_n2269), .CO(
        DP_OP_102J5_124_3590_n1242), .S(DP_OP_102J5_124_3590_n1243) );
  FADDX1_HVT DP_OP_102J5_124_3590_U709 ( .A(DP_OP_102J5_124_3590_n1873), .B(
        DP_OP_102J5_124_3590_n1617), .CI(DP_OP_102J5_124_3590_n2262), .CO(
        DP_OP_102J5_124_3590_n1240), .S(DP_OP_102J5_124_3590_n1241) );
  FADDX1_HVT DP_OP_102J5_124_3590_U708 ( .A(DP_OP_102J5_124_3590_n1880), .B(
        DP_OP_102J5_124_3590_n2232), .CI(DP_OP_102J5_124_3590_n1647), .CO(
        DP_OP_102J5_124_3590_n1238), .S(DP_OP_102J5_124_3590_n1239) );
  FADDX1_HVT DP_OP_102J5_124_3590_U707 ( .A(DP_OP_102J5_124_3590_n2225), .B(
        DP_OP_102J5_124_3590_n1654), .CI(DP_OP_102J5_124_3590_n2218), .CO(
        DP_OP_102J5_124_3590_n1236), .S(DP_OP_102J5_124_3590_n1237) );
  FADDX1_HVT DP_OP_102J5_124_3590_U706 ( .A(DP_OP_102J5_124_3590_n1836), .B(
        DP_OP_102J5_124_3590_n2188), .CI(DP_OP_102J5_124_3590_n1661), .CO(
        DP_OP_102J5_124_3590_n1234), .S(DP_OP_102J5_124_3590_n1235) );
  FADDX1_HVT DP_OP_102J5_124_3590_U705 ( .A(DP_OP_102J5_124_3590_n1866), .B(
        DP_OP_102J5_124_3590_n1691), .CI(DP_OP_102J5_124_3590_n2181), .CO(
        DP_OP_102J5_124_3590_n1232), .S(DP_OP_102J5_124_3590_n1233) );
  FADDX1_HVT DP_OP_102J5_124_3590_U704 ( .A(DP_OP_102J5_124_3590_n1829), .B(
        DP_OP_102J5_124_3590_n1698), .CI(DP_OP_102J5_124_3590_n2174), .CO(
        DP_OP_102J5_124_3590_n1230), .S(DP_OP_102J5_124_3590_n1231) );
  FADDX1_HVT DP_OP_102J5_124_3590_U703 ( .A(DP_OP_102J5_124_3590_n1924), .B(
        DP_OP_102J5_124_3590_n1705), .CI(DP_OP_102J5_124_3590_n2144), .CO(
        DP_OP_102J5_124_3590_n1228), .S(DP_OP_102J5_124_3590_n1229) );
  FADDX1_HVT DP_OP_102J5_124_3590_U702 ( .A(DP_OP_102J5_124_3590_n2137), .B(
        DP_OP_102J5_124_3590_n1735), .CI(DP_OP_102J5_124_3590_n1742), .CO(
        DP_OP_102J5_124_3590_n1226), .S(DP_OP_102J5_124_3590_n1227) );
  FADDX1_HVT DP_OP_102J5_124_3590_U701 ( .A(DP_OP_102J5_124_3590_n1961), .B(
        DP_OP_102J5_124_3590_n2130), .CI(DP_OP_102J5_124_3590_n2100), .CO(
        DP_OP_102J5_124_3590_n1224), .S(DP_OP_102J5_124_3590_n1225) );
  FADDX1_HVT DP_OP_102J5_124_3590_U700 ( .A(DP_OP_102J5_124_3590_n1792), .B(
        DP_OP_102J5_124_3590_n2093), .CI(DP_OP_102J5_124_3590_n2086), .CO(
        DP_OP_102J5_124_3590_n1222), .S(DP_OP_102J5_124_3590_n1223) );
  FADDX1_HVT DP_OP_102J5_124_3590_U699 ( .A(DP_OP_102J5_124_3590_n1778), .B(
        DP_OP_102J5_124_3590_n2056), .CI(DP_OP_102J5_124_3590_n2049), .CO(
        DP_OP_102J5_124_3590_n1220), .S(DP_OP_102J5_124_3590_n1221) );
  FADDX1_HVT DP_OP_102J5_124_3590_U698 ( .A(DP_OP_102J5_124_3590_n1968), .B(
        DP_OP_102J5_124_3590_n2042), .CI(DP_OP_102J5_124_3590_n1749), .CO(
        DP_OP_102J5_124_3590_n1218), .S(DP_OP_102J5_124_3590_n1219) );
  FADDX1_HVT DP_OP_102J5_124_3590_U697 ( .A(DP_OP_102J5_124_3590_n1822), .B(
        DP_OP_102J5_124_3590_n2012), .CI(DP_OP_102J5_124_3590_n2005), .CO(
        DP_OP_102J5_124_3590_n1216), .S(DP_OP_102J5_124_3590_n1217) );
  FADDX1_HVT DP_OP_102J5_124_3590_U696 ( .A(DP_OP_102J5_124_3590_n1998), .B(
        DP_OP_102J5_124_3590_n1785), .CI(DP_OP_102J5_124_3590_n1954), .CO(
        DP_OP_102J5_124_3590_n1214), .S(DP_OP_102J5_124_3590_n1215) );
  FADDX1_HVT DP_OP_102J5_124_3590_U695 ( .A(DP_OP_102J5_124_3590_n1350), .B(
        DP_OP_102J5_124_3590_n1267), .CI(DP_OP_102J5_124_3590_n1312), .CO(
        DP_OP_102J5_124_3590_n1212), .S(DP_OP_102J5_124_3590_n1213) );
  FADDX1_HVT DP_OP_102J5_124_3590_U694 ( .A(DP_OP_102J5_124_3590_n1334), .B(
        DP_OP_102J5_124_3590_n1314), .CI(DP_OP_102J5_124_3590_n1318), .CO(
        DP_OP_102J5_124_3590_n1210), .S(DP_OP_102J5_124_3590_n1211) );
  FADDX1_HVT DP_OP_102J5_124_3590_U693 ( .A(DP_OP_102J5_124_3590_n1332), .B(
        DP_OP_102J5_124_3590_n1320), .CI(DP_OP_102J5_124_3590_n1316), .CO(
        DP_OP_102J5_124_3590_n1208), .S(DP_OP_102J5_124_3590_n1209) );
  FADDX1_HVT DP_OP_102J5_124_3590_U692 ( .A(DP_OP_102J5_124_3590_n1336), .B(
        DP_OP_102J5_124_3590_n1322), .CI(DP_OP_102J5_124_3590_n1326), .CO(
        DP_OP_102J5_124_3590_n1206), .S(DP_OP_102J5_124_3590_n1207) );
  FADDX1_HVT DP_OP_102J5_124_3590_U691 ( .A(DP_OP_102J5_124_3590_n1330), .B(
        DP_OP_102J5_124_3590_n1324), .CI(DP_OP_102J5_124_3590_n1328), .CO(
        DP_OP_102J5_124_3590_n1204), .S(DP_OP_102J5_124_3590_n1205) );
  FADDX1_HVT DP_OP_102J5_124_3590_U690 ( .A(DP_OP_102J5_124_3590_n1340), .B(
        DP_OP_102J5_124_3590_n1342), .CI(DP_OP_102J5_124_3590_n1344), .CO(
        DP_OP_102J5_124_3590_n1202), .S(DP_OP_102J5_124_3590_n1203) );
  FADDX1_HVT DP_OP_102J5_124_3590_U689 ( .A(DP_OP_102J5_124_3590_n1346), .B(
        DP_OP_102J5_124_3590_n1348), .CI(DP_OP_102J5_124_3590_n1338), .CO(
        DP_OP_102J5_124_3590_n1200), .S(DP_OP_102J5_124_3590_n1201) );
  FADDX1_HVT DP_OP_102J5_124_3590_U688 ( .A(DP_OP_102J5_124_3590_n1259), .B(
        DP_OP_102J5_124_3590_n1261), .CI(DP_OP_102J5_124_3590_n1265), .CO(
        DP_OP_102J5_124_3590_n1198), .S(DP_OP_102J5_124_3590_n1199) );
  FADDX1_HVT DP_OP_102J5_124_3590_U687 ( .A(DP_OP_102J5_124_3590_n1263), .B(
        DP_OP_102J5_124_3590_n1255), .CI(DP_OP_102J5_124_3590_n1257), .CO(
        DP_OP_102J5_124_3590_n1196), .S(DP_OP_102J5_124_3590_n1197) );
  FADDX1_HVT DP_OP_102J5_124_3590_U686 ( .A(DP_OP_102J5_124_3590_n1219), .B(
        DP_OP_102J5_124_3590_n1247), .CI(DP_OP_102J5_124_3590_n1249), .CO(
        DP_OP_102J5_124_3590_n1194), .S(DP_OP_102J5_124_3590_n1195) );
  FADDX1_HVT DP_OP_102J5_124_3590_U685 ( .A(DP_OP_102J5_124_3590_n1217), .B(
        DP_OP_102J5_124_3590_n1241), .CI(DP_OP_102J5_124_3590_n1243), .CO(
        DP_OP_102J5_124_3590_n1192), .S(DP_OP_102J5_124_3590_n1193) );
  FADDX1_HVT DP_OP_102J5_124_3590_U684 ( .A(DP_OP_102J5_124_3590_n1239), .B(
        DP_OP_102J5_124_3590_n1245), .CI(DP_OP_102J5_124_3590_n1237), .CO(
        DP_OP_102J5_124_3590_n1190), .S(DP_OP_102J5_124_3590_n1191) );
  FADDX1_HVT DP_OP_102J5_124_3590_U683 ( .A(DP_OP_102J5_124_3590_n1215), .B(
        DP_OP_102J5_124_3590_n1253), .CI(DP_OP_102J5_124_3590_n1233), .CO(
        DP_OP_102J5_124_3590_n1188), .S(DP_OP_102J5_124_3590_n1189) );
  FADDX1_HVT DP_OP_102J5_124_3590_U682 ( .A(DP_OP_102J5_124_3590_n1235), .B(
        DP_OP_102J5_124_3590_n1221), .CI(DP_OP_102J5_124_3590_n1227), .CO(
        DP_OP_102J5_124_3590_n1186), .S(DP_OP_102J5_124_3590_n1187) );
  FADDX1_HVT DP_OP_102J5_124_3590_U681 ( .A(DP_OP_102J5_124_3590_n1229), .B(
        DP_OP_102J5_124_3590_n1251), .CI(DP_OP_102J5_124_3590_n1231), .CO(
        DP_OP_102J5_124_3590_n1184), .S(DP_OP_102J5_124_3590_n1185) );
  FADDX1_HVT DP_OP_102J5_124_3590_U680 ( .A(DP_OP_102J5_124_3590_n1223), .B(
        DP_OP_102J5_124_3590_n1225), .CI(DP_OP_102J5_124_3590_n1310), .CO(
        DP_OP_102J5_124_3590_n1182), .S(DP_OP_102J5_124_3590_n1183) );
  FADDX1_HVT DP_OP_102J5_124_3590_U679 ( .A(DP_OP_102J5_124_3590_n1302), .B(
        DP_OP_102J5_124_3590_n1304), .CI(DP_OP_102J5_124_3590_n1429), .CO(
        DP_OP_102J5_124_3590_n1180), .S(DP_OP_102J5_124_3590_n1181) );
  FADDX1_HVT DP_OP_102J5_124_3590_U678 ( .A(DP_OP_102J5_124_3590_n1308), .B(
        DP_OP_102J5_124_3590_n1306), .CI(DP_OP_102J5_124_3590_n1213), .CO(
        DP_OP_102J5_124_3590_n1178), .S(DP_OP_102J5_124_3590_n1179) );
  FADDX1_HVT DP_OP_102J5_124_3590_U677 ( .A(DP_OP_102J5_124_3590_n1203), .B(
        DP_OP_102J5_124_3590_n1201), .CI(DP_OP_102J5_124_3590_n1205), .CO(
        DP_OP_102J5_124_3590_n1176), .S(DP_OP_102J5_124_3590_n1177) );
  FADDX1_HVT DP_OP_102J5_124_3590_U676 ( .A(DP_OP_102J5_124_3590_n1207), .B(
        DP_OP_102J5_124_3590_n1209), .CI(DP_OP_102J5_124_3590_n1211), .CO(
        DP_OP_102J5_124_3590_n1174), .S(DP_OP_102J5_124_3590_n1175) );
  FADDX1_HVT DP_OP_102J5_124_3590_U675 ( .A(DP_OP_102J5_124_3590_n1300), .B(
        DP_OP_102J5_124_3590_n1290), .CI(DP_OP_102J5_124_3590_n1292), .CO(
        DP_OP_102J5_124_3590_n1172), .S(DP_OP_102J5_124_3590_n1173) );
  FADDX1_HVT DP_OP_102J5_124_3590_U674 ( .A(DP_OP_102J5_124_3590_n1294), .B(
        DP_OP_102J5_124_3590_n1298), .CI(DP_OP_102J5_124_3590_n1296), .CO(
        DP_OP_102J5_124_3590_n1170), .S(DP_OP_102J5_124_3590_n1171) );
  FADDX1_HVT DP_OP_102J5_124_3590_U673 ( .A(DP_OP_102J5_124_3590_n1197), .B(
        DP_OP_102J5_124_3590_n1199), .CI(DP_OP_102J5_124_3590_n1187), .CO(
        DP_OP_102J5_124_3590_n1168), .S(DP_OP_102J5_124_3590_n1169) );
  FADDX1_HVT DP_OP_102J5_124_3590_U672 ( .A(DP_OP_102J5_124_3590_n1193), .B(
        DP_OP_102J5_124_3590_n1195), .CI(DP_OP_102J5_124_3590_n1288), .CO(
        DP_OP_102J5_124_3590_n1166), .S(DP_OP_102J5_124_3590_n1167) );
  FADDX1_HVT DP_OP_102J5_124_3590_U671 ( .A(DP_OP_102J5_124_3590_n1191), .B(
        DP_OP_102J5_124_3590_n1189), .CI(DP_OP_102J5_124_3590_n1185), .CO(
        DP_OP_102J5_124_3590_n1164), .S(DP_OP_102J5_124_3590_n1165) );
  FADDX1_HVT DP_OP_102J5_124_3590_U670 ( .A(DP_OP_102J5_124_3590_n1183), .B(
        DP_OP_102J5_124_3590_n1286), .CI(DP_OP_102J5_124_3590_n1282), .CO(
        DP_OP_102J5_124_3590_n1162), .S(DP_OP_102J5_124_3590_n1163) );
  FADDX1_HVT DP_OP_102J5_124_3590_U669 ( .A(DP_OP_102J5_124_3590_n1284), .B(
        DP_OP_102J5_124_3590_n1181), .CI(DP_OP_102J5_124_3590_n1179), .CO(
        DP_OP_102J5_124_3590_n1160), .S(DP_OP_102J5_124_3590_n1161) );
  FADDX1_HVT DP_OP_102J5_124_3590_U668 ( .A(DP_OP_102J5_124_3590_n1280), .B(
        DP_OP_102J5_124_3590_n1278), .CI(DP_OP_102J5_124_3590_n1173), .CO(
        DP_OP_102J5_124_3590_n1158), .S(DP_OP_102J5_124_3590_n1159) );
  FADDX1_HVT DP_OP_102J5_124_3590_U667 ( .A(DP_OP_102J5_124_3590_n1175), .B(
        DP_OP_102J5_124_3590_n1177), .CI(DP_OP_102J5_124_3590_n1171), .CO(
        DP_OP_102J5_124_3590_n1156), .S(DP_OP_102J5_124_3590_n1157) );
  FADDX1_HVT DP_OP_102J5_124_3590_U666 ( .A(DP_OP_102J5_124_3590_n1169), .B(
        DP_OP_102J5_124_3590_n1276), .CI(DP_OP_102J5_124_3590_n1165), .CO(
        DP_OP_102J5_124_3590_n1154), .S(DP_OP_102J5_124_3590_n1155) );
  FADDX1_HVT DP_OP_102J5_124_3590_U665 ( .A(DP_OP_102J5_124_3590_n1167), .B(
        DP_OP_102J5_124_3590_n1274), .CI(DP_OP_102J5_124_3590_n1163), .CO(
        DP_OP_102J5_124_3590_n1152), .S(DP_OP_102J5_124_3590_n1153) );
  FADDX1_HVT DP_OP_102J5_124_3590_U664 ( .A(DP_OP_102J5_124_3590_n1272), .B(
        DP_OP_102J5_124_3590_n1161), .CI(DP_OP_102J5_124_3590_n1159), .CO(
        DP_OP_102J5_124_3590_n1150), .S(DP_OP_102J5_124_3590_n1151) );
  FADDX1_HVT DP_OP_102J5_124_3590_U663 ( .A(DP_OP_102J5_124_3590_n1157), .B(
        DP_OP_102J5_124_3590_n1270), .CI(DP_OP_102J5_124_3590_n1155), .CO(
        DP_OP_102J5_124_3590_n1148), .S(DP_OP_102J5_124_3590_n1149) );
  FADDX1_HVT DP_OP_102J5_124_3590_U662 ( .A(DP_OP_102J5_124_3590_n1153), .B(
        DP_OP_102J5_124_3590_n1268), .CI(DP_OP_102J5_124_3590_n1151), .CO(
        DP_OP_102J5_124_3590_n1146), .S(DP_OP_102J5_124_3590_n1147) );
  FADDX1_HVT DP_OP_102J5_124_3590_U661 ( .A(DP_OP_102J5_124_3590_n1639), .B(
        DP_OP_102J5_124_3590_n1990), .CI(DP_OP_102J5_124_3590_n1463), .CO(
        DP_OP_102J5_124_3590_n1144), .S(DP_OP_102J5_124_3590_n1145) );
  FADDX1_HVT DP_OP_102J5_124_3590_U660 ( .A(DP_OP_102J5_124_3590_n2122), .B(
        DP_OP_102J5_124_3590_n2166), .CI(DP_OP_102J5_124_3590_n1683), .CO(
        DP_OP_102J5_124_3590_n1142), .S(DP_OP_102J5_124_3590_n1143) );
  FADDX1_HVT DP_OP_102J5_124_3590_U659 ( .A(DP_OP_102J5_124_3590_n2254), .B(
        DP_OP_102J5_124_3590_n1770), .CI(DP_OP_102J5_124_3590_n1814), .CO(
        DP_OP_102J5_124_3590_n1140), .S(DP_OP_102J5_124_3590_n1141) );
  FADDX1_HVT DP_OP_102J5_124_3590_U658 ( .A(DP_OP_102J5_124_3590_n2298), .B(
        DP_OP_102J5_124_3590_n1858), .CI(DP_OP_102J5_124_3590_n1727), .CO(
        DP_OP_102J5_124_3590_n1138), .S(DP_OP_102J5_124_3590_n1139) );
  FADDX1_HVT DP_OP_102J5_124_3590_U657 ( .A(DP_OP_102J5_124_3590_n1946), .B(
        DP_OP_102J5_124_3590_n1551), .CI(DP_OP_102J5_124_3590_n2210), .CO(
        DP_OP_102J5_124_3590_n1136), .S(DP_OP_102J5_124_3590_n1137) );
  FADDX1_HVT DP_OP_102J5_124_3590_U656 ( .A(DP_OP_102J5_124_3590_n2078), .B(
        DP_OP_102J5_124_3590_n2034), .CI(DP_OP_102J5_124_3590_n1595), .CO(
        DP_OP_102J5_124_3590_n1134), .S(DP_OP_102J5_124_3590_n1135) );
  FADDX1_HVT DP_OP_102J5_124_3590_U655 ( .A(DP_OP_102J5_124_3590_n1902), .B(
        DP_OP_102J5_124_3590_n1507), .CI(DP_OP_102J5_124_3590_n1916), .CO(
        DP_OP_102J5_124_3590_n1132), .S(DP_OP_102J5_124_3590_n1133) );
  FADDX1_HVT DP_OP_102J5_124_3590_U654 ( .A(DP_OP_102J5_124_3590_n1909), .B(
        DP_OP_102J5_124_3590_n1477), .CI(DP_OP_102J5_124_3590_n1470), .CO(
        DP_OP_102J5_124_3590_n1130), .S(DP_OP_102J5_124_3590_n1131) );
  FADDX1_HVT DP_OP_102J5_124_3590_U653 ( .A(DP_OP_102J5_124_3590_n2318), .B(
        DP_OP_102J5_124_3590_n1484), .CI(DP_OP_102J5_124_3590_n1514), .CO(
        DP_OP_102J5_124_3590_n1128), .S(DP_OP_102J5_124_3590_n1129) );
  FADDX1_HVT DP_OP_102J5_124_3590_U652 ( .A(DP_OP_102J5_124_3590_n1828), .B(
        DP_OP_102J5_124_3590_n1521), .CI(DP_OP_102J5_124_3590_n2312), .CO(
        DP_OP_102J5_124_3590_n1126), .S(DP_OP_102J5_124_3590_n1127) );
  FADDX1_HVT DP_OP_102J5_124_3590_U651 ( .A(DP_OP_102J5_124_3590_n2305), .B(
        DP_OP_102J5_124_3590_n1528), .CI(DP_OP_102J5_124_3590_n1558), .CO(
        DP_OP_102J5_124_3590_n1124), .S(DP_OP_102J5_124_3590_n1125) );
  FADDX1_HVT DP_OP_102J5_124_3590_U650 ( .A(DP_OP_102J5_124_3590_n1821), .B(
        DP_OP_102J5_124_3590_n1565), .CI(DP_OP_102J5_124_3590_n2275), .CO(
        DP_OP_102J5_124_3590_n1122), .S(DP_OP_102J5_124_3590_n1123) );
  FADDX1_HVT DP_OP_102J5_124_3590_U649 ( .A(DP_OP_102J5_124_3590_n1835), .B(
        DP_OP_102J5_124_3590_n2268), .CI(DP_OP_102J5_124_3590_n1572), .CO(
        DP_OP_102J5_124_3590_n1120), .S(DP_OP_102J5_124_3590_n1121) );
  FADDX1_HVT DP_OP_102J5_124_3590_U648 ( .A(DP_OP_102J5_124_3590_n1865), .B(
        DP_OP_102J5_124_3590_n1602), .CI(DP_OP_102J5_124_3590_n2261), .CO(
        DP_OP_102J5_124_3590_n1118), .S(DP_OP_102J5_124_3590_n1119) );
  FADDX1_HVT DP_OP_102J5_124_3590_U647 ( .A(DP_OP_102J5_124_3590_n1791), .B(
        DP_OP_102J5_124_3590_n2231), .CI(DP_OP_102J5_124_3590_n2224), .CO(
        DP_OP_102J5_124_3590_n1116), .S(DP_OP_102J5_124_3590_n1117) );
  FADDX1_HVT DP_OP_102J5_124_3590_U646 ( .A(DP_OP_102J5_124_3590_n1777), .B(
        DP_OP_102J5_124_3590_n2217), .CI(DP_OP_102J5_124_3590_n2187), .CO(
        DP_OP_102J5_124_3590_n1114), .S(DP_OP_102J5_124_3590_n1115) );
  FADDX1_HVT DP_OP_102J5_124_3590_U645 ( .A(DP_OP_102J5_124_3590_n1748), .B(
        DP_OP_102J5_124_3590_n2180), .CI(DP_OP_102J5_124_3590_n2173), .CO(
        DP_OP_102J5_124_3590_n1112), .S(DP_OP_102J5_124_3590_n1113) );
  FADDX1_HVT DP_OP_102J5_124_3590_U644 ( .A(DP_OP_102J5_124_3590_n1734), .B(
        DP_OP_102J5_124_3590_n1609), .CI(DP_OP_102J5_124_3590_n1616), .CO(
        DP_OP_102J5_124_3590_n1110), .S(DP_OP_102J5_124_3590_n1111) );
  FADDX1_HVT DP_OP_102J5_124_3590_U643 ( .A(DP_OP_102J5_124_3590_n2143), .B(
        DP_OP_102J5_124_3590_n1646), .CI(DP_OP_102J5_124_3590_n1653), .CO(
        DP_OP_102J5_124_3590_n1108), .S(DP_OP_102J5_124_3590_n1109) );
  FADDX1_HVT DP_OP_102J5_124_3590_U642 ( .A(DP_OP_102J5_124_3590_n2136), .B(
        DP_OP_102J5_124_3590_n1660), .CI(DP_OP_102J5_124_3590_n1690), .CO(
        DP_OP_102J5_124_3590_n1106), .S(DP_OP_102J5_124_3590_n1107) );
  FADDX1_HVT DP_OP_102J5_124_3590_U641 ( .A(DP_OP_102J5_124_3590_n2129), .B(
        DP_OP_102J5_124_3590_n1697), .CI(DP_OP_102J5_124_3590_n1704), .CO(
        DP_OP_102J5_124_3590_n1104), .S(DP_OP_102J5_124_3590_n1105) );
  FADDX1_HVT DP_OP_102J5_124_3590_U640 ( .A(DP_OP_102J5_124_3590_n2099), .B(
        DP_OP_102J5_124_3590_n1741), .CI(DP_OP_102J5_124_3590_n1784), .CO(
        DP_OP_102J5_124_3590_n1102), .S(DP_OP_102J5_124_3590_n1103) );
  FADDX1_HVT DP_OP_102J5_124_3590_U639 ( .A(DP_OP_102J5_124_3590_n2092), .B(
        DP_OP_102J5_124_3590_n1872), .CI(DP_OP_102J5_124_3590_n1879), .CO(
        DP_OP_102J5_124_3590_n1100), .S(DP_OP_102J5_124_3590_n1101) );
  FADDX1_HVT DP_OP_102J5_124_3590_U638 ( .A(DP_OP_102J5_124_3590_n2085), .B(
        DP_OP_102J5_124_3590_n1923), .CI(DP_OP_102J5_124_3590_n1953), .CO(
        DP_OP_102J5_124_3590_n1098), .S(DP_OP_102J5_124_3590_n1099) );
  FADDX1_HVT DP_OP_102J5_124_3590_U637 ( .A(DP_OP_102J5_124_3590_n1997), .B(
        DP_OP_102J5_124_3590_n1960), .CI(DP_OP_102J5_124_3590_n2055), .CO(
        DP_OP_102J5_124_3590_n1096), .S(DP_OP_102J5_124_3590_n1097) );
  FADDX1_HVT DP_OP_102J5_124_3590_U636 ( .A(DP_OP_102J5_124_3590_n2048), .B(
        DP_OP_102J5_124_3590_n2041), .CI(DP_OP_102J5_124_3590_n2011), .CO(
        DP_OP_102J5_124_3590_n1094), .S(DP_OP_102J5_124_3590_n1095) );
  FADDX1_HVT DP_OP_102J5_124_3590_U635 ( .A(DP_OP_102J5_124_3590_n2004), .B(
        DP_OP_102J5_124_3590_n1967), .CI(DP_OP_102J5_124_3590_n1266), .CO(
        DP_OP_102J5_124_3590_n1092), .S(DP_OP_102J5_124_3590_n1093) );
  FADDX1_HVT DP_OP_102J5_124_3590_U634 ( .A(DP_OP_102J5_124_3590_n1258), .B(
        DP_OP_102J5_124_3590_n1254), .CI(DP_OP_102J5_124_3590_n1260), .CO(
        DP_OP_102J5_124_3590_n1090), .S(DP_OP_102J5_124_3590_n1091) );
  FADDX1_HVT DP_OP_102J5_124_3590_U633 ( .A(DP_OP_102J5_124_3590_n1264), .B(
        DP_OP_102J5_124_3590_n1256), .CI(DP_OP_102J5_124_3590_n1262), .CO(
        DP_OP_102J5_124_3590_n1088), .S(DP_OP_102J5_124_3590_n1089) );
  FADDX1_HVT DP_OP_102J5_124_3590_U632 ( .A(DP_OP_102J5_124_3590_n1214), .B(
        DP_OP_102J5_124_3590_n1216), .CI(DP_OP_102J5_124_3590_n1220), .CO(
        DP_OP_102J5_124_3590_n1086), .S(DP_OP_102J5_124_3590_n1087) );
  FADDX1_HVT DP_OP_102J5_124_3590_U631 ( .A(DP_OP_102J5_124_3590_n1236), .B(
        DP_OP_102J5_124_3590_n1218), .CI(DP_OP_102J5_124_3590_n1222), .CO(
        DP_OP_102J5_124_3590_n1084), .S(DP_OP_102J5_124_3590_n1085) );
  FADDX1_HVT DP_OP_102J5_124_3590_U630 ( .A(DP_OP_102J5_124_3590_n1238), .B(
        DP_OP_102J5_124_3590_n1224), .CI(DP_OP_102J5_124_3590_n1226), .CO(
        DP_OP_102J5_124_3590_n1082), .S(DP_OP_102J5_124_3590_n1083) );
  FADDX1_HVT DP_OP_102J5_124_3590_U629 ( .A(DP_OP_102J5_124_3590_n1240), .B(
        DP_OP_102J5_124_3590_n1228), .CI(DP_OP_102J5_124_3590_n1230), .CO(
        DP_OP_102J5_124_3590_n1080), .S(DP_OP_102J5_124_3590_n1081) );
  FADDX1_HVT DP_OP_102J5_124_3590_U628 ( .A(DP_OP_102J5_124_3590_n1232), .B(
        DP_OP_102J5_124_3590_n1234), .CI(DP_OP_102J5_124_3590_n1244), .CO(
        DP_OP_102J5_124_3590_n1078), .S(DP_OP_102J5_124_3590_n1079) );
  FADDX1_HVT DP_OP_102J5_124_3590_U627 ( .A(DP_OP_102J5_124_3590_n1248), .B(
        DP_OP_102J5_124_3590_n1242), .CI(DP_OP_102J5_124_3590_n1250), .CO(
        DP_OP_102J5_124_3590_n1076), .S(DP_OP_102J5_124_3590_n1077) );
  FADDX1_HVT DP_OP_102J5_124_3590_U626 ( .A(DP_OP_102J5_124_3590_n1252), .B(
        DP_OP_102J5_124_3590_n1246), .CI(DP_OP_102J5_124_3590_n1139), .CO(
        DP_OP_102J5_124_3590_n1074), .S(DP_OP_102J5_124_3590_n1075) );
  FADDX1_HVT DP_OP_102J5_124_3590_U625 ( .A(DP_OP_102J5_124_3590_n1135), .B(
        DP_OP_102J5_124_3590_n1137), .CI(DP_OP_102J5_124_3590_n1133), .CO(
        DP_OP_102J5_124_3590_n1072), .S(DP_OP_102J5_124_3590_n1073) );
  FADDX1_HVT DP_OP_102J5_124_3590_U624 ( .A(DP_OP_102J5_124_3590_n1143), .B(
        DP_OP_102J5_124_3590_n1141), .CI(DP_OP_102J5_124_3590_n1145), .CO(
        DP_OP_102J5_124_3590_n1070), .S(DP_OP_102J5_124_3590_n1071) );
  FADDX1_HVT DP_OP_102J5_124_3590_U623 ( .A(DP_OP_102J5_124_3590_n1125), .B(
        DP_OP_102J5_124_3590_n1131), .CI(DP_OP_102J5_124_3590_n1129), .CO(
        DP_OP_102J5_124_3590_n1068), .S(DP_OP_102J5_124_3590_n1069) );
  FADDX1_HVT DP_OP_102J5_124_3590_U622 ( .A(DP_OP_102J5_124_3590_n1121), .B(
        DP_OP_102J5_124_3590_n1127), .CI(DP_OP_102J5_124_3590_n1115), .CO(
        DP_OP_102J5_124_3590_n1066), .S(DP_OP_102J5_124_3590_n1067) );
  FADDX1_HVT DP_OP_102J5_124_3590_U621 ( .A(DP_OP_102J5_124_3590_n1113), .B(
        DP_OP_102J5_124_3590_n1109), .CI(DP_OP_102J5_124_3590_n1105), .CO(
        DP_OP_102J5_124_3590_n1064), .S(DP_OP_102J5_124_3590_n1065) );
  FADDX1_HVT DP_OP_102J5_124_3590_U620 ( .A(DP_OP_102J5_124_3590_n1117), .B(
        DP_OP_102J5_124_3590_n1099), .CI(DP_OP_102J5_124_3590_n1097), .CO(
        DP_OP_102J5_124_3590_n1062), .S(DP_OP_102J5_124_3590_n1063) );
  FADDX1_HVT DP_OP_102J5_124_3590_U619 ( .A(DP_OP_102J5_124_3590_n1111), .B(
        DP_OP_102J5_124_3590_n1101), .CI(DP_OP_102J5_124_3590_n1103), .CO(
        DP_OP_102J5_124_3590_n1060), .S(DP_OP_102J5_124_3590_n1061) );
  FADDX1_HVT DP_OP_102J5_124_3590_U618 ( .A(DP_OP_102J5_124_3590_n1107), .B(
        DP_OP_102J5_124_3590_n1123), .CI(DP_OP_102J5_124_3590_n1095), .CO(
        DP_OP_102J5_124_3590_n1058), .S(DP_OP_102J5_124_3590_n1059) );
  FADDX1_HVT DP_OP_102J5_124_3590_U617 ( .A(DP_OP_102J5_124_3590_n1119), .B(
        DP_OP_102J5_124_3590_n1093), .CI(DP_OP_102J5_124_3590_n1212), .CO(
        DP_OP_102J5_124_3590_n1056), .S(DP_OP_102J5_124_3590_n1057) );
  FADDX1_HVT DP_OP_102J5_124_3590_U616 ( .A(DP_OP_102J5_124_3590_n1200), .B(
        DP_OP_102J5_124_3590_n1204), .CI(DP_OP_102J5_124_3590_n1428), .CO(
        DP_OP_102J5_124_3590_n1054), .S(DP_OP_102J5_124_3590_n1055) );
  FADDX1_HVT DP_OP_102J5_124_3590_U615 ( .A(DP_OP_102J5_124_3590_n1210), .B(
        DP_OP_102J5_124_3590_n1208), .CI(DP_OP_102J5_124_3590_n1202), .CO(
        DP_OP_102J5_124_3590_n1052), .S(DP_OP_102J5_124_3590_n1053) );
  FADDX1_HVT DP_OP_102J5_124_3590_U614 ( .A(DP_OP_102J5_124_3590_n1206), .B(
        DP_OP_102J5_124_3590_n1196), .CI(DP_OP_102J5_124_3590_n1198), .CO(
        DP_OP_102J5_124_3590_n1050), .S(DP_OP_102J5_124_3590_n1051) );
  FADDX1_HVT DP_OP_102J5_124_3590_U613 ( .A(DP_OP_102J5_124_3590_n1089), .B(
        DP_OP_102J5_124_3590_n1091), .CI(DP_OP_102J5_124_3590_n1194), .CO(
        DP_OP_102J5_124_3590_n1048), .S(DP_OP_102J5_124_3590_n1049) );
  FADDX1_HVT DP_OP_102J5_124_3590_U612 ( .A(DP_OP_102J5_124_3590_n1083), .B(
        DP_OP_102J5_124_3590_n1192), .CI(DP_OP_102J5_124_3590_n1075), .CO(
        DP_OP_102J5_124_3590_n1046), .S(DP_OP_102J5_124_3590_n1047) );
  FADDX1_HVT DP_OP_102J5_124_3590_U611 ( .A(DP_OP_102J5_124_3590_n1190), .B(
        DP_OP_102J5_124_3590_n1077), .CI(DP_OP_102J5_124_3590_n1085), .CO(
        DP_OP_102J5_124_3590_n1044), .S(DP_OP_102J5_124_3590_n1045) );
  FADDX1_HVT DP_OP_102J5_124_3590_U610 ( .A(DP_OP_102J5_124_3590_n1188), .B(
        DP_OP_102J5_124_3590_n1079), .CI(DP_OP_102J5_124_3590_n1081), .CO(
        DP_OP_102J5_124_3590_n1042), .S(DP_OP_102J5_124_3590_n1043) );
  FADDX1_HVT DP_OP_102J5_124_3590_U609 ( .A(DP_OP_102J5_124_3590_n1186), .B(
        DP_OP_102J5_124_3590_n1087), .CI(DP_OP_102J5_124_3590_n1184), .CO(
        DP_OP_102J5_124_3590_n1040), .S(DP_OP_102J5_124_3590_n1041) );
  FADDX1_HVT DP_OP_102J5_124_3590_U608 ( .A(DP_OP_102J5_124_3590_n1182), .B(
        DP_OP_102J5_124_3590_n1073), .CI(DP_OP_102J5_124_3590_n1071), .CO(
        DP_OP_102J5_124_3590_n1038), .S(DP_OP_102J5_124_3590_n1039) );
  FADDX1_HVT DP_OP_102J5_124_3590_U607 ( .A(DP_OP_102J5_124_3590_n1065), .B(
        DP_OP_102J5_124_3590_n1061), .CI(DP_OP_102J5_124_3590_n1063), .CO(
        DP_OP_102J5_124_3590_n1036), .S(DP_OP_102J5_124_3590_n1037) );
  FADDX1_HVT DP_OP_102J5_124_3590_U606 ( .A(DP_OP_102J5_124_3590_n1059), .B(
        DP_OP_102J5_124_3590_n1069), .CI(DP_OP_102J5_124_3590_n1067), .CO(
        DP_OP_102J5_124_3590_n1034), .S(DP_OP_102J5_124_3590_n1035) );
  FADDX1_HVT DP_OP_102J5_124_3590_U605 ( .A(DP_OP_102J5_124_3590_n1180), .B(
        DP_OP_102J5_124_3590_n1057), .CI(DP_OP_102J5_124_3590_n1178), .CO(
        DP_OP_102J5_124_3590_n1032), .S(DP_OP_102J5_124_3590_n1033) );
  FADDX1_HVT DP_OP_102J5_124_3590_U604 ( .A(DP_OP_102J5_124_3590_n1176), .B(
        DP_OP_102J5_124_3590_n1053), .CI(DP_OP_102J5_124_3590_n1055), .CO(
        DP_OP_102J5_124_3590_n1030), .S(DP_OP_102J5_124_3590_n1031) );
  FADDX1_HVT DP_OP_102J5_124_3590_U603 ( .A(DP_OP_102J5_124_3590_n1174), .B(
        DP_OP_102J5_124_3590_n1170), .CI(DP_OP_102J5_124_3590_n1172), .CO(
        DP_OP_102J5_124_3590_n1028), .S(DP_OP_102J5_124_3590_n1029) );
  FADDX1_HVT DP_OP_102J5_124_3590_U602 ( .A(DP_OP_102J5_124_3590_n1051), .B(
        DP_OP_102J5_124_3590_n1168), .CI(DP_OP_102J5_124_3590_n1049), .CO(
        DP_OP_102J5_124_3590_n1026), .S(DP_OP_102J5_124_3590_n1027) );
  FADDX1_HVT DP_OP_102J5_124_3590_U601 ( .A(DP_OP_102J5_124_3590_n1164), .B(
        DP_OP_102J5_124_3590_n1043), .CI(DP_OP_102J5_124_3590_n1041), .CO(
        DP_OP_102J5_124_3590_n1024), .S(DP_OP_102J5_124_3590_n1025) );
  FADDX1_HVT DP_OP_102J5_124_3590_U600 ( .A(DP_OP_102J5_124_3590_n1166), .B(
        DP_OP_102J5_124_3590_n1047), .CI(DP_OP_102J5_124_3590_n1045), .CO(
        DP_OP_102J5_124_3590_n1022), .S(DP_OP_102J5_124_3590_n1023) );
  FADDX1_HVT DP_OP_102J5_124_3590_U599 ( .A(DP_OP_102J5_124_3590_n1039), .B(
        DP_OP_102J5_124_3590_n1037), .CI(DP_OP_102J5_124_3590_n1035), .CO(
        DP_OP_102J5_124_3590_n1020), .S(DP_OP_102J5_124_3590_n1021) );
  FADDX1_HVT DP_OP_102J5_124_3590_U598 ( .A(DP_OP_102J5_124_3590_n1162), .B(
        DP_OP_102J5_124_3590_n1160), .CI(DP_OP_102J5_124_3590_n1033), .CO(
        DP_OP_102J5_124_3590_n1018), .S(DP_OP_102J5_124_3590_n1019) );
  FADDX1_HVT DP_OP_102J5_124_3590_U597 ( .A(DP_OP_102J5_124_3590_n1158), .B(
        DP_OP_102J5_124_3590_n1156), .CI(DP_OP_102J5_124_3590_n1031), .CO(
        DP_OP_102J5_124_3590_n1016), .S(DP_OP_102J5_124_3590_n1017) );
  FADDX1_HVT DP_OP_102J5_124_3590_U596 ( .A(DP_OP_102J5_124_3590_n1029), .B(
        DP_OP_102J5_124_3590_n1027), .CI(DP_OP_102J5_124_3590_n1154), .CO(
        DP_OP_102J5_124_3590_n1014), .S(DP_OP_102J5_124_3590_n1015) );
  FADDX1_HVT DP_OP_102J5_124_3590_U595 ( .A(DP_OP_102J5_124_3590_n1025), .B(
        DP_OP_102J5_124_3590_n1023), .CI(DP_OP_102J5_124_3590_n1152), .CO(
        DP_OP_102J5_124_3590_n1012), .S(DP_OP_102J5_124_3590_n1013) );
  FADDX1_HVT DP_OP_102J5_124_3590_U594 ( .A(DP_OP_102J5_124_3590_n1021), .B(
        DP_OP_102J5_124_3590_n1019), .CI(DP_OP_102J5_124_3590_n1150), .CO(
        DP_OP_102J5_124_3590_n1010), .S(DP_OP_102J5_124_3590_n1011) );
  FADDX1_HVT DP_OP_102J5_124_3590_U593 ( .A(DP_OP_102J5_124_3590_n1017), .B(
        DP_OP_102J5_124_3590_n1148), .CI(DP_OP_102J5_124_3590_n1015), .CO(
        DP_OP_102J5_124_3590_n1008), .S(DP_OP_102J5_124_3590_n1009) );
  FADDX1_HVT DP_OP_102J5_124_3590_U592 ( .A(DP_OP_102J5_124_3590_n1013), .B(
        DP_OP_102J5_124_3590_n1146), .CI(DP_OP_102J5_124_3590_n1011), .CO(
        DP_OP_102J5_124_3590_n1006), .S(DP_OP_102J5_124_3590_n1007) );
  OR2X1_HVT DP_OP_102J5_124_3590_U591 ( .A1(DP_OP_102J5_124_3590_n2033), .A2(
        DP_OP_102J5_124_3590_n1901), .Y(DP_OP_102J5_124_3590_n1004) );
  FADDX1_HVT DP_OP_102J5_124_3590_U589 ( .A(DP_OP_102J5_124_3590_n2121), .B(
        DP_OP_102J5_124_3590_n1945), .CI(DP_OP_102J5_124_3590_n1462), .CO(
        DP_OP_102J5_124_3590_n1002), .S(DP_OP_102J5_124_3590_n1003) );
  FADDX1_HVT DP_OP_102J5_124_3590_U588 ( .A(DP_OP_102J5_124_3590_n1638), .B(
        DP_OP_102J5_124_3590_n1857), .CI(DP_OP_102J5_124_3590_n1989), .CO(
        DP_OP_102J5_124_3590_n1000), .S(DP_OP_102J5_124_3590_n1001) );
  FADDX1_HVT DP_OP_102J5_124_3590_U587 ( .A(DP_OP_102J5_124_3590_n1506), .B(
        DP_OP_102J5_124_3590_n2209), .CI(DP_OP_102J5_124_3590_n1813), .CO(
        DP_OP_102J5_124_3590_n998), .S(DP_OP_102J5_124_3590_n999) );
  FADDX1_HVT DP_OP_102J5_124_3590_U586 ( .A(DP_OP_102J5_124_3590_n2165), .B(
        DP_OP_102J5_124_3590_n2253), .CI(DP_OP_102J5_124_3590_n1594), .CO(
        DP_OP_102J5_124_3590_n996), .S(DP_OP_102J5_124_3590_n997) );
  FADDX1_HVT DP_OP_102J5_124_3590_U585 ( .A(DP_OP_102J5_124_3590_n1726), .B(
        DP_OP_102J5_124_3590_n1769), .CI(DP_OP_102J5_124_3590_n2297), .CO(
        DP_OP_102J5_124_3590_n994), .S(DP_OP_102J5_124_3590_n995) );
  FADDX1_HVT DP_OP_102J5_124_3590_U584 ( .A(DP_OP_102J5_124_3590_n1550), .B(
        DP_OP_102J5_124_3590_n1682), .CI(DP_OP_102J5_124_3590_n2077), .CO(
        DP_OP_102J5_124_3590_n992), .S(DP_OP_102J5_124_3590_n993) );
  FADDX1_HVT DP_OP_102J5_124_3590_U583 ( .A(DP_OP_102J5_124_3590_n1820), .B(
        DP_OP_102J5_124_3590_n1469), .CI(DP_OP_102J5_124_3590_n1476), .CO(
        DP_OP_102J5_124_3590_n990), .S(DP_OP_102J5_124_3590_n991) );
  FADDX1_HVT DP_OP_102J5_124_3590_U582 ( .A(DP_OP_102J5_124_3590_n1834), .B(
        DP_OP_102J5_124_3590_n2317), .CI(DP_OP_102J5_124_3590_n2311), .CO(
        DP_OP_102J5_124_3590_n988), .S(DP_OP_102J5_124_3590_n989) );
  FADDX1_HVT DP_OP_102J5_124_3590_U581 ( .A(DP_OP_102J5_124_3590_n1790), .B(
        DP_OP_102J5_124_3590_n2304), .CI(DP_OP_102J5_124_3590_n2274), .CO(
        DP_OP_102J5_124_3590_n986), .S(DP_OP_102J5_124_3590_n987) );
  FADDX1_HVT DP_OP_102J5_124_3590_U580 ( .A(DP_OP_102J5_124_3590_n1783), .B(
        DP_OP_102J5_124_3590_n1483), .CI(DP_OP_102J5_124_3590_n2267), .CO(
        DP_OP_102J5_124_3590_n984), .S(DP_OP_102J5_124_3590_n985) );
  FADDX1_HVT DP_OP_102J5_124_3590_U579 ( .A(DP_OP_102J5_124_3590_n1776), .B(
        DP_OP_102J5_124_3590_n2260), .CI(DP_OP_102J5_124_3590_n2230), .CO(
        DP_OP_102J5_124_3590_n982), .S(DP_OP_102J5_124_3590_n983) );
  FADDX1_HVT DP_OP_102J5_124_3590_U578 ( .A(DP_OP_102J5_124_3590_n1740), .B(
        DP_OP_102J5_124_3590_n2223), .CI(DP_OP_102J5_124_3590_n1513), .CO(
        DP_OP_102J5_124_3590_n980), .S(DP_OP_102J5_124_3590_n981) );
  FADDX1_HVT DP_OP_102J5_124_3590_U577 ( .A(DP_OP_102J5_124_3590_n1747), .B(
        DP_OP_102J5_124_3590_n1520), .CI(DP_OP_102J5_124_3590_n1527), .CO(
        DP_OP_102J5_124_3590_n978), .S(DP_OP_102J5_124_3590_n979) );
  FADDX1_HVT DP_OP_102J5_124_3590_U576 ( .A(DP_OP_102J5_124_3590_n1827), .B(
        DP_OP_102J5_124_3590_n1557), .CI(DP_OP_102J5_124_3590_n1564), .CO(
        DP_OP_102J5_124_3590_n976), .S(DP_OP_102J5_124_3590_n977) );
  FADDX1_HVT DP_OP_102J5_124_3590_U575 ( .A(DP_OP_102J5_124_3590_n1864), .B(
        DP_OP_102J5_124_3590_n1571), .CI(DP_OP_102J5_124_3590_n2216), .CO(
        DP_OP_102J5_124_3590_n974), .S(DP_OP_102J5_124_3590_n975) );
  FADDX1_HVT DP_OP_102J5_124_3590_U574 ( .A(DP_OP_102J5_124_3590_n1659), .B(
        DP_OP_102J5_124_3590_n2186), .CI(DP_OP_102J5_124_3590_n1601), .CO(
        DP_OP_102J5_124_3590_n972), .S(DP_OP_102J5_124_3590_n973) );
  FADDX1_HVT DP_OP_102J5_124_3590_U573 ( .A(DP_OP_102J5_124_3590_n2179), .B(
        DP_OP_102J5_124_3590_n1608), .CI(DP_OP_102J5_124_3590_n1615), .CO(
        DP_OP_102J5_124_3590_n970), .S(DP_OP_102J5_124_3590_n971) );
  FADDX1_HVT DP_OP_102J5_124_3590_U572 ( .A(DP_OP_102J5_124_3590_n2172), .B(
        DP_OP_102J5_124_3590_n1645), .CI(DP_OP_102J5_124_3590_n1652), .CO(
        DP_OP_102J5_124_3590_n968), .S(DP_OP_102J5_124_3590_n969) );
  FADDX1_HVT DP_OP_102J5_124_3590_U571 ( .A(DP_OP_102J5_124_3590_n2142), .B(
        DP_OP_102J5_124_3590_n1689), .CI(DP_OP_102J5_124_3590_n1696), .CO(
        DP_OP_102J5_124_3590_n966), .S(DP_OP_102J5_124_3590_n967) );
  FADDX1_HVT DP_OP_102J5_124_3590_U570 ( .A(DP_OP_102J5_124_3590_n2135), .B(
        DP_OP_102J5_124_3590_n1703), .CI(DP_OP_102J5_124_3590_n1733), .CO(
        DP_OP_102J5_124_3590_n964), .S(DP_OP_102J5_124_3590_n965) );
  FADDX1_HVT DP_OP_102J5_124_3590_U569 ( .A(DP_OP_102J5_124_3590_n2128), .B(
        DP_OP_102J5_124_3590_n1871), .CI(DP_OP_102J5_124_3590_n1878), .CO(
        DP_OP_102J5_124_3590_n962), .S(DP_OP_102J5_124_3590_n963) );
  FADDX1_HVT DP_OP_102J5_124_3590_U568 ( .A(DP_OP_102J5_124_3590_n2098), .B(
        DP_OP_102J5_124_3590_n1908), .CI(DP_OP_102J5_124_3590_n1915), .CO(
        DP_OP_102J5_124_3590_n960), .S(DP_OP_102J5_124_3590_n961) );
  FADDX1_HVT DP_OP_102J5_124_3590_U567 ( .A(DP_OP_102J5_124_3590_n2091), .B(
        DP_OP_102J5_124_3590_n1922), .CI(DP_OP_102J5_124_3590_n1952), .CO(
        DP_OP_102J5_124_3590_n958), .S(DP_OP_102J5_124_3590_n959) );
  FADDX1_HVT DP_OP_102J5_124_3590_U566 ( .A(DP_OP_102J5_124_3590_n2084), .B(
        DP_OP_102J5_124_3590_n1959), .CI(DP_OP_102J5_124_3590_n1966), .CO(
        DP_OP_102J5_124_3590_n956), .S(DP_OP_102J5_124_3590_n957) );
  FADDX1_HVT DP_OP_102J5_124_3590_U565 ( .A(DP_OP_102J5_124_3590_n1996), .B(
        DP_OP_102J5_124_3590_n2054), .CI(DP_OP_102J5_124_3590_n2047), .CO(
        DP_OP_102J5_124_3590_n954), .S(DP_OP_102J5_124_3590_n955) );
  FADDX1_HVT DP_OP_102J5_124_3590_U564 ( .A(DP_OP_102J5_124_3590_n2010), .B(
        DP_OP_102J5_124_3590_n2040), .CI(DP_OP_102J5_124_3590_n2003), .CO(
        DP_OP_102J5_124_3590_n952), .S(DP_OP_102J5_124_3590_n953) );
  FADDX1_HVT DP_OP_102J5_124_3590_U563 ( .A(DP_OP_102J5_124_3590_n1138), .B(
        DP_OP_102J5_124_3590_n1132), .CI(DP_OP_102J5_124_3590_n1005), .CO(
        DP_OP_102J5_124_3590_n950), .S(DP_OP_102J5_124_3590_n951) );
  FADDX1_HVT DP_OP_102J5_124_3590_U562 ( .A(DP_OP_102J5_124_3590_n1136), .B(
        DP_OP_102J5_124_3590_n1140), .CI(DP_OP_102J5_124_3590_n1134), .CO(
        DP_OP_102J5_124_3590_n948), .S(DP_OP_102J5_124_3590_n949) );
  FADDX1_HVT DP_OP_102J5_124_3590_U561 ( .A(DP_OP_102J5_124_3590_n1144), .B(
        DP_OP_102J5_124_3590_n1142), .CI(DP_OP_102J5_124_3590_n1114), .CO(
        DP_OP_102J5_124_3590_n946), .S(DP_OP_102J5_124_3590_n947) );
  FADDX1_HVT DP_OP_102J5_124_3590_U560 ( .A(DP_OP_102J5_124_3590_n1112), .B(
        DP_OP_102J5_124_3590_n1096), .CI(DP_OP_102J5_124_3590_n1094), .CO(
        DP_OP_102J5_124_3590_n944), .S(DP_OP_102J5_124_3590_n945) );
  FADDX1_HVT DP_OP_102J5_124_3590_U559 ( .A(DP_OP_102J5_124_3590_n1110), .B(
        DP_OP_102J5_124_3590_n1100), .CI(DP_OP_102J5_124_3590_n1098), .CO(
        DP_OP_102J5_124_3590_n942), .S(DP_OP_102J5_124_3590_n943) );
  FADDX1_HVT DP_OP_102J5_124_3590_U558 ( .A(DP_OP_102J5_124_3590_n1108), .B(
        DP_OP_102J5_124_3590_n1104), .CI(DP_OP_102J5_124_3590_n1102), .CO(
        DP_OP_102J5_124_3590_n940), .S(DP_OP_102J5_124_3590_n941) );
  FADDX1_HVT DP_OP_102J5_124_3590_U557 ( .A(DP_OP_102J5_124_3590_n1106), .B(
        DP_OP_102J5_124_3590_n1118), .CI(DP_OP_102J5_124_3590_n1116), .CO(
        DP_OP_102J5_124_3590_n938), .S(DP_OP_102J5_124_3590_n939) );
  FADDX1_HVT DP_OP_102J5_124_3590_U556 ( .A(DP_OP_102J5_124_3590_n1126), .B(
        DP_OP_102J5_124_3590_n1120), .CI(DP_OP_102J5_124_3590_n1122), .CO(
        DP_OP_102J5_124_3590_n936), .S(DP_OP_102J5_124_3590_n937) );
  FADDX1_HVT DP_OP_102J5_124_3590_U555 ( .A(DP_OP_102J5_124_3590_n1124), .B(
        DP_OP_102J5_124_3590_n1128), .CI(DP_OP_102J5_124_3590_n1130), .CO(
        DP_OP_102J5_124_3590_n934), .S(DP_OP_102J5_124_3590_n935) );
  FADDX1_HVT DP_OP_102J5_124_3590_U554 ( .A(DP_OP_102J5_124_3590_n1092), .B(
        DP_OP_102J5_124_3590_n993), .CI(DP_OP_102J5_124_3590_n995), .CO(
        DP_OP_102J5_124_3590_n932), .S(DP_OP_102J5_124_3590_n933) );
  FADDX1_HVT DP_OP_102J5_124_3590_U553 ( .A(DP_OP_102J5_124_3590_n997), .B(
        DP_OP_102J5_124_3590_n1003), .CI(DP_OP_102J5_124_3590_n1001), .CO(
        DP_OP_102J5_124_3590_n930), .S(DP_OP_102J5_124_3590_n931) );
  FADDX1_HVT DP_OP_102J5_124_3590_U552 ( .A(DP_OP_102J5_124_3590_n999), .B(
        DP_OP_102J5_124_3590_n959), .CI(DP_OP_102J5_124_3590_n957), .CO(
        DP_OP_102J5_124_3590_n928), .S(DP_OP_102J5_124_3590_n929) );
  FADDX1_HVT DP_OP_102J5_124_3590_U551 ( .A(DP_OP_102J5_124_3590_n953), .B(
        DP_OP_102J5_124_3590_n991), .CI(DP_OP_102J5_124_3590_n989), .CO(
        DP_OP_102J5_124_3590_n926), .S(DP_OP_102J5_124_3590_n927) );
  FADDX1_HVT DP_OP_102J5_124_3590_U550 ( .A(DP_OP_102J5_124_3590_n981), .B(
        DP_OP_102J5_124_3590_n979), .CI(DP_OP_102J5_124_3590_n975), .CO(
        DP_OP_102J5_124_3590_n924), .S(DP_OP_102J5_124_3590_n925) );
  FADDX1_HVT DP_OP_102J5_124_3590_U549 ( .A(DP_OP_102J5_124_3590_n983), .B(
        DP_OP_102J5_124_3590_n971), .CI(DP_OP_102J5_124_3590_n969), .CO(
        DP_OP_102J5_124_3590_n922), .S(DP_OP_102J5_124_3590_n923) );
  FADDX1_HVT DP_OP_102J5_124_3590_U548 ( .A(DP_OP_102J5_124_3590_n973), .B(
        DP_OP_102J5_124_3590_n955), .CI(DP_OP_102J5_124_3590_n961), .CO(
        DP_OP_102J5_124_3590_n920), .S(DP_OP_102J5_124_3590_n921) );
  FADDX1_HVT DP_OP_102J5_124_3590_U547 ( .A(DP_OP_102J5_124_3590_n977), .B(
        DP_OP_102J5_124_3590_n963), .CI(DP_OP_102J5_124_3590_n965), .CO(
        DP_OP_102J5_124_3590_n918), .S(DP_OP_102J5_124_3590_n919) );
  FADDX1_HVT DP_OP_102J5_124_3590_U546 ( .A(DP_OP_102J5_124_3590_n967), .B(
        DP_OP_102J5_124_3590_n985), .CI(DP_OP_102J5_124_3590_n987), .CO(
        DP_OP_102J5_124_3590_n916), .S(DP_OP_102J5_124_3590_n917) );
  FADDX1_HVT DP_OP_102J5_124_3590_U545 ( .A(DP_OP_102J5_124_3590_n1088), .B(
        DP_OP_102J5_124_3590_n1090), .CI(DP_OP_102J5_124_3590_n1078), .CO(
        DP_OP_102J5_124_3590_n914), .S(DP_OP_102J5_124_3590_n915) );
  FADDX1_HVT DP_OP_102J5_124_3590_U544 ( .A(DP_OP_102J5_124_3590_n1076), .B(
        DP_OP_102J5_124_3590_n1082), .CI(DP_OP_102J5_124_3590_n1427), .CO(
        DP_OP_102J5_124_3590_n912), .S(DP_OP_102J5_124_3590_n913) );
  FADDX1_HVT DP_OP_102J5_124_3590_U543 ( .A(DP_OP_102J5_124_3590_n1080), .B(
        DP_OP_102J5_124_3590_n1086), .CI(DP_OP_102J5_124_3590_n1074), .CO(
        DP_OP_102J5_124_3590_n910), .S(DP_OP_102J5_124_3590_n911) );
  FADDX1_HVT DP_OP_102J5_124_3590_U542 ( .A(DP_OP_102J5_124_3590_n1084), .B(
        DP_OP_102J5_124_3590_n1072), .CI(DP_OP_102J5_124_3590_n1070), .CO(
        DP_OP_102J5_124_3590_n908), .S(DP_OP_102J5_124_3590_n909) );
  FADDX1_HVT DP_OP_102J5_124_3590_U541 ( .A(DP_OP_102J5_124_3590_n949), .B(
        DP_OP_102J5_124_3590_n951), .CI(DP_OP_102J5_124_3590_n947), .CO(
        DP_OP_102J5_124_3590_n906), .S(DP_OP_102J5_124_3590_n907) );
  FADDX1_HVT DP_OP_102J5_124_3590_U540 ( .A(DP_OP_102J5_124_3590_n1068), .B(
        DP_OP_102J5_124_3590_n935), .CI(DP_OP_102J5_124_3590_n937), .CO(
        DP_OP_102J5_124_3590_n904), .S(DP_OP_102J5_124_3590_n905) );
  FADDX1_HVT DP_OP_102J5_124_3590_U539 ( .A(DP_OP_102J5_124_3590_n941), .B(
        DP_OP_102J5_124_3590_n945), .CI(DP_OP_102J5_124_3590_n943), .CO(
        DP_OP_102J5_124_3590_n902), .S(DP_OP_102J5_124_3590_n903) );
  FADDX1_HVT DP_OP_102J5_124_3590_U538 ( .A(DP_OP_102J5_124_3590_n1066), .B(
        DP_OP_102J5_124_3590_n939), .CI(DP_OP_102J5_124_3590_n1058), .CO(
        DP_OP_102J5_124_3590_n900), .S(DP_OP_102J5_124_3590_n901) );
  FADDX1_HVT DP_OP_102J5_124_3590_U537 ( .A(DP_OP_102J5_124_3590_n1064), .B(
        DP_OP_102J5_124_3590_n1060), .CI(DP_OP_102J5_124_3590_n1062), .CO(
        DP_OP_102J5_124_3590_n898), .S(DP_OP_102J5_124_3590_n899) );
  FADDX1_HVT DP_OP_102J5_124_3590_U536 ( .A(DP_OP_102J5_124_3590_n933), .B(
        DP_OP_102J5_124_3590_n931), .CI(DP_OP_102J5_124_3590_n929), .CO(
        DP_OP_102J5_124_3590_n896), .S(DP_OP_102J5_124_3590_n897) );
  FADDX1_HVT DP_OP_102J5_124_3590_U535 ( .A(DP_OP_102J5_124_3590_n1056), .B(
        DP_OP_102J5_124_3590_n923), .CI(DP_OP_102J5_124_3590_n925), .CO(
        DP_OP_102J5_124_3590_n894), .S(DP_OP_102J5_124_3590_n895) );
  FADDX1_HVT DP_OP_102J5_124_3590_U534 ( .A(DP_OP_102J5_124_3590_n921), .B(
        DP_OP_102J5_124_3590_n927), .CI(DP_OP_102J5_124_3590_n919), .CO(
        DP_OP_102J5_124_3590_n892), .S(DP_OP_102J5_124_3590_n893) );
  FADDX1_HVT DP_OP_102J5_124_3590_U533 ( .A(DP_OP_102J5_124_3590_n917), .B(
        DP_OP_102J5_124_3590_n1054), .CI(DP_OP_102J5_124_3590_n1052), .CO(
        DP_OP_102J5_124_3590_n890), .S(DP_OP_102J5_124_3590_n891) );
  FADDX1_HVT DP_OP_102J5_124_3590_U532 ( .A(DP_OP_102J5_124_3590_n1050), .B(
        DP_OP_102J5_124_3590_n1048), .CI(DP_OP_102J5_124_3590_n915), .CO(
        DP_OP_102J5_124_3590_n888), .S(DP_OP_102J5_124_3590_n889) );
  FADDX1_HVT DP_OP_102J5_124_3590_U531 ( .A(DP_OP_102J5_124_3590_n1046), .B(
        DP_OP_102J5_124_3590_n913), .CI(DP_OP_102J5_124_3590_n911), .CO(
        DP_OP_102J5_124_3590_n886), .S(DP_OP_102J5_124_3590_n887) );
  FADDX1_HVT DP_OP_102J5_124_3590_U530 ( .A(DP_OP_102J5_124_3590_n1044), .B(
        DP_OP_102J5_124_3590_n1040), .CI(DP_OP_102J5_124_3590_n1042), .CO(
        DP_OP_102J5_124_3590_n884), .S(DP_OP_102J5_124_3590_n885) );
  FADDX1_HVT DP_OP_102J5_124_3590_U529 ( .A(DP_OP_102J5_124_3590_n909), .B(
        DP_OP_102J5_124_3590_n1038), .CI(DP_OP_102J5_124_3590_n907), .CO(
        DP_OP_102J5_124_3590_n882), .S(DP_OP_102J5_124_3590_n883) );
  FADDX1_HVT DP_OP_102J5_124_3590_U528 ( .A(DP_OP_102J5_124_3590_n1036), .B(
        DP_OP_102J5_124_3590_n903), .CI(DP_OP_102J5_124_3590_n905), .CO(
        DP_OP_102J5_124_3590_n880), .S(DP_OP_102J5_124_3590_n881) );
  FADDX1_HVT DP_OP_102J5_124_3590_U527 ( .A(DP_OP_102J5_124_3590_n1034), .B(
        DP_OP_102J5_124_3590_n899), .CI(DP_OP_102J5_124_3590_n901), .CO(
        DP_OP_102J5_124_3590_n878), .S(DP_OP_102J5_124_3590_n879) );
  FADDX1_HVT DP_OP_102J5_124_3590_U526 ( .A(DP_OP_102J5_124_3590_n1032), .B(
        DP_OP_102J5_124_3590_n897), .CI(DP_OP_102J5_124_3590_n895), .CO(
        DP_OP_102J5_124_3590_n876), .S(DP_OP_102J5_124_3590_n877) );
  FADDX1_HVT DP_OP_102J5_124_3590_U525 ( .A(DP_OP_102J5_124_3590_n893), .B(
        DP_OP_102J5_124_3590_n891), .CI(DP_OP_102J5_124_3590_n1030), .CO(
        DP_OP_102J5_124_3590_n874), .S(DP_OP_102J5_124_3590_n875) );
  FADDX1_HVT DP_OP_102J5_124_3590_U524 ( .A(DP_OP_102J5_124_3590_n1028), .B(
        DP_OP_102J5_124_3590_n1026), .CI(DP_OP_102J5_124_3590_n889), .CO(
        DP_OP_102J5_124_3590_n872), .S(DP_OP_102J5_124_3590_n873) );
  FADDX1_HVT DP_OP_102J5_124_3590_U523 ( .A(DP_OP_102J5_124_3590_n1024), .B(
        DP_OP_102J5_124_3590_n885), .CI(DP_OP_102J5_124_3590_n887), .CO(
        DP_OP_102J5_124_3590_n870), .S(DP_OP_102J5_124_3590_n871) );
  FADDX1_HVT DP_OP_102J5_124_3590_U522 ( .A(DP_OP_102J5_124_3590_n1022), .B(
        DP_OP_102J5_124_3590_n883), .CI(DP_OP_102J5_124_3590_n1020), .CO(
        DP_OP_102J5_124_3590_n868), .S(DP_OP_102J5_124_3590_n869) );
  FADDX1_HVT DP_OP_102J5_124_3590_U521 ( .A(DP_OP_102J5_124_3590_n881), .B(
        DP_OP_102J5_124_3590_n879), .CI(DP_OP_102J5_124_3590_n1018), .CO(
        DP_OP_102J5_124_3590_n866), .S(DP_OP_102J5_124_3590_n867) );
  FADDX1_HVT DP_OP_102J5_124_3590_U520 ( .A(DP_OP_102J5_124_3590_n877), .B(
        DP_OP_102J5_124_3590_n875), .CI(DP_OP_102J5_124_3590_n1016), .CO(
        DP_OP_102J5_124_3590_n864), .S(DP_OP_102J5_124_3590_n865) );
  FADDX1_HVT DP_OP_102J5_124_3590_U519 ( .A(DP_OP_102J5_124_3590_n1014), .B(
        DP_OP_102J5_124_3590_n873), .CI(DP_OP_102J5_124_3590_n871), .CO(
        DP_OP_102J5_124_3590_n862), .S(DP_OP_102J5_124_3590_n863) );
  FADDX1_HVT DP_OP_102J5_124_3590_U518 ( .A(DP_OP_102J5_124_3590_n1012), .B(
        DP_OP_102J5_124_3590_n869), .CI(DP_OP_102J5_124_3590_n867), .CO(
        DP_OP_102J5_124_3590_n860), .S(DP_OP_102J5_124_3590_n861) );
  FADDX1_HVT DP_OP_102J5_124_3590_U517 ( .A(DP_OP_102J5_124_3590_n1010), .B(
        DP_OP_102J5_124_3590_n865), .CI(DP_OP_102J5_124_3590_n1008), .CO(
        DP_OP_102J5_124_3590_n858), .S(DP_OP_102J5_124_3590_n859) );
  FADDX1_HVT DP_OP_102J5_124_3590_U516 ( .A(DP_OP_102J5_124_3590_n863), .B(
        DP_OP_102J5_124_3590_n861), .CI(DP_OP_102J5_124_3590_n1006), .CO(
        DP_OP_102J5_124_3590_n856), .S(DP_OP_102J5_124_3590_n857) );
  FADDX1_HVT DP_OP_102J5_124_3590_U515 ( .A(DP_OP_102J5_124_3590_n2032), .B(
        DP_OP_102J5_124_3590_n1856), .CI(DP_OP_102J5_124_3590_n1461), .CO(
        DP_OP_102J5_124_3590_n854), .S(DP_OP_102J5_124_3590_n855) );
  FADDX1_HVT DP_OP_102J5_124_3590_U514 ( .A(DP_OP_102J5_124_3590_n2120), .B(
        DP_OP_102J5_124_3590_n1988), .CI(DP_OP_102J5_124_3590_n1944), .CO(
        DP_OP_102J5_124_3590_n852), .S(DP_OP_102J5_124_3590_n853) );
  FADDX1_HVT DP_OP_102J5_124_3590_U513 ( .A(DP_OP_102J5_124_3590_n1900), .B(
        DP_OP_102J5_124_3590_n1681), .CI(DP_OP_102J5_124_3590_n1768), .CO(
        DP_OP_102J5_124_3590_n850), .S(DP_OP_102J5_124_3590_n851) );
  FADDX1_HVT DP_OP_102J5_124_3590_U512 ( .A(DP_OP_102J5_124_3590_n2164), .B(
        DP_OP_102J5_124_3590_n1549), .CI(DP_OP_102J5_124_3590_n2076), .CO(
        DP_OP_102J5_124_3590_n848), .S(DP_OP_102J5_124_3590_n849) );
  FADDX1_HVT DP_OP_102J5_124_3590_U511 ( .A(DP_OP_102J5_124_3590_n1505), .B(
        DP_OP_102J5_124_3590_n2252), .CI(DP_OP_102J5_124_3590_n1637), .CO(
        DP_OP_102J5_124_3590_n846), .S(DP_OP_102J5_124_3590_n847) );
  FADDX1_HVT DP_OP_102J5_124_3590_U510 ( .A(DP_OP_102J5_124_3590_n2296), .B(
        DP_OP_102J5_124_3590_n1725), .CI(DP_OP_102J5_124_3590_n2208), .CO(
        DP_OP_102J5_124_3590_n844), .S(DP_OP_102J5_124_3590_n845) );
  FADDX1_HVT DP_OP_102J5_124_3590_U509 ( .A(DP_OP_102J5_124_3590_n1593), .B(
        DP_OP_102J5_124_3590_n1812), .CI(DP_OP_102J5_124_3590_n1819), .CO(
        DP_OP_102J5_124_3590_n842), .S(DP_OP_102J5_124_3590_n843) );
  FADDX1_HVT DP_OP_102J5_124_3590_U508 ( .A(DP_OP_102J5_124_3590_n1826), .B(
        DP_OP_102J5_124_3590_n2316), .CI(DP_OP_102J5_124_3590_n2310), .CO(
        DP_OP_102J5_124_3590_n840), .S(DP_OP_102J5_124_3590_n841) );
  FADDX1_HVT DP_OP_102J5_124_3590_U507 ( .A(DP_OP_102J5_124_3590_n1782), .B(
        DP_OP_102J5_124_3590_n2303), .CI(DP_OP_102J5_124_3590_n2273), .CO(
        DP_OP_102J5_124_3590_n838), .S(DP_OP_102J5_124_3590_n839) );
  FADDX1_HVT DP_OP_102J5_124_3590_U506 ( .A(DP_OP_102J5_124_3590_n1775), .B(
        DP_OP_102J5_124_3590_n2266), .CI(DP_OP_102J5_124_3590_n1468), .CO(
        DP_OP_102J5_124_3590_n836), .S(DP_OP_102J5_124_3590_n837) );
  FADDX1_HVT DP_OP_102J5_124_3590_U505 ( .A(DP_OP_102J5_124_3590_n1746), .B(
        DP_OP_102J5_124_3590_n2259), .CI(DP_OP_102J5_124_3590_n2229), .CO(
        DP_OP_102J5_124_3590_n834), .S(DP_OP_102J5_124_3590_n835) );
  FADDX1_HVT DP_OP_102J5_124_3590_U504 ( .A(DP_OP_102J5_124_3590_n1739), .B(
        DP_OP_102J5_124_3590_n2222), .CI(DP_OP_102J5_124_3590_n2215), .CO(
        DP_OP_102J5_124_3590_n832), .S(DP_OP_102J5_124_3590_n833) );
  FADDX1_HVT DP_OP_102J5_124_3590_U503 ( .A(DP_OP_102J5_124_3590_n1702), .B(
        DP_OP_102J5_124_3590_n2185), .CI(DP_OP_102J5_124_3590_n2178), .CO(
        DP_OP_102J5_124_3590_n830), .S(DP_OP_102J5_124_3590_n831) );
  FADDX1_HVT DP_OP_102J5_124_3590_U502 ( .A(DP_OP_102J5_124_3590_n1695), .B(
        DP_OP_102J5_124_3590_n2171), .CI(DP_OP_102J5_124_3590_n2141), .CO(
        DP_OP_102J5_124_3590_n828), .S(DP_OP_102J5_124_3590_n829) );
  FADDX1_HVT DP_OP_102J5_124_3590_U501 ( .A(DP_OP_102J5_124_3590_n2134), .B(
        DP_OP_102J5_124_3590_n1475), .CI(DP_OP_102J5_124_3590_n1482), .CO(
        DP_OP_102J5_124_3590_n826), .S(DP_OP_102J5_124_3590_n827) );
  FADDX1_HVT DP_OP_102J5_124_3590_U500 ( .A(DP_OP_102J5_124_3590_n1907), .B(
        DP_OP_102J5_124_3590_n2127), .CI(DP_OP_102J5_124_3590_n2097), .CO(
        DP_OP_102J5_124_3590_n824), .S(DP_OP_102J5_124_3590_n825) );
  FADDX1_HVT DP_OP_102J5_124_3590_U499 ( .A(DP_OP_102J5_124_3590_n2090), .B(
        DP_OP_102J5_124_3590_n1512), .CI(DP_OP_102J5_124_3590_n1519), .CO(
        DP_OP_102J5_124_3590_n822), .S(DP_OP_102J5_124_3590_n823) );
  FADDX1_HVT DP_OP_102J5_124_3590_U498 ( .A(DP_OP_102J5_124_3590_n2083), .B(
        DP_OP_102J5_124_3590_n1526), .CI(DP_OP_102J5_124_3590_n1556), .CO(
        DP_OP_102J5_124_3590_n820), .S(DP_OP_102J5_124_3590_n821) );
  FADDX1_HVT DP_OP_102J5_124_3590_U497 ( .A(DP_OP_102J5_124_3590_n2053), .B(
        DP_OP_102J5_124_3590_n1563), .CI(DP_OP_102J5_124_3590_n1570), .CO(
        DP_OP_102J5_124_3590_n818), .S(DP_OP_102J5_124_3590_n819) );
  FADDX1_HVT DP_OP_102J5_124_3590_U496 ( .A(DP_OP_102J5_124_3590_n2046), .B(
        DP_OP_102J5_124_3590_n1600), .CI(DP_OP_102J5_124_3590_n1607), .CO(
        DP_OP_102J5_124_3590_n816), .S(DP_OP_102J5_124_3590_n817) );
  FADDX1_HVT DP_OP_102J5_124_3590_U495 ( .A(DP_OP_102J5_124_3590_n2039), .B(
        DP_OP_102J5_124_3590_n1614), .CI(DP_OP_102J5_124_3590_n1644), .CO(
        DP_OP_102J5_124_3590_n814), .S(DP_OP_102J5_124_3590_n815) );
  FADDX1_HVT DP_OP_102J5_124_3590_U494 ( .A(DP_OP_102J5_124_3590_n2009), .B(
        DP_OP_102J5_124_3590_n1651), .CI(DP_OP_102J5_124_3590_n1658), .CO(
        DP_OP_102J5_124_3590_n812), .S(DP_OP_102J5_124_3590_n813) );
  FADDX1_HVT DP_OP_102J5_124_3590_U493 ( .A(DP_OP_102J5_124_3590_n2002), .B(
        DP_OP_102J5_124_3590_n1688), .CI(DP_OP_102J5_124_3590_n1732), .CO(
        DP_OP_102J5_124_3590_n810), .S(DP_OP_102J5_124_3590_n811) );
  FADDX1_HVT DP_OP_102J5_124_3590_U492 ( .A(DP_OP_102J5_124_3590_n1995), .B(
        DP_OP_102J5_124_3590_n1789), .CI(DP_OP_102J5_124_3590_n1833), .CO(
        DP_OP_102J5_124_3590_n808), .S(DP_OP_102J5_124_3590_n809) );
  FADDX1_HVT DP_OP_102J5_124_3590_U491 ( .A(DP_OP_102J5_124_3590_n1965), .B(
        DP_OP_102J5_124_3590_n1863), .CI(DP_OP_102J5_124_3590_n1870), .CO(
        DP_OP_102J5_124_3590_n806), .S(DP_OP_102J5_124_3590_n807) );
  FADDX1_HVT DP_OP_102J5_124_3590_U490 ( .A(DP_OP_102J5_124_3590_n1958), .B(
        DP_OP_102J5_124_3590_n1877), .CI(DP_OP_102J5_124_3590_n1914), .CO(
        DP_OP_102J5_124_3590_n804), .S(DP_OP_102J5_124_3590_n805) );
  FADDX1_HVT DP_OP_102J5_124_3590_U489 ( .A(DP_OP_102J5_124_3590_n1951), .B(
        DP_OP_102J5_124_3590_n1921), .CI(DP_OP_102J5_124_3590_n1004), .CO(
        DP_OP_102J5_124_3590_n802), .S(DP_OP_102J5_124_3590_n803) );
  FADDX1_HVT DP_OP_102J5_124_3590_U488 ( .A(DP_OP_102J5_124_3590_n996), .B(
        DP_OP_102J5_124_3590_n992), .CI(DP_OP_102J5_124_3590_n998), .CO(
        DP_OP_102J5_124_3590_n800), .S(DP_OP_102J5_124_3590_n801) );
  FADDX1_HVT DP_OP_102J5_124_3590_U487 ( .A(DP_OP_102J5_124_3590_n1002), .B(
        DP_OP_102J5_124_3590_n994), .CI(DP_OP_102J5_124_3590_n1000), .CO(
        DP_OP_102J5_124_3590_n798), .S(DP_OP_102J5_124_3590_n799) );
  FADDX1_HVT DP_OP_102J5_124_3590_U486 ( .A(DP_OP_102J5_124_3590_n972), .B(
        DP_OP_102J5_124_3590_n952), .CI(DP_OP_102J5_124_3590_n956), .CO(
        DP_OP_102J5_124_3590_n796), .S(DP_OP_102J5_124_3590_n797) );
  FADDX1_HVT DP_OP_102J5_124_3590_U485 ( .A(DP_OP_102J5_124_3590_n974), .B(
        DP_OP_102J5_124_3590_n954), .CI(DP_OP_102J5_124_3590_n958), .CO(
        DP_OP_102J5_124_3590_n794), .S(DP_OP_102J5_124_3590_n795) );
  FADDX1_HVT DP_OP_102J5_124_3590_U484 ( .A(DP_OP_102J5_124_3590_n970), .B(
        DP_OP_102J5_124_3590_n960), .CI(DP_OP_102J5_124_3590_n962), .CO(
        DP_OP_102J5_124_3590_n792), .S(DP_OP_102J5_124_3590_n793) );
  FADDX1_HVT DP_OP_102J5_124_3590_U483 ( .A(DP_OP_102J5_124_3590_n968), .B(
        DP_OP_102J5_124_3590_n964), .CI(DP_OP_102J5_124_3590_n976), .CO(
        DP_OP_102J5_124_3590_n790), .S(DP_OP_102J5_124_3590_n791) );
  FADDX1_HVT DP_OP_102J5_124_3590_U482 ( .A(DP_OP_102J5_124_3590_n984), .B(
        DP_OP_102J5_124_3590_n966), .CI(DP_OP_102J5_124_3590_n980), .CO(
        DP_OP_102J5_124_3590_n788), .S(DP_OP_102J5_124_3590_n789) );
  FADDX1_HVT DP_OP_102J5_124_3590_U481 ( .A(DP_OP_102J5_124_3590_n986), .B(
        DP_OP_102J5_124_3590_n978), .CI(DP_OP_102J5_124_3590_n988), .CO(
        DP_OP_102J5_124_3590_n786), .S(DP_OP_102J5_124_3590_n787) );
  FADDX1_HVT DP_OP_102J5_124_3590_U480 ( .A(DP_OP_102J5_124_3590_n990), .B(
        DP_OP_102J5_124_3590_n982), .CI(DP_OP_102J5_124_3590_n847), .CO(
        DP_OP_102J5_124_3590_n784), .S(DP_OP_102J5_124_3590_n785) );
  FADDX1_HVT DP_OP_102J5_124_3590_U479 ( .A(DP_OP_102J5_124_3590_n849), .B(
        DP_OP_102J5_124_3590_n855), .CI(DP_OP_102J5_124_3590_n843), .CO(
        DP_OP_102J5_124_3590_n782), .S(DP_OP_102J5_124_3590_n783) );
  FADDX1_HVT DP_OP_102J5_124_3590_U478 ( .A(DP_OP_102J5_124_3590_n845), .B(
        DP_OP_102J5_124_3590_n853), .CI(DP_OP_102J5_124_3590_n851), .CO(
        DP_OP_102J5_124_3590_n780), .S(DP_OP_102J5_124_3590_n781) );
  FADDX1_HVT DP_OP_102J5_124_3590_U477 ( .A(DP_OP_102J5_124_3590_n809), .B(
        DP_OP_102J5_124_3590_n835), .CI(DP_OP_102J5_124_3590_n841), .CO(
        DP_OP_102J5_124_3590_n778), .S(DP_OP_102J5_124_3590_n779) );
  FADDX1_HVT DP_OP_102J5_124_3590_U476 ( .A(DP_OP_102J5_124_3590_n831), .B(
        DP_OP_102J5_124_3590_n825), .CI(DP_OP_102J5_124_3590_n823), .CO(
        DP_OP_102J5_124_3590_n776), .S(DP_OP_102J5_124_3590_n777) );
  FADDX1_HVT DP_OP_102J5_124_3590_U475 ( .A(DP_OP_102J5_124_3590_n833), .B(
        DP_OP_102J5_124_3590_n821), .CI(DP_OP_102J5_124_3590_n819), .CO(
        DP_OP_102J5_124_3590_n774), .S(DP_OP_102J5_124_3590_n775) );
  FADDX1_HVT DP_OP_102J5_124_3590_U474 ( .A(DP_OP_102J5_124_3590_n827), .B(
        DP_OP_102J5_124_3590_n817), .CI(DP_OP_102J5_124_3590_n805), .CO(
        DP_OP_102J5_124_3590_n772), .S(DP_OP_102J5_124_3590_n773) );
  FADDX1_HVT DP_OP_102J5_124_3590_U473 ( .A(DP_OP_102J5_124_3590_n829), .B(
        DP_OP_102J5_124_3590_n811), .CI(DP_OP_102J5_124_3590_n807), .CO(
        DP_OP_102J5_124_3590_n770), .S(DP_OP_102J5_124_3590_n771) );
  FADDX1_HVT DP_OP_102J5_124_3590_U472 ( .A(DP_OP_102J5_124_3590_n815), .B(
        DP_OP_102J5_124_3590_n839), .CI(DP_OP_102J5_124_3590_n837), .CO(
        DP_OP_102J5_124_3590_n768), .S(DP_OP_102J5_124_3590_n769) );
  FADDX1_HVT DP_OP_102J5_124_3590_U471 ( .A(DP_OP_102J5_124_3590_n813), .B(
        DP_OP_102J5_124_3590_n803), .CI(DP_OP_102J5_124_3590_n948), .CO(
        DP_OP_102J5_124_3590_n766), .S(DP_OP_102J5_124_3590_n767) );
  FADDX1_HVT DP_OP_102J5_124_3590_U470 ( .A(DP_OP_102J5_124_3590_n946), .B(
        DP_OP_102J5_124_3590_n950), .CI(DP_OP_102J5_124_3590_n936), .CO(
        DP_OP_102J5_124_3590_n764), .S(DP_OP_102J5_124_3590_n765) );
  FADDX1_HVT DP_OP_102J5_124_3590_U469 ( .A(DP_OP_102J5_124_3590_n934), .B(
        DP_OP_102J5_124_3590_n940), .CI(DP_OP_102J5_124_3590_n1426), .CO(
        DP_OP_102J5_124_3590_n762), .S(DP_OP_102J5_124_3590_n763) );
  FADDX1_HVT DP_OP_102J5_124_3590_U468 ( .A(DP_OP_102J5_124_3590_n938), .B(
        DP_OP_102J5_124_3590_n942), .CI(DP_OP_102J5_124_3590_n944), .CO(
        DP_OP_102J5_124_3590_n760), .S(DP_OP_102J5_124_3590_n761) );
  FADDX1_HVT DP_OP_102J5_124_3590_U467 ( .A(DP_OP_102J5_124_3590_n932), .B(
        DP_OP_102J5_124_3590_n930), .CI(DP_OP_102J5_124_3590_n928), .CO(
        DP_OP_102J5_124_3590_n758), .S(DP_OP_102J5_124_3590_n759) );
  FADDX1_HVT DP_OP_102J5_124_3590_U466 ( .A(DP_OP_102J5_124_3590_n799), .B(
        DP_OP_102J5_124_3590_n801), .CI(DP_OP_102J5_124_3590_n795), .CO(
        DP_OP_102J5_124_3590_n756), .S(DP_OP_102J5_124_3590_n757) );
  FADDX1_HVT DP_OP_102J5_124_3590_U465 ( .A(DP_OP_102J5_124_3590_n791), .B(
        DP_OP_102J5_124_3590_n797), .CI(DP_OP_102J5_124_3590_n785), .CO(
        DP_OP_102J5_124_3590_n754), .S(DP_OP_102J5_124_3590_n755) );
  FADDX1_HVT DP_OP_102J5_124_3590_U464 ( .A(DP_OP_102J5_124_3590_n926), .B(
        DP_OP_102J5_124_3590_n793), .CI(DP_OP_102J5_124_3590_n789), .CO(
        DP_OP_102J5_124_3590_n752), .S(DP_OP_102J5_124_3590_n753) );
  FADDX1_HVT DP_OP_102J5_124_3590_U463 ( .A(DP_OP_102J5_124_3590_n924), .B(
        DP_OP_102J5_124_3590_n787), .CI(DP_OP_102J5_124_3590_n916), .CO(
        DP_OP_102J5_124_3590_n750), .S(DP_OP_102J5_124_3590_n751) );
  FADDX1_HVT DP_OP_102J5_124_3590_U462 ( .A(DP_OP_102J5_124_3590_n922), .B(
        DP_OP_102J5_124_3590_n918), .CI(DP_OP_102J5_124_3590_n920), .CO(
        DP_OP_102J5_124_3590_n748), .S(DP_OP_102J5_124_3590_n749) );
  FADDX1_HVT DP_OP_102J5_124_3590_U461 ( .A(DP_OP_102J5_124_3590_n781), .B(
        DP_OP_102J5_124_3590_n783), .CI(DP_OP_102J5_124_3590_n777), .CO(
        DP_OP_102J5_124_3590_n746), .S(DP_OP_102J5_124_3590_n747) );
  FADDX1_HVT DP_OP_102J5_124_3590_U460 ( .A(DP_OP_102J5_124_3590_n775), .B(
        DP_OP_102J5_124_3590_n771), .CI(DP_OP_102J5_124_3590_n914), .CO(
        DP_OP_102J5_124_3590_n744), .S(DP_OP_102J5_124_3590_n745) );
  FADDX1_HVT DP_OP_102J5_124_3590_U459 ( .A(DP_OP_102J5_124_3590_n773), .B(
        DP_OP_102J5_124_3590_n779), .CI(DP_OP_102J5_124_3590_n769), .CO(
        DP_OP_102J5_124_3590_n742), .S(DP_OP_102J5_124_3590_n743) );
  FADDX1_HVT DP_OP_102J5_124_3590_U458 ( .A(DP_OP_102J5_124_3590_n912), .B(
        DP_OP_102J5_124_3590_n910), .CI(DP_OP_102J5_124_3590_n767), .CO(
        DP_OP_102J5_124_3590_n740), .S(DP_OP_102J5_124_3590_n741) );
  FADDX1_HVT DP_OP_102J5_124_3590_U457 ( .A(DP_OP_102J5_124_3590_n908), .B(
        DP_OP_102J5_124_3590_n906), .CI(DP_OP_102J5_124_3590_n765), .CO(
        DP_OP_102J5_124_3590_n738), .S(DP_OP_102J5_124_3590_n739) );
  FADDX1_HVT DP_OP_102J5_124_3590_U456 ( .A(DP_OP_102J5_124_3590_n904), .B(
        DP_OP_102J5_124_3590_n763), .CI(DP_OP_102J5_124_3590_n761), .CO(
        DP_OP_102J5_124_3590_n736), .S(DP_OP_102J5_124_3590_n737) );
  FADDX1_HVT DP_OP_102J5_124_3590_U455 ( .A(DP_OP_102J5_124_3590_n902), .B(
        DP_OP_102J5_124_3590_n898), .CI(DP_OP_102J5_124_3590_n900), .CO(
        DP_OP_102J5_124_3590_n734), .S(DP_OP_102J5_124_3590_n735) );
  FADDX1_HVT DP_OP_102J5_124_3590_U454 ( .A(DP_OP_102J5_124_3590_n896), .B(
        DP_OP_102J5_124_3590_n757), .CI(DP_OP_102J5_124_3590_n894), .CO(
        DP_OP_102J5_124_3590_n732), .S(DP_OP_102J5_124_3590_n733) );
  FADDX1_HVT DP_OP_102J5_124_3590_U453 ( .A(DP_OP_102J5_124_3590_n759), .B(
        DP_OP_102J5_124_3590_n892), .CI(DP_OP_102J5_124_3590_n753), .CO(
        DP_OP_102J5_124_3590_n730), .S(DP_OP_102J5_124_3590_n731) );
  FADDX1_HVT DP_OP_102J5_124_3590_U452 ( .A(DP_OP_102J5_124_3590_n749), .B(
        DP_OP_102J5_124_3590_n755), .CI(DP_OP_102J5_124_3590_n890), .CO(
        DP_OP_102J5_124_3590_n728), .S(DP_OP_102J5_124_3590_n729) );
  FADDX1_HVT DP_OP_102J5_124_3590_U451 ( .A(DP_OP_102J5_124_3590_n751), .B(
        DP_OP_102J5_124_3590_n747), .CI(DP_OP_102J5_124_3590_n888), .CO(
        DP_OP_102J5_124_3590_n726), .S(DP_OP_102J5_124_3590_n727) );
  FADDX1_HVT DP_OP_102J5_124_3590_U450 ( .A(DP_OP_102J5_124_3590_n743), .B(
        DP_OP_102J5_124_3590_n745), .CI(DP_OP_102J5_124_3590_n886), .CO(
        DP_OP_102J5_124_3590_n724), .S(DP_OP_102J5_124_3590_n725) );
  FADDX1_HVT DP_OP_102J5_124_3590_U449 ( .A(DP_OP_102J5_124_3590_n884), .B(
        DP_OP_102J5_124_3590_n741), .CI(DP_OP_102J5_124_3590_n882), .CO(
        DP_OP_102J5_124_3590_n722), .S(DP_OP_102J5_124_3590_n723) );
  FADDX1_HVT DP_OP_102J5_124_3590_U448 ( .A(DP_OP_102J5_124_3590_n739), .B(
        DP_OP_102J5_124_3590_n880), .CI(DP_OP_102J5_124_3590_n878), .CO(
        DP_OP_102J5_124_3590_n720), .S(DP_OP_102J5_124_3590_n721) );
  FADDX1_HVT DP_OP_102J5_124_3590_U447 ( .A(DP_OP_102J5_124_3590_n737), .B(
        DP_OP_102J5_124_3590_n735), .CI(DP_OP_102J5_124_3590_n876), .CO(
        DP_OP_102J5_124_3590_n718), .S(DP_OP_102J5_124_3590_n719) );
  FADDX1_HVT DP_OP_102J5_124_3590_U446 ( .A(DP_OP_102J5_124_3590_n733), .B(
        DP_OP_102J5_124_3590_n731), .CI(DP_OP_102J5_124_3590_n729), .CO(
        DP_OP_102J5_124_3590_n716), .S(DP_OP_102J5_124_3590_n717) );
  FADDX1_HVT DP_OP_102J5_124_3590_U445 ( .A(DP_OP_102J5_124_3590_n874), .B(
        DP_OP_102J5_124_3590_n727), .CI(DP_OP_102J5_124_3590_n872), .CO(
        DP_OP_102J5_124_3590_n714), .S(DP_OP_102J5_124_3590_n715) );
  FADDX1_HVT DP_OP_102J5_124_3590_U444 ( .A(DP_OP_102J5_124_3590_n725), .B(
        DP_OP_102J5_124_3590_n870), .CI(DP_OP_102J5_124_3590_n723), .CO(
        DP_OP_102J5_124_3590_n712), .S(DP_OP_102J5_124_3590_n713) );
  FADDX1_HVT DP_OP_102J5_124_3590_U443 ( .A(DP_OP_102J5_124_3590_n868), .B(
        DP_OP_102J5_124_3590_n721), .CI(DP_OP_102J5_124_3590_n866), .CO(
        DP_OP_102J5_124_3590_n710), .S(DP_OP_102J5_124_3590_n711) );
  FADDX1_HVT DP_OP_102J5_124_3590_U442 ( .A(DP_OP_102J5_124_3590_n719), .B(
        DP_OP_102J5_124_3590_n717), .CI(DP_OP_102J5_124_3590_n864), .CO(
        DP_OP_102J5_124_3590_n708), .S(DP_OP_102J5_124_3590_n709) );
  FADDX1_HVT DP_OP_102J5_124_3590_U441 ( .A(DP_OP_102J5_124_3590_n715), .B(
        DP_OP_102J5_124_3590_n862), .CI(DP_OP_102J5_124_3590_n713), .CO(
        DP_OP_102J5_124_3590_n706), .S(DP_OP_102J5_124_3590_n707) );
  FADDX1_HVT DP_OP_102J5_124_3590_U440 ( .A(DP_OP_102J5_124_3590_n860), .B(
        DP_OP_102J5_124_3590_n711), .CI(DP_OP_102J5_124_3590_n709), .CO(
        DP_OP_102J5_124_3590_n704), .S(DP_OP_102J5_124_3590_n705) );
  FADDX1_HVT DP_OP_102J5_124_3590_U439 ( .A(DP_OP_102J5_124_3590_n858), .B(
        DP_OP_102J5_124_3590_n707), .CI(DP_OP_102J5_124_3590_n856), .CO(
        DP_OP_102J5_124_3590_n702), .S(DP_OP_102J5_124_3590_n703) );
  FADDX1_HVT DP_OP_102J5_124_3590_U437 ( .A(DP_OP_102J5_124_3590_n1832), .B(
        DP_OP_102J5_124_3590_n1481), .CI(DP_OP_102J5_124_3590_n1460), .CO(
        DP_OP_102J5_124_3590_n698), .S(DP_OP_102J5_124_3590_n699) );
  FADDX1_HVT DP_OP_102J5_124_3590_U436 ( .A(DP_OP_102J5_124_3590_n2228), .B(
        DP_OP_102J5_124_3590_n1680), .CI(DP_OP_102J5_124_3590_n1811), .CO(
        DP_OP_102J5_124_3590_n696), .S(DP_OP_102J5_124_3590_n697) );
  FADDX1_HVT DP_OP_102J5_124_3590_U435 ( .A(DP_OP_102J5_124_3590_n1504), .B(
        DP_OP_102J5_124_3590_n1569), .CI(DP_OP_102J5_124_3590_n1701), .CO(
        DP_OP_102J5_124_3590_n694), .S(DP_OP_102J5_124_3590_n695) );
  FADDX1_HVT DP_OP_102J5_124_3590_U434 ( .A(DP_OP_102J5_124_3590_n1943), .B(
        DP_OP_102J5_124_3590_n1899), .CI(DP_OP_102J5_124_3590_n1767), .CO(
        DP_OP_102J5_124_3590_n692), .S(DP_OP_102J5_124_3590_n693) );
  FADDX1_HVT DP_OP_102J5_124_3590_U433 ( .A(DP_OP_102J5_124_3590_n2119), .B(
        DP_OP_102J5_124_3590_n1964), .CI(DP_OP_102J5_124_3590_n2008), .CO(
        DP_OP_102J5_124_3590_n690), .S(DP_OP_102J5_124_3590_n691) );
  FADDX1_HVT DP_OP_102J5_124_3590_U432 ( .A(DP_OP_102J5_124_3590_n1855), .B(
        DP_OP_102J5_124_3590_n1788), .CI(DP_OP_102J5_124_3590_n1548), .CO(
        DP_OP_102J5_124_3590_n688), .S(DP_OP_102J5_124_3590_n689) );
  FADDX1_HVT DP_OP_102J5_124_3590_U431 ( .A(DP_OP_102J5_124_3590_n1613), .B(
        DP_OP_102J5_124_3590_n2031), .CI(DP_OP_102J5_124_3590_n1876), .CO(
        DP_OP_102J5_124_3590_n686), .S(DP_OP_102J5_124_3590_n687) );
  FADDX1_HVT DP_OP_102J5_124_3590_U430 ( .A(DP_OP_102J5_124_3590_n2251), .B(
        DP_OP_102J5_124_3590_n1592), .CI(DP_OP_102J5_124_3590_n1987), .CO(
        DP_OP_102J5_124_3590_n684), .S(DP_OP_102J5_124_3590_n685) );
  FADDX1_HVT DP_OP_102J5_124_3590_U429 ( .A(DP_OP_102J5_124_3590_n2052), .B(
        DP_OP_102J5_124_3590_n1657), .CI(DP_OP_102J5_124_3590_n1636), .CO(
        DP_OP_102J5_124_3590_n682), .S(DP_OP_102J5_124_3590_n683) );
  FADDX1_HVT DP_OP_102J5_124_3590_U428 ( .A(DP_OP_102J5_124_3590_n2163), .B(
        DP_OP_102J5_124_3590_n2140), .CI(DP_OP_102J5_124_3590_n1920), .CO(
        DP_OP_102J5_124_3590_n680), .S(DP_OP_102J5_124_3590_n681) );
  FADDX1_HVT DP_OP_102J5_124_3590_U427 ( .A(DP_OP_102J5_124_3590_n1724), .B(
        DP_OP_102J5_124_3590_n2184), .CI(DP_OP_102J5_124_3590_n2207), .CO(
        DP_OP_102J5_124_3590_n678), .S(DP_OP_102J5_124_3590_n679) );
  FADDX1_HVT DP_OP_102J5_124_3590_U426 ( .A(DP_OP_102J5_124_3590_n2096), .B(
        DP_OP_102J5_124_3590_n2075), .CI(DP_OP_102J5_124_3590_n2272), .CO(
        DP_OP_102J5_124_3590_n676), .S(DP_OP_102J5_124_3590_n677) );
  FADDX1_HVT DP_OP_102J5_124_3590_U425 ( .A(DP_OP_102J5_124_3590_n1745), .B(
        DP_OP_102J5_124_3590_n2295), .CI(DP_OP_102J5_124_3590_n1525), .CO(
        DP_OP_102J5_124_3590_n674), .S(DP_OP_102J5_124_3590_n675) );
  FADDX1_HVT DP_OP_102J5_124_3590_U424 ( .A(DP_OP_102J5_124_3590_n1774), .B(
        DP_OP_102J5_124_3590_n1467), .CI(DP_OP_102J5_124_3590_n701), .CO(
        DP_OP_102J5_124_3590_n672), .S(DP_OP_102J5_124_3590_n673) );
  FADDX1_HVT DP_OP_102J5_124_3590_U423 ( .A(DP_OP_102J5_124_3590_n2309), .B(
        DP_OP_102J5_124_3590_n1474), .CI(DP_OP_102J5_124_3590_n2302), .CO(
        DP_OP_102J5_124_3590_n670), .S(DP_OP_102J5_124_3590_n671) );
  FADDX1_HVT DP_OP_102J5_124_3590_U422 ( .A(DP_OP_102J5_124_3590_n1950), .B(
        DP_OP_102J5_124_3590_n1511), .CI(DP_OP_102J5_124_3590_n2265), .CO(
        DP_OP_102J5_124_3590_n668), .S(DP_OP_102J5_124_3590_n669) );
  FADDX1_HVT DP_OP_102J5_124_3590_U421 ( .A(DP_OP_102J5_124_3590_n2258), .B(
        DP_OP_102J5_124_3590_n1518), .CI(DP_OP_102J5_124_3590_n1555), .CO(
        DP_OP_102J5_124_3590_n666), .S(DP_OP_102J5_124_3590_n667) );
  FADDX1_HVT DP_OP_102J5_124_3590_U420 ( .A(DP_OP_102J5_124_3590_n2221), .B(
        DP_OP_102J5_124_3590_n1562), .CI(DP_OP_102J5_124_3590_n1599), .CO(
        DP_OP_102J5_124_3590_n664), .S(DP_OP_102J5_124_3590_n665) );
  FADDX1_HVT DP_OP_102J5_124_3590_U419 ( .A(DP_OP_102J5_124_3590_n2214), .B(
        DP_OP_102J5_124_3590_n1606), .CI(DP_OP_102J5_124_3590_n1643), .CO(
        DP_OP_102J5_124_3590_n662), .S(DP_OP_102J5_124_3590_n663) );
  FADDX1_HVT DP_OP_102J5_124_3590_U418 ( .A(DP_OP_102J5_124_3590_n2177), .B(
        DP_OP_102J5_124_3590_n1650), .CI(DP_OP_102J5_124_3590_n1687), .CO(
        DP_OP_102J5_124_3590_n660), .S(DP_OP_102J5_124_3590_n661) );
  FADDX1_HVT DP_OP_102J5_124_3590_U417 ( .A(DP_OP_102J5_124_3590_n2170), .B(
        DP_OP_102J5_124_3590_n1694), .CI(DP_OP_102J5_124_3590_n1731), .CO(
        DP_OP_102J5_124_3590_n658), .S(DP_OP_102J5_124_3590_n659) );
  FADDX1_HVT DP_OP_102J5_124_3590_U416 ( .A(DP_OP_102J5_124_3590_n2133), .B(
        DP_OP_102J5_124_3590_n1738), .CI(DP_OP_102J5_124_3590_n1781), .CO(
        DP_OP_102J5_124_3590_n656), .S(DP_OP_102J5_124_3590_n657) );
  FADDX1_HVT DP_OP_102J5_124_3590_U415 ( .A(DP_OP_102J5_124_3590_n2126), .B(
        DP_OP_102J5_124_3590_n1818), .CI(DP_OP_102J5_124_3590_n1825), .CO(
        DP_OP_102J5_124_3590_n654), .S(DP_OP_102J5_124_3590_n655) );
  FADDX1_HVT DP_OP_102J5_124_3590_U414 ( .A(DP_OP_102J5_124_3590_n2089), .B(
        DP_OP_102J5_124_3590_n1862), .CI(DP_OP_102J5_124_3590_n1869), .CO(
        DP_OP_102J5_124_3590_n652), .S(DP_OP_102J5_124_3590_n653) );
  FADDX1_HVT DP_OP_102J5_124_3590_U413 ( .A(DP_OP_102J5_124_3590_n2082), .B(
        DP_OP_102J5_124_3590_n1906), .CI(DP_OP_102J5_124_3590_n1913), .CO(
        DP_OP_102J5_124_3590_n650), .S(DP_OP_102J5_124_3590_n651) );
  FADDX1_HVT DP_OP_102J5_124_3590_U412 ( .A(DP_OP_102J5_124_3590_n2045), .B(
        DP_OP_102J5_124_3590_n1957), .CI(DP_OP_102J5_124_3590_n1994), .CO(
        DP_OP_102J5_124_3590_n648), .S(DP_OP_102J5_124_3590_n649) );
  FADDX1_HVT DP_OP_102J5_124_3590_U411 ( .A(DP_OP_102J5_124_3590_n2038), .B(
        DP_OP_102J5_124_3590_n2001), .CI(DP_OP_102J5_124_3590_n848), .CO(
        DP_OP_102J5_124_3590_n646), .S(DP_OP_102J5_124_3590_n647) );
  FADDX1_HVT DP_OP_102J5_124_3590_U410 ( .A(DP_OP_102J5_124_3590_n846), .B(
        DP_OP_102J5_124_3590_n842), .CI(DP_OP_102J5_124_3590_n850), .CO(
        DP_OP_102J5_124_3590_n644), .S(DP_OP_102J5_124_3590_n645) );
  FADDX1_HVT DP_OP_102J5_124_3590_U409 ( .A(DP_OP_102J5_124_3590_n854), .B(
        DP_OP_102J5_124_3590_n844), .CI(DP_OP_102J5_124_3590_n852), .CO(
        DP_OP_102J5_124_3590_n642), .S(DP_OP_102J5_124_3590_n643) );
  FADDX1_HVT DP_OP_102J5_124_3590_U408 ( .A(DP_OP_102J5_124_3590_n824), .B(
        DP_OP_102J5_124_3590_n806), .CI(DP_OP_102J5_124_3590_n802), .CO(
        DP_OP_102J5_124_3590_n640), .S(DP_OP_102J5_124_3590_n641) );
  FADDX1_HVT DP_OP_102J5_124_3590_U407 ( .A(DP_OP_102J5_124_3590_n822), .B(
        DP_OP_102J5_124_3590_n804), .CI(DP_OP_102J5_124_3590_n808), .CO(
        DP_OP_102J5_124_3590_n638), .S(DP_OP_102J5_124_3590_n639) );
  FADDX1_HVT DP_OP_102J5_124_3590_U406 ( .A(DP_OP_102J5_124_3590_n818), .B(
        DP_OP_102J5_124_3590_n812), .CI(DP_OP_102J5_124_3590_n810), .CO(
        DP_OP_102J5_124_3590_n636), .S(DP_OP_102J5_124_3590_n637) );
  FADDX1_HVT DP_OP_102J5_124_3590_U405 ( .A(DP_OP_102J5_124_3590_n820), .B(
        DP_OP_102J5_124_3590_n814), .CI(DP_OP_102J5_124_3590_n826), .CO(
        DP_OP_102J5_124_3590_n634), .S(DP_OP_102J5_124_3590_n635) );
  FADDX1_HVT DP_OP_102J5_124_3590_U404 ( .A(DP_OP_102J5_124_3590_n816), .B(
        DP_OP_102J5_124_3590_n828), .CI(DP_OP_102J5_124_3590_n832), .CO(
        DP_OP_102J5_124_3590_n632), .S(DP_OP_102J5_124_3590_n633) );
  FADDX1_HVT DP_OP_102J5_124_3590_U403 ( .A(DP_OP_102J5_124_3590_n836), .B(
        DP_OP_102J5_124_3590_n830), .CI(DP_OP_102J5_124_3590_n838), .CO(
        DP_OP_102J5_124_3590_n630), .S(DP_OP_102J5_124_3590_n631) );
  FADDX1_HVT DP_OP_102J5_124_3590_U402 ( .A(DP_OP_102J5_124_3590_n840), .B(
        DP_OP_102J5_124_3590_n834), .CI(DP_OP_102J5_124_3590_n693), .CO(
        DP_OP_102J5_124_3590_n628), .S(DP_OP_102J5_124_3590_n629) );
  FADDX1_HVT DP_OP_102J5_124_3590_U401 ( .A(DP_OP_102J5_124_3590_n689), .B(
        DP_OP_102J5_124_3590_n677), .CI(DP_OP_102J5_124_3590_n675), .CO(
        DP_OP_102J5_124_3590_n626), .S(DP_OP_102J5_124_3590_n627) );
  FADDX1_HVT DP_OP_102J5_124_3590_U400 ( .A(DP_OP_102J5_124_3590_n691), .B(
        DP_OP_102J5_124_3590_n687), .CI(DP_OP_102J5_124_3590_n683), .CO(
        DP_OP_102J5_124_3590_n624), .S(DP_OP_102J5_124_3590_n625) );
  FADDX1_HVT DP_OP_102J5_124_3590_U399 ( .A(DP_OP_102J5_124_3590_n695), .B(
        DP_OP_102J5_124_3590_n679), .CI(DP_OP_102J5_124_3590_n681), .CO(
        DP_OP_102J5_124_3590_n622), .S(DP_OP_102J5_124_3590_n623) );
  FADDX1_HVT DP_OP_102J5_124_3590_U398 ( .A(DP_OP_102J5_124_3590_n697), .B(
        DP_OP_102J5_124_3590_n699), .CI(DP_OP_102J5_124_3590_n685), .CO(
        DP_OP_102J5_124_3590_n620), .S(DP_OP_102J5_124_3590_n621) );
  FADDX1_HVT DP_OP_102J5_124_3590_U397 ( .A(DP_OP_102J5_124_3590_n667), .B(
        DP_OP_102J5_124_3590_n665), .CI(DP_OP_102J5_124_3590_n661), .CO(
        DP_OP_102J5_124_3590_n618), .S(DP_OP_102J5_124_3590_n619) );
  FADDX1_HVT DP_OP_102J5_124_3590_U396 ( .A(DP_OP_102J5_124_3590_n669), .B(
        DP_OP_102J5_124_3590_n651), .CI(DP_OP_102J5_124_3590_n649), .CO(
        DP_OP_102J5_124_3590_n616), .S(DP_OP_102J5_124_3590_n617) );
  FADDX1_HVT DP_OP_102J5_124_3590_U395 ( .A(DP_OP_102J5_124_3590_n659), .B(
        DP_OP_102J5_124_3590_n657), .CI(DP_OP_102J5_124_3590_n653), .CO(
        DP_OP_102J5_124_3590_n614), .S(DP_OP_102J5_124_3590_n615) );
  FADDX1_HVT DP_OP_102J5_124_3590_U394 ( .A(DP_OP_102J5_124_3590_n663), .B(
        DP_OP_102J5_124_3590_n673), .CI(DP_OP_102J5_124_3590_n671), .CO(
        DP_OP_102J5_124_3590_n612), .S(DP_OP_102J5_124_3590_n613) );
  FADDX1_HVT DP_OP_102J5_124_3590_U393 ( .A(DP_OP_102J5_124_3590_n655), .B(
        DP_OP_102J5_124_3590_n798), .CI(DP_OP_102J5_124_3590_n800), .CO(
        DP_OP_102J5_124_3590_n610), .S(DP_OP_102J5_124_3590_n611) );
  FADDX1_HVT DP_OP_102J5_124_3590_U392 ( .A(DP_OP_102J5_124_3590_n788), .B(
        DP_OP_102J5_124_3590_n790), .CI(DP_OP_102J5_124_3590_n647), .CO(
        DP_OP_102J5_124_3590_n608), .S(DP_OP_102J5_124_3590_n609) );
  FADDX1_HVT DP_OP_102J5_124_3590_U391 ( .A(DP_OP_102J5_124_3590_n794), .B(
        DP_OP_102J5_124_3590_n786), .CI(DP_OP_102J5_124_3590_n1425), .CO(
        DP_OP_102J5_124_3590_n606), .S(DP_OP_102J5_124_3590_n607) );
  FADDX1_HVT DP_OP_102J5_124_3590_U390 ( .A(DP_OP_102J5_124_3590_n796), .B(
        DP_OP_102J5_124_3590_n792), .CI(DP_OP_102J5_124_3590_n784), .CO(
        DP_OP_102J5_124_3590_n604), .S(DP_OP_102J5_124_3590_n605) );
  FADDX1_HVT DP_OP_102J5_124_3590_U389 ( .A(DP_OP_102J5_124_3590_n782), .B(
        DP_OP_102J5_124_3590_n780), .CI(DP_OP_102J5_124_3590_n645), .CO(
        DP_OP_102J5_124_3590_n602), .S(DP_OP_102J5_124_3590_n603) );
  FADDX1_HVT DP_OP_102J5_124_3590_U388 ( .A(DP_OP_102J5_124_3590_n643), .B(
        DP_OP_102J5_124_3590_n639), .CI(DP_OP_102J5_124_3590_n635), .CO(
        DP_OP_102J5_124_3590_n600), .S(DP_OP_102J5_124_3590_n601) );
  FADDX1_HVT DP_OP_102J5_124_3590_U387 ( .A(DP_OP_102J5_124_3590_n637), .B(
        DP_OP_102J5_124_3590_n641), .CI(DP_OP_102J5_124_3590_n629), .CO(
        DP_OP_102J5_124_3590_n598), .S(DP_OP_102J5_124_3590_n599) );
  FADDX1_HVT DP_OP_102J5_124_3590_U386 ( .A(DP_OP_102J5_124_3590_n778), .B(
        DP_OP_102J5_124_3590_n633), .CI(DP_OP_102J5_124_3590_n631), .CO(
        DP_OP_102J5_124_3590_n596), .S(DP_OP_102J5_124_3590_n597) );
  FADDX1_HVT DP_OP_102J5_124_3590_U385 ( .A(DP_OP_102J5_124_3590_n768), .B(
        DP_OP_102J5_124_3590_n776), .CI(DP_OP_102J5_124_3590_n770), .CO(
        DP_OP_102J5_124_3590_n594), .S(DP_OP_102J5_124_3590_n595) );
  FADDX1_HVT DP_OP_102J5_124_3590_U384 ( .A(DP_OP_102J5_124_3590_n774), .B(
        DP_OP_102J5_124_3590_n772), .CI(DP_OP_102J5_124_3590_n623), .CO(
        DP_OP_102J5_124_3590_n592), .S(DP_OP_102J5_124_3590_n593) );
  FADDX1_HVT DP_OP_102J5_124_3590_U383 ( .A(DP_OP_102J5_124_3590_n625), .B(
        DP_OP_102J5_124_3590_n627), .CI(DP_OP_102J5_124_3590_n766), .CO(
        DP_OP_102J5_124_3590_n590), .S(DP_OP_102J5_124_3590_n591) );
  FADDX1_HVT DP_OP_102J5_124_3590_U382 ( .A(DP_OP_102J5_124_3590_n621), .B(
        DP_OP_102J5_124_3590_n615), .CI(DP_OP_102J5_124_3590_n617), .CO(
        DP_OP_102J5_124_3590_n588), .S(DP_OP_102J5_124_3590_n589) );
  FADDX1_HVT DP_OP_102J5_124_3590_U381 ( .A(DP_OP_102J5_124_3590_n613), .B(
        DP_OP_102J5_124_3590_n619), .CI(DP_OP_102J5_124_3590_n764), .CO(
        DP_OP_102J5_124_3590_n586), .S(DP_OP_102J5_124_3590_n587) );
  FADDX1_HVT DP_OP_102J5_124_3590_U380 ( .A(DP_OP_102J5_124_3590_n762), .B(
        DP_OP_102J5_124_3590_n760), .CI(DP_OP_102J5_124_3590_n611), .CO(
        DP_OP_102J5_124_3590_n584), .S(DP_OP_102J5_124_3590_n585) );
  FADDX1_HVT DP_OP_102J5_124_3590_U379 ( .A(DP_OP_102J5_124_3590_n758), .B(
        DP_OP_102J5_124_3590_n756), .CI(DP_OP_102J5_124_3590_n754), .CO(
        DP_OP_102J5_124_3590_n582), .S(DP_OP_102J5_124_3590_n583) );
  FADDX1_HVT DP_OP_102J5_124_3590_U378 ( .A(DP_OP_102J5_124_3590_n752), .B(
        DP_OP_102J5_124_3590_n605), .CI(DP_OP_102J5_124_3590_n609), .CO(
        DP_OP_102J5_124_3590_n580), .S(DP_OP_102J5_124_3590_n581) );
  FADDX1_HVT DP_OP_102J5_124_3590_U377 ( .A(DP_OP_102J5_124_3590_n750), .B(
        DP_OP_102J5_124_3590_n607), .CI(DP_OP_102J5_124_3590_n748), .CO(
        DP_OP_102J5_124_3590_n578), .S(DP_OP_102J5_124_3590_n579) );
  FADDX1_HVT DP_OP_102J5_124_3590_U376 ( .A(DP_OP_102J5_124_3590_n746), .B(
        DP_OP_102J5_124_3590_n603), .CI(DP_OP_102J5_124_3590_n601), .CO(
        DP_OP_102J5_124_3590_n576), .S(DP_OP_102J5_124_3590_n577) );
  FADDX1_HVT DP_OP_102J5_124_3590_U375 ( .A(DP_OP_102J5_124_3590_n744), .B(
        DP_OP_102J5_124_3590_n597), .CI(DP_OP_102J5_124_3590_n593), .CO(
        DP_OP_102J5_124_3590_n574), .S(DP_OP_102J5_124_3590_n575) );
  FADDX1_HVT DP_OP_102J5_124_3590_U374 ( .A(DP_OP_102J5_124_3590_n742), .B(
        DP_OP_102J5_124_3590_n595), .CI(DP_OP_102J5_124_3590_n599), .CO(
        DP_OP_102J5_124_3590_n572), .S(DP_OP_102J5_124_3590_n573) );
  FADDX1_HVT DP_OP_102J5_124_3590_U373 ( .A(DP_OP_102J5_124_3590_n740), .B(
        DP_OP_102J5_124_3590_n591), .CI(DP_OP_102J5_124_3590_n589), .CO(
        DP_OP_102J5_124_3590_n570), .S(DP_OP_102J5_124_3590_n571) );
  FADDX1_HVT DP_OP_102J5_124_3590_U372 ( .A(DP_OP_102J5_124_3590_n738), .B(
        DP_OP_102J5_124_3590_n587), .CI(DP_OP_102J5_124_3590_n736), .CO(
        DP_OP_102J5_124_3590_n568), .S(DP_OP_102J5_124_3590_n569) );
  FADDX1_HVT DP_OP_102J5_124_3590_U371 ( .A(DP_OP_102J5_124_3590_n734), .B(
        DP_OP_102J5_124_3590_n585), .CI(DP_OP_102J5_124_3590_n732), .CO(
        DP_OP_102J5_124_3590_n566), .S(DP_OP_102J5_124_3590_n567) );
  FADDX1_HVT DP_OP_102J5_124_3590_U370 ( .A(DP_OP_102J5_124_3590_n583), .B(
        DP_OP_102J5_124_3590_n730), .CI(DP_OP_102J5_124_3590_n728), .CO(
        DP_OP_102J5_124_3590_n564), .S(DP_OP_102J5_124_3590_n565) );
  FADDX1_HVT DP_OP_102J5_124_3590_U369 ( .A(DP_OP_102J5_124_3590_n581), .B(
        DP_OP_102J5_124_3590_n579), .CI(DP_OP_102J5_124_3590_n726), .CO(
        DP_OP_102J5_124_3590_n562), .S(DP_OP_102J5_124_3590_n563) );
  FADDX1_HVT DP_OP_102J5_124_3590_U368 ( .A(DP_OP_102J5_124_3590_n577), .B(
        DP_OP_102J5_124_3590_n573), .CI(DP_OP_102J5_124_3590_n575), .CO(
        DP_OP_102J5_124_3590_n560), .S(DP_OP_102J5_124_3590_n561) );
  FADDX1_HVT DP_OP_102J5_124_3590_U367 ( .A(DP_OP_102J5_124_3590_n724), .B(
        DP_OP_102J5_124_3590_n722), .CI(DP_OP_102J5_124_3590_n571), .CO(
        DP_OP_102J5_124_3590_n558), .S(DP_OP_102J5_124_3590_n559) );
  FADDX1_HVT DP_OP_102J5_124_3590_U366 ( .A(DP_OP_102J5_124_3590_n569), .B(
        DP_OP_102J5_124_3590_n720), .CI(DP_OP_102J5_124_3590_n718), .CO(
        DP_OP_102J5_124_3590_n556), .S(DP_OP_102J5_124_3590_n557) );
  FADDX1_HVT DP_OP_102J5_124_3590_U365 ( .A(DP_OP_102J5_124_3590_n567), .B(
        DP_OP_102J5_124_3590_n716), .CI(DP_OP_102J5_124_3590_n565), .CO(
        DP_OP_102J5_124_3590_n554), .S(DP_OP_102J5_124_3590_n555) );
  FADDX1_HVT DP_OP_102J5_124_3590_U364 ( .A(DP_OP_102J5_124_3590_n563), .B(
        DP_OP_102J5_124_3590_n714), .CI(DP_OP_102J5_124_3590_n561), .CO(
        DP_OP_102J5_124_3590_n552), .S(DP_OP_102J5_124_3590_n553) );
  FADDX1_HVT DP_OP_102J5_124_3590_U363 ( .A(DP_OP_102J5_124_3590_n712), .B(
        DP_OP_102J5_124_3590_n559), .CI(DP_OP_102J5_124_3590_n710), .CO(
        DP_OP_102J5_124_3590_n550), .S(DP_OP_102J5_124_3590_n551) );
  FADDX1_HVT DP_OP_102J5_124_3590_U362 ( .A(DP_OP_102J5_124_3590_n557), .B(
        DP_OP_102J5_124_3590_n555), .CI(DP_OP_102J5_124_3590_n708), .CO(
        DP_OP_102J5_124_3590_n548), .S(DP_OP_102J5_124_3590_n549) );
  FADDX1_HVT DP_OP_102J5_124_3590_U361 ( .A(DP_OP_102J5_124_3590_n553), .B(
        DP_OP_102J5_124_3590_n706), .CI(DP_OP_102J5_124_3590_n551), .CO(
        DP_OP_102J5_124_3590_n546), .S(DP_OP_102J5_124_3590_n547) );
  FADDX1_HVT DP_OP_102J5_124_3590_U360 ( .A(DP_OP_102J5_124_3590_n704), .B(
        DP_OP_102J5_124_3590_n549), .CI(DP_OP_102J5_124_3590_n547), .CO(
        DP_OP_102J5_124_3590_n544), .S(DP_OP_102J5_124_3590_n545) );
  FADDX1_HVT DP_OP_102J5_124_3590_U359 ( .A(DP_OP_102J5_124_3590_n1868), .B(
        DP_OP_102J5_124_3590_n2308), .CI(DP_OP_102J5_124_3590_n1459), .CO(
        DP_OP_102J5_124_3590_n542), .S(DP_OP_102J5_124_3590_n543) );
  FADDX1_HVT DP_OP_102J5_124_3590_U358 ( .A(DP_OP_102J5_124_3590_n700), .B(
        DP_OP_102J5_124_3590_n1547), .CI(DP_OP_102J5_124_3590_n1473), .CO(
        DP_OP_102J5_124_3590_n540), .S(DP_OP_102J5_124_3590_n541) );
  FADDX1_HVT DP_OP_102J5_124_3590_U357 ( .A(DP_OP_102J5_124_3590_n1723), .B(
        DP_OP_102J5_124_3590_n1503), .CI(DP_OP_102J5_124_3590_n1561), .CO(
        DP_OP_102J5_124_3590_n538), .S(DP_OP_102J5_124_3590_n539) );
  FADDX1_HVT DP_OP_102J5_124_3590_U356 ( .A(DP_OP_102J5_124_3590_n2088), .B(
        DP_OP_102J5_124_3590_n1780), .CI(DP_OP_102J5_124_3590_n1635), .CO(
        DP_OP_102J5_124_3590_n536), .S(DP_OP_102J5_124_3590_n537) );
  FADDX1_HVT DP_OP_102J5_124_3590_U355 ( .A(DP_OP_102J5_124_3590_n1824), .B(
        DP_OP_102J5_124_3590_n1737), .CI(DP_OP_102J5_124_3590_n1810), .CO(
        DP_OP_102J5_124_3590_n534), .S(DP_OP_102J5_124_3590_n535) );
  FADDX1_HVT DP_OP_102J5_124_3590_U354 ( .A(DP_OP_102J5_124_3590_n1854), .B(
        DP_OP_102J5_124_3590_n1766), .CI(DP_OP_102J5_124_3590_n1912), .CO(
        DP_OP_102J5_124_3590_n532), .S(DP_OP_102J5_124_3590_n533) );
  FADDX1_HVT DP_OP_102J5_124_3590_U353 ( .A(DP_OP_102J5_124_3590_n1517), .B(
        DP_OP_102J5_124_3590_n1591), .CI(DP_OP_102J5_124_3590_n1693), .CO(
        DP_OP_102J5_124_3590_n530), .S(DP_OP_102J5_124_3590_n531) );
  FADDX1_HVT DP_OP_102J5_124_3590_U352 ( .A(DP_OP_102J5_124_3590_n1898), .B(
        DP_OP_102J5_124_3590_n1986), .CI(DP_OP_102J5_124_3590_n1956), .CO(
        DP_OP_102J5_124_3590_n528), .S(DP_OP_102J5_124_3590_n529) );
  FADDX1_HVT DP_OP_102J5_124_3590_U351 ( .A(DP_OP_102J5_124_3590_n2132), .B(
        DP_OP_102J5_124_3590_n2030), .CI(DP_OP_102J5_124_3590_n1649), .CO(
        DP_OP_102J5_124_3590_n526), .S(DP_OP_102J5_124_3590_n527) );
  FADDX1_HVT DP_OP_102J5_124_3590_U350 ( .A(DP_OP_102J5_124_3590_n2074), .B(
        DP_OP_102J5_124_3590_n2118), .CI(DP_OP_102J5_124_3590_n2000), .CO(
        DP_OP_102J5_124_3590_n524), .S(DP_OP_102J5_124_3590_n525) );
  FADDX1_HVT DP_OP_102J5_124_3590_U349 ( .A(DP_OP_102J5_124_3590_n2044), .B(
        DP_OP_102J5_124_3590_n1679), .CI(DP_OP_102J5_124_3590_n2176), .CO(
        DP_OP_102J5_124_3590_n522), .S(DP_OP_102J5_124_3590_n523) );
  FADDX1_HVT DP_OP_102J5_124_3590_U348 ( .A(DP_OP_102J5_124_3590_n2220), .B(
        DP_OP_102J5_124_3590_n1942), .CI(DP_OP_102J5_124_3590_n1605), .CO(
        DP_OP_102J5_124_3590_n520), .S(DP_OP_102J5_124_3590_n521) );
  FADDX1_HVT DP_OP_102J5_124_3590_U347 ( .A(DP_OP_102J5_124_3590_n2264), .B(
        DP_OP_102J5_124_3590_n2250), .CI(DP_OP_102J5_124_3590_n2162), .CO(
        DP_OP_102J5_124_3590_n518), .S(DP_OP_102J5_124_3590_n519) );
  FADDX1_HVT DP_OP_102J5_124_3590_U346 ( .A(DP_OP_102J5_124_3590_n2206), .B(
        DP_OP_102J5_124_3590_n2294), .CI(DP_OP_102J5_124_3590_n1730), .CO(
        DP_OP_102J5_124_3590_n516), .S(DP_OP_102J5_124_3590_n517) );
  FADDX1_HVT DP_OP_102J5_124_3590_U345 ( .A(DP_OP_102J5_124_3590_n1642), .B(
        DP_OP_102J5_124_3590_n1466), .CI(DP_OP_102J5_124_3590_n1510), .CO(
        DP_OP_102J5_124_3590_n514), .S(DP_OP_102J5_124_3590_n515) );
  FADDX1_HVT DP_OP_102J5_124_3590_U344 ( .A(DP_OP_102J5_124_3590_n2301), .B(
        DP_OP_102J5_124_3590_n1554), .CI(DP_OP_102J5_124_3590_n1598), .CO(
        DP_OP_102J5_124_3590_n512), .S(DP_OP_102J5_124_3590_n513) );
  FADDX1_HVT DP_OP_102J5_124_3590_U343 ( .A(DP_OP_102J5_124_3590_n2257), .B(
        DP_OP_102J5_124_3590_n1686), .CI(DP_OP_102J5_124_3590_n1773), .CO(
        DP_OP_102J5_124_3590_n510), .S(DP_OP_102J5_124_3590_n511) );
  FADDX1_HVT DP_OP_102J5_124_3590_U342 ( .A(DP_OP_102J5_124_3590_n2213), .B(
        DP_OP_102J5_124_3590_n1817), .CI(DP_OP_102J5_124_3590_n1861), .CO(
        DP_OP_102J5_124_3590_n508), .S(DP_OP_102J5_124_3590_n509) );
  FADDX1_HVT DP_OP_102J5_124_3590_U341 ( .A(DP_OP_102J5_124_3590_n2169), .B(
        DP_OP_102J5_124_3590_n1905), .CI(DP_OP_102J5_124_3590_n1949), .CO(
        DP_OP_102J5_124_3590_n506), .S(DP_OP_102J5_124_3590_n507) );
  FADDX1_HVT DP_OP_102J5_124_3590_U340 ( .A(DP_OP_102J5_124_3590_n2125), .B(
        DP_OP_102J5_124_3590_n1993), .CI(DP_OP_102J5_124_3590_n2037), .CO(
        DP_OP_102J5_124_3590_n504), .S(DP_OP_102J5_124_3590_n505) );
  FADDX1_HVT DP_OP_102J5_124_3590_U339 ( .A(DP_OP_102J5_124_3590_n2081), .B(
        DP_OP_102J5_124_3590_n682), .CI(DP_OP_102J5_124_3590_n684), .CO(
        DP_OP_102J5_124_3590_n502), .S(DP_OP_102J5_124_3590_n503) );
  FADDX1_HVT DP_OP_102J5_124_3590_U338 ( .A(DP_OP_102J5_124_3590_n674), .B(
        DP_OP_102J5_124_3590_n678), .CI(DP_OP_102J5_124_3590_n676), .CO(
        DP_OP_102J5_124_3590_n500), .S(DP_OP_102J5_124_3590_n501) );
  FADDX1_HVT DP_OP_102J5_124_3590_U337 ( .A(DP_OP_102J5_124_3590_n692), .B(
        DP_OP_102J5_124_3590_n680), .CI(DP_OP_102J5_124_3590_n686), .CO(
        DP_OP_102J5_124_3590_n498), .S(DP_OP_102J5_124_3590_n499) );
  FADDX1_HVT DP_OP_102J5_124_3590_U336 ( .A(DP_OP_102J5_124_3590_n694), .B(
        DP_OP_102J5_124_3590_n688), .CI(DP_OP_102J5_124_3590_n696), .CO(
        DP_OP_102J5_124_3590_n496), .S(DP_OP_102J5_124_3590_n497) );
  FADDX1_HVT DP_OP_102J5_124_3590_U335 ( .A(DP_OP_102J5_124_3590_n698), .B(
        DP_OP_102J5_124_3590_n690), .CI(DP_OP_102J5_124_3590_n660), .CO(
        DP_OP_102J5_124_3590_n494), .S(DP_OP_102J5_124_3590_n495) );
  FADDX1_HVT DP_OP_102J5_124_3590_U334 ( .A(DP_OP_102J5_124_3590_n656), .B(
        DP_OP_102J5_124_3590_n650), .CI(DP_OP_102J5_124_3590_n648), .CO(
        DP_OP_102J5_124_3590_n492), .S(DP_OP_102J5_124_3590_n493) );
  FADDX1_HVT DP_OP_102J5_124_3590_U333 ( .A(DP_OP_102J5_124_3590_n658), .B(
        DP_OP_102J5_124_3590_n652), .CI(DP_OP_102J5_124_3590_n662), .CO(
        DP_OP_102J5_124_3590_n490), .S(DP_OP_102J5_124_3590_n491) );
  FADDX1_HVT DP_OP_102J5_124_3590_U332 ( .A(DP_OP_102J5_124_3590_n668), .B(
        DP_OP_102J5_124_3590_n654), .CI(DP_OP_102J5_124_3590_n666), .CO(
        DP_OP_102J5_124_3590_n488), .S(DP_OP_102J5_124_3590_n489) );
  FADDX1_HVT DP_OP_102J5_124_3590_U331 ( .A(DP_OP_102J5_124_3590_n670), .B(
        DP_OP_102J5_124_3590_n672), .CI(DP_OP_102J5_124_3590_n664), .CO(
        DP_OP_102J5_124_3590_n486), .S(DP_OP_102J5_124_3590_n487) );
  FADDX1_HVT DP_OP_102J5_124_3590_U330 ( .A(DP_OP_102J5_124_3590_n537), .B(
        DP_OP_102J5_124_3590_n533), .CI(DP_OP_102J5_124_3590_n517), .CO(
        DP_OP_102J5_124_3590_n484), .S(DP_OP_102J5_124_3590_n485) );
  FADDX1_HVT DP_OP_102J5_124_3590_U329 ( .A(DP_OP_102J5_124_3590_n539), .B(
        DP_OP_102J5_124_3590_n531), .CI(DP_OP_102J5_124_3590_n523), .CO(
        DP_OP_102J5_124_3590_n482), .S(DP_OP_102J5_124_3590_n483) );
  FADDX1_HVT DP_OP_102J5_124_3590_U328 ( .A(DP_OP_102J5_124_3590_n535), .B(
        DP_OP_102J5_124_3590_n519), .CI(DP_OP_102J5_124_3590_n527), .CO(
        DP_OP_102J5_124_3590_n480), .S(DP_OP_102J5_124_3590_n481) );
  FADDX1_HVT DP_OP_102J5_124_3590_U327 ( .A(DP_OP_102J5_124_3590_n525), .B(
        DP_OP_102J5_124_3590_n521), .CI(DP_OP_102J5_124_3590_n529), .CO(
        DP_OP_102J5_124_3590_n478), .S(DP_OP_102J5_124_3590_n479) );
  FADDX1_HVT DP_OP_102J5_124_3590_U326 ( .A(DP_OP_102J5_124_3590_n541), .B(
        DP_OP_102J5_124_3590_n543), .CI(DP_OP_102J5_124_3590_n513), .CO(
        DP_OP_102J5_124_3590_n476), .S(DP_OP_102J5_124_3590_n477) );
  FADDX1_HVT DP_OP_102J5_124_3590_U325 ( .A(DP_OP_102J5_124_3590_n507), .B(
        DP_OP_102J5_124_3590_n515), .CI(DP_OP_102J5_124_3590_n511), .CO(
        DP_OP_102J5_124_3590_n474), .S(DP_OP_102J5_124_3590_n475) );
  FADDX1_HVT DP_OP_102J5_124_3590_U324 ( .A(DP_OP_102J5_124_3590_n505), .B(
        DP_OP_102J5_124_3590_n509), .CI(DP_OP_102J5_124_3590_n646), .CO(
        DP_OP_102J5_124_3590_n472), .S(DP_OP_102J5_124_3590_n473) );
  FADDX1_HVT DP_OP_102J5_124_3590_U323 ( .A(DP_OP_102J5_124_3590_n642), .B(
        DP_OP_102J5_124_3590_n644), .CI(DP_OP_102J5_124_3590_n630), .CO(
        DP_OP_102J5_124_3590_n470), .S(DP_OP_102J5_124_3590_n471) );
  FADDX1_HVT DP_OP_102J5_124_3590_U322 ( .A(DP_OP_102J5_124_3590_n636), .B(
        DP_OP_102J5_124_3590_n632), .CI(DP_OP_102J5_124_3590_n1424), .CO(
        DP_OP_102J5_124_3590_n468), .S(DP_OP_102J5_124_3590_n469) );
  FADDX1_HVT DP_OP_102J5_124_3590_U321 ( .A(DP_OP_102J5_124_3590_n638), .B(
        DP_OP_102J5_124_3590_n640), .CI(DP_OP_102J5_124_3590_n628), .CO(
        DP_OP_102J5_124_3590_n466), .S(DP_OP_102J5_124_3590_n467) );
  FADDX1_HVT DP_OP_102J5_124_3590_U320 ( .A(DP_OP_102J5_124_3590_n634), .B(
        DP_OP_102J5_124_3590_n503), .CI(DP_OP_102J5_124_3590_n626), .CO(
        DP_OP_102J5_124_3590_n464), .S(DP_OP_102J5_124_3590_n465) );
  FADDX1_HVT DP_OP_102J5_124_3590_U319 ( .A(DP_OP_102J5_124_3590_n499), .B(
        DP_OP_102J5_124_3590_n624), .CI(DP_OP_102J5_124_3590_n495), .CO(
        DP_OP_102J5_124_3590_n462), .S(DP_OP_102J5_124_3590_n463) );
  FADDX1_HVT DP_OP_102J5_124_3590_U318 ( .A(DP_OP_102J5_124_3590_n497), .B(
        DP_OP_102J5_124_3590_n622), .CI(DP_OP_102J5_124_3590_n620), .CO(
        DP_OP_102J5_124_3590_n460), .S(DP_OP_102J5_124_3590_n461) );
  FADDX1_HVT DP_OP_102J5_124_3590_U317 ( .A(DP_OP_102J5_124_3590_n501), .B(
        DP_OP_102J5_124_3590_n491), .CI(DP_OP_102J5_124_3590_n618), .CO(
        DP_OP_102J5_124_3590_n458), .S(DP_OP_102J5_124_3590_n459) );
  FADDX1_HVT DP_OP_102J5_124_3590_U316 ( .A(DP_OP_102J5_124_3590_n616), .B(
        DP_OP_102J5_124_3590_n489), .CI(DP_OP_102J5_124_3590_n487), .CO(
        DP_OP_102J5_124_3590_n456), .S(DP_OP_102J5_124_3590_n457) );
  FADDX1_HVT DP_OP_102J5_124_3590_U315 ( .A(DP_OP_102J5_124_3590_n614), .B(
        DP_OP_102J5_124_3590_n493), .CI(DP_OP_102J5_124_3590_n612), .CO(
        DP_OP_102J5_124_3590_n454), .S(DP_OP_102J5_124_3590_n455) );
  FADDX1_HVT DP_OP_102J5_124_3590_U314 ( .A(DP_OP_102J5_124_3590_n481), .B(
        DP_OP_102J5_124_3590_n477), .CI(DP_OP_102J5_124_3590_n610), .CO(
        DP_OP_102J5_124_3590_n452), .S(DP_OP_102J5_124_3590_n453) );
  FADDX1_HVT DP_OP_102J5_124_3590_U313 ( .A(DP_OP_102J5_124_3590_n479), .B(
        DP_OP_102J5_124_3590_n485), .CI(DP_OP_102J5_124_3590_n483), .CO(
        DP_OP_102J5_124_3590_n450), .S(DP_OP_102J5_124_3590_n451) );
  FADDX1_HVT DP_OP_102J5_124_3590_U312 ( .A(DP_OP_102J5_124_3590_n475), .B(
        DP_OP_102J5_124_3590_n473), .CI(DP_OP_102J5_124_3590_n608), .CO(
        DP_OP_102J5_124_3590_n448), .S(DP_OP_102J5_124_3590_n449) );
  FADDX1_HVT DP_OP_102J5_124_3590_U311 ( .A(DP_OP_102J5_124_3590_n606), .B(
        DP_OP_102J5_124_3590_n604), .CI(DP_OP_102J5_124_3590_n602), .CO(
        DP_OP_102J5_124_3590_n446), .S(DP_OP_102J5_124_3590_n447) );
  FADDX1_HVT DP_OP_102J5_124_3590_U310 ( .A(DP_OP_102J5_124_3590_n471), .B(
        DP_OP_102J5_124_3590_n600), .CI(DP_OP_102J5_124_3590_n598), .CO(
        DP_OP_102J5_124_3590_n444), .S(DP_OP_102J5_124_3590_n445) );
  FADDX1_HVT DP_OP_102J5_124_3590_U309 ( .A(DP_OP_102J5_124_3590_n596), .B(
        DP_OP_102J5_124_3590_n467), .CI(DP_OP_102J5_124_3590_n465), .CO(
        DP_OP_102J5_124_3590_n442), .S(DP_OP_102J5_124_3590_n443) );
  FADDX1_HVT DP_OP_102J5_124_3590_U308 ( .A(DP_OP_102J5_124_3590_n594), .B(
        DP_OP_102J5_124_3590_n469), .CI(DP_OP_102J5_124_3590_n592), .CO(
        DP_OP_102J5_124_3590_n440), .S(DP_OP_102J5_124_3590_n441) );
  FADDX1_HVT DP_OP_102J5_124_3590_U307 ( .A(DP_OP_102J5_124_3590_n590), .B(
        DP_OP_102J5_124_3590_n463), .CI(DP_OP_102J5_124_3590_n459), .CO(
        DP_OP_102J5_124_3590_n438), .S(DP_OP_102J5_124_3590_n439) );
  FADDX1_HVT DP_OP_102J5_124_3590_U306 ( .A(DP_OP_102J5_124_3590_n461), .B(
        DP_OP_102J5_124_3590_n588), .CI(DP_OP_102J5_124_3590_n586), .CO(
        DP_OP_102J5_124_3590_n436), .S(DP_OP_102J5_124_3590_n437) );
  FADDX1_HVT DP_OP_102J5_124_3590_U305 ( .A(DP_OP_102J5_124_3590_n457), .B(
        DP_OP_102J5_124_3590_n455), .CI(DP_OP_102J5_124_3590_n584), .CO(
        DP_OP_102J5_124_3590_n434), .S(DP_OP_102J5_124_3590_n435) );
  FADDX1_HVT DP_OP_102J5_124_3590_U304 ( .A(DP_OP_102J5_124_3590_n451), .B(
        DP_OP_102J5_124_3590_n453), .CI(DP_OP_102J5_124_3590_n582), .CO(
        DP_OP_102J5_124_3590_n432), .S(DP_OP_102J5_124_3590_n433) );
  FADDX1_HVT DP_OP_102J5_124_3590_U303 ( .A(DP_OP_102J5_124_3590_n449), .B(
        DP_OP_102J5_124_3590_n580), .CI(DP_OP_102J5_124_3590_n578), .CO(
        DP_OP_102J5_124_3590_n430), .S(DP_OP_102J5_124_3590_n431) );
  FADDX1_HVT DP_OP_102J5_124_3590_U302 ( .A(DP_OP_102J5_124_3590_n447), .B(
        DP_OP_102J5_124_3590_n576), .CI(DP_OP_102J5_124_3590_n445), .CO(
        DP_OP_102J5_124_3590_n428), .S(DP_OP_102J5_124_3590_n429) );
  FADDX1_HVT DP_OP_102J5_124_3590_U301 ( .A(DP_OP_102J5_124_3590_n574), .B(
        DP_OP_102J5_124_3590_n443), .CI(DP_OP_102J5_124_3590_n441), .CO(
        DP_OP_102J5_124_3590_n426), .S(DP_OP_102J5_124_3590_n427) );
  FADDX1_HVT DP_OP_102J5_124_3590_U300 ( .A(DP_OP_102J5_124_3590_n572), .B(
        DP_OP_102J5_124_3590_n570), .CI(DP_OP_102J5_124_3590_n439), .CO(
        DP_OP_102J5_124_3590_n424), .S(DP_OP_102J5_124_3590_n425) );
  FADDX1_HVT DP_OP_102J5_124_3590_U299 ( .A(DP_OP_102J5_124_3590_n437), .B(
        DP_OP_102J5_124_3590_n568), .CI(DP_OP_102J5_124_3590_n435), .CO(
        DP_OP_102J5_124_3590_n422), .S(DP_OP_102J5_124_3590_n423) );
  FADDX1_HVT DP_OP_102J5_124_3590_U298 ( .A(DP_OP_102J5_124_3590_n566), .B(
        DP_OP_102J5_124_3590_n433), .CI(DP_OP_102J5_124_3590_n564), .CO(
        DP_OP_102J5_124_3590_n420), .S(DP_OP_102J5_124_3590_n421) );
  FADDX1_HVT DP_OP_102J5_124_3590_U297 ( .A(DP_OP_102J5_124_3590_n431), .B(
        DP_OP_102J5_124_3590_n562), .CI(DP_OP_102J5_124_3590_n429), .CO(
        DP_OP_102J5_124_3590_n418), .S(DP_OP_102J5_124_3590_n419) );
  FADDX1_HVT DP_OP_102J5_124_3590_U296 ( .A(DP_OP_102J5_124_3590_n560), .B(
        DP_OP_102J5_124_3590_n427), .CI(DP_OP_102J5_124_3590_n558), .CO(
        DP_OP_102J5_124_3590_n416), .S(DP_OP_102J5_124_3590_n417) );
  FADDX1_HVT DP_OP_102J5_124_3590_U295 ( .A(DP_OP_102J5_124_3590_n425), .B(
        DP_OP_102J5_124_3590_n423), .CI(DP_OP_102J5_124_3590_n556), .CO(
        DP_OP_102J5_124_3590_n414), .S(DP_OP_102J5_124_3590_n415) );
  FADDX1_HVT DP_OP_102J5_124_3590_U294 ( .A(DP_OP_102J5_124_3590_n421), .B(
        DP_OP_102J5_124_3590_n554), .CI(DP_OP_102J5_124_3590_n419), .CO(
        DP_OP_102J5_124_3590_n412), .S(DP_OP_102J5_124_3590_n413) );
  FADDX1_HVT DP_OP_102J5_124_3590_U293 ( .A(DP_OP_102J5_124_3590_n552), .B(
        DP_OP_102J5_124_3590_n417), .CI(DP_OP_102J5_124_3590_n550), .CO(
        DP_OP_102J5_124_3590_n410), .S(DP_OP_102J5_124_3590_n411) );
  FADDX1_HVT DP_OP_102J5_124_3590_U292 ( .A(DP_OP_102J5_124_3590_n415), .B(
        DP_OP_102J5_124_3590_n548), .CI(DP_OP_102J5_124_3590_n413), .CO(
        DP_OP_102J5_124_3590_n408), .S(DP_OP_102J5_124_3590_n409) );
  FADDX1_HVT DP_OP_102J5_124_3590_U291 ( .A(DP_OP_102J5_124_3590_n546), .B(
        DP_OP_102J5_124_3590_n411), .CI(DP_OP_102J5_124_3590_n409), .CO(
        DP_OP_102J5_124_3590_n406), .S(DP_OP_102J5_124_3590_n407) );
  FADDX1_HVT DP_OP_102J5_124_3590_U289 ( .A(DP_OP_102J5_124_3590_n1729), .B(
        DP_OP_102J5_124_3590_n2300), .CI(DP_OP_102J5_124_3590_n1458), .CO(
        DP_OP_102J5_124_3590_n402), .S(DP_OP_102J5_124_3590_n403) );
  FADDX1_HVT DP_OP_102J5_124_3590_U288 ( .A(DP_OP_102J5_124_3590_n1722), .B(
        DP_OP_102J5_124_3590_n1465), .CI(DP_OP_102J5_124_3590_n2293), .CO(
        DP_OP_102J5_124_3590_n400), .S(DP_OP_102J5_124_3590_n401) );
  FADDX1_HVT DP_OP_102J5_124_3590_U287 ( .A(DP_OP_102J5_124_3590_n1772), .B(
        DP_OP_102J5_124_3590_n1502), .CI(DP_OP_102J5_124_3590_n1509), .CO(
        DP_OP_102J5_124_3590_n398), .S(DP_OP_102J5_124_3590_n399) );
  FADDX1_HVT DP_OP_102J5_124_3590_U286 ( .A(DP_OP_102J5_124_3590_n1634), .B(
        DP_OP_102J5_124_3590_n2256), .CI(DP_OP_102J5_124_3590_n2249), .CO(
        DP_OP_102J5_124_3590_n396), .S(DP_OP_102J5_124_3590_n397) );
  FADDX1_HVT DP_OP_102J5_124_3590_U285 ( .A(DP_OP_102J5_124_3590_n1590), .B(
        DP_OP_102J5_124_3590_n1546), .CI(DP_OP_102J5_124_3590_n1553), .CO(
        DP_OP_102J5_124_3590_n394), .S(DP_OP_102J5_124_3590_n395) );
  FADDX1_HVT DP_OP_102J5_124_3590_U284 ( .A(DP_OP_102J5_124_3590_n2212), .B(
        DP_OP_102J5_124_3590_n2205), .CI(DP_OP_102J5_124_3590_n2168), .CO(
        DP_OP_102J5_124_3590_n392), .S(DP_OP_102J5_124_3590_n393) );
  FADDX1_HVT DP_OP_102J5_124_3590_U283 ( .A(DP_OP_102J5_124_3590_n1941), .B(
        DP_OP_102J5_124_3590_n2161), .CI(DP_OP_102J5_124_3590_n2124), .CO(
        DP_OP_102J5_124_3590_n390), .S(DP_OP_102J5_124_3590_n391) );
  FADDX1_HVT DP_OP_102J5_124_3590_U282 ( .A(DP_OP_102J5_124_3590_n1853), .B(
        DP_OP_102J5_124_3590_n1597), .CI(DP_OP_102J5_124_3590_n2117), .CO(
        DP_OP_102J5_124_3590_n388), .S(DP_OP_102J5_124_3590_n389) );
  FADDX1_HVT DP_OP_102J5_124_3590_U281 ( .A(DP_OP_102J5_124_3590_n1816), .B(
        DP_OP_102J5_124_3590_n1641), .CI(DP_OP_102J5_124_3590_n1678), .CO(
        DP_OP_102J5_124_3590_n386), .S(DP_OP_102J5_124_3590_n387) );
  FADDX1_HVT DP_OP_102J5_124_3590_U280 ( .A(DP_OP_102J5_124_3590_n2080), .B(
        DP_OP_102J5_124_3590_n2073), .CI(DP_OP_102J5_124_3590_n1685), .CO(
        DP_OP_102J5_124_3590_n384), .S(DP_OP_102J5_124_3590_n385) );
  FADDX1_HVT DP_OP_102J5_124_3590_U279 ( .A(DP_OP_102J5_124_3590_n1904), .B(
        DP_OP_102J5_124_3590_n2036), .CI(DP_OP_102J5_124_3590_n2029), .CO(
        DP_OP_102J5_124_3590_n382), .S(DP_OP_102J5_124_3590_n383) );
  FADDX1_HVT DP_OP_102J5_124_3590_U278 ( .A(DP_OP_102J5_124_3590_n1992), .B(
        DP_OP_102J5_124_3590_n1809), .CI(DP_OP_102J5_124_3590_n1860), .CO(
        DP_OP_102J5_124_3590_n380), .S(DP_OP_102J5_124_3590_n381) );
  FADDX1_HVT DP_OP_102J5_124_3590_U277 ( .A(DP_OP_102J5_124_3590_n1985), .B(
        DP_OP_102J5_124_3590_n1897), .CI(DP_OP_102J5_124_3590_n1948), .CO(
        DP_OP_102J5_124_3590_n378), .S(DP_OP_102J5_124_3590_n379) );
  FADDX1_HVT DP_OP_102J5_124_3590_U276 ( .A(DP_OP_102J5_124_3590_n405), .B(
        DP_OP_102J5_124_3590_n516), .CI(DP_OP_102J5_124_3590_n532), .CO(
        DP_OP_102J5_124_3590_n376), .S(DP_OP_102J5_124_3590_n377) );
  FADDX1_HVT DP_OP_102J5_124_3590_U275 ( .A(DP_OP_102J5_124_3590_n526), .B(
        DP_OP_102J5_124_3590_n520), .CI(DP_OP_102J5_124_3590_n522), .CO(
        DP_OP_102J5_124_3590_n374), .S(DP_OP_102J5_124_3590_n375) );
  FADDX1_HVT DP_OP_102J5_124_3590_U274 ( .A(DP_OP_102J5_124_3590_n528), .B(
        DP_OP_102J5_124_3590_n518), .CI(DP_OP_102J5_124_3590_n530), .CO(
        DP_OP_102J5_124_3590_n372), .S(DP_OP_102J5_124_3590_n373) );
  FADDX1_HVT DP_OP_102J5_124_3590_U273 ( .A(DP_OP_102J5_124_3590_n538), .B(
        DP_OP_102J5_124_3590_n524), .CI(DP_OP_102J5_124_3590_n536), .CO(
        DP_OP_102J5_124_3590_n370), .S(DP_OP_102J5_124_3590_n371) );
  FADDX1_HVT DP_OP_102J5_124_3590_U272 ( .A(DP_OP_102J5_124_3590_n540), .B(
        DP_OP_102J5_124_3590_n542), .CI(DP_OP_102J5_124_3590_n534), .CO(
        DP_OP_102J5_124_3590_n368), .S(DP_OP_102J5_124_3590_n369) );
  FADDX1_HVT DP_OP_102J5_124_3590_U271 ( .A(DP_OP_102J5_124_3590_n504), .B(
        DP_OP_102J5_124_3590_n506), .CI(DP_OP_102J5_124_3590_n510), .CO(
        DP_OP_102J5_124_3590_n366), .S(DP_OP_102J5_124_3590_n367) );
  FADDX1_HVT DP_OP_102J5_124_3590_U270 ( .A(DP_OP_102J5_124_3590_n512), .B(
        DP_OP_102J5_124_3590_n508), .CI(DP_OP_102J5_124_3590_n514), .CO(
        DP_OP_102J5_124_3590_n364), .S(DP_OP_102J5_124_3590_n365) );
  FADDX1_HVT DP_OP_102J5_124_3590_U269 ( .A(DP_OP_102J5_124_3590_n379), .B(
        DP_OP_102J5_124_3590_n403), .CI(DP_OP_102J5_124_3590_n401), .CO(
        DP_OP_102J5_124_3590_n362), .S(DP_OP_102J5_124_3590_n363) );
  FADDX1_HVT DP_OP_102J5_124_3590_U268 ( .A(DP_OP_102J5_124_3590_n381), .B(
        DP_OP_102J5_124_3590_n397), .CI(DP_OP_102J5_124_3590_n389), .CO(
        DP_OP_102J5_124_3590_n360), .S(DP_OP_102J5_124_3590_n361) );
  FADDX1_HVT DP_OP_102J5_124_3590_U267 ( .A(DP_OP_102J5_124_3590_n391), .B(
        DP_OP_102J5_124_3590_n387), .CI(DP_OP_102J5_124_3590_n383), .CO(
        DP_OP_102J5_124_3590_n358), .S(DP_OP_102J5_124_3590_n359) );
  FADDX1_HVT DP_OP_102J5_124_3590_U266 ( .A(DP_OP_102J5_124_3590_n385), .B(
        DP_OP_102J5_124_3590_n399), .CI(DP_OP_102J5_124_3590_n395), .CO(
        DP_OP_102J5_124_3590_n356), .S(DP_OP_102J5_124_3590_n357) );
  FADDX1_HVT DP_OP_102J5_124_3590_U265 ( .A(DP_OP_102J5_124_3590_n393), .B(
        DP_OP_102J5_124_3590_n502), .CI(DP_OP_102J5_124_3590_n498), .CO(
        DP_OP_102J5_124_3590_n354), .S(DP_OP_102J5_124_3590_n355) );
  FADDX1_HVT DP_OP_102J5_124_3590_U264 ( .A(DP_OP_102J5_124_3590_n496), .B(
        DP_OP_102J5_124_3590_n500), .CI(DP_OP_102J5_124_3590_n494), .CO(
        DP_OP_102J5_124_3590_n352), .S(DP_OP_102J5_124_3590_n353) );
  FADDX1_HVT DP_OP_102J5_124_3590_U263 ( .A(DP_OP_102J5_124_3590_n490), .B(
        DP_OP_102J5_124_3590_n486), .CI(DP_OP_102J5_124_3590_n1423), .CO(
        DP_OP_102J5_124_3590_n350), .S(DP_OP_102J5_124_3590_n351) );
  FADDX1_HVT DP_OP_102J5_124_3590_U262 ( .A(DP_OP_102J5_124_3590_n492), .B(
        DP_OP_102J5_124_3590_n488), .CI(DP_OP_102J5_124_3590_n377), .CO(
        DP_OP_102J5_124_3590_n348), .S(DP_OP_102J5_124_3590_n349) );
  FADDX1_HVT DP_OP_102J5_124_3590_U261 ( .A(DP_OP_102J5_124_3590_n371), .B(
        DP_OP_102J5_124_3590_n375), .CI(DP_OP_102J5_124_3590_n369), .CO(
        DP_OP_102J5_124_3590_n346), .S(DP_OP_102J5_124_3590_n347) );
  FADDX1_HVT DP_OP_102J5_124_3590_U260 ( .A(DP_OP_102J5_124_3590_n484), .B(
        DP_OP_102J5_124_3590_n373), .CI(DP_OP_102J5_124_3590_n476), .CO(
        DP_OP_102J5_124_3590_n344), .S(DP_OP_102J5_124_3590_n345) );
  FADDX1_HVT DP_OP_102J5_124_3590_U259 ( .A(DP_OP_102J5_124_3590_n482), .B(
        DP_OP_102J5_124_3590_n478), .CI(DP_OP_102J5_124_3590_n480), .CO(
        DP_OP_102J5_124_3590_n342), .S(DP_OP_102J5_124_3590_n343) );
  FADDX1_HVT DP_OP_102J5_124_3590_U258 ( .A(DP_OP_102J5_124_3590_n367), .B(
        DP_OP_102J5_124_3590_n365), .CI(DP_OP_102J5_124_3590_n472), .CO(
        DP_OP_102J5_124_3590_n340), .S(DP_OP_102J5_124_3590_n341) );
  FADDX1_HVT DP_OP_102J5_124_3590_U257 ( .A(DP_OP_102J5_124_3590_n474), .B(
        DP_OP_102J5_124_3590_n359), .CI(DP_OP_102J5_124_3590_n361), .CO(
        DP_OP_102J5_124_3590_n338), .S(DP_OP_102J5_124_3590_n339) );
  FADDX1_HVT DP_OP_102J5_124_3590_U256 ( .A(DP_OP_102J5_124_3590_n357), .B(
        DP_OP_102J5_124_3590_n363), .CI(DP_OP_102J5_124_3590_n470), .CO(
        DP_OP_102J5_124_3590_n336), .S(DP_OP_102J5_124_3590_n337) );
  FADDX1_HVT DP_OP_102J5_124_3590_U255 ( .A(DP_OP_102J5_124_3590_n468), .B(
        DP_OP_102J5_124_3590_n466), .CI(DP_OP_102J5_124_3590_n355), .CO(
        DP_OP_102J5_124_3590_n334), .S(DP_OP_102J5_124_3590_n335) );
  FADDX1_HVT DP_OP_102J5_124_3590_U254 ( .A(DP_OP_102J5_124_3590_n464), .B(
        DP_OP_102J5_124_3590_n462), .CI(DP_OP_102J5_124_3590_n353), .CO(
        DP_OP_102J5_124_3590_n332), .S(DP_OP_102J5_124_3590_n333) );
  FADDX1_HVT DP_OP_102J5_124_3590_U253 ( .A(DP_OP_102J5_124_3590_n460), .B(
        DP_OP_102J5_124_3590_n458), .CI(DP_OP_102J5_124_3590_n456), .CO(
        DP_OP_102J5_124_3590_n330), .S(DP_OP_102J5_124_3590_n331) );
  FADDX1_HVT DP_OP_102J5_124_3590_U252 ( .A(DP_OP_102J5_124_3590_n351), .B(
        DP_OP_102J5_124_3590_n454), .CI(DP_OP_102J5_124_3590_n349), .CO(
        DP_OP_102J5_124_3590_n328), .S(DP_OP_102J5_124_3590_n329) );
  FADDX1_HVT DP_OP_102J5_124_3590_U251 ( .A(DP_OP_102J5_124_3590_n452), .B(
        DP_OP_102J5_124_3590_n345), .CI(DP_OP_102J5_124_3590_n347), .CO(
        DP_OP_102J5_124_3590_n326), .S(DP_OP_102J5_124_3590_n327) );
  FADDX1_HVT DP_OP_102J5_124_3590_U250 ( .A(DP_OP_102J5_124_3590_n450), .B(
        DP_OP_102J5_124_3590_n343), .CI(DP_OP_102J5_124_3590_n341), .CO(
        DP_OP_102J5_124_3590_n324), .S(DP_OP_102J5_124_3590_n325) );
  FADDX1_HVT DP_OP_102J5_124_3590_U249 ( .A(DP_OP_102J5_124_3590_n448), .B(
        DP_OP_102J5_124_3590_n339), .CI(DP_OP_102J5_124_3590_n446), .CO(
        DP_OP_102J5_124_3590_n322), .S(DP_OP_102J5_124_3590_n323) );
  FADDX1_HVT DP_OP_102J5_124_3590_U248 ( .A(DP_OP_102J5_124_3590_n337), .B(
        DP_OP_102J5_124_3590_n444), .CI(DP_OP_102J5_124_3590_n442), .CO(
        DP_OP_102J5_124_3590_n320), .S(DP_OP_102J5_124_3590_n321) );
  FADDX1_HVT DP_OP_102J5_124_3590_U247 ( .A(DP_OP_102J5_124_3590_n440), .B(
        DP_OP_102J5_124_3590_n335), .CI(DP_OP_102J5_124_3590_n333), .CO(
        DP_OP_102J5_124_3590_n318), .S(DP_OP_102J5_124_3590_n319) );
  FADDX1_HVT DP_OP_102J5_124_3590_U246 ( .A(DP_OP_102J5_124_3590_n438), .B(
        DP_OP_102J5_124_3590_n436), .CI(DP_OP_102J5_124_3590_n331), .CO(
        DP_OP_102J5_124_3590_n316), .S(DP_OP_102J5_124_3590_n317) );
  FADDX1_HVT DP_OP_102J5_124_3590_U245 ( .A(DP_OP_102J5_124_3590_n329), .B(
        DP_OP_102J5_124_3590_n434), .CI(DP_OP_102J5_124_3590_n432), .CO(
        DP_OP_102J5_124_3590_n314), .S(DP_OP_102J5_124_3590_n315) );
  FADDX1_HVT DP_OP_102J5_124_3590_U244 ( .A(DP_OP_102J5_124_3590_n327), .B(
        DP_OP_102J5_124_3590_n325), .CI(DP_OP_102J5_124_3590_n430), .CO(
        DP_OP_102J5_124_3590_n312), .S(DP_OP_102J5_124_3590_n313) );
  FADDX1_HVT DP_OP_102J5_124_3590_U243 ( .A(DP_OP_102J5_124_3590_n323), .B(
        DP_OP_102J5_124_3590_n428), .CI(DP_OP_102J5_124_3590_n321), .CO(
        DP_OP_102J5_124_3590_n310), .S(DP_OP_102J5_124_3590_n311) );
  FADDX1_HVT DP_OP_102J5_124_3590_U242 ( .A(DP_OP_102J5_124_3590_n426), .B(
        DP_OP_102J5_124_3590_n319), .CI(DP_OP_102J5_124_3590_n424), .CO(
        DP_OP_102J5_124_3590_n308), .S(DP_OP_102J5_124_3590_n309) );
  FADDX1_HVT DP_OP_102J5_124_3590_U241 ( .A(DP_OP_102J5_124_3590_n317), .B(
        DP_OP_102J5_124_3590_n422), .CI(DP_OP_102J5_124_3590_n315), .CO(
        DP_OP_102J5_124_3590_n306), .S(DP_OP_102J5_124_3590_n307) );
  FADDX1_HVT DP_OP_102J5_124_3590_U240 ( .A(DP_OP_102J5_124_3590_n420), .B(
        DP_OP_102J5_124_3590_n313), .CI(DP_OP_102J5_124_3590_n418), .CO(
        DP_OP_102J5_124_3590_n304), .S(DP_OP_102J5_124_3590_n305) );
  FADDX1_HVT DP_OP_102J5_124_3590_U239 ( .A(DP_OP_102J5_124_3590_n311), .B(
        DP_OP_102J5_124_3590_n416), .CI(DP_OP_102J5_124_3590_n309), .CO(
        DP_OP_102J5_124_3590_n302), .S(DP_OP_102J5_124_3590_n303) );
  FADDX1_HVT DP_OP_102J5_124_3590_U238 ( .A(DP_OP_102J5_124_3590_n414), .B(
        DP_OP_102J5_124_3590_n307), .CI(DP_OP_102J5_124_3590_n412), .CO(
        DP_OP_102J5_124_3590_n300), .S(DP_OP_102J5_124_3590_n301) );
  FADDX1_HVT DP_OP_102J5_124_3590_U237 ( .A(DP_OP_102J5_124_3590_n305), .B(
        DP_OP_102J5_124_3590_n303), .CI(DP_OP_102J5_124_3590_n410), .CO(
        DP_OP_102J5_124_3590_n298), .S(DP_OP_102J5_124_3590_n299) );
  FADDX1_HVT DP_OP_102J5_124_3590_U236 ( .A(DP_OP_102J5_124_3590_n408), .B(
        DP_OP_102J5_124_3590_n301), .CI(DP_OP_102J5_124_3590_n299), .CO(
        DP_OP_102J5_124_3590_n296), .S(DP_OP_102J5_124_3590_n297) );
  FADDX1_HVT DP_OP_102J5_124_3590_U235 ( .A(DP_OP_102J5_124_3590_n404), .B(
        DP_OP_102J5_124_3590_n2292), .CI(DP_OP_102J5_124_3590_n2248), .CO(
        DP_OP_102J5_124_3590_n221), .S(DP_OP_102J5_124_3590_n295) );
  FADDX1_HVT DP_OP_102J5_124_3590_U234 ( .A(DP_OP_102J5_124_3590_n1896), .B(
        DP_OP_102J5_124_3590_n2204), .CI(DP_OP_102J5_124_3590_n1457), .CO(
        DP_OP_102J5_124_3590_n293), .S(DP_OP_102J5_124_3590_n294) );
  FADDX1_HVT DP_OP_102J5_124_3590_U233 ( .A(DP_OP_102J5_124_3590_n1808), .B(
        DP_OP_102J5_124_3590_n2160), .CI(DP_OP_102J5_124_3590_n1501), .CO(
        DP_OP_102J5_124_3590_n291), .S(DP_OP_102J5_124_3590_n292) );
  FADDX1_HVT DP_OP_102J5_124_3590_U232 ( .A(DP_OP_102J5_124_3590_n1721), .B(
        DP_OP_102J5_124_3590_n2116), .CI(DP_OP_102J5_124_3590_n2072), .CO(
        DP_OP_102J5_124_3590_n289), .S(DP_OP_102J5_124_3590_n290) );
  FADDX1_HVT DP_OP_102J5_124_3590_U231 ( .A(DP_OP_102J5_124_3590_n2028), .B(
        DP_OP_102J5_124_3590_n1984), .CI(DP_OP_102J5_124_3590_n1940), .CO(
        DP_OP_102J5_124_3590_n287), .S(DP_OP_102J5_124_3590_n288) );
  FADDX1_HVT DP_OP_102J5_124_3590_U230 ( .A(DP_OP_102J5_124_3590_n1633), .B(
        DP_OP_102J5_124_3590_n1545), .CI(DP_OP_102J5_124_3590_n1589), .CO(
        DP_OP_102J5_124_3590_n285), .S(DP_OP_102J5_124_3590_n286) );
  FADDX1_HVT DP_OP_102J5_124_3590_U229 ( .A(DP_OP_102J5_124_3590_n1765), .B(
        DP_OP_102J5_124_3590_n1852), .CI(DP_OP_102J5_124_3590_n1677), .CO(
        DP_OP_102J5_124_3590_n283), .S(DP_OP_102J5_124_3590_n284) );
  FADDX1_HVT DP_OP_102J5_124_3590_U228 ( .A(DP_OP_102J5_124_3590_n390), .B(
        DP_OP_102J5_124_3590_n380), .CI(DP_OP_102J5_124_3590_n378), .CO(
        DP_OP_102J5_124_3590_n281), .S(DP_OP_102J5_124_3590_n282) );
  FADDX1_HVT DP_OP_102J5_124_3590_U227 ( .A(DP_OP_102J5_124_3590_n394), .B(
        DP_OP_102J5_124_3590_n382), .CI(DP_OP_102J5_124_3590_n386), .CO(
        DP_OP_102J5_124_3590_n279), .S(DP_OP_102J5_124_3590_n280) );
  FADDX1_HVT DP_OP_102J5_124_3590_U226 ( .A(DP_OP_102J5_124_3590_n396), .B(
        DP_OP_102J5_124_3590_n384), .CI(DP_OP_102J5_124_3590_n388), .CO(
        DP_OP_102J5_124_3590_n277), .S(DP_OP_102J5_124_3590_n278) );
  FADDX1_HVT DP_OP_102J5_124_3590_U225 ( .A(DP_OP_102J5_124_3590_n392), .B(
        DP_OP_102J5_124_3590_n398), .CI(DP_OP_102J5_124_3590_n400), .CO(
        DP_OP_102J5_124_3590_n275), .S(DP_OP_102J5_124_3590_n276) );
  FADDX1_HVT DP_OP_102J5_124_3590_U224 ( .A(DP_OP_102J5_124_3590_n402), .B(
        DP_OP_102J5_124_3590_n295), .CI(DP_OP_102J5_124_3590_n290), .CO(
        DP_OP_102J5_124_3590_n273), .S(DP_OP_102J5_124_3590_n274) );
  FADDX1_HVT DP_OP_102J5_124_3590_U223 ( .A(DP_OP_102J5_124_3590_n292), .B(
        DP_OP_102J5_124_3590_n284), .CI(DP_OP_102J5_124_3590_n286), .CO(
        DP_OP_102J5_124_3590_n271), .S(DP_OP_102J5_124_3590_n272) );
  FADDX1_HVT DP_OP_102J5_124_3590_U222 ( .A(DP_OP_102J5_124_3590_n288), .B(
        DP_OP_102J5_124_3590_n294), .CI(DP_OP_102J5_124_3590_n376), .CO(
        DP_OP_102J5_124_3590_n269), .S(DP_OP_102J5_124_3590_n270) );
  FADDX1_HVT DP_OP_102J5_124_3590_U221 ( .A(DP_OP_102J5_124_3590_n368), .B(
        DP_OP_102J5_124_3590_n370), .CI(DP_OP_102J5_124_3590_n372), .CO(
        DP_OP_102J5_124_3590_n267), .S(DP_OP_102J5_124_3590_n268) );
  FADDX1_HVT DP_OP_102J5_124_3590_U220 ( .A(DP_OP_102J5_124_3590_n374), .B(
        DP_OP_102J5_124_3590_n366), .CI(DP_OP_102J5_124_3590_n364), .CO(
        DP_OP_102J5_124_3590_n265), .S(DP_OP_102J5_124_3590_n266) );
  FADDX1_HVT DP_OP_102J5_124_3590_U219 ( .A(DP_OP_102J5_124_3590_n1422), .B(
        DP_OP_102J5_124_3590_n362), .CI(DP_OP_102J5_124_3590_n360), .CO(
        DP_OP_102J5_124_3590_n263), .S(DP_OP_102J5_124_3590_n264) );
  FADDX1_HVT DP_OP_102J5_124_3590_U218 ( .A(DP_OP_102J5_124_3590_n358), .B(
        DP_OP_102J5_124_3590_n278), .CI(DP_OP_102J5_124_3590_n276), .CO(
        DP_OP_102J5_124_3590_n261), .S(DP_OP_102J5_124_3590_n262) );
  FADDX1_HVT DP_OP_102J5_124_3590_U217 ( .A(DP_OP_102J5_124_3590_n356), .B(
        DP_OP_102J5_124_3590_n280), .CI(DP_OP_102J5_124_3590_n282), .CO(
        DP_OP_102J5_124_3590_n259), .S(DP_OP_102J5_124_3590_n260) );
  FADDX1_HVT DP_OP_102J5_124_3590_U216 ( .A(DP_OP_102J5_124_3590_n354), .B(
        DP_OP_102J5_124_3590_n274), .CI(DP_OP_102J5_124_3590_n272), .CO(
        DP_OP_102J5_124_3590_n257), .S(DP_OP_102J5_124_3590_n258) );
  FADDX1_HVT DP_OP_102J5_124_3590_U215 ( .A(DP_OP_102J5_124_3590_n352), .B(
        DP_OP_102J5_124_3590_n350), .CI(DP_OP_102J5_124_3590_n348), .CO(
        DP_OP_102J5_124_3590_n255), .S(DP_OP_102J5_124_3590_n256) );
  FADDX1_HVT DP_OP_102J5_124_3590_U214 ( .A(DP_OP_102J5_124_3590_n270), .B(
        DP_OP_102J5_124_3590_n346), .CI(DP_OP_102J5_124_3590_n344), .CO(
        DP_OP_102J5_124_3590_n253), .S(DP_OP_102J5_124_3590_n254) );
  FADDX1_HVT DP_OP_102J5_124_3590_U213 ( .A(DP_OP_102J5_124_3590_n342), .B(
        DP_OP_102J5_124_3590_n268), .CI(DP_OP_102J5_124_3590_n266), .CO(
        DP_OP_102J5_124_3590_n251), .S(DP_OP_102J5_124_3590_n252) );
  FADDX1_HVT DP_OP_102J5_124_3590_U212 ( .A(DP_OP_102J5_124_3590_n340), .B(
        DP_OP_102J5_124_3590_n338), .CI(DP_OP_102J5_124_3590_n264), .CO(
        DP_OP_102J5_124_3590_n249), .S(DP_OP_102J5_124_3590_n250) );
  FADDX1_HVT DP_OP_102J5_124_3590_U211 ( .A(DP_OP_102J5_124_3590_n262), .B(
        DP_OP_102J5_124_3590_n260), .CI(DP_OP_102J5_124_3590_n336), .CO(
        DP_OP_102J5_124_3590_n247), .S(DP_OP_102J5_124_3590_n248) );
  FADDX1_HVT DP_OP_102J5_124_3590_U210 ( .A(DP_OP_102J5_124_3590_n334), .B(
        DP_OP_102J5_124_3590_n258), .CI(DP_OP_102J5_124_3590_n332), .CO(
        DP_OP_102J5_124_3590_n245), .S(DP_OP_102J5_124_3590_n246) );
  FADDX1_HVT DP_OP_102J5_124_3590_U209 ( .A(DP_OP_102J5_124_3590_n330), .B(
        DP_OP_102J5_124_3590_n256), .CI(DP_OP_102J5_124_3590_n328), .CO(
        DP_OP_102J5_124_3590_n243), .S(DP_OP_102J5_124_3590_n244) );
  FADDX1_HVT DP_OP_102J5_124_3590_U208 ( .A(DP_OP_102J5_124_3590_n254), .B(
        DP_OP_102J5_124_3590_n324), .CI(DP_OP_102J5_124_3590_n252), .CO(
        DP_OP_102J5_124_3590_n241), .S(DP_OP_102J5_124_3590_n242) );
  FADDX1_HVT DP_OP_102J5_124_3590_U207 ( .A(DP_OP_102J5_124_3590_n326), .B(
        DP_OP_102J5_124_3590_n322), .CI(DP_OP_102J5_124_3590_n250), .CO(
        DP_OP_102J5_124_3590_n239), .S(DP_OP_102J5_124_3590_n240) );
  FADDX1_HVT DP_OP_102J5_124_3590_U206 ( .A(DP_OP_102J5_124_3590_n248), .B(
        DP_OP_102J5_124_3590_n320), .CI(DP_OP_102J5_124_3590_n318), .CO(
        DP_OP_102J5_124_3590_n237), .S(DP_OP_102J5_124_3590_n238) );
  FADDX1_HVT DP_OP_102J5_124_3590_U205 ( .A(DP_OP_102J5_124_3590_n246), .B(
        DP_OP_102J5_124_3590_n316), .CI(DP_OP_102J5_124_3590_n244), .CO(
        DP_OP_102J5_124_3590_n235), .S(DP_OP_102J5_124_3590_n236) );
  FADDX1_HVT DP_OP_102J5_124_3590_U204 ( .A(DP_OP_102J5_124_3590_n314), .B(
        DP_OP_102J5_124_3590_n242), .CI(DP_OP_102J5_124_3590_n312), .CO(
        DP_OP_102J5_124_3590_n233), .S(DP_OP_102J5_124_3590_n234) );
  FADDX1_HVT DP_OP_102J5_124_3590_U203 ( .A(DP_OP_102J5_124_3590_n240), .B(
        DP_OP_102J5_124_3590_n310), .CI(DP_OP_102J5_124_3590_n238), .CO(
        DP_OP_102J5_124_3590_n231), .S(DP_OP_102J5_124_3590_n232) );
  FADDX1_HVT DP_OP_102J5_124_3590_U202 ( .A(DP_OP_102J5_124_3590_n308), .B(
        DP_OP_102J5_124_3590_n236), .CI(DP_OP_102J5_124_3590_n306), .CO(
        DP_OP_102J5_124_3590_n229), .S(DP_OP_102J5_124_3590_n230) );
  FADDX1_HVT DP_OP_102J5_124_3590_U201 ( .A(DP_OP_102J5_124_3590_n234), .B(
        DP_OP_102J5_124_3590_n304), .CI(DP_OP_102J5_124_3590_n232), .CO(
        DP_OP_102J5_124_3590_n227), .S(DP_OP_102J5_124_3590_n228) );
  FADDX1_HVT DP_OP_102J5_124_3590_U200 ( .A(DP_OP_102J5_124_3590_n302), .B(
        DP_OP_102J5_124_3590_n230), .CI(DP_OP_102J5_124_3590_n300), .CO(
        DP_OP_102J5_124_3590_n225), .S(DP_OP_102J5_124_3590_n226) );
  FADDX1_HVT DP_OP_102J5_124_3590_U199 ( .A(DP_OP_102J5_124_3590_n228), .B(
        DP_OP_102J5_124_3590_n298), .CI(DP_OP_102J5_124_3590_n226), .CO(
        DP_OP_102J5_124_3590_n223), .S(DP_OP_102J5_124_3590_n224) );
  FADDX1_HVT DP_OP_102J5_124_3590_U197 ( .A(DP_OP_102J5_124_3590_n287), .B(
        DP_OP_102J5_124_3590_n283), .CI(DP_OP_102J5_124_3590_n222), .CO(
        DP_OP_102J5_124_3590_n219), .S(DP_OP_102J5_124_3590_n220) );
  FADDX1_HVT DP_OP_102J5_124_3590_U196 ( .A(DP_OP_102J5_124_3590_n289), .B(
        DP_OP_102J5_124_3590_n291), .CI(DP_OP_102J5_124_3590_n285), .CO(
        DP_OP_102J5_124_3590_n217), .S(DP_OP_102J5_124_3590_n218) );
  FADDX1_HVT DP_OP_102J5_124_3590_U195 ( .A(DP_OP_102J5_124_3590_n293), .B(
        DP_OP_102J5_124_3590_n277), .CI(DP_OP_102J5_124_3590_n275), .CO(
        DP_OP_102J5_124_3590_n215), .S(DP_OP_102J5_124_3590_n216) );
  FADDX1_HVT DP_OP_102J5_124_3590_U194 ( .A(DP_OP_102J5_124_3590_n281), .B(
        DP_OP_102J5_124_3590_n279), .CI(DP_OP_102J5_124_3590_n1421), .CO(
        DP_OP_102J5_124_3590_n213), .S(DP_OP_102J5_124_3590_n214) );
  FADDX1_HVT DP_OP_102J5_124_3590_U193 ( .A(DP_OP_102J5_124_3590_n273), .B(
        DP_OP_102J5_124_3590_n271), .CI(DP_OP_102J5_124_3590_n218), .CO(
        DP_OP_102J5_124_3590_n211), .S(DP_OP_102J5_124_3590_n212) );
  FADDX1_HVT DP_OP_102J5_124_3590_U192 ( .A(DP_OP_102J5_124_3590_n220), .B(
        DP_OP_102J5_124_3590_n269), .CI(DP_OP_102J5_124_3590_n267), .CO(
        DP_OP_102J5_124_3590_n209), .S(DP_OP_102J5_124_3590_n210) );
  FADDX1_HVT DP_OP_102J5_124_3590_U191 ( .A(DP_OP_102J5_124_3590_n265), .B(
        DP_OP_102J5_124_3590_n263), .CI(DP_OP_102J5_124_3590_n216), .CO(
        DP_OP_102J5_124_3590_n207), .S(DP_OP_102J5_124_3590_n208) );
  FADDX1_HVT DP_OP_102J5_124_3590_U190 ( .A(DP_OP_102J5_124_3590_n261), .B(
        DP_OP_102J5_124_3590_n259), .CI(DP_OP_102J5_124_3590_n214), .CO(
        DP_OP_102J5_124_3590_n205), .S(DP_OP_102J5_124_3590_n206) );
  FADDX1_HVT DP_OP_102J5_124_3590_U189 ( .A(DP_OP_102J5_124_3590_n257), .B(
        DP_OP_102J5_124_3590_n212), .CI(DP_OP_102J5_124_3590_n255), .CO(
        DP_OP_102J5_124_3590_n203), .S(DP_OP_102J5_124_3590_n204) );
  FADDX1_HVT DP_OP_102J5_124_3590_U188 ( .A(DP_OP_102J5_124_3590_n210), .B(
        DP_OP_102J5_124_3590_n253), .CI(DP_OP_102J5_124_3590_n251), .CO(
        DP_OP_102J5_124_3590_n201), .S(DP_OP_102J5_124_3590_n202) );
  FADDX1_HVT DP_OP_102J5_124_3590_U187 ( .A(DP_OP_102J5_124_3590_n249), .B(
        DP_OP_102J5_124_3590_n208), .CI(DP_OP_102J5_124_3590_n247), .CO(
        DP_OP_102J5_124_3590_n199), .S(DP_OP_102J5_124_3590_n200) );
  FADDX1_HVT DP_OP_102J5_124_3590_U186 ( .A(DP_OP_102J5_124_3590_n206), .B(
        DP_OP_102J5_124_3590_n245), .CI(DP_OP_102J5_124_3590_n204), .CO(
        DP_OP_102J5_124_3590_n197), .S(DP_OP_102J5_124_3590_n198) );
  FADDX1_HVT DP_OP_102J5_124_3590_U185 ( .A(DP_OP_102J5_124_3590_n243), .B(
        DP_OP_102J5_124_3590_n202), .CI(DP_OP_102J5_124_3590_n241), .CO(
        DP_OP_102J5_124_3590_n195), .S(DP_OP_102J5_124_3590_n196) );
  FADDX1_HVT DP_OP_102J5_124_3590_U184 ( .A(DP_OP_102J5_124_3590_n239), .B(
        DP_OP_102J5_124_3590_n200), .CI(DP_OP_102J5_124_3590_n237), .CO(
        DP_OP_102J5_124_3590_n193), .S(DP_OP_102J5_124_3590_n194) );
  FADDX1_HVT DP_OP_102J5_124_3590_U183 ( .A(DP_OP_102J5_124_3590_n198), .B(
        DP_OP_102J5_124_3590_n235), .CI(DP_OP_102J5_124_3590_n196), .CO(
        DP_OP_102J5_124_3590_n191), .S(DP_OP_102J5_124_3590_n192) );
  FADDX1_HVT DP_OP_102J5_124_3590_U182 ( .A(DP_OP_102J5_124_3590_n233), .B(
        DP_OP_102J5_124_3590_n231), .CI(DP_OP_102J5_124_3590_n194), .CO(
        DP_OP_102J5_124_3590_n189), .S(DP_OP_102J5_124_3590_n190) );
  FADDX1_HVT DP_OP_102J5_124_3590_U181 ( .A(DP_OP_102J5_124_3590_n229), .B(
        DP_OP_102J5_124_3590_n192), .CI(DP_OP_102J5_124_3590_n227), .CO(
        DP_OP_102J5_124_3590_n187), .S(DP_OP_102J5_124_3590_n188) );
  FADDX1_HVT DP_OP_102J5_124_3590_U180 ( .A(DP_OP_102J5_124_3590_n190), .B(
        DP_OP_102J5_124_3590_n225), .CI(DP_OP_102J5_124_3590_n188), .CO(
        DP_OP_102J5_124_3590_n185), .S(DP_OP_102J5_124_3590_n186) );
  FADDX1_HVT DP_OP_102J5_124_3590_U179 ( .A(DP_OP_102J5_124_3590_n221), .B(
        DP_OP_102J5_124_3590_n219), .CI(DP_OP_102J5_124_3590_n217), .CO(
        DP_OP_102J5_124_3590_n183), .S(DP_OP_102J5_124_3590_n184) );
  FADDX1_HVT DP_OP_102J5_124_3590_U178 ( .A(DP_OP_102J5_124_3590_n1420), .B(
        DP_OP_102J5_124_3590_n215), .CI(DP_OP_102J5_124_3590_n213), .CO(
        DP_OP_102J5_124_3590_n181), .S(DP_OP_102J5_124_3590_n182) );
  FADDX1_HVT DP_OP_102J5_124_3590_U177 ( .A(DP_OP_102J5_124_3590_n211), .B(
        DP_OP_102J5_124_3590_n184), .CI(DP_OP_102J5_124_3590_n209), .CO(
        DP_OP_102J5_124_3590_n179), .S(DP_OP_102J5_124_3590_n180) );
  FADDX1_HVT DP_OP_102J5_124_3590_U176 ( .A(DP_OP_102J5_124_3590_n207), .B(
        DP_OP_102J5_124_3590_n182), .CI(DP_OP_102J5_124_3590_n205), .CO(
        DP_OP_102J5_124_3590_n177), .S(DP_OP_102J5_124_3590_n178) );
  FADDX1_HVT DP_OP_102J5_124_3590_U175 ( .A(DP_OP_102J5_124_3590_n203), .B(
        DP_OP_102J5_124_3590_n180), .CI(DP_OP_102J5_124_3590_n201), .CO(
        DP_OP_102J5_124_3590_n175), .S(DP_OP_102J5_124_3590_n176) );
  FADDX1_HVT DP_OP_102J5_124_3590_U174 ( .A(DP_OP_102J5_124_3590_n199), .B(
        DP_OP_102J5_124_3590_n178), .CI(DP_OP_102J5_124_3590_n197), .CO(
        DP_OP_102J5_124_3590_n173), .S(DP_OP_102J5_124_3590_n174) );
  FADDX1_HVT DP_OP_102J5_124_3590_U173 ( .A(DP_OP_102J5_124_3590_n176), .B(
        DP_OP_102J5_124_3590_n195), .CI(DP_OP_102J5_124_3590_n193), .CO(
        DP_OP_102J5_124_3590_n171), .S(DP_OP_102J5_124_3590_n172) );
  FADDX1_HVT DP_OP_102J5_124_3590_U172 ( .A(DP_OP_102J5_124_3590_n174), .B(
        DP_OP_102J5_124_3590_n191), .CI(DP_OP_102J5_124_3590_n172), .CO(
        DP_OP_102J5_124_3590_n169), .S(DP_OP_102J5_124_3590_n170) );
  FADDX1_HVT DP_OP_102J5_124_3590_U171 ( .A(DP_OP_102J5_124_3590_n189), .B(
        DP_OP_102J5_124_3590_n187), .CI(DP_OP_102J5_124_3590_n170), .CO(
        DP_OP_102J5_124_3590_n167), .S(DP_OP_102J5_124_3590_n168) );
  FADDX1_HVT DP_OP_102J5_124_3590_U169 ( .A(DP_OP_102J5_124_3590_n166), .B(
        DP_OP_102J5_124_3590_n183), .CI(DP_OP_102J5_124_3590_n181), .CO(
        DP_OP_102J5_124_3590_n163), .S(DP_OP_102J5_124_3590_n164) );
  FADDX1_HVT DP_OP_102J5_124_3590_U168 ( .A(DP_OP_102J5_124_3590_n179), .B(
        DP_OP_102J5_124_3590_n164), .CI(DP_OP_102J5_124_3590_n177), .CO(
        DP_OP_102J5_124_3590_n161), .S(DP_OP_102J5_124_3590_n162) );
  FADDX1_HVT DP_OP_102J5_124_3590_U167 ( .A(DP_OP_102J5_124_3590_n175), .B(
        DP_OP_102J5_124_3590_n162), .CI(DP_OP_102J5_124_3590_n173), .CO(
        DP_OP_102J5_124_3590_n159), .S(DP_OP_102J5_124_3590_n160) );
  FADDX1_HVT DP_OP_102J5_124_3590_U166 ( .A(DP_OP_102J5_124_3590_n171), .B(
        DP_OP_102J5_124_3590_n160), .CI(DP_OP_102J5_124_3590_n169), .CO(
        DP_OP_102J5_124_3590_n157), .S(DP_OP_102J5_124_3590_n158) );
  FADDX1_HVT DP_OP_102J5_124_3590_U164 ( .A(DP_OP_102J5_124_3590_n165), .B(
        DP_OP_102J5_124_3590_n156), .CI(DP_OP_102J5_124_3590_n163), .CO(
        DP_OP_102J5_124_3590_n153), .S(DP_OP_102J5_124_3590_n154) );
  FADDX1_HVT DP_OP_102J5_124_3590_U163 ( .A(DP_OP_102J5_124_3590_n154), .B(
        DP_OP_102J5_124_3590_n161), .CI(DP_OP_102J5_124_3590_n159), .CO(
        DP_OP_102J5_124_3590_n151), .S(DP_OP_102J5_124_3590_n152) );
  FADDX1_HVT DP_OP_102J5_124_3590_U162 ( .A(DP_OP_102J5_124_3590_n1419), .B(
        DP_OP_102J5_124_3590_n155), .CI(DP_OP_102J5_124_3590_n153), .CO(
        DP_OP_102J5_124_3590_n149), .S(DP_OP_102J5_124_3590_n150) );
  FADDX1_HVT DP_OP_102J5_124_3590_U154 ( .A(DP_OP_102J5_124_3590_n1405), .B(
        DP_OP_102J5_124_3590_n1403), .CI(DP_OP_102J5_124_3590_n1401), .CO(
        DP_OP_102J5_124_3590_n116), .S(n_accumulator_sum[0]) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U153 ( .A1(DP_OP_102J5_124_3590_n1353), 
        .A2(DP_OP_102J5_124_3590_n1355), .Y(DP_OP_102J5_124_3590_n115) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U152 ( .A1(DP_OP_102J5_124_3590_n1355), .A2(
        DP_OP_102J5_124_3590_n1353), .Y(DP_OP_102J5_124_3590_n114) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U146 ( .A1(DP_OP_102J5_124_3590_n1269), 
        .A2(DP_OP_102J5_124_3590_n1271), .Y(DP_OP_102J5_124_3590_n112) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U137 ( .A1(DP_OP_102J5_124_3590_n1147), 
        .A2(DP_OP_102J5_124_3590_n1149), .Y(DP_OP_102J5_124_3590_n106) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U129 ( .A1(DP_OP_102J5_124_3590_n1007), 
        .A2(DP_OP_102J5_124_3590_n1009), .Y(DP_OP_102J5_124_3590_n101) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U128 ( .A1(DP_OP_102J5_124_3590_n1009), .A2(
        DP_OP_102J5_124_3590_n1007), .Y(DP_OP_102J5_124_3590_n100) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U123 ( .A1(DP_OP_102J5_124_3590_n857), .A2(
        DP_OP_102J5_124_3590_n859), .Y(DP_OP_102J5_124_3590_n98) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U115 ( .A1(DP_OP_102J5_124_3590_n703), .A2(
        DP_OP_102J5_124_3590_n705), .Y(DP_OP_102J5_124_3590_n93) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U114 ( .A1(DP_OP_102J5_124_3590_n705), .A2(
        DP_OP_102J5_124_3590_n703), .Y(DP_OP_102J5_124_3590_n92) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U108 ( .A1(DP_OP_102J5_124_3590_n545), .A2(
        DP_OP_102J5_124_3590_n702), .Y(DP_OP_102J5_124_3590_n89) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U107 ( .A1(DP_OP_102J5_124_3590_n702), .A2(
        DP_OP_102J5_124_3590_n545), .Y(DP_OP_102J5_124_3590_n88) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U102 ( .A1(DP_OP_102J5_124_3590_n407), .A2(
        DP_OP_102J5_124_3590_n544), .Y(DP_OP_102J5_124_3590_n86) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U101 ( .A1(DP_OP_102J5_124_3590_n544), .A2(
        DP_OP_102J5_124_3590_n407), .Y(DP_OP_102J5_124_3590_n85) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U93 ( .A1(DP_OP_102J5_124_3590_n297), .A2(
        DP_OP_102J5_124_3590_n406), .Y(DP_OP_102J5_124_3590_n80) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U92 ( .A1(DP_OP_102J5_124_3590_n406), .A2(
        DP_OP_102J5_124_3590_n297), .Y(DP_OP_102J5_124_3590_n79) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U85 ( .A1(DP_OP_102J5_124_3590_n224), .A2(
        DP_OP_102J5_124_3590_n296), .Y(DP_OP_102J5_124_3590_n75) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U84 ( .A1(DP_OP_102J5_124_3590_n296), .A2(
        DP_OP_102J5_124_3590_n224), .Y(DP_OP_102J5_124_3590_n74) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U80 ( .A1(DP_OP_102J5_124_3590_n79), .A2(
        DP_OP_102J5_124_3590_n74), .Y(DP_OP_102J5_124_3590_n72) );
  AOI21X1_HVT DP_OP_102J5_124_3590_U79 ( .A1(DP_OP_102J5_124_3590_n81), .A2(
        DP_OP_102J5_124_3590_n72), .A3(DP_OP_102J5_124_3590_n73), .Y(
        DP_OP_102J5_124_3590_n71) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U77 ( .A1(DP_OP_102J5_124_3590_n186), .A2(
        DP_OP_102J5_124_3590_n223), .Y(DP_OP_102J5_124_3590_n70) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U76 ( .A1(DP_OP_102J5_124_3590_n223), .A2(
        DP_OP_102J5_124_3590_n186), .Y(DP_OP_102J5_124_3590_n69) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U71 ( .A1(DP_OP_102J5_124_3590_n168), .A2(
        DP_OP_102J5_124_3590_n185), .Y(DP_OP_102J5_124_3590_n67) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U70 ( .A1(DP_OP_102J5_124_3590_n185), .A2(
        DP_OP_102J5_124_3590_n168), .Y(DP_OP_102J5_124_3590_n66) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U60 ( .A1(DP_OP_102J5_124_3590_n167), .A2(
        DP_OP_102J5_124_3590_n158), .Y(DP_OP_102J5_124_3590_n59) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U59 ( .A1(DP_OP_102J5_124_3590_n158), .A2(
        DP_OP_102J5_124_3590_n167), .Y(DP_OP_102J5_124_3590_n58) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U54 ( .A1(DP_OP_102J5_124_3590_n157), .A2(
        DP_OP_102J5_124_3590_n152), .Y(DP_OP_102J5_124_3590_n56) );
  AOI21X1_HVT DP_OP_102J5_124_3590_U48 ( .A1(DP_OP_102J5_124_3590_n57), .A2(
        n250), .A3(DP_OP_102J5_124_3590_n54), .Y(DP_OP_102J5_124_3590_n52) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U46 ( .A1(DP_OP_102J5_124_3590_n151), .A2(
        DP_OP_102J5_124_3590_n150), .Y(DP_OP_102J5_124_3590_n51) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U45 ( .A1(DP_OP_102J5_124_3590_n150), .A2(
        DP_OP_102J5_124_3590_n151), .Y(DP_OP_102J5_124_3590_n50) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U40 ( .A1(DP_OP_102J5_124_3590_n149), .A2(
        DP_OP_102J5_124_3590_n148), .Y(DP_OP_102J5_124_3590_n48) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U39 ( .A1(DP_OP_102J5_124_3590_n148), .A2(
        DP_OP_102J5_124_3590_n149), .Y(DP_OP_102J5_124_3590_n47) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U35 ( .A1(DP_OP_102J5_124_3590_n47), .A2(
        DP_OP_102J5_124_3590_n50), .Y(DP_OP_102J5_124_3590_n45) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U33 ( .A1(n250), .A2(
        DP_OP_102J5_124_3590_n45), .Y(DP_OP_102J5_124_3590_n43) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U31 ( .A1(DP_OP_102J5_124_3590_n43), .A2(
        DP_OP_102J5_124_3590_n58), .Y(DP_OP_102J5_124_3590_n41) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U26 ( .A1(DP_OP_102J5_124_3590_n146), .A2(
        DP_OP_102J5_124_3590_n147), .Y(DP_OP_102J5_124_3590_n37) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U19 ( .A1(DP_OP_102J5_124_3590_n41), .A2(
        n259), .Y(DP_OP_102J5_124_3590_n32) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U16 ( .A1(DP_OP_102J5_124_3590_n144), .A2(
        DP_OP_102J5_124_3590_n145), .Y(DP_OP_102J5_124_3590_n30) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U15 ( .A1(DP_OP_102J5_124_3590_n145), .A2(
        DP_OP_102J5_124_3590_n144), .Y(DP_OP_102J5_124_3590_n29) );
  FADDX1_HVT DP_OP_102J5_124_3590_U7 ( .A(DP_OP_102J5_124_3590_n143), .B(
        DP_OP_102J5_124_3590_n142), .CI(n249), .CO(DP_OP_102J5_124_3590_n25), 
        .S(n_accumulator_sum[19]) );
  FADDX1_HVT DP_OP_102J5_124_3590_U6 ( .A(DP_OP_102J5_124_3590_n141), .B(
        DP_OP_102J5_124_3590_n140), .CI(DP_OP_102J5_124_3590_n25), .CO(
        DP_OP_102J5_124_3590_n24), .S(n_accumulator_sum[20]) );
  FADDX1_HVT DP_OP_102J5_124_3590_U5 ( .A(DP_OP_102J5_124_3590_n139), .B(
        DP_OP_102J5_124_3590_n138), .CI(DP_OP_102J5_124_3590_n24), .CO(
        DP_OP_102J5_124_3590_n23), .S(n_accumulator_sum[21]) );
  XNOR2X1_HVT DP_OP_102J5_124_3590_U590 ( .A1(DP_OP_102J5_124_3590_n1901), 
        .A2(DP_OP_102J5_124_3590_n2033), .Y(DP_OP_102J5_124_3590_n1005) );
  OAI21X1_HVT DP_OP_102J5_124_3590_U148 ( .A1(DP_OP_102J5_124_3590_n4), .A2(
        DP_OP_102J5_124_3590_n114), .A3(DP_OP_102J5_124_3590_n115), .Y(
        DP_OP_102J5_124_3590_n113) );
  OAI21X1_HVT DP_OP_102J5_124_3590_U125 ( .A1(DP_OP_102J5_124_3590_n102), .A2(
        DP_OP_102J5_124_3590_n100), .A3(DP_OP_102J5_124_3590_n101), .Y(
        DP_OP_102J5_124_3590_n99) );
  OAI21X1_HVT DP_OP_102J5_124_3590_U111 ( .A1(DP_OP_102J5_124_3590_n94), .A2(
        DP_OP_102J5_124_3590_n92), .A3(DP_OP_102J5_124_3590_n93), .Y(
        DP_OP_102J5_124_3590_n91) );
  OAI21X1_HVT DP_OP_102J5_124_3590_U12 ( .A1(DP_OP_102J5_124_3590_n29), .A2(
        DP_OP_102J5_124_3590_n33), .A3(DP_OP_102J5_124_3590_n30), .Y(
        DP_OP_102J5_124_3590_n28) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U1178 ( .A1(n211), .A2(
        DP_OP_102J5_124_3590_n1797), .Y(DP_OP_102J5_124_3590_n1789) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U814 ( .A1(n264), .A2(
        DP_OP_102J5_124_3590_n2), .Y(DP_OP_102J5_124_3590_n1426) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U815 ( .A1(n265), .A2(
        DP_OP_102J5_124_3590_n2), .Y(DP_OP_102J5_124_3590_n1427) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U811 ( .A1(n266), .A2(
        DP_OP_102J5_124_3590_n2), .Y(DP_OP_102J5_124_3590_n1423) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U808 ( .A1(n163), .A2(accumulate_reset), .Y(
        DP_OP_102J5_124_3590_n1420) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U820 ( .A1(n254), .A2(
        DP_OP_102J5_124_3590_n2), .Y(DP_OP_102J5_124_3590_n1432) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U801 ( .A1(n269), .A2(accumulate_reset), .Y(
        DP_OP_102J5_124_3590_n141) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U818 ( .A1(n252), .A2(
        DP_OP_102J5_124_3590_n2), .Y(DP_OP_102J5_124_3590_n1430) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U817 ( .A1(n251), .A2(
        DP_OP_102J5_124_3590_n2), .Y(DP_OP_102J5_124_3590_n1429) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U813 ( .A1(n267), .A2(
        DP_OP_102J5_124_3590_n2), .Y(DP_OP_102J5_124_3590_n1425) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U819 ( .A1(n253), .A2(
        DP_OP_102J5_124_3590_n2), .Y(DP_OP_102J5_124_3590_n1431) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U807 ( .A1(n268), .A2(accumulate_reset), .Y(
        DP_OP_102J5_124_3590_n165) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U806 ( .A1(n258), .A2(accumulate_reset), .Y(
        DP_OP_102J5_124_3590_n155) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U805 ( .A1(n165), .A2(accumulate_reset), .Y(
        DP_OP_102J5_124_3590_n1419) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U816 ( .A1(n248), .A2(
        DP_OP_102J5_124_3590_n2), .Y(DP_OP_102J5_124_3590_n1428) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U799 ( .A1(n270), .A2(accumulate_reset), .Y(
        DP_OP_102J5_124_3590_n137) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U803 ( .A1(n262), .A2(accumulate_reset), .Y(
        DP_OP_102J5_124_3590_n145) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U802 ( .A1(n261), .A2(accumulate_reset), .Y(
        DP_OP_102J5_124_3590_n143) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U804 ( .A1(n260), .A2(accumulate_reset), .Y(
        DP_OP_102J5_124_3590_n147) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U809 ( .A1(n164), .A2(
        DP_OP_102J5_124_3590_n2), .Y(DP_OP_102J5_124_3590_n1421) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U812 ( .A1(n166), .A2(
        DP_OP_102J5_124_3590_n2), .Y(DP_OP_102J5_124_3590_n1424) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U810 ( .A1(n263), .A2(
        DP_OP_102J5_124_3590_n2), .Y(DP_OP_102J5_124_3590_n1422) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U800 ( .A1(n167), .A2(accumulate_reset), .Y(
        DP_OP_102J5_124_3590_n139) );
  OAI21X1_HVT DP_OP_102J5_124_3590_U81 ( .A1(DP_OP_102J5_124_3590_n80), .A2(
        DP_OP_102J5_124_3590_n74), .A3(DP_OP_102J5_124_3590_n75), .Y(
        DP_OP_102J5_124_3590_n73) );
  OAI21X1_HVT DP_OP_102J5_124_3590_U56 ( .A1(DP_OP_102J5_124_3590_n58), .A2(
        DP_OP_102J5_124_3590_n60), .A3(DP_OP_102J5_124_3590_n59), .Y(
        DP_OP_102J5_124_3590_n57) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U11 ( .A1(DP_OP_102J5_124_3590_n29), .A2(
        DP_OP_102J5_124_3590_n32), .Y(DP_OP_102J5_124_3590_n27) );
  OA221X1_HVT U106 ( .A1(1'b0), .A2(DP_OP_102J5_124_3590_n48), .A3(
        DP_OP_102J5_124_3590_n47), .A4(DP_OP_102J5_124_3590_n51), .A5(n107), 
        .Y(n109) );
  OA221X1_HVT U107 ( .A1(1'b0), .A2(DP_OP_102J5_124_3590_n86), .A3(
        DP_OP_102J5_124_3590_n85), .A4(DP_OP_102J5_124_3590_n89), .A5(n105), 
        .Y(DP_OP_102J5_124_3590_n82) );
  OR3X1_HVT U108 ( .A1(n104), .A2(DP_OP_102J5_124_3590_n88), .A3(
        DP_OP_102J5_124_3590_n85), .Y(n105) );
  INVX0_HVT U110 ( .A(DP_OP_102J5_124_3590_n91), .Y(n104) );
  NAND2X0_HVT U111 ( .A1(DP_OP_102J5_124_3590_n45), .A2(
        DP_OP_102J5_124_3590_n54), .Y(n107) );
  OAI21X1_HVT U113 ( .A1(DP_OP_102J5_124_3590_n59), .A2(
        DP_OP_102J5_124_3590_n43), .A3(n109), .Y(DP_OP_102J5_124_3590_n42) );
  NOR2X0_HVT U114 ( .A1(DP_OP_102J5_124_3590_n66), .A2(
        DP_OP_102J5_124_3590_n69), .Y(n110) );
  INVX0_HVT U115 ( .A(DP_OP_102J5_124_3590_n82), .Y(n111) );
  NAND3X0_HVT U116 ( .A1(DP_OP_102J5_124_3590_n72), .A2(n110), .A3(n111), .Y(
        n112) );
  NAND2X0_HVT U117 ( .A1(n110), .A2(DP_OP_102J5_124_3590_n73), .Y(n113) );
  OR2X1_HVT U118 ( .A1(DP_OP_102J5_124_3590_n66), .A2(DP_OP_102J5_124_3590_n70), .Y(n114) );
  NAND4X0_HVT U119 ( .A1(DP_OP_102J5_124_3590_n67), .A2(n112), .A3(n113), .A4(
        n114), .Y(DP_OP_102J5_124_3590_n61) );
  OA21X1_HVT U120 ( .A1(DP_OP_102J5_124_3590_n69), .A2(
        DP_OP_102J5_124_3590_n71), .A3(DP_OP_102J5_124_3590_n70), .Y(n115) );
  INVX0_HVT U121 ( .A(DP_OP_102J5_124_3590_n66), .Y(n116) );
  NAND2X0_HVT U122 ( .A1(n116), .A2(DP_OP_102J5_124_3590_n67), .Y(n117) );
  HADDX1_HVT U123 ( .A0(n115), .B0(n117), .SO(n_accumulator_sum[12]) );
  NAND2X0_HVT U124 ( .A1(DP_OP_102J5_124_3590_n113), .A2(n256), .Y(n118) );
  NAND2X0_HVT U125 ( .A1(DP_OP_102J5_124_3590_n112), .A2(n118), .Y(n162) );
  INVX0_HVT U126 ( .A(DP_OP_102J5_124_3590_n58), .Y(n119) );
  NAND2X0_HVT U127 ( .A1(n119), .A2(DP_OP_102J5_124_3590_n59), .Y(n120) );
  HADDX1_HVT U128 ( .A0(DP_OP_102J5_124_3590_n60), .B0(n120), .SO(
        n_accumulator_sum[13]) );
  NAND2X0_HVT U129 ( .A1(n255), .A2(n162), .Y(n121) );
  AND2X1_HVT U130 ( .A1(n121), .A2(DP_OP_102J5_124_3590_n106), .Y(
        DP_OP_102J5_124_3590_n102) );
  AND2X1_HVT U131 ( .A1(n250), .A2(DP_OP_102J5_124_3590_n56), .Y(n122) );
  HADDX1_HVT U132 ( .A0(n122), .B0(DP_OP_102J5_124_3590_n57), .SO(
        n_accumulator_sum[14]) );
  NAND2X0_HVT U133 ( .A1(DP_OP_102J5_124_3590_n99), .A2(n257), .Y(n123) );
  AND2X1_HVT U134 ( .A1(n123), .A2(DP_OP_102J5_124_3590_n98), .Y(
        DP_OP_102J5_124_3590_n94) );
  NAND2X0_HVT U135 ( .A1(DP_OP_102J5_124_3590_n42), .A2(n259), .Y(n124) );
  AND2X1_HVT U136 ( .A1(n124), .A2(DP_OP_102J5_124_3590_n37), .Y(
        DP_OP_102J5_124_3590_n33) );
  INVX0_HVT U137 ( .A(DP_OP_102J5_124_3590_n50), .Y(n125) );
  NAND2X0_HVT U138 ( .A1(n125), .A2(DP_OP_102J5_124_3590_n51), .Y(n126) );
  HADDX1_HVT U139 ( .A0(DP_OP_102J5_124_3590_n52), .B0(n126), .SO(
        n_accumulator_sum[15]) );
  INVX0_HVT U140 ( .A(DP_OP_102J5_124_3590_n92), .Y(n127) );
  NAND2X0_HVT U141 ( .A1(n127), .A2(DP_OP_102J5_124_3590_n93), .Y(n128) );
  HADDX1_HVT U142 ( .A0(DP_OP_102J5_124_3590_n94), .B0(n128), .SO(
        n_accumulator_sum[6]) );
  AND2X1_HVT U143 ( .A1(DP_OP_102J5_124_3590_n77), .A2(
        DP_OP_102J5_124_3590_n80), .Y(n129) );
  HADDX1_HVT U144 ( .A0(n129), .B0(DP_OP_102J5_124_3590_n81), .SO(
        n_accumulator_sum[9]) );
  OA21X1_HVT U145 ( .A1(DP_OP_102J5_124_3590_n50), .A2(
        DP_OP_102J5_124_3590_n52), .A3(DP_OP_102J5_124_3590_n51), .Y(n130) );
  INVX0_HVT U146 ( .A(DP_OP_102J5_124_3590_n47), .Y(n131) );
  NAND2X0_HVT U147 ( .A1(n131), .A2(DP_OP_102J5_124_3590_n48), .Y(n132) );
  HADDX1_HVT U148 ( .A0(n130), .B0(n132), .SO(n_accumulator_sum[16]) );
  OR2X1_HVT U149 ( .A1(accumulate_reset), .A2(n271), .Y(n133) );
  FADDX1_HVT U150 ( .A(DP_OP_102J5_124_3590_n23), .B(DP_OP_102J5_124_3590_n137), .CI(n133), .S(n_accumulator_sum[22]) );
  AND2X1_HVT U151 ( .A1(DP_OP_102J5_124_3590_n112), .A2(n256), .Y(n134) );
  HADDX1_HVT U152 ( .A0(n134), .B0(DP_OP_102J5_124_3590_n113), .SO(
        n_accumulator_sum[2]) );
  INVX0_HVT U153 ( .A(DP_OP_102J5_124_3590_n100), .Y(n135) );
  NAND2X0_HVT U154 ( .A1(n135), .A2(DP_OP_102J5_124_3590_n101), .Y(n136) );
  HADDX1_HVT U155 ( .A0(DP_OP_102J5_124_3590_n102), .B0(n136), .SO(
        n_accumulator_sum[4]) );
  INVX0_HVT U156 ( .A(DP_OP_102J5_124_3590_n88), .Y(n137) );
  NAND2X0_HVT U157 ( .A1(n137), .A2(DP_OP_102J5_124_3590_n89), .Y(n138) );
  HADDX1_HVT U158 ( .A0(DP_OP_102J5_124_3590_n90), .B0(n138), .SO(
        n_accumulator_sum[7]) );
  INVX0_HVT U159 ( .A(DP_OP_102J5_124_3590_n74), .Y(n139) );
  NAND2X0_HVT U160 ( .A1(DP_OP_102J5_124_3590_n81), .A2(
        DP_OP_102J5_124_3590_n77), .Y(n140) );
  AO22X1_HVT U161 ( .A1(n139), .A2(DP_OP_102J5_124_3590_n75), .A3(
        DP_OP_102J5_124_3590_n80), .A4(n140), .Y(n141) );
  NAND4X0_HVT U162 ( .A1(n139), .A2(DP_OP_102J5_124_3590_n75), .A3(
        DP_OP_102J5_124_3590_n80), .A4(n140), .Y(n142) );
  NAND2X0_HVT U163 ( .A1(n141), .A2(n142), .Y(n_accumulator_sum[10]) );
  INVX0_HVT U164 ( .A(DP_OP_102J5_124_3590_n60), .Y(n143) );
  AOI21X1_HVT U165 ( .A1(DP_OP_102J5_124_3590_n41), .A2(n143), .A3(
        DP_OP_102J5_124_3590_n42), .Y(n144) );
  NAND2X0_HVT U166 ( .A1(n259), .A2(DP_OP_102J5_124_3590_n37), .Y(n145) );
  HADDX1_HVT U167 ( .A0(n144), .B0(n145), .SO(n_accumulator_sum[17]) );
  INVX0_HVT U168 ( .A(DP_OP_102J5_124_3590_n114), .Y(n146) );
  AND2X1_HVT U169 ( .A1(n146), .A2(DP_OP_102J5_124_3590_n115), .Y(n147) );
  HADDX1_HVT U170 ( .A0(n147), .B0(DP_OP_102J5_124_3590_n116), .SO(
        n_accumulator_sum[1]) );
  AND2X1_HVT U171 ( .A1(DP_OP_102J5_124_3590_n106), .A2(n255), .Y(n148) );
  HADDX1_HVT U172 ( .A0(n148), .B0(n162), .SO(n_accumulator_sum[3]) );
  AND2X1_HVT U173 ( .A1(DP_OP_102J5_124_3590_n98), .A2(n257), .Y(n149) );
  HADDX1_HVT U174 ( .A0(n149), .B0(DP_OP_102J5_124_3590_n99), .SO(
        n_accumulator_sum[5]) );
  OA21X1_HVT U175 ( .A1(DP_OP_102J5_124_3590_n88), .A2(
        DP_OP_102J5_124_3590_n90), .A3(DP_OP_102J5_124_3590_n89), .Y(n150) );
  INVX0_HVT U176 ( .A(DP_OP_102J5_124_3590_n85), .Y(n151) );
  NAND2X0_HVT U177 ( .A1(n151), .A2(DP_OP_102J5_124_3590_n86), .Y(n152) );
  HADDX1_HVT U178 ( .A0(n150), .B0(n152), .SO(n_accumulator_sum[8]) );
  INVX0_HVT U179 ( .A(DP_OP_102J5_124_3590_n69), .Y(n153) );
  NAND2X0_HVT U180 ( .A1(n153), .A2(DP_OP_102J5_124_3590_n70), .Y(n154) );
  HADDX1_HVT U181 ( .A0(DP_OP_102J5_124_3590_n71), .B0(n154), .SO(
        n_accumulator_sum[11]) );
  OA21X1_HVT U182 ( .A1(DP_OP_102J5_124_3590_n32), .A2(
        DP_OP_102J5_124_3590_n60), .A3(DP_OP_102J5_124_3590_n33), .Y(n155) );
  INVX0_HVT U183 ( .A(DP_OP_102J5_124_3590_n29), .Y(n156) );
  NAND2X0_HVT U184 ( .A1(n156), .A2(DP_OP_102J5_124_3590_n30), .Y(n157) );
  HADDX1_HVT U185 ( .A0(n155), .B0(n157), .SO(n_accumulator_sum[18]) );
  INVX0_HVT U186 ( .A(DP_OP_102J5_124_3590_n79), .Y(DP_OP_102J5_124_3590_n77)
         );
  INVX2_HVT U187 ( .A(srstn), .Y(n272) );
  INVX1_HVT U188 ( .A(DP_OP_102J5_124_3590_n61), .Y(DP_OP_102J5_124_3590_n60)
         );
  INVX0_HVT U189 ( .A(DP_OP_102J5_124_3590_n116), .Y(DP_OP_102J5_124_3590_n4)
         );
  INVX1_HVT U190 ( .A(n272), .Y(n158) );
  INVX2_HVT U191 ( .A(n158), .Y(n159) );
  INVX2_HVT U192 ( .A(n158), .Y(n160) );
  INVX2_HVT U193 ( .A(n158), .Y(n161) );
  INVX1_HVT U194 ( .A(DP_OP_102J5_124_3590_n2362), .Y(DP_OP_102J5_124_3590_n2)
         );
  INVX1_HVT U195 ( .A(DP_OP_102J5_124_3590_n91), .Y(DP_OP_102J5_124_3590_n90)
         );
  INVX1_HVT U196 ( .A(DP_OP_102J5_124_3590_n82), .Y(DP_OP_102J5_124_3590_n81)
         );
  INVX1_HVT U197 ( .A(accumulate_reset), .Y(DP_OP_102J5_124_3590_n2362) );
  AO21X1_HVT U198 ( .A1(DP_OP_102J5_124_3590_n61), .A2(
        DP_OP_102J5_124_3590_n27), .A3(DP_OP_102J5_124_3590_n28), .Y(n249) );
  OR2X1_HVT U199 ( .A1(DP_OP_102J5_124_3590_n152), .A2(
        DP_OP_102J5_124_3590_n157), .Y(n250) );
  OR2X1_HVT U200 ( .A1(DP_OP_102J5_124_3590_n1149), .A2(
        DP_OP_102J5_124_3590_n1147), .Y(n255) );
  OR2X1_HVT U201 ( .A1(DP_OP_102J5_124_3590_n1271), .A2(
        DP_OP_102J5_124_3590_n1269), .Y(n256) );
  OR2X1_HVT U202 ( .A1(DP_OP_102J5_124_3590_n859), .A2(
        DP_OP_102J5_124_3590_n857), .Y(n257) );
  OR2X1_HVT U203 ( .A1(DP_OP_102J5_124_3590_n147), .A2(
        DP_OP_102J5_124_3590_n146), .Y(n259) );
  INVX1_HVT U204 ( .A(DP_OP_102J5_124_3590_n137), .Y(DP_OP_102J5_124_3590_n138) );
  INVX1_HVT U205 ( .A(DP_OP_102J5_124_3590_n139), .Y(DP_OP_102J5_124_3590_n140) );
  INVX1_HVT U206 ( .A(DP_OP_102J5_124_3590_n141), .Y(DP_OP_102J5_124_3590_n142) );
  INVX1_HVT U207 ( .A(DP_OP_102J5_124_3590_n143), .Y(DP_OP_102J5_124_3590_n144) );
  INVX1_HVT U208 ( .A(DP_OP_102J5_124_3590_n145), .Y(DP_OP_102J5_124_3590_n146) );
  INVX1_HVT U209 ( .A(DP_OP_102J5_124_3590_n147), .Y(DP_OP_102J5_124_3590_n148) );
  INVX1_HVT U210 ( .A(src_window[15]), .Y(DP_OP_102J5_124_3590_n1489) );
  INVX1_HVT U211 ( .A(src_window[14]), .Y(DP_OP_102J5_124_3590_n1490) );
  INVX1_HVT U212 ( .A(src_window[13]), .Y(DP_OP_102J5_124_3590_n1491) );
  INVX1_HVT U213 ( .A(src_window[12]), .Y(DP_OP_102J5_124_3590_n1492) );
  INVX1_HVT U214 ( .A(src_window[11]), .Y(DP_OP_102J5_124_3590_n1493) );
  INVX1_HVT U215 ( .A(src_window[10]), .Y(DP_OP_102J5_124_3590_n1494) );
  INVX1_HVT U216 ( .A(src_window[9]), .Y(DP_OP_102J5_124_3590_n1495) );
  INVX1_HVT U217 ( .A(src_window[8]), .Y(DP_OP_102J5_124_3590_n1496) );
  INVX1_HVT U218 ( .A(src_window[31]), .Y(DP_OP_102J5_124_3590_n1533) );
  INVX1_HVT U219 ( .A(src_window[30]), .Y(DP_OP_102J5_124_3590_n1534) );
  INVX1_HVT U220 ( .A(src_window[29]), .Y(DP_OP_102J5_124_3590_n1535) );
  INVX1_HVT U221 ( .A(src_window[28]), .Y(DP_OP_102J5_124_3590_n1536) );
  INVX1_HVT U222 ( .A(src_window[27]), .Y(DP_OP_102J5_124_3590_n1537) );
  INVX1_HVT U223 ( .A(src_window[26]), .Y(DP_OP_102J5_124_3590_n1538) );
  INVX1_HVT U224 ( .A(src_window[25]), .Y(DP_OP_102J5_124_3590_n1539) );
  INVX1_HVT U225 ( .A(src_window[24]), .Y(DP_OP_102J5_124_3590_n1540) );
  INVX1_HVT U226 ( .A(DP_OP_102J5_124_3590_n155), .Y(DP_OP_102J5_124_3590_n156) );
  INVX1_HVT U227 ( .A(src_window[47]), .Y(DP_OP_102J5_124_3590_n1577) );
  INVX1_HVT U228 ( .A(src_window[46]), .Y(DP_OP_102J5_124_3590_n1578) );
  INVX1_HVT U229 ( .A(src_window[45]), .Y(DP_OP_102J5_124_3590_n1579) );
  INVX1_HVT U230 ( .A(src_window[44]), .Y(DP_OP_102J5_124_3590_n1580) );
  INVX1_HVT U231 ( .A(src_window[43]), .Y(DP_OP_102J5_124_3590_n1581) );
  INVX1_HVT U232 ( .A(src_window[42]), .Y(DP_OP_102J5_124_3590_n1582) );
  INVX1_HVT U233 ( .A(src_window[41]), .Y(DP_OP_102J5_124_3590_n1583) );
  INVX1_HVT U234 ( .A(src_window[40]), .Y(DP_OP_102J5_124_3590_n1584) );
  INVX1_HVT U235 ( .A(src_window[63]), .Y(DP_OP_102J5_124_3590_n1621) );
  INVX1_HVT U236 ( .A(src_window[62]), .Y(DP_OP_102J5_124_3590_n1622) );
  INVX1_HVT U237 ( .A(src_window[61]), .Y(DP_OP_102J5_124_3590_n1623) );
  INVX1_HVT U238 ( .A(src_window[60]), .Y(DP_OP_102J5_124_3590_n1624) );
  INVX1_HVT U239 ( .A(src_window[59]), .Y(DP_OP_102J5_124_3590_n1625) );
  INVX1_HVT U240 ( .A(src_window[58]), .Y(DP_OP_102J5_124_3590_n1626) );
  INVX1_HVT U241 ( .A(src_window[57]), .Y(DP_OP_102J5_124_3590_n1627) );
  INVX1_HVT U242 ( .A(src_window[56]), .Y(DP_OP_102J5_124_3590_n1628) );
  INVX1_HVT U243 ( .A(DP_OP_102J5_124_3590_n165), .Y(DP_OP_102J5_124_3590_n166) );
  INVX1_HVT U244 ( .A(src_window[79]), .Y(DP_OP_102J5_124_3590_n1665) );
  INVX1_HVT U245 ( .A(src_window[78]), .Y(DP_OP_102J5_124_3590_n1666) );
  INVX1_HVT U246 ( .A(src_window[77]), .Y(DP_OP_102J5_124_3590_n1667) );
  INVX1_HVT U247 ( .A(src_window[76]), .Y(DP_OP_102J5_124_3590_n1668) );
  INVX1_HVT U248 ( .A(src_window[75]), .Y(DP_OP_102J5_124_3590_n1669) );
  INVX1_HVT U249 ( .A(src_window[74]), .Y(DP_OP_102J5_124_3590_n1670) );
  INVX1_HVT U250 ( .A(src_window[73]), .Y(DP_OP_102J5_124_3590_n1671) );
  INVX1_HVT U251 ( .A(src_window[72]), .Y(DP_OP_102J5_124_3590_n1672) );
  INVX1_HVT U252 ( .A(src_window[95]), .Y(DP_OP_102J5_124_3590_n1709) );
  INVX1_HVT U253 ( .A(src_window[94]), .Y(DP_OP_102J5_124_3590_n1710) );
  INVX1_HVT U254 ( .A(src_window[93]), .Y(DP_OP_102J5_124_3590_n1711) );
  INVX1_HVT U255 ( .A(src_window[92]), .Y(DP_OP_102J5_124_3590_n1712) );
  INVX1_HVT U256 ( .A(src_window[91]), .Y(DP_OP_102J5_124_3590_n1713) );
  INVX1_HVT U257 ( .A(src_window[90]), .Y(DP_OP_102J5_124_3590_n1714) );
  INVX1_HVT U258 ( .A(src_window[89]), .Y(DP_OP_102J5_124_3590_n1715) );
  INVX1_HVT U259 ( .A(src_window[88]), .Y(DP_OP_102J5_124_3590_n1716) );
  INVX1_HVT U260 ( .A(src_window[111]), .Y(DP_OP_102J5_124_3590_n1753) );
  INVX1_HVT U261 ( .A(src_window[110]), .Y(DP_OP_102J5_124_3590_n1754) );
  INVX1_HVT U262 ( .A(src_window[109]), .Y(DP_OP_102J5_124_3590_n1755) );
  INVX1_HVT U263 ( .A(src_window[108]), .Y(DP_OP_102J5_124_3590_n1756) );
  INVX1_HVT U264 ( .A(src_window[107]), .Y(DP_OP_102J5_124_3590_n1757) );
  INVX1_HVT U265 ( .A(src_window[106]), .Y(DP_OP_102J5_124_3590_n1758) );
  INVX1_HVT U266 ( .A(src_window[105]), .Y(DP_OP_102J5_124_3590_n1759) );
  INVX1_HVT U267 ( .A(src_window[104]), .Y(DP_OP_102J5_124_3590_n1760) );
  INVX1_HVT U268 ( .A(src_window[127]), .Y(DP_OP_102J5_124_3590_n1796) );
  INVX1_HVT U269 ( .A(src_window[126]), .Y(DP_OP_102J5_124_3590_n1797) );
  INVX1_HVT U270 ( .A(src_window[125]), .Y(DP_OP_102J5_124_3590_n1798) );
  INVX1_HVT U271 ( .A(src_window[124]), .Y(DP_OP_102J5_124_3590_n1799) );
  INVX1_HVT U272 ( .A(src_window[123]), .Y(DP_OP_102J5_124_3590_n1800) );
  INVX1_HVT U273 ( .A(src_window[122]), .Y(DP_OP_102J5_124_3590_n1801) );
  INVX1_HVT U274 ( .A(src_window[121]), .Y(DP_OP_102J5_124_3590_n1802) );
  INVX1_HVT U275 ( .A(src_window[120]), .Y(DP_OP_102J5_124_3590_n1803) );
  INVX1_HVT U276 ( .A(src_window[143]), .Y(DP_OP_102J5_124_3590_n1840) );
  INVX1_HVT U277 ( .A(src_window[142]), .Y(DP_OP_102J5_124_3590_n1841) );
  INVX1_HVT U278 ( .A(src_window[141]), .Y(DP_OP_102J5_124_3590_n1842) );
  INVX1_HVT U279 ( .A(src_window[140]), .Y(DP_OP_102J5_124_3590_n1843) );
  INVX1_HVT U280 ( .A(src_window[139]), .Y(DP_OP_102J5_124_3590_n1844) );
  INVX1_HVT U281 ( .A(src_window[138]), .Y(DP_OP_102J5_124_3590_n1845) );
  INVX1_HVT U282 ( .A(src_window[137]), .Y(DP_OP_102J5_124_3590_n1846) );
  INVX1_HVT U283 ( .A(src_window[136]), .Y(DP_OP_102J5_124_3590_n1847) );
  INVX1_HVT U284 ( .A(src_window[159]), .Y(DP_OP_102J5_124_3590_n1884) );
  INVX1_HVT U285 ( .A(src_window[158]), .Y(DP_OP_102J5_124_3590_n1885) );
  INVX1_HVT U286 ( .A(src_window[157]), .Y(DP_OP_102J5_124_3590_n1886) );
  INVX1_HVT U287 ( .A(src_window[156]), .Y(DP_OP_102J5_124_3590_n1887) );
  INVX1_HVT U288 ( .A(src_window[155]), .Y(DP_OP_102J5_124_3590_n1888) );
  INVX1_HVT U289 ( .A(src_window[154]), .Y(DP_OP_102J5_124_3590_n1889) );
  INVX1_HVT U290 ( .A(src_window[153]), .Y(DP_OP_102J5_124_3590_n1890) );
  INVX1_HVT U291 ( .A(src_window[152]), .Y(DP_OP_102J5_124_3590_n1891) );
  INVX1_HVT U292 ( .A(src_window[151]), .Y(DP_OP_102J5_124_3590_n1928) );
  INVX1_HVT U293 ( .A(src_window[150]), .Y(DP_OP_102J5_124_3590_n1929) );
  INVX1_HVT U294 ( .A(src_window[149]), .Y(DP_OP_102J5_124_3590_n1930) );
  INVX1_HVT U295 ( .A(src_window[148]), .Y(DP_OP_102J5_124_3590_n1931) );
  INVX1_HVT U296 ( .A(src_window[147]), .Y(DP_OP_102J5_124_3590_n1932) );
  INVX1_HVT U297 ( .A(src_window[146]), .Y(DP_OP_102J5_124_3590_n1933) );
  INVX1_HVT U298 ( .A(src_window[145]), .Y(DP_OP_102J5_124_3590_n1934) );
  INVX1_HVT U299 ( .A(src_window[144]), .Y(DP_OP_102J5_124_3590_n1935) );
  INVX1_HVT U300 ( .A(src_window[135]), .Y(DP_OP_102J5_124_3590_n1972) );
  INVX1_HVT U301 ( .A(src_window[134]), .Y(DP_OP_102J5_124_3590_n1973) );
  INVX1_HVT U302 ( .A(src_window[133]), .Y(DP_OP_102J5_124_3590_n1974) );
  INVX1_HVT U303 ( .A(src_window[132]), .Y(DP_OP_102J5_124_3590_n1975) );
  INVX1_HVT U304 ( .A(src_window[131]), .Y(DP_OP_102J5_124_3590_n1976) );
  INVX1_HVT U305 ( .A(src_window[130]), .Y(DP_OP_102J5_124_3590_n1977) );
  INVX1_HVT U306 ( .A(src_window[129]), .Y(DP_OP_102J5_124_3590_n1978) );
  INVX1_HVT U307 ( .A(src_window[128]), .Y(DP_OP_102J5_124_3590_n1979) );
  INVX1_HVT U308 ( .A(src_window[119]), .Y(DP_OP_102J5_124_3590_n2016) );
  INVX1_HVT U309 ( .A(src_window[118]), .Y(DP_OP_102J5_124_3590_n2017) );
  INVX1_HVT U310 ( .A(src_window[117]), .Y(DP_OP_102J5_124_3590_n2018) );
  INVX1_HVT U311 ( .A(src_window[116]), .Y(DP_OP_102J5_124_3590_n2019) );
  INVX1_HVT U312 ( .A(src_window[115]), .Y(DP_OP_102J5_124_3590_n2020) );
  INVX1_HVT U313 ( .A(src_window[114]), .Y(DP_OP_102J5_124_3590_n2021) );
  INVX1_HVT U314 ( .A(src_window[113]), .Y(DP_OP_102J5_124_3590_n2022) );
  INVX1_HVT U315 ( .A(src_window[112]), .Y(DP_OP_102J5_124_3590_n2023) );
  INVX1_HVT U316 ( .A(src_window[103]), .Y(DP_OP_102J5_124_3590_n2060) );
  INVX1_HVT U317 ( .A(src_window[102]), .Y(DP_OP_102J5_124_3590_n2061) );
  INVX1_HVT U318 ( .A(src_window[101]), .Y(DP_OP_102J5_124_3590_n2062) );
  INVX1_HVT U319 ( .A(src_window[100]), .Y(DP_OP_102J5_124_3590_n2063) );
  INVX1_HVT U320 ( .A(src_window[99]), .Y(DP_OP_102J5_124_3590_n2064) );
  INVX1_HVT U321 ( .A(src_window[98]), .Y(DP_OP_102J5_124_3590_n2065) );
  INVX1_HVT U322 ( .A(src_window[97]), .Y(DP_OP_102J5_124_3590_n2066) );
  INVX1_HVT U323 ( .A(src_window[96]), .Y(DP_OP_102J5_124_3590_n2067) );
  INVX1_HVT U324 ( .A(src_window[87]), .Y(DP_OP_102J5_124_3590_n2104) );
  INVX1_HVT U325 ( .A(src_window[86]), .Y(DP_OP_102J5_124_3590_n2105) );
  INVX1_HVT U326 ( .A(src_window[85]), .Y(DP_OP_102J5_124_3590_n2106) );
  INVX1_HVT U327 ( .A(src_window[84]), .Y(DP_OP_102J5_124_3590_n2107) );
  INVX1_HVT U328 ( .A(src_window[83]), .Y(DP_OP_102J5_124_3590_n2108) );
  INVX1_HVT U329 ( .A(src_window[82]), .Y(DP_OP_102J5_124_3590_n2109) );
  INVX1_HVT U330 ( .A(src_window[81]), .Y(DP_OP_102J5_124_3590_n2110) );
  INVX1_HVT U331 ( .A(src_window[80]), .Y(DP_OP_102J5_124_3590_n2111) );
  INVX1_HVT U332 ( .A(src_window[71]), .Y(DP_OP_102J5_124_3590_n2148) );
  INVX1_HVT U333 ( .A(src_window[70]), .Y(DP_OP_102J5_124_3590_n2149) );
  INVX1_HVT U334 ( .A(src_window[69]), .Y(DP_OP_102J5_124_3590_n2150) );
  INVX1_HVT U335 ( .A(src_window[68]), .Y(DP_OP_102J5_124_3590_n2151) );
  INVX1_HVT U336 ( .A(src_window[67]), .Y(DP_OP_102J5_124_3590_n2152) );
  INVX1_HVT U337 ( .A(src_window[66]), .Y(DP_OP_102J5_124_3590_n2153) );
  INVX1_HVT U338 ( .A(src_window[65]), .Y(DP_OP_102J5_124_3590_n2154) );
  INVX1_HVT U339 ( .A(src_window[64]), .Y(DP_OP_102J5_124_3590_n2155) );
  INVX1_HVT U340 ( .A(src_window[55]), .Y(DP_OP_102J5_124_3590_n2192) );
  INVX1_HVT U341 ( .A(src_window[54]), .Y(DP_OP_102J5_124_3590_n2193) );
  INVX1_HVT U342 ( .A(src_window[53]), .Y(DP_OP_102J5_124_3590_n2194) );
  INVX1_HVT U343 ( .A(src_window[52]), .Y(DP_OP_102J5_124_3590_n2195) );
  INVX1_HVT U344 ( .A(src_window[51]), .Y(DP_OP_102J5_124_3590_n2196) );
  INVX1_HVT U345 ( .A(src_window[50]), .Y(DP_OP_102J5_124_3590_n2197) );
  INVX1_HVT U346 ( .A(src_window[49]), .Y(DP_OP_102J5_124_3590_n2198) );
  INVX1_HVT U347 ( .A(src_window[48]), .Y(DP_OP_102J5_124_3590_n2199) );
  INVX1_HVT U348 ( .A(DP_OP_102J5_124_3590_n221), .Y(DP_OP_102J5_124_3590_n222) );
  INVX1_HVT U349 ( .A(src_window[39]), .Y(DP_OP_102J5_124_3590_n2236) );
  INVX1_HVT U350 ( .A(src_window[38]), .Y(DP_OP_102J5_124_3590_n2237) );
  INVX1_HVT U351 ( .A(src_window[37]), .Y(DP_OP_102J5_124_3590_n2238) );
  INVX1_HVT U352 ( .A(src_window[36]), .Y(DP_OP_102J5_124_3590_n2239) );
  INVX1_HVT U353 ( .A(src_window[35]), .Y(DP_OP_102J5_124_3590_n2240) );
  INVX1_HVT U354 ( .A(src_window[34]), .Y(DP_OP_102J5_124_3590_n2241) );
  INVX1_HVT U355 ( .A(src_window[33]), .Y(DP_OP_102J5_124_3590_n2242) );
  INVX1_HVT U356 ( .A(src_window[32]), .Y(DP_OP_102J5_124_3590_n2243) );
  INVX1_HVT U357 ( .A(src_window[23]), .Y(DP_OP_102J5_124_3590_n2280) );
  INVX1_HVT U358 ( .A(src_window[22]), .Y(DP_OP_102J5_124_3590_n2281) );
  INVX1_HVT U359 ( .A(src_window[21]), .Y(DP_OP_102J5_124_3590_n2282) );
  INVX1_HVT U360 ( .A(src_window[20]), .Y(DP_OP_102J5_124_3590_n2283) );
  INVX1_HVT U361 ( .A(src_window[19]), .Y(DP_OP_102J5_124_3590_n2284) );
  INVX1_HVT U362 ( .A(src_window[18]), .Y(DP_OP_102J5_124_3590_n2285) );
  INVX1_HVT U363 ( .A(src_window[17]), .Y(DP_OP_102J5_124_3590_n2286) );
  INVX1_HVT U364 ( .A(src_window[16]), .Y(DP_OP_102J5_124_3590_n2287) );
  INVX1_HVT U365 ( .A(src_window[7]), .Y(DP_OP_102J5_124_3590_n2323) );
  INVX1_HVT U366 ( .A(src_window[6]), .Y(DP_OP_102J5_124_3590_n2324) );
  INVX1_HVT U367 ( .A(src_window[5]), .Y(DP_OP_102J5_124_3590_n2325) );
  INVX1_HVT U368 ( .A(src_window[4]), .Y(DP_OP_102J5_124_3590_n2326) );
  INVX1_HVT U369 ( .A(src_window[3]), .Y(DP_OP_102J5_124_3590_n2327) );
  INVX1_HVT U370 ( .A(src_window[2]), .Y(DP_OP_102J5_124_3590_n2328) );
  INVX1_HVT U371 ( .A(src_window[1]), .Y(DP_OP_102J5_124_3590_n2329) );
  INVX1_HVT U372 ( .A(src_window[0]), .Y(DP_OP_102J5_124_3590_n2330) );
  INVX1_HVT U373 ( .A(DP_OP_102J5_124_3590_n404), .Y(DP_OP_102J5_124_3590_n405) );
  INVX1_HVT U374 ( .A(DP_OP_102J5_124_3590_n56), .Y(DP_OP_102J5_124_3590_n54)
         );
  INVX1_HVT U375 ( .A(DP_OP_102J5_124_3590_n700), .Y(DP_OP_102J5_124_3590_n701) );
endmodule


module fc_quantize ( clk, srstn, fc_state, quantized_data, 
        unquautized_data_22_, unquautized_data_21_, unquautized_data_20_, 
        unquautized_data_19_, unquautized_data_18_, unquautized_data_17_, 
        unquautized_data_16_, unquautized_data_15_, unquautized_data_14_, 
        unquautized_data_13_, unquautized_data_12_, unquautized_data_11_, 
        unquautized_data_10_, unquautized_data_9_, unquautized_data_8_, 
        unquautized_data_7_, unquautized_data_6_, unquautized_data_5_, 
        unquautized_data_4_ );
  output [7:0] quantized_data;
  input clk, srstn, fc_state, unquautized_data_22_, unquautized_data_21_,
         unquautized_data_20_, unquautized_data_19_, unquautized_data_18_,
         unquautized_data_17_, unquautized_data_16_, unquautized_data_15_,
         unquautized_data_14_, unquautized_data_13_, unquautized_data_12_,
         unquautized_data_11_, unquautized_data_10_, unquautized_data_9_,
         unquautized_data_8_, unquautized_data_7_, unquautized_data_6_,
         unquautized_data_5_, unquautized_data_4_;
  wire   n13, n1, n2, n4, n5, n6, n7, n10, n11, n12, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82;
  wire   [7:0] n_quantized_data;

  DFFSSRX1_HVT quantized_data_reg_7_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[7]), .CLK(clk), .Q(quantized_data[7]) );
  DFFSSRX1_HVT quantized_data_reg_6_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[6]), .CLK(clk), .Q(quantized_data[6]) );
  DFFSSRX1_HVT quantized_data_reg_5_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[5]), .CLK(clk), .Q(quantized_data[5]) );
  DFFSSRX1_HVT quantized_data_reg_4_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[4]), .CLK(clk), .Q(quantized_data[4]) );
  DFFSSRX1_HVT quantized_data_reg_3_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[3]), .CLK(clk), .Q(quantized_data[3]) );
  DFFSSRX1_HVT quantized_data_reg_2_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[2]), .CLK(clk), .Q(quantized_data[2]) );
  DFFSSRX1_HVT quantized_data_reg_1_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[1]), .CLK(clk), .Q(quantized_data[1]) );
  DFFSSRX1_HVT quantized_data_reg_0_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[0]), .CLK(clk), .Q(quantized_data[0]) );
  AO221X1_HVT U3 ( .A1(1'b1), .A2(n67), .A3(n59), .A4(n6), .A5(n7), .Y(n10) );
  AO221X1_HVT U4 ( .A1(1'b1), .A2(n58), .A3(n49), .A4(n1), .A5(n2), .Y(n4) );
  NAND3X0_HVT U5 ( .A1(unquautized_data_6_), .A2(unquautized_data_5_), .A3(
        unquautized_data_4_), .Y(n1) );
  INVX0_HVT U6 ( .A(n66), .Y(n2) );
  AO21X1_HVT U8 ( .A1(n55), .A2(n50), .A3(n53), .Y(n5) );
  NAND3X0_HVT U9 ( .A1(n81), .A2(n4), .A3(n5), .Y(n_quantized_data[2]) );
  NAND2X0_HVT U10 ( .A1(unquautized_data_8_), .A2(n58), .Y(n6) );
  INVX0_HVT U11 ( .A(n66), .Y(n7) );
  AO21X1_HVT U13 ( .A1(n65), .A2(n60), .A3(n63), .Y(n11) );
  NAND3X0_HVT U14 ( .A1(n81), .A2(n10), .A3(n11), .Y(n_quantized_data[4]) );
  INVX1_HVT U15 ( .A(n33), .Y(n78) );
  INVX0_HVT U16 ( .A(n21), .Y(n73) );
  INVX0_HVT U17 ( .A(unquautized_data_15_), .Y(n25) );
  INVX0_HVT U18 ( .A(unquautized_data_19_), .Y(n27) );
  INVX0_HVT U19 ( .A(unquautized_data_20_), .Y(n23) );
  INVX0_HVT U20 ( .A(unquautized_data_21_), .Y(n24) );
  INVX0_HVT U21 ( .A(unquautized_data_13_), .Y(n22) );
  INVX0_HVT U22 ( .A(unquautized_data_9_), .Y(n59) );
  INVX0_HVT U23 ( .A(unquautized_data_7_), .Y(n49) );
  INVX0_HVT U24 ( .A(unquautized_data_6_), .Y(n45) );
  INVX0_HVT U25 ( .A(unquautized_data_5_), .Y(n39) );
  INVX1_HVT U26 ( .A(srstn), .Y(n13) );
  INVX1_HVT U27 ( .A(n70), .Y(n66) );
  INVX1_HVT U28 ( .A(n41), .Y(n81) );
  OR2X1_HVT U29 ( .A1(n72), .A2(n71), .Y(n21) );
  INVX1_HVT U30 ( .A(unquautized_data_22_), .Y(n36) );
  INVX1_HVT U31 ( .A(unquautized_data_10_), .Y(n65) );
  INVX1_HVT U32 ( .A(unquautized_data_8_), .Y(n55) );
  INVX1_HVT U33 ( .A(n75), .Y(n61) );
  INVX1_HVT U34 ( .A(fc_state), .Y(n20) );
  INVX1_HVT U35 ( .A(unquautized_data_17_), .Y(n34) );
  INVX1_HVT U36 ( .A(n60), .Y(n74) );
  INVX1_HVT U37 ( .A(n50), .Y(n51) );
  INVX1_HVT U38 ( .A(unquautized_data_12_), .Y(n77) );
  INVX1_HVT U39 ( .A(unquautized_data_11_), .Y(n71) );
  NAND2X0_HVT U40 ( .A1(n77), .A2(n76), .Y(n12) );
  NAND3X0_HVT U41 ( .A1(n61), .A2(n33), .A3(n12), .Y(n79) );
  NAND2X0_HVT U42 ( .A1(n72), .A2(n71), .Y(n14) );
  NAND3X0_HVT U43 ( .A1(n66), .A2(n21), .A3(n14), .Y(n80) );
  AND4X1_HVT U44 ( .A1(unquautized_data_20_), .A2(unquautized_data_19_), .A3(
        unquautized_data_18_), .A4(unquautized_data_17_), .Y(n15) );
  AND4X1_HVT U45 ( .A1(unquautized_data_16_), .A2(unquautized_data_14_), .A3(
        unquautized_data_21_), .A4(n15), .Y(n16) );
  NAND3X0_HVT U46 ( .A1(unquautized_data_13_), .A2(unquautized_data_15_), .A3(
        n16), .Y(n19) );
  AND4X1_HVT U47 ( .A1(unquautized_data_6_), .A2(unquautized_data_5_), .A3(
        unquautized_data_4_), .A4(unquautized_data_7_), .Y(n58) );
  AND3X1_HVT U48 ( .A1(n58), .A2(unquautized_data_8_), .A3(unquautized_data_9_), .Y(n67) );
  NAND2X0_HVT U49 ( .A1(n67), .A2(unquautized_data_10_), .Y(n72) );
  OR3X1_HVT U50 ( .A1(n19), .A2(n21), .A3(n77), .Y(n17) );
  HADDX1_HVT U51 ( .A0(n36), .B0(n17), .SO(n82) );
  HADDX1_HVT U52 ( .A0(unquautized_data_12_), .B0(n21), .SO(n18) );
  AO221X1_HVT U53 ( .A1(n82), .A2(n19), .A3(n82), .A4(n18), .A5(n20), .Y(n70)
         );
  NAND2X0_HVT U54 ( .A1(n36), .A2(n20), .Y(n75) );
  OAI22X1_HVT U55 ( .A1(unquautized_data_4_), .A2(n70), .A3(
        unquautized_data_6_), .A4(n75), .Y(n40) );
  AO22X1_HVT U56 ( .A1(unquautized_data_6_), .A2(n61), .A3(unquautized_data_4_), .A4(n66), .Y(n38) );
  OA221X1_HVT U57 ( .A1(unquautized_data_12_), .A2(n73), .A3(n77), .A4(n21), 
        .A5(n36), .Y(n37) );
  NAND3X0_HVT U58 ( .A1(unquautized_data_6_), .A2(unquautized_data_5_), .A3(
        unquautized_data_7_), .Y(n50) );
  NAND3X0_HVT U59 ( .A1(unquautized_data_8_), .A2(unquautized_data_9_), .A3(
        n51), .Y(n60) );
  NAND4X0_HVT U60 ( .A1(unquautized_data_10_), .A2(unquautized_data_12_), .A3(
        unquautized_data_11_), .A4(n74), .Y(n33) );
  OA222X1_HVT U61 ( .A1(n22), .A2(n78), .A3(n22), .A4(unquautized_data_15_), 
        .A5(n33), .A6(unquautized_data_13_), .Y(n31) );
  OA222X1_HVT U62 ( .A1(unquautized_data_20_), .A2(n24), .A3(n23), .A4(n78), 
        .A5(unquautized_data_21_), .A6(n33), .Y(n30) );
  OA22X1_HVT U63 ( .A1(unquautized_data_16_), .A2(n34), .A3(
        unquautized_data_14_), .A4(n25), .Y(n26) );
  OA221X1_HVT U64 ( .A1(unquautized_data_19_), .A2(n33), .A3(n27), .A4(
        unquautized_data_18_), .A5(n26), .Y(n29) );
  OAI21X1_HVT U65 ( .A1(unquautized_data_18_), .A2(unquautized_data_16_), .A3(
        n33), .Y(n28) );
  NAND4X0_HVT U66 ( .A1(n31), .A2(n30), .A3(n29), .A4(n28), .Y(n32) );
  AO221X1_HVT U67 ( .A1(n78), .A2(n34), .A3(n33), .A4(unquautized_data_14_), 
        .A5(n32), .Y(n35) );
  AO22X1_HVT U68 ( .A1(n37), .A2(fc_state), .A3(n36), .A4(n35), .Y(n41) );
  AO221X1_HVT U69 ( .A1(unquautized_data_5_), .A2(n40), .A3(n39), .A4(n38), 
        .A5(n41), .Y(n_quantized_data[0]) );
  NAND3X0_HVT U70 ( .A1(unquautized_data_5_), .A2(n61), .A3(n49), .Y(n44) );
  NAND2X0_HVT U71 ( .A1(unquautized_data_5_), .A2(unquautized_data_4_), .Y(n42) );
  HADDX1_HVT U72 ( .A0(unquautized_data_6_), .B0(n42), .SO(n43) );
  OA22X1_HVT U73 ( .A1(n45), .A2(n44), .A3(n70), .A4(n43), .Y(n48) );
  NAND2X0_HVT U74 ( .A1(unquautized_data_6_), .A2(unquautized_data_5_), .Y(n46) );
  NAND3X0_HVT U75 ( .A1(unquautized_data_7_), .A2(n61), .A3(n46), .Y(n47) );
  NAND3X0_HVT U76 ( .A1(n81), .A2(n48), .A3(n47), .Y(n_quantized_data[1]) );
  AO21X1_HVT U77 ( .A1(unquautized_data_8_), .A2(n51), .A3(n75), .Y(n53) );
  NAND2X0_HVT U78 ( .A1(n51), .A2(n61), .Y(n52) );
  OA22X1_HVT U79 ( .A1(unquautized_data_9_), .A2(n52), .A3(n58), .A4(n70), .Y(
        n54) );
  OA22X1_HVT U80 ( .A1(n54), .A2(n55), .A3(n59), .A4(n53), .Y(n57) );
  NAND3X0_HVT U81 ( .A1(n58), .A2(n66), .A3(n55), .Y(n56) );
  NAND3X0_HVT U82 ( .A1(n81), .A2(n57), .A3(n56), .Y(n_quantized_data[3]) );
  AO21X1_HVT U83 ( .A1(unquautized_data_10_), .A2(n74), .A3(n75), .Y(n63) );
  NAND2X0_HVT U84 ( .A1(n74), .A2(n61), .Y(n62) );
  OA22X1_HVT U85 ( .A1(unquautized_data_11_), .A2(n62), .A3(n67), .A4(n70), 
        .Y(n64) );
  OA22X1_HVT U86 ( .A1(n64), .A2(n65), .A3(n71), .A4(n63), .Y(n69) );
  NAND3X0_HVT U87 ( .A1(n67), .A2(n66), .A3(n65), .Y(n68) );
  NAND3X0_HVT U88 ( .A1(n81), .A2(n69), .A3(n68), .Y(n_quantized_data[5]) );
  NAND3X0_HVT U89 ( .A1(unquautized_data_10_), .A2(unquautized_data_11_), .A3(
        n74), .Y(n76) );
  NAND3X0_HVT U90 ( .A1(n81), .A2(n80), .A3(n79), .Y(n_quantized_data[6]) );
  AND2X1_HVT U91 ( .A1(n82), .A2(fc_state), .Y(n_quantized_data[7]) );
endmodule


module fc_top ( clk, srstn, conv_done, mem_sel, sram_rdata_c0, sram_rdata_c1, 
        sram_rdata_c2, sram_rdata_c3, sram_rdata_c4, sram_raddr_c0, 
        sram_raddr_c1, sram_raddr_c2, sram_raddr_c3, sram_raddr_c4, 
        sram_rdata_d0, sram_rdata_d1, sram_rdata_d2, sram_rdata_d3, 
        sram_rdata_d4, sram_raddr_d0, sram_raddr_d1, sram_raddr_d2, 
        sram_raddr_d3, sram_raddr_d4, sram_rdata_e0, sram_rdata_e1, 
        sram_rdata_e2, sram_rdata_e3, sram_rdata_e4, sram_raddr_e0, 
        sram_raddr_e1, sram_raddr_e2, sram_raddr_e3, sram_raddr_e4, 
        sram_write_enable_e0, sram_write_enable_e1, sram_write_enable_e2, 
        sram_write_enable_e3, sram_write_enable_e4, sram_bytemask_e, 
        sram_waddr_e, sram_wdata_e, sram_write_enable_f, sram_bytemask_f, 
        sram_waddr_f, sram_wdata_f, sram_rdata_weight, sram_raddr_weight, 
        fc1_done, fc2_done );
  input [31:0] sram_rdata_c0;
  input [31:0] sram_rdata_c1;
  input [31:0] sram_rdata_c2;
  input [31:0] sram_rdata_c3;
  input [31:0] sram_rdata_c4;
  output [5:0] sram_raddr_c0;
  output [5:0] sram_raddr_c1;
  output [5:0] sram_raddr_c2;
  output [5:0] sram_raddr_c3;
  output [5:0] sram_raddr_c4;
  input [31:0] sram_rdata_d0;
  input [31:0] sram_rdata_d1;
  input [31:0] sram_rdata_d2;
  input [31:0] sram_rdata_d3;
  input [31:0] sram_rdata_d4;
  output [5:0] sram_raddr_d0;
  output [5:0] sram_raddr_d1;
  output [5:0] sram_raddr_d2;
  output [5:0] sram_raddr_d3;
  output [5:0] sram_raddr_d4;
  input [31:0] sram_rdata_e0;
  input [31:0] sram_rdata_e1;
  input [31:0] sram_rdata_e2;
  input [31:0] sram_rdata_e3;
  input [31:0] sram_rdata_e4;
  output [4:0] sram_raddr_e0;
  output [4:0] sram_raddr_e1;
  output [4:0] sram_raddr_e2;
  output [4:0] sram_raddr_e3;
  output [4:0] sram_raddr_e4;
  output [3:0] sram_bytemask_e;
  output [4:0] sram_waddr_e;
  output [7:0] sram_wdata_e;
  output [3:0] sram_bytemask_f;
  output [1:0] sram_waddr_f;
  output [7:0] sram_wdata_f;
  input [79:0] sram_rdata_weight;
  output [14:0] sram_raddr_weight;
  input clk, srstn, conv_done, mem_sel;
  output sram_write_enable_e0, sram_write_enable_e1, sram_write_enable_e2,
         sram_write_enable_e3, sram_write_enable_e4, sram_write_enable_f,
         fc1_done, fc2_done;
  wire   accumulate_reset, fc_state, data_out_22_, data_out_21_, data_out_20_,
         data_out_19_, data_out_18_, data_out_17_, data_out_16_, data_out_15_,
         data_out_14_, data_out_13_, data_out_12_, data_out_11_, data_out_10_,
         data_out_9_, data_out_8_, data_out_7_, data_out_6_, data_out_5_,
         data_out_4_, data_out_3_, data_out_2_, data_out_1_, data_out_0_,
         SYNOPSYS_UNCONNECTED_1;
  wire   [1:0] sram_sel;
  wire   [159:0] src_window;

  fc_controller fc_controller ( .clk(clk), .srstn(srstn), .conv_done(conv_done), .mem_sel(mem_sel), .accumulate_reset(accumulate_reset), .fc_state(fc_state), 
        .sram_sel(sram_sel), .sram_raddr_c0(sram_raddr_c0), .sram_raddr_c1(
        sram_raddr_c1), .sram_raddr_c2(sram_raddr_c2), .sram_raddr_c3(
        sram_raddr_c3), .sram_raddr_c4(sram_raddr_c4), .sram_raddr_d0(
        sram_raddr_d0), .sram_raddr_d1(sram_raddr_d1), .sram_raddr_d2(
        sram_raddr_d2), .sram_raddr_d3(sram_raddr_d3), .sram_raddr_d4(
        sram_raddr_d4), .sram_raddr_e0(sram_raddr_e0), .sram_raddr_e1(
        sram_raddr_e1), .sram_raddr_e2(sram_raddr_e2), .sram_raddr_e3(
        sram_raddr_e3), .sram_raddr_e4(sram_raddr_e4), .sram_write_enable_e0(
        sram_write_enable_e0), .sram_write_enable_e1(sram_write_enable_e1), 
        .sram_write_enable_e2(sram_write_enable_e2), .sram_write_enable_e3(
        sram_write_enable_e3), .sram_write_enable_e4(sram_write_enable_e4), 
        .sram_write_enable_f(sram_write_enable_f), .sram_waddr({
        SYNOPSYS_UNCONNECTED_1, sram_waddr_e}), .sram_bytemask(sram_bytemask_e), .sram_raddr_weight(sram_raddr_weight), .fc1_done(fc1_done), .fc2_done(
        fc2_done) );
  fc_data_reg fc_data_reg ( .clk(clk), .srstn(srstn), .sram_rdata_c0(
        sram_rdata_c0), .sram_rdata_c1(sram_rdata_c1), .sram_rdata_c2(
        sram_rdata_c2), .sram_rdata_c3(sram_rdata_c3), .sram_rdata_c4(
        sram_rdata_c4), .sram_rdata_d0(sram_rdata_d0), .sram_rdata_d1(
        sram_rdata_d1), .sram_rdata_d2(sram_rdata_d2), .sram_rdata_d3(
        sram_rdata_d3), .sram_rdata_d4(sram_rdata_d4), .sram_rdata_e0(
        sram_rdata_e0), .sram_rdata_e1(sram_rdata_e1), .sram_rdata_e2(
        sram_rdata_e2), .sram_rdata_e3(sram_rdata_e3), .sram_rdata_e4(
        sram_rdata_e4), .sram_sel(sram_sel), .src_window(src_window) );
  fc_multiplier_accumulator fc_multiplier_accumulator ( .clk(clk), .srstn(
        srstn), .src_window(src_window), .sram_rdata_weight(sram_rdata_weight), 
        .accumulate_reset(accumulate_reset), .data_out({data_out_22_, 
        data_out_21_, data_out_20_, data_out_19_, data_out_18_, data_out_17_, 
        data_out_16_, data_out_15_, data_out_14_, data_out_13_, data_out_12_, 
        data_out_11_, data_out_10_, data_out_9_, data_out_8_, data_out_7_, 
        data_out_6_, data_out_5_, data_out_4_, data_out_3_, data_out_2_, 
        data_out_1_, data_out_0_}) );
  fc_quantize fc_quantize ( .clk(clk), .srstn(srstn), .fc_state(fc_state), 
        .quantized_data(sram_wdata_e), .unquautized_data_22_(data_out_22_), 
        .unquautized_data_21_(data_out_21_), .unquautized_data_20_(
        data_out_20_), .unquautized_data_19_(data_out_19_), 
        .unquautized_data_18_(data_out_18_), .unquautized_data_17_(
        data_out_17_), .unquautized_data_16_(data_out_16_), 
        .unquautized_data_15_(data_out_15_), .unquautized_data_14_(
        data_out_14_), .unquautized_data_13_(data_out_13_), 
        .unquautized_data_12_(data_out_12_), .unquautized_data_11_(
        data_out_11_), .unquautized_data_10_(data_out_10_), 
        .unquautized_data_9_(data_out_9_), .unquautized_data_8_(data_out_8_), 
        .unquautized_data_7_(data_out_7_), .unquautized_data_6_(data_out_6_), 
        .unquautized_data_5_(data_out_5_), .unquautized_data_4_(data_out_4_)
         );
  NBUFFX2_HVT U1 ( .A(sram_wdata_e[1]), .Y(sram_wdata_f[1]) );
  NBUFFX2_HVT U2 ( .A(sram_wdata_e[7]), .Y(sram_wdata_f[7]) );
  NBUFFX2_HVT U3 ( .A(sram_wdata_e[4]), .Y(sram_wdata_f[4]) );
  NBUFFX2_HVT U4 ( .A(sram_wdata_e[6]), .Y(sram_wdata_f[6]) );
  NBUFFX2_HVT U5 ( .A(sram_wdata_e[2]), .Y(sram_wdata_f[2]) );
  NBUFFX2_HVT U6 ( .A(sram_wdata_e[3]), .Y(sram_wdata_f[3]) );
  NBUFFX2_HVT U7 ( .A(sram_wdata_e[0]), .Y(sram_wdata_f[0]) );
  NBUFFX2_HVT U8 ( .A(sram_wdata_e[5]), .Y(sram_wdata_f[5]) );
  NBUFFX2_HVT U9 ( .A(sram_bytemask_e[3]), .Y(sram_bytemask_f[3]) );
  NBUFFX2_HVT U10 ( .A(sram_waddr_e[1]), .Y(sram_waddr_f[1]) );
  NBUFFX2_HVT U11 ( .A(sram_waddr_e[0]), .Y(sram_waddr_f[0]) );
  NBUFFX2_HVT U12 ( .A(sram_bytemask_e[1]), .Y(sram_bytemask_f[1]) );
  NBUFFX2_HVT U13 ( .A(sram_bytemask_e[0]), .Y(sram_bytemask_f[0]) );
  NBUFFX2_HVT U14 ( .A(sram_bytemask_e[2]), .Y(sram_bytemask_f[2]) );
endmodule


module lenet ( clk, srstn, conv_start, fc_done, sram_rdata_a0, sram_rdata_a1, 
        sram_rdata_a2, sram_rdata_a3, sram_rdata_a4, sram_rdata_a5, 
        sram_rdata_a6, sram_rdata_a7, sram_rdata_a8, sram_rdata_b0, 
        sram_rdata_b1, sram_rdata_b2, sram_rdata_b3, sram_rdata_b4, 
        sram_rdata_b5, sram_rdata_b6, sram_rdata_b7, sram_rdata_b8, 
        conv_sram_rdata_weight, conv_sram_raddr_weight, sram_raddr_a0, 
        sram_raddr_a1, sram_raddr_a2, sram_raddr_a3, sram_raddr_a4, 
        sram_raddr_a5, sram_raddr_a6, sram_raddr_a7, sram_raddr_a8, 
        sram_write_enable_b0, sram_write_enable_b1, sram_write_enable_b2, 
        sram_write_enable_b3, sram_write_enable_b4, sram_write_enable_b5, 
        sram_write_enable_b6, sram_write_enable_b7, sram_write_enable_b8, 
        sram_bytemask_b, sram_waddr_b, sram_wdata_b, sram_raddr_b0, 
        sram_raddr_b1, sram_raddr_b2, sram_raddr_b3, sram_raddr_b4, 
        sram_raddr_b5, sram_raddr_b6, sram_raddr_b7, sram_raddr_b8, 
        sram_write_enable_c0, sram_write_enable_c1, sram_write_enable_c2, 
        sram_write_enable_c3, sram_write_enable_c4, sram_bytemask_c, 
        sram_waddr_c, sram_wdata_c, sram_write_enable_d0, sram_write_enable_d1, 
        sram_write_enable_d2, sram_write_enable_d3, sram_write_enable_d4, 
        sram_bytemask_d, sram_waddr_d, sram_wdata_d, conv_done, mem_sel, 
        sram_rdata_c0, sram_rdata_c1, sram_rdata_c2, sram_rdata_c3, 
        sram_rdata_c4, sram_raddr_c0, sram_raddr_c1, sram_raddr_c2, 
        sram_raddr_c3, sram_raddr_c4, sram_rdata_d0, sram_rdata_d1, 
        sram_rdata_d2, sram_rdata_d3, sram_rdata_d4, sram_raddr_d0, 
        sram_raddr_d1, sram_raddr_d2, sram_raddr_d3, sram_raddr_d4, 
        sram_rdata_e0, sram_rdata_e1, sram_rdata_e2, sram_rdata_e3, 
        sram_rdata_e4, sram_raddr_e0, sram_raddr_e1, sram_raddr_e2, 
        sram_raddr_e3, sram_raddr_e4, sram_write_enable_e0, 
        sram_write_enable_e1, sram_write_enable_e2, sram_write_enable_e3, 
        sram_write_enable_e4, sram_bytemask_e, sram_waddr_e, sram_wdata_e, 
        sram_write_enable_f, sram_bytemask_f, sram_waddr_f, sram_wdata_f, 
        fc_sram_rdata_weight, fc_sram_raddr_weight, fc1_done, fc2_done );
  input [31:0] sram_rdata_a0;
  input [31:0] sram_rdata_a1;
  input [31:0] sram_rdata_a2;
  input [31:0] sram_rdata_a3;
  input [31:0] sram_rdata_a4;
  input [31:0] sram_rdata_a5;
  input [31:0] sram_rdata_a6;
  input [31:0] sram_rdata_a7;
  input [31:0] sram_rdata_a8;
  input [31:0] sram_rdata_b0;
  input [31:0] sram_rdata_b1;
  input [31:0] sram_rdata_b2;
  input [31:0] sram_rdata_b3;
  input [31:0] sram_rdata_b4;
  input [31:0] sram_rdata_b5;
  input [31:0] sram_rdata_b6;
  input [31:0] sram_rdata_b7;
  input [31:0] sram_rdata_b8;
  input [99:0] conv_sram_rdata_weight;
  output [16:0] conv_sram_raddr_weight;
  output [9:0] sram_raddr_a0;
  output [9:0] sram_raddr_a1;
  output [9:0] sram_raddr_a2;
  output [9:0] sram_raddr_a3;
  output [9:0] sram_raddr_a4;
  output [9:0] sram_raddr_a5;
  output [9:0] sram_raddr_a6;
  output [9:0] sram_raddr_a7;
  output [9:0] sram_raddr_a8;
  output [3:0] sram_bytemask_b;
  output [9:0] sram_waddr_b;
  output [7:0] sram_wdata_b;
  output [9:0] sram_raddr_b0;
  output [9:0] sram_raddr_b1;
  output [9:0] sram_raddr_b2;
  output [9:0] sram_raddr_b3;
  output [9:0] sram_raddr_b4;
  output [9:0] sram_raddr_b5;
  output [9:0] sram_raddr_b6;
  output [9:0] sram_raddr_b7;
  output [9:0] sram_raddr_b8;
  output [3:0] sram_bytemask_c;
  output [9:0] sram_waddr_c;
  output [7:0] sram_wdata_c;
  output [3:0] sram_bytemask_d;
  output [9:0] sram_waddr_d;
  output [7:0] sram_wdata_d;
  input [31:0] sram_rdata_c0;
  input [31:0] sram_rdata_c1;
  input [31:0] sram_rdata_c2;
  input [31:0] sram_rdata_c3;
  input [31:0] sram_rdata_c4;
  output [5:0] sram_raddr_c0;
  output [5:0] sram_raddr_c1;
  output [5:0] sram_raddr_c2;
  output [5:0] sram_raddr_c3;
  output [5:0] sram_raddr_c4;
  input [31:0] sram_rdata_d0;
  input [31:0] sram_rdata_d1;
  input [31:0] sram_rdata_d2;
  input [31:0] sram_rdata_d3;
  input [31:0] sram_rdata_d4;
  output [5:0] sram_raddr_d0;
  output [5:0] sram_raddr_d1;
  output [5:0] sram_raddr_d2;
  output [5:0] sram_raddr_d3;
  output [5:0] sram_raddr_d4;
  input [31:0] sram_rdata_e0;
  input [31:0] sram_rdata_e1;
  input [31:0] sram_rdata_e2;
  input [31:0] sram_rdata_e3;
  input [31:0] sram_rdata_e4;
  output [4:0] sram_raddr_e0;
  output [4:0] sram_raddr_e1;
  output [4:0] sram_raddr_e2;
  output [4:0] sram_raddr_e3;
  output [4:0] sram_raddr_e4;
  output [3:0] sram_bytemask_e;
  output [4:0] sram_waddr_e;
  output [7:0] sram_wdata_e;
  output [3:0] sram_bytemask_f;
  output [1:0] sram_waddr_f;
  output [7:0] sram_wdata_f;
  input [79:0] fc_sram_rdata_weight;
  output [14:0] fc_sram_raddr_weight;
  input clk, srstn, conv_start, fc_done;
  output sram_write_enable_b0, sram_write_enable_b1, sram_write_enable_b2,
         sram_write_enable_b3, sram_write_enable_b4, sram_write_enable_b5,
         sram_write_enable_b6, sram_write_enable_b7, sram_write_enable_b8,
         sram_write_enable_c0, sram_write_enable_c1, sram_write_enable_c2,
         sram_write_enable_c3, sram_write_enable_c4, sram_write_enable_d0,
         sram_write_enable_d1, sram_write_enable_d2, sram_write_enable_d3,
         sram_write_enable_d4, conv_done, mem_sel, sram_write_enable_e0,
         sram_write_enable_e1, sram_write_enable_e2, sram_write_enable_e3,
         sram_write_enable_e4, sram_write_enable_f, fc1_done, fc2_done;


  conv_top conv_top ( .clk(clk), .srstn(srstn), .conv_start(conv_start), 
        .fc_done(fc2_done), .sram_rdata_a0(sram_rdata_a0), .sram_rdata_a1(
        sram_rdata_a1), .sram_rdata_a2(sram_rdata_a2), .sram_rdata_a3(
        sram_rdata_a3), .sram_rdata_a4(sram_rdata_a4), .sram_rdata_a5(
        sram_rdata_a5), .sram_rdata_a6(sram_rdata_a6), .sram_rdata_a7(
        sram_rdata_a7), .sram_rdata_a8(sram_rdata_a8), .sram_rdata_b0(
        sram_rdata_b0), .sram_rdata_b1(sram_rdata_b1), .sram_rdata_b2(
        sram_rdata_b2), .sram_rdata_b3(sram_rdata_b3), .sram_rdata_b4(
        sram_rdata_b4), .sram_rdata_b5(sram_rdata_b5), .sram_rdata_b6(
        sram_rdata_b6), .sram_rdata_b7(sram_rdata_b7), .sram_rdata_b8(
        sram_rdata_b8), .sram_rdata_weight(conv_sram_rdata_weight), 
        .sram_raddr_weight(conv_sram_raddr_weight), .sram_raddr_a0(
        sram_raddr_a0), .sram_raddr_a1(sram_raddr_a1), .sram_raddr_a2(
        sram_raddr_a2), .sram_raddr_a3(sram_raddr_a3), .sram_raddr_a4(
        sram_raddr_a4), .sram_raddr_a5(sram_raddr_a5), .sram_raddr_a6(
        sram_raddr_a6), .sram_raddr_a7(sram_raddr_a7), .sram_raddr_a8(
        sram_raddr_a8), .sram_write_enable_b0(sram_write_enable_b0), 
        .sram_write_enable_b1(sram_write_enable_b1), .sram_write_enable_b2(
        sram_write_enable_b2), .sram_write_enable_b3(sram_write_enable_b3), 
        .sram_write_enable_b4(sram_write_enable_b4), .sram_write_enable_b5(
        sram_write_enable_b5), .sram_write_enable_b6(sram_write_enable_b6), 
        .sram_write_enable_b7(sram_write_enable_b7), .sram_write_enable_b8(
        sram_write_enable_b8), .sram_bytemask_b(sram_bytemask_b), 
        .sram_waddr_b(sram_waddr_b), .sram_wdata_b(sram_wdata_b), 
        .sram_raddr_b0(sram_raddr_b0), .sram_raddr_b1(sram_raddr_b1), 
        .sram_raddr_b2(sram_raddr_b2), .sram_raddr_b3(sram_raddr_b3), 
        .sram_raddr_b4(sram_raddr_b4), .sram_raddr_b5(sram_raddr_b5), 
        .sram_raddr_b6(sram_raddr_b6), .sram_raddr_b7(sram_raddr_b7), 
        .sram_raddr_b8(sram_raddr_b8), .sram_write_enable_c0(
        sram_write_enable_c0), .sram_write_enable_c1(sram_write_enable_c1), 
        .sram_write_enable_c2(sram_write_enable_c2), .sram_write_enable_c3(
        sram_write_enable_c3), .sram_write_enable_c4(sram_write_enable_c4), 
        .sram_bytemask_c(sram_bytemask_c), .sram_waddr_c(sram_waddr_c), 
        .sram_wdata_c(sram_wdata_c), .sram_write_enable_d0(
        sram_write_enable_d0), .sram_write_enable_d1(sram_write_enable_d1), 
        .sram_write_enable_d2(sram_write_enable_d2), .sram_write_enable_d3(
        sram_write_enable_d3), .sram_write_enable_d4(sram_write_enable_d4), 
        .sram_bytemask_d(sram_bytemask_d), .sram_waddr_d(sram_waddr_d), 
        .sram_wdata_d(sram_wdata_d), .conv_done(conv_done), .mem_sel(mem_sel)
         );
  fc_top fc_top ( .clk(clk), .srstn(srstn), .conv_done(conv_done), .mem_sel(
        mem_sel), .sram_rdata_c0(sram_rdata_c0), .sram_rdata_c1(sram_rdata_c1), 
        .sram_rdata_c2(sram_rdata_c2), .sram_rdata_c3(sram_rdata_c3), 
        .sram_rdata_c4(sram_rdata_c4), .sram_raddr_c0(sram_raddr_c0), 
        .sram_raddr_c1(sram_raddr_c1), .sram_raddr_c2(sram_raddr_c2), 
        .sram_raddr_c3(sram_raddr_c3), .sram_raddr_c4(sram_raddr_c4), 
        .sram_rdata_d0(sram_rdata_d0), .sram_rdata_d1(sram_rdata_d1), 
        .sram_rdata_d2(sram_rdata_d2), .sram_rdata_d3(sram_rdata_d3), 
        .sram_rdata_d4(sram_rdata_d4), .sram_raddr_d0(sram_raddr_d0), 
        .sram_raddr_d1(sram_raddr_d1), .sram_raddr_d2(sram_raddr_d2), 
        .sram_raddr_d3(sram_raddr_d3), .sram_raddr_d4(sram_raddr_d4), 
        .sram_rdata_e0(sram_rdata_e0), .sram_rdata_e1(sram_rdata_e1), 
        .sram_rdata_e2(sram_rdata_e2), .sram_rdata_e3(sram_rdata_e3), 
        .sram_rdata_e4(sram_rdata_e4), .sram_raddr_e0(sram_raddr_e0), 
        .sram_raddr_e1(sram_raddr_e1), .sram_raddr_e2(sram_raddr_e2), 
        .sram_raddr_e3(sram_raddr_e3), .sram_raddr_e4(sram_raddr_e4), 
        .sram_write_enable_e0(sram_write_enable_e0), .sram_write_enable_e1(
        sram_write_enable_e1), .sram_write_enable_e2(sram_write_enable_e2), 
        .sram_write_enable_e3(sram_write_enable_e3), .sram_write_enable_e4(
        sram_write_enable_e4), .sram_bytemask_e(sram_bytemask_e), 
        .sram_waddr_e(sram_waddr_e), .sram_wdata_e(sram_wdata_e), 
        .sram_write_enable_f(sram_write_enable_f), .sram_bytemask_f(
        sram_bytemask_f), .sram_waddr_f(sram_waddr_f), .sram_wdata_f(
        sram_wdata_f), .sram_rdata_weight(fc_sram_rdata_weight), 
        .sram_raddr_weight(fc_sram_raddr_weight), .fc1_done(fc1_done), 
        .fc2_done(fc2_done) );
endmodule

