
module fsm ( clk, srstn, conv_start, conv1_done, conv_done, fc_done, mode, 
        mem_sel );
  output [1:0] mode;
  input clk, srstn, conv_start, conv1_done, conv_done, fc_done;
  output mem_sel;
  wire   n_mem_sel, done_control, n2, n6, n8, n3, n5, n7, n9, n10, n11, n13,
         n14, n15, n16;
  wire   [1:0] n_mode;

  DFFSSRX1_HVT mode_reg_1_ ( .D(1'b0), .SETB(n8), .RSTB(n_mode[1]), .CLK(clk), 
        .Q(mode[1]), .QN(n11) );
  DFFSSRX1_HVT done_control_reg ( .D(done_control), .SETB(n2), .RSTB(srstn), 
        .CLK(clk), .Q(done_control), .QN(n10) );
  DFFSSRX1_HVT mem_sel_reg ( .D(n_mem_sel), .SETB(srstn), .RSTB(1'b1), .CLK(
        clk), .Q(mem_sel) );
  DFFSSRX2_HVT mode_reg_0_ ( .D(1'b0), .SETB(n8), .RSTB(n_mode[0]), .CLK(clk), 
        .Q(n5), .QN(n6) );
  OR2X1_HVT U4 ( .A1(n15), .A2(n3), .Y(n_mode[1]) );
  AND3X2_HVT U5 ( .A1(n11), .A2(conv1_done), .A3(mode[0]), .Y(n3) );
  INVX4_HVT U6 ( .A(n6), .Y(mode[0]) );
  INVX0_HVT U7 ( .A(srstn), .Y(n8) );
  INVX0_HVT U8 ( .A(conv_done), .Y(n2) );
  INVX1_HVT U9 ( .A(n5), .Y(n7) );
  AND2X1_HVT U10 ( .A1(n9), .A2(n7), .Y(n15) );
  INVX1_HVT U11 ( .A(n11), .Y(n9) );
  INVX1_HVT U12 ( .A(conv1_done), .Y(n13) );
  MUX21X1_HVT U13 ( .A1(n13), .A2(conv_start), .S0(n7), .Y(n14) );
  AO22X1_HVT U14 ( .A1(n15), .A2(conv_done), .A3(n14), .A4(n11), .Y(n_mode[0])
         );
  AO22X1_HVT U15 ( .A1(done_control), .A2(fc_done), .A3(n10), .A4(conv_done), 
        .Y(n16) );
  HADDX1_HVT U16 ( .A0(mem_sel), .B0(n16), .SO(n_mem_sel) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_0 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n1;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n1), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n1) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_26 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_25 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_24 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_23 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_22 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_21 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_20 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_19 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_18 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_17 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_16 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_15 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_14 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_13 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_12 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_11 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_10 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_9 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_8 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_7 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_6 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_5 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_4 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_3 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_2 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_1 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22627, n2;

  AND2X1_HVT main_gate ( .A1(net22627), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22627) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module conv_control ( clk, srstn, mode, mem_sel, conv1_done, sram_raddr_weight, 
        box_sel, load_conv1_bias_enable, conv1_bias_set, sram_raddr_a0, 
        sram_raddr_a1, sram_raddr_a2, sram_raddr_a3, sram_raddr_a4, 
        sram_raddr_a5, sram_raddr_a6, sram_raddr_a7, sram_raddr_a8, 
        sram_write_enable_b0, sram_write_enable_b1, sram_write_enable_b2, 
        sram_write_enable_b3, sram_write_enable_b4, sram_write_enable_b5, 
        sram_write_enable_b6, sram_write_enable_b7, sram_write_enable_b8, 
        sram_bytemask_b, sram_waddr_b, conv_done, channel, set, 
        load_conv2_bias0_enable, load_conv2_bias1_enable, sram_raddr_b0, 
        sram_raddr_b1, sram_raddr_b2, sram_raddr_b3, sram_raddr_b4, 
        sram_raddr_b5, sram_raddr_b6, sram_raddr_b7, sram_raddr_b8, 
        sram_write_enable_c0, sram_write_enable_c1, sram_write_enable_c2, 
        sram_write_enable_c3, sram_write_enable_c4, sram_bytemask_c, 
        sram_waddr_c, sram_write_enable_d0, sram_write_enable_d1, 
        sram_write_enable_d2, sram_write_enable_d3, sram_write_enable_d4, 
        sram_bytemask_d, sram_waddr_d );
  input [1:0] mode;
  output [16:0] sram_raddr_weight;
  output [3:0] box_sel;
  output [16:0] conv1_bias_set;
  output [9:0] sram_raddr_a0;
  output [9:0] sram_raddr_a1;
  output [9:0] sram_raddr_a2;
  output [9:0] sram_raddr_a3;
  output [9:0] sram_raddr_a4;
  output [9:0] sram_raddr_a5;
  output [9:0] sram_raddr_a6;
  output [9:0] sram_raddr_a7;
  output [9:0] sram_raddr_a8;
  output [3:0] sram_bytemask_b;
  output [9:0] sram_waddr_b;
  output [4:0] channel;
  output [7:0] set;
  output [9:0] sram_raddr_b0;
  output [9:0] sram_raddr_b1;
  output [9:0] sram_raddr_b2;
  output [9:0] sram_raddr_b3;
  output [9:0] sram_raddr_b4;
  output [9:0] sram_raddr_b5;
  output [9:0] sram_raddr_b6;
  output [9:0] sram_raddr_b7;
  output [9:0] sram_raddr_b8;
  output [3:0] sram_bytemask_c;
  output [9:0] sram_waddr_c;
  output [3:0] sram_bytemask_d;
  output [9:0] sram_waddr_d;
  input clk, srstn, mem_sel;
  output conv1_done, load_conv1_bias_enable, sram_write_enable_b0,
         sram_write_enable_b1, sram_write_enable_b2, sram_write_enable_b3,
         sram_write_enable_b4, sram_write_enable_b5, sram_write_enable_b6,
         sram_write_enable_b7, sram_write_enable_b8, conv_done,
         load_conv2_bias0_enable, load_conv2_bias1_enable,
         sram_write_enable_c0, sram_write_enable_c1, sram_write_enable_c2,
         sram_write_enable_c3, sram_write_enable_c4, sram_write_enable_d0,
         sram_write_enable_d1, sram_write_enable_d2, sram_write_enable_d3,
         sram_write_enable_d4;
  wire   n_conv1_done, n_conv_done, conv1_weight_done, conv2_weight_done,
         delay3_write_enable, load_data_enable, n_conv1_weight_done,
         n_write_enable, write_enable, delay_write_enable, delay2_write_enable,
         n_load_data_enable, n_box_sel_1_, n_addr_row_sel_cnt_0_,
         n_sram_write_enable_b0, n_sram_write_enable_b1,
         n_sram_write_enable_b2, n_sram_write_enable_b3,
         n_sram_write_enable_b4, n_sram_write_enable_b5,
         n_sram_write_enable_b6, n_sram_write_enable_b7,
         n_sram_write_enable_b8, n_sram_write_enable_c0,
         n_sram_write_enable_c1, n_sram_write_enable_c2,
         n_sram_write_enable_c3, n_sram_write_enable_c4,
         n_sram_write_enable_d0, n_sram_write_enable_d1,
         n_sram_write_enable_d2, n_sram_write_enable_d3,
         n_sram_write_enable_d4, N2914, net22461, net22638, net22643, net22648,
         net22653, net22654, net22657, net22662, net22691, net22698, net22705,
         net22712, net22719, net22726, net22733, net22747, net22754, net22757,
         net22775, net22782, net22789, net22796, net22810, net22817, net22824,
         net22838, net22852, net22855, net22860, net22863, net22866, net22869,
         net22872, net22875, net22878, net22881, net22884, net22887, net22890,
         net22893, net22898, net22900, net22901, net22902, net22903, net22904,
         net22905, net22906, net22907, net22908, net22909, net22912, net22916,
         net22917, net22918, net22919, net22920, net22921, net22922, net22923,
         net22924, net22925, net22928, net22932, net22933, net22934, net22935,
         net22936, net22937, net22940, net22943, net22945, net22946, net22947,
         net22948, net22949, net22952, net23433, net23878, net23892, net24315,
         net24760, net25205, net25219, net25642, net26088, net26534, net26549,
         net26972, net27506, net28021, net28536, net29051, net29566, net30081,
         net30596, net31111, net31203, net31626, n368, n369, n371, n392, n1020,
         n1021, n1022, n1023, n1024, n1027, n1051, n1052, n1053, n1061, n1062,
         n1063, n1070, n1655, n1662, n1667, n1, n2, n3, n4, n5, n6, n8, n9,
         n10, n12, n13, n14, n15, n17, n18, n21, n22, n23, n25, n26, n27, n28,
         n30, n31, n32, n33, n34, n35, n36, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n55, n56, n57, n58, n59, n60, n61, n66, n67, n68,
         n69, n70, n71, n72, n73, n75, n77, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n91, n92, n93, n95, n97, n98, n99, n101, n103,
         n104, n107, n108, n110, n112, n114, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n134, n137, n138, n139, n140, n143, n145, n146, n147, n148,
         n149, n150, n152, n153, n156, n158, n159, n160, n161, n163, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n370, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1025, n1026, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1064, n1065, n1066, n1067, n1068, n1069,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1656, n1657, n1658, n1659, n1660, n1661,
         n1663, n1664, n1665, n1666, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004;
  wire   [7:0] conv1_weight_cnt;
  wire   [7:0] conv2_weight_cnt;
  wire   [3:0] state;
  wire   [3:0] n_state;
  wire   [4:0] channel_cnt;
  wire   [1:0] data_sel_col;
  wire   [1:0] data_sel_row;
  wire   [9:0] delay1_sram_waddr_b;
  wire   [3:0] write_row_conv1;
  wire   [1:0] write_col_conv1;
  wire   [4:0] delay3_addr_change;
  wire   [2:0] delay3_state;
  wire   [3:0] n_row;
  wire   [7:0] n_weight_cnt;
  wire   [7:0] weight_cnt;
  wire   [7:0] delay_set;
  wire   [1:0] n_addr_col_sel_cnt;
  wire   [1:0] addr_col_sel_cnt;
  wire   [1:0] addr_row_sel_cnt;
  wire   [3:0] n_sram_bytemask_b;
  wire   [3:0] row;
  wire   [3:0] col;
  wire   [3:0] row_delay;
  wire   [3:0] col_delay;
  wire   [3:0] write_row;
  wire   [3:0] write_col;
  wire   [3:0] row_enable;
  wire   [3:0] col_enable;
  wire   [9:0] delay1_sram_waddr_c;
  wire   [9:0] delay1_sram_waddr_d;
  wire   [3:0] n_sram_bytemask_c;
  wire   [3:0] n_sram_bytemask_d;
  wire   [4:0] addr_change;
  wire   [4:0] delay_addr_change;
  wire   [4:0] delay2_addr_change;
  wire   [4:0] delay_channel;
  wire   [4:0] delay2_channel;
  wire   [3:0] delay1_state;
  wire   [3:0] delay2_state;
  wire   [9:0] n_sram_raddr_a0;
  wire   [9:0] n_sram_raddr_a1;
  wire   [9:0] n_sram_raddr_a2;
  wire   [9:0] n_sram_raddr_a3;
  wire   [9:0] n_sram_raddr_a4;
  wire   [9:0] n_sram_raddr_a5;
  wire   [9:0] n_sram_raddr_a6;
  wire   [9:0] n_sram_raddr_a7;
  wire   [9:0] n_sram_raddr_a8;
  wire   [9:0] n_sram_raddr_b0;
  wire   [9:0] n_sram_raddr_b1;
  wire   [9:0] n_sram_raddr_b2;
  wire   [9:0] n_sram_raddr_b3;
  wire   [9:0] n_sram_raddr_b4;
  wire   [9:0] n_sram_raddr_b5;
  wire   [9:0] n_sram_raddr_b6;
  wire   [9:0] n_sram_raddr_b7;
  wire   [9:0] n_sram_raddr_b8;

  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_0 clk_gate_col_reg ( .CLK(clk), 
        .EN(net22461), .ENCLK(net22657) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_26 clk_gate_weight_cnt_reg ( 
        .CLK(clk), .EN(net22461), .ENCLK(net22662) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_25 clk_gate_sram_raddr_weight_reg ( 
        .CLK(clk), .EN(net22775), .ENCLK(net22757) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_24 clk_gate_sram_raddr_weight_reg_0 ( 
        .CLK(clk), .EN(net22775), .ENCLK(net22855) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_23 clk_gate_delay1_sram_waddr_b_reg ( 
        .CLK(clk), .EN(net22860), .ENCLK(net22893) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_22 clk_gate_delay1_sram_waddr_c_reg ( 
        .CLK(clk), .EN(net22898), .ENCLK(net22912) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_21 clk_gate_delay1_sram_waddr_d_reg ( 
        .CLK(clk), .EN(net22898), .ENCLK(net22928) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_20 clk_gate_channel_cnt_reg ( 
        .CLK(clk), .EN(net22932), .ENCLK(net22940) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_19 clk_gate_addr_change_reg ( 
        .CLK(clk), .EN(net22943), .ENCLK(net22952) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_18 clk_gate_sram_raddr_a7_reg ( 
        .CLK(clk), .EN(net23892), .ENCLK(net23433) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_17 clk_gate_sram_raddr_a1_reg ( 
        .CLK(clk), .EN(net23892), .ENCLK(net23878) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_16 clk_gate_sram_raddr_a4_reg ( 
        .CLK(clk), .EN(net23892), .ENCLK(net24315) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_15 clk_gate_sram_raddr_a8_reg ( 
        .CLK(clk), .EN(net25219), .ENCLK(net24760) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_14 clk_gate_sram_raddr_a2_reg ( 
        .CLK(clk), .EN(net25219), .ENCLK(net25205) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_13 clk_gate_sram_raddr_a5_reg ( 
        .CLK(clk), .EN(net25219), .ENCLK(net25642) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_12 clk_gate_sram_raddr_a0_reg ( 
        .CLK(clk), .EN(net26549), .ENCLK(net26088) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_11 clk_gate_sram_raddr_a3_reg ( 
        .CLK(clk), .EN(net26549), .ENCLK(net26534) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_10 clk_gate_sram_raddr_a6_reg ( 
        .CLK(clk), .EN(net26549), .ENCLK(net26972) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_9 clk_gate_sram_raddr_b7_reg ( 
        .CLK(clk), .EN(net31203), .ENCLK(net27506) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_8 clk_gate_sram_raddr_b8_reg ( 
        .CLK(clk), .EN(net31203), .ENCLK(net28021) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_7 clk_gate_sram_raddr_b0_reg ( 
        .CLK(clk), .EN(net31203), .ENCLK(net28536) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_6 clk_gate_sram_raddr_b1_reg ( 
        .CLK(clk), .EN(net31203), .ENCLK(net29051) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_5 clk_gate_sram_raddr_b2_reg ( 
        .CLK(clk), .EN(net31203), .ENCLK(net29566) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_4 clk_gate_sram_raddr_b3_reg ( 
        .CLK(clk), .EN(net31203), .ENCLK(net30081) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_3 clk_gate_sram_raddr_b4_reg ( 
        .CLK(clk), .EN(net31203), .ENCLK(net30596) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_2 clk_gate_sram_raddr_b5_reg ( 
        .CLK(clk), .EN(net31203), .ENCLK(net31111) );
  SNPS_CLOCK_GATE_HIGH_conv_control_mydesign_1 clk_gate_sram_raddr_b6_reg ( 
        .CLK(clk), .EN(net31203), .ENCLK(net31626) );
  DFFSSRX1_HVT channel_cnt_reg_0_ ( .D(1'b0), .SETB(n197), .RSTB(net22937), 
        .CLK(net22940), .Q(channel_cnt[0]) );
  DFFSSRX1_HVT state_reg_0_ ( .D(1'b0), .SETB(n193), .RSTB(n_state[0]), .CLK(
        clk), .Q(state[0]), .QN(n310) );
  DFFSSRX1_HVT weight_cnt_reg_0_ ( .D(1'b0), .SETB(n199), .RSTB(
        n_weight_cnt[0]), .CLK(net22662), .Q(weight_cnt[0]), .QN(n299) );
  DFFSSRX1_HVT delay_set_reg_0_ ( .D(1'b0), .SETB(n195), .RSTB(weight_cnt[0]), 
        .CLK(clk), .Q(delay_set[0]) );
  DFFSSRX1_HVT set_reg_0_ ( .D(1'b0), .SETB(n229), .RSTB(delay_set[0]), .CLK(
        clk), .Q(set[0]) );
  DFFSSRX1_HVT conv2_weight_cnt_reg_0_ ( .D(1'b0), .SETB(n208), .RSTB(set[0]), 
        .CLK(clk), .Q(conv2_weight_cnt[0]) );
  DFFSSRX1_HVT conv1_weight_cnt_reg_0_ ( .D(1'b0), .SETB(n186), .RSTB(
        conv2_weight_cnt[0]), .CLK(clk), .Q(conv1_weight_cnt[0]) );
  DFFSSRX1_HVT conv_done_reg ( .D(1'b0), .SETB(n183), .RSTB(n_conv_done), 
        .CLK(clk), .Q(conv_done) );
  DFFSSRX1_HVT state_reg_1_ ( .D(1'b0), .SETB(n198), .RSTB(n_state[1]), .CLK(
        clk), .Q(state[1]), .QN(n251) );
  DFFSSRX1_HVT weight_cnt_reg_7_ ( .D(1'b0), .SETB(n194), .RSTB(
        n_weight_cnt[7]), .CLK(net22662), .Q(weight_cnt[7]), .QN(n448) );
  DFFSSRX1_HVT delay_set_reg_7_ ( .D(1'b0), .SETB(n200), .RSTB(weight_cnt[7]), 
        .CLK(clk), .Q(delay_set[7]) );
  DFFSSRX1_HVT set_reg_7_ ( .D(1'b0), .SETB(n196), .RSTB(delay_set[7]), .CLK(
        clk), .Q(set[7]) );
  DFFSSRX1_HVT conv2_weight_cnt_reg_7_ ( .D(1'b0), .SETB(n186), .RSTB(set[7]), 
        .CLK(clk), .Q(conv2_weight_cnt[7]) );
  DFFSSRX1_HVT conv1_weight_cnt_reg_7_ ( .D(1'b0), .SETB(n207), .RSTB(
        conv2_weight_cnt[7]), .CLK(clk), .Q(conv1_weight_cnt[7]) );
  DFFSSRX1_HVT weight_cnt_reg_6_ ( .D(1'b0), .SETB(n185), .RSTB(
        n_weight_cnt[6]), .CLK(net22662), .Q(weight_cnt[6]) );
  DFFSSRX1_HVT delay_set_reg_6_ ( .D(1'b0), .SETB(n182), .RSTB(weight_cnt[6]), 
        .CLK(clk), .Q(delay_set[6]) );
  DFFSSRX1_HVT set_reg_6_ ( .D(1'b0), .SETB(n175), .RSTB(delay_set[6]), .CLK(
        clk), .Q(set[6]) );
  DFFSSRX1_HVT conv2_weight_cnt_reg_6_ ( .D(1'b0), .SETB(n177), .RSTB(set[6]), 
        .CLK(clk), .Q(conv2_weight_cnt[6]) );
  DFFSSRX1_HVT conv1_weight_cnt_reg_6_ ( .D(1'b0), .SETB(n176), .RSTB(
        conv2_weight_cnt[6]), .CLK(clk), .Q(conv1_weight_cnt[6]) );
  DFFSSRX1_HVT weight_cnt_reg_5_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_weight_cnt[5]), .CLK(net22662), .Q(weight_cnt[5]), .QN(n439) );
  DFFSSRX1_HVT delay_set_reg_5_ ( .D(1'b0), .SETB(n182), .RSTB(weight_cnt[5]), 
        .CLK(clk), .Q(delay_set[5]) );
  DFFSSRX1_HVT set_reg_5_ ( .D(1'b0), .SETB(n208), .RSTB(delay_set[5]), .CLK(
        clk), .Q(set[5]) );
  DFFSSRX1_HVT conv2_weight_cnt_reg_5_ ( .D(1'b0), .SETB(n187), .RSTB(set[5]), 
        .CLK(clk), .Q(conv2_weight_cnt[5]) );
  DFFSSRX1_HVT conv1_weight_cnt_reg_5_ ( .D(1'b0), .SETB(n184), .RSTB(
        conv2_weight_cnt[5]), .CLK(clk), .Q(conv1_weight_cnt[5]) );
  DFFSSRX1_HVT weight_cnt_reg_4_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_weight_cnt[4]), .CLK(net22662), .Q(weight_cnt[4]) );
  DFFSSRX1_HVT delay_set_reg_4_ ( .D(1'b0), .SETB(n177), .RSTB(weight_cnt[4]), 
        .CLK(clk), .Q(delay_set[4]) );
  DFFSSRX1_HVT set_reg_4_ ( .D(1'b0), .SETB(n176), .RSTB(delay_set[4]), .CLK(
        clk), .Q(set[4]) );
  DFFSSRX1_HVT conv2_weight_cnt_reg_4_ ( .D(1'b0), .SETB(n174), .RSTB(set[4]), 
        .CLK(clk), .Q(conv2_weight_cnt[4]) );
  DFFSSRX1_HVT conv1_weight_cnt_reg_4_ ( .D(1'b0), .SETB(n187), .RSTB(
        conv2_weight_cnt[4]), .CLK(clk), .Q(conv1_weight_cnt[4]) );
  DFFSSRX1_HVT weight_cnt_reg_3_ ( .D(1'b0), .SETB(n207), .RSTB(
        n_weight_cnt[3]), .CLK(net22662), .Q(weight_cnt[3]), .QN(n424) );
  DFFSSRX1_HVT delay_set_reg_3_ ( .D(1'b0), .SETB(n186), .RSTB(weight_cnt[3]), 
        .CLK(clk), .Q(delay_set[3]) );
  DFFSSRX1_HVT set_reg_3_ ( .D(1'b0), .SETB(n183), .RSTB(delay_set[3]), .CLK(
        clk), .Q(set[3]) );
  DFFSSRX1_HVT conv2_weight_cnt_reg_3_ ( .D(1'b0), .SETB(n197), .RSTB(set[3]), 
        .CLK(clk), .Q(conv2_weight_cnt[3]) );
  DFFSSRX1_HVT conv1_weight_cnt_reg_3_ ( .D(1'b0), .SETB(n193), .RSTB(
        conv2_weight_cnt[3]), .CLK(clk), .Q(conv1_weight_cnt[3]) );
  DFFSSRX1_HVT weight_cnt_reg_2_ ( .D(1'b0), .SETB(n199), .RSTB(
        n_weight_cnt[2]), .CLK(net22662), .Q(weight_cnt[2]) );
  DFFSSRX1_HVT delay_set_reg_2_ ( .D(1'b0), .SETB(n195), .RSTB(weight_cnt[2]), 
        .CLK(clk), .Q(delay_set[2]) );
  DFFSSRX1_HVT set_reg_2_ ( .D(1'b0), .SETB(n184), .RSTB(delay_set[2]), .CLK(
        clk), .Q(set[2]) );
  DFFSSRX1_HVT conv2_weight_cnt_reg_2_ ( .D(1'b0), .SETB(n208), .RSTB(set[2]), 
        .CLK(clk), .Q(conv2_weight_cnt[2]) );
  DFFSSRX1_HVT conv1_weight_cnt_reg_2_ ( .D(1'b0), .SETB(n185), .RSTB(
        conv2_weight_cnt[2]), .CLK(clk), .Q(conv1_weight_cnt[2]) );
  DFFSSRX1_HVT weight_cnt_reg_1_ ( .D(1'b0), .SETB(n182), .RSTB(
        n_weight_cnt[1]), .CLK(net22662), .Q(weight_cnt[1]), .QN(n430) );
  DFFSSRX1_HVT delay_set_reg_1_ ( .D(1'b0), .SETB(n198), .RSTB(weight_cnt[1]), 
        .CLK(clk), .Q(delay_set[1]) );
  DFFSSRX1_HVT set_reg_1_ ( .D(1'b0), .SETB(n194), .RSTB(delay_set[1]), .CLK(
        clk), .Q(set[1]) );
  DFFSSRX1_HVT conv2_weight_cnt_reg_1_ ( .D(1'b0), .SETB(n200), .RSTB(set[1]), 
        .CLK(clk), .Q(conv2_weight_cnt[1]) );
  DFFSSRX1_HVT conv1_weight_cnt_reg_1_ ( .D(1'b0), .SETB(n196), .RSTB(
        conv2_weight_cnt[1]), .CLK(clk), .Q(conv1_weight_cnt[1]) );
  DFFSSRX1_HVT conv1_done_reg ( .D(1'b0), .SETB(n186), .RSTB(n_conv1_done), 
        .CLK(clk), .Q(conv1_done), .QN(n449) );
  DFFSSRX1_HVT col_reg_0_ ( .D(1'b0), .SETB(n207), .RSTB(net22653), .CLK(
        net22657), .Q(col[0]), .QN(n254) );
  DFFSSRX1_HVT col_delay_reg_0_ ( .D(1'b0), .SETB(n187), .RSTB(col[0]), .CLK(
        clk), .Q(col_delay[0]) );
  DFFSSRX1_HVT write_col_reg_0_ ( .D(1'b0), .SETB(n184), .RSTB(col_delay[0]), 
        .CLK(clk), .Q(write_col[0]) );
  DFFSSRX1_HVT col_enable_reg_0_ ( .D(1'b0), .SETB(n175), .RSTB(write_col[0]), 
        .CLK(clk), .Q(col_enable[0]) );
  DFFSSRX1_HVT write_col_conv1_reg_0_ ( .D(1'b0), .SETB(n177), .RSTB(
        col_enable[0]), .CLK(clk), .Q(write_col_conv1[0]) );
  DFFSSRX1_HVT col_reg_1_ ( .D(1'b0), .SETB(n176), .RSTB(net22648), .CLK(
        net22657), .Q(col[1]), .QN(n312) );
  DFFSSRX1_HVT col_delay_reg_1_ ( .D(1'b0), .SETB(n174), .RSTB(col[1]), .CLK(
        clk), .Q(col_delay[1]) );
  DFFSSRX1_HVT write_col_reg_1_ ( .D(1'b0), .SETB(n183), .RSTB(col_delay[1]), 
        .CLK(clk), .Q(write_col[1]) );
  DFFSSRX1_HVT col_enable_reg_1_ ( .D(1'b0), .SETB(n208), .RSTB(write_col[1]), 
        .CLK(clk), .Q(col_enable[1]) );
  DFFSSRX1_HVT write_col_conv1_reg_1_ ( .D(1'b0), .SETB(n186), .RSTB(
        col_enable[1]), .CLK(clk), .Q(write_col_conv1[1]), .QN(n320) );
  DFFSSRX1_HVT col_reg_2_ ( .D(1'b0), .SETB(n183), .RSTB(net22643), .CLK(
        net22657), .Q(col[2]), .QN(n233) );
  DFFSSRX1_HVT col_delay_reg_2_ ( .D(1'b0), .SETB(n175), .RSTB(col[2]), .CLK(
        clk), .Q(col_delay[2]) );
  DFFSSRX1_HVT write_col_reg_2_ ( .D(1'b0), .SETB(n177), .RSTB(col_delay[2]), 
        .CLK(clk), .Q(write_col[2]) );
  DFFSSRX1_HVT col_enable_reg_2_ ( .D(1'b0), .SETB(n176), .RSTB(write_col[2]), 
        .CLK(clk), .Q(col_enable[2]) );
  DFFSSRX1_HVT write_col_conv1_reg_2_ ( .D(1'b0), .SETB(n174), .RSTB(
        col_enable[2]), .CLK(clk), .Q(n261), .QN(n1063) );
  DFFSSRX1_HVT col_reg_3_ ( .D(1'b0), .SETB(n200), .RSTB(net22638), .CLK(
        net22657), .Q(col[3]), .QN(n238) );
  DFFSSRX1_HVT col_delay_reg_3_ ( .D(1'b0), .SETB(n207), .RSTB(col[3]), .CLK(
        clk), .Q(col_delay[3]) );
  DFFSSRX1_HVT write_col_reg_3_ ( .D(1'b0), .SETB(n185), .RSTB(col_delay[3]), 
        .CLK(clk), .Q(write_col[3]) );
  DFFSSRX1_HVT col_enable_reg_3_ ( .D(1'b0), .SETB(n182), .RSTB(write_col[3]), 
        .CLK(clk), .Q(col_enable[3]) );
  DFFSSRX1_HVT write_col_conv1_reg_3_ ( .D(1'b0), .SETB(n197), .RSTB(
        col_enable[3]), .CLK(clk), .Q(n262), .QN(n1062) );
  DFFSSRX1_HVT addr_col_sel_cnt_reg_0_ ( .D(1'b0), .SETB(n193), .RSTB(
        n_addr_col_sel_cnt[0]), .CLK(clk), .Q(addr_col_sel_cnt[0]), .QN(n1052)
         );
  DFFSSRX1_HVT data_sel_col_reg_0_ ( .D(1'b0), .SETB(n199), .RSTB(
        addr_col_sel_cnt[0]), .CLK(clk), .Q(data_sel_col[0]) );
  DFFSSRX1_HVT addr_col_sel_cnt_reg_1_ ( .D(1'b0), .SETB(n195), .RSTB(
        n_addr_col_sel_cnt[1]), .CLK(clk), .Q(addr_col_sel_cnt[1]), .QN(n1051)
         );
  DFFSSRX1_HVT data_sel_col_reg_1_ ( .D(1'b0), .SETB(n229), .RSTB(
        addr_col_sel_cnt[1]), .CLK(clk), .Q(data_sel_col[1]) );
  DFFSSRX1_HVT addr_row_sel_cnt_reg_0_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_addr_row_sel_cnt_0_), .CLK(clk), .Q(addr_row_sel_cnt[0]), .QN(n317)
         );
  DFFSSRX1_HVT data_sel_row_reg_0_ ( .D(1'b0), .SETB(n187), .RSTB(
        addr_row_sel_cnt[0]), .CLK(clk), .Q(data_sel_row[0]) );
  DFFSSRX1_HVT addr_row_sel_cnt_reg_1_ ( .D(n392), .SETB(n1667), .RSTB(n181), 
        .CLK(clk), .Q(addr_row_sel_cnt[1]), .QN(n1053) );
  DFFSSRX1_HVT data_sel_row_reg_1_ ( .D(1'b0), .SETB(n184), .RSTB(
        addr_row_sel_cnt[1]), .CLK(clk), .Q(data_sel_row[1]) );
  DFFSSRX1_HVT conv2_weight_done_reg ( .D(1'b0), .SETB(n198), .RSTB(net22654), 
        .CLK(net22657), .Q(conv2_weight_done) );
  DFFSSRX1_HVT row_reg_0_ ( .D(1'b0), .SETB(n194), .RSTB(n_row[0]), .CLK(
        net22657), .Q(row[0]), .QN(n253) );
  DFFSSRX1_HVT row_delay_reg_0_ ( .D(1'b0), .SETB(n200), .RSTB(row[0]), .CLK(
        clk), .Q(row_delay[0]) );
  DFFSSRX1_HVT write_row_reg_0_ ( .D(1'b0), .SETB(n196), .RSTB(row_delay[0]), 
        .CLK(clk), .Q(write_row[0]) );
  DFFSSRX1_HVT row_enable_reg_0_ ( .D(1'b0), .SETB(n199), .RSTB(write_row[0]), 
        .CLK(clk), .Q(row_enable[0]) );
  DFFSSRX1_HVT write_row_conv1_reg_0_ ( .D(1'b0), .SETB(n207), .RSTB(
        row_enable[0]), .CLK(clk), .Q(write_row_conv1[0]) );
  DFFSSRX1_HVT sram_bytemask_d_reg_1_ ( .D(1'b0), .SETB(n186), .RSTB(
        n_sram_bytemask_d[1]), .CLK(clk), .Q(sram_bytemask_d[1]) );
  DFFSSRX1_HVT sram_bytemask_c_reg_1_ ( .D(1'b0), .SETB(n183), .RSTB(
        n_sram_bytemask_c[1]), .CLK(clk), .Q(sram_bytemask_c[1]) );
  DFFSSRX1_HVT sram_bytemask_d_reg_0_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_bytemask_d[0]), .CLK(clk), .Q(sram_bytemask_d[0]) );
  DFFSSRX1_HVT sram_bytemask_c_reg_0_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_bytemask_c[0]), .CLK(clk), .Q(sram_bytemask_c[0]) );
  DFFSSRX1_HVT sram_bytemask_c_reg_2_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_bytemask_c[2]), .CLK(clk), .Q(sram_bytemask_c[2]) );
  DFFSSRX1_HVT sram_bytemask_c_reg_3_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_bytemask_c[3]), .CLK(clk), .Q(sram_bytemask_c[3]) );
  DFFSSRX1_HVT sram_bytemask_d_reg_2_ ( .D(1'b0), .SETB(n207), .RSTB(
        n_sram_bytemask_d[2]), .CLK(clk), .Q(sram_bytemask_d[2]) );
  DFFSSRX1_HVT sram_bytemask_d_reg_3_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_bytemask_d[3]), .CLK(clk), .Q(sram_bytemask_d[3]) );
  DFFSSRX1_HVT row_reg_1_ ( .D(1'b0), .SETB(n185), .RSTB(n_row[1]), .CLK(
        net22657), .Q(row[1]), .QN(n319) );
  DFFSSRX1_HVT row_delay_reg_1_ ( .D(1'b0), .SETB(n182), .RSTB(row[1]), .CLK(
        clk), .Q(row_delay[1]) );
  DFFSSRX1_HVT write_row_reg_1_ ( .D(1'b0), .SETB(n175), .RSTB(row_delay[1]), 
        .CLK(clk), .Q(write_row[1]) );
  DFFSSRX1_HVT row_enable_reg_1_ ( .D(1'b0), .SETB(n177), .RSTB(write_row[1]), 
        .CLK(clk), .Q(row_enable[1]) );
  DFFSSRX1_HVT write_row_conv1_reg_1_ ( .D(1'b0), .SETB(n176), .RSTB(
        row_enable[1]), .CLK(clk), .Q(n249), .QN(n1061) );
  DFFSSRX1_HVT box_sel_reg_2_ ( .D(n371), .SETB(n1655), .RSTB(n181), .CLK(clk), 
        .Q(box_sel[2]) );
  DFFSSRX1_HVT box_sel_reg_1_ ( .D(1'b0), .SETB(n174), .RSTB(n_box_sel_1_), 
        .CLK(clk), .Q(box_sel[1]) );
  DFFSSRX1_HVT box_sel_reg_0_ ( .D(n369), .SETB(n1662), .RSTB(n181), .CLK(clk), 
        .Q(box_sel[0]) );
  DFFSSRX1_HVT box_sel_reg_3_ ( .D(n368), .SETB(n1655), .RSTB(n181), .CLK(clk), 
        .Q(box_sel[3]) );
  DFFSSRX1_HVT row_reg_2_ ( .D(1'b0), .SETB(n193), .RSTB(n_row[2]), .CLK(
        net22657), .Q(row[2]), .QN(n252) );
  DFFSSRX1_HVT row_delay_reg_2_ ( .D(1'b0), .SETB(n207), .RSTB(row[2]), .CLK(
        clk), .Q(row_delay[2]) );
  DFFSSRX1_HVT write_row_reg_2_ ( .D(1'b0), .SETB(n187), .RSTB(row_delay[2]), 
        .CLK(clk), .Q(write_row[2]) );
  DFFSSRX1_HVT row_enable_reg_2_ ( .D(1'b0), .SETB(n184), .RSTB(write_row[2]), 
        .CLK(clk), .Q(row_enable[2]) );
  DFFSSRX1_HVT write_row_conv1_reg_2_ ( .D(1'b0), .SETB(n197), .RSTB(
        row_enable[2]), .CLK(clk), .Q(write_row_conv1[2]), .QN(n296) );
  DFFSSRX1_HVT row_reg_3_ ( .D(1'b0), .SETB(n193), .RSTB(n_row[3]), .CLK(
        net22657), .Q(row[3]), .QN(n321) );
  DFFSSRX1_HVT row_delay_reg_3_ ( .D(1'b0), .SETB(n199), .RSTB(row[3]), .CLK(
        clk), .Q(row_delay[3]) );
  DFFSSRX1_HVT write_row_reg_3_ ( .D(1'b0), .SETB(n195), .RSTB(row_delay[3]), 
        .CLK(clk), .Q(write_row[3]) );
  DFFSSRX1_HVT row_enable_reg_3_ ( .D(1'b0), .SETB(n208), .RSTB(write_row[3]), 
        .CLK(clk), .Q(row_enable[3]) );
  DFFSSRX1_HVT write_row_conv1_reg_3_ ( .D(1'b0), .SETB(n208), .RSTB(
        row_enable[3]), .CLK(clk), .Q(write_row_conv1[3]), .QN(n405) );
  DFFSSRX1_HVT channel_cnt_reg_4_ ( .D(1'b0), .SETB(n186), .RSTB(net22933), 
        .CLK(net22940), .Q(channel_cnt[4]), .QN(n311) );
  DFFSSRX1_HVT channel_cnt_reg_3_ ( .D(1'b0), .SETB(n183), .RSTB(net22934), 
        .CLK(net22940), .Q(channel_cnt[3]) );
  DFFSSRX1_HVT channel_cnt_reg_2_ ( .D(1'b0), .SETB(n198), .RSTB(net22935), 
        .CLK(net22940), .Q(channel_cnt[2]), .QN(n420) );
  DFFSSRX1_HVT channel_cnt_reg_1_ ( .D(1'b0), .SETB(n194), .RSTB(net22936), 
        .CLK(net22940), .Q(channel_cnt[1]) );
  DFFSSRX1_HVT load_conv1_bias_enable_reg ( .D(1'b0), .SETB(n200), .RSTB(n1020), .CLK(clk), .Q(load_conv1_bias_enable) );
  DFFSSRX1_HVT sram_raddr_weight_reg_7_ ( .D(1'b0), .SETB(n196), .RSTB(
        net22782), .CLK(net22855), .Q(sram_raddr_weight[7]), .QN(n410) );
  DFFSSRX1_HVT conv1_bias_set_reg_7_ ( .D(1'b0), .SETB(n229), .RSTB(
        sram_raddr_weight[7]), .CLK(clk), .Q(conv1_bias_set[7]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_6_ ( .D(1'b0), .SETB(n207), .RSTB(
        net22789), .CLK(net22855), .Q(sram_raddr_weight[6]), .QN(n407) );
  DFFSSRX1_HVT conv1_bias_set_reg_6_ ( .D(1'b0), .SETB(n185), .RSTB(
        sram_raddr_weight[6]), .CLK(clk), .Q(conv1_bias_set[6]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_5_ ( .D(1'b0), .SETB(n182), .RSTB(
        net22796), .CLK(net22855), .Q(sram_raddr_weight[5]), .QN(n422) );
  DFFSSRX1_HVT conv1_bias_set_reg_5_ ( .D(1'b0), .SETB(n175), .RSTB(
        sram_raddr_weight[5]), .CLK(clk), .Q(conv1_bias_set[5]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_3_ ( .D(1'b0), .SETB(n177), .RSTB(
        net22817), .CLK(net22855), .Q(sram_raddr_weight[3]), .QN(n417) );
  DFFSSRX1_HVT conv1_bias_set_reg_3_ ( .D(1'b0), .SETB(n176), .RSTB(
        sram_raddr_weight[3]), .CLK(clk), .Q(conv1_bias_set[3]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_16_ ( .D(1'b0), .SETB(n174), .RSTB(
        net22691), .CLK(net22757), .Q(sram_raddr_weight[16]), .QN(n451) );
  DFFSSRX1_HVT conv1_bias_set_reg_16_ ( .D(1'b0), .SETB(n175), .RSTB(
        sram_raddr_weight[16]), .CLK(clk), .Q(conv1_bias_set[16]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_15_ ( .D(1'b0), .SETB(n208), .RSTB(
        net22698), .CLK(net22757), .Q(sram_raddr_weight[15]), .QN(n292) );
  DFFSSRX1_HVT conv1_bias_set_reg_15_ ( .D(1'b0), .SETB(n187), .RSTB(
        sram_raddr_weight[15]), .CLK(clk), .Q(conv1_bias_set[15]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_14_ ( .D(1'b0), .SETB(n184), .RSTB(
        net22705), .CLK(net22757), .Q(sram_raddr_weight[14]), .QN(n362) );
  DFFSSRX1_HVT conv1_bias_set_reg_14_ ( .D(1'b0), .SETB(n175), .RSTB(
        sram_raddr_weight[14]), .CLK(clk), .Q(conv1_bias_set[14]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_13_ ( .D(1'b0), .SETB(n177), .RSTB(
        net22712), .CLK(net22757), .Q(sram_raddr_weight[13]) );
  DFFSSRX1_HVT conv1_bias_set_reg_13_ ( .D(1'b0), .SETB(n176), .RSTB(
        sram_raddr_weight[13]), .CLK(clk), .Q(conv1_bias_set[13]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_12_ ( .D(1'b0), .SETB(n174), .RSTB(
        net22719), .CLK(net22757), .Q(sram_raddr_weight[12]), .QN(n414) );
  DFFSSRX1_HVT conv1_bias_set_reg_12_ ( .D(1'b0), .SETB(n229), .RSTB(
        sram_raddr_weight[12]), .CLK(clk), .Q(conv1_bias_set[12]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_11_ ( .D(1'b0), .SETB(n207), .RSTB(
        net22726), .CLK(net22757), .Q(sram_raddr_weight[11]) );
  DFFSSRX1_HVT conv1_bias_set_reg_11_ ( .D(1'b0), .SETB(n186), .RSTB(
        sram_raddr_weight[11]), .CLK(clk), .Q(conv1_bias_set[11]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_10_ ( .D(1'b0), .SETB(n183), .RSTB(
        net22733), .CLK(net22757), .Q(sram_raddr_weight[10]), .QN(n415) );
  DFFSSRX1_HVT conv1_bias_set_reg_10_ ( .D(1'b0), .SETB(n197), .RSTB(
        sram_raddr_weight[10]), .CLK(clk), .Q(conv1_bias_set[10]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_9_ ( .D(1'b0), .SETB(n193), .RSTB(
        net22747), .CLK(net22757), .Q(sram_raddr_weight[9]), .QN(n293) );
  DFFSSRX1_HVT conv1_bias_set_reg_9_ ( .D(1'b0), .SETB(n199), .RSTB(
        sram_raddr_weight[9]), .CLK(clk), .Q(conv1_bias_set[9]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_8_ ( .D(1'b0), .SETB(n195), .RSTB(
        net22754), .CLK(net22757), .Q(sram_raddr_weight[8]), .QN(n395) );
  DFFSSRX1_HVT conv1_bias_set_reg_8_ ( .D(1'b0), .SETB(n174), .RSTB(
        sram_raddr_weight[8]), .CLK(clk), .Q(conv1_bias_set[8]) );
  DFFSSRX1_HVT load_conv2_bias0_enable_reg ( .D(1'b0), .SETB(n208), .RSTB(
        n1021), .CLK(clk), .Q(load_conv2_bias0_enable) );
  DFFSSRX1_HVT conv1_weight_done_reg ( .D(1'b0), .SETB(n185), .RSTB(
        n_conv1_weight_done), .CLK(clk), .Q(conv1_weight_done), .QN(n250) );
  DFFSSRX1_HVT load_data_enable_reg ( .D(1'b0), .SETB(n182), .RSTB(
        n_load_data_enable), .CLK(clk), .Q(load_data_enable) );
  DFFSSRX1_HVT write_enable_reg ( .D(1'b0), .SETB(n198), .RSTB(n_write_enable), 
        .CLK(clk), .Q(write_enable) );
  DFFSSRX1_HVT delay_write_enable_reg ( .D(1'b0), .SETB(n194), .RSTB(
        write_enable), .CLK(clk), .Q(delay_write_enable) );
  DFFSSRX1_HVT delay2_write_enable_reg ( .D(1'b0), .SETB(n200), .RSTB(
        delay_write_enable), .CLK(clk), .Q(delay2_write_enable) );
  DFFSSRX1_HVT delay3_write_enable_reg ( .D(1'b0), .SETB(n196), .RSTB(
        delay2_write_enable), .CLK(clk), .Q(delay3_write_enable) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_9_ ( .D(1'b0), .SETB(N2914), .RSTB(
        net22863), .CLK(net22893), .Q(delay1_sram_waddr_b[9]) );
  DFFSSRX1_HVT sram_waddr_b_reg_9_ ( .D(1'b0), .SETB(n229), .RSTB(
        delay1_sram_waddr_b[9]), .CLK(clk), .Q(sram_waddr_b[9]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_8_ ( .D(1'b0), .SETB(N2914), .RSTB(
        net22866), .CLK(net22893), .Q(delay1_sram_waddr_b[8]), .QN(n431) );
  DFFSSRX1_HVT sram_waddr_b_reg_8_ ( .D(1'b0), .SETB(n207), .RSTB(
        delay1_sram_waddr_b[8]), .CLK(clk), .Q(sram_waddr_b[8]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_7_ ( .D(1'b0), .SETB(N2914), .RSTB(
        net22869), .CLK(net22893), .Q(delay1_sram_waddr_b[7]) );
  DFFSSRX1_HVT sram_waddr_b_reg_7_ ( .D(1'b0), .SETB(n187), .RSTB(
        delay1_sram_waddr_b[7]), .CLK(clk), .Q(sram_waddr_b[7]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_6_ ( .D(1'b0), .SETB(N2914), .RSTB(
        net22872), .CLK(net22893), .Q(delay1_sram_waddr_b[6]), .QN(n375) );
  DFFSSRX1_HVT sram_waddr_b_reg_6_ ( .D(1'b0), .SETB(n184), .RSTB(
        delay1_sram_waddr_b[6]), .CLK(clk), .Q(sram_waddr_b[6]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_5_ ( .D(1'b0), .SETB(N2914), .RSTB(
        net22875), .CLK(net22893), .Q(delay1_sram_waddr_b[5]) );
  DFFSSRX1_HVT sram_waddr_b_reg_5_ ( .D(1'b0), .SETB(n175), .RSTB(
        delay1_sram_waddr_b[5]), .CLK(clk), .Q(sram_waddr_b[5]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_4_ ( .D(1'b0), .SETB(N2914), .RSTB(
        net22878), .CLK(net22893), .Q(delay1_sram_waddr_b[4]), .QN(n376) );
  DFFSSRX1_HVT sram_waddr_b_reg_4_ ( .D(1'b0), .SETB(n177), .RSTB(
        delay1_sram_waddr_b[4]), .CLK(clk), .Q(sram_waddr_b[4]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_3_ ( .D(1'b0), .SETB(N2914), .RSTB(
        net22881), .CLK(net22893), .Q(delay1_sram_waddr_b[3]) );
  DFFSSRX1_HVT sram_waddr_b_reg_3_ ( .D(1'b0), .SETB(n176), .RSTB(
        delay1_sram_waddr_b[3]), .CLK(clk), .Q(sram_waddr_b[3]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_2_ ( .D(1'b0), .SETB(N2914), .RSTB(
        net22884), .CLK(net22893), .Q(delay1_sram_waddr_b[2]), .QN(n409) );
  DFFSSRX1_HVT sram_waddr_b_reg_2_ ( .D(1'b0), .SETB(n174), .RSTB(
        delay1_sram_waddr_b[2]), .CLK(clk), .Q(sram_waddr_b[2]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_1_ ( .D(1'b0), .SETB(N2914), .RSTB(
        net22887), .CLK(net22893), .Q(delay1_sram_waddr_b[1]) );
  DFFSSRX1_HVT sram_waddr_b_reg_1_ ( .D(1'b0), .SETB(n182), .RSTB(
        delay1_sram_waddr_b[1]), .CLK(clk), .Q(sram_waddr_b[1]) );
  DFFSSRX1_HVT delay1_sram_waddr_b_reg_0_ ( .D(1'b0), .SETB(N2914), .RSTB(
        net22890), .CLK(net22893), .Q(delay1_sram_waddr_b[0]) );
  DFFSSRX1_HVT sram_waddr_b_reg_0_ ( .D(1'b0), .SETB(n208), .RSTB(
        delay1_sram_waddr_b[0]), .CLK(clk), .Q(sram_waddr_b[0]) );
  DFFSSRX1_HVT sram_bytemask_b_reg_3_ ( .D(1'b0), .SETB(n186), .RSTB(
        n_sram_bytemask_b[3]), .CLK(clk), .Q(sram_bytemask_b[3]) );
  DFFSSRX1_HVT sram_bytemask_b_reg_2_ ( .D(1'b0), .SETB(n183), .RSTB(
        n_sram_bytemask_b[2]), .CLK(clk), .Q(sram_bytemask_b[2]) );
  DFFSSRX1_HVT sram_bytemask_b_reg_1_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_bytemask_b[1]), .CLK(clk), .Q(sram_bytemask_b[1]) );
  DFFSSRX1_HVT sram_bytemask_b_reg_0_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_bytemask_b[0]), .CLK(clk), .Q(sram_bytemask_b[0]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_1_ ( .D(1'b0), .SETB(n176), .RSTB(
        net22838), .CLK(net22855), .Q(sram_raddr_weight[1]), .QN(n421) );
  DFFSSRX1_HVT conv1_bias_set_reg_1_ ( .D(1'b0), .SETB(n174), .RSTB(
        sram_raddr_weight[1]), .CLK(clk), .Q(conv1_bias_set[1]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_0_ ( .D(1'b0), .SETB(n229), .RSTB(
        net22852), .CLK(net22855), .Q(sram_raddr_weight[0]), .QN(n300) );
  DFFSSRX1_HVT conv1_bias_set_reg_0_ ( .D(1'b0), .SETB(n207), .RSTB(
        sram_raddr_weight[0]), .CLK(clk), .Q(conv1_bias_set[0]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_2_ ( .D(1'b0), .SETB(n185), .RSTB(
        net22824), .CLK(net22855), .Q(sram_raddr_weight[2]), .QN(n294) );
  DFFSSRX1_HVT conv1_bias_set_reg_2_ ( .D(1'b0), .SETB(n182), .RSTB(
        sram_raddr_weight[2]), .CLK(clk), .Q(conv1_bias_set[2]) );
  DFFSSRX1_HVT sram_raddr_weight_reg_4_ ( .D(1'b0), .SETB(n197), .RSTB(
        net22810), .CLK(net22855), .Q(sram_raddr_weight[4]), .QN(n433) );
  DFFSSRX1_HVT conv1_bias_set_reg_4_ ( .D(1'b0), .SETB(n193), .RSTB(
        sram_raddr_weight[4]), .CLK(clk), .Q(conv1_bias_set[4]) );
  DFFSSRX1_HVT load_conv2_bias1_enable_reg ( .D(1'b0), .SETB(n199), .RSTB(
        n1022), .CLK(clk), .Q(load_conv2_bias1_enable) );
  DFFSSRX1_HVT addr_change_reg_0_ ( .D(1'b0), .SETB(n195), .RSTB(net22949), 
        .CLK(net22952), .Q(addr_change[0]) );
  DFFSSRX1_HVT addr_change_reg_1_ ( .D(1'b0), .SETB(n184), .RSTB(net22948), 
        .CLK(net22952), .Q(addr_change[1]) );
  DFFSSRX1_HVT addr_change_reg_2_ ( .D(1'b0), .SETB(n208), .RSTB(net22947), 
        .CLK(net22952), .Q(addr_change[2]) );
  DFFSSRX1_HVT addr_change_reg_3_ ( .D(1'b0), .SETB(n187), .RSTB(net22946), 
        .CLK(net22952), .Q(addr_change[3]), .QN(n441) );
  DFFSSRX1_HVT addr_change_reg_4_ ( .D(1'b0), .SETB(n184), .RSTB(net22945), 
        .CLK(net22952), .Q(addr_change[4]), .QN(n447) );
  DFFSSRX1_HVT delay_addr_change_reg_4_ ( .D(1'b0), .SETB(n198), .RSTB(
        addr_change[4]), .CLK(clk), .Q(delay_addr_change[4]) );
  DFFSSRX1_HVT delay_addr_change_reg_3_ ( .D(1'b0), .SETB(n194), .RSTB(
        addr_change[3]), .CLK(clk), .Q(delay_addr_change[3]) );
  DFFSSRX1_HVT delay_addr_change_reg_2_ ( .D(1'b0), .SETB(n200), .RSTB(
        addr_change[2]), .CLK(clk), .Q(delay_addr_change[2]) );
  DFFSSRX1_HVT delay_addr_change_reg_1_ ( .D(1'b0), .SETB(n196), .RSTB(
        addr_change[1]), .CLK(clk), .Q(delay_addr_change[1]) );
  DFFSSRX1_HVT delay_addr_change_reg_0_ ( .D(1'b0), .SETB(n229), .RSTB(
        addr_change[0]), .CLK(clk), .Q(delay_addr_change[0]) );
  DFFSSRX1_HVT delay2_addr_change_reg_4_ ( .D(1'b0), .SETB(n207), .RSTB(
        delay_addr_change[4]), .CLK(clk), .Q(delay2_addr_change[4]) );
  DFFSSRX1_HVT delay2_addr_change_reg_3_ ( .D(1'b0), .SETB(n186), .RSTB(
        delay_addr_change[3]), .CLK(clk), .Q(delay2_addr_change[3]) );
  DFFSSRX1_HVT delay2_addr_change_reg_2_ ( .D(1'b0), .SETB(n183), .RSTB(
        delay_addr_change[2]), .CLK(clk), .Q(delay2_addr_change[2]) );
  DFFSSRX1_HVT delay2_addr_change_reg_1_ ( .D(1'b0), .SETB(n175), .RSTB(
        delay_addr_change[1]), .CLK(clk), .Q(delay2_addr_change[1]) );
  DFFSSRX1_HVT delay2_addr_change_reg_0_ ( .D(1'b0), .SETB(n177), .RSTB(
        delay_addr_change[0]), .CLK(clk), .Q(delay2_addr_change[0]) );
  DFFSSRX1_HVT delay3_addr_change_reg_4_ ( .D(1'b0), .SETB(n176), .RSTB(
        delay2_addr_change[4]), .CLK(clk), .Q(delay3_addr_change[4]), .QN(n460) );
  DFFSSRX1_HVT delay3_addr_change_reg_3_ ( .D(1'b0), .SETB(n174), .RSTB(
        delay2_addr_change[3]), .CLK(clk), .Q(delay3_addr_change[3]), .QN(n318) );
  DFFSSRX1_HVT delay3_addr_change_reg_2_ ( .D(1'b0), .SETB(n183), .RSTB(
        delay2_addr_change[2]), .CLK(clk), .Q(delay3_addr_change[2]), .QN(n257) );
  DFFSSRX1_HVT delay3_addr_change_reg_1_ ( .D(1'b0), .SETB(n208), .RSTB(
        delay2_addr_change[1]), .CLK(clk), .Q(delay3_addr_change[1]) );
  DFFSSRX1_HVT delay3_addr_change_reg_0_ ( .D(1'b0), .SETB(n185), .RSTB(
        delay2_addr_change[0]), .CLK(clk), .Q(delay3_addr_change[0]) );
  DFFSSRX1_HVT delay_channel_reg_4_ ( .D(1'b0), .SETB(n206), .RSTB(
        channel_cnt[4]), .CLK(clk), .Q(delay_channel[4]) );
  DFFSSRX1_HVT delay_channel_reg_3_ ( .D(1'b0), .SETB(n199), .RSTB(
        channel_cnt[3]), .CLK(clk), .Q(delay_channel[3]) );
  DFFSSRX1_HVT delay_channel_reg_2_ ( .D(1'b0), .SETB(n184), .RSTB(
        channel_cnt[2]), .CLK(clk), .Q(delay_channel[2]) );
  DFFSSRX1_HVT delay_channel_reg_1_ ( .D(1'b0), .SETB(n198), .RSTB(
        channel_cnt[1]), .CLK(clk), .Q(delay_channel[1]) );
  DFFSSRX1_HVT delay_channel_reg_0_ ( .D(1'b0), .SETB(n196), .RSTB(
        channel_cnt[0]), .CLK(clk), .Q(delay_channel[0]) );
  DFFSSRX1_HVT delay2_channel_reg_4_ ( .D(1'b0), .SETB(n197), .RSTB(
        delay_channel[4]), .CLK(clk), .Q(delay2_channel[4]) );
  DFFSSRX1_HVT delay2_channel_reg_3_ ( .D(1'b0), .SETB(n195), .RSTB(
        delay_channel[3]), .CLK(clk), .Q(delay2_channel[3]) );
  DFFSSRX1_HVT delay2_channel_reg_2_ ( .D(1'b0), .SETB(n210), .RSTB(
        delay_channel[2]), .CLK(clk), .Q(delay2_channel[2]) );
  DFFSSRX1_HVT delay2_channel_reg_1_ ( .D(1'b0), .SETB(n194), .RSTB(
        delay_channel[1]), .CLK(clk), .Q(delay2_channel[1]) );
  DFFSSRX1_HVT delay2_channel_reg_0_ ( .D(1'b0), .SETB(n185), .RSTB(
        delay_channel[0]), .CLK(clk), .Q(delay2_channel[0]) );
  DFFSSRX1_HVT channel_reg_4_ ( .D(1'b0), .SETB(n193), .RSTB(delay2_channel[4]), .CLK(clk), .Q(channel[4]) );
  DFFSSRX1_HVT channel_reg_3_ ( .D(1'b0), .SETB(n187), .RSTB(delay2_channel[3]), .CLK(clk), .Q(channel[3]) );
  DFFSSRX1_HVT channel_reg_2_ ( .D(1'b0), .SETB(n206), .RSTB(delay2_channel[2]), .CLK(clk), .Q(channel[2]) );
  DFFSSRX1_HVT channel_reg_1_ ( .D(1'b0), .SETB(n200), .RSTB(delay2_channel[1]), .CLK(clk), .Q(channel[1]) );
  DFFSSRX1_HVT channel_reg_0_ ( .D(1'b0), .SETB(n182), .RSTB(delay2_channel[0]), .CLK(clk), .Q(channel[0]) );
  DFFSSRX1_HVT delay1_state_reg_3_ ( .D(1'b0), .SETB(n182), .RSTB(state[3]), 
        .CLK(clk), .Q(delay1_state[3]) );
  DFFSSRX1_HVT delay2_state_reg_3_ ( .D(1'b0), .SETB(n175), .RSTB(
        delay1_state[3]), .CLK(clk), .Q(delay2_state[3]) );
  DFFSSRX1_HVT delay3_state_reg_3_ ( .D(1'b0), .SETB(n177), .RSTB(
        delay2_state[3]), .CLK(clk), .QN(n1027) );
  DFFSSRX1_HVT delay1_state_reg_2_ ( .D(1'b0), .SETB(n176), .RSTB(state[2]), 
        .CLK(clk), .Q(delay1_state[2]) );
  DFFSSRX1_HVT delay2_state_reg_2_ ( .D(1'b0), .SETB(n174), .RSTB(
        delay1_state[2]), .CLK(clk), .Q(delay2_state[2]) );
  DFFSSRX1_HVT delay3_state_reg_2_ ( .D(1'b0), .SETB(n229), .RSTB(
        delay2_state[2]), .CLK(clk), .Q(delay3_state[2]) );
  DFFSSRX1_HVT delay1_state_reg_1_ ( .D(1'b0), .SETB(n207), .RSTB(state[1]), 
        .CLK(clk), .Q(delay1_state[1]) );
  DFFSSRX1_HVT delay2_state_reg_1_ ( .D(1'b0), .SETB(n187), .RSTB(
        delay1_state[1]), .CLK(clk), .Q(delay2_state[1]) );
  DFFSSRX1_HVT delay3_state_reg_1_ ( .D(1'b0), .SETB(n184), .RSTB(
        delay2_state[1]), .CLK(clk), .Q(delay3_state[1]) );
  DFFSSRX1_HVT delay1_state_reg_0_ ( .D(1'b0), .SETB(n197), .RSTB(state[0]), 
        .CLK(clk), .Q(delay1_state[0]) );
  DFFSSRX1_HVT delay2_state_reg_0_ ( .D(1'b0), .SETB(n193), .RSTB(
        delay1_state[0]), .CLK(clk), .Q(delay2_state[0]) );
  DFFSSRX1_HVT delay3_state_reg_0_ ( .D(1'b0), .SETB(n199), .RSTB(
        delay2_state[0]), .CLK(clk), .Q(delay3_state[0]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_9_ ( .D(1'b0), .SETB(n195), .RSTB(
        net22916), .CLK(net22928), .Q(delay1_sram_waddr_d[9]), .QN(n455) );
  DFFSSRX1_HVT sram_waddr_d_reg_9_ ( .D(1'b0), .SETB(n207), .RSTB(
        delay1_sram_waddr_d[9]), .CLK(clk), .Q(sram_waddr_d[9]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_8_ ( .D(1'b0), .SETB(n208), .RSTB(
        net22917), .CLK(net22928), .Q(delay1_sram_waddr_d[8]) );
  DFFSSRX1_HVT sram_waddr_d_reg_8_ ( .D(1'b0), .SETB(n186), .RSTB(
        delay1_sram_waddr_d[8]), .CLK(clk), .Q(sram_waddr_d[8]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_7_ ( .D(1'b0), .SETB(n183), .RSTB(
        net22918), .CLK(net22928), .Q(delay1_sram_waddr_d[7]) );
  DFFSSRX1_HVT sram_waddr_d_reg_7_ ( .D(1'b0), .SETB(n198), .RSTB(
        delay1_sram_waddr_d[7]), .CLK(clk), .Q(sram_waddr_d[7]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_6_ ( .D(1'b0), .SETB(n194), .RSTB(
        net22919), .CLK(net22928), .Q(delay1_sram_waddr_d[6]) );
  DFFSSRX1_HVT sram_waddr_d_reg_6_ ( .D(1'b0), .SETB(n200), .RSTB(
        delay1_sram_waddr_d[6]), .CLK(clk), .Q(sram_waddr_d[6]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_5_ ( .D(1'b0), .SETB(n196), .RSTB(
        net22920), .CLK(net22928), .Q(delay1_sram_waddr_d[5]) );
  DFFSSRX1_HVT sram_waddr_d_reg_5_ ( .D(1'b0), .SETB(n229), .RSTB(
        delay1_sram_waddr_d[5]), .CLK(clk), .Q(sram_waddr_d[5]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_4_ ( .D(1'b0), .SETB(n207), .RSTB(
        net22921), .CLK(net22928), .Q(delay1_sram_waddr_d[4]) );
  DFFSSRX1_HVT sram_waddr_d_reg_4_ ( .D(1'b0), .SETB(n185), .RSTB(
        delay1_sram_waddr_d[4]), .CLK(clk), .Q(sram_waddr_d[4]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_3_ ( .D(1'b0), .SETB(n182), .RSTB(
        net22922), .CLK(net22928), .Q(delay1_sram_waddr_d[3]) );
  DFFSSRX1_HVT sram_waddr_d_reg_3_ ( .D(1'b0), .SETB(n175), .RSTB(
        delay1_sram_waddr_d[3]), .CLK(clk), .Q(sram_waddr_d[3]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_2_ ( .D(1'b0), .SETB(n177), .RSTB(
        net22923), .CLK(net22928), .Q(delay1_sram_waddr_d[2]) );
  DFFSSRX1_HVT sram_waddr_d_reg_2_ ( .D(1'b0), .SETB(n176), .RSTB(
        delay1_sram_waddr_d[2]), .CLK(clk), .Q(sram_waddr_d[2]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_1_ ( .D(1'b0), .SETB(n174), .RSTB(
        net22924), .CLK(net22928), .Q(delay1_sram_waddr_d[1]) );
  DFFSSRX1_HVT sram_waddr_d_reg_1_ ( .D(1'b0), .SETB(n208), .RSTB(
        delay1_sram_waddr_d[1]), .CLK(clk), .Q(sram_waddr_d[1]) );
  DFFSSRX1_HVT delay1_sram_waddr_d_reg_0_ ( .D(1'b0), .SETB(n208), .RSTB(
        net22925), .CLK(net22928), .Q(delay1_sram_waddr_d[0]), .QN(n426) );
  DFFSSRX1_HVT sram_waddr_d_reg_0_ ( .D(1'b0), .SETB(n210), .RSTB(
        delay1_sram_waddr_d[0]), .CLK(clk), .Q(sram_waddr_d[0]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_9_ ( .D(1'b0), .SETB(n206), .RSTB(
        net22900), .CLK(net22912), .Q(delay1_sram_waddr_c[9]), .QN(n454) );
  DFFSSRX1_HVT sram_waddr_c_reg_9_ ( .D(1'b0), .SETB(n175), .RSTB(
        delay1_sram_waddr_c[9]), .CLK(clk), .Q(sram_waddr_c[9]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_8_ ( .D(1'b0), .SETB(n177), .RSTB(
        net22901), .CLK(net22912), .Q(delay1_sram_waddr_c[8]) );
  DFFSSRX1_HVT sram_waddr_c_reg_8_ ( .D(1'b0), .SETB(n176), .RSTB(
        delay1_sram_waddr_c[8]), .CLK(clk), .Q(sram_waddr_c[8]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_7_ ( .D(1'b0), .SETB(n174), .RSTB(
        net22902), .CLK(net22912), .Q(delay1_sram_waddr_c[7]) );
  DFFSSRX1_HVT sram_waddr_c_reg_7_ ( .D(1'b0), .SETB(n184), .RSTB(
        delay1_sram_waddr_c[7]), .CLK(clk), .Q(sram_waddr_c[7]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_6_ ( .D(1'b0), .SETB(n207), .RSTB(
        net22903), .CLK(net22912), .Q(delay1_sram_waddr_c[6]) );
  DFFSSRX1_HVT sram_waddr_c_reg_6_ ( .D(1'b0), .SETB(n210), .RSTB(
        delay1_sram_waddr_c[6]), .CLK(clk), .Q(sram_waddr_c[6]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_5_ ( .D(1'b0), .SETB(n206), .RSTB(
        net22904), .CLK(net22912), .Q(delay1_sram_waddr_c[5]) );
  DFFSSRX1_HVT sram_waddr_c_reg_5_ ( .D(1'b0), .SETB(n197), .RSTB(
        delay1_sram_waddr_c[5]), .CLK(clk), .Q(sram_waddr_c[5]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_4_ ( .D(1'b0), .SETB(n193), .RSTB(
        net22905), .CLK(net22912), .Q(delay1_sram_waddr_c[4]) );
  DFFSSRX1_HVT sram_waddr_c_reg_4_ ( .D(1'b0), .SETB(n199), .RSTB(
        delay1_sram_waddr_c[4]), .CLK(clk), .Q(sram_waddr_c[4]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_3_ ( .D(1'b0), .SETB(n195), .RSTB(
        net22906), .CLK(net22912), .Q(delay1_sram_waddr_c[3]) );
  DFFSSRX1_HVT sram_waddr_c_reg_3_ ( .D(1'b0), .SETB(n229), .RSTB(
        delay1_sram_waddr_c[3]), .CLK(clk), .Q(sram_waddr_c[3]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_2_ ( .D(1'b0), .SETB(n208), .RSTB(
        net22907), .CLK(net22912), .Q(delay1_sram_waddr_c[2]) );
  DFFSSRX1_HVT sram_waddr_c_reg_2_ ( .D(1'b0), .SETB(n210), .RSTB(
        delay1_sram_waddr_c[2]), .CLK(clk), .Q(sram_waddr_c[2]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_1_ ( .D(1'b0), .SETB(n206), .RSTB(
        net22908), .CLK(net22912), .Q(delay1_sram_waddr_c[1]) );
  DFFSSRX1_HVT sram_waddr_c_reg_1_ ( .D(1'b0), .SETB(n198), .RSTB(
        delay1_sram_waddr_c[1]), .CLK(clk), .Q(sram_waddr_c[1]) );
  DFFSSRX1_HVT delay1_sram_waddr_c_reg_0_ ( .D(1'b0), .SETB(n194), .RSTB(
        net22909), .CLK(net22912), .Q(delay1_sram_waddr_c[0]), .QN(n425) );
  DFFSSRX1_HVT sram_waddr_c_reg_0_ ( .D(1'b0), .SETB(n200), .RSTB(
        delay1_sram_waddr_c[0]), .CLK(clk), .Q(sram_waddr_c[0]) );
  DFFSSRX1_HVT sram_raddr_a7_reg_9_ ( .D(1'b0), .SETB(n196), .RSTB(
        n_sram_raddr_a7[9]), .CLK(net23433), .Q(sram_raddr_a7[9]) );
  DFFSSRX1_HVT sram_raddr_a7_reg_8_ ( .D(1'b0), .SETB(n183), .RSTB(
        n_sram_raddr_a7[8]), .CLK(net23433), .Q(sram_raddr_a7[8]) );
  DFFSSRX1_HVT sram_raddr_a7_reg_7_ ( .D(1'b0), .SETB(n207), .RSTB(
        n_sram_raddr_a7[7]), .CLK(net23433), .Q(sram_raddr_a7[7]) );
  DFFSSRX1_HVT sram_raddr_a7_reg_6_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_a7[6]), .CLK(net23433), .Q(sram_raddr_a7[6]) );
  DFFSSRX1_HVT sram_raddr_a7_reg_5_ ( .D(1'b0), .SETB(n206), .RSTB(
        n_sram_raddr_a7[5]), .CLK(net23433), .Q(sram_raddr_a7[5]) );
  DFFSSRX1_HVT sram_raddr_a7_reg_4_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_a7[4]), .CLK(net23433), .Q(sram_raddr_a7[4]) );
  DFFSSRX1_HVT sram_raddr_a7_reg_3_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_a7[3]), .CLK(net23433), .Q(sram_raddr_a7[3]), .QN(n453)
         );
  DFFSSRX1_HVT sram_raddr_a7_reg_2_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_a7[2]), .CLK(net23433), .Q(sram_raddr_a7[2]) );
  DFFSSRX1_HVT sram_raddr_a7_reg_1_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_raddr_a7[1]), .CLK(net23433), .Q(sram_raddr_a7[1]), .QN(n429)
         );
  DFFSSRX1_HVT sram_raddr_a7_reg_0_ ( .D(1'b0), .SETB(n229), .RSTB(
        n_sram_raddr_a7[0]), .CLK(net23433), .Q(sram_raddr_a7[0]), .QN(n289)
         );
  DFFSSRX1_HVT sram_raddr_a8_reg_9_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_a8[9]), .CLK(net24760), .Q(sram_raddr_a8[9]) );
  DFFSSRX1_HVT sram_raddr_a8_reg_8_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_a8[8]), .CLK(net24760), .Q(sram_raddr_a8[8]) );
  DFFSSRX1_HVT sram_raddr_a8_reg_7_ ( .D(1'b0), .SETB(n206), .RSTB(
        n_sram_raddr_a8[7]), .CLK(net24760), .Q(sram_raddr_a8[7]) );
  DFFSSRX1_HVT sram_raddr_a8_reg_6_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_a8[6]), .CLK(net24760), .Q(sram_raddr_a8[6]) );
  DFFSSRX1_HVT sram_raddr_a8_reg_5_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_a8[5]), .CLK(net24760), .Q(sram_raddr_a8[5]) );
  DFFSSRX1_HVT sram_raddr_a8_reg_4_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_a8[4]), .CLK(net24760), .Q(sram_raddr_a8[4]) );
  DFFSSRX1_HVT sram_raddr_a8_reg_3_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_raddr_a8[3]), .CLK(net24760), .Q(sram_raddr_a8[3]) );
  DFFSSRX1_HVT sram_raddr_a8_reg_2_ ( .D(1'b0), .SETB(n229), .RSTB(
        n_sram_raddr_a8[2]), .CLK(net24760), .Q(sram_raddr_a8[2]), .QN(n438)
         );
  DFFSSRX1_HVT sram_raddr_a8_reg_1_ ( .D(1'b0), .SETB(n207), .RSTB(
        n_sram_raddr_a8[1]), .CLK(net24760), .Q(sram_raddr_a8[1]), .QN(n437)
         );
  DFFSSRX1_HVT sram_raddr_a8_reg_0_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_a8[0]), .CLK(net24760), .Q(sram_raddr_a8[0]), .QN(n288)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_9_ ( .D(1'b0), .SETB(n206), .RSTB(
        n_sram_raddr_a0[9]), .CLK(net26088), .Q(sram_raddr_a0[9]), .QN(n444)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_8_ ( .D(1'b0), .SETB(n197), .RSTB(
        n_sram_raddr_a0[8]), .CLK(net26088), .Q(sram_raddr_a0[8]), .QN(n402)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_7_ ( .D(1'b0), .SETB(n193), .RSTB(
        n_sram_raddr_a0[7]), .CLK(net26088), .Q(sram_raddr_a0[7]), .QN(n355)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_6_ ( .D(1'b0), .SETB(n199), .RSTB(
        n_sram_raddr_a0[6]), .CLK(net26088), .Q(sram_raddr_a0[6]), .QN(n432)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_5_ ( .D(1'b0), .SETB(n195), .RSTB(
        n_sram_raddr_a0[5]), .CLK(net26088), .Q(sram_raddr_a0[5]), .QN(n291)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_4_ ( .D(1'b0), .SETB(n229), .RSTB(
        n_sram_raddr_a0[4]), .CLK(net26088), .Q(sram_raddr_a0[4]), .QN(n367)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_3_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_a0[3]), .CLK(net26088), .Q(sram_raddr_a0[3]), .QN(n237)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_2_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_a0[2]), .CLK(net26088), .Q(sram_raddr_a0[2]), .QN(n248)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_1_ ( .D(1'b0), .SETB(n206), .RSTB(
        n_sram_raddr_a0[1]), .CLK(net26088), .Q(sram_raddr_a0[1]), .QN(n297)
         );
  DFFSSRX1_HVT sram_raddr_a0_reg_0_ ( .D(1'b0), .SETB(n198), .RSTB(
        n_sram_raddr_a0[0]), .CLK(net26088), .Q(sram_raddr_a0[0]), .QN(n416)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_9_ ( .D(1'b0), .SETB(n194), .RSTB(
        n_sram_raddr_a1[9]), .CLK(net23878), .Q(sram_raddr_a1[9]), .QN(n445)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_8_ ( .D(1'b0), .SETB(n200), .RSTB(
        n_sram_raddr_a1[8]), .CLK(net23878), .Q(sram_raddr_a1[8]), .QN(n403)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_7_ ( .D(1'b0), .SETB(n196), .RSTB(
        n_sram_raddr_a1[7]), .CLK(net23878), .Q(sram_raddr_a1[7]), .QN(n423)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_6_ ( .D(1'b0), .SETB(n187), .RSTB(
        n_sram_raddr_a1[6]), .CLK(net23878), .Q(sram_raddr_a1[6]), .QN(n434)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_5_ ( .D(1'b0), .SETB(n207), .RSTB(
        n_sram_raddr_a1[5]), .CLK(net23878), .Q(sram_raddr_a1[5]), .QN(n380)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_4_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_a1[4]), .CLK(net23878), .Q(sram_raddr_a1[4]), .QN(n282)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_3_ ( .D(1'b0), .SETB(n206), .RSTB(
        n_sram_raddr_a1[3]), .CLK(net23878), .Q(sram_raddr_a1[3]), .QN(n236)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_2_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_a1[2]), .CLK(net23878), .Q(sram_raddr_a1[2]), .QN(n247)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_1_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_a1[1]), .CLK(net23878), .Q(sram_raddr_a1[1]), .QN(n436)
         );
  DFFSSRX1_HVT sram_raddr_a1_reg_0_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_a1[0]), .CLK(net23878), .Q(sram_raddr_a1[0]), .QN(n301)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_9_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_raddr_a2[9]), .CLK(net25205), .Q(sram_raddr_a2[9]), .QN(n446)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_8_ ( .D(1'b0), .SETB(n187), .RSTB(
        n_sram_raddr_a2[8]), .CLK(net25205), .Q(sram_raddr_a2[8]), .QN(n435)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_7_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_a2[7]), .CLK(net25205), .Q(sram_raddr_a2[7]), .QN(n356)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_6_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_a2[6]), .CLK(net25205), .Q(sram_raddr_a2[6]), .QN(n378)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_5_ ( .D(1'b0), .SETB(n206), .RSTB(
        n_sram_raddr_a2[5]), .CLK(net25205), .Q(sram_raddr_a2[5]), .QN(n385)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_4_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_a2[4]), .CLK(net25205), .Q(sram_raddr_a2[4]), .QN(n366)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_3_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_a2[3]), .CLK(net25205), .Q(sram_raddr_a2[3]), .QN(n370)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_2_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_a2[2]), .CLK(net25205), .Q(sram_raddr_a2[2]), .QN(n440)
         );
  DFFSSRX1_HVT sram_raddr_a2_reg_1_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_raddr_a2[1]), .CLK(net25205), .Q(sram_raddr_a2[1]) );
  DFFSSRX1_HVT sram_raddr_a2_reg_0_ ( .D(1'b0), .SETB(n186), .RSTB(
        n_sram_raddr_a2[0]), .CLK(net25205), .Q(sram_raddr_a2[0]), .QN(n427)
         );
  DFFSSRX1_HVT sram_raddr_a3_reg_9_ ( .D(1'b0), .SETB(n207), .RSTB(
        n_sram_raddr_a3[9]), .CLK(net26534), .Q(sram_raddr_a3[9]) );
  DFFSSRX1_HVT sram_raddr_a3_reg_8_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_a3[8]), .CLK(net26534), .Q(sram_raddr_a3[8]) );
  DFFSSRX1_HVT sram_raddr_a3_reg_7_ ( .D(1'b0), .SETB(n206), .RSTB(
        n_sram_raddr_a3[7]), .CLK(net26534), .Q(sram_raddr_a3[7]), .QN(n383)
         );
  DFFSSRX1_HVT sram_raddr_a3_reg_6_ ( .D(1'b0), .SETB(n197), .RSTB(
        n_sram_raddr_a3[6]), .CLK(net26534), .Q(sram_raddr_a3[6]), .QN(n349)
         );
  DFFSSRX1_HVT sram_raddr_a3_reg_5_ ( .D(1'b0), .SETB(n193), .RSTB(
        n_sram_raddr_a3[5]), .CLK(net26534), .Q(sram_raddr_a3[5]), .QN(n428)
         );
  DFFSSRX1_HVT sram_raddr_a3_reg_4_ ( .D(1'b0), .SETB(n199), .RSTB(
        n_sram_raddr_a3[4]), .CLK(net26534), .Q(sram_raddr_a3[4]), .QN(n279)
         );
  DFFSSRX1_HVT sram_raddr_a3_reg_3_ ( .D(1'b0), .SETB(n195), .RSTB(
        n_sram_raddr_a3[3]), .CLK(net26534), .Q(sram_raddr_a3[3]), .QN(n245)
         );
  DFFSSRX1_HVT sram_raddr_a3_reg_2_ ( .D(1'b0), .SETB(n186), .RSTB(
        n_sram_raddr_a3[2]), .CLK(net26534), .Q(sram_raddr_a3[2]), .QN(n234)
         );
  DFFSSRX1_HVT sram_raddr_a3_reg_1_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_a3[1]), .CLK(net26534), .Q(sram_raddr_a3[1]) );
  DFFSSRX1_HVT sram_raddr_a3_reg_0_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_a3[0]), .CLK(net26534), .Q(sram_raddr_a3[0]), .QN(n418)
         );
  DFFSSRX1_HVT sram_raddr_a4_reg_9_ ( .D(1'b0), .SETB(n206), .RSTB(
        n_sram_raddr_a4[9]), .CLK(net24315), .Q(sram_raddr_a4[9]) );
  DFFSSRX1_HVT sram_raddr_a4_reg_8_ ( .D(1'b0), .SETB(n198), .RSTB(
        n_sram_raddr_a4[8]), .CLK(net24315), .Q(sram_raddr_a4[8]) );
  DFFSSRX1_HVT sram_raddr_a4_reg_7_ ( .D(1'b0), .SETB(n194), .RSTB(
        n_sram_raddr_a4[7]), .CLK(net24315), .Q(sram_raddr_a4[7]) );
  DFFSSRX1_HVT sram_raddr_a4_reg_6_ ( .D(1'b0), .SETB(n200), .RSTB(
        n_sram_raddr_a4[6]), .CLK(net24315), .Q(sram_raddr_a4[6]), .QN(n353)
         );
  DFFSSRX1_HVT sram_raddr_a4_reg_5_ ( .D(1'b0), .SETB(n196), .RSTB(
        n_sram_raddr_a4[5]), .CLK(net24315), .Q(sram_raddr_a4[5]), .QN(n404)
         );
  DFFSSRX1_HVT sram_raddr_a4_reg_4_ ( .D(1'b0), .SETB(n182), .RSTB(
        n_sram_raddr_a4[4]), .CLK(net24315), .Q(sram_raddr_a4[4]), .QN(n246)
         );
  DFFSSRX1_HVT sram_raddr_a4_reg_3_ ( .D(1'b0), .SETB(n207), .RSTB(
        n_sram_raddr_a4[3]), .CLK(net24315), .Q(sram_raddr_a4[3]), .QN(n290)
         );
  DFFSSRX1_HVT sram_raddr_a4_reg_2_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_a4[2]), .CLK(net24315), .Q(sram_raddr_a4[2]), .QN(n235)
         );
  DFFSSRX1_HVT sram_raddr_a4_reg_1_ ( .D(1'b0), .SETB(n206), .RSTB(
        n_sram_raddr_a4[1]), .CLK(net24315), .Q(sram_raddr_a4[1]), .QN(n298)
         );
  DFFSSRX1_HVT sram_raddr_a4_reg_0_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_a4[0]), .CLK(net24315), .Q(sram_raddr_a4[0]), .QN(n396)
         );
  DFFSSRX1_HVT sram_raddr_a5_reg_9_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_a5[9]), .CLK(net25642), .Q(sram_raddr_a5[9]), .QN(n442)
         );
  DFFSSRX1_HVT sram_raddr_a5_reg_8_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_a5[8]), .CLK(net25642), .Q(sram_raddr_a5[8]) );
  DFFSSRX1_HVT sram_raddr_a5_reg_7_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_raddr_a5[7]), .CLK(net25642), .Q(sram_raddr_a5[7]), .QN(n352)
         );
  DFFSSRX1_HVT sram_raddr_a5_reg_6_ ( .D(1'b0), .SETB(n197), .RSTB(
        n_sram_raddr_a5[6]), .CLK(net25642), .Q(sram_raddr_a5[6]), .QN(n413)
         );
  DFFSSRX1_HVT sram_raddr_a5_reg_5_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_a5[5]), .CLK(net25642), .Q(sram_raddr_a5[5]), .QN(n350)
         );
  DFFSSRX1_HVT sram_raddr_a5_reg_4_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_a5[4]), .CLK(net25642), .Q(sram_raddr_a5[4]), .QN(n412)
         );
  DFFSSRX1_HVT sram_raddr_a5_reg_3_ ( .D(1'b0), .SETB(n206), .RSTB(
        n_sram_raddr_a5[3]), .CLK(net25642), .Q(sram_raddr_a5[3]), .QN(n278)
         );
  DFFSSRX1_HVT sram_raddr_a5_reg_2_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_a5[2]), .CLK(net25642), .Q(sram_raddr_a5[2]), .QN(n411)
         );
  DFFSSRX1_HVT sram_raddr_a5_reg_1_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_a5[1]), .CLK(net25642), .Q(sram_raddr_a5[1]) );
  DFFSSRX1_HVT sram_raddr_a5_reg_0_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_a5[0]), .CLK(net25642), .Q(sram_raddr_a5[0]), .QN(n394)
         );
  DFFSSRX1_HVT sram_raddr_a6_reg_9_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_raddr_a6[9]), .CLK(net26972), .Q(sram_raddr_a6[9]) );
  DFFSSRX1_HVT sram_raddr_a6_reg_8_ ( .D(1'b0), .SETB(n184), .RSTB(
        n_sram_raddr_a6[8]), .CLK(net26972), .Q(sram_raddr_a6[8]) );
  DFFSSRX1_HVT sram_raddr_a6_reg_7_ ( .D(1'b0), .SETB(n207), .RSTB(
        n_sram_raddr_a6[7]), .CLK(net26972), .Q(sram_raddr_a6[7]) );
  DFFSSRX1_HVT sram_raddr_a6_reg_6_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_a6[6]), .CLK(net26972), .Q(sram_raddr_a6[6]), .QN(n452)
         );
  DFFSSRX1_HVT sram_raddr_a6_reg_5_ ( .D(1'b0), .SETB(n206), .RSTB(
        n_sram_raddr_a6[5]), .CLK(net26972), .Q(sram_raddr_a6[5]) );
  DFFSSRX1_HVT sram_raddr_a6_reg_4_ ( .D(1'b0), .SETB(n197), .RSTB(
        n_sram_raddr_a6[4]), .CLK(net26972), .Q(sram_raddr_a6[4]) );
  DFFSSRX1_HVT sram_raddr_a6_reg_3_ ( .D(1'b0), .SETB(n193), .RSTB(
        n_sram_raddr_a6[3]), .CLK(net26972), .Q(sram_raddr_a6[3]) );
  DFFSSRX1_HVT sram_raddr_a6_reg_2_ ( .D(1'b0), .SETB(n199), .RSTB(
        n_sram_raddr_a6[2]), .CLK(net26972), .Q(sram_raddr_a6[2]), .QN(n443)
         );
  DFFSSRX1_HVT sram_raddr_a6_reg_1_ ( .D(1'b0), .SETB(n195), .RSTB(
        n_sram_raddr_a6[1]), .CLK(net26972), .Q(sram_raddr_a6[1]) );
  DFFSSRX1_HVT sram_raddr_a6_reg_0_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_a6[0]), .CLK(net26972), .Q(sram_raddr_a6[0]), .QN(n295)
         );
  DFFSSRX1_HVT sram_raddr_b7_reg_9_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_b7[9]), .CLK(net27506), .Q(sram_raddr_b7[9]), .QN(n372)
         );
  DFFSSRX1_HVT sram_raddr_b7_reg_8_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_b7[8]), .CLK(net27506), .Q(sram_raddr_b7[8]), .QN(n391)
         );
  DFFSSRX1_HVT sram_raddr_b7_reg_7_ ( .D(1'b0), .SETB(n206), .RSTB(
        n_sram_raddr_b7[7]), .CLK(net27506), .Q(sram_raddr_b7[7]), .QN(n347)
         );
  DFFSSRX1_HVT sram_raddr_b7_reg_6_ ( .D(1'b0), .SETB(n198), .RSTB(
        n_sram_raddr_b7[6]), .CLK(net27506), .Q(sram_raddr_b7[6]) );
  DFFSSRX1_HVT sram_raddr_b7_reg_5_ ( .D(1'b0), .SETB(n194), .RSTB(
        n_sram_raddr_b7[5]), .CLK(net27506), .Q(sram_raddr_b7[5]), .QN(n364)
         );
  DFFSSRX1_HVT sram_raddr_b7_reg_4_ ( .D(1'b0), .SETB(n200), .RSTB(
        n_sram_raddr_b7[4]), .CLK(net27506), .Q(sram_raddr_b7[4]), .QN(n281)
         );
  DFFSSRX1_HVT sram_raddr_b7_reg_3_ ( .D(1'b0), .SETB(n196), .RSTB(
        n_sram_raddr_b7[3]), .CLK(net27506), .Q(sram_raddr_b7[3]), .QN(n382)
         );
  DFFSSRX1_HVT sram_raddr_b7_reg_2_ ( .D(1'b0), .SETB(n183), .RSTB(
        n_sram_raddr_b7[2]), .CLK(net27506), .Q(sram_raddr_b7[2]), .QN(n240)
         );
  DFFSSRX1_HVT sram_raddr_b7_reg_1_ ( .D(1'b0), .SETB(n207), .RSTB(
        n_sram_raddr_b7[1]), .CLK(net27506), .Q(sram_raddr_b7[1]) );
  DFFSSRX1_HVT sram_raddr_b7_reg_0_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_b7[0]), .CLK(net27506), .Q(sram_raddr_b7[0]), .QN(n398)
         );
  DFFSSRX1_HVT sram_raddr_b8_reg_9_ ( .D(1'b0), .SETB(n206), .RSTB(
        n_sram_raddr_b8[9]), .CLK(net28021), .Q(sram_raddr_b8[9]), .QN(n374)
         );
  DFFSSRX1_HVT sram_raddr_b8_reg_8_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_b8[8]), .CLK(net28021), .Q(sram_raddr_b8[8]), .QN(n359)
         );
  DFFSSRX1_HVT sram_raddr_b8_reg_7_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_b8[7]), .CLK(net28021), .Q(sram_raddr_b8[7]), .QN(n275)
         );
  DFFSSRX1_HVT sram_raddr_b8_reg_6_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_b8[6]), .CLK(net28021), .Q(sram_raddr_b8[6]) );
  DFFSSRX1_HVT sram_raddr_b8_reg_5_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_raddr_b8[5]), .CLK(net28021), .Q(sram_raddr_b8[5]), .QN(n342)
         );
  DFFSSRX1_HVT sram_raddr_b8_reg_4_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_b8[4]), .CLK(net28021), .Q(sram_raddr_b8[4]), .QN(n381)
         );
  DFFSSRX1_HVT sram_raddr_b8_reg_3_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_b8[3]), .CLK(net28021), .Q(sram_raddr_b8[3]), .QN(n287)
         );
  DFFSSRX1_HVT sram_raddr_b8_reg_2_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_b8[2]), .CLK(net28021), .Q(sram_raddr_b8[2]), .QN(n241)
         );
  DFFSSRX1_HVT sram_raddr_b8_reg_1_ ( .D(1'b0), .SETB(n206), .RSTB(
        n_sram_raddr_b8[1]), .CLK(net28021), .Q(sram_raddr_b8[1]) );
  DFFSSRX1_HVT sram_raddr_b8_reg_0_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_b8[0]), .CLK(net28021), .Q(sram_raddr_b8[0]), .QN(n399)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_9_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_b0[9]), .CLK(net28536), .Q(sram_raddr_b0[9]), .QN(n401)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_8_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_b0[8]), .CLK(net28536), .Q(sram_raddr_b0[8]), .QN(n346)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_7_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_raddr_b0[7]), .CLK(net28536), .Q(sram_raddr_b0[7]), .QN(n269)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_6_ ( .D(1'b0), .SETB(n182), .RSTB(
        n_sram_raddr_b0[6]), .CLK(net28536), .Q(sram_raddr_b0[6]), .QN(n339)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_5_ ( .D(1'b0), .SETB(n207), .RSTB(
        n_sram_raddr_b0[5]), .CLK(net28536), .Q(sram_raddr_b0[5]), .QN(n340)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_4_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_b0[4]), .CLK(net28536), .Q(sram_raddr_b0[4]), .QN(n256)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_3_ ( .D(1'b0), .SETB(n206), .RSTB(
        n_sram_raddr_b0[3]), .CLK(net28536), .Q(sram_raddr_b0[3]), .QN(n379)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_2_ ( .D(1'b0), .SETB(n197), .RSTB(
        n_sram_raddr_b0[2]), .CLK(net28536), .Q(sram_raddr_b0[2]), .QN(n284)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_1_ ( .D(1'b0), .SETB(n193), .RSTB(
        n_sram_raddr_b0[1]), .CLK(net28536), .Q(sram_raddr_b0[1]), .QN(n322)
         );
  DFFSSRX1_HVT sram_raddr_b0_reg_0_ ( .D(1'b0), .SETB(n199), .RSTB(
        n_sram_raddr_b0[0]), .CLK(net28536), .Q(sram_raddr_b0[0]), .QN(n242)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_9_ ( .D(1'b0), .SETB(n195), .RSTB(
        n_sram_raddr_b1[9]), .CLK(net29051), .Q(sram_raddr_b1[9]), .QN(n377)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_8_ ( .D(1'b0), .SETB(n194), .RSTB(
        n_sram_raddr_b1[8]), .CLK(net29051), .Q(sram_raddr_b1[8]), .QN(n272)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_7_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_b1[7]), .CLK(net29051), .Q(sram_raddr_b1[7]), .QN(n333)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_6_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_b1[6]), .CLK(net29051), .Q(sram_raddr_b1[6]), .QN(n344)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_5_ ( .D(1'b0), .SETB(n206), .RSTB(
        n_sram_raddr_b1[5]), .CLK(net29051), .Q(sram_raddr_b1[5]), .QN(n270)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_4_ ( .D(1'b0), .SETB(n198), .RSTB(
        n_sram_raddr_b1[4]), .CLK(net29051), .Q(sram_raddr_b1[4]), .QN(n316)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_3_ ( .D(1'b0), .SETB(n194), .RSTB(
        n_sram_raddr_b1[3]), .CLK(net29051), .Q(sram_raddr_b1[3]), .QN(n386)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_2_ ( .D(1'b0), .SETB(n200), .RSTB(
        n_sram_raddr_b1[2]), .CLK(net29051), .Q(sram_raddr_b1[2]), .QN(n277)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_1_ ( .D(1'b0), .SETB(n196), .RSTB(
        n_sram_raddr_b1[1]), .CLK(net29051), .Q(sram_raddr_b1[1]), .QN(n323)
         );
  DFFSSRX1_HVT sram_raddr_b1_reg_0_ ( .D(1'b0), .SETB(n184), .RSTB(
        n_sram_raddr_b1[0]), .CLK(net29051), .Q(sram_raddr_b1[0]), .QN(n243)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_9_ ( .D(1'b0), .SETB(n207), .RSTB(
        n_sram_raddr_b2[9]), .CLK(net29566), .Q(sram_raddr_b2[9]), .QN(n419)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_8_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_b2[8]), .CLK(net29566), .Q(sram_raddr_b2[8]), .QN(n360)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_7_ ( .D(1'b0), .SETB(n206), .RSTB(
        n_sram_raddr_b2[7]), .CLK(net29566), .Q(sram_raddr_b2[7]), .QN(n267)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_6_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_b2[6]), .CLK(net29566), .Q(sram_raddr_b2[6]), .QN(n337)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_5_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_b2[5]), .CLK(net29566), .Q(sram_raddr_b2[5]), .QN(n334)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_4_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_b2[4]), .CLK(net29566), .Q(sram_raddr_b2[4]), .QN(n255)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_3_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_raddr_b2[3]), .CLK(net29566), .Q(sram_raddr_b2[3]), .QN(n406)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_2_ ( .D(1'b0), .SETB(n196), .RSTB(
        n_sram_raddr_b2[2]), .CLK(net29566), .Q(sram_raddr_b2[2]), .QN(n354)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_1_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_b2[1]), .CLK(net29566), .Q(sram_raddr_b2[1]), .QN(n325)
         );
  DFFSSRX1_HVT sram_raddr_b2_reg_0_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_b2[0]), .CLK(net29566), .Q(sram_raddr_b2[0]), .QN(n260)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_9_ ( .D(1'b0), .SETB(n206), .RSTB(
        n_sram_raddr_b3[9]), .CLK(net30081), .Q(sram_raddr_b3[9]), .QN(n361)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_8_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_b3[8]), .CLK(net30081), .Q(sram_raddr_b3[8]), .QN(n273)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_7_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_b3[7]), .CLK(net30081), .Q(sram_raddr_b3[7]), .QN(n388)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_6_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_b3[6]), .CLK(net30081), .Q(sram_raddr_b3[6]), .QN(n358)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_5_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_raddr_b3[5]), .CLK(net30081), .Q(sram_raddr_b3[5]), .QN(n268)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_4_ ( .D(1'b0), .SETB(n183), .RSTB(
        n_sram_raddr_b3[4]), .CLK(net30081), .Q(sram_raddr_b3[4]), .QN(n335)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_3_ ( .D(1'b0), .SETB(n207), .RSTB(
        n_sram_raddr_b3[3]), .CLK(net30081), .Q(sram_raddr_b3[3]), .QN(n343)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_2_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_b3[2]), .CLK(net30081), .Q(sram_raddr_b3[2]), .QN(n315)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_1_ ( .D(1'b0), .SETB(n206), .RSTB(
        n_sram_raddr_b3[1]), .CLK(net30081), .Q(sram_raddr_b3[1]), .QN(n324)
         );
  DFFSSRX1_HVT sram_raddr_b3_reg_0_ ( .D(1'b0), .SETB(n197), .RSTB(
        n_sram_raddr_b3[0]), .CLK(net30081), .Q(sram_raddr_b3[0]), .QN(n258)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_9_ ( .D(1'b0), .SETB(n193), .RSTB(
        n_sram_raddr_b4[9]), .CLK(net30596), .Q(sram_raddr_b4[9]), .QN(n351)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_8_ ( .D(1'b0), .SETB(n199), .RSTB(
        n_sram_raddr_b4[8]), .CLK(net30596), .Q(sram_raddr_b4[8]), .QN(n345)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_7_ ( .D(1'b0), .SETB(n195), .RSTB(
        n_sram_raddr_b4[7]), .CLK(net30596), .Q(sram_raddr_b4[7]), .QN(n332)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_6_ ( .D(1'b0), .SETB(n195), .RSTB(
        n_sram_raddr_b4[6]), .CLK(net30596), .Q(sram_raddr_b4[6]), .QN(n387)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_5_ ( .D(1'b0), .SETB(n208), .RSTB(
        n_sram_raddr_b4[5]), .CLK(net30596), .Q(sram_raddr_b4[5]), .QN(n276)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_4_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_b4[4]), .CLK(net30596), .Q(sram_raddr_b4[4]), .QN(n357)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_3_ ( .D(1'b0), .SETB(n206), .RSTB(
        n_sram_raddr_b4[3]), .CLK(net30596), .Q(sram_raddr_b4[3]), .QN(n336)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_2_ ( .D(1'b0), .SETB(n198), .RSTB(
        n_sram_raddr_b4[2]), .CLK(net30596), .Q(sram_raddr_b4[2]), .QN(n314)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_1_ ( .D(1'b0), .SETB(n194), .RSTB(
        n_sram_raddr_b4[1]), .CLK(net30596), .Q(sram_raddr_b4[1]), .QN(n326)
         );
  DFFSSRX1_HVT sram_raddr_b4_reg_0_ ( .D(1'b0), .SETB(n200), .RSTB(
        n_sram_raddr_b4[0]), .CLK(net30596), .Q(sram_raddr_b4[0]), .QN(n259)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_9_ ( .D(1'b0), .SETB(n196), .RSTB(
        n_sram_raddr_b5[9]), .CLK(net31111), .Q(sram_raddr_b5[9]), .QN(n348)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_8_ ( .D(1'b0), .SETB(n198), .RSTB(
        n_sram_raddr_b5[8]), .CLK(net31111), .Q(sram_raddr_b5[8]), .QN(n286)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_7_ ( .D(1'b0), .SETB(n207), .RSTB(
        n_sram_raddr_b5[7]), .CLK(net31111), .Q(sram_raddr_b5[7]), .QN(n393)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_6_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_b5[6]), .CLK(net31111), .Q(sram_raddr_b5[6]), .QN(n365)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_5_ ( .D(1'b0), .SETB(n206), .RSTB(
        n_sram_raddr_b5[5]), .CLK(net31111), .Q(sram_raddr_b5[5]), .QN(n271)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_4_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_b5[4]), .CLK(net31111), .Q(sram_raddr_b5[4]), .QN(n341)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_3_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_b5[3]), .CLK(net31111), .Q(sram_raddr_b5[3]), .QN(n384)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_2_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_b5[2]), .CLK(net31111), .Q(sram_raddr_b5[2]), .QN(n313)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_1_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_raddr_b5[1]), .CLK(net31111), .Q(sram_raddr_b5[1]), .QN(n327)
         );
  DFFSSRX1_HVT sram_raddr_b5_reg_0_ ( .D(1'b0), .SETB(n185), .RSTB(
        n_sram_raddr_b5[0]), .CLK(net31111), .Q(sram_raddr_b5[0]), .QN(n244)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_9_ ( .D(1'b0), .SETB(n182), .RSTB(
        n_sram_raddr_b6[9]), .CLK(net31626), .Q(sram_raddr_b6[9]), .QN(n373)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_8_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_b6[8]), .CLK(net31626), .Q(sram_raddr_b6[8]), .QN(n274)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_7_ ( .D(1'b0), .SETB(n206), .RSTB(
        n_sram_raddr_b6[7]), .CLK(net31626), .Q(sram_raddr_b6[7]), .QN(n338)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_6_ ( .D(1'b0), .SETB(n175), .RSTB(
        n_sram_raddr_b6[6]), .CLK(net31626), .Q(sram_raddr_b6[6]), .QN(n408)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_5_ ( .D(1'b0), .SETB(n177), .RSTB(
        n_sram_raddr_b6[5]), .CLK(net31626), .Q(sram_raddr_b6[5]), .QN(n363)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_4_ ( .D(1'b0), .SETB(n176), .RSTB(
        n_sram_raddr_b6[4]), .CLK(net31626), .Q(sram_raddr_b6[4]), .QN(n280)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_3_ ( .D(1'b0), .SETB(n174), .RSTB(
        n_sram_raddr_b6[3]), .CLK(net31626), .Q(sram_raddr_b6[3]), .QN(n389)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_2_ ( .D(1'b0), .SETB(n186), .RSTB(
        n_sram_raddr_b6[2]), .CLK(net31626), .Q(sram_raddr_b6[2]), .QN(n239)
         );
  DFFSSRX1_HVT sram_raddr_b6_reg_1_ ( .D(1'b0), .SETB(n183), .RSTB(
        n_sram_raddr_b6[1]), .CLK(net31626), .Q(sram_raddr_b6[1]) );
  DFFSSRX1_HVT sram_raddr_b6_reg_0_ ( .D(1'b0), .SETB(n210), .RSTB(
        n_sram_raddr_b6[0]), .CLK(net31626), .Q(sram_raddr_b6[0]), .QN(n397)
         );
  DFFSSRX1_HVT sram_write_enable_b7_reg ( .D(n_sram_write_enable_b7), .SETB(
        n181), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b7) );
  DFFSSRX1_HVT sram_write_enable_b8_reg ( .D(n_sram_write_enable_b8), .SETB(
        n181), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b8) );
  DFFSSRX1_HVT sram_write_enable_b0_reg ( .D(n_sram_write_enable_b0), .SETB(
        srstn), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b0) );
  DFFSSRX1_HVT sram_write_enable_b1_reg ( .D(n_sram_write_enable_b1), .SETB(
        n181), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b1) );
  DFFSSRX1_HVT sram_write_enable_b2_reg ( .D(n_sram_write_enable_b2), .SETB(
        n181), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b2) );
  DFFSSRX1_HVT sram_write_enable_b3_reg ( .D(n_sram_write_enable_b3), .SETB(
        srstn), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b3) );
  DFFSSRX1_HVT sram_write_enable_b4_reg ( .D(n_sram_write_enable_b4), .SETB(
        n181), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b4) );
  DFFSSRX1_HVT sram_write_enable_b5_reg ( .D(n_sram_write_enable_b5), .SETB(
        srstn), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b5) );
  DFFSSRX1_HVT sram_write_enable_b6_reg ( .D(n_sram_write_enable_b6), .SETB(
        n227), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_b6) );
  DFFSSRX1_HVT sram_write_enable_d3_reg ( .D(n_sram_write_enable_d3), .SETB(
        n181), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_d3) );
  DFFSSRX1_HVT sram_write_enable_d4_reg ( .D(n_sram_write_enable_d4), .SETB(
        srstn), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_d4) );
  DFFSSRX1_HVT sram_write_enable_c0_reg ( .D(n_sram_write_enable_c0), .SETB(
        n227), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_c0) );
  DFFSSRX1_HVT sram_write_enable_c1_reg ( .D(n_sram_write_enable_c1), .SETB(
        n181), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_c1) );
  DFFSSRX1_HVT sram_write_enable_c2_reg ( .D(n_sram_write_enable_c2), .SETB(
        srstn), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_c2) );
  DFFSSRX1_HVT sram_write_enable_c3_reg ( .D(n_sram_write_enable_c3), .SETB(
        n227), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_c3) );
  DFFSSRX1_HVT sram_write_enable_c4_reg ( .D(n_sram_write_enable_c4), .SETB(
        n181), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_c4) );
  DFFSSRX1_HVT sram_write_enable_d0_reg ( .D(n_sram_write_enable_d0), .SETB(
        srstn), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_d0) );
  DFFSSRX1_HVT sram_write_enable_d1_reg ( .D(n_sram_write_enable_d1), .SETB(
        n181), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_d1) );
  DFFSSRX1_HVT sram_write_enable_d2_reg ( .D(n_sram_write_enable_d2), .SETB(
        srstn), .RSTB(1'b1), .CLK(clk), .Q(sram_write_enable_d2) );
  DFFSSRX1_HVT state_reg_3_ ( .D(1'b0), .SETB(n184), .RSTB(n_state[3]), .CLK(
        clk), .Q(state[3]), .QN(n1023) );
  DFFSSRX1_HVT state_reg_2_ ( .D(1'b0), .SETB(n187), .RSTB(n_state[2]), .CLK(
        clk), .Q(state[2]), .QN(n1024) );
  AO221X1_HVT U3 ( .A1(1'b1), .A2(n1488), .A3(n1490), .A4(n375), .A5(n156), 
        .Y(n158) );
  AO221X1_HVT U4 ( .A1(1'b1), .A2(n1929), .A3(n1926), .A4(n168), .A5(n150), 
        .Y(n_sram_raddr_a4[8]) );
  AO221X1_HVT U5 ( .A1(1'b1), .A2(n1494), .A3(n1496), .A4(n376), .A5(n137), 
        .Y(n138) );
  AO221X1_HVT U6 ( .A1(1'b1), .A2(n1502), .A3(n409), .A4(n1503), .A5(n114), 
        .Y(n116) );
  AO221X1_HVT U7 ( .A1(1'b1), .A2(n1638), .A3(n436), .A4(n301), .A5(n108), .Y(
        n110) );
  AO222X1_HVT U8 ( .A1(sram_raddr_b7[7]), .A2(n231), .A3(n68), .A4(n1233), 
        .A5(1'b1), .A6(n73), .Y(n_sram_raddr_b7[7]) );
  AO221X1_HVT U9 ( .A1(1'b1), .A2(n908), .A3(n914), .A4(n277), .A5(n104), .Y(
        n1185) );
  AO221X1_HVT U10 ( .A1(1'b1), .A2(n1435), .A3(n407), .A4(n98), .A5(n99), .Y(
        n101) );
  AO221X1_HVT U11 ( .A1(1'b1), .A2(n1884), .A3(n1881), .A4(n1839), .A5(n95), 
        .Y(n_sram_raddr_a3[8]) );
  AO221X1_HVT U12 ( .A1(1'b1), .A2(n86), .A3(n1338), .A4(n1310), .A5(n89), .Y(
        n91) );
  AO221X1_HVT U13 ( .A1(1'b1), .A2(n1924), .A3(n1923), .A4(n168), .A5(n77), 
        .Y(n_sram_raddr_a4[7]) );
  AO222X1_HVT U14 ( .A1(sram_raddr_b7[5]), .A2(n230), .A3(n55), .A4(n1221), 
        .A5(1'b1), .A6(n61), .Y(n_sram_raddr_b7[5]) );
  AO222X1_HVT U15 ( .A1(sram_raddr_b8[7]), .A2(n232), .A3(n44), .A4(n1318), 
        .A5(1'b1), .A6(n50), .Y(n_sram_raddr_b8[7]) );
  AO22X1_HVT U16 ( .A1(n342), .A2(n1306), .A3(n1311), .A4(1'b1), .Y(n31) );
  OA221X1_HVT U17 ( .A1(1'b0), .A2(n1567), .A3(n1566), .A4(col[2]), .A5(n1565), 
        .Y(net22643) );
  OA221X1_HVT U18 ( .A1(1'b0), .A2(n541), .A3(row[2]), .A4(n540), .A5(n539), 
        .Y(n_row[2]) );
  OA221X1_HVT U19 ( .A1(1'b0), .A2(n1550), .A3(channel_cnt[1]), .A4(
        channel_cnt[0]), .A5(n1549), .Y(net22936) );
  OA221X1_HVT U20 ( .A1(1'b0), .A2(sram_raddr_weight[13]), .A3(
        sram_raddr_weight[12]), .A4(n1406), .A5(n203), .Y(n163) );
  OA221X1_HVT U21 ( .A1(1'b0), .A2(n1557), .A3(addr_change[0]), .A4(
        addr_change[1]), .A5(n1556), .Y(net22948) );
  OA221X1_HVT U22 ( .A1(1'b0), .A2(n1544), .A3(n1532), .A4(
        delay1_sram_waddr_d[8]), .A5(n1531), .Y(net22917) );
  OA221X1_HVT U23 ( .A1(1'b0), .A2(n586), .A3(n256), .A4(n622), .A5(n143), .Y(
        n145) );
  OA221X1_HVT U24 ( .A1(1'b0), .A2(n1262), .A3(sram_raddr_b1[6]), .A4(n929), 
        .A5(n938), .Y(n1226) );
  OA221X1_HVT U25 ( .A1(1'b0), .A2(n192), .A3(sram_raddr_b8[3]), .A4(n1277), 
        .A5(n1276), .Y(n993) );
  OA221X1_HVT U26 ( .A1(1'b0), .A2(n1557), .A3(addr_change[2]), .A4(n134), 
        .A5(n1555), .Y(net22947) );
  OA221X1_HVT U27 ( .A1(1'b0), .A2(n1544), .A3(n1534), .A4(
        delay1_sram_waddr_d[7]), .A5(n1533), .Y(net22918) );
  OA221X1_HVT U28 ( .A1(1'b0), .A2(n1557), .A3(addr_change[3]), .A4(n112), 
        .A5(n1554), .Y(net22946) );
  OA221X1_HVT U29 ( .A1(1'b0), .A2(n1544), .A3(n1536), .A4(
        delay1_sram_waddr_d[6]), .A5(n1535), .Y(net22919) );
  OA21X1_HVT U30 ( .A1(n1234), .A2(sram_raddr_b7[7]), .A3(n179), .Y(n68) );
  OA221X1_HVT U31 ( .A1(1'b0), .A2(n1470), .A3(n249), .A4(n296), .A5(n405), 
        .Y(n103) );
  OA221X1_HVT U32 ( .A1(1'b0), .A2(n1544), .A3(n1538), .A4(
        delay1_sram_waddr_d[5]), .A5(n1537), .Y(net22920) );
  OA221X1_HVT U33 ( .A1(1'b0), .A2(n1544), .A3(n1540), .A4(
        delay1_sram_waddr_d[4]), .A5(n1539), .Y(net22921) );
  OA221X1_HVT U34 ( .A1(1'b0), .A2(n1544), .A3(delay1_sram_waddr_d[3]), .A4(
        n75), .A5(n1541), .Y(net22922) );
  OA221X1_HVT U35 ( .A1(1'b0), .A2(n1544), .A3(delay1_sram_waddr_d[2]), .A4(
        n66), .A5(n1542), .Y(net22923) );
  OA21X1_HVT U36 ( .A1(n1215), .A2(sram_raddr_b7[5]), .A3(n223), .Y(n55) );
  OA221X1_HVT U37 ( .A1(1'b0), .A2(n1305), .A3(sram_raddr_b4[8]), .A4(n1368), 
        .A5(n949), .Y(n973) );
  OA221X1_HVT U38 ( .A1(1'b0), .A2(n1544), .A3(delay1_sram_waddr_d[0]), .A4(
        delay1_sram_waddr_d[1]), .A5(n1543), .Y(net22924) );
  OA221X1_HVT U39 ( .A1(1'b0), .A2(n1528), .A3(n1516), .A4(
        delay1_sram_waddr_c[8]), .A5(n1515), .Y(net22901) );
  OA21X1_HVT U40 ( .A1(n1319), .A2(sram_raddr_b8[7]), .A3(n222), .Y(n44) );
  OA221X1_HVT U41 ( .A1(1'b0), .A2(n695), .A3(sram_raddr_b1[8]), .A4(n1368), 
        .A5(n1305), .Y(n700) );
  OA221X1_HVT U42 ( .A1(1'b0), .A2(n1528), .A3(n1518), .A4(
        delay1_sram_waddr_c[7]), .A5(n1517), .Y(net22902) );
  OA221X1_HVT U43 ( .A1(1'b0), .A2(n1528), .A3(n1520), .A4(
        delay1_sram_waddr_c[6]), .A5(n1519), .Y(net22903) );
  OA221X1_HVT U44 ( .A1(1'b0), .A2(n1528), .A3(n1522), .A4(
        delay1_sram_waddr_c[5]), .A5(n1521), .Y(net22904) );
  OA221X1_HVT U45 ( .A1(1'b0), .A2(n1528), .A3(n1524), .A4(
        delay1_sram_waddr_c[4]), .A5(n1523), .Y(net22905) );
  OA221X1_HVT U46 ( .A1(1'b0), .A2(n1528), .A3(delay1_sram_waddr_c[3]), .A4(
        n25), .A5(n1525), .Y(net22906) );
  OA221X1_HVT U47 ( .A1(1'b0), .A2(n1401), .A3(n226), .A4(n362), .A5(n18), .Y(
        n1397) );
  OA221X1_HVT U48 ( .A1(1'b0), .A2(n1528), .A3(delay1_sram_waddr_c[2]), .A4(
        n17), .A5(n1526), .Y(net22907) );
  OA221X1_HVT U49 ( .A1(1'b0), .A2(n10), .A3(n173), .A4(n930), .A5(n934), .Y(
        n12) );
  OA221X1_HVT U50 ( .A1(1'b0), .A2(n1528), .A3(delay1_sram_waddr_c[0]), .A4(
        delay1_sram_waddr_c[1]), .A5(n1527), .Y(net22908) );
  INVX1_HVT U51 ( .A(n1833), .Y(n172) );
  INVX1_HVT U52 ( .A(n1268), .Y(n169) );
  INVX1_HVT U53 ( .A(n1322), .Y(n173) );
  INVX0_HVT U54 ( .A(n663), .Y(n1) );
  OA221X1_HVT U55 ( .A1(n1), .A2(col[0]), .A3(n1), .A4(n706), .A5(n664), .Y(n2) );
  OA22X1_HVT U56 ( .A1(n270), .A2(n2), .A3(n925), .A4(n224), .Y(n3) );
  NAND3X0_HVT U57 ( .A1(n924), .A2(n669), .A3(n3), .Y(n4) );
  NAND2X0_HVT U58 ( .A1(n913), .A2(n270), .Y(n5) );
  AND2X1_HVT U59 ( .A1(n5), .A2(n672), .Y(n6) );
  AO222X1_HVT U60 ( .A1(n4), .A2(n202), .A3(sram_raddr_b1[5]), .A4(n232), .A5(
        n188), .A6(n6), .Y(n_sram_raddr_b1[5]) );
  AND2X1_HVT U62 ( .A1(n669), .A2(n213), .Y(n8) );
  AO222X1_HVT U63 ( .A1(n706), .A2(n675), .A3(n706), .A4(n1200), .A5(n675), 
        .A6(n674), .Y(n9) );
  OA22X1_HVT U64 ( .A1(n344), .A2(n8), .A3(sram_raddr_b1[6]), .A4(n9), .Y(n10)
         );
  OA22X1_HVT U66 ( .A1(n344), .A2(n1305), .A3(n12), .A4(n219), .Y(n13) );
  NAND2X0_HVT U67 ( .A1(n672), .A2(n344), .Y(n14) );
  NAND3X0_HVT U68 ( .A1(n14), .A2(n683), .A3(n179), .Y(n15) );
  NAND2X0_HVT U69 ( .A1(n13), .A2(n15), .Y(n_sram_raddr_b1[6]) );
  INVX0_HVT U71 ( .A(n1527), .Y(n17) );
  NAND2X0_HVT U72 ( .A1(n1394), .A2(n1456), .Y(n18) );
  INVX0_HVT U74 ( .A(n566), .Y(n21) );
  NAND2X0_HVT U75 ( .A1(sram_raddr_b0[2]), .A2(n21), .Y(n22) );
  NAND3X0_HVT U76 ( .A1(n567), .A2(n812), .A3(n22), .Y(n23) );
  AO222X1_HVT U77 ( .A1(n23), .A2(n201), .A3(sram_raddr_b0[2]), .A4(n231), 
        .A5(n284), .A6(n222), .Y(n_sram_raddr_b0[2]) );
  INVX0_HVT U79 ( .A(n1526), .Y(n25) );
  OA22X1_HVT U80 ( .A1(n269), .A2(n609), .A3(n861), .A4(n173), .Y(n26) );
  NAND2X0_HVT U81 ( .A1(n269), .A2(n610), .Y(n27) );
  NAND3X0_HVT U82 ( .A1(n27), .A2(n26), .A3(n859), .Y(n28) );
  AO222X1_HVT U83 ( .A1(n28), .A2(n203), .A3(n613), .A4(sram_raddr_b0[7]), 
        .A5(n269), .A6(n630), .Y(n_sram_raddr_b0[7]) );
  INVX0_HVT U85 ( .A(n179), .Y(n30) );
  OA21X1_HVT U86 ( .A1(n1300), .A2(col[1]), .A3(n214), .Y(n32) );
  OA22X1_HVT U87 ( .A1(n342), .A2(n32), .A3(n1301), .A4(n1307), .Y(n33) );
  NAND2X0_HVT U88 ( .A1(n1338), .A2(n1302), .Y(n34) );
  AO221X1_HVT U89 ( .A1(n1312), .A2(n1303), .A3(n1312), .A4(n271), .A5(n225), 
        .Y(n35) );
  AND4X1_HVT U90 ( .A1(n33), .A2(n1304), .A3(n34), .A4(n35), .Y(n36) );
  OAI222X1_HVT U91 ( .A1(n30), .A2(n31), .A3(n36), .A4(n226), .A5(n342), .A6(
        n1305), .Y(n_sram_raddr_b8[5]) );
  NAND4X0_HVT U95 ( .A1(row[0]), .A2(col[2]), .A3(row[1]), .A4(col[3]), .Y(n40) );
  NAND3X0_HVT U96 ( .A1(row[0]), .A2(n233), .A3(n534), .Y(n41) );
  NAND3X0_HVT U97 ( .A1(n533), .A2(n40), .A3(n41), .Y(n42) );
  AO221X1_HVT U98 ( .A1(n42), .A2(n253), .A3(n42), .A4(n552), .A5(n1571), .Y(
        n43) );
  NAND3X0_HVT U99 ( .A1(row[3]), .A2(n539), .A3(n43), .Y(n535) );
  OA21X1_HVT U100 ( .A1(n393), .A2(n1313), .A3(n1321), .Y(n45) );
  AO22X1_HVT U101 ( .A1(n1324), .A2(n213), .A3(n211), .A4(col[1]), .Y(n46) );
  OA22X1_HVT U102 ( .A1(n173), .A2(n45), .A3(n275), .A4(n46), .Y(n47) );
  NAND3X0_HVT U103 ( .A1(n275), .A2(n1320), .A3(n1324), .Y(n48) );
  NAND3X0_HVT U104 ( .A1(n47), .A2(n1314), .A3(n48), .Y(n49) );
  OA221X1_HVT U105 ( .A1(n49), .A2(n1315), .A3(n49), .A4(n1338), .A5(n205), 
        .Y(n50) );
  OA21X1_HVT U110 ( .A1(n1212), .A2(n276), .A3(n1216), .Y(n56) );
  AO22X1_HVT U111 ( .A1(n1217), .A2(n212), .A3(n213), .A4(col[0]), .Y(n57) );
  OA22X1_HVT U112 ( .A1(n224), .A2(n56), .A3(n364), .A4(n57), .Y(n58) );
  NAND3X0_HVT U113 ( .A1(n364), .A2(n1228), .A3(n1217), .Y(n59) );
  NAND3X0_HVT U114 ( .A1(n58), .A2(n1213), .A3(n59), .Y(n60) );
  OA221X1_HVT U115 ( .A1(n60), .A2(n1214), .A3(n60), .A4(n1250), .A5(n204), 
        .Y(n61) );
  INVX0_HVT U120 ( .A(n1543), .Y(n66) );
  OA21X1_HVT U121 ( .A1(n912), .A2(n914), .A3(n1262), .Y(n67) );
  OA21X1_HVT U122 ( .A1(sram_raddr_b1[3]), .A2(n908), .A3(n67), .Y(n1195) );
  OA21X1_HVT U123 ( .A1(n332), .A2(n1229), .A3(n1235), .Y(n69) );
  AO22X1_HVT U124 ( .A1(n1246), .A2(n211), .A3(n212), .A4(col[0]), .Y(n70) );
  OA22X1_HVT U125 ( .A1(n225), .A2(n69), .A3(n347), .A4(n70), .Y(n71) );
  NAND3X0_HVT U126 ( .A1(n1230), .A2(n71), .A3(n1237), .Y(n72) );
  OA221X1_HVT U127 ( .A1(n72), .A2(n1231), .A3(n72), .A4(n1250), .A5(n203), 
        .Y(n73) );
  INVX0_HVT U129 ( .A(n1542), .Y(n75) );
  AO22X1_HVT U131 ( .A1(n1935), .A2(sram_raddr_a4[7]), .A3(n1804), .A4(n1798), 
        .Y(n77) );
  OA222X1_HVT U133 ( .A1(sram_raddr_weight[11]), .A2(sram_raddr_weight[9]), 
        .A3(sram_raddr_weight[11]), .A4(sram_raddr_weight[10]), .A5(
        sram_raddr_weight[11]), .A6(n1418), .Y(n79) );
  AND2X1_HVT U134 ( .A1(n1410), .A2(n1456), .Y(n80) );
  OA21X1_HVT U135 ( .A1(sram_raddr_weight[10]), .A2(n1413), .A3(
        sram_raddr_weight[11]), .Y(n81) );
  AO222X1_HVT U136 ( .A1(n79), .A2(n80), .A3(n81), .A4(n205), .A5(n1411), .A6(
        n202), .Y(net22726) );
  NAND2X0_HVT U137 ( .A1(n668), .A2(n281), .Y(n82) );
  NAND2X0_HVT U138 ( .A1(n82), .A2(sram_raddr_b7[5]), .Y(n83) );
  NAND2X0_HVT U139 ( .A1(n83), .A2(n671), .Y(n1214) );
  NAND4X0_HVT U140 ( .A1(state[0]), .A2(n1024), .A3(state[3]), .A4(n251), .Y(
        n84) );
  AO21X1_HVT U141 ( .A1(n1391), .A2(n84), .A3(n1070), .Y(net22775) );
  AND2X1_HVT U142 ( .A1(n1324), .A2(n1320), .Y(n85) );
  AO222X1_HVT U143 ( .A1(n85), .A2(sram_raddr_b8[6]), .A3(n85), .A4(n1307), 
        .A5(sram_raddr_b8[6]), .A6(n1308), .Y(n86) );
  INVX0_HVT U144 ( .A(n1312), .Y(n87) );
  AO221X1_HVT U145 ( .A1(n1312), .A2(sram_raddr_b5[6]), .A3(n87), .A4(n365), 
        .A5(n225), .Y(n88) );
  NAND2X0_HVT U146 ( .A1(n1309), .A2(n88), .Y(n89) );
  OR2X1_HVT U148 ( .A1(sram_raddr_b8[6]), .A2(n1311), .Y(n92) );
  AND2X1_HVT U149 ( .A1(n222), .A2(n1316), .Y(n93) );
  AO222X1_HVT U150 ( .A1(n91), .A2(n201), .A3(n92), .A4(n93), .A5(n231), .A6(
        sram_raddr_b8[6]), .Y(n_sram_raddr_b8[6]) );
  AO22X1_HVT U152 ( .A1(n1888), .A2(sram_raddr_a3[8]), .A3(n1770), .A4(n1766), 
        .Y(n95) );
  AO221X1_HVT U154 ( .A1(n1434), .A2(n1440), .A3(n1434), .A4(n407), .A5(n226), 
        .Y(n97) );
  NAND2X0_HVT U155 ( .A1(sram_raddr_weight[5]), .A2(n1439), .Y(n98) );
  INVX0_HVT U156 ( .A(n1456), .Y(n99) );
  NAND3X0_HVT U158 ( .A1(n283), .A2(n97), .A3(n101), .Y(net22789) );
  OA21X1_HVT U160 ( .A1(write_row_conv1[2]), .A2(n1061), .A3(n103), .Y(n1349)
         );
  INVX0_HVT U161 ( .A(n1262), .Y(n104) );
  OA22X1_HVT U164 ( .A1(n436), .A2(n1893), .A3(n189), .A4(n1775), .Y(n107) );
  INVX0_HVT U165 ( .A(n1665), .Y(n108) );
  NAND3X0_HVT U167 ( .A1(n107), .A2(n1776), .A3(n110), .Y(n_sram_raddr_a1[1])
         );
  INVX0_HVT U169 ( .A(n1555), .Y(n112) );
  INVX0_HVT U171 ( .A(n1507), .Y(n114) );
  INVX0_HVT U173 ( .A(n1504), .Y(n117) );
  AO221X1_HVT U174 ( .A1(n1500), .A2(n409), .A3(n1500), .A4(n117), .A5(n1499), 
        .Y(n118) );
  NAND2X0_HVT U175 ( .A1(n116), .A2(n118), .Y(net22884) );
  AO21X1_HVT U176 ( .A1(channel_cnt[2]), .A2(n1548), .A3(channel_cnt[3]), .Y(
        n119) );
  AND3X1_HVT U177 ( .A1(n1550), .A2(n1547), .A3(n119), .Y(net22934) );
  NAND2X0_HVT U178 ( .A1(n590), .A2(n280), .Y(n120) );
  NAND2X0_HVT U179 ( .A1(n120), .A2(sram_raddr_b6[5]), .Y(n121) );
  NAND2X0_HVT U180 ( .A1(n121), .A2(n592), .Y(n1123) );
  INVX0_HVT U181 ( .A(n1195), .Y(n122) );
  OA21X1_HVT U182 ( .A1(n909), .A2(n970), .A3(n122), .Y(n123) );
  AO21X1_HVT U183 ( .A1(n907), .A2(n214), .A3(n336), .Y(n124) );
  NAND3X0_HVT U184 ( .A1(n336), .A2(n1228), .A3(sram_raddr_b4[2]), .Y(n125) );
  NAND4X0_HVT U185 ( .A1(n910), .A2(n123), .A3(n124), .A4(n125), .Y(n126) );
  NAND2X0_HVT U186 ( .A1(n314), .A2(n223), .Y(n127) );
  NAND2X0_HVT U187 ( .A1(n1305), .A2(n127), .Y(n128) );
  AND2X1_HVT U188 ( .A1(n336), .A2(sram_raddr_b4[2]), .Y(n129) );
  AO222X1_HVT U189 ( .A1(n126), .A2(n1558), .A3(n128), .A4(sram_raddr_b4[3]), 
        .A5(n188), .A6(n129), .Y(n_sram_raddr_b4[3]) );
  NAND2X0_HVT U190 ( .A1(n1922), .A2(sram_raddr_a4[7]), .Y(n130) );
  NAND2X0_HVT U191 ( .A1(n1925), .A2(n130), .Y(n131) );
  AO222X1_HVT U192 ( .A1(n131), .A2(n1975), .A3(n1932), .A4(n1923), .A5(
        sram_raddr_a7[7]), .A6(n1935), .Y(n132) );
  OR2X1_HVT U193 ( .A1(n1924), .A2(n132), .Y(n_sram_raddr_a7[7]) );
  INVX0_HVT U195 ( .A(n1556), .Y(n134) );
  INVX0_HVT U198 ( .A(n1507), .Y(n137) );
  AO221X1_HVT U199 ( .A1(n1493), .A2(n376), .A3(n1493), .A4(n1495), .A5(n1499), 
        .Y(n139) );
  NAND2X0_HVT U200 ( .A1(n138), .A2(n139), .Y(net22878) );
  AOI22X1_HVT U201 ( .A1(n1996), .A2(n1998), .A3(n2002), .A4(n1997), .Y(n140)
         );
  OAI221X1_HVT U202 ( .A1(n140), .A2(n1996), .A3(n140), .A4(n1997), .A5(n1662), 
        .Y(n_box_sel_1_) );
  NAND2X0_HVT U205 ( .A1(n585), .A2(n1150), .Y(n143) );
  OA22X1_HVT U207 ( .A1(n340), .A2(n145), .A3(n837), .A4(n225), .Y(n146) );
  NAND3X0_HVT U208 ( .A1(n840), .A2(n593), .A3(n146), .Y(n147) );
  NAND2X0_HVT U209 ( .A1(n597), .A2(n340), .Y(n148) );
  AND2X1_HVT U210 ( .A1(n148), .A2(n596), .Y(n149) );
  AO222X1_HVT U211 ( .A1(n147), .A2(n201), .A3(sram_raddr_b0[5]), .A4(n230), 
        .A5(n222), .A6(n149), .Y(n_sram_raddr_b0[5]) );
  AO22X1_HVT U212 ( .A1(n1935), .A2(sram_raddr_a4[8]), .A3(n1804), .A4(n1800), 
        .Y(n150) );
  INVX0_HVT U214 ( .A(n1586), .Y(n152) );
  OR2X1_HVT U215 ( .A1(n1582), .A2(sram_raddr_a0[2]), .Y(n153) );
  AO222X1_HVT U216 ( .A1(n152), .A2(n153), .A3(n1975), .A4(n1739), .A5(n521), 
        .A6(n1852), .Y(n_sram_raddr_a0[2]) );
  INVX0_HVT U219 ( .A(n1507), .Y(n156) );
  AO221X1_HVT U221 ( .A1(n1487), .A2(n375), .A3(n1487), .A4(n1489), .A5(n1499), 
        .Y(n159) );
  NAND2X0_HVT U222 ( .A1(n158), .A2(n159), .Y(net22872) );
  INVX0_HVT U223 ( .A(n1404), .Y(n160) );
  OA221X1_HVT U224 ( .A1(sram_raddr_weight[13]), .A2(sram_raddr_weight[12]), 
        .A3(sram_raddr_weight[13]), .A4(n1407), .A5(n160), .Y(n161) );
  OR3X1_HVT U226 ( .A1(n1405), .A2(n161), .A3(n163), .Y(net22712) );
  AND3X1_HVT U230 ( .A1(n1384), .A2(weight_cnt[0]), .A3(weight_cnt[1]), .Y(
        n167) );
  OA21X1_HVT U231 ( .A1(n167), .A2(weight_cnt[2]), .A3(n1374), .Y(
        n_weight_cnt[2]) );
  INVX1_HVT U232 ( .A(n229), .Y(n209) );
  INVX4_HVT U233 ( .A(srstn), .Y(n180) );
  INVX4_HVT U234 ( .A(n180), .Y(n181) );
  NBUFFX2_HVT U235 ( .A(n227), .Y(n228) );
  INVX1_HVT U236 ( .A(n1070), .Y(n227) );
  INVX1_HVT U237 ( .A(srstn), .Y(n1070) );
  INVX1_HVT U238 ( .A(n189), .Y(n170) );
  INVX1_HVT U239 ( .A(n1943), .Y(n168) );
  INVX1_HVT U240 ( .A(mode[0]), .Y(n523) );
  INVX1_HVT U241 ( .A(n1847), .Y(n477) );
  NOR2X0_HVT U242 ( .A1(n1390), .A2(n1389), .Y(net22648) );
  INVX0_HVT U243 ( .A(n1936), .Y(n468) );
  INVX0_HVT U244 ( .A(n209), .Y(n185) );
  INVX1_HVT U245 ( .A(n224), .Y(n178) );
  INVX0_HVT U246 ( .A(n1659), .Y(n1660) );
  NOR2X0_HVT U247 ( .A1(n1483), .A2(n1501), .Y(n1486) );
  INVX1_HVT U248 ( .A(n1670), .Y(n1671) );
  NOR2X1_HVT U249 ( .A1(n352), .A2(n1714), .Y(n1726) );
  NOR2X1_HVT U250 ( .A1(n1880), .A2(sram_raddr_a3[8]), .Y(n1885) );
  INVX2_HVT U251 ( .A(n1975), .Y(n171) );
  INVX0_HVT U252 ( .A(n1652), .Y(n1653) );
  INVX0_HVT U253 ( .A(n903), .Y(n904) );
  INVX1_HVT U254 ( .A(n673), .Y(n675) );
  INVX1_HVT U255 ( .A(n1221), .Y(n1222) );
  INVX1_HVT U256 ( .A(n1111), .Y(n1109) );
  INVX1_HVT U257 ( .A(n1558), .Y(n226) );
  INVX1_HVT U258 ( .A(n1441), .Y(n1445) );
  INVX0_HVT U259 ( .A(n1917), .Y(n1921) );
  INVX1_HVT U260 ( .A(n1558), .Y(n219) );
  INVX0_HVT U261 ( .A(n1773), .Y(n482) );
  INVX0_HVT U262 ( .A(n1807), .Y(n479) );
  AOI22X1_HVT U263 ( .A1(n1933), .A2(n1932), .A3(n170), .A4(n1931), .Y(n1934)
         );
  INVX0_HVT U264 ( .A(n1728), .Y(n1729) );
  INVX0_HVT U265 ( .A(n1406), .Y(n1411) );
  INVX0_HVT U266 ( .A(n1531), .Y(n1530) );
  INVX0_HVT U267 ( .A(n1515), .Y(n1514) );
  INVX0_HVT U268 ( .A(n1075), .Y(n1059) );
  INVX0_HVT U269 ( .A(n888), .Y(n877) );
  INVX0_HVT U270 ( .A(n993), .Y(n493) );
  INVX0_HVT U271 ( .A(n1673), .Y(n1674) );
  INVX0_HVT U272 ( .A(n1621), .Y(n1622) );
  INVX0_HVT U273 ( .A(n1724), .Y(n1725) );
  INVX0_HVT U274 ( .A(n700), .Y(n698) );
  INVX0_HVT U275 ( .A(n861), .Y(n862) );
  INVX0_HVT U276 ( .A(n1890), .Y(n471) );
  INVX0_HVT U277 ( .A(n1166), .Y(n1167) );
  INVX0_HVT U278 ( .A(n1668), .Y(n1669) );
  INVX0_HVT U279 ( .A(n1457), .Y(net22654) );
  INVX0_HVT U280 ( .A(n1458), .Y(n1444) );
  INVX1_HVT U281 ( .A(n226), .Y(n203) );
  INVX1_HVT U282 ( .A(n219), .Y(n201) );
  INVX1_HVT U283 ( .A(n219), .Y(n202) );
  INVX0_HVT U284 ( .A(n964), .Y(n965) );
  INVX0_HVT U285 ( .A(n1988), .Y(n1945) );
  INVX0_HVT U286 ( .A(n1623), .Y(n1624) );
  INVX0_HVT U287 ( .A(n1617), .Y(n1618) );
  INVX0_HVT U288 ( .A(n1615), .Y(n1578) );
  INVX0_HVT U289 ( .A(n880), .Y(n881) );
  INVX0_HVT U290 ( .A(n1722), .Y(n1693) );
  INVX1_HVT U291 ( .A(n228), .Y(n197) );
  INVX1_HVT U292 ( .A(n209), .Y(n193) );
  INVX1_HVT U293 ( .A(n209), .Y(n187) );
  INVX1_HVT U294 ( .A(n228), .Y(n184) );
  INVX1_HVT U295 ( .A(n209), .Y(n199) );
  INVX1_HVT U296 ( .A(n227), .Y(n195) );
  INVX1_HVT U297 ( .A(n209), .Y(n186) );
  INVX1_HVT U298 ( .A(n228), .Y(n183) );
  INVX1_HVT U299 ( .A(n228), .Y(n198) );
  INVX1_HVT U300 ( .A(n228), .Y(n194) );
  INVX1_HVT U301 ( .A(n209), .Y(n200) );
  INVX1_HVT U302 ( .A(n227), .Y(n196) );
  INVX1_HVT U303 ( .A(n228), .Y(n182) );
  INVX0_HVT U304 ( .A(n667), .Y(n659) );
  INVX0_HVT U305 ( .A(n925), .Y(n926) );
  INVX0_HVT U306 ( .A(n1066), .Y(n1067) );
  INVX1_HVT U307 ( .A(n1261), .Y(n191) );
  INVX0_HVT U308 ( .A(n1715), .Y(n1716) );
  INVX0_HVT U309 ( .A(n589), .Y(n581) );
  INVX1_HVT U310 ( .A(n1261), .Y(n190) );
  INVX1_HVT U311 ( .A(n1261), .Y(n192) );
  INVX1_HVT U312 ( .A(n220), .Y(n188) );
  INVX0_HVT U313 ( .A(n695), .Y(n685) );
  AND2X1_HVT U314 ( .A1(n1368), .A2(n1305), .Y(n1268) );
  INVX0_HVT U315 ( .A(n1675), .Y(n1676) );
  INVX0_HVT U316 ( .A(n1370), .Y(n536) );
  INVX0_HVT U317 ( .A(n949), .Y(n946) );
  INVX0_HVT U318 ( .A(n749), .Y(n738) );
  INVX2_HVT U319 ( .A(n228), .Y(n174) );
  INVX2_HVT U320 ( .A(n228), .Y(n175) );
  INVX2_HVT U321 ( .A(n209), .Y(n176) );
  INVX2_HVT U322 ( .A(n209), .Y(n177) );
  INVX0_HVT U323 ( .A(n689), .Y(n707) );
  INVX0_HVT U324 ( .A(n1850), .Y(n1869) );
  INVX0_HVT U325 ( .A(n1768), .Y(n1769) );
  INVX0_HVT U326 ( .A(n1334), .Y(n978) );
  INVX0_HVT U327 ( .A(n1238), .Y(n895) );
  INVX1_HVT U328 ( .A(n226), .Y(n205) );
  INVX1_HVT U329 ( .A(n1975), .Y(n189) );
  INVX0_HVT U330 ( .A(n1942), .Y(n1982) );
  INVX0_HVT U331 ( .A(n1730), .Y(n1731) );
  INVX1_HVT U332 ( .A(n226), .Y(n204) );
  INVX0_HVT U333 ( .A(n1602), .Y(n1608) );
  INVX1_HVT U334 ( .A(n1317), .Y(n230) );
  INVX0_HVT U335 ( .A(n1336), .Y(n1342) );
  INVX0_HVT U336 ( .A(n1914), .Y(n1916) );
  INVX1_HVT U337 ( .A(n1317), .Y(n231) );
  INVX0_HVT U338 ( .A(n1802), .Y(n1803) );
  INVX0_HVT U339 ( .A(n2000), .Y(n2003) );
  INVX0_HVT U340 ( .A(n1996), .Y(n1999) );
  INVX0_HVT U341 ( .A(n1997), .Y(n526) );
  INVX0_HVT U342 ( .A(n1035), .Y(n1018) );
  INVX0_HVT U343 ( .A(n846), .Y(n848) );
  INVX0_HVT U344 ( .A(n1382), .Y(n1385) );
  NOR2X0_HVT U345 ( .A1(conv1_weight_done), .A2(n1667), .Y(n1975) );
  NOR2X1_HVT U346 ( .A1(n1925), .A2(sram_raddr_a4[8]), .Y(n1930) );
  AND2X1_HVT U347 ( .A1(n1568), .A2(n250), .Y(n1833) );
  INVX0_HVT U348 ( .A(n1765), .Y(n1767) );
  INVX0_HVT U349 ( .A(n1569), .Y(n1680) );
  INVX0_HVT U350 ( .A(n1139), .Y(n1128) );
  INVX0_HVT U351 ( .A(n1376), .Y(n1377) );
  INVX0_HVT U352 ( .A(n1091), .Y(n1092) );
  INVX0_HVT U353 ( .A(n668), .Y(n657) );
  INVX0_HVT U354 ( .A(n660), .Y(n661) );
  INVX0_HVT U355 ( .A(n558), .Y(n551) );
  INVX0_HVT U356 ( .A(n1328), .Y(n1330) );
  NOR2X1_HVT U357 ( .A1(n353), .A2(n1650), .Y(n1661) );
  INVX0_HVT U358 ( .A(n1547), .Y(n1546) );
  INVX0_HVT U359 ( .A(n1080), .Y(n1134) );
  INVX0_HVT U360 ( .A(n582), .Y(n583) );
  INVX0_HVT U361 ( .A(n590), .Y(n579) );
  INVX0_HVT U362 ( .A(n739), .Y(n740) );
  AOI22X1_HVT U363 ( .A1(sram_raddr_b7[6]), .A2(n1308), .A3(n1218), .A4(n1228), 
        .Y(n1219) );
  INVX0_HVT U364 ( .A(n920), .Y(n915) );
  INVX0_HVT U365 ( .A(n1565), .Y(n1388) );
  INVX0_HVT U366 ( .A(n1508), .Y(n1471) );
  INVX0_HVT U367 ( .A(n1026), .Y(n1028) );
  AND4X1_HVT U368 ( .A1(n554), .A2(row[0]), .A3(n553), .A4(n552), .Y(n1322) );
  INVX0_HVT U369 ( .A(n1952), .Y(n1957) );
  INVX1_HVT U370 ( .A(n1368), .Y(n179) );
  AND4X1_HVT U371 ( .A1(n554), .A2(n553), .A3(n319), .A4(n253), .Y(n1065) );
  INVX0_HVT U372 ( .A(n1293), .Y(n1291) );
  INVX0_HVT U373 ( .A(n1579), .Y(n1583) );
  INVX0_HVT U374 ( .A(n1581), .Y(n1580) );
  INVX0_HVT U375 ( .A(n575), .Y(n721) );
  INVX0_HVT U376 ( .A(n796), .Y(n799) );
  INVX0_HVT U377 ( .A(n1904), .Y(n1905) );
  INVX0_HVT U378 ( .A(n548), .Y(n554) );
  INVX0_HVT U379 ( .A(n1205), .Y(n1203) );
  INVX0_HVT U380 ( .A(n1549), .Y(n1548) );
  INVX0_HVT U381 ( .A(n646), .Y(n641) );
  INVX0_HVT U382 ( .A(n1858), .Y(n1859) );
  INVX0_HVT U383 ( .A(n1783), .Y(n1784) );
  INVX0_HVT U384 ( .A(n1554), .Y(n1553) );
  INVX0_HVT U385 ( .A(n728), .Y(n722) );
  INVX0_HVT U386 ( .A(n1749), .Y(n1750) );
  INVX0_HVT U387 ( .A(n731), .Y(n724) );
  AND2X2_HVT U388 ( .A1(mode[1]), .A2(n523), .Y(n1356) );
  INVX0_HVT U389 ( .A(mode[1]), .Y(n524) );
  INVX0_HVT U390 ( .A(n1632), .Y(n1633) );
  INVX0_HVT U391 ( .A(n1300), .Y(n1288) );
  INVX0_HVT U392 ( .A(n1472), .Y(n1474) );
  INVX0_HVT U393 ( .A(n1563), .Y(n1021) );
  AND4X1_HVT U394 ( .A1(state[1]), .A2(state[0]), .A3(n1023), .A4(state[2]), 
        .Y(n1558) );
  INVX1_HVT U395 ( .A(n227), .Y(n229) );
  INVX2_HVT U396 ( .A(n228), .Y(n206) );
  INVX2_HVT U397 ( .A(n228), .Y(n208) );
  INVX2_HVT U398 ( .A(n228), .Y(n207) );
  INVX2_HVT U399 ( .A(n209), .Y(n210) );
  NAND2X2_HVT U400 ( .A1(n556), .A2(n1357), .Y(n1456) );
  INVX1_HVT U401 ( .A(n1308), .Y(n211) );
  INVX1_HVT U402 ( .A(n1308), .Y(n212) );
  INVX2_HVT U403 ( .A(n1308), .Y(n213) );
  INVX2_HVT U404 ( .A(n1308), .Y(n214) );
  INVX1_HVT U405 ( .A(n1268), .Y(n215) );
  INVX1_HVT U406 ( .A(n1833), .Y(n216) );
  INVX1_HVT U407 ( .A(n1065), .Y(n217) );
  INVX1_HVT U408 ( .A(n1065), .Y(n218) );
  INVX1_HVT U409 ( .A(n179), .Y(n220) );
  INVX1_HVT U410 ( .A(n220), .Y(n221) );
  INVX1_HVT U411 ( .A(n220), .Y(n222) );
  INVX1_HVT U412 ( .A(n220), .Y(n223) );
  INVX1_HVT U413 ( .A(n1322), .Y(n224) );
  INVX1_HVT U414 ( .A(n1322), .Y(n225) );
  OAI21X1_HVT U415 ( .A1(n559), .A2(n558), .A3(n1545), .Y(n1317) );
  INVX0_HVT U416 ( .A(n1317), .Y(n232) );
  INVX1_HVT U417 ( .A(n1391), .Y(n2004) );
  INVX1_HVT U418 ( .A(n231), .Y(n1305) );
  OR2X1_HVT U419 ( .A1(n556), .A2(n557), .Y(n1368) );
  INVX1_HVT U420 ( .A(n1200), .Y(n1228) );
  INVX1_HVT U421 ( .A(n1946), .Y(n1990) );
  NAND4X0_HVT U422 ( .A1(state[0]), .A2(state[1]), .A3(n1023), .A4(n1024), .Y(
        n1391) );
  INVX1_HVT U423 ( .A(n216), .Y(n1897) );
  INVX1_HVT U424 ( .A(n677), .Y(n706) );
  INVX1_HVT U425 ( .A(n1359), .Y(n1365) );
  OA221X1_HVT U426 ( .A1(n1569), .A2(n1052), .A3(n1569), .A4(
        addr_col_sel_cnt[1]), .A5(n1560), .Y(n1946) );
  INVX1_HVT U427 ( .A(n1456), .Y(n1466) );
  INVX1_HVT U428 ( .A(n217), .Y(n1262) );
  INVX1_HVT U429 ( .A(n1301), .Y(n1320) );
  OAI21X1_HVT U430 ( .A1(n250), .A2(n1357), .A3(n1371), .Y(n_conv1_weight_done) );
  INVX1_HVT U431 ( .A(n1501), .Y(n1507) );
  OAI21X1_HVT U432 ( .A1(n769), .A2(n275), .A3(n792), .Y(n1315) );
  OA221X1_HVT U433 ( .A1(n1569), .A2(n1052), .A3(n1569), .A4(n1051), .A5(n1560), .Y(n1760) );
  INVX1_HVT U434 ( .A(n556), .Y(n1550) );
  NAND3X0_HVT U435 ( .A1(n1024), .A2(n1446), .A3(state[3]), .Y(n556) );
  INVX1_HVT U436 ( .A(n544), .Y(n546) );
  INVX1_HVT U437 ( .A(n545), .Y(n547) );
  INVX1_HVT U438 ( .A(mem_sel), .Y(n1513) );
  INVX1_HVT U439 ( .A(n1799), .Y(n1801) );
  INVX1_HVT U440 ( .A(n1245), .Y(n1260) );
  INVX1_HVT U441 ( .A(n1333), .Y(n1348) );
  OAI21X1_HVT U442 ( .A1(n1276), .A2(n381), .A3(n750), .Y(n1289) );
  AO221X1_HVT U443 ( .A1(sram_raddr_b1[9]), .A2(n965), .A3(n377), .A4(n964), 
        .A5(n218), .Y(n1245) );
  OAI21X1_HVT U444 ( .A1(sram_raddr_a4[5]), .A2(n1643), .A3(n1650), .Y(n1787)
         );
  OAI21X1_HVT U445 ( .A1(n680), .A2(n347), .A3(n689), .Y(n1231) );
  OAI21X1_HVT U446 ( .A1(sram_raddr_a5[4]), .A2(n1694), .A3(n1700), .Y(n1817)
         );
  AO221X1_HVT U447 ( .A1(sram_raddr_b2[9]), .A2(n1067), .A3(n419), .A4(n1066), 
        .A5(n217), .Y(n1333) );
  OAI21X1_HVT U448 ( .A1(sram_raddr_b4[6]), .A2(n670), .A3(n679), .Y(n930) );
  OAI21X1_HVT U449 ( .A1(sram_raddr_a5[6]), .A2(n1707), .A3(n1714), .Y(n1826)
         );
  OAI21X1_HVT U450 ( .A1(n603), .A2(n338), .A3(n623), .Y(n1145) );
  AO22X1_HVT U451 ( .A1(write_row_conv1[0]), .A2(n1365), .A3(n1356), .A4(
        col_enable[1]), .Y(n544) );
  AO22X1_HVT U452 ( .A1(write_col_conv1[0]), .A2(n1365), .A3(n1356), .A4(
        col_enable[0]), .Y(n545) );
  AND2X1_HVT U453 ( .A1(n1529), .A2(n1513), .Y(n1528) );
  AND2X1_HVT U454 ( .A1(n1529), .A2(mem_sel), .Y(n1544) );
  INVX1_HVT U455 ( .A(n1499), .Y(n1506) );
  AO21X1_HVT U456 ( .A1(n1477), .A2(n1476), .A3(n1508), .Y(n1501) );
  AND4X1_HVT U457 ( .A1(n1570), .A2(n1053), .A3(n2004), .A4(n317), .Y(n1568)
         );
  INVX2_HVT U458 ( .A(n1760), .Y(n1888) );
  AND2X1_HVT U459 ( .A1(n1365), .A2(delay2_write_enable), .Y(n1470) );
  NAND2X0_HVT U460 ( .A1(mode[0]), .A2(n524), .Y(n1359) );
  INVX2_HVT U461 ( .A(n1893), .Y(n1935) );
  INVX1_HVT U462 ( .A(n522), .Y(n1570) );
  NAND2X0_HVT U463 ( .A1(n1994), .A2(n250), .Y(n1569) );
  AND2X1_HVT U464 ( .A1(n2004), .A2(n522), .Y(n1994) );
  NAND3X0_HVT U465 ( .A1(n553), .A2(n252), .A3(n321), .Y(n558) );
  AND3X1_HVT U466 ( .A1(n1566), .A2(n238), .A3(n233), .Y(n553) );
  NAND2X0_HVT U467 ( .A1(row[1]), .A2(row[0]), .Y(n559) );
  INVX1_HVT U468 ( .A(n1363), .Y(n1545) );
  NAND2X0_HVT U469 ( .A1(channel_cnt[1]), .A2(channel_cnt[0]), .Y(n1549) );
  NAND4X0_HVT U470 ( .A1(n1053), .A2(n1570), .A3(n2004), .A4(
        addr_row_sel_cnt[0]), .Y(n1667) );
  INVX1_HVT U471 ( .A(n1564), .Y(n1020) );
  NOR4X1_HVT U472 ( .A1(conv2_weight_cnt[7]), .A2(conv2_weight_cnt[6]), .A3(
        n530), .A4(n529), .Y(n_conv_done) );
  NOR4X1_HVT U473 ( .A1(conv1_weight_cnt[7]), .A2(conv1_weight_cnt[6]), .A3(
        conv1_weight_cnt[5]), .A4(n1359), .Y(n527) );
  NOR4X1_HVT U474 ( .A1(conv1_done), .A2(conv1_weight_cnt[1]), .A3(
        conv1_weight_cnt[0]), .A4(conv1_weight_cnt[3]), .Y(n528) );
  NOR4X1_HVT U475 ( .A1(channel_cnt[1]), .A2(channel_cnt[4]), .A3(
        conv2_weight_done), .A4(n531), .Y(n532) );
  INVX1_HVT U476 ( .A(n2001), .Y(n1995) );
  INVX1_HVT U477 ( .A(n1517), .Y(n1516) );
  INVX1_HVT U478 ( .A(n1519), .Y(n1518) );
  INVX1_HVT U479 ( .A(n1521), .Y(n1520) );
  INVX1_HVT U480 ( .A(n1523), .Y(n1522) );
  INVX1_HVT U481 ( .A(n1525), .Y(n1524) );
  INVX1_HVT U482 ( .A(n1533), .Y(n1532) );
  INVX1_HVT U483 ( .A(n1535), .Y(n1534) );
  INVX1_HVT U484 ( .A(n1537), .Y(n1536) );
  INVX1_HVT U485 ( .A(n1539), .Y(n1538) );
  INVX1_HVT U486 ( .A(n1541), .Y(n1540) );
  NOR4X1_HVT U487 ( .A1(delay1_sram_waddr_b[0]), .A2(delay1_sram_waddr_b[1]), 
        .A3(delay1_sram_waddr_b[2]), .A4(delay1_sram_waddr_b[3]), .Y(n1495) );
  INVX1_HVT U488 ( .A(n1390), .Y(n1567) );
  INVX1_HVT U489 ( .A(n1373), .Y(n1379) );
  INVX1_HVT U490 ( .A(n1804), .Y(n1795) );
  INVX1_HVT U491 ( .A(n1870), .Y(n1875) );
  INVX1_HVT U492 ( .A(n1629), .Y(n1630) );
  INVX1_HVT U493 ( .A(n973), .Y(n960) );
  INVX1_HVT U494 ( .A(n1844), .Y(n1831) );
  INVX1_HVT U495 ( .A(n1392), .Y(n1442) );
  INVX1_HVT U496 ( .A(n1839), .Y(n1943) );
  INVX1_HVT U497 ( .A(n1986), .Y(n1987) );
  INVX1_HVT U498 ( .A(n1974), .Y(n1976) );
  INVX1_HVT U499 ( .A(n1963), .Y(n1968) );
  INVX1_HVT U500 ( .A(n1842), .Y(n1843) );
  INVX1_HVT U501 ( .A(n1827), .Y(n1832) );
  INVX1_HVT U502 ( .A(n1818), .Y(n1822) );
  INVX1_HVT U503 ( .A(n1761), .Y(n1762) );
  INVX1_HVT U504 ( .A(n1770), .Y(n1759) );
  INVX1_HVT U505 ( .A(n1151), .Y(n1152) );
  INVX1_HVT U506 ( .A(n1147), .Y(n1149) );
  INVX1_HVT U507 ( .A(n1136), .Y(n1137) );
  INVX1_HVT U508 ( .A(n1232), .Y(n1234) );
  INVX1_HVT U509 ( .A(n1235), .Y(n1236) );
  INVX1_HVT U510 ( .A(n1248), .Y(n1254) );
  NAND2X0_HVT U511 ( .A1(n1261), .A2(n1080), .Y(n1164) );
  NAND2X0_HVT U512 ( .A1(n1261), .A2(n1176), .Y(n1250) );
  NAND2X0_HVT U513 ( .A1(n1261), .A2(n1328), .Y(n1338) );
  INVX1_HVT U514 ( .A(n951), .Y(n952) );
  INVX1_HVT U515 ( .A(n683), .Y(n696) );
  INVX1_HVT U516 ( .A(n692), .Y(n711) );
  INVX1_HVT U517 ( .A(n944), .Y(n950) );
  INVX1_HVT U518 ( .A(n928), .Y(n1204) );
  INVX1_HVT U519 ( .A(n901), .Y(n914) );
  INVX1_HVT U520 ( .A(n957), .Y(n970) );
  NAND2X0_HVT U521 ( .A1(col[1]), .A2(n211), .Y(n1334) );
  INVX1_HVT U522 ( .A(n1321), .Y(n1323) );
  INVX1_HVT U523 ( .A(n1316), .Y(n1319) );
  INVX1_HVT U524 ( .A(n1042), .Y(n1057) );
  INVX1_HVT U525 ( .A(n1015), .Y(n1292) );
  INVX1_HVT U526 ( .A(n1019), .Y(n1073) );
  INVX1_HVT U527 ( .A(n1001), .Y(n999) );
  INVX1_HVT U528 ( .A(n843), .Y(n1110) );
  INVX1_HVT U529 ( .A(n863), .Y(n886) );
  INVX1_HVT U530 ( .A(n867), .Y(n868) );
  INVX1_HVT U531 ( .A(n829), .Y(n827) );
  INVX1_HVT U532 ( .A(n1086), .Y(n1160) );
  INVX1_HVT U533 ( .A(n763), .Y(n1000) );
  INVX1_HVT U534 ( .A(n750), .Y(n758) );
  NAND2X0_HVT U535 ( .A1(n721), .A2(n312), .Y(n1301) );
  INVX1_HVT U536 ( .A(n746), .Y(n747) );
  INVX1_HVT U537 ( .A(n787), .Y(n744) );
  NAND2X0_HVT U538 ( .A1(n217), .A2(n1328), .Y(n787) );
  INVX1_HVT U539 ( .A(n665), .Y(n666) );
  INVX1_HVT U540 ( .A(n1150), .Y(n1127) );
  INVX1_HVT U541 ( .A(n607), .Y(n605) );
  INVX1_HVT U542 ( .A(n597), .Y(n828) );
  INVX1_HVT U543 ( .A(n777), .Y(n690) );
  INVX1_HVT U544 ( .A(n1645), .Y(n1646) );
  INVX1_HVT U545 ( .A(n587), .Y(n588) );
  INVX1_HVT U546 ( .A(n608), .Y(n622) );
  NAND3X0_HVT U547 ( .A1(n238), .A2(n254), .A3(n233), .Y(n1200) );
  NAND2X0_HVT U548 ( .A1(n1176), .A2(n1328), .Y(n1150) );
  INVX1_HVT U549 ( .A(n1430), .Y(n1425) );
  INVX1_HVT U550 ( .A(n1434), .Y(n1429) );
  INVX1_HVT U551 ( .A(n1410), .Y(n1407) );
  INVX1_HVT U552 ( .A(n1412), .Y(n1418) );
  INVX1_HVT U553 ( .A(n1436), .Y(n1439) );
  INVX1_HVT U554 ( .A(n1709), .Y(n1710) );
  INVX1_HVT U555 ( .A(n1702), .Y(n1703) );
  INVX1_HVT U556 ( .A(n1695), .Y(n1696) );
  NAND2X0_HVT U557 ( .A1(n172), .A2(n1942), .Y(n1722) );
  INVX1_HVT U558 ( .A(n1607), .Y(n1606) );
  INVX1_HVT U559 ( .A(n1588), .Y(n1587) );
  INVX1_HVT U560 ( .A(n1593), .Y(n1594) );
  INVX1_HVT U561 ( .A(n1589), .Y(n1590) );
  NAND2X0_HVT U562 ( .A1(n172), .A2(n1850), .Y(n1615) );
  NAND2X0_HVT U563 ( .A1(n181), .A2(n1561), .Y(net31203) );
  NOR4X1_HVT U564 ( .A1(n1549), .A2(n311), .A3(channel_cnt[3]), .A4(
        channel_cnt[2]), .Y(n557) );
  OAI221X1_HVT U565 ( .A1(n1135), .A2(n1134), .A3(n1135), .A4(n1133), .A5(n204), .Y(n263) );
  OAI221X1_HVT U566 ( .A1(n1146), .A2(n1164), .A3(n1146), .A4(n1145), .A5(n201), .Y(n264) );
  OAI221X1_HVT U567 ( .A1(n1124), .A2(n1164), .A3(n1124), .A4(n1123), .A5(n202), .Y(n265) );
  OAI221X1_HVT U568 ( .A1(n733), .A2(n1322), .A3(n733), .A4(n992), .A5(n204), 
        .Y(n266) );
  AND3X1_HVT U569 ( .A1(n1417), .A2(n1467), .A3(n1563), .Y(n283) );
  AND4X1_HVT U570 ( .A1(n1358), .A2(n1447), .A3(n1363), .A4(n1367), .Y(n285)
         );
  OAI221X1_HVT U571 ( .A1(sram_raddr_b4[5]), .A2(n1204), .A3(n276), .A4(n928), 
        .A5(n223), .Y(n302) );
  AOI22X1_HVT U572 ( .A1(n178), .A2(n1085), .A3(n1084), .A4(n1164), .Y(n303)
         );
  AOI22X1_HVT U573 ( .A1(n1778), .A2(n1804), .A3(sram_raddr_a4[2]), .A4(n1935), 
        .Y(n304) );
  AOI22X1_HVT U574 ( .A1(sram_raddr_b7[1]), .A2(n1238), .A3(n1180), .A4(n1250), 
        .Y(n305) );
  AOI22X1_HVT U575 ( .A1(n1975), .A2(n235), .A3(n1898), .A4(n1932), .Y(n306)
         );
  AOI22X1_HVT U576 ( .A1(sram_raddr_a6[2]), .A2(n1888), .A3(n1852), .A4(n1886), 
        .Y(n307) );
  AOI22X1_HVT U577 ( .A1(sram_raddr_a6[1]), .A2(n1888), .A3(n1869), .A4(n1851), 
        .Y(n308) );
  AOI22X1_HVT U578 ( .A1(sram_raddr_b8[1]), .A2(n1334), .A3(n1266), .A4(n1338), 
        .Y(n309) );
  AOI22X1_HVT U579 ( .A1(n1739), .A2(n1770), .A3(sram_raddr_a3[2]), .A4(n1888), 
        .Y(n328) );
  AOI22X1_HVT U580 ( .A1(sram_raddr_a2[9]), .A2(n1734), .A3(n1733), .A4(n1732), 
        .Y(n329) );
  AOI22X1_HVT U581 ( .A1(sram_raddr_a1[9]), .A2(n1679), .A3(n1678), .A4(n1677), 
        .Y(n330) );
  AOI22X1_HVT U582 ( .A1(sram_raddr_a0[9]), .A2(n1627), .A3(n1626), .A4(n1625), 
        .Y(n331) );
  AND3X1_HVT U583 ( .A1(n1282), .A2(n991), .A3(n990), .Y(n390) );
  AND2X1_HVT U584 ( .A1(n1357), .A2(n1564), .Y(n400) );
  OAI222X1_HVT U585 ( .A1(sram_raddr_weight[5]), .A2(n1439), .A3(
        sram_raddr_weight[5]), .A4(n1456), .A5(n422), .A6(n1438), .Y(n450) );
  OAI221X1_HVT U586 ( .A1(sram_raddr_a1[2]), .A2(n1638), .A3(sram_raddr_a1[2]), 
        .A4(n1665), .A5(n1631), .Y(n456) );
  OAI221X1_HVT U587 ( .A1(n927), .A2(n957), .A3(n927), .A4(n926), .A5(n202), 
        .Y(n457) );
  AOI22X1_HVT U588 ( .A1(sram_raddr_a6[9]), .A2(n1888), .A3(n1887), .A4(n1886), 
        .Y(n458) );
  NAND2X0_HVT U589 ( .A1(n168), .A2(n1898), .Y(n459) );
  NAND2X0_HVT U590 ( .A1(n1897), .A2(n248), .Y(n461) );
  NAND2X0_HVT U591 ( .A1(n172), .A2(n1914), .Y(n1665) );
  NAND2X0_HVT U592 ( .A1(n517), .A2(n518), .Y(n462) );
  NAND2X0_HVT U593 ( .A1(n503), .A2(n504), .Y(n463) );
  NAND2X0_HVT U594 ( .A1(n499), .A2(n500), .Y(n464) );
  NAND2X0_HVT U595 ( .A1(n501), .A2(n502), .Y(n466) );
  NAND2X0_HVT U596 ( .A1(n497), .A2(n498), .Y(n467) );
  NAND2X0_HVT U597 ( .A1(sram_raddr_a7[9]), .A2(n1935), .Y(n469) );
  NAND3X0_HVT U598 ( .A1(n1934), .A2(n468), .A3(n469), .Y(n_sram_raddr_a7[9])
         );
  NAND2X0_HVT U599 ( .A1(sram_raddr_a7[2]), .A2(n1935), .Y(n470) );
  NAND3X0_HVT U600 ( .A1(n306), .A2(n475), .A3(n470), .Y(n_sram_raddr_a7[2])
         );
  NAND2X0_HVT U601 ( .A1(n1975), .A2(n1889), .Y(n472) );
  NAND3X0_HVT U602 ( .A1(n458), .A2(n471), .A3(n472), .Y(n_sram_raddr_a6[9])
         );
  NAND2X0_HVT U603 ( .A1(n1975), .A2(n234), .Y(n473) );
  NAND3X0_HVT U604 ( .A1(n307), .A2(n461), .A3(n473), .Y(n_sram_raddr_a6[2])
         );
  NAND2X0_HVT U605 ( .A1(n170), .A2(sram_raddr_a3[1]), .Y(n474) );
  NAND3X0_HVT U606 ( .A1(n308), .A2(n1849), .A3(n474), .Y(n_sram_raddr_a6[1])
         );
  NAND2X0_HVT U607 ( .A1(n1897), .A2(n247), .Y(n475) );
  NAND3X0_HVT U608 ( .A1(n304), .A2(n459), .A3(n475), .Y(n_sram_raddr_a4[2])
         );
  NAND2X0_HVT U609 ( .A1(n1852), .A2(n168), .Y(n476) );
  NAND3X0_HVT U610 ( .A1(n328), .A2(n461), .A3(n476), .Y(n_sram_raddr_a3[2])
         );
  NAND2X0_HVT U611 ( .A1(n170), .A2(n1845), .Y(n478) );
  NAND3X0_HVT U612 ( .A1(n329), .A2(n477), .A3(n478), .Y(n_sram_raddr_a2[9])
         );
  NAND2X0_HVT U613 ( .A1(n170), .A2(n1805), .Y(n480) );
  NAND3X0_HVT U614 ( .A1(n330), .A2(n479), .A3(n480), .Y(n_sram_raddr_a1[9])
         );
  NAND2X0_HVT U615 ( .A1(n1975), .A2(n1778), .Y(n481) );
  NAND3X0_HVT U616 ( .A1(n459), .A2(n456), .A3(n481), .Y(n_sram_raddr_a1[2])
         );
  NAND2X0_HVT U617 ( .A1(n170), .A2(n1771), .Y(n483) );
  NAND3X0_HVT U618 ( .A1(n331), .A2(n482), .A3(n483), .Y(n_sram_raddr_a0[9])
         );
  NAND2X0_HVT U619 ( .A1(n203), .A2(n1440), .Y(n484) );
  NAND3X0_HVT U620 ( .A1(n450), .A2(n283), .A3(n484), .Y(net22796) );
  NAND2X0_HVT U621 ( .A1(n1559), .A2(n449), .Y(n485) );
  NAND3X0_HVT U622 ( .A1(n285), .A2(n400), .A3(n485), .Y(n_state[0]) );
  NAND2X0_HVT U623 ( .A1(n178), .A2(n1267), .Y(n486) );
  NAND3X0_HVT U624 ( .A1(n309), .A2(n1265), .A3(n486), .Y(n1269) );
  NAND2X0_HVT U625 ( .A1(n1220), .A2(n1250), .Y(n487) );
  NAND3X0_HVT U626 ( .A1(n1219), .A2(n467), .A3(n487), .Y(n1225) );
  NAND2X0_HVT U627 ( .A1(n178), .A2(n1181), .Y(n488) );
  NAND3X0_HVT U628 ( .A1(n305), .A2(n1179), .A3(n488), .Y(n1182) );
  NAND2X0_HVT U629 ( .A1(sram_raddr_b6[7]), .A2(n230), .Y(n489) );
  NAND3X0_HVT U630 ( .A1(n464), .A2(n264), .A3(n489), .Y(n_sram_raddr_b6[7])
         );
  NAND2X0_HVT U631 ( .A1(sram_raddr_b6[6]), .A2(n231), .Y(n490) );
  NAND3X0_HVT U632 ( .A1(n466), .A2(n263), .A3(n490), .Y(n_sram_raddr_b6[6])
         );
  NAND2X0_HVT U633 ( .A1(sram_raddr_b6[5]), .A2(n231), .Y(n491) );
  NAND3X0_HVT U634 ( .A1(n463), .A2(n265), .A3(n491), .Y(n_sram_raddr_b6[5])
         );
  NAND2X0_HVT U635 ( .A1(sram_raddr_b6[1]), .A2(n1086), .Y(n492) );
  NAND3X0_HVT U636 ( .A1(n303), .A2(n1083), .A3(n492), .Y(n1087) );
  NAND2X0_HVT U637 ( .A1(n992), .A2(n1019), .Y(n494) );
  NAND3X0_HVT U638 ( .A1(n390), .A2(n493), .A3(n494), .Y(n997) );
  NAND2X0_HVT U639 ( .A1(sram_raddr_b4[5]), .A2(n232), .Y(n495) );
  NAND3X0_HVT U640 ( .A1(n302), .A2(n457), .A3(n495), .Y(n_sram_raddr_b4[5])
         );
  NAND2X0_HVT U641 ( .A1(sram_raddr_b2[3]), .A2(n231), .Y(n496) );
  NAND3X0_HVT U642 ( .A1(n462), .A2(n266), .A3(n496), .Y(n_sram_raddr_b2[3])
         );
  AND2X1_HVT U643 ( .A1(n519), .A2(n520), .Y(n1839) );
  AND2X1_HVT U644 ( .A1(n1229), .A2(n178), .Y(n497) );
  OR2X1_HVT U645 ( .A1(n1216), .A2(sram_raddr_b4[6]), .Y(n498) );
  AND2X1_HVT U646 ( .A1(n1148), .A2(n223), .Y(n499) );
  OR2X1_HVT U647 ( .A1(n1149), .A2(sram_raddr_b6[7]), .Y(n500) );
  AND2X1_HVT U648 ( .A1(n1147), .A2(n221), .Y(n501) );
  OR2X1_HVT U649 ( .A1(n1137), .A2(sram_raddr_b6[6]), .Y(n502) );
  AND2X1_HVT U650 ( .A1(n1136), .A2(n223), .Y(n503) );
  OR2X1_HVT U651 ( .A1(n1125), .A2(sram_raddr_b6[5]), .Y(n504) );
  AND2X1_HVT U652 ( .A1(n1071), .A2(n1074), .Y(n505) );
  OR2X1_HVT U653 ( .A1(n1072), .A2(n1073), .Y(n506) );
  AND2X1_HVT U654 ( .A1(n505), .A2(n506), .Y(n1076) );
  AND2X1_HVT U655 ( .A1(n1011), .A2(n1013), .Y(n507) );
  OR2X1_HVT U656 ( .A1(n1012), .A2(n1073), .Y(n508) );
  AND2X1_HVT U657 ( .A1(n507), .A2(n508), .Y(n1014) );
  AND2X1_HVT U658 ( .A1(n1010), .A2(n1304), .Y(n509) );
  OR2X1_HVT U659 ( .A1(n1301), .A2(n1026), .Y(n510) );
  AND2X1_HVT U660 ( .A1(n509), .A2(n510), .Y(n1013) );
  AND2X1_HVT U661 ( .A1(n968), .A2(n971), .Y(n511) );
  OR2X1_HVT U662 ( .A1(n969), .A2(n970), .Y(n512) );
  AND2X1_HVT U663 ( .A1(n511), .A2(n512), .Y(n972) );
  AND2X1_HVT U664 ( .A1(n884), .A2(n887), .Y(n513) );
  OR2X1_HVT U665 ( .A1(n885), .A2(n886), .Y(n514) );
  AND2X1_HVT U666 ( .A1(n513), .A2(n514), .Y(n889) );
  AND2X1_HVT U667 ( .A1(n743), .A2(n745), .Y(n515) );
  OR2X1_HVT U668 ( .A1(n255), .A2(n744), .Y(n516) );
  AND2X1_HVT U669 ( .A1(n515), .A2(n516), .Y(n748) );
  AND2X1_HVT U670 ( .A1(n998), .A2(n188), .Y(n517) );
  OR2X1_HVT U671 ( .A1(sram_raddr_b2[2]), .A2(sram_raddr_b2[3]), .Y(n518) );
  AND2X1_HVT U672 ( .A1(n317), .A2(n1572), .Y(n519) );
  OR2X1_HVT U673 ( .A1(n1571), .A2(n253), .Y(n520) );
  AND2X1_HVT U674 ( .A1(n519), .A2(n520), .Y(n521) );
  AO21X1_HVT U675 ( .A1(n523), .A2(n524), .A3(n1070), .Y(N2914) );
  AND2X1_HVT U676 ( .A1(col[1]), .A2(col[0]), .Y(n1566) );
  NAND3X0_HVT U677 ( .A1(n1566), .A2(col[3]), .A3(n233), .Y(n522) );
  AND3X1_HVT U678 ( .A1(n1994), .A2(n1051), .A3(n1052), .Y(
        n_addr_col_sel_cnt[0]) );
  AND3X1_HVT U679 ( .A1(n1051), .A2(n1994), .A3(addr_col_sel_cnt[0]), .Y(
        n_addr_col_sel_cnt[1]) );
  AO21X1_HVT U680 ( .A1(addr_row_sel_cnt[0]), .A2(n1994), .A3(n1568), .Y(
        n_addr_row_sel_cnt_0_) );
  AO22X1_HVT U681 ( .A1(col[1]), .A2(n1356), .A3(n1365), .A4(data_sel_col[1]), 
        .Y(n1997) );
  AO22X1_HVT U682 ( .A1(row[1]), .A2(n1356), .A3(n1365), .A4(data_sel_row[1]), 
        .Y(n2001) );
  AO22X1_HVT U683 ( .A1(row[0]), .A2(n1356), .A3(n1365), .A4(data_sel_row[0]), 
        .Y(n2000) );
  NAND2X0_HVT U684 ( .A1(n2004), .A2(n2000), .Y(n525) );
  OA22X1_HVT U685 ( .A1(n526), .A2(n1391), .A3(n1995), .A4(n525), .Y(n1662) );
  AO22X1_HVT U686 ( .A1(col[0]), .A2(n1356), .A3(n1365), .A4(data_sel_col[0]), 
        .Y(n1996) );
  AND2X1_HVT U687 ( .A1(n310), .A2(n251), .Y(n1446) );
  NAND3X0_HVT U688 ( .A1(n226), .A2(n556), .A3(n1391), .Y(n1998) );
  NAND2X0_HVT U689 ( .A1(n219), .A2(n556), .Y(n2002) );
  NAND3X0_HVT U690 ( .A1(n2004), .A2(n1997), .A3(n1996), .Y(n1655) );
  AND4X1_HVT U691 ( .A1(conv1_weight_cnt[2]), .A2(conv1_weight_cnt[4]), .A3(
        n528), .A4(n527), .Y(n_conv1_done) );
  NAND4X0_HVT U692 ( .A1(state[1]), .A2(n1023), .A3(n1024), .A4(n310), .Y(
        n1357) );
  AO22X1_HVT U693 ( .A1(row[1]), .A2(col[3]), .A3(row[0]), .A4(col[2]), .Y(
        n533) );
  OA21X1_HVT U694 ( .A1(row[0]), .A2(col[2]), .A3(n1566), .Y(n534) );
  NAND2X0_HVT U695 ( .A1(n319), .A2(n238), .Y(n550) );
  NAND2X0_HVT U696 ( .A1(row[1]), .A2(col[3]), .Y(n549) );
  NAND2X0_HVT U697 ( .A1(n550), .A2(n549), .Y(n552) );
  NAND3X0_HVT U698 ( .A1(row[1]), .A2(row[3]), .A3(n252), .Y(n1571) );
  NAND2X0_HVT U699 ( .A1(n252), .A2(n559), .Y(n539) );
  OR2X1_HVT U700 ( .A1(n1391), .A2(n535), .Y(n1371) );
  OR4X1_HVT U701 ( .A1(conv_done), .A2(conv2_weight_cnt[3]), .A3(
        conv2_weight_cnt[0]), .A4(conv2_weight_cnt[2]), .Y(n530) );
  NAND4X0_HVT U702 ( .A1(n1356), .A2(conv2_weight_cnt[5]), .A3(
        conv2_weight_cnt[1]), .A4(conv2_weight_cnt[4]), .Y(n529) );
  AND2X1_HVT U703 ( .A1(n2004), .A2(n250), .Y(n1559) );
  NAND2X0_HVT U704 ( .A1(n1228), .A2(n312), .Y(n1080) );
  NOR2X0_HVT U705 ( .A1(n556), .A2(channel_cnt[0]), .Y(net22937) );
  OR2X1_HVT U706 ( .A1(channel_cnt[2]), .A2(channel_cnt[3]), .Y(n531) );
  AO22X1_HVT U707 ( .A1(n1559), .A2(n1134), .A3(net22937), .A4(n532), .Y(
        n_load_data_enable) );
  NAND2X0_HVT U708 ( .A1(n252), .A2(n321), .Y(n548) );
  AO221X1_HVT U709 ( .A1(n550), .A2(n534), .A3(n550), .A4(n533), .A5(n548), 
        .Y(n1392) );
  NAND2X0_HVT U710 ( .A1(n205), .A2(n1442), .Y(n1458) );
  NAND2X0_HVT U711 ( .A1(n2004), .A2(n535), .Y(n1370) );
  OA22X1_HVT U712 ( .A1(n553), .A2(n1458), .A3(n1570), .A4(n1370), .Y(n1390)
         );
  NAND2X0_HVT U713 ( .A1(n1466), .A2(n1390), .Y(n538) );
  AO22X1_HVT U714 ( .A1(n1570), .A2(n536), .A3(n553), .A4(n1444), .Y(n540) );
  AO22X1_HVT U715 ( .A1(row[0]), .A2(n538), .A3(n253), .A4(n540), .Y(n_row[0])
         );
  AO21X1_HVT U716 ( .A1(row[0]), .A2(n540), .A3(row[1]), .Y(n537) );
  OA221X1_HVT U717 ( .A1(n538), .A2(n559), .A3(n538), .A4(n540), .A5(n537), 
        .Y(n_row[1]) );
  AO221X1_HVT U719 ( .A1(n540), .A2(n252), .A3(n540), .A4(n559), .A5(n538), 
        .Y(n541) );
  AND3X1_HVT U720 ( .A1(row[0]), .A2(row[1]), .A3(n540), .Y(n542) );
  AO22X1_HVT U721 ( .A1(row[2]), .A2(n542), .A3(row[3]), .A4(n541), .Y(
        n_row[3]) );
  AND2X1_HVT U722 ( .A1(n545), .A2(n544), .Y(n543) );
  AND2X1_HVT U723 ( .A1(n1470), .A2(n543), .Y(n_sram_bytemask_b[0]) );
  AND3X1_HVT U724 ( .A1(n547), .A2(n1470), .A3(n544), .Y(n_sram_bytemask_b[1])
         );
  AND3X1_HVT U725 ( .A1(n1470), .A2(n546), .A3(n545), .Y(n_sram_bytemask_b[2])
         );
  AND3X1_HVT U726 ( .A1(n1470), .A2(n547), .A3(n546), .Y(n_sram_bytemask_b[3])
         );
  AND3X1_HVT U727 ( .A1(n1356), .A2(n543), .A3(n1513), .Y(n_sram_bytemask_c[0]) );
  AND4X1_HVT U728 ( .A1(n1356), .A2(n547), .A3(n1513), .A4(n544), .Y(
        n_sram_bytemask_c[1]) );
  AND4X1_HVT U729 ( .A1(n1356), .A2(n546), .A3(n1513), .A4(n545), .Y(
        n_sram_bytemask_c[2]) );
  AND4X1_HVT U730 ( .A1(n1356), .A2(n547), .A3(n546), .A4(n1513), .Y(
        n_sram_bytemask_c[3]) );
  AND3X1_HVT U731 ( .A1(mem_sel), .A2(n1356), .A3(n543), .Y(
        n_sram_bytemask_d[0]) );
  AND4X1_HVT U732 ( .A1(n1356), .A2(mem_sel), .A3(n547), .A4(n544), .Y(
        n_sram_bytemask_d[1]) );
  AND4X1_HVT U733 ( .A1(n1356), .A2(mem_sel), .A3(n546), .A4(n545), .Y(
        n_sram_bytemask_d[2]) );
  AND4X1_HVT U734 ( .A1(mem_sel), .A2(n1356), .A3(n547), .A4(n546), .Y(
        n_sram_bytemask_d[3]) );
  NAND2X0_HVT U735 ( .A1(n238), .A2(n233), .Y(n575) );
  AO21X1_HVT U736 ( .A1(n1566), .A2(n548), .A3(n575), .Y(n1308) );
  AO22X1_HVT U737 ( .A1(col[1]), .A2(col[0]), .A3(n312), .A4(n254), .Y(n1389)
         );
  NAND2X0_HVT U738 ( .A1(n212), .A2(n1389), .Y(n1086) );
  NAND2X0_HVT U739 ( .A1(n217), .A2(n1080), .Y(n608) );
  NAND4X0_HVT U740 ( .A1(n551), .A2(n550), .A3(n253), .A4(n549), .Y(n1261) );
  AO22X1_HVT U741 ( .A1(n191), .A2(n397), .A3(n178), .A4(n258), .Y(n555) );
  AO221X1_HVT U742 ( .A1(sram_raddr_b0[0]), .A2(n1086), .A3(n242), .A4(n608), 
        .A5(n555), .Y(n560) );
  NAND2X0_HVT U743 ( .A1(n1550), .A2(n557), .Y(n1363) );
  AO22X1_HVT U744 ( .A1(n201), .A2(n560), .A3(sram_raddr_b0[0]), .A4(n169), 
        .Y(n_sram_raddr_b0[0]) );
  NAND2X0_HVT U745 ( .A1(sram_raddr_b3[0]), .A2(sram_raddr_b3[1]), .Y(n565) );
  NAND2X0_HVT U746 ( .A1(n258), .A2(n324), .Y(n1111) );
  NAND2X0_HVT U747 ( .A1(n565), .A2(n1111), .Y(n1085) );
  OA22X1_HVT U748 ( .A1(n1160), .A2(n322), .A3(n173), .A4(n1085), .Y(n562) );
  NAND2X0_HVT U749 ( .A1(sram_raddr_b6[1]), .A2(sram_raddr_b6[0]), .Y(n564) );
  OA21X1_HVT U750 ( .A1(sram_raddr_b6[1]), .A2(sram_raddr_b6[0]), .A3(n564), 
        .Y(n1084) );
  NAND2X0_HVT U751 ( .A1(n192), .A2(n1084), .Y(n806) );
  NAND2X0_HVT U752 ( .A1(sram_raddr_b0[0]), .A2(sram_raddr_b0[1]), .Y(n804) );
  NAND2X0_HVT U753 ( .A1(n242), .A2(n322), .Y(n829) );
  NAND3X0_HVT U754 ( .A1(n804), .A2(n608), .A3(n829), .Y(n561) );
  NAND3X0_HVT U755 ( .A1(n562), .A2(n806), .A3(n561), .Y(n563) );
  AO22X1_HVT U756 ( .A1(n204), .A2(n563), .A3(sram_raddr_b0[1]), .A4(n215), 
        .Y(n_sram_raddr_b0[1]) );
  NAND2X0_HVT U757 ( .A1(n239), .A2(n564), .Y(n568) );
  OA21X1_HVT U758 ( .A1(n564), .A2(n239), .A3(n568), .Y(n1091) );
  NAND2X0_HVT U759 ( .A1(n315), .A2(n565), .Y(n577) );
  OA21X1_HVT U760 ( .A1(n565), .A2(n315), .A3(n577), .Y(n809) );
  OA22X1_HVT U761 ( .A1(n1091), .A2(n1261), .A3(n809), .A4(n224), .Y(n812) );
  OA21X1_HVT U762 ( .A1(n622), .A2(n804), .A3(n213), .Y(n566) );
  NAND4X0_HVT U763 ( .A1(col[0]), .A2(n238), .A3(n312), .A4(n233), .Y(n1176)
         );
  NAND2X0_HVT U764 ( .A1(n217), .A2(n1176), .Y(n677) );
  NAND2X0_HVT U765 ( .A1(n706), .A2(n1200), .Y(n777) );
  NAND3X0_HVT U766 ( .A1(n566), .A2(n284), .A3(n777), .Y(n567) );
  NAND2X0_HVT U767 ( .A1(sram_raddr_b0[3]), .A2(n232), .Y(n574) );
  AND2X1_HVT U768 ( .A1(n214), .A2(n567), .Y(n569) );
  NAND2X0_HVT U769 ( .A1(n379), .A2(n569), .Y(n570) );
  NAND2X0_HVT U770 ( .A1(sram_raddr_b6[3]), .A2(n568), .Y(n590) );
  OA21X1_HVT U771 ( .A1(sram_raddr_b6[3]), .A2(n568), .A3(n590), .Y(n1097) );
  NAND2X0_HVT U772 ( .A1(n192), .A2(n1097), .Y(n820) );
  OA221X1_HVT U773 ( .A1(n690), .A2(n570), .A3(n569), .A4(n379), .A5(n820), 
        .Y(n571) );
  HADDX1_HVT U774 ( .A0(n343), .B0(n577), .SO(n817) );
  AO221X1_HVT U775 ( .A1(n571), .A2(n225), .A3(n571), .A4(n817), .A5(n219), 
        .Y(n573) );
  AO221X1_HVT U776 ( .A1(sram_raddr_b0[3]), .A2(sram_raddr_b0[2]), .A3(n379), 
        .A4(n284), .A5(n1368), .Y(n572) );
  NAND3X0_HVT U777 ( .A1(n574), .A2(n573), .A3(n572), .Y(n_sram_raddr_b0[3])
         );
  NAND2X0_HVT U778 ( .A1(sram_raddr_b0[3]), .A2(sram_raddr_b0[2]), .Y(n826) );
  NAND3X0_HVT U779 ( .A1(sram_raddr_b0[3]), .A2(sram_raddr_b0[0]), .A3(
        sram_raddr_b0[1]), .Y(n604) );
  AND3X1_HVT U780 ( .A1(n826), .A2(n256), .A3(n604), .Y(n576) );
  NAND3X0_HVT U781 ( .A1(col[1]), .A2(n721), .A3(n254), .Y(n1328) );
  NAND2X0_HVT U782 ( .A1(n826), .A2(n256), .Y(n585) );
  NAND3X0_HVT U783 ( .A1(sram_raddr_b0[3]), .A2(sram_raddr_b0[2]), .A3(
        sram_raddr_b0[4]), .Y(n597) );
  NAND2X0_HVT U784 ( .A1(n585), .A2(n597), .Y(n582) );
  AO22X1_HVT U785 ( .A1(n576), .A2(n608), .A3(n1150), .A4(n582), .Y(n589) );
  OA221X1_HVT U786 ( .A1(n622), .A2(n826), .A3(n622), .A4(n604), .A5(n211), 
        .Y(n586) );
  NAND2X0_HVT U787 ( .A1(sram_raddr_b3[3]), .A2(n577), .Y(n578) );
  NAND2X0_HVT U788 ( .A1(n578), .A2(n335), .Y(n587) );
  OA21X1_HVT U789 ( .A1(n335), .A2(n578), .A3(n587), .Y(n830) );
  OA22X1_HVT U790 ( .A1(n586), .A2(n256), .A3(n830), .A4(n224), .Y(n580) );
  AO22X1_HVT U791 ( .A1(n579), .A2(sram_raddr_b6[4]), .A3(n590), .A4(n280), 
        .Y(n1107) );
  NAND2X0_HVT U792 ( .A1(n190), .A2(n1107), .Y(n832) );
  NAND3X0_HVT U793 ( .A1(n581), .A2(n580), .A3(n832), .Y(n584) );
  AO222X1_HVT U794 ( .A1(n584), .A2(n203), .A3(n231), .A4(sram_raddr_b0[4]), 
        .A5(n223), .A6(n583), .Y(n_sram_raddr_b0[4]) );
  NAND2X0_HVT U795 ( .A1(n588), .A2(n268), .Y(n591) );
  OA21X1_HVT U796 ( .A1(n588), .A2(n268), .A3(n591), .Y(n837) );
  NAND3X0_HVT U797 ( .A1(n340), .A2(n597), .A3(n589), .Y(n593) );
  NAND3X0_HVT U798 ( .A1(n590), .A2(n363), .A3(n280), .Y(n592) );
  NAND2X0_HVT U799 ( .A1(n191), .A2(n1123), .Y(n840) );
  NAND4X0_HVT U800 ( .A1(sram_raddr_b0[3]), .A2(sram_raddr_b0[2]), .A3(
        sram_raddr_b0[5]), .A4(sram_raddr_b0[4]), .Y(n596) );
  NAND2X0_HVT U801 ( .A1(sram_raddr_b3[6]), .A2(n591), .Y(n602) );
  OA21X1_HVT U802 ( .A1(sram_raddr_b3[6]), .A2(n591), .A3(n602), .Y(n850) );
  NAND2X0_HVT U803 ( .A1(n850), .A2(n178), .Y(n595) );
  NAND2X0_HVT U804 ( .A1(sram_raddr_b6[6]), .A2(n592), .Y(n603) );
  OA21X1_HVT U805 ( .A1(sram_raddr_b6[6]), .A2(n592), .A3(n603), .Y(n1133) );
  NAND2X0_HVT U806 ( .A1(n190), .A2(n1133), .Y(n847) );
  NAND3X0_HVT U807 ( .A1(n826), .A2(n340), .A3(n256), .Y(n607) );
  AO222X1_HVT U808 ( .A1(n622), .A2(n605), .A3(n622), .A4(n1127), .A5(n605), 
        .A6(n604), .Y(n601) );
  OA222X1_HVT U809 ( .A1(n339), .A2(n213), .A3(n339), .A4(n593), .A5(
        sram_raddr_b0[6]), .A6(n601), .Y(n594) );
  NAND3X0_HVT U810 ( .A1(n595), .A2(n847), .A3(n594), .Y(n600) );
  AO221X1_HVT U811 ( .A1(n188), .A2(n339), .A3(n188), .A4(n596), .A5(n231), 
        .Y(n613) );
  NAND3X0_HVT U812 ( .A1(n223), .A2(sram_raddr_b0[5]), .A3(n828), .Y(n598) );
  NAND2X0_HVT U813 ( .A1(n339), .A2(n598), .Y(n599) );
  AO22X1_HVT U814 ( .A1(n202), .A2(n600), .A3(n613), .A4(n599), .Y(
        n_sram_raddr_b0[6]) );
  AND4X1_HVT U815 ( .A1(n188), .A2(sram_raddr_b0[6]), .A3(sram_raddr_b0[5]), 
        .A4(n828), .Y(n630) );
  OA21X1_HVT U816 ( .A1(n601), .A2(n339), .A3(n212), .Y(n609) );
  NAND2X0_HVT U817 ( .A1(n388), .A2(n602), .Y(n627) );
  OA21X1_HVT U818 ( .A1(n602), .A2(n388), .A3(n627), .Y(n861) );
  NAND2X0_HVT U819 ( .A1(n338), .A2(n603), .Y(n623) );
  NAND2X0_HVT U820 ( .A1(n192), .A2(n1145), .Y(n859) );
  NAND2X0_HVT U821 ( .A1(n605), .A2(n604), .Y(n606) );
  NAND2X0_HVT U822 ( .A1(sram_raddr_b0[6]), .A2(n606), .Y(n620) );
  NAND2X0_HVT U823 ( .A1(sram_raddr_b0[6]), .A2(n607), .Y(n618) );
  AO22X1_HVT U824 ( .A1(n608), .A2(n620), .A3(n1150), .A4(n618), .Y(n610) );
  HADDX1_HVT U825 ( .A0(sram_raddr_b3[8]), .B0(n627), .SO(n869) );
  OA22X1_HVT U826 ( .A1(n609), .A2(n346), .A3(n869), .A4(n225), .Y(n612) );
  HADDX1_HVT U827 ( .A0(n274), .B0(n623), .SO(n1157) );
  NAND2X0_HVT U828 ( .A1(n190), .A2(n1157), .Y(n872) );
  NAND3X0_HVT U829 ( .A1(n346), .A2(n269), .A3(n610), .Y(n626) );
  NAND3X0_HVT U830 ( .A1(sram_raddr_b0[8]), .A2(sram_raddr_b0[7]), .A3(n777), 
        .Y(n611) );
  NAND4X0_HVT U831 ( .A1(n612), .A2(n872), .A3(n626), .A4(n611), .Y(n616) );
  AO21X1_HVT U832 ( .A1(sram_raddr_b0[7]), .A2(n630), .A3(sram_raddr_b0[8]), 
        .Y(n615) );
  NAND2X0_HVT U833 ( .A1(sram_raddr_b0[8]), .A2(sram_raddr_b0[7]), .Y(n614) );
  AO21X1_HVT U834 ( .A1(n614), .A2(n169), .A3(n613), .Y(n617) );
  AO22X1_HVT U835 ( .A1(n204), .A2(n616), .A3(n615), .A4(n617), .Y(
        n_sram_raddr_b0[8]) );
  NAND2X0_HVT U836 ( .A1(sram_raddr_b0[9]), .A2(n617), .Y(n633) );
  AND2X1_HVT U837 ( .A1(n346), .A2(n269), .Y(n621) );
  OA221X1_HVT U838 ( .A1(n1127), .A2(n621), .A3(n1127), .A4(n618), .A5(n214), 
        .Y(n619) );
  OA221X1_HVT U839 ( .A1(n622), .A2(n621), .A3(n622), .A4(n620), .A5(n619), 
        .Y(n625) );
  OR2X1_HVT U840 ( .A1(n623), .A2(sram_raddr_b6[8]), .Y(n624) );
  HADDX1_HVT U841 ( .A0(n624), .B0(n373), .SO(n1165) );
  NAND2X0_HVT U842 ( .A1(n190), .A2(n1165), .Y(n884) );
  OA221X1_HVT U843 ( .A1(sram_raddr_b0[9]), .A2(n626), .A3(n401), .A4(n625), 
        .A5(n884), .Y(n629) );
  OR2X1_HVT U844 ( .A1(n627), .A2(sram_raddr_b3[8]), .Y(n628) );
  HADDX1_HVT U845 ( .A0(sram_raddr_b3[9]), .B0(n628), .SO(n885) );
  AO221X1_HVT U846 ( .A1(n629), .A2(n224), .A3(n629), .A4(n885), .A5(n226), 
        .Y(n632) );
  NAND4X0_HVT U847 ( .A1(sram_raddr_b0[7]), .A2(sram_raddr_b0[8]), .A3(n630), 
        .A4(n401), .Y(n631) );
  NAND3X0_HVT U848 ( .A1(n633), .A2(n632), .A3(n631), .Y(n_sram_raddr_b0[9])
         );
  NAND2X0_HVT U849 ( .A1(col[0]), .A2(n212), .Y(n1238) );
  AO22X1_HVT U850 ( .A1(n192), .A2(n398), .A3(n178), .A4(n259), .Y(n634) );
  AO221X1_HVT U851 ( .A1(sram_raddr_b1[0]), .A2(n1238), .A3(n243), .A4(n677), 
        .A5(n634), .Y(n635) );
  AO22X1_HVT U852 ( .A1(n204), .A2(n635), .A3(sram_raddr_b1[0]), .A4(n169), 
        .Y(n_sram_raddr_b1[0]) );
  NAND2X0_HVT U853 ( .A1(sram_raddr_b4[0]), .A2(sram_raddr_b4[1]), .Y(n639) );
  NAND2X0_HVT U854 ( .A1(n259), .A2(n326), .Y(n1205) );
  NAND2X0_HVT U855 ( .A1(n639), .A2(n1205), .Y(n1181) );
  OA22X1_HVT U856 ( .A1(n895), .A2(n323), .A3(n224), .A4(n1181), .Y(n637) );
  NAND2X0_HVT U857 ( .A1(sram_raddr_b7[1]), .A2(sram_raddr_b7[0]), .Y(n646) );
  OA21X1_HVT U858 ( .A1(sram_raddr_b7[1]), .A2(sram_raddr_b7[0]), .A3(n646), 
        .Y(n1180) );
  NAND2X0_HVT U859 ( .A1(n192), .A2(n1180), .Y(n898) );
  NAND2X0_HVT U860 ( .A1(sram_raddr_b1[0]), .A2(sram_raddr_b1[1]), .Y(n896) );
  NAND2X0_HVT U861 ( .A1(n243), .A2(n323), .Y(n901) );
  NAND3X0_HVT U862 ( .A1(n677), .A2(n896), .A3(n901), .Y(n636) );
  NAND3X0_HVT U863 ( .A1(n637), .A2(n898), .A3(n636), .Y(n638) );
  AO22X1_HVT U864 ( .A1(n203), .A2(n638), .A3(sram_raddr_b1[1]), .A4(n215), 
        .Y(n_sram_raddr_b1[1]) );
  OA21X1_HVT U865 ( .A1(n706), .A2(n896), .A3(n214), .Y(n640) );
  NAND2X0_HVT U866 ( .A1(n314), .A2(n639), .Y(n655) );
  OA21X1_HVT U867 ( .A1(n639), .A2(n314), .A3(n655), .Y(n903) );
  OA22X1_HVT U868 ( .A1(n640), .A2(n277), .A3(n903), .A4(n224), .Y(n642) );
  NAND3X0_HVT U869 ( .A1(n640), .A2(n777), .A3(n277), .Y(n645) );
  AO22X1_HVT U870 ( .A1(sram_raddr_b7[2]), .A2(n641), .A3(n240), .A4(n646), 
        .Y(n1186) );
  NAND2X0_HVT U871 ( .A1(n191), .A2(n1186), .Y(n902) );
  NAND3X0_HVT U872 ( .A1(n642), .A2(n645), .A3(n902), .Y(n643) );
  AO22X1_HVT U873 ( .A1(n201), .A2(n643), .A3(n221), .A4(n277), .Y(n644) );
  AO21X1_HVT U874 ( .A1(n230), .A2(sram_raddr_b1[2]), .A3(n644), .Y(
        n_sram_raddr_b1[2]) );
  NAND2X0_HVT U875 ( .A1(sram_raddr_b1[3]), .A2(n231), .Y(n653) );
  AO221X1_HVT U876 ( .A1(sram_raddr_b1[3]), .A2(sram_raddr_b1[2]), .A3(n386), 
        .A4(n277), .A5(n1368), .Y(n652) );
  AND2X1_HVT U877 ( .A1(n213), .A2(n645), .Y(n648) );
  NAND2X0_HVT U878 ( .A1(n386), .A2(n648), .Y(n649) );
  NAND2X0_HVT U879 ( .A1(n240), .A2(n646), .Y(n647) );
  NAND2X0_HVT U880 ( .A1(sram_raddr_b7[3]), .A2(n647), .Y(n668) );
  OA21X1_HVT U881 ( .A1(sram_raddr_b7[3]), .A2(n647), .A3(n668), .Y(n1191) );
  NAND2X0_HVT U882 ( .A1(n190), .A2(n1191), .Y(n910) );
  OA221X1_HVT U883 ( .A1(n690), .A2(n649), .A3(n648), .A4(n386), .A5(n910), 
        .Y(n650) );
  HADDX1_HVT U884 ( .A0(n336), .B0(n655), .SO(n909) );
  AO221X1_HVT U885 ( .A1(n650), .A2(n173), .A3(n650), .A4(n909), .A5(n226), 
        .Y(n651) );
  NAND3X0_HVT U886 ( .A1(n653), .A2(n652), .A3(n651), .Y(n_sram_raddr_b1[3])
         );
  NAND3X0_HVT U887 ( .A1(sram_raddr_b1[3]), .A2(sram_raddr_b1[2]), .A3(
        sram_raddr_b1[4]), .Y(n913) );
  NAND2X0_HVT U888 ( .A1(sram_raddr_b1[3]), .A2(sram_raddr_b1[2]), .Y(n912) );
  NAND2X0_HVT U889 ( .A1(n912), .A2(n316), .Y(n663) );
  NAND2X0_HVT U890 ( .A1(n913), .A2(n663), .Y(n660) );
  NAND3X0_HVT U891 ( .A1(sram_raddr_b1[3]), .A2(sram_raddr_b1[0]), .A3(
        sram_raddr_b1[1]), .Y(n674) );
  AND3X1_HVT U892 ( .A1(n912), .A2(n316), .A3(n674), .Y(n654) );
  AO22X1_HVT U893 ( .A1(n1228), .A2(n660), .A3(n654), .A4(n677), .Y(n667) );
  OA221X1_HVT U894 ( .A1(n706), .A2(n912), .A3(n706), .A4(n674), .A5(n211), 
        .Y(n664) );
  NAND2X0_HVT U895 ( .A1(sram_raddr_b4[3]), .A2(n655), .Y(n656) );
  NAND2X0_HVT U896 ( .A1(n656), .A2(n357), .Y(n665) );
  OA21X1_HVT U897 ( .A1(n357), .A2(n656), .A3(n665), .Y(n911) );
  OA22X1_HVT U898 ( .A1(n664), .A2(n316), .A3(n911), .A4(n225), .Y(n658) );
  AO22X1_HVT U899 ( .A1(n657), .A2(sram_raddr_b7[4]), .A3(n668), .A4(n281), 
        .Y(n1201) );
  NAND2X0_HVT U900 ( .A1(n192), .A2(n1201), .Y(n916) );
  NAND3X0_HVT U901 ( .A1(n659), .A2(n658), .A3(n916), .Y(n662) );
  AO222X1_HVT U902 ( .A1(n662), .A2(n204), .A3(n232), .A4(sram_raddr_b1[4]), 
        .A5(n221), .A6(n661), .Y(n_sram_raddr_b1[4]) );
  NAND2X0_HVT U903 ( .A1(n666), .A2(n276), .Y(n670) );
  OA21X1_HVT U904 ( .A1(n666), .A2(n276), .A3(n670), .Y(n925) );
  NAND3X0_HVT U905 ( .A1(n270), .A2(n913), .A3(n667), .Y(n669) );
  NAND3X0_HVT U906 ( .A1(n668), .A2(n364), .A3(n281), .Y(n671) );
  NAND2X0_HVT U907 ( .A1(n190), .A2(n1214), .Y(n924) );
  NAND4X0_HVT U908 ( .A1(sram_raddr_b1[3]), .A2(sram_raddr_b1[2]), .A3(
        sram_raddr_b1[5]), .A4(sram_raddr_b1[4]), .Y(n672) );
  NAND3X0_HVT U909 ( .A1(n912), .A2(n270), .A3(n316), .Y(n673) );
  NAND2X0_HVT U910 ( .A1(sram_raddr_b4[6]), .A2(n670), .Y(n679) );
  NAND2X0_HVT U911 ( .A1(sram_raddr_b7[6]), .A2(n671), .Y(n680) );
  OA21X1_HVT U912 ( .A1(sram_raddr_b7[6]), .A2(n671), .A3(n680), .Y(n1220) );
  NAND2X0_HVT U913 ( .A1(n190), .A2(n1220), .Y(n934) );
  OR3X1_HVT U915 ( .A1(n344), .A2(n270), .A3(n913), .Y(n683) );
  NAND2X0_HVT U916 ( .A1(sram_raddr_b1[6]), .A2(n673), .Y(n702) );
  NAND2X0_HVT U917 ( .A1(n675), .A2(n674), .Y(n676) );
  NAND2X0_HVT U918 ( .A1(sram_raddr_b1[6]), .A2(n676), .Y(n704) );
  AO22X1_HVT U919 ( .A1(n1228), .A2(n702), .A3(n677), .A4(n704), .Y(n688) );
  NAND2X0_HVT U920 ( .A1(n688), .A2(n333), .Y(n682) );
  AND2X1_HVT U921 ( .A1(n1228), .A2(n702), .Y(n678) );
  OA22X1_HVT U922 ( .A1(n895), .A2(n678), .A3(n706), .A4(n704), .Y(n691) );
  NAND2X0_HVT U923 ( .A1(n332), .A2(n679), .Y(n692) );
  OA21X1_HVT U924 ( .A1(n679), .A2(n332), .A3(n692), .Y(n939) );
  OA22X1_HVT U925 ( .A1(n691), .A2(n333), .A3(n939), .A4(n173), .Y(n681) );
  NAND2X0_HVT U926 ( .A1(n347), .A2(n680), .Y(n689) );
  NAND2X0_HVT U927 ( .A1(n192), .A2(n1231), .Y(n942) );
  NAND3X0_HVT U928 ( .A1(n682), .A2(n681), .A3(n942), .Y(n687) );
  NAND2X0_HVT U929 ( .A1(n333), .A2(n683), .Y(n686) );
  NAND2X0_HVT U930 ( .A1(sram_raddr_b1[7]), .A2(n696), .Y(n684) );
  NAND2X0_HVT U931 ( .A1(n221), .A2(n684), .Y(n695) );
  AO222X1_HVT U932 ( .A1(n687), .A2(n201), .A3(n686), .A4(n685), .A5(
        sram_raddr_b1[7]), .A6(n231), .Y(n_sram_raddr_b1[7]) );
  NAND3X0_HVT U933 ( .A1(n333), .A2(n272), .A3(n688), .Y(n710) );
  AO22X1_HVT U934 ( .A1(sram_raddr_b7[8]), .A2(n689), .A3(n391), .A4(n707), 
        .Y(n1242) );
  NAND2X0_HVT U935 ( .A1(n190), .A2(n1242), .Y(n955) );
  AO221X1_HVT U936 ( .A1(n691), .A2(n690), .A3(n691), .A4(n333), .A5(n272), 
        .Y(n694) );
  AO22X1_HVT U937 ( .A1(sram_raddr_b4[8]), .A2(n692), .A3(n345), .A4(n711), 
        .Y(n956) );
  NAND2X0_HVT U938 ( .A1(n178), .A2(n956), .Y(n693) );
  NAND4X0_HVT U939 ( .A1(n710), .A2(n955), .A3(n694), .A4(n693), .Y(n699) );
  NAND3X0_HVT U940 ( .A1(n223), .A2(sram_raddr_b1[7]), .A3(n696), .Y(n701) );
  NAND2X0_HVT U941 ( .A1(n272), .A2(n701), .Y(n697) );
  AO22X1_HVT U942 ( .A1(n205), .A2(n699), .A3(n698), .A4(n697), .Y(
        n_sram_raddr_b1[8]) );
  AO222X1_HVT U943 ( .A1(n377), .A2(n272), .A3(n377), .A4(n701), .A5(
        sram_raddr_b1[9]), .A6(n700), .Y(n715) );
  AND2X1_HVT U944 ( .A1(n333), .A2(n272), .Y(n705) );
  OA221X1_HVT U945 ( .A1(col[0]), .A2(n705), .A3(col[0]), .A4(n702), .A5(n212), 
        .Y(n703) );
  OA221X1_HVT U946 ( .A1(n706), .A2(n705), .A3(n706), .A4(n704), .A5(n703), 
        .Y(n709) );
  NAND2X0_HVT U947 ( .A1(n707), .A2(n391), .Y(n708) );
  HADDX1_HVT U948 ( .A0(n372), .B0(n708), .SO(n1251) );
  NAND2X0_HVT U949 ( .A1(n192), .A2(n1251), .Y(n968) );
  OA221X1_HVT U950 ( .A1(sram_raddr_b1[9]), .A2(n710), .A3(n377), .A4(n709), 
        .A5(n968), .Y(n713) );
  NAND2X0_HVT U951 ( .A1(n711), .A2(n345), .Y(n712) );
  HADDX1_HVT U952 ( .A0(sram_raddr_b4[9]), .B0(n712), .SO(n969) );
  AO221X1_HVT U953 ( .A1(n713), .A2(n224), .A3(n713), .A4(n969), .A5(n219), 
        .Y(n714) );
  NAND2X0_HVT U954 ( .A1(n715), .A2(n714), .Y(n_sram_raddr_b1[9]) );
  AO22X1_HVT U955 ( .A1(n191), .A2(n399), .A3(n1322), .A4(n244), .Y(n716) );
  AO221X1_HVT U956 ( .A1(sram_raddr_b2[0]), .A2(n1334), .A3(n260), .A4(n787), 
        .A5(n716), .Y(n717) );
  AO22X1_HVT U957 ( .A1(n205), .A2(n717), .A3(sram_raddr_b2[0]), .A4(n169), 
        .Y(n_sram_raddr_b2[0]) );
  NAND2X0_HVT U958 ( .A1(sram_raddr_b5[0]), .A2(sram_raddr_b5[1]), .Y(n731) );
  NAND2X0_HVT U959 ( .A1(n244), .A2(n327), .Y(n1293) );
  NAND2X0_HVT U960 ( .A1(n731), .A2(n1293), .Y(n1267) );
  OA22X1_HVT U961 ( .A1(n978), .A2(n325), .A3(n225), .A4(n1267), .Y(n719) );
  NAND2X0_HVT U962 ( .A1(sram_raddr_b8[1]), .A2(sram_raddr_b8[0]), .Y(n728) );
  OA21X1_HVT U963 ( .A1(sram_raddr_b8[1]), .A2(sram_raddr_b8[0]), .A3(n728), 
        .Y(n1266) );
  NAND2X0_HVT U964 ( .A1(n191), .A2(n1266), .Y(n981) );
  NAND2X0_HVT U965 ( .A1(sram_raddr_b2[0]), .A2(sram_raddr_b2[1]), .Y(n979) );
  NAND2X0_HVT U966 ( .A1(n260), .A2(n325), .Y(n1001) );
  NAND3X0_HVT U967 ( .A1(n787), .A2(n979), .A3(n1001), .Y(n718) );
  NAND3X0_HVT U968 ( .A1(n719), .A2(n981), .A3(n718), .Y(n720) );
  AO22X1_HVT U969 ( .A1(n1558), .A2(n720), .A3(sram_raddr_b2[1]), .A4(n215), 
        .Y(n_sram_raddr_b2[1]) );
  NAND2X0_HVT U970 ( .A1(n354), .A2(n979), .Y(n734) );
  OA22X1_HVT U971 ( .A1(sram_raddr_b2[2]), .A2(n1301), .A3(n744), .A4(n734), 
        .Y(n727) );
  AO22X1_HVT U972 ( .A1(sram_raddr_b8[2]), .A2(n722), .A3(n241), .A4(n728), 
        .Y(n1273) );
  NAND2X0_HVT U973 ( .A1(n190), .A2(n1273), .Y(n984) );
  AO221X1_HVT U974 ( .A1(n211), .A2(n744), .A3(n212), .A4(n979), .A5(n354), 
        .Y(n723) );
  NAND3X0_HVT U975 ( .A1(n727), .A2(n984), .A3(n723), .Y(n725) );
  AO22X1_HVT U976 ( .A1(sram_raddr_b5[2]), .A2(n724), .A3(n313), .A4(n731), 
        .Y(n986) );
  OA221X1_HVT U977 ( .A1(n725), .A2(n178), .A3(n725), .A4(n986), .A5(n205), 
        .Y(n726) );
  AO221X1_HVT U978 ( .A1(sram_raddr_b2[2]), .A2(n230), .A3(n354), .A4(n222), 
        .A5(n726), .Y(n_sram_raddr_b2[2]) );
  NAND2X0_HVT U979 ( .A1(n213), .A2(n727), .Y(n730) );
  OA221X1_HVT U980 ( .A1(n787), .A2(sram_raddr_b2[2]), .A3(n787), .A4(n1320), 
        .A5(n734), .Y(n729) );
  NAND2X0_HVT U981 ( .A1(n241), .A2(n728), .Y(n1277) );
  NAND2X0_HVT U982 ( .A1(sram_raddr_b8[3]), .A2(n1277), .Y(n1276) );
  AO221X1_HVT U983 ( .A1(sram_raddr_b2[3]), .A2(n730), .A3(n406), .A4(n729), 
        .A5(n993), .Y(n733) );
  NAND2X0_HVT U984 ( .A1(n313), .A2(n731), .Y(n732) );
  NAND2X0_HVT U985 ( .A1(sram_raddr_b5[3]), .A2(n732), .Y(n736) );
  OA21X1_HVT U986 ( .A1(sram_raddr_b5[3]), .A2(n732), .A3(n736), .Y(n992) );
  NAND2X0_HVT U987 ( .A1(sram_raddr_b2[3]), .A2(sram_raddr_b2[2]), .Y(n998) );
  NAND2X0_HVT U988 ( .A1(n255), .A2(n998), .Y(n742) );
  NAND3X0_HVT U989 ( .A1(sram_raddr_b2[4]), .A2(sram_raddr_b2[3]), .A3(
        sram_raddr_b2[2]), .Y(n763) );
  NAND2X0_HVT U990 ( .A1(n742), .A2(n763), .Y(n739) );
  NAND2X0_HVT U991 ( .A1(sram_raddr_b2[3]), .A2(n734), .Y(n756) );
  AND2X1_HVT U992 ( .A1(n255), .A2(n756), .Y(n735) );
  AO22X1_HVT U993 ( .A1(n1320), .A2(n739), .A3(n735), .A4(n787), .Y(n749) );
  OA21X1_HVT U994 ( .A1(n744), .A2(n756), .A3(n211), .Y(n745) );
  NAND2X0_HVT U995 ( .A1(n341), .A2(n736), .Y(n746) );
  OA21X1_HVT U996 ( .A1(n736), .A2(n341), .A3(n746), .Y(n1002) );
  OA22X1_HVT U997 ( .A1(n745), .A2(n255), .A3(n1002), .A4(n173), .Y(n737) );
  NAND2X0_HVT U998 ( .A1(n381), .A2(n1276), .Y(n750) );
  NAND2X0_HVT U999 ( .A1(n191), .A2(n1289), .Y(n1004) );
  NAND3X0_HVT U1000 ( .A1(n738), .A2(n737), .A3(n1004), .Y(n741) );
  AO222X1_HVT U1001 ( .A1(n741), .A2(n205), .A3(n232), .A4(sram_raddr_b2[4]), 
        .A5(n222), .A6(n740), .Y(n_sram_raddr_b2[4]) );
  NAND2X0_HVT U1002 ( .A1(n312), .A2(n742), .Y(n743) );
  NAND2X0_HVT U1003 ( .A1(n747), .A2(n271), .Y(n755) );
  OA21X1_HVT U1004 ( .A1(n747), .A2(n271), .A3(n755), .Y(n1012) );
  OA22X1_HVT U1005 ( .A1(n748), .A2(n334), .A3(n1012), .A4(n173), .Y(n751) );
  NAND3X0_HVT U1006 ( .A1(n334), .A2(n763), .A3(n749), .Y(n757) );
  AO22X1_HVT U1007 ( .A1(sram_raddr_b8[5]), .A2(n750), .A3(n342), .A4(n758), 
        .Y(n1302) );
  NAND2X0_HVT U1008 ( .A1(n190), .A2(n1302), .Y(n1011) );
  NAND3X0_HVT U1009 ( .A1(n751), .A2(n757), .A3(n1011), .Y(n752) );
  AO22X1_HVT U1010 ( .A1(n203), .A2(n752), .A3(n231), .A4(sram_raddr_b2[5]), 
        .Y(n754) );
  NAND4X0_HVT U1011 ( .A1(sram_raddr_b2[5]), .A2(sram_raddr_b2[4]), .A3(
        sram_raddr_b2[3]), .A4(sram_raddr_b2[2]), .Y(n762) );
  NAND2X0_HVT U1012 ( .A1(n334), .A2(n763), .Y(n753) );
  OA222X1_HVT U1013 ( .A1(n754), .A2(n223), .A3(n754), .A4(n762), .A5(n754), 
        .A6(n753), .Y(n_sram_raddr_b2[5]) );
  NAND2X0_HVT U1014 ( .A1(sram_raddr_b5[6]), .A2(n755), .Y(n768) );
  OA21X1_HVT U1015 ( .A1(sram_raddr_b5[6]), .A2(n755), .A3(n768), .Y(n1025) );
  NAND2X0_HVT U1016 ( .A1(n1025), .A2(n1322), .Y(n761) );
  NAND3X0_HVT U1017 ( .A1(n334), .A2(n255), .A3(n998), .Y(n771) );
  NAND3X0_HVT U1018 ( .A1(n334), .A2(n255), .A3(n756), .Y(n772) );
  AOI22X1_HVT U1019 ( .A1(n1320), .A2(n771), .A3(n787), .A4(n772), .Y(n767) );
  OA222X1_HVT U1020 ( .A1(n337), .A2(n211), .A3(n337), .A4(n757), .A5(
        sram_raddr_b2[6]), .A6(n767), .Y(n760) );
  NAND2X0_HVT U1021 ( .A1(n758), .A2(n342), .Y(n759) );
  NAND2X0_HVT U1022 ( .A1(sram_raddr_b8[6]), .A2(n759), .Y(n769) );
  OA21X1_HVT U1023 ( .A1(sram_raddr_b8[6]), .A2(n759), .A3(n769), .Y(n1310) );
  NAND2X0_HVT U1024 ( .A1(n190), .A2(n1310), .Y(n1032) );
  NAND3X0_HVT U1025 ( .A1(n761), .A2(n760), .A3(n1032), .Y(n766) );
  AO221X1_HVT U1026 ( .A1(n223), .A2(n337), .A3(n188), .A4(n762), .A5(n232), 
        .Y(n780) );
  NAND3X0_HVT U1027 ( .A1(n221), .A2(sram_raddr_b2[5]), .A3(n1000), .Y(n764)
         );
  NAND2X0_HVT U1028 ( .A1(n337), .A2(n764), .Y(n765) );
  AO22X1_HVT U1029 ( .A1(n205), .A2(n766), .A3(n780), .A4(n765), .Y(
        n_sram_raddr_b2[6]) );
  AND4X1_HVT U1030 ( .A1(n188), .A2(sram_raddr_b2[6]), .A3(sram_raddr_b2[5]), 
        .A4(n1000), .Y(n798) );
  OA21X1_HVT U1031 ( .A1(n767), .A2(n337), .A3(n214), .Y(n775) );
  NAND2X0_HVT U1032 ( .A1(n393), .A2(n768), .Y(n789) );
  OA21X1_HVT U1033 ( .A1(n768), .A2(n393), .A3(n789), .Y(n1037) );
  OA22X1_HVT U1034 ( .A1(n775), .A2(n267), .A3(n1037), .A4(n224), .Y(n770) );
  NAND2X0_HVT U1035 ( .A1(n275), .A2(n769), .Y(n792) );
  NAND2X0_HVT U1036 ( .A1(n191), .A2(n1315), .Y(n1039) );
  NAND2X0_HVT U1037 ( .A1(n770), .A2(n1039), .Y(n773) );
  NAND2X0_HVT U1038 ( .A1(sram_raddr_b2[6]), .A2(n771), .Y(n784) );
  NAND2X0_HVT U1039 ( .A1(sram_raddr_b2[6]), .A2(n772), .Y(n783) );
  AO22X1_HVT U1040 ( .A1(n1320), .A2(n784), .A3(n787), .A4(n783), .Y(n776) );
  OA221X1_HVT U1041 ( .A1(n773), .A2(n267), .A3(n773), .A4(n776), .A5(n201), 
        .Y(n774) );
  AO221X1_HVT U1042 ( .A1(sram_raddr_b2[7]), .A2(n780), .A3(n267), .A4(n798), 
        .A5(n774), .Y(n_sram_raddr_b2[7]) );
  HADDX1_HVT U1043 ( .A0(sram_raddr_b5[8]), .B0(n789), .SO(n1049) );
  OA22X1_HVT U1044 ( .A1(n1049), .A2(n224), .A3(n775), .A4(n360), .Y(n779) );
  HADDX1_HVT U1045 ( .A0(n359), .B0(n792), .SO(n1329) );
  NAND2X0_HVT U1046 ( .A1(n191), .A2(n1329), .Y(n1047) );
  NAND3X0_HVT U1047 ( .A1(n360), .A2(n267), .A3(n776), .Y(n791) );
  NAND3X0_HVT U1048 ( .A1(sram_raddr_b2[8]), .A2(sram_raddr_b2[7]), .A3(n777), 
        .Y(n778) );
  NAND4X0_HVT U1049 ( .A1(n779), .A2(n1047), .A3(n791), .A4(n778), .Y(n782) );
  AO21X1_HVT U1050 ( .A1(sram_raddr_b2[7]), .A2(n798), .A3(sram_raddr_b2[8]), 
        .Y(n781) );
  NAND2X0_HVT U1051 ( .A1(sram_raddr_b2[8]), .A2(sram_raddr_b2[7]), .Y(n796)
         );
  AO21X1_HVT U1052 ( .A1(n188), .A2(n796), .A3(n780), .Y(n797) );
  AO22X1_HVT U1053 ( .A1(n1558), .A2(n782), .A3(n781), .A4(n797), .Y(
        n_sram_raddr_b2[8]) );
  NAND3X0_HVT U1054 ( .A1(n360), .A2(n267), .A3(n783), .Y(n786) );
  NAND4X0_HVT U1055 ( .A1(n212), .A2(n267), .A3(n360), .A4(n784), .Y(n785) );
  AO22X1_HVT U1056 ( .A1(n787), .A2(n786), .A3(n1334), .A4(n785), .Y(n788) );
  NAND2X0_HVT U1057 ( .A1(sram_raddr_b2[9]), .A2(n788), .Y(n795) );
  OR2X1_HVT U1058 ( .A1(n789), .A2(sram_raddr_b5[8]), .Y(n790) );
  HADDX1_HVT U1059 ( .A0(sram_raddr_b5[9]), .B0(n790), .SO(n1072) );
  OA22X1_HVT U1060 ( .A1(sram_raddr_b2[9]), .A2(n791), .A3(n225), .A4(n1072), 
        .Y(n794) );
  OR2X1_HVT U1061 ( .A1(n792), .A2(sram_raddr_b8[8]), .Y(n793) );
  HADDX1_HVT U1062 ( .A0(n793), .B0(n374), .SO(n1339) );
  NAND2X0_HVT U1063 ( .A1(n190), .A2(n1339), .Y(n1071) );
  NAND3X0_HVT U1064 ( .A1(n795), .A2(n794), .A3(n1071), .Y(n801) );
  OA222X1_HVT U1065 ( .A1(sram_raddr_b2[9]), .A2(n799), .A3(sram_raddr_b2[9]), 
        .A4(n798), .A5(n419), .A6(n797), .Y(n800) );
  AO21X1_HVT U1066 ( .A1(n204), .A2(n801), .A3(n800), .Y(n_sram_raddr_b2[9])
         );
  NAND2X0_HVT U1067 ( .A1(n1080), .A2(n173), .Y(n863) );
  AO22X1_HVT U1068 ( .A1(n192), .A2(n397), .A3(n1262), .A4(n242), .Y(n802) );
  AO221X1_HVT U1069 ( .A1(sram_raddr_b3[0]), .A2(n1086), .A3(n258), .A4(n863), 
        .A5(n802), .Y(n803) );
  AO22X1_HVT U1070 ( .A1(n1558), .A2(n803), .A3(sram_raddr_b3[0]), .A4(n215), 
        .Y(n_sram_raddr_b3[0]) );
  OA22X1_HVT U1071 ( .A1(n886), .A2(n1085), .A3(n1160), .A4(n324), .Y(n807) );
  NAND2X0_HVT U1072 ( .A1(n804), .A2(n829), .Y(n805) );
  NAND2X0_HVT U1073 ( .A1(n1262), .A2(n805), .Y(n1083) );
  NAND3X0_HVT U1074 ( .A1(n807), .A2(n806), .A3(n1083), .Y(n808) );
  AO22X1_HVT U1075 ( .A1(n201), .A2(n808), .A3(sram_raddr_b3[1]), .A4(n169), 
        .Y(n_sram_raddr_b3[1]) );
  OA22X1_HVT U1076 ( .A1(sram_raddr_b3[2]), .A2(n1127), .A3(n809), .A4(n1080), 
        .Y(n811) );
  NAND2X0_HVT U1077 ( .A1(sram_raddr_b3[2]), .A2(n1308), .Y(n810) );
  AO221X1_HVT U1078 ( .A1(sram_raddr_b0[2]), .A2(n829), .A3(n284), .A4(n827), 
        .A5(n218), .Y(n1088) );
  NAND4X0_HVT U1079 ( .A1(n812), .A2(n811), .A3(n810), .A4(n1088), .Y(n815) );
  NAND2X0_HVT U1080 ( .A1(n188), .A2(n315), .Y(n813) );
  NAND2X0_HVT U1081 ( .A1(n1305), .A2(n813), .Y(n824) );
  NAND2X0_HVT U1082 ( .A1(n315), .A2(n1368), .Y(n814) );
  AO22X1_HVT U1083 ( .A1(n1558), .A2(n815), .A3(n824), .A4(n814), .Y(
        n_sram_raddr_b3[2]) );
  OA21X1_HVT U1084 ( .A1(sram_raddr_b3[2]), .A2(n1127), .A3(n213), .Y(n816) );
  OA22X1_HVT U1085 ( .A1(n886), .A2(n817), .A3(n816), .A4(n343), .Y(n821) );
  OA222X1_HVT U1086 ( .A1(sram_raddr_b0[3]), .A2(sram_raddr_b0[2]), .A3(
        sram_raddr_b0[3]), .A4(n829), .A5(n827), .A6(n826), .Y(n818) );
  NAND2X0_HVT U1087 ( .A1(n1262), .A2(n818), .Y(n1102) );
  NAND3X0_HVT U1088 ( .A1(sram_raddr_b3[2]), .A2(n343), .A3(n1150), .Y(n819)
         );
  NAND4X0_HVT U1089 ( .A1(n821), .A2(n820), .A3(n1102), .A4(n819), .Y(n823) );
  AND2X1_HVT U1090 ( .A1(sram_raddr_b3[2]), .A2(n343), .Y(n822) );
  AO222X1_HVT U1091 ( .A1(n824), .A2(sram_raddr_b3[3]), .A3(n823), .A4(n204), 
        .A5(n822), .A6(n222), .Y(n_sram_raddr_b3[3]) );
  NAND3X0_HVT U1092 ( .A1(sram_raddr_b3[3]), .A2(sram_raddr_b3[2]), .A3(
        sram_raddr_b3[4]), .Y(n843) );
  NAND2X0_HVT U1093 ( .A1(sram_raddr_b3[3]), .A2(sram_raddr_b3[2]), .Y(n1108)
         );
  NAND2X0_HVT U1094 ( .A1(n335), .A2(n1108), .Y(n825) );
  AND2X1_HVT U1095 ( .A1(n843), .A2(n825), .Y(n834) );
  OA22X1_HVT U1096 ( .A1(n1127), .A2(n834), .A3(n213), .A4(n335), .Y(n833) );
  OA21X1_HVT U1097 ( .A1(n827), .A2(n826), .A3(n256), .Y(n838) );
  OAI221X1_HVT U1098 ( .A1(n838), .A2(n829), .A3(n838), .A4(n828), .A5(n1262), 
        .Y(n1114) );
  OR2X1_HVT U1099 ( .A1(n886), .A2(n830), .Y(n831) );
  NAND4X0_HVT U1100 ( .A1(n833), .A2(n832), .A3(n1114), .A4(n831), .Y(n835) );
  AO222X1_HVT U1101 ( .A1(n835), .A2(n204), .A3(n230), .A4(sram_raddr_b3[4]), 
        .A5(n223), .A6(n834), .Y(n_sram_raddr_b3[4]) );
  OA221X1_HVT U1102 ( .A1(n1389), .A2(n335), .A3(n1389), .A4(n1108), .A5(n213), 
        .Y(n836) );
  OA22X1_HVT U1103 ( .A1(n886), .A2(n837), .A3(n268), .A4(n836), .Y(n841) );
  NAND3X0_HVT U1104 ( .A1(n268), .A2(n335), .A3(n1108), .Y(n856) );
  OR2X1_HVT U1105 ( .A1(n856), .A2(n1127), .Y(n839) );
  NAND2X0_HVT U1106 ( .A1(n838), .A2(n340), .Y(n846) );
  AO221X1_HVT U1107 ( .A1(n846), .A2(n838), .A3(n846), .A4(n340), .A5(n218), 
        .Y(n1121) );
  AND4X1_HVT U1108 ( .A1(n841), .A2(n840), .A3(n839), .A4(n1121), .Y(n842) );
  OA22X1_HVT U1109 ( .A1(n842), .A2(n219), .A3(n1305), .A4(n268), .Y(n845) );
  AO221X1_HVT U1110 ( .A1(sram_raddr_b3[5]), .A2(n1110), .A3(n268), .A4(n843), 
        .A5(n1368), .Y(n844) );
  NAND2X0_HVT U1111 ( .A1(n845), .A2(n844), .Y(n_sram_raddr_b3[5]) );
  NAND2X0_HVT U1112 ( .A1(sram_raddr_b0[6]), .A2(n846), .Y(n857) );
  NAND2X0_HVT U1113 ( .A1(n1262), .A2(n857), .Y(n849) );
  OA221X1_HVT U1114 ( .A1(n849), .A2(n848), .A3(n849), .A4(n339), .A5(n847), 
        .Y(n1132) );
  AO221X1_HVT U1115 ( .A1(n211), .A2(n1127), .A3(n214), .A4(n856), .A5(n358), 
        .Y(n853) );
  NAND2X0_HVT U1116 ( .A1(n850), .A2(n863), .Y(n852) );
  NAND3X0_HVT U1117 ( .A1(n1150), .A2(n358), .A3(n856), .Y(n851) );
  NAND4X0_HVT U1118 ( .A1(n1132), .A2(n853), .A3(n852), .A4(n851), .Y(n855) );
  NAND4X0_HVT U1119 ( .A1(sram_raddr_b3[6]), .A2(sram_raddr_b3[5]), .A3(n1110), 
        .A4(n1305), .Y(n874) );
  AND2X1_HVT U1120 ( .A1(n169), .A2(n874), .Y(n866) );
  OA222X1_HVT U1121 ( .A1(sram_raddr_b3[6]), .A2(n223), .A3(sram_raddr_b3[6]), 
        .A4(sram_raddr_b3[5]), .A5(sram_raddr_b3[6]), .A6(n1110), .Y(n854) );
  AO22X1_HVT U1122 ( .A1(n204), .A2(n855), .A3(n866), .A4(n854), .Y(
        n_sram_raddr_b3[6]) );
  AND4X1_HVT U1123 ( .A1(n222), .A2(sram_raddr_b3[6]), .A3(sram_raddr_b3[5]), 
        .A4(n1110), .Y(n890) );
  NAND2X0_HVT U1124 ( .A1(sram_raddr_b3[6]), .A2(n856), .Y(n870) );
  NAND3X0_HVT U1125 ( .A1(n1150), .A2(n388), .A3(n870), .Y(n860) );
  NAND2X0_HVT U1126 ( .A1(n269), .A2(n857), .Y(n867) );
  AO221X1_HVT U1127 ( .A1(n867), .A2(n857), .A3(n867), .A4(n269), .A5(n218), 
        .Y(n1143) );
  AO221X1_HVT U1128 ( .A1(n212), .A2(n1389), .A3(n211), .A4(n870), .A5(n388), 
        .Y(n858) );
  NAND4X0_HVT U1129 ( .A1(n860), .A2(n859), .A3(n1143), .A4(n858), .Y(n864) );
  OA221X1_HVT U1130 ( .A1(n864), .A2(n863), .A3(n864), .A4(n862), .A5(n201), 
        .Y(n865) );
  AO221X1_HVT U1131 ( .A1(sram_raddr_b3[7]), .A2(n866), .A3(n388), .A4(n890), 
        .A5(n865), .Y(n_sram_raddr_b3[7]) );
  NAND2X0_HVT U1132 ( .A1(n868), .A2(n346), .Y(n880) );
  AO221X1_HVT U1133 ( .A1(n880), .A2(n868), .A3(n880), .A4(n346), .A5(n218), 
        .Y(n1156) );
  OA21X1_HVT U1134 ( .A1(n869), .A2(n886), .A3(n1156), .Y(n873) );
  NAND4X0_HVT U1135 ( .A1(n1150), .A2(n273), .A3(n388), .A4(n870), .Y(n883) );
  AND3X1_HVT U1136 ( .A1(n212), .A2(n388), .A3(n870), .Y(n879) );
  OR3X1_HVT U1137 ( .A1(n1160), .A2(n879), .A3(n273), .Y(n871) );
  NAND4X0_HVT U1138 ( .A1(n873), .A2(n872), .A3(n883), .A4(n871), .Y(n878) );
  OR3X1_HVT U1139 ( .A1(n388), .A2(n874), .A3(n273), .Y(n875) );
  NAND2X0_HVT U1140 ( .A1(n875), .A2(n169), .Y(n888) );
  AO21X1_HVT U1141 ( .A1(sram_raddr_b3[7]), .A2(n890), .A3(sram_raddr_b3[8]), 
        .Y(n876) );
  AO22X1_HVT U1142 ( .A1(n204), .A2(n878), .A3(n877), .A4(n876), .Y(
        n_sram_raddr_b3[8]) );
  AO21X1_HVT U1143 ( .A1(n879), .A2(n273), .A3(n1160), .Y(n882) );
  AO221X1_HVT U1144 ( .A1(sram_raddr_b0[9]), .A2(n881), .A3(n401), .A4(n880), 
        .A5(n217), .Y(n1170) );
  OA221X1_HVT U1145 ( .A1(sram_raddr_b3[9]), .A2(n883), .A3(n361), .A4(n882), 
        .A5(n1170), .Y(n887) );
  OA22X1_HVT U1146 ( .A1(n889), .A2(n226), .A3(n361), .A4(n888), .Y(n892) );
  NAND4X0_HVT U1147 ( .A1(sram_raddr_b3[7]), .A2(sram_raddr_b3[8]), .A3(n890), 
        .A4(n361), .Y(n891) );
  NAND2X0_HVT U1148 ( .A1(n892), .A2(n891), .Y(n_sram_raddr_b3[9]) );
  NAND2X0_HVT U1149 ( .A1(n1176), .A2(n173), .Y(n957) );
  AO22X1_HVT U1150 ( .A1(n190), .A2(n398), .A3(n1262), .A4(n243), .Y(n893) );
  AO221X1_HVT U1151 ( .A1(sram_raddr_b4[0]), .A2(n1238), .A3(n259), .A4(n957), 
        .A5(n893), .Y(n894) );
  AO22X1_HVT U1152 ( .A1(n205), .A2(n894), .A3(sram_raddr_b4[0]), .A4(n169), 
        .Y(n_sram_raddr_b4[0]) );
  OA22X1_HVT U1153 ( .A1(n895), .A2(n326), .A3(n970), .A4(n1181), .Y(n899) );
  NAND2X0_HVT U1154 ( .A1(n896), .A2(n901), .Y(n897) );
  NAND2X0_HVT U1155 ( .A1(n1262), .A2(n897), .Y(n1179) );
  NAND3X0_HVT U1156 ( .A1(n899), .A2(n898), .A3(n1179), .Y(n900) );
  AO22X1_HVT U1157 ( .A1(n205), .A2(n900), .A3(sram_raddr_b4[1]), .A4(n169), 
        .Y(n_sram_raddr_b4[1]) );
  AO21X1_HVT U1158 ( .A1(n204), .A2(n1308), .A3(n230), .Y(n1561) );
  AND2X1_HVT U1159 ( .A1(sram_raddr_b1[2]), .A2(n901), .Y(n908) );
  NAND2X0_HVT U1160 ( .A1(n1228), .A2(n314), .Y(n907) );
  NAND3X0_HVT U1161 ( .A1(n902), .A2(n1185), .A3(n907), .Y(n905) );
  OA221X1_HVT U1162 ( .A1(n905), .A2(n957), .A3(n905), .A4(n904), .A5(n203), 
        .Y(n906) );
  AO221X1_HVT U1163 ( .A1(sram_raddr_b4[2]), .A2(n1561), .A3(n314), .A4(n221), 
        .A5(n906), .Y(n_sram_raddr_b4[2]) );
  NAND3X0_HVT U1164 ( .A1(sram_raddr_b4[3]), .A2(sram_raddr_b4[2]), .A3(
        sram_raddr_b4[4]), .Y(n928) );
  NAND2X0_HVT U1165 ( .A1(sram_raddr_b4[3]), .A2(sram_raddr_b4[2]), .Y(n1202)
         );
  NAND2X0_HVT U1166 ( .A1(n357), .A2(n1202), .Y(n921) );
  AND2X1_HVT U1167 ( .A1(n928), .A2(n921), .Y(n918) );
  OA22X1_HVT U1168 ( .A1(n970), .A2(n911), .A3(n918), .A4(n1200), .Y(n917) );
  OA21X1_HVT U1169 ( .A1(n914), .A2(n912), .A3(n316), .Y(n920) );
  AO221X1_HVT U1170 ( .A1(n915), .A2(n914), .A3(n915), .A4(n913), .A5(n218), 
        .Y(n1208) );
  NAND3X0_HVT U1171 ( .A1(n917), .A2(n916), .A3(n1208), .Y(n919) );
  AO222X1_HVT U1172 ( .A1(n919), .A2(n1558), .A3(n1561), .A4(sram_raddr_b4[4]), 
        .A5(n918), .A6(n223), .Y(n_sram_raddr_b4[4]) );
  NAND3X0_HVT U1173 ( .A1(n276), .A2(n357), .A3(n1202), .Y(n940) );
  OR2X1_HVT U1174 ( .A1(n1200), .A2(n940), .Y(n923) );
  NAND2X0_HVT U1175 ( .A1(n920), .A2(n270), .Y(n929) );
  AO221X1_HVT U1176 ( .A1(n929), .A2(n920), .A3(n929), .A4(n270), .A5(n218), 
        .Y(n1213) );
  OAI221X1_HVT U1177 ( .A1(n1308), .A2(n254), .A3(n1308), .A4(n921), .A5(
        sram_raddr_b4[5]), .Y(n922) );
  NAND4X0_HVT U1178 ( .A1(n924), .A2(n923), .A3(n1213), .A4(n922), .Y(n927) );
  NAND2X0_HVT U1179 ( .A1(sram_raddr_b1[6]), .A2(n929), .Y(n938) );
  OR2X1_HVT U1180 ( .A1(n970), .A2(n930), .Y(n933) );
  AO221X1_HVT U1181 ( .A1(n213), .A2(n1200), .A3(n212), .A4(n940), .A5(n387), 
        .Y(n932) );
  NAND3X0_HVT U1182 ( .A1(n1228), .A2(n387), .A3(n940), .Y(n931) );
  NAND4X0_HVT U1183 ( .A1(n934), .A2(n933), .A3(n932), .A4(n931), .Y(n937) );
  NAND3X0_HVT U1184 ( .A1(sram_raddr_b4[6]), .A2(sram_raddr_b4[5]), .A3(n1204), 
        .Y(n944) );
  OA221X1_HVT U1185 ( .A1(sram_raddr_b4[6]), .A2(sram_raddr_b4[5]), .A3(
        sram_raddr_b4[6]), .A4(n1204), .A5(n944), .Y(n935) );
  AO22X1_HVT U1186 ( .A1(n222), .A2(n935), .A3(n232), .A4(sram_raddr_b4[6]), 
        .Y(n936) );
  AO221X1_HVT U1187 ( .A1(n205), .A2(n1226), .A3(n202), .A4(n937), .A5(n936), 
        .Y(n_sram_raddr_b4[6]) );
  NAND2X0_HVT U1188 ( .A1(n333), .A2(n938), .Y(n951) );
  AO221X1_HVT U1189 ( .A1(n951), .A2(n938), .A3(n951), .A4(n333), .A5(n218), 
        .Y(n1230) );
  OA21X1_HVT U1190 ( .A1(n970), .A2(n939), .A3(n1230), .Y(n943) );
  NAND2X0_HVT U1191 ( .A1(sram_raddr_b4[6]), .A2(n940), .Y(n962) );
  NAND3X0_HVT U1192 ( .A1(n1228), .A2(n332), .A3(n962), .Y(n953) );
  AO221X1_HVT U1193 ( .A1(n211), .A2(col[0]), .A3(n211), .A4(n962), .A5(n332), 
        .Y(n941) );
  NAND4X0_HVT U1194 ( .A1(n943), .A2(n953), .A3(n942), .A4(n941), .Y(n948) );
  NAND2X0_HVT U1195 ( .A1(n332), .A2(n944), .Y(n947) );
  NAND2X0_HVT U1196 ( .A1(sram_raddr_b4[7]), .A2(n950), .Y(n945) );
  NAND2X0_HVT U1197 ( .A1(n222), .A2(n945), .Y(n949) );
  AO222X1_HVT U1198 ( .A1(n948), .A2(n201), .A3(n947), .A4(n946), .A5(
        sram_raddr_b4[7]), .A6(n230), .Y(n_sram_raddr_b4[7]) );
  AND3X1_HVT U1199 ( .A1(n221), .A2(sram_raddr_b4[7]), .A3(n950), .Y(n961) );
  OR2X1_HVT U1200 ( .A1(n953), .A2(sram_raddr_b4[8]), .Y(n967) );
  NAND2X0_HVT U1201 ( .A1(n952), .A2(n272), .Y(n964) );
  AO221X1_HVT U1202 ( .A1(n964), .A2(n952), .A3(n964), .A4(n272), .A5(n218), 
        .Y(n1241) );
  NAND3X0_HVT U1203 ( .A1(n1238), .A2(n953), .A3(sram_raddr_b4[8]), .Y(n954)
         );
  NAND4X0_HVT U1204 ( .A1(n967), .A2(n955), .A3(n1241), .A4(n954), .Y(n958) );
  OA221X1_HVT U1205 ( .A1(n958), .A2(n957), .A3(n958), .A4(n956), .A5(n203), 
        .Y(n959) );
  AO221X1_HVT U1206 ( .A1(n960), .A2(sram_raddr_b4[8]), .A3(n960), .A4(n961), 
        .A5(n959), .Y(n_sram_raddr_b4[8]) );
  NAND3X0_HVT U1207 ( .A1(n351), .A2(n961), .A3(sram_raddr_b4[8]), .Y(n975) );
  AND2X1_HVT U1208 ( .A1(n332), .A2(n962), .Y(n963) );
  OA221X1_HVT U1209 ( .A1(n1200), .A2(n963), .A3(n1200), .A4(n345), .A5(n211), 
        .Y(n966) );
  OA221X1_HVT U1210 ( .A1(sram_raddr_b4[9]), .A2(n967), .A3(n351), .A4(n966), 
        .A5(n1245), .Y(n971) );
  OA22X1_HVT U1211 ( .A1(n973), .A2(n351), .A3(n972), .A4(n226), .Y(n974) );
  NAND2X0_HVT U1212 ( .A1(n975), .A2(n974), .Y(n_sram_raddr_b4[9]) );
  NAND2X0_HVT U1213 ( .A1(n225), .A2(n1328), .Y(n1019) );
  AO22X1_HVT U1214 ( .A1(n190), .A2(n399), .A3(n1262), .A4(n260), .Y(n976) );
  AO221X1_HVT U1215 ( .A1(sram_raddr_b5[0]), .A2(n1334), .A3(n244), .A4(n1019), 
        .A5(n976), .Y(n977) );
  AO22X1_HVT U1216 ( .A1(n202), .A2(n977), .A3(sram_raddr_b5[0]), .A4(n215), 
        .Y(n_sram_raddr_b5[0]) );
  OA22X1_HVT U1217 ( .A1(n978), .A2(n327), .A3(n1073), .A4(n1267), .Y(n982) );
  NAND2X0_HVT U1218 ( .A1(n979), .A2(n1001), .Y(n980) );
  NAND2X0_HVT U1219 ( .A1(n1262), .A2(n980), .Y(n1265) );
  NAND3X0_HVT U1220 ( .A1(n982), .A2(n981), .A3(n1265), .Y(n983) );
  AO22X1_HVT U1221 ( .A1(n205), .A2(n983), .A3(sram_raddr_b5[1]), .A4(n215), 
        .Y(n_sram_raddr_b5[1]) );
  AO22X1_HVT U1222 ( .A1(sram_raddr_b5[2]), .A2(n213), .A3(n313), .A4(n1301), 
        .Y(n985) );
  AO221X1_HVT U1223 ( .A1(sram_raddr_b2[2]), .A2(n1001), .A3(n354), .A4(n999), 
        .A5(n218), .Y(n1271) );
  NAND3X0_HVT U1224 ( .A1(n985), .A2(n984), .A3(n1271), .Y(n987) );
  OA221X1_HVT U1225 ( .A1(n987), .A2(n1019), .A3(n987), .A4(n986), .A5(n202), 
        .Y(n988) );
  AO221X1_HVT U1226 ( .A1(sram_raddr_b5[2]), .A2(n232), .A3(n313), .A4(n188), 
        .A5(n988), .Y(n_sram_raddr_b5[2]) );
  OA222X1_HVT U1227 ( .A1(sram_raddr_b2[3]), .A2(sram_raddr_b2[2]), .A3(
        sram_raddr_b2[3]), .A4(n1001), .A5(n999), .A6(n998), .Y(n989) );
  NAND2X0_HVT U1228 ( .A1(n1262), .A2(n989), .Y(n1282) );
  AO221X1_HVT U1229 ( .A1(n212), .A2(sram_raddr_b5[2]), .A3(n214), .A4(n1301), 
        .A5(n384), .Y(n991) );
  NAND3X0_HVT U1230 ( .A1(sram_raddr_b5[2]), .A2(n1320), .A3(n384), .Y(n990)
         );
  NAND2X0_HVT U1231 ( .A1(n222), .A2(n313), .Y(n994) );
  NAND2X0_HVT U1232 ( .A1(n1305), .A2(n994), .Y(n996) );
  AND2X1_HVT U1233 ( .A1(sram_raddr_b5[2]), .A2(n384), .Y(n995) );
  AO222X1_HVT U1234 ( .A1(n997), .A2(n203), .A3(n996), .A4(sram_raddr_b5[3]), 
        .A5(n995), .A6(n222), .Y(n_sram_raddr_b5[3]) );
  NAND3X0_HVT U1235 ( .A1(sram_raddr_b5[4]), .A2(sram_raddr_b5[3]), .A3(
        sram_raddr_b5[2]), .Y(n1015) );
  NAND2X0_HVT U1236 ( .A1(sram_raddr_b5[3]), .A2(sram_raddr_b5[2]), .Y(n1290)
         );
  NAND2X0_HVT U1237 ( .A1(n341), .A2(n1290), .Y(n1009) );
  AND2X1_HVT U1238 ( .A1(n1015), .A2(n1009), .Y(n1006) );
  OA22X1_HVT U1239 ( .A1(n211), .A2(n341), .A3(n1006), .A4(n1301), .Y(n1005)
         );
  OA21X1_HVT U1240 ( .A1(n999), .A2(n998), .A3(n255), .Y(n1008) );
  OAI221X1_HVT U1241 ( .A1(n1008), .A2(n1001), .A3(n1008), .A4(n1000), .A5(
        n1262), .Y(n1296) );
  OR2X1_HVT U1242 ( .A1(n1073), .A2(n1002), .Y(n1003) );
  NAND4X0_HVT U1243 ( .A1(n1005), .A2(n1004), .A3(n1296), .A4(n1003), .Y(n1007) );
  AO222X1_HVT U1244 ( .A1(n1007), .A2(n205), .A3(n231), .A4(sram_raddr_b5[4]), 
        .A5(n221), .A6(n1006), .Y(n_sram_raddr_b5[4]) );
  NAND2X0_HVT U1245 ( .A1(n1008), .A2(n334), .Y(n1035) );
  AO221X1_HVT U1246 ( .A1(n1035), .A2(n1008), .A3(n1035), .A4(n334), .A5(n217), 
        .Y(n1304) );
  NAND3X0_HVT U1247 ( .A1(n271), .A2(n341), .A3(n1290), .Y(n1026) );
  OAI221X1_HVT U1248 ( .A1(n1308), .A2(n312), .A3(n1308), .A4(n1009), .A5(
        sram_raddr_b5[5]), .Y(n1010) );
  OA22X1_HVT U1249 ( .A1(n1014), .A2(n219), .A3(n1305), .A4(n271), .Y(n1017)
         );
  AO221X1_HVT U1250 ( .A1(sram_raddr_b5[5]), .A2(n1292), .A3(n271), .A4(n1015), 
        .A5(n1368), .Y(n1016) );
  NAND2X0_HVT U1251 ( .A1(n1017), .A2(n1016), .Y(n_sram_raddr_b5[5]) );
  AO221X1_HVT U1252 ( .A1(sram_raddr_b2[6]), .A2(n1035), .A3(n337), .A4(n1018), 
        .A5(n218), .Y(n1309) );
  NAND2X0_HVT U1253 ( .A1(n1025), .A2(n1019), .Y(n1031) );
  NAND2X0_HVT U1254 ( .A1(sram_raddr_b5[6]), .A2(n1026), .Y(n1054) );
  NAND2X0_HVT U1255 ( .A1(n1320), .A2(n1054), .Y(n1029) );
  AO222X1_HVT U1256 ( .A1(n365), .A2(n1029), .A3(n365), .A4(n1028), .A5(n1029), 
        .A6(n213), .Y(n1030) );
  NAND4X0_HVT U1257 ( .A1(n1032), .A2(n1309), .A3(n1031), .A4(n1030), .Y(n1034) );
  NAND3X0_HVT U1258 ( .A1(sram_raddr_b5[6]), .A2(sram_raddr_b5[5]), .A3(n1292), 
        .Y(n1042) );
  AO21X1_HVT U1259 ( .A1(n221), .A2(n1042), .A3(n232), .Y(n1043) );
  OA222X1_HVT U1260 ( .A1(sram_raddr_b5[6]), .A2(n222), .A3(sram_raddr_b5[6]), 
        .A4(sram_raddr_b5[5]), .A5(sram_raddr_b5[6]), .A6(n1292), .Y(n1033) );
  AO22X1_HVT U1261 ( .A1(n1558), .A2(n1034), .A3(n1043), .A4(n1033), .Y(
        n_sram_raddr_b5[6]) );
  NAND2X0_HVT U1262 ( .A1(sram_raddr_b2[6]), .A2(n1035), .Y(n1036) );
  NAND2X0_HVT U1263 ( .A1(n267), .A2(n1036), .Y(n1046) );
  AO221X1_HVT U1264 ( .A1(n1046), .A2(n1036), .A3(n1046), .A4(n267), .A5(n218), 
        .Y(n1314) );
  OA21X1_HVT U1265 ( .A1(n1073), .A2(n1037), .A3(n1314), .Y(n1041) );
  NAND3X0_HVT U1266 ( .A1(n1320), .A2(n393), .A3(n1054), .Y(n1040) );
  AO221X1_HVT U1267 ( .A1(n214), .A2(col[1]), .A3(n212), .A4(n1054), .A5(n393), 
        .Y(n1038) );
  NAND4X0_HVT U1268 ( .A1(n1041), .A2(n1040), .A3(n1039), .A4(n1038), .Y(n1045) );
  OA222X1_HVT U1269 ( .A1(sram_raddr_b5[7]), .A2(n221), .A3(sram_raddr_b5[7]), 
        .A4(n1057), .A5(n1043), .A6(n393), .Y(n1044) );
  AO21X1_HVT U1270 ( .A1(n201), .A2(n1045), .A3(n1044), .Y(n_sram_raddr_b5[7])
         );
  OR2X1_HVT U1271 ( .A1(n1046), .A2(sram_raddr_b2[8]), .Y(n1066) );
  NAND2X0_HVT U1272 ( .A1(sram_raddr_b2[8]), .A2(n1046), .Y(n1048) );
  OA221X1_HVT U1273 ( .A1(n218), .A2(n1066), .A3(n218), .A4(n1048), .A5(n1047), 
        .Y(n1327) );
  AND3X1_HVT U1274 ( .A1(n212), .A2(n393), .A3(n1054), .Y(n1064) );
  NAND2X0_HVT U1275 ( .A1(sram_raddr_b5[8]), .A2(n1334), .Y(n1050) );
  OA22X1_HVT U1276 ( .A1(n1064), .A2(n1050), .A3(n1049), .A4(n1073), .Y(n1055)
         );
  NAND4X0_HVT U1277 ( .A1(n1320), .A2(n286), .A3(n393), .A4(n1054), .Y(n1069)
         );
  NAND3X0_HVT U1278 ( .A1(n1327), .A2(n1055), .A3(n1069), .Y(n1060) );
  NAND4X0_HVT U1279 ( .A1(sram_raddr_b5[8]), .A2(sram_raddr_b5[7]), .A3(n1057), 
        .A4(n1305), .Y(n1056) );
  NAND2X0_HVT U1280 ( .A1(n169), .A2(n1056), .Y(n1075) );
  AND3X1_HVT U1281 ( .A1(n221), .A2(sram_raddr_b5[7]), .A3(n1057), .Y(n1077)
         );
  OR2X1_HVT U1282 ( .A1(sram_raddr_b5[8]), .A2(n1077), .Y(n1058) );
  AO22X1_HVT U1283 ( .A1(n204), .A2(n1060), .A3(n1059), .A4(n1058), .Y(
        n_sram_raddr_b5[8]) );
  AO22X1_HVT U1284 ( .A1(col[1]), .A2(n211), .A3(n1064), .A4(n286), .Y(n1068)
         );
  OA221X1_HVT U1285 ( .A1(sram_raddr_b5[9]), .A2(n1069), .A3(n348), .A4(n1068), 
        .A5(n1333), .Y(n1074) );
  OA22X1_HVT U1286 ( .A1(n1076), .A2(n219), .A3(n348), .A4(n1075), .Y(n1079)
         );
  NAND3X0_HVT U1287 ( .A1(sram_raddr_b5[8]), .A2(n1077), .A3(n348), .Y(n1078)
         );
  NAND2X0_HVT U1288 ( .A1(n1079), .A2(n1078), .Y(n_sram_raddr_b5[9]) );
  AO22X1_HVT U1289 ( .A1(n1262), .A2(n242), .A3(n1322), .A4(n258), .Y(n1081)
         );
  AO221X1_HVT U1290 ( .A1(sram_raddr_b6[0]), .A2(n1086), .A3(n397), .A4(n1164), 
        .A5(n1081), .Y(n1082) );
  AO22X1_HVT U1291 ( .A1(n203), .A2(n1082), .A3(sram_raddr_b6[0]), .A4(n169), 
        .Y(n_sram_raddr_b6[0]) );
  AO22X1_HVT U1292 ( .A1(n1558), .A2(n1087), .A3(sram_raddr_b6[1]), .A4(n215), 
        .Y(n_sram_raddr_b6[1]) );
  AO22X1_HVT U1293 ( .A1(sram_raddr_b6[2]), .A2(n214), .A3(n239), .A4(n1127), 
        .Y(n1090) );
  AO221X1_HVT U1294 ( .A1(sram_raddr_b3[2]), .A2(n1111), .A3(n315), .A4(n1109), 
        .A5(n173), .Y(n1089) );
  NAND3X0_HVT U1295 ( .A1(n1090), .A2(n1089), .A3(n1088), .Y(n1093) );
  OA221X1_HVT U1296 ( .A1(n1093), .A2(n1164), .A3(n1093), .A4(n1092), .A5(n202), .Y(n1094) );
  AO221X1_HVT U1297 ( .A1(sram_raddr_b6[2]), .A2(n231), .A3(n239), .A4(n222), 
        .A5(n1094), .Y(n_sram_raddr_b6[2]) );
  NAND2X0_HVT U1298 ( .A1(n223), .A2(n239), .Y(n1095) );
  NAND2X0_HVT U1299 ( .A1(n1305), .A2(n1095), .Y(n1106) );
  NAND2X0_HVT U1300 ( .A1(n239), .A2(n1150), .Y(n1096) );
  NAND2X0_HVT U1301 ( .A1(n211), .A2(n1096), .Y(n1098) );
  AOI22X1_HVT U1302 ( .A1(sram_raddr_b6[3]), .A2(n1098), .A3(n1097), .A4(n1164), .Y(n1103) );
  NAND3X0_HVT U1303 ( .A1(sram_raddr_b6[2]), .A2(n389), .A3(n1150), .Y(n1101)
         );
  OA222X1_HVT U1304 ( .A1(sram_raddr_b3[3]), .A2(sram_raddr_b3[2]), .A3(
        sram_raddr_b3[3]), .A4(n1111), .A5(n1109), .A6(n1108), .Y(n1099) );
  NAND2X0_HVT U1305 ( .A1(n1322), .A2(n1099), .Y(n1100) );
  NAND4X0_HVT U1306 ( .A1(n1103), .A2(n1102), .A3(n1101), .A4(n1100), .Y(n1105) );
  AND2X1_HVT U1307 ( .A1(sram_raddr_b6[2]), .A2(n389), .Y(n1104) );
  AO222X1_HVT U1308 ( .A1(n1106), .A2(sram_raddr_b6[3]), .A3(n1105), .A4(n1558), .A5(n1104), .A6(n221), .Y(n_sram_raddr_b6[3]) );
  AND3X1_HVT U1309 ( .A1(sram_raddr_b6[3]), .A2(sram_raddr_b6[2]), .A3(
        sram_raddr_b6[4]), .Y(n1125) );
  OA21X1_HVT U1310 ( .A1(n239), .A2(n389), .A3(n280), .Y(n1126) );
  NOR2X0_HVT U1311 ( .A1(n1125), .A2(n1126), .Y(n1116) );
  OA22X1_HVT U1312 ( .A1(n1127), .A2(n1116), .A3(n214), .A4(n280), .Y(n1115)
         );
  NAND2X0_HVT U1313 ( .A1(n1164), .A2(n1107), .Y(n1113) );
  OA21X1_HVT U1314 ( .A1(n1109), .A2(n1108), .A3(n335), .Y(n1118) );
  OAI221X1_HVT U1315 ( .A1(n1118), .A2(n1111), .A3(n1118), .A4(n1110), .A5(
        n178), .Y(n1112) );
  NAND4X0_HVT U1316 ( .A1(n1115), .A2(n1114), .A3(n1113), .A4(n1112), .Y(n1117) );
  AO222X1_HVT U1317 ( .A1(n1117), .A2(n202), .A3(n232), .A4(sram_raddr_b6[4]), 
        .A5(n179), .A6(n1116), .Y(n_sram_raddr_b6[4]) );
  NAND3X0_HVT U1318 ( .A1(n1126), .A2(n363), .A3(n1150), .Y(n1122) );
  AO221X1_HVT U1319 ( .A1(n214), .A2(n1127), .A3(n214), .A4(n1126), .A5(n363), 
        .Y(n1120) );
  NAND2X0_HVT U1320 ( .A1(n1118), .A2(n268), .Y(n1139) );
  AO221X1_HVT U1321 ( .A1(n1139), .A2(n1118), .A3(n1139), .A4(n268), .A5(n224), 
        .Y(n1119) );
  NAND4X0_HVT U1322 ( .A1(n1122), .A2(n1121), .A3(n1120), .A4(n1119), .Y(n1124) );
  NAND4X0_HVT U1323 ( .A1(sram_raddr_b6[3]), .A2(sram_raddr_b6[2]), .A3(
        sram_raddr_b6[5]), .A4(sram_raddr_b6[4]), .Y(n1136) );
  NAND2X0_HVT U1324 ( .A1(n1126), .A2(n363), .Y(n1138) );
  AO221X1_HVT U1325 ( .A1(n213), .A2(n1127), .A3(n213), .A4(n1138), .A5(n408), 
        .Y(n1131) );
  AO221X1_HVT U1326 ( .A1(sram_raddr_b3[6]), .A2(n1139), .A3(n358), .A4(n1128), 
        .A5(n225), .Y(n1130) );
  NAND3X0_HVT U1327 ( .A1(n408), .A2(n1150), .A3(n1138), .Y(n1129) );
  NAND4X0_HVT U1328 ( .A1(n1132), .A2(n1131), .A3(n1130), .A4(n1129), .Y(n1135) );
  NAND2X0_HVT U1329 ( .A1(sram_raddr_b6[6]), .A2(n1137), .Y(n1147) );
  NAND2X0_HVT U1330 ( .A1(sram_raddr_b6[6]), .A2(n1138), .Y(n1153) );
  NAND3X0_HVT U1331 ( .A1(n338), .A2(n1150), .A3(n1153), .Y(n1144) );
  NAND2X0_HVT U1332 ( .A1(sram_raddr_b3[6]), .A2(n1139), .Y(n1140) );
  NAND2X0_HVT U1333 ( .A1(n388), .A2(n1140), .Y(n1151) );
  AO221X1_HVT U1334 ( .A1(n1151), .A2(n1140), .A3(n1151), .A4(n388), .A5(n173), 
        .Y(n1142) );
  AO221X1_HVT U1335 ( .A1(n214), .A2(n1389), .A3(n214), .A4(n1153), .A5(n338), 
        .Y(n1141) );
  NAND4X0_HVT U1336 ( .A1(n1144), .A2(n1143), .A3(n1142), .A4(n1141), .Y(n1146) );
  NAND2X0_HVT U1337 ( .A1(sram_raddr_b6[7]), .A2(n1149), .Y(n1148) );
  AO221X1_HVT U1338 ( .A1(n188), .A2(n274), .A3(n221), .A4(n1148), .A5(n232), 
        .Y(n1172) );
  AND3X1_HVT U1339 ( .A1(n221), .A2(sram_raddr_b6[7]), .A3(n1149), .Y(n1173)
         );
  NAND4X0_HVT U1340 ( .A1(n274), .A2(n338), .A3(n1150), .A4(n1153), .Y(n1162)
         );
  NAND2X0_HVT U1341 ( .A1(n1152), .A2(n273), .Y(n1166) );
  AO221X1_HVT U1342 ( .A1(n1166), .A2(n1152), .A3(n1166), .A4(n273), .A5(n173), 
        .Y(n1155) );
  AND3X1_HVT U1343 ( .A1(n213), .A2(n338), .A3(n1153), .Y(n1161) );
  OR3X1_HVT U1344 ( .A1(n1160), .A2(n1161), .A3(n274), .Y(n1154) );
  NAND4X0_HVT U1345 ( .A1(n1162), .A2(n1156), .A3(n1155), .A4(n1154), .Y(n1158) );
  OA221X1_HVT U1346 ( .A1(n1158), .A2(n1157), .A3(n1158), .A4(n1164), .A5(n202), .Y(n1159) );
  AO221X1_HVT U1347 ( .A1(n1172), .A2(sram_raddr_b6[8]), .A3(n1172), .A4(n1173), .A5(n1159), .Y(n_sram_raddr_b6[8]) );
  AO21X1_HVT U1348 ( .A1(n1161), .A2(n274), .A3(n1160), .Y(n1163) );
  AO22X1_HVT U1349 ( .A1(sram_raddr_b6[9]), .A2(n1163), .A3(n373), .A4(n1162), 
        .Y(n1171) );
  NAND2X0_HVT U1350 ( .A1(n1165), .A2(n1164), .Y(n1169) );
  AO221X1_HVT U1351 ( .A1(sram_raddr_b3[9]), .A2(n1167), .A3(n361), .A4(n1166), 
        .A5(n225), .Y(n1168) );
  NAND4X0_HVT U1352 ( .A1(n1171), .A2(n1170), .A3(n1169), .A4(n1168), .Y(n1175) );
  OA222X1_HVT U1353 ( .A1(sram_raddr_b6[9]), .A2(sram_raddr_b6[8]), .A3(
        sram_raddr_b6[9]), .A4(n1173), .A5(n373), .A6(n1172), .Y(n1174) );
  AO21X1_HVT U1354 ( .A1(n205), .A2(n1175), .A3(n1174), .Y(n_sram_raddr_b6[9])
         );
  AO22X1_HVT U1355 ( .A1(n1262), .A2(n243), .A3(n178), .A4(n259), .Y(n1177) );
  AO221X1_HVT U1356 ( .A1(sram_raddr_b7[0]), .A2(n1238), .A3(n398), .A4(n1250), 
        .A5(n1177), .Y(n1178) );
  AO22X1_HVT U1357 ( .A1(n204), .A2(n1178), .A3(sram_raddr_b7[0]), .A4(n169), 
        .Y(n_sram_raddr_b7[0]) );
  AO22X1_HVT U1358 ( .A1(n204), .A2(n1182), .A3(sram_raddr_b7[1]), .A4(n215), 
        .Y(n_sram_raddr_b7[1]) );
  NAND2X0_HVT U1359 ( .A1(n1228), .A2(n240), .Y(n1189) );
  OA21X1_HVT U1360 ( .A1(n212), .A2(n240), .A3(n1189), .Y(n1184) );
  AO221X1_HVT U1361 ( .A1(sram_raddr_b4[2]), .A2(n1205), .A3(n314), .A4(n1203), 
        .A5(n173), .Y(n1183) );
  NAND3X0_HVT U1362 ( .A1(n1185), .A2(n1184), .A3(n1183), .Y(n1187) );
  OA221X1_HVT U1363 ( .A1(n1187), .A2(n1250), .A3(n1187), .A4(n1186), .A5(n203), .Y(n1188) );
  AO221X1_HVT U1364 ( .A1(sram_raddr_b7[2]), .A2(n232), .A3(n240), .A4(n223), 
        .A5(n1188), .Y(n_sram_raddr_b7[2]) );
  NAND2X0_HVT U1365 ( .A1(n214), .A2(n1189), .Y(n1190) );
  OA222X1_HVT U1366 ( .A1(sram_raddr_b7[3]), .A2(n1228), .A3(sram_raddr_b7[3]), 
        .A4(sram_raddr_b7[2]), .A5(n382), .A6(n1190), .Y(n1194) );
  OA222X1_HVT U1367 ( .A1(sram_raddr_b4[3]), .A2(sram_raddr_b4[2]), .A3(
        sram_raddr_b4[3]), .A4(n1205), .A5(n1203), .A6(n1202), .Y(n1192) );
  AO22X1_HVT U1368 ( .A1(n178), .A2(n1192), .A3(n1191), .A4(n1250), .Y(n1193)
         );
  OR3X1_HVT U1369 ( .A1(n1195), .A2(n1194), .A3(n1193), .Y(n1199) );
  NAND2X0_HVT U1370 ( .A1(n221), .A2(n240), .Y(n1196) );
  NAND2X0_HVT U1371 ( .A1(n1305), .A2(n1196), .Y(n1198) );
  AND2X1_HVT U1372 ( .A1(sram_raddr_b7[2]), .A2(n382), .Y(n1197) );
  AO222X1_HVT U1373 ( .A1(n1199), .A2(n201), .A3(n1198), .A4(sram_raddr_b7[3]), 
        .A5(n1197), .A6(n221), .Y(n_sram_raddr_b7[3]) );
  AND3X1_HVT U1374 ( .A1(sram_raddr_b7[3]), .A2(sram_raddr_b7[2]), .A3(
        sram_raddr_b7[4]), .Y(n1215) );
  OA21X1_HVT U1375 ( .A1(n240), .A2(n382), .A3(n281), .Y(n1217) );
  NOR2X0_HVT U1376 ( .A1(n1215), .A2(n1217), .Y(n1210) );
  OA22X1_HVT U1377 ( .A1(n213), .A2(n281), .A3(n1210), .A4(n1200), .Y(n1209)
         );
  NAND2X0_HVT U1378 ( .A1(n1250), .A2(n1201), .Y(n1207) );
  OA21X1_HVT U1379 ( .A1(n1203), .A2(n1202), .A3(n357), .Y(n1212) );
  OAI221X1_HVT U1380 ( .A1(n1212), .A2(n1205), .A3(n1212), .A4(n1204), .A5(
        n178), .Y(n1206) );
  NAND4X0_HVT U1381 ( .A1(n1209), .A2(n1208), .A3(n1207), .A4(n1206), .Y(n1211) );
  AO222X1_HVT U1382 ( .A1(n1211), .A2(n202), .A3(n232), .A4(sram_raddr_b7[4]), 
        .A5(n179), .A6(n1210), .Y(n_sram_raddr_b7[4]) );
  NAND2X0_HVT U1383 ( .A1(n1212), .A2(n276), .Y(n1216) );
  NAND4X0_HVT U1384 ( .A1(sram_raddr_b7[3]), .A2(sram_raddr_b7[2]), .A3(
        sram_raddr_b7[5]), .A4(sram_raddr_b7[4]), .Y(n1221) );
  NAND2X0_HVT U1385 ( .A1(sram_raddr_b4[6]), .A2(n1216), .Y(n1229) );
  NAND2X0_HVT U1386 ( .A1(n1217), .A2(n364), .Y(n1227) );
  HADDX1_HVT U1387 ( .A0(sram_raddr_b7[6]), .B0(n1227), .SO(n1218) );
  NAND2X0_HVT U1388 ( .A1(sram_raddr_b7[6]), .A2(n1222), .Y(n1232) );
  OA21X1_HVT U1389 ( .A1(sram_raddr_b7[6]), .A2(n1222), .A3(n1232), .Y(n1223)
         );
  AO22X1_HVT U1390 ( .A1(n188), .A2(n1223), .A3(n230), .A4(sram_raddr_b7[6]), 
        .Y(n1224) );
  AO221X1_HVT U1391 ( .A1(n204), .A2(n1226), .A3(n1558), .A4(n1225), .A5(n1224), .Y(n_sram_raddr_b7[6]) );
  NAND2X0_HVT U1392 ( .A1(sram_raddr_b7[6]), .A2(n1227), .Y(n1246) );
  NAND3X0_HVT U1393 ( .A1(n1228), .A2(n347), .A3(n1246), .Y(n1237) );
  NAND2X0_HVT U1394 ( .A1(n332), .A2(n1229), .Y(n1235) );
  NAND2X0_HVT U1395 ( .A1(sram_raddr_b7[7]), .A2(n1234), .Y(n1233) );
  AO221X1_HVT U1396 ( .A1(n222), .A2(n391), .A3(n188), .A4(n1233), .A5(n232), 
        .Y(n1256) );
  AND3X1_HVT U1397 ( .A1(n188), .A2(sram_raddr_b7[7]), .A3(n1234), .Y(n1257)
         );
  OR2X1_HVT U1398 ( .A1(n1237), .A2(sram_raddr_b7[8]), .Y(n1248) );
  NAND2X0_HVT U1399 ( .A1(n1236), .A2(n345), .Y(n1249) );
  AO221X1_HVT U1400 ( .A1(n1249), .A2(n1236), .A3(n1249), .A4(n345), .A5(n173), 
        .Y(n1240) );
  NAND3X0_HVT U1401 ( .A1(n1238), .A2(n1237), .A3(sram_raddr_b7[8]), .Y(n1239)
         );
  NAND4X0_HVT U1402 ( .A1(n1248), .A2(n1241), .A3(n1240), .A4(n1239), .Y(n1243) );
  OA221X1_HVT U1403 ( .A1(n1243), .A2(n1250), .A3(n1243), .A4(n1242), .A5(n203), .Y(n1244) );
  AO221X1_HVT U1404 ( .A1(n1256), .A2(sram_raddr_b7[8]), .A3(n1256), .A4(n1257), .A5(n1244), .Y(n_sram_raddr_b7[8]) );
  NAND2X0_HVT U1405 ( .A1(n347), .A2(n1246), .Y(n1247) );
  AO221X1_HVT U1406 ( .A1(n254), .A2(sram_raddr_b7[8]), .A3(n254), .A4(n1247), 
        .A5(n1308), .Y(n1255) );
  HADDX1_HVT U1407 ( .A0(n351), .B0(n1249), .SO(n1252) );
  AO22X1_HVT U1408 ( .A1(n178), .A2(n1252), .A3(n1251), .A4(n1250), .Y(n1253)
         );
  AO221X1_HVT U1409 ( .A1(sram_raddr_b7[9]), .A2(n1255), .A3(n372), .A4(n1254), 
        .A5(n1253), .Y(n1259) );
  OA222X1_HVT U1410 ( .A1(sram_raddr_b7[9]), .A2(sram_raddr_b7[8]), .A3(
        sram_raddr_b7[9]), .A4(n1257), .A5(n372), .A6(n1256), .Y(n1258) );
  AO221X1_HVT U1411 ( .A1(n202), .A2(n1260), .A3(n205), .A4(n1259), .A5(n1258), 
        .Y(n_sram_raddr_b7[9]) );
  AO22X1_HVT U1412 ( .A1(n1262), .A2(n260), .A3(n178), .A4(n244), .Y(n1263) );
  AO221X1_HVT U1413 ( .A1(sram_raddr_b8[0]), .A2(n1334), .A3(n399), .A4(n1338), 
        .A5(n1263), .Y(n1264) );
  AO22X1_HVT U1414 ( .A1(n202), .A2(n1264), .A3(sram_raddr_b8[0]), .A4(n169), 
        .Y(n_sram_raddr_b8[0]) );
  AO22X1_HVT U1415 ( .A1(n205), .A2(n1269), .A3(sram_raddr_b8[1]), .A4(n215), 
        .Y(n_sram_raddr_b8[1]) );
  AO22X1_HVT U1416 ( .A1(sram_raddr_b8[2]), .A2(n214), .A3(n241), .A4(n1301), 
        .Y(n1272) );
  AO221X1_HVT U1417 ( .A1(sram_raddr_b5[2]), .A2(n1293), .A3(n313), .A4(n1291), 
        .A5(n225), .Y(n1270) );
  NAND3X0_HVT U1418 ( .A1(n1272), .A2(n1271), .A3(n1270), .Y(n1274) );
  OA221X1_HVT U1419 ( .A1(n1274), .A2(n1338), .A3(n1274), .A4(n1273), .A5(n202), .Y(n1275) );
  AO221X1_HVT U1420 ( .A1(sram_raddr_b8[2]), .A2(n232), .A3(n241), .A4(n223), 
        .A5(n1275), .Y(n_sram_raddr_b8[2]) );
  OA222X1_HVT U1421 ( .A1(sram_raddr_b5[3]), .A2(sram_raddr_b5[2]), .A3(
        sram_raddr_b5[3]), .A4(n1293), .A5(n1291), .A6(n1290), .Y(n1279) );
  OA21X1_HVT U1422 ( .A1(sram_raddr_b8[3]), .A2(n1277), .A3(n1276), .Y(n1278)
         );
  AOI22X1_HVT U1423 ( .A1(n178), .A2(n1279), .A3(n1278), .A4(n1338), .Y(n1283)
         );
  AO221X1_HVT U1424 ( .A1(n214), .A2(sram_raddr_b8[2]), .A3(n214), .A4(n1301), 
        .A5(n287), .Y(n1281) );
  NAND3X0_HVT U1425 ( .A1(sram_raddr_b8[2]), .A2(n1320), .A3(n287), .Y(n1280)
         );
  NAND4X0_HVT U1426 ( .A1(n1283), .A2(n1282), .A3(n1281), .A4(n1280), .Y(n1287) );
  NAND2X0_HVT U1427 ( .A1(n221), .A2(n241), .Y(n1284) );
  NAND2X0_HVT U1428 ( .A1(n1305), .A2(n1284), .Y(n1286) );
  AND2X1_HVT U1429 ( .A1(sram_raddr_b8[2]), .A2(n287), .Y(n1285) );
  AO222X1_HVT U1430 ( .A1(n1287), .A2(n201), .A3(n1286), .A4(sram_raddr_b8[3]), 
        .A5(n1285), .A6(n179), .Y(n_sram_raddr_b8[3]) );
  NAND3X0_HVT U1431 ( .A1(sram_raddr_b8[4]), .A2(sram_raddr_b8[3]), .A3(
        sram_raddr_b8[2]), .Y(n1306) );
  OA21X1_HVT U1432 ( .A1(n287), .A2(n241), .A3(n381), .Y(n1300) );
  AND2X1_HVT U1433 ( .A1(n1306), .A2(n1288), .Y(n1298) );
  OA22X1_HVT U1434 ( .A1(n213), .A2(n381), .A3(n1298), .A4(n1301), .Y(n1297)
         );
  NAND2X0_HVT U1435 ( .A1(n1338), .A2(n1289), .Y(n1295) );
  OA21X1_HVT U1436 ( .A1(n1291), .A2(n1290), .A3(n341), .Y(n1303) );
  OAI221X1_HVT U1437 ( .A1(n1303), .A2(n1293), .A3(n1303), .A4(n1292), .A5(
        n178), .Y(n1294) );
  NAND4X0_HVT U1438 ( .A1(n1297), .A2(n1296), .A3(n1295), .A4(n1294), .Y(n1299) );
  AO222X1_HVT U1439 ( .A1(n1299), .A2(n203), .A3(n230), .A4(sram_raddr_b8[4]), 
        .A5(n222), .A6(n1298), .Y(n_sram_raddr_b8[4]) );
  NAND2X0_HVT U1440 ( .A1(n1300), .A2(n342), .Y(n1307) );
  NAND2X0_HVT U1441 ( .A1(n1303), .A2(n271), .Y(n1312) );
  AND4X1_HVT U1442 ( .A1(sram_raddr_b8[5]), .A2(sram_raddr_b8[4]), .A3(
        sram_raddr_b8[3]), .A4(sram_raddr_b8[2]), .Y(n1311) );
  NAND2X0_HVT U1443 ( .A1(sram_raddr_b8[6]), .A2(n1307), .Y(n1324) );
  NAND2X0_HVT U1444 ( .A1(sram_raddr_b8[6]), .A2(n1311), .Y(n1316) );
  NAND2X0_HVT U1445 ( .A1(sram_raddr_b5[6]), .A2(n1312), .Y(n1313) );
  NAND2X0_HVT U1446 ( .A1(n393), .A2(n1313), .Y(n1321) );
  NAND2X0_HVT U1447 ( .A1(sram_raddr_b8[7]), .A2(n1319), .Y(n1318) );
  AO221X1_HVT U1448 ( .A1(n188), .A2(n359), .A3(n222), .A4(n1318), .A5(n230), 
        .Y(n1344) );
  AND3X1_HVT U1449 ( .A1(n188), .A2(sram_raddr_b8[7]), .A3(n1319), .Y(n1345)
         );
  NAND4X0_HVT U1450 ( .A1(n1320), .A2(n359), .A3(n275), .A4(n1324), .Y(n1336)
         );
  NAND2X0_HVT U1451 ( .A1(n1323), .A2(n286), .Y(n1337) );
  AO221X1_HVT U1452 ( .A1(n1337), .A2(n1323), .A3(n1337), .A4(n286), .A5(n225), 
        .Y(n1326) );
  NAND3X0_HVT U1453 ( .A1(n213), .A2(n275), .A3(n1324), .Y(n1335) );
  NAND3X0_HVT U1454 ( .A1(sram_raddr_b8[8]), .A2(n1334), .A3(n1335), .Y(n1325)
         );
  NAND4X0_HVT U1455 ( .A1(n1327), .A2(n1336), .A3(n1326), .A4(n1325), .Y(n1331) );
  OA221X1_HVT U1456 ( .A1(n1331), .A2(n1330), .A3(n1331), .A4(n1329), .A5(n202), .Y(n1332) );
  AO221X1_HVT U1457 ( .A1(n1344), .A2(sram_raddr_b8[8]), .A3(n1344), .A4(n1345), .A5(n1332), .Y(n_sram_raddr_b8[8]) );
  OA21X1_HVT U1458 ( .A1(sram_raddr_b8[8]), .A2(n1335), .A3(n1334), .Y(n1343)
         );
  HADDX1_HVT U1459 ( .A0(n348), .B0(n1337), .SO(n1340) );
  AO22X1_HVT U1460 ( .A1(n178), .A2(n1340), .A3(n1339), .A4(n1338), .Y(n1341)
         );
  AO221X1_HVT U1461 ( .A1(sram_raddr_b8[9]), .A2(n1343), .A3(n374), .A4(n1342), 
        .A5(n1341), .Y(n1347) );
  OA222X1_HVT U1462 ( .A1(sram_raddr_b8[9]), .A2(sram_raddr_b8[8]), .A3(
        sram_raddr_b8[9]), .A4(n1345), .A5(n374), .A6(n1344), .Y(n1346) );
  AO221X1_HVT U1463 ( .A1(n1558), .A2(n1348), .A3(n1558), .A4(n1347), .A5(
        n1346), .Y(n_sram_raddr_b8[9]) );
  OA221X1_HVT U1464 ( .A1(n1063), .A2(write_col_conv1[1]), .A3(n261), .A4(n320), .A5(n1062), .Y(n1352) );
  NAND2X0_HVT U1465 ( .A1(n1352), .A2(n1349), .Y(n_sram_write_enable_b0) );
  OA221X1_HVT U1466 ( .A1(write_col_conv1[1]), .A2(n262), .A3(n320), .A4(n1062), .A5(n1063), .Y(n1353) );
  NAND2X0_HVT U1467 ( .A1(n1353), .A2(n1349), .Y(n_sram_write_enable_b1) );
  NAND3X0_HVT U1468 ( .A1(write_col_conv1[1]), .A2(n1063), .A3(n262), .Y(n1472) );
  NAND3X0_HVT U1469 ( .A1(n1062), .A2(n261), .A3(n320), .Y(n1476) );
  NAND2X0_HVT U1470 ( .A1(n1472), .A2(n1476), .Y(n1469) );
  NAND2X0_HVT U1471 ( .A1(n1349), .A2(n1469), .Y(n_sram_write_enable_b2) );
  AO222X1_HVT U1472 ( .A1(write_row_conv1[3]), .A2(n1061), .A3(
        write_row_conv1[3]), .A4(write_row_conv1[2]), .A5(n249), .A6(n405), 
        .Y(n1350) );
  AND3X1_HVT U1473 ( .A1(n1350), .A2(n1470), .A3(n296), .Y(n1351) );
  NAND2X0_HVT U1474 ( .A1(n1352), .A2(n1351), .Y(n_sram_write_enable_b3) );
  NAND2X0_HVT U1475 ( .A1(n1353), .A2(n1351), .Y(n_sram_write_enable_b4) );
  NAND2X0_HVT U1476 ( .A1(n1351), .A2(n1469), .Y(n_sram_write_enable_b5) );
  OA222X1_HVT U1477 ( .A1(n1061), .A2(write_row_conv1[3]), .A3(n249), .A4(
        write_row_conv1[2]), .A5(n405), .A6(n296), .Y(n1473) );
  NAND4X0_HVT U1478 ( .A1(n1473), .A2(n1365), .A3(delay2_write_enable), .A4(
        n1352), .Y(n_sram_write_enable_b6) );
  NAND4X0_HVT U1479 ( .A1(n1473), .A2(n1365), .A3(delay2_write_enable), .A4(
        n1353), .Y(n_sram_write_enable_b7) );
  NAND4X0_HVT U1480 ( .A1(n1473), .A2(n1365), .A3(delay2_write_enable), .A4(
        n1469), .Y(n_sram_write_enable_b8) );
  AND3X1_HVT U1481 ( .A1(n1356), .A2(delay3_write_enable), .A3(n460), .Y(n1355) );
  NAND4X0_HVT U1482 ( .A1(n1355), .A2(n1513), .A3(n318), .A4(n257), .Y(
        n_sram_write_enable_c0) );
  AND3X1_HVT U1483 ( .A1(delay3_addr_change[2]), .A2(n1355), .A3(n318), .Y(
        n1354) );
  NAND2X0_HVT U1484 ( .A1(n1354), .A2(n1513), .Y(n_sram_write_enable_c1) );
  NAND4X0_HVT U1485 ( .A1(delay3_addr_change[3]), .A2(n1355), .A3(n1513), .A4(
        n257), .Y(n_sram_write_enable_c2) );
  NAND4X0_HVT U1486 ( .A1(delay3_addr_change[3]), .A2(delay3_addr_change[2]), 
        .A3(n1355), .A4(n1513), .Y(n_sram_write_enable_c3) );
  AND3X1_HVT U1487 ( .A1(delay3_addr_change[4]), .A2(n318), .A3(n257), .Y(
        n1509) );
  NAND4X0_HVT U1488 ( .A1(n1356), .A2(delay3_write_enable), .A3(n1509), .A4(
        n1513), .Y(n_sram_write_enable_c4) );
  NAND4X0_HVT U1489 ( .A1(mem_sel), .A2(n1355), .A3(n257), .A4(n318), .Y(
        n_sram_write_enable_d0) );
  NAND2X0_HVT U1490 ( .A1(mem_sel), .A2(n1354), .Y(n_sram_write_enable_d1) );
  NAND4X0_HVT U1491 ( .A1(delay3_addr_change[3]), .A2(mem_sel), .A3(n1355), 
        .A4(n257), .Y(n_sram_write_enable_d2) );
  NAND4X0_HVT U1492 ( .A1(mem_sel), .A2(delay3_addr_change[3]), .A3(
        delay3_addr_change[2]), .A4(n1355), .Y(n_sram_write_enable_d3) );
  NAND4X0_HVT U1493 ( .A1(mem_sel), .A2(n1356), .A3(delay3_write_enable), .A4(
        n1509), .Y(n_sram_write_enable_d4) );
  NAND4X0_HVT U1494 ( .A1(state[0]), .A2(n1023), .A3(n1024), .A4(n251), .Y(
        n1564) );
  NAND3X0_HVT U1495 ( .A1(n1023), .A2(n1446), .A3(state[2]), .Y(n1358) );
  NAND3X0_HVT U1496 ( .A1(state[1]), .A2(n1024), .A3(state[3]), .Y(n1447) );
  NAND2X0_HVT U1497 ( .A1(n1550), .A2(conv_done), .Y(n1367) );
  NAND3X0_HVT U1498 ( .A1(n1023), .A2(n1024), .A3(n310), .Y(n1360) );
  OA22X1_HVT U1499 ( .A1(conv_done), .A2(n1363), .A3(n1360), .A4(n1359), .Y(
        n1362) );
  NAND2X0_HVT U1500 ( .A1(n1446), .A2(state[2]), .Y(n1417) );
  NAND2X0_HVT U1501 ( .A1(n2004), .A2(n449), .Y(n1361) );
  NAND4X0_HVT U1502 ( .A1(n400), .A2(n1362), .A3(n1417), .A4(n1361), .Y(
        n_state[1]) );
  NAND4X0_HVT U1503 ( .A1(state[0]), .A2(n1023), .A3(n251), .A4(state[2]), .Y(
        n1563) );
  OA21X1_HVT U1504 ( .A1(n1023), .A2(n1417), .A3(n1563), .Y(n1465) );
  OA22X1_HVT U1505 ( .A1(conv_done), .A2(n1363), .A3(n1391), .A4(n449), .Y(
        n1364) );
  NAND4X0_HVT U1506 ( .A1(state[1]), .A2(state[0]), .A3(n1024), .A4(state[3]), 
        .Y(n1467) );
  NAND3X0_HVT U1507 ( .A1(n1465), .A2(n1364), .A3(n1467), .Y(n_state[2]) );
  NAND2X0_HVT U1508 ( .A1(n1023), .A2(state[2]), .Y(n1369) );
  NAND3X0_HVT U1509 ( .A1(n1023), .A2(n1446), .A3(n1365), .Y(n1366) );
  NAND4X0_HVT U1510 ( .A1(n1369), .A2(n1368), .A3(n1367), .A4(n1366), .Y(
        n_state[3]) );
  NAND2X0_HVT U1511 ( .A1(n205), .A2(n1392), .Y(n1457) );
  NAND3X0_HVT U1512 ( .A1(n1466), .A2(n1458), .A3(n1370), .Y(n1380) );
  NAND2X0_HVT U1513 ( .A1(n1457), .A2(n1371), .Y(n1384) );
  AO22X1_HVT U1514 ( .A1(weight_cnt[0]), .A2(n1380), .A3(n299), .A4(n1384), 
        .Y(n_weight_cnt[0]) );
  AO22X1_HVT U1515 ( .A1(weight_cnt[1]), .A2(n299), .A3(n430), .A4(
        weight_cnt[0]), .Y(n1372) );
  AO22X1_HVT U1516 ( .A1(n1372), .A2(n1384), .A3(weight_cnt[1]), .A4(n1380), 
        .Y(n_weight_cnt[1]) );
  NAND3X0_HVT U1517 ( .A1(weight_cnt[1]), .A2(weight_cnt[0]), .A3(
        weight_cnt[2]), .Y(n1373) );
  AO21X1_HVT U1518 ( .A1(n1384), .A2(n1373), .A3(n1380), .Y(n1374) );
  OA222X1_HVT U1519 ( .A1(weight_cnt[3]), .A2(n1379), .A3(weight_cnt[3]), .A4(
        n1384), .A5(n424), .A6(n1374), .Y(n_weight_cnt[3]) );
  NAND3X0_HVT U1520 ( .A1(weight_cnt[3]), .A2(n1379), .A3(weight_cnt[4]), .Y(
        n1376) );
  OA221X1_HVT U1521 ( .A1(weight_cnt[4]), .A2(n1379), .A3(weight_cnt[4]), .A4(
        weight_cnt[3]), .A5(n1376), .Y(n1375) );
  AO22X1_HVT U1522 ( .A1(n1375), .A2(n1384), .A3(weight_cnt[4]), .A4(n1380), 
        .Y(n_weight_cnt[4]) );
  AO22X1_HVT U1523 ( .A1(n1377), .A2(n439), .A3(n1376), .A4(weight_cnt[5]), 
        .Y(n1378) );
  AO22X1_HVT U1524 ( .A1(n1378), .A2(n1384), .A3(weight_cnt[5]), .A4(n1380), 
        .Y(n_weight_cnt[5]) );
  AND4X1_HVT U1525 ( .A1(weight_cnt[3]), .A2(n1379), .A3(weight_cnt[4]), .A4(
        weight_cnt[5]), .Y(n1381) );
  NAND2X0_HVT U1526 ( .A1(n1381), .A2(weight_cnt[6]), .Y(n1382) );
  AO21X1_HVT U1527 ( .A1(n1384), .A2(n1382), .A3(n1380), .Y(n1383) );
  OA221X1_HVT U1528 ( .A1(weight_cnt[6]), .A2(n1381), .A3(weight_cnt[6]), .A4(
        n1384), .A5(n1383), .Y(n_weight_cnt[6]) );
  OA222X1_HVT U1529 ( .A1(weight_cnt[7]), .A2(n1385), .A3(weight_cnt[7]), .A4(
        n1384), .A5(n448), .A6(n1383), .Y(n_weight_cnt[7]) );
  OR3X1_HVT U1530 ( .A1(conv2_weight_done), .A2(write_enable), .A3(
        load_data_enable), .Y(n1387) );
  OR3X1_HVT U1531 ( .A1(conv1_weight_done), .A2(write_enable), .A3(
        load_data_enable), .Y(n1386) );
  AO22X1_HVT U1532 ( .A1(n1550), .A2(n1387), .A3(n2004), .A4(n1386), .Y(
        n_write_enable) );
  NAND2X0_HVT U1533 ( .A1(n1550), .A2(srstn), .Y(net22461) );
  NAND2X0_HVT U1534 ( .A1(n1566), .A2(col[2]), .Y(n1565) );
  OA221X1_HVT U1535 ( .A1(n1388), .A2(col[3]), .A3(n1565), .A4(n238), .A5(
        n1567), .Y(net22638) );
  AND2X1_HVT U1536 ( .A1(n254), .A2(n1567), .Y(net22653) );
  AO221X1_HVT U1537 ( .A1(sram_raddr_weight[4]), .A2(sram_raddr_weight[3]), 
        .A3(sram_raddr_weight[4]), .A4(sram_raddr_weight[2]), .A5(n1392), .Y(
        n1437) );
  NOR2X0_HVT U1538 ( .A1(n1437), .A2(sram_raddr_weight[5]), .Y(n1440) );
  NAND2X0_HVT U1539 ( .A1(n1440), .A2(n407), .Y(n1434) );
  NAND2X0_HVT U1540 ( .A1(n1429), .A2(n410), .Y(n1430) );
  NAND3X0_HVT U1541 ( .A1(n293), .A2(n395), .A3(n1425), .Y(n1413) );
  OR3X1_HVT U1542 ( .A1(sram_raddr_weight[11]), .A2(sram_raddr_weight[10]), 
        .A3(n1413), .Y(n1406) );
  OR3X1_HVT U1543 ( .A1(sram_raddr_weight[13]), .A2(sram_raddr_weight[12]), 
        .A3(n1406), .Y(n1393) );
  NAND2X0_HVT U1544 ( .A1(n205), .A2(n1393), .Y(n1401) );
  NAND4X0_HVT U1545 ( .A1(sram_raddr_weight[3]), .A2(sram_raddr_weight[2]), 
        .A3(sram_raddr_weight[0]), .A4(sram_raddr_weight[1]), .Y(n1441) );
  NAND2X0_HVT U1546 ( .A1(sram_raddr_weight[4]), .A2(n1445), .Y(n1436) );
  AND3X1_HVT U1547 ( .A1(sram_raddr_weight[5]), .A2(sram_raddr_weight[6]), 
        .A3(n1439), .Y(n1435) );
  AND2X1_HVT U1548 ( .A1(sram_raddr_weight[7]), .A2(n1435), .Y(n1424) );
  NAND2X0_HVT U1549 ( .A1(sram_raddr_weight[8]), .A2(n1424), .Y(n1412) );
  NAND4X0_HVT U1550 ( .A1(sram_raddr_weight[11]), .A2(sram_raddr_weight[9]), 
        .A3(sram_raddr_weight[10]), .A4(n1418), .Y(n1410) );
  AND4X1_HVT U1551 ( .A1(sram_raddr_weight[12]), .A2(sram_raddr_weight[13]), 
        .A3(n1407), .A4(n1456), .Y(n1403) );
  NAND2X0_HVT U1552 ( .A1(sram_raddr_weight[14]), .A2(n1403), .Y(n1399) );
  OR2X1_HVT U1553 ( .A1(n292), .A2(n1399), .Y(n1394) );
  AO221X1_HVT U1554 ( .A1(n1397), .A2(n292), .A3(n1397), .A4(n219), .A5(n451), 
        .Y(n1396) );
  NOR2X0_HVT U1555 ( .A1(n226), .A2(n1393), .Y(n1405) );
  NAND2X0_HVT U1556 ( .A1(n1405), .A2(n362), .Y(n1398) );
  AO221X1_HVT U1557 ( .A1(n1394), .A2(sram_raddr_weight[15]), .A3(n1394), .A4(
        n1398), .A5(sram_raddr_weight[16]), .Y(n1395) );
  NAND2X0_HVT U1558 ( .A1(n1396), .A2(n1395), .Y(net22691) );
  OAI222X1_HVT U1559 ( .A1(sram_raddr_weight[15]), .A2(n1399), .A3(
        sram_raddr_weight[15]), .A4(n1398), .A5(n292), .A6(n1397), .Y(net22698) );
  NAND3X0_HVT U1560 ( .A1(sram_raddr_weight[13]), .A2(sram_raddr_weight[12]), 
        .A3(n1407), .Y(n1400) );
  NAND2X0_HVT U1561 ( .A1(n1456), .A2(n1400), .Y(n1404) );
  NAND2X0_HVT U1562 ( .A1(n1401), .A2(n1404), .Y(n1402) );
  AO222X1_HVT U1563 ( .A1(n362), .A2(n1403), .A3(n362), .A4(n1405), .A5(
        sram_raddr_weight[14]), .A6(n1402), .Y(net22705) );
  AO22X1_HVT U1564 ( .A1(n203), .A2(n1406), .A3(n1456), .A4(n1410), .Y(n1409)
         );
  AO22X1_HVT U1565 ( .A1(n201), .A2(n1411), .A3(n1407), .A4(n1456), .Y(n1408)
         );
  AO22X1_HVT U1566 ( .A1(sram_raddr_weight[12]), .A2(n1409), .A3(n414), .A4(
        n1408), .Y(net22719) );
  AND2X1_HVT U1567 ( .A1(n1456), .A2(n1412), .Y(n1423) );
  AO22X1_HVT U1568 ( .A1(n203), .A2(n1413), .A3(n293), .A4(n1456), .Y(n1416)
         );
  OR2X1_HVT U1569 ( .A1(n219), .A2(n1413), .Y(n1422) );
  NAND3X0_HVT U1570 ( .A1(sram_raddr_weight[9]), .A2(n1418), .A3(n1456), .Y(
        n1414) );
  NAND2X0_HVT U1571 ( .A1(n1422), .A2(n1414), .Y(n1415) );
  AO222X1_HVT U1572 ( .A1(sram_raddr_weight[10]), .A2(n1423), .A3(
        sram_raddr_weight[10]), .A4(n1416), .A5(n415), .A6(n1415), .Y(net22733) );
  NAND3X0_HVT U1573 ( .A1(n1418), .A2(n293), .A3(n1456), .Y(n1421) );
  AO221X1_HVT U1574 ( .A1(n203), .A2(sram_raddr_weight[8]), .A3(n201), .A4(
        n1430), .A5(n1423), .Y(n1419) );
  NAND2X0_HVT U1575 ( .A1(sram_raddr_weight[9]), .A2(n1419), .Y(n1420) );
  NAND4X0_HVT U1576 ( .A1(n283), .A2(n1422), .A3(n1421), .A4(n1420), .Y(
        net22747) );
  NAND2X0_HVT U1577 ( .A1(n1423), .A2(n1424), .Y(n1428) );
  OA22X1_HVT U1578 ( .A1(n1425), .A2(n226), .A3(n1466), .A4(n1424), .Y(n1426)
         );
  AO222X1_HVT U1579 ( .A1(n395), .A2(n219), .A3(n395), .A4(n1430), .A5(
        sram_raddr_weight[8]), .A6(n1426), .Y(n1427) );
  NAND3X0_HVT U1580 ( .A1(n1428), .A2(n1427), .A3(n283), .Y(net22754) );
  OA22X1_HVT U1581 ( .A1(n1429), .A2(n226), .A3(n1466), .A4(n1435), .Y(n1431)
         );
  OA22X1_HVT U1582 ( .A1(n1431), .A2(n410), .A3(n219), .A4(n1430), .Y(n1433)
         );
  NAND3X0_HVT U1583 ( .A1(n1435), .A2(n410), .A3(n1456), .Y(n1432) );
  NAND3X0_HVT U1584 ( .A1(n283), .A2(n1433), .A3(n1432), .Y(net22782) );
  AO22X1_HVT U1585 ( .A1(n203), .A2(n1437), .A3(n1456), .A4(n1436), .Y(n1438)
         );
  NAND2X0_HVT U1586 ( .A1(n1456), .A2(n1441), .Y(n1451) );
  NAND4X0_HVT U1587 ( .A1(n201), .A2(n1442), .A3(n417), .A4(n294), .Y(n1454)
         );
  NAND3X0_HVT U1588 ( .A1(n1457), .A2(n1451), .A3(n1454), .Y(n1449) );
  NAND2X0_HVT U1589 ( .A1(n1442), .A2(n294), .Y(n1450) );
  OR2X1_HVT U1590 ( .A1(sram_raddr_weight[3]), .A2(n1450), .Y(n1443) );
  AO22X1_HVT U1591 ( .A1(n1445), .A2(n1456), .A3(n1444), .A4(n1443), .Y(n1448)
         );
  NAND3X0_HVT U1592 ( .A1(n1023), .A2(n310), .A3(state[2]), .Y(n1562) );
  NAND3X0_HVT U1593 ( .A1(n1023), .A2(n1024), .A3(n1446), .Y(n1551) );
  NAND4X0_HVT U1594 ( .A1(n1465), .A2(n1447), .A3(n1562), .A4(n1551), .Y(n1460) );
  AO221X1_HVT U1595 ( .A1(sram_raddr_weight[4]), .A2(n1449), .A3(n433), .A4(
        n1448), .A5(n1460), .Y(net22810) );
  NAND3X0_HVT U1596 ( .A1(sram_raddr_weight[2]), .A2(sram_raddr_weight[0]), 
        .A3(sram_raddr_weight[1]), .Y(n1452) );
  AOI22X1_HVT U1597 ( .A1(n202), .A2(n1450), .A3(n1456), .A4(n1452), .Y(n1453)
         );
  OA22X1_HVT U1598 ( .A1(n1453), .A2(n417), .A3(n1452), .A4(n1451), .Y(n1455)
         );
  NAND3X0_HVT U1599 ( .A1(n283), .A2(n1455), .A3(n1454), .Y(net22817) );
  NAND2X0_HVT U1600 ( .A1(sram_raddr_weight[0]), .A2(sram_raddr_weight[1]), 
        .Y(n1459) );
  NAND2X0_HVT U1601 ( .A1(n1456), .A2(n1459), .Y(n1463) );
  NAND2X0_HVT U1602 ( .A1(n1457), .A2(n1463), .Y(n1462) );
  OAI21X1_HVT U1603 ( .A1(n1459), .A2(n1466), .A3(n1458), .Y(n1461) );
  AO221X1_HVT U1604 ( .A1(sram_raddr_weight[2]), .A2(n1462), .A3(n294), .A4(
        n1461), .A5(n1460), .Y(net22824) );
  AO222X1_HVT U1605 ( .A1(n421), .A2(n1463), .A3(n421), .A4(n300), .A5(n1463), 
        .A6(n226), .Y(n1464) );
  NAND2X0_HVT U1606 ( .A1(n1465), .A2(n1464), .Y(net22838) );
  AO22X1_HVT U1607 ( .A1(sram_raddr_weight[0]), .A2(n219), .A3(n300), .A4(
        n1466), .Y(n1468) );
  NAND3X0_HVT U1608 ( .A1(n1468), .A2(n1467), .A3(n1562), .Y(net22852) );
  NAND2X0_HVT U1609 ( .A1(write_col_conv1[0]), .A2(n1469), .Y(n1508) );
  AO21X1_HVT U1610 ( .A1(n1471), .A2(n1470), .A3(N2914), .Y(net22860) );
  NAND2X0_HVT U1611 ( .A1(n1473), .A2(write_row_conv1[0]), .Y(n1477) );
  NAND3X0_HVT U1612 ( .A1(write_col_conv1[0]), .A2(n1474), .A3(n1477), .Y(
        n1499) );
  NAND2X0_HVT U1613 ( .A1(n1495), .A2(n376), .Y(n1493) );
  NOR2X0_HVT U1614 ( .A1(n1493), .A2(delay1_sram_waddr_b[5]), .Y(n1489) );
  NAND2X0_HVT U1615 ( .A1(n1489), .A2(n375), .Y(n1487) );
  NOR2X0_HVT U1616 ( .A1(n1487), .A2(delay1_sram_waddr_b[7]), .Y(n1484) );
  NAND2X0_HVT U1617 ( .A1(n1484), .A2(n431), .Y(n1475) );
  HADDX1_HVT U1618 ( .A0(delay1_sram_waddr_b[9]), .B0(n1475), .SO(n1480) );
  NAND4X0_HVT U1619 ( .A1(delay1_sram_waddr_b[0]), .A2(delay1_sram_waddr_b[1]), 
        .A3(delay1_sram_waddr_b[2]), .A4(delay1_sram_waddr_b[3]), .Y(n1496) );
  NOR2X0_HVT U1620 ( .A1(n376), .A2(n1496), .Y(n1494) );
  NAND2X0_HVT U1621 ( .A1(delay1_sram_waddr_b[5]), .A2(n1494), .Y(n1490) );
  NOR2X0_HVT U1622 ( .A1(n375), .A2(n1490), .Y(n1488) );
  AND2X1_HVT U1623 ( .A1(delay1_sram_waddr_b[7]), .A2(n1488), .Y(n1483) );
  NAND2X0_HVT U1624 ( .A1(delay1_sram_waddr_b[8]), .A2(n1483), .Y(n1478) );
  HADDX1_HVT U1625 ( .A0(delay1_sram_waddr_b[9]), .B0(n1478), .SO(n1479) );
  OAI22X1_HVT U1626 ( .A1(n1499), .A2(n1480), .A3(n1501), .A4(n1479), .Y(
        net22863) );
  OAI22X1_HVT U1627 ( .A1(n1484), .A2(n1499), .A3(n1483), .A4(n1501), .Y(n1482) );
  AO22X1_HVT U1628 ( .A1(n1506), .A2(n1484), .A3(n1507), .A4(n1483), .Y(n1481)
         );
  AO22X1_HVT U1629 ( .A1(delay1_sram_waddr_b[8]), .A2(n1482), .A3(n431), .A4(
        n1481), .Y(net22866) );
  OA221X1_HVT U1630 ( .A1(n1484), .A2(delay1_sram_waddr_b[7]), .A3(n1484), 
        .A4(n1487), .A5(n1506), .Y(n1485) );
  AO221X1_HVT U1631 ( .A1(n1486), .A2(delay1_sram_waddr_b[7]), .A3(n1486), 
        .A4(n1488), .A5(n1485), .Y(net22869) );
  AO21X1_HVT U1632 ( .A1(delay1_sram_waddr_b[5]), .A2(n1493), .A3(n1489), .Y(
        n1492) );
  OA21X1_HVT U1633 ( .A1(delay1_sram_waddr_b[5]), .A2(n1494), .A3(n1490), .Y(
        n1491) );
  AO22X1_HVT U1634 ( .A1(n1506), .A2(n1492), .A3(n1507), .A4(n1491), .Y(
        net22875) );
  OR3X1_HVT U1635 ( .A1(delay1_sram_waddr_b[0]), .A2(delay1_sram_waddr_b[1]), 
        .A3(delay1_sram_waddr_b[2]), .Y(n1500) );
  AO21X1_HVT U1636 ( .A1(delay1_sram_waddr_b[3]), .A2(n1500), .A3(n1495), .Y(
        n1498) );
  AND3X1_HVT U1637 ( .A1(delay1_sram_waddr_b[0]), .A2(delay1_sram_waddr_b[1]), 
        .A3(delay1_sram_waddr_b[2]), .Y(n1502) );
  OA21X1_HVT U1638 ( .A1(delay1_sram_waddr_b[3]), .A2(n1502), .A3(n1496), .Y(
        n1497) );
  AO22X1_HVT U1639 ( .A1(n1506), .A2(n1498), .A3(n1507), .A4(n1497), .Y(
        net22881) );
  OR2X1_HVT U1640 ( .A1(delay1_sram_waddr_b[0]), .A2(delay1_sram_waddr_b[1]), 
        .Y(n1504) );
  NAND2X0_HVT U1641 ( .A1(delay1_sram_waddr_b[0]), .A2(delay1_sram_waddr_b[1]), 
        .Y(n1503) );
  NAND2X0_HVT U1642 ( .A1(n1504), .A2(n1503), .Y(n1505) );
  MUX21X1_HVT U1643 ( .A1(n1507), .A2(n1506), .S0(n1505), .Y(net22887) );
  NOR2X0_HVT U1644 ( .A1(n1508), .A2(delay1_sram_waddr_b[0]), .Y(net22890) );
  AND4X1_HVT U1645 ( .A1(delay3_state[2]), .A2(n1027), .A3(delay3_state[0]), 
        .A4(delay3_state[1]), .Y(n1529) );
  NAND4X0_HVT U1646 ( .A1(n1529), .A2(delay3_addr_change[0]), .A3(
        delay3_addr_change[1]), .A4(n1509), .Y(n1512) );
  NAND2X0_HVT U1647 ( .A1(delay3_state[2]), .A2(n1027), .Y(n1510) );
  OR3X1_HVT U1648 ( .A1(delay3_state[0]), .A2(delay3_state[1]), .A3(n1510), 
        .Y(n1511) );
  NAND3X0_HVT U1649 ( .A1(srstn), .A2(n1512), .A3(n1511), .Y(net22898) );
  NAND4X0_HVT U1650 ( .A1(delay1_sram_waddr_c[0]), .A2(delay1_sram_waddr_c[1]), 
        .A3(delay1_sram_waddr_c[2]), .A4(delay1_sram_waddr_c[3]), .Y(n1525) );
  NAND2X0_HVT U1651 ( .A1(n1524), .A2(delay1_sram_waddr_c[4]), .Y(n1523) );
  NAND2X0_HVT U1652 ( .A1(n1522), .A2(delay1_sram_waddr_c[5]), .Y(n1521) );
  NAND2X0_HVT U1653 ( .A1(n1520), .A2(delay1_sram_waddr_c[6]), .Y(n1519) );
  NAND2X0_HVT U1654 ( .A1(n1518), .A2(delay1_sram_waddr_c[7]), .Y(n1517) );
  NAND2X0_HVT U1655 ( .A1(n1516), .A2(delay1_sram_waddr_c[8]), .Y(n1515) );
  OA221X1_HVT U1656 ( .A1(n1514), .A2(delay1_sram_waddr_c[9]), .A3(n1515), 
        .A4(n454), .A5(n1528), .Y(net22900) );
  NAND3X0_HVT U1657 ( .A1(delay1_sram_waddr_c[0]), .A2(delay1_sram_waddr_c[1]), 
        .A3(delay1_sram_waddr_c[2]), .Y(n1526) );
  NAND2X0_HVT U1658 ( .A1(delay1_sram_waddr_c[0]), .A2(delay1_sram_waddr_c[1]), 
        .Y(n1527) );
  AND2X1_HVT U1659 ( .A1(n1528), .A2(n425), .Y(net22909) );
  NAND4X0_HVT U1660 ( .A1(delay1_sram_waddr_d[0]), .A2(delay1_sram_waddr_d[1]), 
        .A3(delay1_sram_waddr_d[2]), .A4(delay1_sram_waddr_d[3]), .Y(n1541) );
  NAND2X0_HVT U1661 ( .A1(n1540), .A2(delay1_sram_waddr_d[4]), .Y(n1539) );
  NAND2X0_HVT U1662 ( .A1(n1538), .A2(delay1_sram_waddr_d[5]), .Y(n1537) );
  NAND2X0_HVT U1663 ( .A1(n1536), .A2(delay1_sram_waddr_d[6]), .Y(n1535) );
  NAND2X0_HVT U1664 ( .A1(n1534), .A2(delay1_sram_waddr_d[7]), .Y(n1533) );
  NAND2X0_HVT U1665 ( .A1(n1532), .A2(delay1_sram_waddr_d[8]), .Y(n1531) );
  OA221X1_HVT U1666 ( .A1(n1530), .A2(delay1_sram_waddr_d[9]), .A3(n1531), 
        .A4(n455), .A5(n1544), .Y(net22916) );
  NAND3X0_HVT U1667 ( .A1(delay1_sram_waddr_d[0]), .A2(delay1_sram_waddr_d[1]), 
        .A3(delay1_sram_waddr_d[2]), .Y(n1542) );
  NAND2X0_HVT U1668 ( .A1(delay1_sram_waddr_d[0]), .A2(delay1_sram_waddr_d[1]), 
        .Y(n1543) );
  AND2X1_HVT U1669 ( .A1(n1544), .A2(n426), .Y(net22925) );
  NAND2X0_HVT U1670 ( .A1(n1545), .A2(srstn), .Y(net22932) );
  NAND3X0_HVT U1671 ( .A1(n1548), .A2(channel_cnt[2]), .A3(channel_cnt[3]), 
        .Y(n1547) );
  OA221X1_HVT U1672 ( .A1(channel_cnt[4]), .A2(n1546), .A3(n311), .A4(n1547), 
        .A5(n1550), .Y(net22933) );
  OA221X1_HVT U1673 ( .A1(n1548), .A2(channel_cnt[2]), .A3(n1549), .A4(n420), 
        .A5(n1550), .Y(net22935) );
  NAND3X0_HVT U1674 ( .A1(srstn), .A2(n219), .A3(n1551), .Y(net22943) );
  NAND4X0_HVT U1675 ( .A1(addr_change[0]), .A2(addr_change[1]), .A3(
        addr_change[2]), .A4(addr_change[3]), .Y(n1554) );
  NAND4X0_HVT U1676 ( .A1(addr_change[1]), .A2(addr_change[0]), .A3(
        addr_change[4]), .A4(n441), .Y(n1552) );
  OA21X1_HVT U1677 ( .A1(addr_change[2]), .A2(n1552), .A3(n202), .Y(n1557) );
  OA221X1_HVT U1678 ( .A1(addr_change[4]), .A2(n1553), .A3(n447), .A4(n1554), 
        .A5(n1557), .Y(net22945) );
  NAND3X0_HVT U1679 ( .A1(addr_change[0]), .A2(addr_change[1]), .A3(
        addr_change[2]), .Y(n1555) );
  NAND2X0_HVT U1680 ( .A1(addr_change[0]), .A2(addr_change[1]), .Y(n1556) );
  NOR2X0_HVT U1681 ( .A1(n219), .A2(addr_change[0]), .Y(net22949) );
  NAND4X0_HVT U1682 ( .A1(n1570), .A2(n1559), .A3(addr_row_sel_cnt[0]), .A4(
        addr_row_sel_cnt[1]), .Y(n1560) );
  OA221X1_HVT U1683 ( .A1(n1569), .A2(n1051), .A3(n1569), .A4(
        addr_col_sel_cnt[0]), .A5(n1560), .Y(n1893) );
  NAND2X0_HVT U1684 ( .A1(srstn), .A2(n1935), .Y(net23892) );
  NAND2X0_HVT U1685 ( .A1(srstn), .A2(n1990), .Y(net25219) );
  NAND2X0_HVT U1686 ( .A1(n181), .A2(n1888), .Y(net26549) );
  NOR2X0_HVT U1687 ( .A1(n251), .A2(n1562), .Y(n1022) );
  NAND3X0_HVT U1688 ( .A1(n1051), .A2(n1052), .A3(n1680), .Y(n1850) );
  AND4X1_HVT U1689 ( .A1(n1570), .A2(n2004), .A3(addr_row_sel_cnt[1]), .A4(
        n250), .Y(n1572) );
  AO22X1_HVT U1690 ( .A1(n1839), .A2(n295), .A3(n170), .A4(n418), .Y(n1573) );
  AO221X1_HVT U1691 ( .A1(sram_raddr_a0[0]), .A2(n1888), .A3(n416), .A4(n1615), 
        .A5(n1573), .Y(n_sram_raddr_a0[0]) );
  NAND2X0_HVT U1692 ( .A1(sram_raddr_a6[1]), .A2(sram_raddr_a6[0]), .Y(n1579)
         );
  OA21X1_HVT U1693 ( .A1(sram_raddr_a6[1]), .A2(sram_raddr_a6[0]), .A3(n1579), 
        .Y(n1851) );
  NAND2X0_HVT U1694 ( .A1(n521), .A2(n1851), .Y(n1736) );
  AO221X1_HVT U1695 ( .A1(n1760), .A2(n1578), .A3(n1760), .A4(sram_raddr_a0[0]), .A5(n297), .Y(n1576) );
  NAND3X0_HVT U1696 ( .A1(sram_raddr_a0[0]), .A2(n1615), .A3(n297), .Y(n1575)
         );
  NAND2X0_HVT U1697 ( .A1(sram_raddr_a3[1]), .A2(sram_raddr_a3[0]), .Y(n1581)
         );
  OA21X1_HVT U1698 ( .A1(sram_raddr_a3[1]), .A2(sram_raddr_a3[0]), .A3(n1581), 
        .Y(n1737) );
  NAND2X0_HVT U1699 ( .A1(n1975), .A2(n1737), .Y(n1574) );
  NAND4X0_HVT U1700 ( .A1(n1736), .A2(n1576), .A3(n1575), .A4(n1574), .Y(
        n_sram_raddr_a0[1]) );
  AND3X1_HVT U1701 ( .A1(sram_raddr_a0[2]), .A2(sram_raddr_a0[1]), .A3(
        sram_raddr_a0[0]), .Y(n1577) );
  OA21X1_HVT U1702 ( .A1(n1578), .A2(n1577), .A3(n1760), .Y(n1586) );
  AND3X1_HVT U1703 ( .A1(sram_raddr_a0[1]), .A2(sram_raddr_a0[0]), .A3(n1615), 
        .Y(n1582) );
  AO22X1_HVT U1704 ( .A1(n1583), .A2(n443), .A3(n1579), .A4(sram_raddr_a6[2]), 
        .Y(n1852) );
  AO22X1_HVT U1705 ( .A1(sram_raddr_a3[2]), .A2(n1581), .A3(n234), .A4(n1580), 
        .Y(n1739) );
  NAND4X0_HVT U1706 ( .A1(sram_raddr_a3[2]), .A2(sram_raddr_a3[3]), .A3(
        sram_raddr_a3[1]), .A4(sram_raddr_a3[0]), .Y(n1588) );
  AO221X1_HVT U1707 ( .A1(n245), .A2(n234), .A3(n245), .A4(n1581), .A5(n1587), 
        .Y(n1740) );
  OA22X1_HVT U1708 ( .A1(n1586), .A2(n237), .A3(n171), .A4(n1740), .Y(n1584)
         );
  NAND3X0_HVT U1709 ( .A1(sram_raddr_a0[2]), .A2(n1582), .A3(n237), .Y(n1585)
         );
  NAND4X0_HVT U1710 ( .A1(sram_raddr_a6[1]), .A2(sram_raddr_a6[0]), .A3(
        sram_raddr_a6[2]), .A4(sram_raddr_a6[3]), .Y(n1589) );
  OA221X1_HVT U1711 ( .A1(sram_raddr_a6[3]), .A2(sram_raddr_a6[2]), .A3(
        sram_raddr_a6[3]), .A4(n1583), .A5(n1589), .Y(n1853) );
  NAND2X0_HVT U1712 ( .A1(n168), .A2(n1853), .Y(n1741) );
  NAND3X0_HVT U1713 ( .A1(n1584), .A2(n1585), .A3(n1741), .Y(
        n_sram_raddr_a0[3]) );
  AND2X1_HVT U1714 ( .A1(n1586), .A2(n1585), .Y(n1596) );
  AND2X1_HVT U1715 ( .A1(sram_raddr_a3[4]), .A2(n1587), .Y(n1592) );
  AO21X1_HVT U1716 ( .A1(n279), .A2(n1588), .A3(n1592), .Y(n1746) );
  OA22X1_HVT U1717 ( .A1(n1596), .A2(n367), .A3(n189), .A4(n1746), .Y(n1591)
         );
  AND4X1_HVT U1718 ( .A1(sram_raddr_a0[3]), .A2(sram_raddr_a0[2]), .A3(
        sram_raddr_a0[1]), .A4(sram_raddr_a0[0]), .Y(n1601) );
  NAND3X0_HVT U1719 ( .A1(n1601), .A2(n1615), .A3(n367), .Y(n1595) );
  NAND2X0_HVT U1720 ( .A1(n1590), .A2(sram_raddr_a6[4]), .Y(n1593) );
  OA21X1_HVT U1721 ( .A1(n1590), .A2(sram_raddr_a6[4]), .A3(n1593), .Y(n1857)
         );
  NAND2X0_HVT U1722 ( .A1(n521), .A2(n1857), .Y(n1744) );
  NAND3X0_HVT U1723 ( .A1(n1591), .A2(n1595), .A3(n1744), .Y(
        n_sram_raddr_a0[4]) );
  NAND2X0_HVT U1724 ( .A1(sram_raddr_a3[5]), .A2(n1592), .Y(n1600) );
  OA21X1_HVT U1725 ( .A1(sram_raddr_a3[5]), .A2(n1592), .A3(n1600), .Y(n1748)
         );
  NAND2X0_HVT U1726 ( .A1(n170), .A2(n1748), .Y(n1599) );
  NAND2X0_HVT U1727 ( .A1(n1594), .A2(sram_raddr_a6[5]), .Y(n1602) );
  OA21X1_HVT U1728 ( .A1(n1594), .A2(sram_raddr_a6[5]), .A3(n1602), .Y(n1863)
         );
  NAND2X0_HVT U1729 ( .A1(n168), .A2(n1863), .Y(n1751) );
  NAND4X0_HVT U1730 ( .A1(sram_raddr_a0[4]), .A2(n1601), .A3(n1615), .A4(n291), 
        .Y(n1597) );
  AND3X1_HVT U1731 ( .A1(n1596), .A2(n1597), .A3(n1595), .Y(n1605) );
  AO21X1_HVT U1732 ( .A1(n291), .A2(n1597), .A3(n1605), .Y(n1598) );
  NAND3X0_HVT U1733 ( .A1(n1599), .A2(n1751), .A3(n1598), .Y(
        n_sram_raddr_a0[5]) );
  OR2X1_HVT U1734 ( .A1(n349), .A2(n1600), .Y(n1607) );
  AO21X1_HVT U1735 ( .A1(n349), .A2(n1600), .A3(n1606), .Y(n1756) );
  OA22X1_HVT U1736 ( .A1(n1605), .A2(n432), .A3(n189), .A4(n1756), .Y(n1603)
         );
  AND3X1_HVT U1737 ( .A1(sram_raddr_a0[5]), .A2(sram_raddr_a0[4]), .A3(n1601), 
        .Y(n1610) );
  NAND3X0_HVT U1738 ( .A1(n1610), .A2(n1615), .A3(n432), .Y(n1604) );
  AO22X1_HVT U1739 ( .A1(n1608), .A2(n452), .A3(n1602), .A4(sram_raddr_a6[6]), 
        .Y(n1868) );
  NAND2X0_HVT U1740 ( .A1(n1839), .A2(n1868), .Y(n1754) );
  NAND3X0_HVT U1741 ( .A1(n1603), .A2(n1604), .A3(n1754), .Y(
        n_sram_raddr_a0[6]) );
  AND2X1_HVT U1742 ( .A1(n1605), .A2(n1604), .Y(n1614) );
  AND2X1_HVT U1743 ( .A1(sram_raddr_a3[7]), .A2(n1606), .Y(n1619) );
  AO21X1_HVT U1744 ( .A1(n383), .A2(n1607), .A3(n1619), .Y(n1758) );
  OA22X1_HVT U1745 ( .A1(n1614), .A2(n355), .A3(n189), .A4(n1758), .Y(n1612)
         );
  AND2X1_HVT U1746 ( .A1(n1608), .A2(sram_raddr_a6[6]), .Y(n1609) );
  NAND2X0_HVT U1747 ( .A1(n1609), .A2(sram_raddr_a6[7]), .Y(n1617) );
  OA21X1_HVT U1748 ( .A1(n1609), .A2(sram_raddr_a6[7]), .A3(n1617), .Y(n1874)
         );
  NAND2X0_HVT U1749 ( .A1(n168), .A2(n1874), .Y(n1763) );
  AND2X1_HVT U1750 ( .A1(sram_raddr_a0[6]), .A2(n1610), .Y(n1616) );
  NAND3X0_HVT U1751 ( .A1(n1616), .A2(n355), .A3(n1615), .Y(n1611) );
  NAND3X0_HVT U1752 ( .A1(n1612), .A2(n1763), .A3(n1611), .Y(
        n_sram_raddr_a0[7]) );
  NAND2X0_HVT U1753 ( .A1(n355), .A2(n1615), .Y(n1613) );
  NAND2X0_HVT U1754 ( .A1(n1614), .A2(n1613), .Y(n1627) );
  AND3X1_HVT U1755 ( .A1(sram_raddr_a0[7]), .A2(n1616), .A3(n1615), .Y(n1625)
         );
  NAND2X0_HVT U1756 ( .A1(n1618), .A2(sram_raddr_a6[8]), .Y(n1621) );
  OA21X1_HVT U1757 ( .A1(n1618), .A2(sram_raddr_a6[8]), .A3(n1621), .Y(n1881)
         );
  NAND2X0_HVT U1758 ( .A1(sram_raddr_a3[8]), .A2(n1619), .Y(n1623) );
  OA21X1_HVT U1759 ( .A1(sram_raddr_a3[8]), .A2(n1619), .A3(n1623), .Y(n1766)
         );
  AO22X1_HVT U1760 ( .A1(n521), .A2(n1881), .A3(n170), .A4(n1766), .Y(n1620)
         );
  AO221X1_HVT U1761 ( .A1(sram_raddr_a0[8]), .A2(n1627), .A3(n402), .A4(n1625), 
        .A5(n1620), .Y(n_sram_raddr_a0[8]) );
  HADDX1_HVT U1762 ( .A0(sram_raddr_a6[9]), .B0(n1622), .SO(n1887) );
  AND2X1_HVT U1763 ( .A1(n521), .A2(n1887), .Y(n1773) );
  HADDX1_HVT U1764 ( .A0(sram_raddr_a3[9]), .B0(n1624), .SO(n1771) );
  HADDX1_HVT U1765 ( .A0(sram_raddr_a0[9]), .B0(sram_raddr_a0[8]), .SO(n1626)
         );
  NAND2X0_HVT U1766 ( .A1(n_addr_col_sel_cnt[1]), .A2(n250), .Y(n1914) );
  AO22X1_HVT U1767 ( .A1(n1839), .A2(n289), .A3(n170), .A4(n396), .Y(n1628) );
  AO221X1_HVT U1768 ( .A1(sram_raddr_a1[0]), .A2(n1935), .A3(n301), .A4(n1665), 
        .A5(n1628), .Y(n_sram_raddr_a1[0]) );
  NAND2X0_HVT U1769 ( .A1(sram_raddr_a4[1]), .A2(sram_raddr_a4[0]), .Y(n1629)
         );
  AO21X1_HVT U1770 ( .A1(n298), .A2(n396), .A3(n1630), .Y(n1775) );
  AO22X1_HVT U1771 ( .A1(sram_raddr_a7[1]), .A2(n289), .A3(n429), .A4(
        sram_raddr_a7[0]), .Y(n1892) );
  NAND2X0_HVT U1772 ( .A1(n168), .A2(n1892), .Y(n1776) );
  AND2X1_HVT U1773 ( .A1(sram_raddr_a1[1]), .A2(sram_raddr_a1[0]), .Y(n1638)
         );
  NAND3X0_HVT U1774 ( .A1(sram_raddr_a1[2]), .A2(sram_raddr_a1[1]), .A3(
        sram_raddr_a1[0]), .Y(n1636) );
  AO21X1_HVT U1775 ( .A1(n1665), .A2(n1636), .A3(n1935), .Y(n1631) );
  AO22X1_HVT U1776 ( .A1(sram_raddr_a4[2]), .A2(n1629), .A3(n235), .A4(n1630), 
        .Y(n1778) );
  NAND3X0_HVT U1777 ( .A1(sram_raddr_a7[1]), .A2(sram_raddr_a7[0]), .A3(
        sram_raddr_a7[2]), .Y(n1632) );
  OA221X1_HVT U1778 ( .A1(sram_raddr_a7[2]), .A2(sram_raddr_a7[0]), .A3(
        sram_raddr_a7[2]), .A4(sram_raddr_a7[1]), .A5(n1632), .Y(n1898) );
  NAND4X0_HVT U1779 ( .A1(sram_raddr_a4[2]), .A2(sram_raddr_a4[3]), .A3(
        sram_raddr_a4[1]), .A4(sram_raddr_a4[0]), .Y(n1637) );
  OA221X1_HVT U1780 ( .A1(sram_raddr_a4[3]), .A2(sram_raddr_a4[2]), .A3(
        sram_raddr_a4[3]), .A4(n1630), .A5(n1637), .Y(n1779) );
  AOI22X1_HVT U1781 ( .A1(sram_raddr_a1[3]), .A2(n1631), .A3(n170), .A4(n1779), 
        .Y(n1635) );
  NAND4X0_HVT U1782 ( .A1(sram_raddr_a1[2]), .A2(n1638), .A3(n1665), .A4(n236), 
        .Y(n1634) );
  AO22X1_HVT U1783 ( .A1(n1633), .A2(n453), .A3(n1632), .A4(sram_raddr_a7[3]), 
        .Y(n1899) );
  NAND2X0_HVT U1784 ( .A1(n1839), .A2(n1899), .Y(n1780) );
  NAND3X0_HVT U1785 ( .A1(n1635), .A2(n1634), .A3(n1780), .Y(
        n_sram_raddr_a1[3]) );
  AOI221X1_HVT U1786 ( .A1(n1665), .A2(n236), .A3(n1665), .A4(n1636), .A5(
        n1935), .Y(n1642) );
  NOR2X0_HVT U1787 ( .A1(n246), .A2(n1637), .Y(n1643) );
  AO21X1_HVT U1788 ( .A1(n246), .A2(n1637), .A3(n1643), .Y(n1782) );
  OA22X1_HVT U1789 ( .A1(n1642), .A2(n282), .A3(n171), .A4(n1782), .Y(n1640)
         );
  AND4X1_HVT U1790 ( .A1(sram_raddr_a1[3]), .A2(sram_raddr_a1[2]), .A3(n1638), 
        .A4(n1665), .Y(n1644) );
  NAND2X0_HVT U1791 ( .A1(n1644), .A2(n282), .Y(n1641) );
  AND4X1_HVT U1792 ( .A1(sram_raddr_a7[1]), .A2(sram_raddr_a7[0]), .A3(
        sram_raddr_a7[2]), .A4(sram_raddr_a7[3]), .Y(n1639) );
  NAND2X0_HVT U1793 ( .A1(n1639), .A2(sram_raddr_a7[4]), .Y(n1645) );
  OA21X1_HVT U1794 ( .A1(n1639), .A2(sram_raddr_a7[4]), .A3(n1645), .Y(n1903)
         );
  NAND2X0_HVT U1795 ( .A1(n168), .A2(n1903), .Y(n1785) );
  NAND3X0_HVT U1796 ( .A1(n1640), .A2(n1641), .A3(n1785), .Y(
        n_sram_raddr_a1[4]) );
  AND2X1_HVT U1797 ( .A1(n1642), .A2(n1641), .Y(n1649) );
  NAND2X0_HVT U1798 ( .A1(sram_raddr_a4[5]), .A2(n1643), .Y(n1650) );
  OA22X1_HVT U1799 ( .A1(n1649), .A2(n380), .A3(n189), .A4(n1787), .Y(n1647)
         );
  AND2X1_HVT U1800 ( .A1(sram_raddr_a1[4]), .A2(n1644), .Y(n1651) );
  NAND2X0_HVT U1801 ( .A1(n1651), .A2(n380), .Y(n1648) );
  NAND2X0_HVT U1802 ( .A1(n1646), .A2(sram_raddr_a7[5]), .Y(n1652) );
  OA21X1_HVT U1803 ( .A1(n1646), .A2(sram_raddr_a7[5]), .A3(n1652), .Y(n1909)
         );
  NAND2X0_HVT U1804 ( .A1(n168), .A2(n1909), .Y(n1789) );
  NAND3X0_HVT U1805 ( .A1(n1647), .A2(n1648), .A3(n1789), .Y(
        n_sram_raddr_a1[5]) );
  AND2X1_HVT U1806 ( .A1(n1649), .A2(n1648), .Y(n1657) );
  AO21X1_HVT U1807 ( .A1(n353), .A2(n1650), .A3(n1661), .Y(n1794) );
  OA22X1_HVT U1808 ( .A1(n1657), .A2(n434), .A3(n189), .A4(n1794), .Y(n1654)
         );
  AND2X1_HVT U1809 ( .A1(sram_raddr_a1[5]), .A2(n1651), .Y(n1658) );
  NAND2X0_HVT U1810 ( .A1(n1658), .A2(n434), .Y(n1656) );
  NAND2X0_HVT U1811 ( .A1(n1653), .A2(sram_raddr_a7[6]), .Y(n1659) );
  OA21X1_HVT U1812 ( .A1(n1653), .A2(sram_raddr_a7[6]), .A3(n1659), .Y(n1915)
         );
  NAND2X0_HVT U1813 ( .A1(n1839), .A2(n1915), .Y(n1792) );
  NAND3X0_HVT U1814 ( .A1(n1654), .A2(n1656), .A3(n1792), .Y(
        n_sram_raddr_a1[6]) );
  NAND2X0_HVT U1815 ( .A1(n1657), .A2(n1656), .Y(n1664) );
  AND2X1_HVT U1816 ( .A1(sram_raddr_a1[6]), .A2(n1658), .Y(n1666) );
  NAND2X0_HVT U1817 ( .A1(n1660), .A2(sram_raddr_a7[7]), .Y(n1668) );
  OA21X1_HVT U1818 ( .A1(n1660), .A2(sram_raddr_a7[7]), .A3(n1668), .Y(n1923)
         );
  NAND2X0_HVT U1819 ( .A1(sram_raddr_a4[7]), .A2(n1661), .Y(n1670) );
  OA21X1_HVT U1820 ( .A1(sram_raddr_a4[7]), .A2(n1661), .A3(n1670), .Y(n1798)
         );
  AO22X1_HVT U1821 ( .A1(n521), .A2(n1923), .A3(n1975), .A4(n1798), .Y(n1663)
         );
  AO221X1_HVT U1822 ( .A1(sram_raddr_a1[7]), .A2(n1664), .A3(n423), .A4(n1666), 
        .A5(n1663), .Y(n_sram_raddr_a1[7]) );
  AO21X1_HVT U1823 ( .A1(n423), .A2(n1665), .A3(n1664), .Y(n1679) );
  AND2X1_HVT U1824 ( .A1(sram_raddr_a1[7]), .A2(n1666), .Y(n1677) );
  NAND2X0_HVT U1825 ( .A1(n1669), .A2(sram_raddr_a7[8]), .Y(n1673) );
  OA21X1_HVT U1826 ( .A1(n1669), .A2(sram_raddr_a7[8]), .A3(n1673), .Y(n1926)
         );
  NAND2X0_HVT U1827 ( .A1(sram_raddr_a4[8]), .A2(n1671), .Y(n1675) );
  OA21X1_HVT U1828 ( .A1(sram_raddr_a4[8]), .A2(n1671), .A3(n1675), .Y(n1800)
         );
  AO22X1_HVT U1829 ( .A1(n521), .A2(n1926), .A3(n170), .A4(n1800), .Y(n1672)
         );
  AO221X1_HVT U1830 ( .A1(sram_raddr_a1[8]), .A2(n1679), .A3(n403), .A4(n1677), 
        .A5(n1672), .Y(n_sram_raddr_a1[8]) );
  HADDX1_HVT U1831 ( .A0(sram_raddr_a7[9]), .B0(n1674), .SO(n1933) );
  AND2X1_HVT U1832 ( .A1(n1839), .A2(n1933), .Y(n1807) );
  HADDX1_HVT U1833 ( .A0(sram_raddr_a4[9]), .B0(n1676), .SO(n1805) );
  HADDX1_HVT U1834 ( .A0(sram_raddr_a1[9]), .B0(sram_raddr_a1[8]), .SO(n1678)
         );
  NAND3X0_HVT U1835 ( .A1(n1052), .A2(n1680), .A3(addr_col_sel_cnt[1]), .Y(
        n1942) );
  AO22X1_HVT U1836 ( .A1(n1839), .A2(n288), .A3(n1975), .A4(n394), .Y(n1681)
         );
  AO221X1_HVT U1837 ( .A1(sram_raddr_a2[0]), .A2(n1990), .A3(n427), .A4(n1722), 
        .A5(n1681), .Y(n_sram_raddr_a2[0]) );
  AO22X1_HVT U1838 ( .A1(sram_raddr_a8[1]), .A2(n288), .A3(n437), .A4(
        sram_raddr_a8[0]), .Y(n1939) );
  NAND2X0_HVT U1839 ( .A1(sram_raddr_a5[1]), .A2(sram_raddr_a5[0]), .Y(n1688)
         );
  OA21X1_HVT U1840 ( .A1(sram_raddr_a5[1]), .A2(sram_raddr_a5[0]), .A3(n1688), 
        .Y(n1808) );
  NAND2X0_HVT U1841 ( .A1(sram_raddr_a2[1]), .A2(sram_raddr_a2[0]), .Y(n1686)
         );
  OA21X1_HVT U1842 ( .A1(sram_raddr_a2[1]), .A2(sram_raddr_a2[0]), .A3(n1686), 
        .Y(n1682) );
  AO222X1_HVT U1843 ( .A1(n1839), .A2(n1939), .A3(n170), .A4(n1808), .A5(n1682), .A6(n1897), .Y(n1941) );
  AO22X1_HVT U1844 ( .A1(n1982), .A2(n1682), .A3(sram_raddr_a2[1]), .A4(n1990), 
        .Y(n1683) );
  OR2X1_HVT U1845 ( .A1(n1941), .A2(n1683), .Y(n_sram_raddr_a2[1]) );
  NAND2X0_HVT U1846 ( .A1(sram_raddr_a8[1]), .A2(sram_raddr_a8[0]), .Y(n1684)
         );
  AND3X1_HVT U1847 ( .A1(sram_raddr_a8[1]), .A2(sram_raddr_a8[0]), .A3(
        sram_raddr_a8[2]), .Y(n1690) );
  AO21X1_HVT U1848 ( .A1(n1684), .A2(n438), .A3(n1690), .Y(n1944) );
  NAND3X0_HVT U1849 ( .A1(sram_raddr_a5[2]), .A2(sram_raddr_a5[1]), .A3(
        sram_raddr_a5[0]), .Y(n1685) );
  NAND2X0_HVT U1850 ( .A1(n411), .A2(n1688), .Y(n1952) );
  NAND2X0_HVT U1851 ( .A1(n1685), .A2(n1952), .Y(n1947) );
  OA22X1_HVT U1852 ( .A1(n1943), .A2(n1944), .A3(n171), .A4(n1947), .Y(n1812)
         );
  AND3X1_HVT U1853 ( .A1(sram_raddr_a2[2]), .A2(sram_raddr_a2[1]), .A3(
        sram_raddr_a2[0]), .Y(n1708) );
  AND2X1_HVT U1854 ( .A1(n440), .A2(n1686), .Y(n1814) );
  OR2X1_HVT U1855 ( .A1(n1708), .A2(n1814), .Y(n1810) );
  OA22X1_HVT U1856 ( .A1(n1693), .A2(n1810), .A3(n1946), .A4(n440), .Y(n1687)
         );
  NAND2X0_HVT U1857 ( .A1(n1812), .A2(n1687), .Y(n_sram_raddr_a2[2]) );
  OA21X1_HVT U1858 ( .A1(n1693), .A2(n1708), .A3(n1946), .Y(n1689) );
  AND4X1_HVT U1859 ( .A1(sram_raddr_a5[3]), .A2(sram_raddr_a5[2]), .A3(
        sram_raddr_a5[1]), .A4(sram_raddr_a5[0]), .Y(n1694) );
  AO221X1_HVT U1860 ( .A1(n278), .A2(n411), .A3(n278), .A4(n1688), .A5(n1694), 
        .Y(n1813) );
  OA22X1_HVT U1861 ( .A1(n1689), .A2(n370), .A3(n171), .A4(n1813), .Y(n1692)
         );
  NAND3X0_HVT U1862 ( .A1(n1708), .A2(n1722), .A3(n370), .Y(n1691) );
  NAND4X0_HVT U1863 ( .A1(sram_raddr_a8[1]), .A2(sram_raddr_a8[0]), .A3(
        sram_raddr_a8[2]), .A4(sram_raddr_a8[3]), .Y(n1695) );
  OA21X1_HVT U1864 ( .A1(n1690), .A2(sram_raddr_a8[3]), .A3(n1695), .Y(n1951)
         );
  NAND2X0_HVT U1865 ( .A1(n168), .A2(n1951), .Y(n1815) );
  NAND3X0_HVT U1866 ( .A1(n1692), .A2(n1691), .A3(n1815), .Y(
        n_sram_raddr_a2[3]) );
  OA221X1_HVT U1867 ( .A1(n1693), .A2(sram_raddr_a2[3]), .A3(n1693), .A4(n1708), .A5(n1946), .Y(n1699) );
  NAND2X0_HVT U1868 ( .A1(sram_raddr_a5[4]), .A2(n1694), .Y(n1700) );
  OA22X1_HVT U1869 ( .A1(n1699), .A2(n366), .A3(n171), .A4(n1817), .Y(n1697)
         );
  NAND4X0_HVT U1870 ( .A1(sram_raddr_a2[3]), .A2(n1708), .A3(n1722), .A4(n366), 
        .Y(n1698) );
  NAND2X0_HVT U1871 ( .A1(n1696), .A2(sram_raddr_a8[4]), .Y(n1702) );
  OA21X1_HVT U1872 ( .A1(n1696), .A2(sram_raddr_a8[4]), .A3(n1702), .Y(n1956)
         );
  NAND2X0_HVT U1873 ( .A1(n521), .A2(n1956), .Y(n1819) );
  NAND3X0_HVT U1874 ( .A1(n1697), .A2(n1698), .A3(n1819), .Y(
        n_sram_raddr_a2[4]) );
  AND2X1_HVT U1875 ( .A1(n1699), .A2(n1698), .Y(n1706) );
  NOR2X0_HVT U1876 ( .A1(n350), .A2(n1700), .Y(n1707) );
  AO21X1_HVT U1877 ( .A1(n350), .A2(n1700), .A3(n1707), .Y(n1821) );
  OA22X1_HVT U1878 ( .A1(n1706), .A2(n385), .A3(n171), .A4(n1821), .Y(n1704)
         );
  AND3X1_HVT U1879 ( .A1(sram_raddr_a2[4]), .A2(sram_raddr_a2[3]), .A3(n1708), 
        .Y(n1701) );
  NAND3X0_HVT U1880 ( .A1(n1701), .A2(n1722), .A3(n385), .Y(n1705) );
  NAND2X0_HVT U1881 ( .A1(n1703), .A2(sram_raddr_a8[5]), .Y(n1709) );
  OA21X1_HVT U1882 ( .A1(n1703), .A2(sram_raddr_a8[5]), .A3(n1709), .Y(n1962)
         );
  NAND2X0_HVT U1883 ( .A1(n1839), .A2(n1962), .Y(n1824) );
  NAND3X0_HVT U1884 ( .A1(n1704), .A2(n1705), .A3(n1824), .Y(
        n_sram_raddr_a2[5]) );
  AND2X1_HVT U1885 ( .A1(n1706), .A2(n1705), .Y(n1713) );
  NAND2X0_HVT U1886 ( .A1(sram_raddr_a5[6]), .A2(n1707), .Y(n1714) );
  OA22X1_HVT U1887 ( .A1(n1713), .A2(n378), .A3(n189), .A4(n1826), .Y(n1711)
         );
  AND4X1_HVT U1888 ( .A1(sram_raddr_a2[5]), .A2(sram_raddr_a2[4]), .A3(
        sram_raddr_a2[3]), .A4(n1708), .Y(n1717) );
  NAND3X0_HVT U1889 ( .A1(n1717), .A2(n1722), .A3(n378), .Y(n1712) );
  NAND2X0_HVT U1890 ( .A1(n1710), .A2(sram_raddr_a8[6]), .Y(n1715) );
  OA21X1_HVT U1891 ( .A1(n1710), .A2(sram_raddr_a8[6]), .A3(n1715), .Y(n1967)
         );
  NAND2X0_HVT U1892 ( .A1(n521), .A2(n1967), .Y(n1828) );
  NAND3X0_HVT U1893 ( .A1(n1711), .A2(n1712), .A3(n1828), .Y(
        n_sram_raddr_a2[6]) );
  AND2X1_HVT U1894 ( .A1(n1713), .A2(n1712), .Y(n1721) );
  AO21X1_HVT U1895 ( .A1(n352), .A2(n1714), .A3(n1726), .Y(n1830) );
  OA22X1_HVT U1896 ( .A1(n1721), .A2(n356), .A3(n171), .A4(n1830), .Y(n1719)
         );
  NAND2X0_HVT U1897 ( .A1(n1716), .A2(sram_raddr_a8[7]), .Y(n1724) );
  OA21X1_HVT U1898 ( .A1(n1716), .A2(sram_raddr_a8[7]), .A3(n1724), .Y(n1973)
         );
  NAND2X0_HVT U1899 ( .A1(n168), .A2(n1973), .Y(n1835) );
  AND2X1_HVT U1900 ( .A1(sram_raddr_a2[6]), .A2(n1717), .Y(n1723) );
  NAND3X0_HVT U1901 ( .A1(n1723), .A2(n356), .A3(n1722), .Y(n1718) );
  NAND3X0_HVT U1902 ( .A1(n1719), .A2(n1835), .A3(n1718), .Y(
        n_sram_raddr_a2[7]) );
  NAND2X0_HVT U1903 ( .A1(n356), .A2(n1722), .Y(n1720) );
  NAND2X0_HVT U1904 ( .A1(n1721), .A2(n1720), .Y(n1734) );
  AND3X1_HVT U1905 ( .A1(sram_raddr_a2[7]), .A2(n1723), .A3(n1722), .Y(n1732)
         );
  NAND2X0_HVT U1906 ( .A1(n1725), .A2(sram_raddr_a8[8]), .Y(n1728) );
  OA21X1_HVT U1907 ( .A1(n1725), .A2(sram_raddr_a8[8]), .A3(n1728), .Y(n1981)
         );
  NAND2X0_HVT U1908 ( .A1(sram_raddr_a5[8]), .A2(n1726), .Y(n1730) );
  OA21X1_HVT U1909 ( .A1(sram_raddr_a5[8]), .A2(n1726), .A3(n1730), .Y(n1840)
         );
  AO22X1_HVT U1910 ( .A1(n521), .A2(n1981), .A3(n1975), .A4(n1840), .Y(n1727)
         );
  AO221X1_HVT U1911 ( .A1(sram_raddr_a2[8]), .A2(n1734), .A3(n435), .A4(n1732), 
        .A5(n1727), .Y(n_sram_raddr_a2[8]) );
  HADDX1_HVT U1912 ( .A0(sram_raddr_a8[9]), .B0(n1729), .SO(n1989) );
  AND2X1_HVT U1913 ( .A1(n521), .A2(n1989), .Y(n1847) );
  HADDX1_HVT U1914 ( .A0(sram_raddr_a5[9]), .B0(n1731), .SO(n1845) );
  HADDX1_HVT U1915 ( .A0(sram_raddr_a2[9]), .B0(sram_raddr_a2[8]), .SO(n1733)
         );
  NAND2X0_HVT U1916 ( .A1(n189), .A2(n1850), .Y(n1770) );
  AO22X1_HVT U1917 ( .A1(n521), .A2(n295), .A3(n1897), .A4(sram_raddr_a0[0]), 
        .Y(n1735) );
  AO221X1_HVT U1918 ( .A1(sram_raddr_a3[0]), .A2(n1888), .A3(n418), .A4(n1770), 
        .A5(n1735), .Y(n_sram_raddr_a3[0]) );
  OA21X1_HVT U1919 ( .A1(n297), .A2(n216), .A3(n1736), .Y(n1849) );
  AOI22X1_HVT U1920 ( .A1(n1737), .A2(n1770), .A3(sram_raddr_a3[1]), .A4(n1888), .Y(n1738) );
  NAND2X0_HVT U1921 ( .A1(n1849), .A2(n1738), .Y(n_sram_raddr_a3[1]) );
  OA22X1_HVT U1922 ( .A1(n1760), .A2(n245), .A3(n1759), .A4(n1740), .Y(n1742)
         );
  AO221X1_HVT U1923 ( .A1(sram_raddr_a0[3]), .A2(n248), .A3(n237), .A4(
        sram_raddr_a0[2]), .A5(n216), .Y(n1855) );
  NAND3X0_HVT U1924 ( .A1(n1742), .A2(n1741), .A3(n1855), .Y(
        n_sram_raddr_a3[3]) );
  NAND3X0_HVT U1925 ( .A1(n367), .A2(n237), .A3(n248), .Y(n1749) );
  NAND2X0_HVT U1926 ( .A1(n237), .A2(n248), .Y(n1743) );
  NAND2X0_HVT U1927 ( .A1(sram_raddr_a0[4]), .A2(n1743), .Y(n1745) );
  OA221X1_HVT U1928 ( .A1(n172), .A2(n1749), .A3(n216), .A4(n1745), .A5(n1744), 
        .Y(n1862) );
  OA22X1_HVT U1929 ( .A1(n1760), .A2(n279), .A3(n1759), .A4(n1746), .Y(n1747)
         );
  NAND2X0_HVT U1930 ( .A1(n1862), .A2(n1747), .Y(n_sram_raddr_a3[4]) );
  AOI22X1_HVT U1931 ( .A1(n1748), .A2(n1770), .A3(sram_raddr_a3[5]), .A4(n1888), .Y(n1752) );
  AO221X1_HVT U1932 ( .A1(sram_raddr_a0[5]), .A2(n1750), .A3(n291), .A4(n1749), 
        .A5(n172), .Y(n1866) );
  NAND3X0_HVT U1933 ( .A1(n1752), .A2(n1751), .A3(n1866), .Y(
        n_sram_raddr_a3[5]) );
  NAND4X0_HVT U1934 ( .A1(n291), .A2(n367), .A3(n237), .A4(n248), .Y(n1753) );
  OR2X1_HVT U1935 ( .A1(n1753), .A2(sram_raddr_a0[6]), .Y(n1761) );
  NAND2X0_HVT U1936 ( .A1(sram_raddr_a0[6]), .A2(n1753), .Y(n1755) );
  OA221X1_HVT U1937 ( .A1(n172), .A2(n1761), .A3(n216), .A4(n1755), .A5(n1754), 
        .Y(n1873) );
  OA22X1_HVT U1938 ( .A1(n1760), .A2(n349), .A3(n1759), .A4(n1756), .Y(n1757)
         );
  NAND2X0_HVT U1939 ( .A1(n1873), .A2(n1757), .Y(n_sram_raddr_a3[6]) );
  OA22X1_HVT U1940 ( .A1(n1760), .A2(n383), .A3(n1759), .A4(n1758), .Y(n1764)
         );
  NAND2X0_HVT U1941 ( .A1(n1762), .A2(n355), .Y(n1765) );
  AO221X1_HVT U1942 ( .A1(n1765), .A2(n1762), .A3(n1765), .A4(n355), .A5(n172), 
        .Y(n1878) );
  NAND3X0_HVT U1943 ( .A1(n1764), .A2(n1763), .A3(n1878), .Y(
        n_sram_raddr_a3[7]) );
  OA221X1_HVT U1944 ( .A1(sram_raddr_a0[8]), .A2(n1767), .A3(n402), .A4(n1765), 
        .A5(n1897), .Y(n1884) );
  NAND2X0_HVT U1945 ( .A1(n1767), .A2(n402), .Y(n1768) );
  OA221X1_HVT U1946 ( .A1(sram_raddr_a0[9]), .A2(n1769), .A3(n444), .A4(n1768), 
        .A5(n1897), .Y(n1890) );
  AO22X1_HVT U1947 ( .A1(n1771), .A2(n1770), .A3(sram_raddr_a3[9]), .A4(n1888), 
        .Y(n1772) );
  OR3X1_HVT U1948 ( .A1(n1773), .A2(n1890), .A3(n1772), .Y(n_sram_raddr_a3[9])
         );
  NAND2X0_HVT U1949 ( .A1(n1914), .A2(n171), .Y(n1804) );
  AO22X1_HVT U1950 ( .A1(n1839), .A2(n289), .A3(n1897), .A4(sram_raddr_a1[0]), 
        .Y(n1774) );
  AO221X1_HVT U1951 ( .A1(sram_raddr_a4[0]), .A2(n1935), .A3(n396), .A4(n1804), 
        .A5(n1774), .Y(n_sram_raddr_a4[0]) );
  OA22X1_HVT U1952 ( .A1(n1795), .A2(n1775), .A3(n1893), .A4(n298), .Y(n1777)
         );
  NAND2X0_HVT U1953 ( .A1(n1897), .A2(sram_raddr_a1[1]), .Y(n1894) );
  NAND3X0_HVT U1954 ( .A1(n1777), .A2(n1776), .A3(n1894), .Y(
        n_sram_raddr_a4[1]) );
  AOI22X1_HVT U1955 ( .A1(n1779), .A2(n1804), .A3(sram_raddr_a4[3]), .A4(n1935), .Y(n1781) );
  AO221X1_HVT U1956 ( .A1(sram_raddr_a1[2]), .A2(n236), .A3(n247), .A4(
        sram_raddr_a1[3]), .A5(n172), .Y(n1901) );
  NAND3X0_HVT U1957 ( .A1(n1781), .A2(n1780), .A3(n1901), .Y(
        n_sram_raddr_a4[3]) );
  OA22X1_HVT U1958 ( .A1(n1893), .A2(n246), .A3(n1795), .A4(n1782), .Y(n1786)
         );
  NAND2X0_HVT U1959 ( .A1(n247), .A2(n236), .Y(n1783) );
  AO221X1_HVT U1960 ( .A1(sram_raddr_a1[4]), .A2(n1784), .A3(n282), .A4(n1783), 
        .A5(n216), .Y(n1907) );
  NAND3X0_HVT U1961 ( .A1(n1786), .A2(n1785), .A3(n1907), .Y(
        n_sram_raddr_a4[4]) );
  OA22X1_HVT U1962 ( .A1(n1893), .A2(n404), .A3(n1795), .A4(n1787), .Y(n1790)
         );
  NAND4X0_HVT U1963 ( .A1(n380), .A2(n282), .A3(n247), .A4(n236), .Y(n1791) );
  AND3X1_HVT U1964 ( .A1(n282), .A2(n247), .A3(n236), .Y(n1788) );
  AO221X1_HVT U1965 ( .A1(n1791), .A2(n1788), .A3(n1791), .A4(n380), .A5(n172), 
        .Y(n1912) );
  NAND3X0_HVT U1966 ( .A1(n1790), .A2(n1789), .A3(n1912), .Y(
        n_sram_raddr_a4[5]) );
  OR2X1_HVT U1967 ( .A1(n1791), .A2(sram_raddr_a1[6]), .Y(n1797) );
  NAND2X0_HVT U1968 ( .A1(sram_raddr_a1[6]), .A2(n1791), .Y(n1793) );
  OA221X1_HVT U1969 ( .A1(n216), .A2(n1797), .A3(n216), .A4(n1793), .A5(n1792), 
        .Y(n1920) );
  OA22X1_HVT U1970 ( .A1(n1893), .A2(n353), .A3(n1795), .A4(n1794), .Y(n1796)
         );
  NAND2X0_HVT U1971 ( .A1(n1920), .A2(n1796), .Y(n_sram_raddr_a4[6]) );
  OR2X1_HVT U1972 ( .A1(n1797), .A2(sram_raddr_a1[7]), .Y(n1799) );
  OA221X1_HVT U1973 ( .A1(n1801), .A2(sram_raddr_a1[7]), .A3(n1801), .A4(n1797), .A5(n1897), .Y(n1924) );
  OA221X1_HVT U1974 ( .A1(sram_raddr_a1[8]), .A2(n1801), .A3(n403), .A4(n1799), 
        .A5(n1897), .Y(n1929) );
  NAND2X0_HVT U1975 ( .A1(n1801), .A2(n403), .Y(n1802) );
  OA221X1_HVT U1976 ( .A1(sram_raddr_a1[9]), .A2(n1803), .A3(n445), .A4(n1802), 
        .A5(n1897), .Y(n1936) );
  AO22X1_HVT U1977 ( .A1(n1805), .A2(n1804), .A3(sram_raddr_a4[9]), .A4(n1935), 
        .Y(n1806) );
  OR3X1_HVT U1978 ( .A1(n1807), .A2(n1936), .A3(n1806), .Y(n_sram_raddr_a4[9])
         );
  NAND2X0_HVT U1979 ( .A1(n171), .A2(n1942), .Y(n1844) );
  AO22X1_HVT U1980 ( .A1(n521), .A2(n288), .A3(n1897), .A4(n427), .Y(n1937) );
  AO221X1_HVT U1981 ( .A1(sram_raddr_a5[0]), .A2(n1990), .A3(n394), .A4(n1844), 
        .A5(n1937), .Y(n_sram_raddr_a5[0]) );
  AO22X1_HVT U1982 ( .A1(n1982), .A2(n1808), .A3(sram_raddr_a5[1]), .A4(n1990), 
        .Y(n1809) );
  OR2X1_HVT U1983 ( .A1(n1941), .A2(n1809), .Y(n_sram_raddr_a5[1]) );
  OA22X1_HVT U1984 ( .A1(n1946), .A2(n411), .A3(n1942), .A4(n1947), .Y(n1811)
         );
  NAND2X0_HVT U1985 ( .A1(n1897), .A2(n1810), .Y(n1949) );
  NAND3X0_HVT U1986 ( .A1(n1812), .A2(n1811), .A3(n1949), .Y(
        n_sram_raddr_a5[2]) );
  OA22X1_HVT U1987 ( .A1(n1831), .A2(n1813), .A3(n1946), .A4(n278), .Y(n1816)
         );
  NAND2X0_HVT U1988 ( .A1(n1814), .A2(n370), .Y(n1818) );
  AO221X1_HVT U1989 ( .A1(n1818), .A2(n1814), .A3(n1818), .A4(n370), .A5(n172), 
        .Y(n1954) );
  NAND3X0_HVT U1990 ( .A1(n1816), .A2(n1815), .A3(n1954), .Y(
        n_sram_raddr_a5[3]) );
  OA22X1_HVT U1991 ( .A1(n1946), .A2(n412), .A3(n1831), .A4(n1817), .Y(n1820)
         );
  AO221X1_HVT U1992 ( .A1(sram_raddr_a2[4]), .A2(n1822), .A3(n366), .A4(n1818), 
        .A5(n216), .Y(n1960) );
  NAND3X0_HVT U1993 ( .A1(n1820), .A2(n1819), .A3(n1960), .Y(
        n_sram_raddr_a5[4]) );
  OA22X1_HVT U1994 ( .A1(n1946), .A2(n350), .A3(n1831), .A4(n1821), .Y(n1825)
         );
  AND2X1_HVT U1995 ( .A1(n1822), .A2(n366), .Y(n1823) );
  NAND2X0_HVT U1996 ( .A1(n1823), .A2(n385), .Y(n1827) );
  AO221X1_HVT U1997 ( .A1(n1827), .A2(n1823), .A3(n1827), .A4(n385), .A5(n216), 
        .Y(n1965) );
  NAND3X0_HVT U1998 ( .A1(n1825), .A2(n1824), .A3(n1965), .Y(
        n_sram_raddr_a5[5]) );
  OA22X1_HVT U1999 ( .A1(n1946), .A2(n413), .A3(n1831), .A4(n1826), .Y(n1829)
         );
  AO221X1_HVT U2000 ( .A1(sram_raddr_a2[6]), .A2(n1832), .A3(n378), .A4(n1827), 
        .A5(n172), .Y(n1971) );
  NAND3X0_HVT U2001 ( .A1(n1829), .A2(n1828), .A3(n1971), .Y(
        n_sram_raddr_a5[6]) );
  OA22X1_HVT U2002 ( .A1(n1946), .A2(n352), .A3(n1831), .A4(n1830), .Y(n1836)
         );
  AND2X1_HVT U2003 ( .A1(n1832), .A2(n378), .Y(n1834) );
  NAND2X0_HVT U2004 ( .A1(n1834), .A2(n356), .Y(n1837) );
  AO221X1_HVT U2005 ( .A1(n1837), .A2(n1834), .A3(n1837), .A4(n356), .A5(n172), 
        .Y(n1978) );
  NAND3X0_HVT U2006 ( .A1(n1836), .A2(n1835), .A3(n1978), .Y(
        n_sram_raddr_a5[7]) );
  OR2X1_HVT U2007 ( .A1(n1837), .A2(sram_raddr_a2[8]), .Y(n1842) );
  AO21X1_HVT U2008 ( .A1(sram_raddr_a2[8]), .A2(n1837), .A3(n1843), .Y(n1838)
         );
  AO22X1_HVT U2009 ( .A1(n521), .A2(n1981), .A3(n1897), .A4(n1838), .Y(n1984)
         );
  AO22X1_HVT U2010 ( .A1(n1840), .A2(n1844), .A3(sram_raddr_a5[8]), .A4(n1990), 
        .Y(n1841) );
  OR2X1_HVT U2011 ( .A1(n1984), .A2(n1841), .Y(n_sram_raddr_a5[8]) );
  OA221X1_HVT U2012 ( .A1(sram_raddr_a2[9]), .A2(n1843), .A3(n446), .A4(n1842), 
        .A5(n1897), .Y(n1993) );
  AO22X1_HVT U2013 ( .A1(n1845), .A2(n1844), .A3(sram_raddr_a5[9]), .A4(n1990), 
        .Y(n1846) );
  OR3X1_HVT U2014 ( .A1(n1847), .A2(n1993), .A3(n1846), .Y(n_sram_raddr_a5[9])
         );
  NAND2X0_HVT U2015 ( .A1(n1943), .A2(n1850), .Y(n1886) );
  AO22X1_HVT U2016 ( .A1(n1897), .A2(sram_raddr_a0[0]), .A3(n1975), .A4(
        sram_raddr_a3[0]), .Y(n1848) );
  AO221X1_HVT U2017 ( .A1(sram_raddr_a6[0]), .A2(n1888), .A3(n295), .A4(n1886), 
        .A5(n1848), .Y(n_sram_raddr_a6[0]) );
  AOI22X1_HVT U2018 ( .A1(sram_raddr_a6[3]), .A2(n1888), .A3(n1853), .A4(n1886), .Y(n1856) );
  AO221X1_HVT U2019 ( .A1(sram_raddr_a3[2]), .A2(n245), .A3(n234), .A4(
        sram_raddr_a3[3]), .A5(n189), .Y(n1854) );
  NAND3X0_HVT U2020 ( .A1(n1856), .A2(n1855), .A3(n1854), .Y(
        n_sram_raddr_a6[3]) );
  AOI22X1_HVT U2021 ( .A1(sram_raddr_a6[4]), .A2(n1888), .A3(n1869), .A4(n1857), .Y(n1861) );
  NAND2X0_HVT U2022 ( .A1(n234), .A2(n245), .Y(n1858) );
  AO221X1_HVT U2023 ( .A1(sram_raddr_a3[4]), .A2(n1859), .A3(n279), .A4(n1858), 
        .A5(n189), .Y(n1860) );
  NAND3X0_HVT U2024 ( .A1(n1862), .A2(n1861), .A3(n1860), .Y(
        n_sram_raddr_a6[4]) );
  AOI22X1_HVT U2025 ( .A1(sram_raddr_a6[5]), .A2(n1888), .A3(n1863), .A4(n1886), .Y(n1867) );
  NAND4X0_HVT U2026 ( .A1(n428), .A2(n279), .A3(n234), .A4(n245), .Y(n1870) );
  AND3X1_HVT U2027 ( .A1(n279), .A2(n234), .A3(n245), .Y(n1864) );
  AO221X1_HVT U2028 ( .A1(n1870), .A2(n1864), .A3(n1870), .A4(n428), .A5(n171), 
        .Y(n1865) );
  NAND3X0_HVT U2029 ( .A1(n1867), .A2(n1866), .A3(n1865), .Y(
        n_sram_raddr_a6[5]) );
  AOI22X1_HVT U2030 ( .A1(sram_raddr_a6[6]), .A2(n1888), .A3(n1869), .A4(n1868), .Y(n1872) );
  AO221X1_HVT U2031 ( .A1(sram_raddr_a3[6]), .A2(n1875), .A3(n349), .A4(n1870), 
        .A5(n189), .Y(n1871) );
  NAND3X0_HVT U2032 ( .A1(n1873), .A2(n1872), .A3(n1871), .Y(
        n_sram_raddr_a6[6]) );
  AOI22X1_HVT U2033 ( .A1(sram_raddr_a6[7]), .A2(n1888), .A3(n1874), .A4(n1886), .Y(n1879) );
  AND2X1_HVT U2034 ( .A1(n1875), .A2(n349), .Y(n1876) );
  NAND2X0_HVT U2035 ( .A1(n1876), .A2(n383), .Y(n1880) );
  AO221X1_HVT U2036 ( .A1(n1880), .A2(n1876), .A3(n1880), .A4(n383), .A5(n189), 
        .Y(n1877) );
  NAND3X0_HVT U2037 ( .A1(n1879), .A2(n1878), .A3(n1877), .Y(
        n_sram_raddr_a6[7]) );
  OA221X1_HVT U2038 ( .A1(n1885), .A2(sram_raddr_a3[8]), .A3(n1885), .A4(n1880), .A5(n170), .Y(n1883) );
  AO22X1_HVT U2039 ( .A1(sram_raddr_a6[8]), .A2(n1888), .A3(n1881), .A4(n1886), 
        .Y(n1882) );
  OR3X1_HVT U2040 ( .A1(n1884), .A2(n1883), .A3(n1882), .Y(n_sram_raddr_a6[8])
         );
  HADDX1_HVT U2041 ( .A0(sram_raddr_a3[9]), .B0(n1885), .SO(n1889) );
  NAND2X0_HVT U2042 ( .A1(n1943), .A2(n1914), .Y(n1932) );
  AO22X1_HVT U2043 ( .A1(n1897), .A2(sram_raddr_a1[0]), .A3(n1975), .A4(
        sram_raddr_a4[0]), .Y(n1891) );
  AO221X1_HVT U2044 ( .A1(sram_raddr_a7[0]), .A2(n1935), .A3(n289), .A4(n1932), 
        .A5(n1891), .Y(n_sram_raddr_a7[0]) );
  NAND2X0_HVT U2045 ( .A1(n1892), .A2(n1932), .Y(n1896) );
  OA22X1_HVT U2046 ( .A1(n1893), .A2(n429), .A3(n171), .A4(n298), .Y(n1895) );
  NAND3X0_HVT U2047 ( .A1(n1896), .A2(n1895), .A3(n1894), .Y(
        n_sram_raddr_a7[1]) );
  AOI22X1_HVT U2048 ( .A1(sram_raddr_a7[3]), .A2(n1935), .A3(n1899), .A4(n1932), .Y(n1902) );
  AO221X1_HVT U2049 ( .A1(sram_raddr_a4[2]), .A2(n290), .A3(n235), .A4(
        sram_raddr_a4[3]), .A5(n171), .Y(n1900) );
  NAND3X0_HVT U2050 ( .A1(n1902), .A2(n1901), .A3(n1900), .Y(
        n_sram_raddr_a7[3]) );
  AOI22X1_HVT U2051 ( .A1(sram_raddr_a7[4]), .A2(n1935), .A3(n1903), .A4(n1932), .Y(n1908) );
  NAND2X0_HVT U2052 ( .A1(n235), .A2(n290), .Y(n1904) );
  AO221X1_HVT U2053 ( .A1(sram_raddr_a4[4]), .A2(n1905), .A3(n246), .A4(n1904), 
        .A5(n189), .Y(n1906) );
  NAND3X0_HVT U2054 ( .A1(n1908), .A2(n1907), .A3(n1906), .Y(
        n_sram_raddr_a7[4]) );
  AOI22X1_HVT U2055 ( .A1(sram_raddr_a7[5]), .A2(n1935), .A3(n1909), .A4(n1932), .Y(n1913) );
  NAND4X0_HVT U2056 ( .A1(n404), .A2(n246), .A3(n235), .A4(n290), .Y(n1917) );
  AND3X1_HVT U2057 ( .A1(n246), .A2(n235), .A3(n290), .Y(n1910) );
  AO221X1_HVT U2058 ( .A1(n1917), .A2(n1910), .A3(n1917), .A4(n404), .A5(n189), 
        .Y(n1911) );
  NAND3X0_HVT U2059 ( .A1(n1913), .A2(n1912), .A3(n1911), .Y(
        n_sram_raddr_a7[5]) );
  AOI22X1_HVT U2060 ( .A1(sram_raddr_a7[6]), .A2(n1935), .A3(n1916), .A4(n1915), .Y(n1919) );
  AO221X1_HVT U2061 ( .A1(sram_raddr_a4[6]), .A2(n1921), .A3(n353), .A4(n1917), 
        .A5(n171), .Y(n1918) );
  NAND3X0_HVT U2062 ( .A1(n1920), .A2(n1919), .A3(n1918), .Y(
        n_sram_raddr_a7[6]) );
  NAND2X0_HVT U2063 ( .A1(n1921), .A2(n353), .Y(n1922) );
  OR2X1_HVT U2064 ( .A1(n1922), .A2(sram_raddr_a4[7]), .Y(n1925) );
  OA221X1_HVT U2065 ( .A1(n1930), .A2(sram_raddr_a4[8]), .A3(n1930), .A4(n1925), .A5(n170), .Y(n1928) );
  AO22X1_HVT U2066 ( .A1(sram_raddr_a7[8]), .A2(n1935), .A3(n1926), .A4(n1932), 
        .Y(n1927) );
  OR3X1_HVT U2067 ( .A1(n1929), .A2(n1928), .A3(n1927), .Y(n_sram_raddr_a7[8])
         );
  HADDX1_HVT U2068 ( .A0(sram_raddr_a4[9]), .B0(n1930), .SO(n1931) );
  AO221X1_HVT U2069 ( .A1(sram_raddr_a8[0]), .A2(n1990), .A3(n288), .A4(n1982), 
        .A5(n1937), .Y(n1938) );
  AO21X1_HVT U2070 ( .A1(n170), .A2(n394), .A3(n1938), .Y(n_sram_raddr_a8[0])
         );
  AO22X1_HVT U2071 ( .A1(sram_raddr_a8[1]), .A2(n1990), .A3(n1982), .A4(n1939), 
        .Y(n1940) );
  OR2X1_HVT U2072 ( .A1(n1941), .A2(n1940), .Y(n_sram_raddr_a8[1]) );
  NAND2X0_HVT U2073 ( .A1(n1943), .A2(n1942), .Y(n1988) );
  OA22X1_HVT U2074 ( .A1(n1946), .A2(n438), .A3(n1945), .A4(n1944), .Y(n1950)
         );
  NAND2X0_HVT U2075 ( .A1(n170), .A2(n1947), .Y(n1948) );
  NAND3X0_HVT U2076 ( .A1(n1950), .A2(n1949), .A3(n1948), .Y(
        n_sram_raddr_a8[2]) );
  AOI22X1_HVT U2077 ( .A1(sram_raddr_a8[3]), .A2(n1990), .A3(n1951), .A4(n1988), .Y(n1955) );
  AO221X1_HVT U2078 ( .A1(sram_raddr_a5[3]), .A2(n1957), .A3(n278), .A4(n1952), 
        .A5(n171), .Y(n1953) );
  NAND3X0_HVT U2079 ( .A1(n1955), .A2(n1954), .A3(n1953), .Y(
        n_sram_raddr_a8[3]) );
  AOI22X1_HVT U2080 ( .A1(sram_raddr_a8[4]), .A2(n1990), .A3(n1956), .A4(n1988), .Y(n1961) );
  AND2X1_HVT U2081 ( .A1(n1957), .A2(n278), .Y(n1958) );
  NAND2X0_HVT U2082 ( .A1(n1958), .A2(n412), .Y(n1963) );
  AO221X1_HVT U2083 ( .A1(n1963), .A2(n1958), .A3(n1963), .A4(n412), .A5(n171), 
        .Y(n1959) );
  NAND3X0_HVT U2084 ( .A1(n1961), .A2(n1960), .A3(n1959), .Y(
        n_sram_raddr_a8[4]) );
  AOI22X1_HVT U2085 ( .A1(sram_raddr_a8[5]), .A2(n1990), .A3(n1962), .A4(n1988), .Y(n1966) );
  AO221X1_HVT U2086 ( .A1(sram_raddr_a5[5]), .A2(n1968), .A3(n350), .A4(n1963), 
        .A5(n171), .Y(n1964) );
  NAND3X0_HVT U2087 ( .A1(n1966), .A2(n1965), .A3(n1964), .Y(
        n_sram_raddr_a8[5]) );
  AOI22X1_HVT U2088 ( .A1(sram_raddr_a8[6]), .A2(n1990), .A3(n1967), .A4(n1988), .Y(n1972) );
  AND2X1_HVT U2089 ( .A1(n1968), .A2(n350), .Y(n1969) );
  NAND2X0_HVT U2090 ( .A1(n1969), .A2(n413), .Y(n1974) );
  AO221X1_HVT U2091 ( .A1(n1974), .A2(n1969), .A3(n1974), .A4(n413), .A5(n189), 
        .Y(n1970) );
  NAND3X0_HVT U2092 ( .A1(n1972), .A2(n1971), .A3(n1970), .Y(
        n_sram_raddr_a8[6]) );
  AOI22X1_HVT U2093 ( .A1(sram_raddr_a8[7]), .A2(n1990), .A3(n1973), .A4(n1988), .Y(n1979) );
  NAND2X0_HVT U2094 ( .A1(n1976), .A2(n352), .Y(n1980) );
  AO221X1_HVT U2095 ( .A1(n1980), .A2(n1976), .A3(n1980), .A4(n352), .A5(n171), 
        .Y(n1977) );
  NAND3X0_HVT U2096 ( .A1(n1979), .A2(n1978), .A3(n1977), .Y(
        n_sram_raddr_a8[7]) );
  OR2X1_HVT U2097 ( .A1(n1980), .A2(sram_raddr_a5[8]), .Y(n1986) );
  OA221X1_HVT U2098 ( .A1(n1987), .A2(sram_raddr_a5[8]), .A3(n1987), .A4(n1980), .A5(n170), .Y(n1985) );
  AO22X1_HVT U2099 ( .A1(sram_raddr_a8[8]), .A2(n1990), .A3(n1982), .A4(n1981), 
        .Y(n1983) );
  OR3X1_HVT U2100 ( .A1(n1985), .A2(n1984), .A3(n1983), .Y(n_sram_raddr_a8[8])
         );
  OA221X1_HVT U2101 ( .A1(sram_raddr_a5[9]), .A2(n1987), .A3(n442), .A4(n1986), 
        .A5(n170), .Y(n1992) );
  AO22X1_HVT U2102 ( .A1(sram_raddr_a8[9]), .A2(n1990), .A3(n1989), .A4(n1988), 
        .Y(n1991) );
  OR3X1_HVT U2103 ( .A1(n1993), .A2(n1992), .A3(n1991), .Y(n_sram_raddr_a8[9])
         );
  AND2X1_HVT U2104 ( .A1(n1994), .A2(addr_row_sel_cnt[1]), .Y(n392) );
  OA221X1_HVT U2105 ( .A1(n2004), .A2(n1995), .A3(n2004), .A4(n2002), .A5(
        n2000), .Y(n371) );
  AO22X1_HVT U2106 ( .A1(n1999), .A2(n1998), .A3(n1997), .A4(n2002), .Y(n369)
         );
  OA221X1_HVT U2107 ( .A1(n2004), .A2(n2003), .A3(n2004), .A4(n2002), .A5(
        n2001), .Y(n368) );
endmodule


module data_reg ( clk, srstn, mode, box_sel, sram_rdata_a0, sram_rdata_a1, 
        sram_rdata_a2, sram_rdata_a3, sram_rdata_a4, sram_rdata_a5, 
        sram_rdata_a6, sram_rdata_a7, sram_rdata_a8, sram_rdata_b0, 
        sram_rdata_b1, sram_rdata_b2, sram_rdata_b3, sram_rdata_b4, 
        sram_rdata_b5, sram_rdata_b6, sram_rdata_b7, sram_rdata_b8, 
        sram_rdata_weight, conv1_weight, weight, src_window );
  input [1:0] mode;
  input [3:0] box_sel;
  input [31:0] sram_rdata_a0;
  input [31:0] sram_rdata_a1;
  input [31:0] sram_rdata_a2;
  input [31:0] sram_rdata_a3;
  input [31:0] sram_rdata_a4;
  input [31:0] sram_rdata_a5;
  input [31:0] sram_rdata_a6;
  input [31:0] sram_rdata_a7;
  input [31:0] sram_rdata_a8;
  input [31:0] sram_rdata_b0;
  input [31:0] sram_rdata_b1;
  input [31:0] sram_rdata_b2;
  input [31:0] sram_rdata_b3;
  input [31:0] sram_rdata_b4;
  input [31:0] sram_rdata_b5;
  input [31:0] sram_rdata_b6;
  input [31:0] sram_rdata_b7;
  input [31:0] sram_rdata_b8;
  input [99:0] sram_rdata_weight;
  output [99:0] conv1_weight;
  output [99:0] weight;
  output [287:0] src_window;
  input clk, srstn;
  wire   N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52,
         N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66,
         N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80,
         N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94,
         N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106,
         N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139,
         N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161,
         N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172,
         N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183,
         N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194,
         N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205,
         N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216,
         N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227,
         N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238,
         N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249,
         N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260,
         N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271,
         N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282,
         N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293,
         N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304,
         N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315,
         N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326,
         N346, n2, n3, n5, n6, n8, n9, n11, n12, n14, n15, n17, n18, n20, n21,
         n23, n24, n26, n27, n29, n30, n32, n33, n35, n36, n37, n3900, n4000,
         n4200, n4300, n4500, n4600, n4800, n4900, n5100, n5200, n5400, n5500,
         n5700, n5800, n6000, n6100, n6300, n6400, n6600, n6700, n6900, n7000,
         n7200, n7300, n7500, n7600, n7800, n7900, n8100, n8200, n8400, n8500,
         n8700, n8800, n9000, n9100, n9300, n9400, n9600, n9700, n9800, n9900,
         n10000, n10100, n10200, n10300, n10400, n10500, n10600, n10700,
         n10800, n10900, n11000, n11100, n11200, n11300, n11400, n11500,
         n11600, n11700, n11800, n11900, n12000, n12100, n12200, n12300,
         n12400, n12500, n12600, n12700, n12800, n12900, n13000, n13100,
         n13200, n13300, n13400, n13500, n13600, n13700, n13800, n13900,
         n14000, n14100, n14200, n14300, n14400, n14500, n14600, n14700,
         n14800, n14900, n15000, n15100, n15200, n15300, n15400, n15500,
         n15600, n15700, n15800, n15900, n16000, n16100, n16200, n16300,
         n16400, n16500, n16600, n1670, n1680, n1690, n1700, n1710, n1720,
         n1730, n1740, n1750, n1760, n1770, n1780, n1790, n1800, n1810, n1820,
         n1830, n1840, n1850, n1860, n1870, n1880, n1890, n1900, n1910, n1920,
         n1930, n1940, n1950, n1960, n1970, n1980, n1990, n2000, n2010, n2020,
         n2030, n2040, n2050, n2060, n2070, n2080, n2090, n2100, n2110, n2120,
         n2130, n2140, n2150, n2160, n2170, n2180, n2190, n2200, n2210, n2220,
         n2230, n2240, n2250, n2260, n2270, n2280, n2290, n2300, n2310, n2320,
         n2330, n2340, n2350, n2360, n2370, n2380, n2390, n2400, n2410, n2420,
         n2430, n2440, n2450, n2460, n2470, n2480, n2490, n2500, n2510, n2520,
         n2530, n2540, n2550, n2560, n2570, n2580, n2590, n2600, n2610, n2620,
         n2630, n2640, n2650, n2660, n2670, n2680, n2690, n2700, n2710, n2720,
         n2730, n2740, n2750, n2760, n2770, n2780, n2790, n2800, n2810, n2820,
         n2830, n2840, n2850, n2860, n2870, n2880, n2890, n2900, n2910, n2920,
         n2930, n2940, n2950, n2960, n2970, n2980, n2990, n3000, n3010, n3020,
         n3030, n3040, n3050, n3060, n3070, n3080, n3090, n3100, n3110, n3120,
         n3130, n3140, n3150, n3160, n3170, n3180, n3190, n3200, n3210, n3220,
         n3230, n3240, n3250, n3260, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n3460, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n3901, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n4001, n401, n402, n403, n404, n405, n406, n407, n408, n409, n4101,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n4201, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n4301, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n4401, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n4501, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n4601, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n4701, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n4801, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n4901, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n5001, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n5101, n511, n512, n513, n514, n515, n516, n517, n518, n519, n5201,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n5301, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n5401, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n5501, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n5601, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n5701, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n5801, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n5901, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n6001, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n6101, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n6201, n621, n622, n623, n624, n625, n626, n627, n628, n629, n6301,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n6401, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n6501, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n6601, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n6701, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n6801, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n6901, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n7001, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n7101, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n7201, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n7301, n731, n732, n733, n734, n735, n736, n737, n738, n739, n7401,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n7501, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n7601, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n7701, n771, n772, n773,
         n774, n775, n777, n778, n779, n7801, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n7901, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n8001, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n8101, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n8201, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n8301, n831, n832, n833, n834, n835, n836, n837, n838, n839, n8401,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n8501, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n8601, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n8701, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n8801, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n8901, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n9001, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n9101, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n9201, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n9301, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n9401, n941, n942, n943, n944, n945, n946, n947, n948, n949, n9501,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n9601, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n9701, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n9801, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n9901, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n10001, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n10101, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n10201, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n10301, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n10401, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n10501, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n10601, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n10701, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n10801, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n10901, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n11001, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n11101, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n11201, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n11301, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n11401, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n11501, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n11601, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n11701, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n11801, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n11901, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n12001, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n12101, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n12201, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n12301, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n12401, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n12501, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n12601, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n12701, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n12801, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n12901, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n13001, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n13101, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n13201, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n13301, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n13401, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n13501, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n13601, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n13701, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n13801, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n13901, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n14001, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n14101, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n14201, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n14301, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n14401, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n14501, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n14601, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n14701, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n14801, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n14901, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n15001, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n15101, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n15201, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n15301, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n15401, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n15501, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n15601, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n15701, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n15801, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n15901, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n16001, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n16101, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n16201, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n16301, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n16401, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n16501, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n16601, n1661, n1662, n1663, n1664
;
  wire   [287:0] n_src_aox;
  wire   [31:0] sram_rdata_0;
  wire   [31:0] sram_rdata_1;
  wire   [31:0] sram_rdata_2;
  wire   [31:0] sram_rdata_3;
  wire   [31:0] sram_rdata_4;
  wire   [31:0] sram_rdata_5;
  wire   [31:0] sram_rdata_6;
  wire   [31:0] sram_rdata_7;
  wire   [31:0] sram_rdata_8;

  DFFSSRX1_HVT src_aox_reg_0__7_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[287]), .CLK(clk), .Q(src_window[287]) );
  DFFSSRX1_HVT src_aox_reg_0__6_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[286]), .CLK(clk), .Q(src_window[286]) );
  DFFSSRX1_HVT src_aox_reg_0__5_ ( .D(1'b0), .SETB(n13000), .RSTB(
        n_src_aox[285]), .CLK(clk), .Q(src_window[285]) );
  DFFSSRX1_HVT src_aox_reg_0__4_ ( .D(1'b0), .SETB(n577), .RSTB(n_src_aox[284]), .CLK(clk), .Q(src_window[284]) );
  DFFSSRX1_HVT src_aox_reg_0__3_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[283]), .CLK(clk), .Q(src_window[283]) );
  DFFSSRX1_HVT src_aox_reg_0__2_ ( .D(1'b0), .SETB(n11400), .RSTB(
        n_src_aox[282]), .CLK(clk), .Q(src_window[282]) );
  DFFSSRX1_HVT src_aox_reg_0__1_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[281]), .CLK(clk), .Q(src_window[281]) );
  DFFSSRX1_HVT src_aox_reg_0__0_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[280]), .CLK(clk), .Q(src_window[280]) );
  DFFSSRX1_HVT src_aox_reg_1__7_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[279]), .CLK(clk), .Q(src_window[279]) );
  DFFSSRX1_HVT src_aox_reg_1__6_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[278]), .CLK(clk), .Q(src_window[278]) );
  DFFSSRX1_HVT src_aox_reg_1__5_ ( .D(1'b0), .SETB(n11400), .RSTB(
        n_src_aox[277]), .CLK(clk), .Q(src_window[277]) );
  DFFSSRX1_HVT src_aox_reg_1__4_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[276]), .CLK(clk), .Q(src_window[276]) );
  DFFSSRX1_HVT src_aox_reg_1__3_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[275]), .CLK(clk), .Q(src_window[275]) );
  DFFSSRX1_HVT src_aox_reg_1__2_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[274]), .CLK(clk), .Q(src_window[274]) );
  DFFSSRX1_HVT src_aox_reg_1__1_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[273]), .CLK(clk), .Q(src_window[273]) );
  DFFSSRX1_HVT src_aox_reg_1__0_ ( .D(1'b0), .SETB(n577), .RSTB(n_src_aox[272]), .CLK(clk), .Q(src_window[272]) );
  DFFSSRX1_HVT src_aox_reg_2__7_ ( .D(1'b0), .SETB(N346), .RSTB(n_src_aox[271]), .CLK(clk), .Q(src_window[271]) );
  DFFSSRX1_HVT src_aox_reg_2__6_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[270]), .CLK(clk), .Q(src_window[270]) );
  DFFSSRX1_HVT src_aox_reg_2__5_ ( .D(1'b0), .SETB(n577), .RSTB(n_src_aox[269]), .CLK(clk), .Q(src_window[269]) );
  DFFSSRX1_HVT src_aox_reg_2__4_ ( .D(1'b0), .SETB(n13000), .RSTB(
        n_src_aox[268]), .CLK(clk), .Q(src_window[268]) );
  DFFSSRX1_HVT src_aox_reg_2__3_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[267]), .CLK(clk), .Q(src_window[267]) );
  DFFSSRX1_HVT src_aox_reg_2__2_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[266]), .CLK(clk), .Q(src_window[266]) );
  DFFSSRX1_HVT src_aox_reg_2__1_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[265]), .CLK(clk), .Q(src_window[265]) );
  DFFSSRX1_HVT src_aox_reg_2__0_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[264]), .CLK(clk), .Q(src_window[264]) );
  DFFSSRX1_HVT src_aox_reg_3__7_ ( .D(1'b0), .SETB(n11400), .RSTB(
        n_src_aox[263]), .CLK(clk), .Q(src_window[263]) );
  DFFSSRX1_HVT src_aox_reg_3__6_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[262]), .CLK(clk), .Q(src_window[262]) );
  DFFSSRX1_HVT src_aox_reg_3__5_ ( .D(1'b0), .SETB(N346), .RSTB(n_src_aox[261]), .CLK(clk), .Q(src_window[261]) );
  DFFSSRX1_HVT src_aox_reg_3__4_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[260]), .CLK(clk), .Q(src_window[260]) );
  DFFSSRX1_HVT src_aox_reg_3__3_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[259]), .CLK(clk), .Q(src_window[259]) );
  DFFSSRX1_HVT src_aox_reg_3__2_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[258]), .CLK(clk), .Q(src_window[258]) );
  DFFSSRX1_HVT src_aox_reg_3__1_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[257]), .CLK(clk), .Q(src_window[257]) );
  DFFSSRX1_HVT src_aox_reg_3__0_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[256]), .CLK(clk), .Q(src_window[256]) );
  DFFSSRX1_HVT src_aox_reg_4__7_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[255]), .CLK(clk), .Q(src_window[255]) );
  DFFSSRX1_HVT src_aox_reg_4__6_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[254]), .CLK(clk), .Q(src_window[254]) );
  DFFSSRX1_HVT src_aox_reg_4__5_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[253]), .CLK(clk), .Q(src_window[253]) );
  DFFSSRX1_HVT src_aox_reg_4__4_ ( .D(1'b0), .SETB(n577), .RSTB(n_src_aox[252]), .CLK(clk), .Q(src_window[252]) );
  DFFSSRX1_HVT src_aox_reg_4__3_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[251]), .CLK(clk), .Q(src_window[251]) );
  DFFSSRX1_HVT src_aox_reg_4__2_ ( .D(1'b0), .SETB(n11400), .RSTB(
        n_src_aox[250]), .CLK(clk), .Q(src_window[250]) );
  DFFSSRX1_HVT src_aox_reg_4__1_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[249]), .CLK(clk), .Q(src_window[249]) );
  DFFSSRX1_HVT src_aox_reg_4__0_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[248]), .CLK(clk), .Q(src_window[248]) );
  DFFSSRX1_HVT src_aox_reg_5__7_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[247]), .CLK(clk), .Q(src_window[247]) );
  DFFSSRX1_HVT src_aox_reg_5__6_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[246]), .CLK(clk), .Q(src_window[246]) );
  DFFSSRX1_HVT src_aox_reg_5__5_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[245]), .CLK(clk), .Q(src_window[245]) );
  DFFSSRX1_HVT src_aox_reg_5__4_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[244]), .CLK(clk), .Q(src_window[244]) );
  DFFSSRX1_HVT src_aox_reg_5__3_ ( .D(1'b0), .SETB(n2600), .RSTB(
        n_src_aox[243]), .CLK(clk), .Q(src_window[243]) );
  DFFSSRX1_HVT src_aox_reg_5__2_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[242]), .CLK(clk), .Q(src_window[242]) );
  DFFSSRX1_HVT src_aox_reg_5__1_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[241]), .CLK(clk), .Q(src_window[241]) );
  DFFSSRX1_HVT src_aox_reg_5__0_ ( .D(1'b0), .SETB(n577), .RSTB(n_src_aox[240]), .CLK(clk), .Q(src_window[240]) );
  DFFSSRX1_HVT src_aox_reg_6__7_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[239]), .CLK(clk), .Q(src_window[239]) );
  DFFSSRX1_HVT src_aox_reg_6__6_ ( .D(1'b0), .SETB(N346), .RSTB(n_src_aox[238]), .CLK(clk), .Q(src_window[238]) );
  DFFSSRX1_HVT src_aox_reg_6__5_ ( .D(1'b0), .SETB(n577), .RSTB(n_src_aox[237]), .CLK(clk), .Q(src_window[237]) );
  DFFSSRX1_HVT src_aox_reg_6__4_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[236]), .CLK(clk), .Q(src_window[236]) );
  DFFSSRX1_HVT src_aox_reg_6__3_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[235]), .CLK(clk), .Q(src_window[235]) );
  DFFSSRX1_HVT src_aox_reg_6__2_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[234]), .CLK(clk), .Q(src_window[234]) );
  DFFSSRX1_HVT src_aox_reg_6__1_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[233]), .CLK(clk), .Q(src_window[233]) );
  DFFSSRX1_HVT src_aox_reg_6__0_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[232]), .CLK(clk), .Q(src_window[232]) );
  DFFSSRX1_HVT src_aox_reg_7__7_ ( .D(1'b0), .SETB(n11400), .RSTB(
        n_src_aox[231]), .CLK(clk), .Q(src_window[231]) );
  DFFSSRX1_HVT src_aox_reg_7__6_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[230]), .CLK(clk), .Q(src_window[230]) );
  DFFSSRX1_HVT src_aox_reg_7__5_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[229]), .CLK(clk), .Q(src_window[229]) );
  DFFSSRX1_HVT src_aox_reg_7__4_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[228]), .CLK(clk), .Q(src_window[228]) );
  DFFSSRX1_HVT src_aox_reg_7__3_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[227]), .CLK(clk), .Q(src_window[227]) );
  DFFSSRX1_HVT src_aox_reg_7__2_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[226]), .CLK(clk), .Q(src_window[226]) );
  DFFSSRX1_HVT src_aox_reg_7__1_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[225]), .CLK(clk), .Q(src_window[225]) );
  DFFSSRX1_HVT src_aox_reg_7__0_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[224]), .CLK(clk), .Q(src_window[224]) );
  DFFSSRX1_HVT src_aox_reg_8__7_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[223]), .CLK(clk), .Q(src_window[223]) );
  DFFSSRX1_HVT src_aox_reg_8__6_ ( .D(1'b0), .SETB(n13000), .RSTB(
        n_src_aox[222]), .CLK(clk), .Q(src_window[222]) );
  DFFSSRX1_HVT src_aox_reg_8__5_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[221]), .CLK(clk), .Q(src_window[221]) );
  DFFSSRX1_HVT src_aox_reg_8__4_ ( .D(1'b0), .SETB(n577), .RSTB(n_src_aox[220]), .CLK(clk), .Q(src_window[220]) );
  DFFSSRX1_HVT src_aox_reg_8__3_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[219]), .CLK(clk), .Q(src_window[219]) );
  DFFSSRX1_HVT src_aox_reg_8__2_ ( .D(1'b0), .SETB(n11400), .RSTB(
        n_src_aox[218]), .CLK(clk), .Q(src_window[218]) );
  DFFSSRX1_HVT src_aox_reg_8__1_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[217]), .CLK(clk), .Q(src_window[217]) );
  DFFSSRX1_HVT src_aox_reg_8__0_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[216]), .CLK(clk), .Q(src_window[216]) );
  DFFSSRX1_HVT src_aox_reg_9__7_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[215]), .CLK(clk), .Q(src_window[215]) );
  DFFSSRX1_HVT src_aox_reg_9__6_ ( .D(1'b0), .SETB(n13000), .RSTB(
        n_src_aox[214]), .CLK(clk), .Q(src_window[214]) );
  DFFSSRX1_HVT src_aox_reg_9__5_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[213]), .CLK(clk), .Q(src_window[213]) );
  DFFSSRX1_HVT src_aox_reg_9__4_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[212]), .CLK(clk), .Q(src_window[212]) );
  DFFSSRX1_HVT src_aox_reg_9__3_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[211]), .CLK(clk), .Q(src_window[211]) );
  DFFSSRX1_HVT src_aox_reg_9__2_ ( .D(1'b0), .SETB(n11400), .RSTB(
        n_src_aox[210]), .CLK(clk), .Q(src_window[210]) );
  DFFSSRX1_HVT src_aox_reg_9__1_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[209]), .CLK(clk), .Q(src_window[209]) );
  DFFSSRX1_HVT src_aox_reg_9__0_ ( .D(1'b0), .SETB(n577), .RSTB(n_src_aox[208]), .CLK(clk), .Q(src_window[208]) );
  DFFSSRX1_HVT src_aox_reg_10__7_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[207]), .CLK(clk), .Q(src_window[207]) );
  DFFSSRX1_HVT src_aox_reg_10__6_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[206]), .CLK(clk), .Q(src_window[206]) );
  DFFSSRX1_HVT src_aox_reg_10__5_ ( .D(1'b0), .SETB(n577), .RSTB(
        n_src_aox[205]), .CLK(clk), .Q(src_window[205]) );
  DFFSSRX1_HVT src_aox_reg_10__4_ ( .D(1'b0), .SETB(n11400), .RSTB(
        n_src_aox[204]), .CLK(clk), .Q(src_window[204]) );
  DFFSSRX1_HVT src_aox_reg_10__3_ ( .D(1'b0), .SETB(n11400), .RSTB(
        n_src_aox[203]), .CLK(clk), .Q(src_window[203]) );
  DFFSSRX1_HVT src_aox_reg_10__2_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[202]), .CLK(clk), .Q(src_window[202]) );
  DFFSSRX1_HVT src_aox_reg_10__1_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[201]), .CLK(clk), .Q(src_window[201]) );
  DFFSSRX1_HVT src_aox_reg_10__0_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[200]), .CLK(clk), .Q(src_window[200]) );
  DFFSSRX1_HVT src_aox_reg_11__7_ ( .D(1'b0), .SETB(n11400), .RSTB(
        n_src_aox[199]), .CLK(clk), .Q(src_window[199]) );
  DFFSSRX1_HVT src_aox_reg_11__6_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[198]), .CLK(clk), .Q(src_window[198]) );
  DFFSSRX1_HVT src_aox_reg_11__5_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[197]), .CLK(clk), .Q(src_window[197]) );
  DFFSSRX1_HVT src_aox_reg_11__4_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[196]), .CLK(clk), .Q(src_window[196]) );
  DFFSSRX1_HVT src_aox_reg_11__3_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[195]), .CLK(clk), .Q(src_window[195]) );
  DFFSSRX1_HVT src_aox_reg_11__2_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[194]), .CLK(clk), .Q(src_window[194]) );
  DFFSSRX1_HVT src_aox_reg_11__1_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[193]), .CLK(clk), .Q(src_window[193]) );
  DFFSSRX1_HVT src_aox_reg_11__0_ ( .D(1'b0), .SETB(n13000), .RSTB(
        n_src_aox[192]), .CLK(clk), .Q(src_window[192]) );
  DFFSSRX1_HVT src_aox_reg_12__7_ ( .D(1'b0), .SETB(N346), .RSTB(
        n_src_aox[191]), .CLK(clk), .Q(src_window[191]) );
  DFFSSRX1_HVT src_aox_reg_12__6_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[190]), .CLK(clk), .Q(src_window[190]) );
  DFFSSRX1_HVT src_aox_reg_12__5_ ( .D(1'b0), .SETB(n13000), .RSTB(
        n_src_aox[189]), .CLK(clk), .Q(src_window[189]) );
  DFFSSRX1_HVT src_aox_reg_12__4_ ( .D(1'b0), .SETB(n577), .RSTB(
        n_src_aox[188]), .CLK(clk), .Q(src_window[188]) );
  DFFSSRX1_HVT src_aox_reg_12__3_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[187]), .CLK(clk), .Q(src_window[187]) );
  DFFSSRX1_HVT src_aox_reg_12__2_ ( .D(1'b0), .SETB(n11400), .RSTB(
        n_src_aox[186]), .CLK(clk), .Q(src_window[186]) );
  DFFSSRX1_HVT src_aox_reg_12__1_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[185]), .CLK(clk), .Q(src_window[185]) );
  DFFSSRX1_HVT src_aox_reg_12__0_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[184]), .CLK(clk), .Q(src_window[184]) );
  DFFSSRX1_HVT src_aox_reg_13__7_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[183]), .CLK(clk), .Q(src_window[183]) );
  DFFSSRX1_HVT src_aox_reg_13__6_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[182]), .CLK(clk), .Q(src_window[182]) );
  DFFSSRX1_HVT src_aox_reg_13__5_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[181]), .CLK(clk), .Q(src_window[181]) );
  DFFSSRX1_HVT src_aox_reg_13__4_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[180]), .CLK(clk), .Q(src_window[180]) );
  DFFSSRX1_HVT src_aox_reg_13__3_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[179]), .CLK(clk), .Q(src_window[179]) );
  DFFSSRX1_HVT src_aox_reg_13__2_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[178]), .CLK(clk), .Q(src_window[178]) );
  DFFSSRX1_HVT src_aox_reg_13__1_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[177]), .CLK(clk), .Q(src_window[177]) );
  DFFSSRX1_HVT src_aox_reg_13__0_ ( .D(1'b0), .SETB(n577), .RSTB(
        n_src_aox[176]), .CLK(clk), .Q(src_window[176]) );
  DFFSSRX1_HVT src_aox_reg_14__7_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[175]), .CLK(clk), .Q(src_window[175]) );
  DFFSSRX1_HVT src_aox_reg_14__6_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[174]), .CLK(clk), .Q(src_window[174]) );
  DFFSSRX1_HVT src_aox_reg_14__5_ ( .D(1'b0), .SETB(n577), .RSTB(
        n_src_aox[173]), .CLK(clk), .Q(src_window[173]) );
  DFFSSRX1_HVT src_aox_reg_14__4_ ( .D(1'b0), .SETB(n13000), .RSTB(
        n_src_aox[172]), .CLK(clk), .Q(src_window[172]) );
  DFFSSRX1_HVT src_aox_reg_14__3_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[171]), .CLK(clk), .Q(src_window[171]) );
  DFFSSRX1_HVT src_aox_reg_14__2_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[170]), .CLK(clk), .Q(src_window[170]) );
  DFFSSRX1_HVT src_aox_reg_14__1_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[169]), .CLK(clk), .Q(src_window[169]) );
  DFFSSRX1_HVT src_aox_reg_14__0_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[168]), .CLK(clk), .Q(src_window[168]) );
  DFFSSRX1_HVT src_aox_reg_15__7_ ( .D(1'b0), .SETB(n11400), .RSTB(
        n_src_aox[167]), .CLK(clk), .Q(src_window[167]) );
  DFFSSRX1_HVT src_aox_reg_15__6_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[166]), .CLK(clk), .Q(src_window[166]) );
  DFFSSRX1_HVT src_aox_reg_15__5_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[165]), .CLK(clk), .Q(src_window[165]) );
  DFFSSRX1_HVT src_aox_reg_15__4_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[164]), .CLK(clk), .Q(src_window[164]) );
  DFFSSRX1_HVT src_aox_reg_15__3_ ( .D(1'b0), .SETB(n2600), .RSTB(
        n_src_aox[163]), .CLK(clk), .Q(src_window[163]) );
  DFFSSRX1_HVT src_aox_reg_15__2_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[162]), .CLK(clk), .Q(src_window[162]) );
  DFFSSRX1_HVT src_aox_reg_15__1_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[161]), .CLK(clk), .Q(src_window[161]) );
  DFFSSRX1_HVT src_aox_reg_15__0_ ( .D(1'b0), .SETB(n11400), .RSTB(
        n_src_aox[160]), .CLK(clk), .Q(src_window[160]) );
  DFFSSRX1_HVT src_aox_reg_16__7_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[159]), .CLK(clk), .Q(src_window[159]) );
  DFFSSRX1_HVT src_aox_reg_16__6_ ( .D(1'b0), .SETB(N346), .RSTB(
        n_src_aox[158]), .CLK(clk), .Q(src_window[158]) );
  DFFSSRX1_HVT src_aox_reg_16__5_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[157]), .CLK(clk), .Q(src_window[157]) );
  DFFSSRX1_HVT src_aox_reg_16__4_ ( .D(1'b0), .SETB(n577), .RSTB(
        n_src_aox[156]), .CLK(clk), .Q(src_window[156]) );
  DFFSSRX1_HVT src_aox_reg_16__3_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[155]), .CLK(clk), .Q(src_window[155]) );
  DFFSSRX1_HVT src_aox_reg_16__2_ ( .D(1'b0), .SETB(n11400), .RSTB(
        n_src_aox[154]), .CLK(clk), .Q(src_window[154]) );
  DFFSSRX1_HVT src_aox_reg_16__1_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[153]), .CLK(clk), .Q(src_window[153]) );
  DFFSSRX1_HVT src_aox_reg_16__0_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[152]), .CLK(clk), .Q(src_window[152]) );
  DFFSSRX1_HVT src_aox_reg_17__7_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[151]), .CLK(clk), .Q(src_window[151]) );
  DFFSSRX1_HVT src_aox_reg_17__6_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[150]), .CLK(clk), .Q(src_window[150]) );
  DFFSSRX1_HVT src_aox_reg_17__5_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[149]), .CLK(clk), .Q(src_window[149]) );
  DFFSSRX1_HVT src_aox_reg_17__4_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[148]), .CLK(clk), .Q(src_window[148]) );
  DFFSSRX1_HVT src_aox_reg_17__3_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[147]), .CLK(clk), .Q(src_window[147]) );
  DFFSSRX1_HVT src_aox_reg_17__2_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[146]), .CLK(clk), .Q(src_window[146]) );
  DFFSSRX1_HVT src_aox_reg_17__1_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[145]), .CLK(clk), .Q(src_window[145]) );
  DFFSSRX1_HVT src_aox_reg_17__0_ ( .D(1'b0), .SETB(n577), .RSTB(
        n_src_aox[144]), .CLK(clk), .Q(src_window[144]) );
  DFFSSRX1_HVT src_aox_reg_18__7_ ( .D(1'b0), .SETB(n2600), .RSTB(
        n_src_aox[143]), .CLK(clk), .Q(src_window[143]) );
  DFFSSRX1_HVT src_aox_reg_18__6_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[142]), .CLK(clk), .Q(src_window[142]) );
  DFFSSRX1_HVT src_aox_reg_18__5_ ( .D(1'b0), .SETB(n577), .RSTB(
        n_src_aox[141]), .CLK(clk), .Q(src_window[141]) );
  DFFSSRX1_HVT src_aox_reg_18__4_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[140]), .CLK(clk), .Q(src_window[140]) );
  DFFSSRX1_HVT src_aox_reg_18__3_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[139]), .CLK(clk), .Q(src_window[139]) );
  DFFSSRX1_HVT src_aox_reg_18__2_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[138]), .CLK(clk), .Q(src_window[138]) );
  DFFSSRX1_HVT src_aox_reg_18__1_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[137]), .CLK(clk), .Q(src_window[137]) );
  DFFSSRX1_HVT src_aox_reg_18__0_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[136]), .CLK(clk), .Q(src_window[136]) );
  DFFSSRX1_HVT src_aox_reg_19__7_ ( .D(1'b0), .SETB(n11400), .RSTB(
        n_src_aox[135]), .CLK(clk), .Q(src_window[135]) );
  DFFSSRX1_HVT src_aox_reg_19__6_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[134]), .CLK(clk), .Q(src_window[134]) );
  DFFSSRX1_HVT src_aox_reg_19__5_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[133]), .CLK(clk), .Q(src_window[133]) );
  DFFSSRX1_HVT src_aox_reg_19__4_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[132]), .CLK(clk), .Q(src_window[132]) );
  DFFSSRX1_HVT src_aox_reg_19__3_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[131]), .CLK(clk), .Q(src_window[131]) );
  DFFSSRX1_HVT src_aox_reg_19__2_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[130]), .CLK(clk), .Q(src_window[130]) );
  DFFSSRX1_HVT src_aox_reg_19__1_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[129]), .CLK(clk), .Q(src_window[129]) );
  DFFSSRX1_HVT src_aox_reg_19__0_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[128]), .CLK(clk), .Q(src_window[128]) );
  DFFSSRX1_HVT src_aox_reg_20__7_ ( .D(1'b0), .SETB(n2600), .RSTB(
        n_src_aox[127]), .CLK(clk), .Q(src_window[127]) );
  DFFSSRX1_HVT src_aox_reg_20__6_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[126]), .CLK(clk), .Q(src_window[126]) );
  DFFSSRX1_HVT src_aox_reg_20__5_ ( .D(1'b0), .SETB(n2600), .RSTB(
        n_src_aox[125]), .CLK(clk), .Q(src_window[125]) );
  DFFSSRX1_HVT src_aox_reg_20__4_ ( .D(1'b0), .SETB(n577), .RSTB(
        n_src_aox[124]), .CLK(clk), .Q(src_window[124]) );
  DFFSSRX1_HVT src_aox_reg_20__3_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[123]), .CLK(clk), .Q(src_window[123]) );
  DFFSSRX1_HVT src_aox_reg_20__2_ ( .D(1'b0), .SETB(n11400), .RSTB(
        n_src_aox[122]), .CLK(clk), .Q(src_window[122]) );
  DFFSSRX1_HVT src_aox_reg_20__1_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[121]), .CLK(clk), .Q(src_window[121]) );
  DFFSSRX1_HVT src_aox_reg_20__0_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[120]), .CLK(clk), .Q(src_window[120]) );
  DFFSSRX1_HVT src_aox_reg_21__7_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[119]), .CLK(clk), .Q(src_window[119]) );
  DFFSSRX1_HVT src_aox_reg_21__6_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[118]), .CLK(clk), .Q(src_window[118]) );
  DFFSSRX1_HVT src_aox_reg_21__5_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[117]), .CLK(clk), .Q(src_window[117]) );
  DFFSSRX1_HVT src_aox_reg_21__4_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[116]), .CLK(clk), .Q(src_window[116]) );
  DFFSSRX1_HVT src_aox_reg_21__3_ ( .D(1'b0), .SETB(n2600), .RSTB(
        n_src_aox[115]), .CLK(clk), .Q(src_window[115]) );
  DFFSSRX1_HVT src_aox_reg_21__2_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[114]), .CLK(clk), .Q(src_window[114]) );
  DFFSSRX1_HVT src_aox_reg_21__1_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[113]), .CLK(clk), .Q(src_window[113]) );
  DFFSSRX1_HVT src_aox_reg_21__0_ ( .D(1'b0), .SETB(n577), .RSTB(
        n_src_aox[112]), .CLK(clk), .Q(src_window[112]) );
  DFFSSRX1_HVT src_aox_reg_22__7_ ( .D(1'b0), .SETB(N346), .RSTB(
        n_src_aox[111]), .CLK(clk), .Q(src_window[111]) );
  DFFSSRX1_HVT src_aox_reg_22__6_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[110]), .CLK(clk), .Q(src_window[110]) );
  DFFSSRX1_HVT src_aox_reg_22__5_ ( .D(1'b0), .SETB(n577), .RSTB(
        n_src_aox[109]), .CLK(clk), .Q(src_window[109]) );
  DFFSSRX1_HVT src_aox_reg_22__4_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[108]), .CLK(clk), .Q(src_window[108]) );
  DFFSSRX1_HVT src_aox_reg_22__3_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[107]), .CLK(clk), .Q(src_window[107]) );
  DFFSSRX1_HVT src_aox_reg_22__2_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[106]), .CLK(clk), .Q(src_window[106]) );
  DFFSSRX1_HVT src_aox_reg_22__1_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[105]), .CLK(clk), .Q(src_window[105]) );
  DFFSSRX1_HVT src_aox_reg_22__0_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[104]), .CLK(clk), .Q(src_window[104]) );
  DFFSSRX1_HVT src_aox_reg_23__7_ ( .D(1'b0), .SETB(n11400), .RSTB(
        n_src_aox[103]), .CLK(clk), .Q(src_window[103]) );
  DFFSSRX1_HVT src_aox_reg_23__6_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[102]), .CLK(clk), .Q(src_window[102]) );
  DFFSSRX1_HVT src_aox_reg_23__5_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[101]), .CLK(clk), .Q(src_window[101]) );
  DFFSSRX1_HVT src_aox_reg_23__4_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[100]), .CLK(clk), .Q(src_window[100]) );
  DFFSSRX1_HVT src_aox_reg_23__3_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[99]), .CLK(clk), .Q(src_window[99]) );
  DFFSSRX1_HVT src_aox_reg_23__2_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[98]), .CLK(clk), .Q(src_window[98]) );
  DFFSSRX1_HVT src_aox_reg_23__1_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[97]), .CLK(clk), .Q(src_window[97]) );
  DFFSSRX1_HVT src_aox_reg_23__0_ ( .D(1'b0), .SETB(n13000), .RSTB(
        n_src_aox[96]), .CLK(clk), .Q(src_window[96]) );
  DFFSSRX1_HVT src_aox_reg_24__7_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[95]), .CLK(clk), .Q(src_window[95]) );
  DFFSSRX1_HVT src_aox_reg_24__6_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[94]), .CLK(clk), .Q(src_window[94]) );
  DFFSSRX1_HVT src_aox_reg_24__5_ ( .D(1'b0), .SETB(n13000), .RSTB(
        n_src_aox[93]), .CLK(clk), .Q(src_window[93]) );
  DFFSSRX1_HVT src_aox_reg_24__4_ ( .D(1'b0), .SETB(n577), .RSTB(n_src_aox[92]), .CLK(clk), .Q(src_window[92]) );
  DFFSSRX1_HVT src_aox_reg_24__3_ ( .D(1'b0), .SETB(n2600), .RSTB(
        n_src_aox[91]), .CLK(clk), .Q(src_window[91]) );
  DFFSSRX1_HVT src_aox_reg_24__2_ ( .D(1'b0), .SETB(n11400), .RSTB(
        n_src_aox[90]), .CLK(clk), .Q(src_window[90]) );
  DFFSSRX1_HVT src_aox_reg_24__1_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[89]), .CLK(clk), .Q(src_window[89]) );
  DFFSSRX1_HVT src_aox_reg_24__0_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[88]), .CLK(clk), .Q(src_window[88]) );
  DFFSSRX1_HVT src_aox_reg_25__7_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[87]), .CLK(clk), .Q(src_window[87]) );
  DFFSSRX1_HVT src_aox_reg_25__6_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[86]), .CLK(clk), .Q(src_window[86]) );
  DFFSSRX1_HVT src_aox_reg_25__5_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[85]), .CLK(clk), .Q(src_window[85]) );
  DFFSSRX1_HVT src_aox_reg_25__4_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[84]), .CLK(clk), .Q(src_window[84]) );
  DFFSSRX1_HVT src_aox_reg_25__3_ ( .D(1'b0), .SETB(n2600), .RSTB(
        n_src_aox[83]), .CLK(clk), .Q(src_window[83]) );
  DFFSSRX1_HVT src_aox_reg_25__2_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[82]), .CLK(clk), .Q(src_window[82]) );
  DFFSSRX1_HVT src_aox_reg_25__1_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[81]), .CLK(clk), .Q(src_window[81]) );
  DFFSSRX1_HVT src_aox_reg_25__0_ ( .D(1'b0), .SETB(n577), .RSTB(n_src_aox[80]), .CLK(clk), .Q(src_window[80]) );
  DFFSSRX1_HVT src_aox_reg_26__7_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[79]), .CLK(clk), .Q(src_window[79]) );
  DFFSSRX1_HVT src_aox_reg_26__6_ ( .D(1'b0), .SETB(n2600), .RSTB(
        n_src_aox[78]), .CLK(clk), .Q(src_window[78]) );
  DFFSSRX1_HVT src_aox_reg_26__5_ ( .D(1'b0), .SETB(n577), .RSTB(n_src_aox[77]), .CLK(clk), .Q(src_window[77]) );
  DFFSSRX1_HVT src_aox_reg_26__4_ ( .D(1'b0), .SETB(n13000), .RSTB(
        n_src_aox[76]), .CLK(clk), .Q(src_window[76]) );
  DFFSSRX1_HVT src_aox_reg_26__3_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[75]), .CLK(clk), .Q(src_window[75]) );
  DFFSSRX1_HVT src_aox_reg_26__2_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[74]), .CLK(clk), .Q(src_window[74]) );
  DFFSSRX1_HVT src_aox_reg_26__1_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[73]), .CLK(clk), .Q(src_window[73]) );
  DFFSSRX1_HVT src_aox_reg_26__0_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[72]), .CLK(clk), .Q(src_window[72]) );
  DFFSSRX1_HVT src_aox_reg_27__7_ ( .D(1'b0), .SETB(n11400), .RSTB(
        n_src_aox[71]), .CLK(clk), .Q(src_window[71]) );
  DFFSSRX1_HVT src_aox_reg_27__6_ ( .D(1'b0), .SETB(n13000), .RSTB(
        n_src_aox[70]), .CLK(clk), .Q(src_window[70]) );
  DFFSSRX1_HVT src_aox_reg_27__5_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[69]), .CLK(clk), .Q(src_window[69]) );
  DFFSSRX1_HVT src_aox_reg_27__4_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[68]), .CLK(clk), .Q(src_window[68]) );
  DFFSSRX1_HVT src_aox_reg_27__3_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[67]), .CLK(clk), .Q(src_window[67]) );
  DFFSSRX1_HVT src_aox_reg_27__2_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[66]), .CLK(clk), .Q(src_window[66]) );
  DFFSSRX1_HVT src_aox_reg_27__1_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[65]), .CLK(clk), .Q(src_window[65]) );
  DFFSSRX1_HVT src_aox_reg_27__0_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[64]), .CLK(clk), .Q(src_window[64]) );
  DFFSSRX1_HVT src_aox_reg_28__7_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[63]), .CLK(clk), .Q(src_window[63]) );
  DFFSSRX1_HVT src_aox_reg_28__6_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[62]), .CLK(clk), .Q(src_window[62]) );
  DFFSSRX1_HVT src_aox_reg_28__5_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[61]), .CLK(clk), .Q(src_window[61]) );
  DFFSSRX1_HVT src_aox_reg_28__4_ ( .D(1'b0), .SETB(N346), .RSTB(n_src_aox[60]), .CLK(clk), .Q(src_window[60]) );
  DFFSSRX1_HVT src_aox_reg_28__3_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[59]), .CLK(clk), .Q(src_window[59]) );
  DFFSSRX1_HVT src_aox_reg_28__2_ ( .D(1'b0), .SETB(n11400), .RSTB(
        n_src_aox[58]), .CLK(clk), .Q(src_window[58]) );
  DFFSSRX1_HVT src_aox_reg_28__1_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[57]), .CLK(clk), .Q(src_window[57]) );
  DFFSSRX1_HVT src_aox_reg_28__0_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[56]), .CLK(clk), .Q(src_window[56]) );
  DFFSSRX1_HVT src_aox_reg_29__7_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[55]), .CLK(clk), .Q(src_window[55]) );
  DFFSSRX1_HVT src_aox_reg_29__6_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[54]), .CLK(clk), .Q(src_window[54]) );
  DFFSSRX1_HVT src_aox_reg_29__5_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[53]), .CLK(clk), .Q(src_window[53]) );
  DFFSSRX1_HVT src_aox_reg_29__4_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[52]), .CLK(clk), .Q(src_window[52]) );
  DFFSSRX1_HVT src_aox_reg_29__3_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[51]), .CLK(clk), .Q(src_window[51]) );
  DFFSSRX1_HVT src_aox_reg_29__2_ ( .D(1'b0), .SETB(n11400), .RSTB(
        n_src_aox[50]), .CLK(clk), .Q(src_window[50]) );
  DFFSSRX1_HVT src_aox_reg_29__1_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[49]), .CLK(clk), .Q(src_window[49]) );
  DFFSSRX1_HVT src_aox_reg_29__0_ ( .D(1'b0), .SETB(n577), .RSTB(n_src_aox[48]), .CLK(clk), .Q(src_window[48]) );
  DFFSSRX1_HVT src_aox_reg_30__7_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[47]), .CLK(clk), .Q(src_window[47]) );
  DFFSSRX1_HVT src_aox_reg_30__6_ ( .D(1'b0), .SETB(n13000), .RSTB(
        n_src_aox[46]), .CLK(clk), .Q(src_window[46]) );
  DFFSSRX1_HVT src_aox_reg_30__5_ ( .D(1'b0), .SETB(n577), .RSTB(n_src_aox[45]), .CLK(clk), .Q(src_window[45]) );
  DFFSSRX1_HVT src_aox_reg_30__4_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[44]), .CLK(clk), .Q(src_window[44]) );
  DFFSSRX1_HVT src_aox_reg_30__3_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[43]), .CLK(clk), .Q(src_window[43]) );
  DFFSSRX1_HVT src_aox_reg_30__2_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[42]), .CLK(clk), .Q(src_window[42]) );
  DFFSSRX1_HVT src_aox_reg_30__1_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[41]), .CLK(clk), .Q(src_window[41]) );
  DFFSSRX1_HVT src_aox_reg_30__0_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[40]), .CLK(clk), .Q(src_window[40]) );
  DFFSSRX1_HVT src_aox_reg_31__7_ ( .D(1'b0), .SETB(n11400), .RSTB(
        n_src_aox[39]), .CLK(clk), .Q(src_window[39]) );
  DFFSSRX1_HVT src_aox_reg_31__6_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[38]), .CLK(clk), .Q(src_window[38]) );
  DFFSSRX1_HVT src_aox_reg_31__5_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[37]), .CLK(clk), .Q(src_window[37]) );
  DFFSSRX1_HVT src_aox_reg_31__4_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[36]), .CLK(clk), .Q(src_window[36]) );
  DFFSSRX1_HVT src_aox_reg_31__3_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[35]), .CLK(clk), .Q(src_window[35]) );
  DFFSSRX1_HVT src_aox_reg_31__2_ ( .D(1'b0), .SETB(n13000), .RSTB(
        n_src_aox[34]), .CLK(clk), .Q(src_window[34]) );
  DFFSSRX1_HVT src_aox_reg_31__1_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[33]), .CLK(clk), .Q(src_window[33]) );
  DFFSSRX1_HVT src_aox_reg_31__0_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[32]), .CLK(clk), .Q(src_window[32]) );
  DFFSSRX1_HVT src_aox_reg_32__7_ ( .D(1'b0), .SETB(n2600), .RSTB(
        n_src_aox[31]), .CLK(clk), .Q(src_window[31]) );
  DFFSSRX1_HVT src_aox_reg_32__6_ ( .D(1'b0), .SETB(n2580), .RSTB(
        n_src_aox[30]), .CLK(clk), .Q(src_window[30]) );
  DFFSSRX1_HVT src_aox_reg_32__5_ ( .D(1'b0), .SETB(n2600), .RSTB(
        n_src_aox[29]), .CLK(clk), .Q(src_window[29]) );
  DFFSSRX1_HVT src_aox_reg_32__4_ ( .D(1'b0), .SETB(N346), .RSTB(n_src_aox[28]), .CLK(clk), .Q(src_window[28]) );
  DFFSSRX1_HVT src_aox_reg_32__3_ ( .D(1'b0), .SETB(n2600), .RSTB(
        n_src_aox[27]), .CLK(clk), .Q(src_window[27]) );
  DFFSSRX1_HVT src_aox_reg_32__2_ ( .D(1'b0), .SETB(n11400), .RSTB(
        n_src_aox[26]), .CLK(clk), .Q(src_window[26]) );
  DFFSSRX1_HVT src_aox_reg_32__1_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[25]), .CLK(clk), .Q(src_window[25]) );
  DFFSSRX1_HVT src_aox_reg_32__0_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[24]), .CLK(clk), .Q(src_window[24]) );
  DFFSSRX1_HVT src_aox_reg_33__7_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[23]), .CLK(clk), .Q(src_window[23]) );
  DFFSSRX1_HVT src_aox_reg_33__6_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[22]), .CLK(clk), .Q(src_window[22]) );
  DFFSSRX1_HVT src_aox_reg_33__5_ ( .D(1'b0), .SETB(n2630), .RSTB(
        n_src_aox[21]), .CLK(clk), .Q(src_window[21]) );
  DFFSSRX1_HVT src_aox_reg_33__4_ ( .D(1'b0), .SETB(n9900), .RSTB(
        n_src_aox[20]), .CLK(clk), .Q(src_window[20]) );
  DFFSSRX1_HVT src_aox_reg_33__3_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[19]), .CLK(clk), .Q(src_window[19]) );
  DFFSSRX1_HVT src_aox_reg_33__2_ ( .D(1'b0), .SETB(n13000), .RSTB(
        n_src_aox[18]), .CLK(clk), .Q(src_window[18]) );
  DFFSSRX1_HVT src_aox_reg_33__1_ ( .D(1'b0), .SETB(n2620), .RSTB(
        n_src_aox[17]), .CLK(clk), .Q(src_window[17]) );
  DFFSSRX1_HVT src_aox_reg_33__0_ ( .D(1'b0), .SETB(n577), .RSTB(n_src_aox[16]), .CLK(clk), .Q(src_window[16]) );
  DFFSSRX1_HVT src_aox_reg_34__7_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[15]), .CLK(clk), .Q(src_window[15]) );
  DFFSSRX1_HVT src_aox_reg_34__6_ ( .D(1'b0), .SETB(n2590), .RSTB(
        n_src_aox[14]), .CLK(clk), .Q(src_window[14]) );
  DFFSSRX1_HVT src_aox_reg_34__5_ ( .D(1'b0), .SETB(n577), .RSTB(n_src_aox[13]), .CLK(clk), .Q(src_window[13]) );
  DFFSSRX1_HVT src_aox_reg_34__4_ ( .D(1'b0), .SETB(n2600), .RSTB(
        n_src_aox[12]), .CLK(clk), .Q(src_window[12]) );
  DFFSSRX1_HVT src_aox_reg_34__3_ ( .D(1'b0), .SETB(n13100), .RSTB(
        n_src_aox[11]), .CLK(clk), .Q(src_window[11]) );
  DFFSSRX1_HVT src_aox_reg_34__2_ ( .D(1'b0), .SETB(n9800), .RSTB(
        n_src_aox[10]), .CLK(clk), .Q(src_window[10]) );
  DFFSSRX1_HVT src_aox_reg_34__1_ ( .D(1'b0), .SETB(n9900), .RSTB(n_src_aox[9]), .CLK(clk), .Q(src_window[9]) );
  DFFSSRX1_HVT src_aox_reg_34__0_ ( .D(1'b0), .SETB(n2630), .RSTB(n_src_aox[8]), .CLK(clk), .Q(src_window[8]) );
  DFFSSRX1_HVT src_aox_reg_35__7_ ( .D(1'b0), .SETB(n11400), .RSTB(
        n_src_aox[7]), .CLK(clk), .Q(src_window[7]) );
  DFFSSRX1_HVT src_aox_reg_35__6_ ( .D(1'b0), .SETB(n2580), .RSTB(n_src_aox[6]), .CLK(clk), .Q(src_window[6]) );
  DFFSSRX1_HVT src_aox_reg_35__5_ ( .D(1'b0), .SETB(n2630), .RSTB(n_src_aox[5]), .CLK(clk), .Q(src_window[5]) );
  DFFSSRX1_HVT src_aox_reg_35__4_ ( .D(1'b0), .SETB(n11300), .RSTB(
        n_src_aox[4]), .CLK(clk), .Q(src_window[4]) );
  DFFSSRX1_HVT src_aox_reg_35__3_ ( .D(1'b0), .SETB(n2600), .RSTB(n_src_aox[3]), .CLK(clk), .Q(src_window[3]) );
  DFFSSRX1_HVT src_aox_reg_35__2_ ( .D(1'b0), .SETB(n2580), .RSTB(n_src_aox[2]), .CLK(clk), .Q(src_window[2]) );
  DFFSSRX1_HVT src_aox_reg_35__1_ ( .D(1'b0), .SETB(n2620), .RSTB(n_src_aox[1]), .CLK(clk), .Q(src_window[1]) );
  DFFSSRX1_HVT src_aox_reg_35__0_ ( .D(1'b0), .SETB(n13000), .RSTB(
        n_src_aox[0]), .CLK(clk), .Q(src_window[0]) );
  DFFSSRX1_HVT conv1_weight_reg_99_ ( .D(1'b0), .SETB(n13300), .RSTB(
        sram_rdata_weight[99]), .CLK(clk), .Q(conv1_weight[99]) );
  DFFSSRX1_HVT weight_reg_99_ ( .D(1'b0), .SETB(n13400), .RSTB(
        conv1_weight[99]), .CLK(clk), .Q(weight[99]) );
  DFFSSRX1_HVT conv1_weight_reg_98_ ( .D(1'b0), .SETB(n13200), .RSTB(
        sram_rdata_weight[98]), .CLK(clk), .Q(conv1_weight[98]) );
  DFFSSRX1_HVT weight_reg_98_ ( .D(1'b0), .SETB(n2450), .RSTB(conv1_weight[98]), .CLK(clk), .Q(weight[98]) );
  DFFSSRX1_HVT conv1_weight_reg_97_ ( .D(1'b0), .SETB(n2490), .RSTB(
        sram_rdata_weight[97]), .CLK(clk), .Q(conv1_weight[97]) );
  DFFSSRX1_HVT weight_reg_97_ ( .D(1'b0), .SETB(n2540), .RSTB(conv1_weight[97]), .CLK(clk), .Q(weight[97]) );
  DFFSSRX1_HVT conv1_weight_reg_96_ ( .D(1'b0), .SETB(n2420), .RSTB(
        sram_rdata_weight[96]), .CLK(clk), .Q(conv1_weight[96]) );
  DFFSSRX1_HVT weight_reg_96_ ( .D(1'b0), .SETB(n2830), .RSTB(conv1_weight[96]), .CLK(clk), .Q(weight[96]) );
  DFFSSRX1_HVT conv1_weight_reg_95_ ( .D(1'b0), .SETB(n2480), .RSTB(
        sram_rdata_weight[95]), .CLK(clk), .Q(conv1_weight[95]) );
  DFFSSRX1_HVT weight_reg_95_ ( .D(1'b0), .SETB(n2530), .RSTB(conv1_weight[95]), .CLK(clk), .Q(weight[95]) );
  DFFSSRX1_HVT conv1_weight_reg_94_ ( .D(1'b0), .SETB(n2410), .RSTB(
        sram_rdata_weight[94]), .CLK(clk), .Q(conv1_weight[94]) );
  DFFSSRX1_HVT weight_reg_94_ ( .D(1'b0), .SETB(n2460), .RSTB(conv1_weight[94]), .CLK(clk), .Q(weight[94]) );
  DFFSSRX1_HVT conv1_weight_reg_93_ ( .D(1'b0), .SETB(n2500), .RSTB(
        sram_rdata_weight[93]), .CLK(clk), .Q(conv1_weight[93]) );
  DFFSSRX1_HVT weight_reg_93_ ( .D(1'b0), .SETB(n2550), .RSTB(conv1_weight[93]), .CLK(clk), .Q(weight[93]) );
  DFFSSRX1_HVT conv1_weight_reg_92_ ( .D(1'b0), .SETB(n2430), .RSTB(
        sram_rdata_weight[92]), .CLK(clk), .Q(conv1_weight[92]) );
  DFFSSRX1_HVT weight_reg_92_ ( .D(1'b0), .SETB(n2500), .RSTB(conv1_weight[92]), .CLK(clk), .Q(weight[92]) );
  DFFSSRX1_HVT conv1_weight_reg_91_ ( .D(1'b0), .SETB(n12400), .RSTB(
        sram_rdata_weight[91]), .CLK(clk), .Q(conv1_weight[91]) );
  DFFSSRX1_HVT weight_reg_91_ ( .D(1'b0), .SETB(n12200), .RSTB(
        conv1_weight[91]), .CLK(clk), .Q(weight[91]) );
  DFFSSRX1_HVT conv1_weight_reg_90_ ( .D(1'b0), .SETB(n12300), .RSTB(
        sram_rdata_weight[90]), .CLK(clk), .Q(conv1_weight[90]) );
  DFFSSRX1_HVT weight_reg_90_ ( .D(1'b0), .SETB(n2450), .RSTB(conv1_weight[90]), .CLK(clk), .Q(weight[90]) );
  DFFSSRX1_HVT conv1_weight_reg_89_ ( .D(1'b0), .SETB(n2490), .RSTB(
        sram_rdata_weight[89]), .CLK(clk), .Q(conv1_weight[89]) );
  DFFSSRX1_HVT weight_reg_89_ ( .D(1'b0), .SETB(n2540), .RSTB(conv1_weight[89]), .CLK(clk), .Q(weight[89]) );
  DFFSSRX1_HVT conv1_weight_reg_88_ ( .D(1'b0), .SETB(n2420), .RSTB(
        sram_rdata_weight[88]), .CLK(clk), .Q(conv1_weight[88]) );
  DFFSSRX1_HVT weight_reg_88_ ( .D(1'b0), .SETB(n13400), .RSTB(
        conv1_weight[88]), .CLK(clk), .Q(weight[88]) );
  DFFSSRX1_HVT conv1_weight_reg_87_ ( .D(1'b0), .SETB(n2510), .RSTB(
        sram_rdata_weight[87]), .CLK(clk), .Q(conv1_weight[87]) );
  DFFSSRX1_HVT weight_reg_87_ ( .D(1'b0), .SETB(n2560), .RSTB(conv1_weight[87]), .CLK(clk), .Q(weight[87]) );
  DFFSSRX1_HVT conv1_weight_reg_86_ ( .D(1'b0), .SETB(n2440), .RSTB(
        sram_rdata_weight[86]), .CLK(clk), .Q(conv1_weight[86]) );
  DFFSSRX1_HVT weight_reg_86_ ( .D(1'b0), .SETB(n2460), .RSTB(conv1_weight[86]), .CLK(clk), .Q(weight[86]) );
  DFFSSRX1_HVT conv1_weight_reg_85_ ( .D(1'b0), .SETB(n2500), .RSTB(
        sram_rdata_weight[85]), .CLK(clk), .Q(conv1_weight[85]) );
  DFFSSRX1_HVT weight_reg_85_ ( .D(1'b0), .SETB(n2550), .RSTB(conv1_weight[85]), .CLK(clk), .Q(weight[85]) );
  DFFSSRX1_HVT conv1_weight_reg_84_ ( .D(1'b0), .SETB(n2430), .RSTB(
        sram_rdata_weight[84]), .CLK(clk), .Q(conv1_weight[84]) );
  DFFSSRX1_HVT weight_reg_84_ ( .D(1'b0), .SETB(n2460), .RSTB(conv1_weight[84]), .CLK(clk), .Q(weight[84]) );
  DFFSSRX1_HVT conv1_weight_reg_83_ ( .D(1'b0), .SETB(n12400), .RSTB(
        sram_rdata_weight[83]), .CLK(clk), .Q(conv1_weight[83]) );
  DFFSSRX1_HVT weight_reg_83_ ( .D(1'b0), .SETB(n12200), .RSTB(
        conv1_weight[83]), .CLK(clk), .Q(weight[83]) );
  DFFSSRX1_HVT conv1_weight_reg_82_ ( .D(1'b0), .SETB(n12300), .RSTB(
        sram_rdata_weight[82]), .CLK(clk), .Q(conv1_weight[82]) );
  DFFSSRX1_HVT weight_reg_82_ ( .D(1'b0), .SETB(n13400), .RSTB(
        conv1_weight[82]), .CLK(clk), .Q(weight[82]) );
  DFFSSRX1_HVT conv1_weight_reg_81_ ( .D(1'b0), .SETB(n2480), .RSTB(
        sram_rdata_weight[81]), .CLK(clk), .Q(conv1_weight[81]) );
  DFFSSRX1_HVT weight_reg_81_ ( .D(1'b0), .SETB(n2530), .RSTB(conv1_weight[81]), .CLK(clk), .Q(weight[81]) );
  DFFSSRX1_HVT conv1_weight_reg_80_ ( .D(1'b0), .SETB(n2410), .RSTB(
        sram_rdata_weight[80]), .CLK(clk), .Q(conv1_weight[80]) );
  DFFSSRX1_HVT weight_reg_80_ ( .D(1'b0), .SETB(n2840), .RSTB(conv1_weight[80]), .CLK(clk), .Q(weight[80]) );
  DFFSSRX1_HVT conv1_weight_reg_79_ ( .D(1'b0), .SETB(n2480), .RSTB(
        sram_rdata_weight[79]), .CLK(clk), .Q(conv1_weight[79]) );
  DFFSSRX1_HVT weight_reg_79_ ( .D(1'b0), .SETB(n2530), .RSTB(conv1_weight[79]), .CLK(clk), .Q(weight[79]) );
  DFFSSRX1_HVT conv1_weight_reg_78_ ( .D(1'b0), .SETB(n2410), .RSTB(
        sram_rdata_weight[78]), .CLK(clk), .Q(conv1_weight[78]) );
  DFFSSRX1_HVT weight_reg_78_ ( .D(1'b0), .SETB(n2460), .RSTB(conv1_weight[78]), .CLK(clk), .Q(weight[78]) );
  DFFSSRX1_HVT conv1_weight_reg_77_ ( .D(1'b0), .SETB(n2500), .RSTB(
        sram_rdata_weight[77]), .CLK(clk), .Q(conv1_weight[77]) );
  DFFSSRX1_HVT weight_reg_77_ ( .D(1'b0), .SETB(n2550), .RSTB(conv1_weight[77]), .CLK(clk), .Q(weight[77]) );
  DFFSSRX1_HVT conv1_weight_reg_76_ ( .D(1'b0), .SETB(n2430), .RSTB(
        sram_rdata_weight[76]), .CLK(clk), .Q(conv1_weight[76]) );
  DFFSSRX1_HVT weight_reg_76_ ( .D(1'b0), .SETB(n12300), .RSTB(
        conv1_weight[76]), .CLK(clk), .Q(weight[76]) );
  DFFSSRX1_HVT conv1_weight_reg_75_ ( .D(1'b0), .SETB(n13300), .RSTB(
        sram_rdata_weight[75]), .CLK(clk), .Q(conv1_weight[75]) );
  DFFSSRX1_HVT weight_reg_75_ ( .D(1'b0), .SETB(n13400), .RSTB(
        conv1_weight[75]), .CLK(clk), .Q(weight[75]) );
  DFFSSRX1_HVT conv1_weight_reg_74_ ( .D(1'b0), .SETB(n13200), .RSTB(
        sram_rdata_weight[74]), .CLK(clk), .Q(conv1_weight[74]) );
  DFFSSRX1_HVT weight_reg_74_ ( .D(1'b0), .SETB(n2840), .RSTB(conv1_weight[74]), .CLK(clk), .Q(weight[74]) );
  DFFSSRX1_HVT conv1_weight_reg_73_ ( .D(1'b0), .SETB(n2510), .RSTB(
        sram_rdata_weight[73]), .CLK(clk), .Q(conv1_weight[73]) );
  DFFSSRX1_HVT weight_reg_73_ ( .D(1'b0), .SETB(n2560), .RSTB(conv1_weight[73]), .CLK(clk), .Q(weight[73]) );
  DFFSSRX1_HVT conv1_weight_reg_72_ ( .D(1'b0), .SETB(n2440), .RSTB(
        sram_rdata_weight[72]), .CLK(clk), .Q(conv1_weight[72]) );
  DFFSSRX1_HVT weight_reg_72_ ( .D(1'b0), .SETB(n2550), .RSTB(conv1_weight[72]), .CLK(clk), .Q(weight[72]) );
  DFFSSRX1_HVT conv1_weight_reg_71_ ( .D(1'b0), .SETB(n2510), .RSTB(
        sram_rdata_weight[71]), .CLK(clk), .Q(conv1_weight[71]) );
  DFFSSRX1_HVT weight_reg_71_ ( .D(1'b0), .SETB(n2560), .RSTB(conv1_weight[71]), .CLK(clk), .Q(weight[71]) );
  DFFSSRX1_HVT conv1_weight_reg_70_ ( .D(1'b0), .SETB(n2440), .RSTB(
        sram_rdata_weight[70]), .CLK(clk), .Q(conv1_weight[70]) );
  DFFSSRX1_HVT weight_reg_70_ ( .D(1'b0), .SETB(n2460), .RSTB(conv1_weight[70]), .CLK(clk), .Q(weight[70]) );
  DFFSSRX1_HVT conv1_weight_reg_69_ ( .D(1'b0), .SETB(n2500), .RSTB(
        sram_rdata_weight[69]), .CLK(clk), .Q(conv1_weight[69]) );
  DFFSSRX1_HVT weight_reg_69_ ( .D(1'b0), .SETB(n2550), .RSTB(conv1_weight[69]), .CLK(clk), .Q(weight[69]) );
  DFFSSRX1_HVT conv1_weight_reg_68_ ( .D(1'b0), .SETB(n2430), .RSTB(
        sram_rdata_weight[68]), .CLK(clk), .Q(conv1_weight[68]) );
  DFFSSRX1_HVT weight_reg_68_ ( .D(1'b0), .SETB(n13200), .RSTB(
        conv1_weight[68]), .CLK(clk), .Q(weight[68]) );
  DFFSSRX1_HVT conv1_weight_reg_67_ ( .D(1'b0), .SETB(n12400), .RSTB(
        sram_rdata_weight[67]), .CLK(clk), .Q(conv1_weight[67]) );
  DFFSSRX1_HVT weight_reg_67_ ( .D(1'b0), .SETB(n12200), .RSTB(
        conv1_weight[67]), .CLK(clk), .Q(weight[67]) );
  DFFSSRX1_HVT conv1_weight_reg_66_ ( .D(1'b0), .SETB(n12300), .RSTB(
        sram_rdata_weight[66]), .CLK(clk), .Q(conv1_weight[66]) );
  DFFSSRX1_HVT weight_reg_66_ ( .D(1'b0), .SETB(n2450), .RSTB(conv1_weight[66]), .CLK(clk), .Q(weight[66]) );
  DFFSSRX1_HVT conv1_weight_reg_65_ ( .D(1'b0), .SETB(n2490), .RSTB(
        sram_rdata_weight[65]), .CLK(clk), .Q(conv1_weight[65]) );
  DFFSSRX1_HVT weight_reg_65_ ( .D(1'b0), .SETB(n2540), .RSTB(conv1_weight[65]), .CLK(clk), .Q(weight[65]) );
  DFFSSRX1_HVT conv1_weight_reg_64_ ( .D(1'b0), .SETB(n2420), .RSTB(
        sram_rdata_weight[64]), .CLK(clk), .Q(conv1_weight[64]) );
  DFFSSRX1_HVT weight_reg_64_ ( .D(1'b0), .SETB(n2850), .RSTB(conv1_weight[64]), .CLK(clk), .Q(weight[64]) );
  DFFSSRX1_HVT conv1_weight_reg_63_ ( .D(1'b0), .SETB(n2480), .RSTB(
        sram_rdata_weight[63]), .CLK(clk), .Q(conv1_weight[63]) );
  DFFSSRX1_HVT weight_reg_63_ ( .D(1'b0), .SETB(n2530), .RSTB(conv1_weight[63]), .CLK(clk), .Q(weight[63]) );
  DFFSSRX1_HVT conv1_weight_reg_62_ ( .D(1'b0), .SETB(n2410), .RSTB(
        sram_rdata_weight[62]), .CLK(clk), .Q(conv1_weight[62]) );
  DFFSSRX1_HVT weight_reg_62_ ( .D(1'b0), .SETB(n2460), .RSTB(conv1_weight[62]), .CLK(clk), .Q(weight[62]) );
  DFFSSRX1_HVT conv1_weight_reg_61_ ( .D(1'b0), .SETB(n2500), .RSTB(
        sram_rdata_weight[61]), .CLK(clk), .Q(conv1_weight[61]) );
  DFFSSRX1_HVT weight_reg_61_ ( .D(1'b0), .SETB(n2550), .RSTB(conv1_weight[61]), .CLK(clk), .Q(weight[61]) );
  DFFSSRX1_HVT conv1_weight_reg_60_ ( .D(1'b0), .SETB(n2430), .RSTB(
        sram_rdata_weight[60]), .CLK(clk), .Q(conv1_weight[60]) );
  DFFSSRX1_HVT weight_reg_60_ ( .D(1'b0), .SETB(n2460), .RSTB(conv1_weight[60]), .CLK(clk), .Q(weight[60]) );
  DFFSSRX1_HVT conv1_weight_reg_59_ ( .D(1'b0), .SETB(n12400), .RSTB(
        sram_rdata_weight[59]), .CLK(clk), .Q(conv1_weight[59]) );
  DFFSSRX1_HVT weight_reg_59_ ( .D(1'b0), .SETB(n12200), .RSTB(
        conv1_weight[59]), .CLK(clk), .Q(weight[59]) );
  DFFSSRX1_HVT conv1_weight_reg_58_ ( .D(1'b0), .SETB(n12300), .RSTB(
        sram_rdata_weight[58]), .CLK(clk), .Q(conv1_weight[58]) );
  DFFSSRX1_HVT weight_reg_58_ ( .D(1'b0), .SETB(n2450), .RSTB(conv1_weight[58]), .CLK(clk), .Q(weight[58]) );
  DFFSSRX1_HVT conv1_weight_reg_57_ ( .D(1'b0), .SETB(n2490), .RSTB(
        sram_rdata_weight[57]), .CLK(clk), .Q(conv1_weight[57]) );
  DFFSSRX1_HVT weight_reg_57_ ( .D(1'b0), .SETB(n2540), .RSTB(conv1_weight[57]), .CLK(clk), .Q(weight[57]) );
  DFFSSRX1_HVT conv1_weight_reg_56_ ( .D(1'b0), .SETB(n2420), .RSTB(
        sram_rdata_weight[56]), .CLK(clk), .Q(conv1_weight[56]) );
  DFFSSRX1_HVT weight_reg_56_ ( .D(1'b0), .SETB(n2850), .RSTB(conv1_weight[56]), .CLK(clk), .Q(weight[56]) );
  DFFSSRX1_HVT conv1_weight_reg_55_ ( .D(1'b0), .SETB(n2510), .RSTB(
        sram_rdata_weight[55]), .CLK(clk), .Q(conv1_weight[55]) );
  DFFSSRX1_HVT weight_reg_55_ ( .D(1'b0), .SETB(n2560), .RSTB(conv1_weight[55]), .CLK(clk), .Q(weight[55]) );
  DFFSSRX1_HVT conv1_weight_reg_54_ ( .D(1'b0), .SETB(n2440), .RSTB(
        sram_rdata_weight[54]), .CLK(clk), .Q(conv1_weight[54]) );
  DFFSSRX1_HVT weight_reg_54_ ( .D(1'b0), .SETB(n2460), .RSTB(conv1_weight[54]), .CLK(clk), .Q(weight[54]) );
  DFFSSRX1_HVT conv1_weight_reg_53_ ( .D(1'b0), .SETB(n2500), .RSTB(
        sram_rdata_weight[53]), .CLK(clk), .Q(conv1_weight[53]) );
  DFFSSRX1_HVT weight_reg_53_ ( .D(1'b0), .SETB(n2550), .RSTB(conv1_weight[53]), .CLK(clk), .Q(weight[53]) );
  DFFSSRX1_HVT conv1_weight_reg_52_ ( .D(1'b0), .SETB(n2430), .RSTB(
        sram_rdata_weight[52]), .CLK(clk), .Q(conv1_weight[52]) );
  DFFSSRX1_HVT weight_reg_52_ ( .D(1'b0), .SETB(n2460), .RSTB(conv1_weight[52]), .CLK(clk), .Q(weight[52]) );
  DFFSSRX1_HVT conv1_weight_reg_51_ ( .D(1'b0), .SETB(n13300), .RSTB(
        sram_rdata_weight[51]), .CLK(clk), .Q(conv1_weight[51]) );
  DFFSSRX1_HVT weight_reg_51_ ( .D(1'b0), .SETB(n13400), .RSTB(
        conv1_weight[51]), .CLK(clk), .Q(weight[51]) );
  DFFSSRX1_HVT conv1_weight_reg_50_ ( .D(1'b0), .SETB(n13200), .RSTB(
        sram_rdata_weight[50]), .CLK(clk), .Q(conv1_weight[50]) );
  DFFSSRX1_HVT weight_reg_50_ ( .D(1'b0), .SETB(n2550), .RSTB(conv1_weight[50]), .CLK(clk), .Q(weight[50]) );
  DFFSSRX1_HVT conv1_weight_reg_49_ ( .D(1'b0), .SETB(n2480), .RSTB(
        sram_rdata_weight[49]), .CLK(clk), .Q(conv1_weight[49]) );
  DFFSSRX1_HVT weight_reg_49_ ( .D(1'b0), .SETB(n2530), .RSTB(conv1_weight[49]), .CLK(clk), .Q(weight[49]) );
  DFFSSRX1_HVT conv1_weight_reg_48_ ( .D(1'b0), .SETB(n2410), .RSTB(
        sram_rdata_weight[48]), .CLK(clk), .Q(conv1_weight[48]) );
  DFFSSRX1_HVT weight_reg_48_ ( .D(1'b0), .SETB(n2830), .RSTB(conv1_weight[48]), .CLK(clk), .Q(weight[48]) );
  DFFSSRX1_HVT conv1_weight_reg_47_ ( .D(1'b0), .SETB(n2480), .RSTB(
        sram_rdata_weight[47]), .CLK(clk), .Q(conv1_weight[47]) );
  DFFSSRX1_HVT weight_reg_47_ ( .D(1'b0), .SETB(n2530), .RSTB(conv1_weight[47]), .CLK(clk), .Q(weight[47]) );
  DFFSSRX1_HVT conv1_weight_reg_46_ ( .D(1'b0), .SETB(n2410), .RSTB(
        sram_rdata_weight[46]), .CLK(clk), .Q(conv1_weight[46]) );
  DFFSSRX1_HVT weight_reg_46_ ( .D(1'b0), .SETB(n2460), .RSTB(conv1_weight[46]), .CLK(clk), .Q(weight[46]) );
  DFFSSRX1_HVT conv1_weight_reg_45_ ( .D(1'b0), .SETB(n2500), .RSTB(
        sram_rdata_weight[45]), .CLK(clk), .Q(conv1_weight[45]) );
  DFFSSRX1_HVT weight_reg_45_ ( .D(1'b0), .SETB(n2550), .RSTB(conv1_weight[45]), .CLK(clk), .Q(weight[45]) );
  DFFSSRX1_HVT conv1_weight_reg_44_ ( .D(1'b0), .SETB(n2430), .RSTB(
        sram_rdata_weight[44]), .CLK(clk), .Q(conv1_weight[44]) );
  DFFSSRX1_HVT weight_reg_44_ ( .D(1'b0), .SETB(n13400), .RSTB(
        conv1_weight[44]), .CLK(clk), .Q(weight[44]) );
  DFFSSRX1_HVT conv1_weight_reg_43_ ( .D(1'b0), .SETB(n12400), .RSTB(
        sram_rdata_weight[43]), .CLK(clk), .Q(conv1_weight[43]) );
  DFFSSRX1_HVT weight_reg_43_ ( .D(1'b0), .SETB(n12200), .RSTB(
        conv1_weight[43]), .CLK(clk), .Q(weight[43]) );
  DFFSSRX1_HVT conv1_weight_reg_42_ ( .D(1'b0), .SETB(n12300), .RSTB(
        sram_rdata_weight[42]), .CLK(clk), .Q(conv1_weight[42]) );
  DFFSSRX1_HVT weight_reg_42_ ( .D(1'b0), .SETB(n2830), .RSTB(conv1_weight[42]), .CLK(clk), .Q(weight[42]) );
  DFFSSRX1_HVT conv1_weight_reg_41_ ( .D(1'b0), .SETB(n2510), .RSTB(
        sram_rdata_weight[41]), .CLK(clk), .Q(conv1_weight[41]) );
  DFFSSRX1_HVT weight_reg_41_ ( .D(1'b0), .SETB(n2560), .RSTB(conv1_weight[41]), .CLK(clk), .Q(weight[41]) );
  DFFSSRX1_HVT conv1_weight_reg_40_ ( .D(1'b0), .SETB(n2440), .RSTB(
        sram_rdata_weight[40]), .CLK(clk), .Q(conv1_weight[40]) );
  DFFSSRX1_HVT weight_reg_40_ ( .D(1'b0), .SETB(n2850), .RSTB(conv1_weight[40]), .CLK(clk), .Q(weight[40]) );
  DFFSSRX1_HVT conv1_weight_reg_39_ ( .D(1'b0), .SETB(n2510), .RSTB(
        sram_rdata_weight[39]), .CLK(clk), .Q(conv1_weight[39]) );
  DFFSSRX1_HVT weight_reg_39_ ( .D(1'b0), .SETB(n2560), .RSTB(conv1_weight[39]), .CLK(clk), .Q(weight[39]) );
  DFFSSRX1_HVT conv1_weight_reg_38_ ( .D(1'b0), .SETB(n2440), .RSTB(
        sram_rdata_weight[38]), .CLK(clk), .Q(conv1_weight[38]) );
  DFFSSRX1_HVT weight_reg_38_ ( .D(1'b0), .SETB(n2460), .RSTB(conv1_weight[38]), .CLK(clk), .Q(weight[38]) );
  DFFSSRX1_HVT conv1_weight_reg_37_ ( .D(1'b0), .SETB(n2500), .RSTB(
        sram_rdata_weight[37]), .CLK(clk), .Q(conv1_weight[37]) );
  DFFSSRX1_HVT weight_reg_37_ ( .D(1'b0), .SETB(n2550), .RSTB(conv1_weight[37]), .CLK(clk), .Q(weight[37]) );
  DFFSSRX1_HVT conv1_weight_reg_36_ ( .D(1'b0), .SETB(n2430), .RSTB(
        sram_rdata_weight[36]), .CLK(clk), .Q(conv1_weight[36]) );
  DFFSSRX1_HVT weight_reg_36_ ( .D(1'b0), .SETB(n2460), .RSTB(conv1_weight[36]), .CLK(clk), .Q(weight[36]) );
  DFFSSRX1_HVT conv1_weight_reg_35_ ( .D(1'b0), .SETB(n12400), .RSTB(
        sram_rdata_weight[35]), .CLK(clk), .Q(conv1_weight[35]) );
  DFFSSRX1_HVT weight_reg_35_ ( .D(1'b0), .SETB(n12200), .RSTB(
        conv1_weight[35]), .CLK(clk), .Q(weight[35]) );
  DFFSSRX1_HVT conv1_weight_reg_34_ ( .D(1'b0), .SETB(n12300), .RSTB(
        sram_rdata_weight[34]), .CLK(clk), .Q(conv1_weight[34]) );
  DFFSSRX1_HVT weight_reg_34_ ( .D(1'b0), .SETB(n2450), .RSTB(conv1_weight[34]), .CLK(clk), .Q(weight[34]) );
  DFFSSRX1_HVT conv1_weight_reg_33_ ( .D(1'b0), .SETB(n2490), .RSTB(
        sram_rdata_weight[33]), .CLK(clk), .Q(conv1_weight[33]) );
  DFFSSRX1_HVT weight_reg_33_ ( .D(1'b0), .SETB(n2540), .RSTB(conv1_weight[33]), .CLK(clk), .Q(weight[33]) );
  DFFSSRX1_HVT conv1_weight_reg_32_ ( .D(1'b0), .SETB(n2420), .RSTB(
        sram_rdata_weight[32]), .CLK(clk), .Q(conv1_weight[32]) );
  DFFSSRX1_HVT weight_reg_32_ ( .D(1'b0), .SETB(n2840), .RSTB(conv1_weight[32]), .CLK(clk), .Q(weight[32]) );
  DFFSSRX1_HVT conv1_weight_reg_31_ ( .D(1'b0), .SETB(n2480), .RSTB(
        sram_rdata_weight[31]), .CLK(clk), .Q(conv1_weight[31]) );
  DFFSSRX1_HVT weight_reg_31_ ( .D(1'b0), .SETB(n2530), .RSTB(conv1_weight[31]), .CLK(clk), .Q(weight[31]) );
  DFFSSRX1_HVT conv1_weight_reg_30_ ( .D(1'b0), .SETB(n2410), .RSTB(
        sram_rdata_weight[30]), .CLK(clk), .Q(conv1_weight[30]) );
  DFFSSRX1_HVT weight_reg_30_ ( .D(1'b0), .SETB(n2460), .RSTB(conv1_weight[30]), .CLK(clk), .Q(weight[30]) );
  DFFSSRX1_HVT conv1_weight_reg_29_ ( .D(1'b0), .SETB(n2500), .RSTB(
        sram_rdata_weight[29]), .CLK(clk), .Q(conv1_weight[29]) );
  DFFSSRX1_HVT weight_reg_29_ ( .D(1'b0), .SETB(n2550), .RSTB(conv1_weight[29]), .CLK(clk), .Q(weight[29]) );
  DFFSSRX1_HVT conv1_weight_reg_28_ ( .D(1'b0), .SETB(n2430), .RSTB(
        sram_rdata_weight[28]), .CLK(clk), .Q(conv1_weight[28]) );
  DFFSSRX1_HVT weight_reg_28_ ( .D(1'b0), .SETB(n2850), .RSTB(conv1_weight[28]), .CLK(clk), .Q(weight[28]) );
  DFFSSRX1_HVT conv1_weight_reg_27_ ( .D(1'b0), .SETB(n13300), .RSTB(
        sram_rdata_weight[27]), .CLK(clk), .Q(conv1_weight[27]) );
  DFFSSRX1_HVT weight_reg_27_ ( .D(1'b0), .SETB(n13400), .RSTB(
        conv1_weight[27]), .CLK(clk), .Q(weight[27]) );
  DFFSSRX1_HVT conv1_weight_reg_26_ ( .D(1'b0), .SETB(n13200), .RSTB(
        sram_rdata_weight[26]), .CLK(clk), .Q(conv1_weight[26]) );
  DFFSSRX1_HVT weight_reg_26_ ( .D(1'b0), .SETB(n2450), .RSTB(conv1_weight[26]), .CLK(clk), .Q(weight[26]) );
  DFFSSRX1_HVT conv1_weight_reg_25_ ( .D(1'b0), .SETB(n2490), .RSTB(
        sram_rdata_weight[25]), .CLK(clk), .Q(conv1_weight[25]) );
  DFFSSRX1_HVT weight_reg_25_ ( .D(1'b0), .SETB(n2540), .RSTB(conv1_weight[25]), .CLK(clk), .Q(weight[25]) );
  DFFSSRX1_HVT conv1_weight_reg_24_ ( .D(1'b0), .SETB(n2420), .RSTB(
        sram_rdata_weight[24]), .CLK(clk), .Q(conv1_weight[24]) );
  DFFSSRX1_HVT weight_reg_24_ ( .D(1'b0), .SETB(n13300), .RSTB(
        conv1_weight[24]), .CLK(clk), .Q(weight[24]) );
  DFFSSRX1_HVT conv1_weight_reg_23_ ( .D(1'b0), .SETB(n2510), .RSTB(
        sram_rdata_weight[23]), .CLK(clk), .Q(conv1_weight[23]) );
  DFFSSRX1_HVT weight_reg_23_ ( .D(1'b0), .SETB(n2560), .RSTB(conv1_weight[23]), .CLK(clk), .Q(weight[23]) );
  DFFSSRX1_HVT conv1_weight_reg_22_ ( .D(1'b0), .SETB(n2440), .RSTB(
        sram_rdata_weight[22]), .CLK(clk), .Q(conv1_weight[22]) );
  DFFSSRX1_HVT weight_reg_22_ ( .D(1'b0), .SETB(n2460), .RSTB(conv1_weight[22]), .CLK(clk), .Q(weight[22]) );
  DFFSSRX1_HVT conv1_weight_reg_21_ ( .D(1'b0), .SETB(n2500), .RSTB(
        sram_rdata_weight[21]), .CLK(clk), .Q(conv1_weight[21]) );
  DFFSSRX1_HVT weight_reg_21_ ( .D(1'b0), .SETB(n2550), .RSTB(conv1_weight[21]), .CLK(clk), .Q(weight[21]) );
  DFFSSRX1_HVT conv1_weight_reg_20_ ( .D(1'b0), .SETB(n2430), .RSTB(
        sram_rdata_weight[20]), .CLK(clk), .Q(conv1_weight[20]) );
  DFFSSRX1_HVT weight_reg_20_ ( .D(1'b0), .SETB(n13300), .RSTB(
        conv1_weight[20]), .CLK(clk), .Q(weight[20]) );
  DFFSSRX1_HVT conv1_weight_reg_19_ ( .D(1'b0), .SETB(n12400), .RSTB(
        sram_rdata_weight[19]), .CLK(clk), .Q(conv1_weight[19]) );
  DFFSSRX1_HVT weight_reg_19_ ( .D(1'b0), .SETB(n12200), .RSTB(
        conv1_weight[19]), .CLK(clk), .Q(weight[19]) );
  DFFSSRX1_HVT conv1_weight_reg_18_ ( .D(1'b0), .SETB(n12300), .RSTB(
        sram_rdata_weight[18]), .CLK(clk), .Q(conv1_weight[18]) );
  DFFSSRX1_HVT weight_reg_18_ ( .D(1'b0), .SETB(n12400), .RSTB(
        conv1_weight[18]), .CLK(clk), .Q(weight[18]) );
  DFFSSRX1_HVT conv1_weight_reg_17_ ( .D(1'b0), .SETB(n2480), .RSTB(
        sram_rdata_weight[17]), .CLK(clk), .Q(conv1_weight[17]) );
  DFFSSRX1_HVT weight_reg_17_ ( .D(1'b0), .SETB(n2530), .RSTB(conv1_weight[17]), .CLK(clk), .Q(weight[17]) );
  DFFSSRX1_HVT conv1_weight_reg_16_ ( .D(1'b0), .SETB(n2410), .RSTB(
        sram_rdata_weight[16]), .CLK(clk), .Q(conv1_weight[16]) );
  DFFSSRX1_HVT weight_reg_16_ ( .D(1'b0), .SETB(n2450), .RSTB(conv1_weight[16]), .CLK(clk), .Q(weight[16]) );
  DFFSSRX1_HVT conv1_weight_reg_15_ ( .D(1'b0), .SETB(n2490), .RSTB(
        sram_rdata_weight[15]), .CLK(clk), .Q(conv1_weight[15]) );
  DFFSSRX1_HVT weight_reg_15_ ( .D(1'b0), .SETB(n2540), .RSTB(conv1_weight[15]), .CLK(clk), .Q(weight[15]) );
  DFFSSRX1_HVT conv1_weight_reg_14_ ( .D(1'b0), .SETB(n2420), .RSTB(
        sram_rdata_weight[14]), .CLK(clk), .Q(conv1_weight[14]) );
  DFFSSRX1_HVT weight_reg_14_ ( .D(1'b0), .SETB(n12400), .RSTB(
        conv1_weight[14]), .CLK(clk), .Q(weight[14]) );
  DFFSSRX1_HVT conv1_weight_reg_13_ ( .D(1'b0), .SETB(n2480), .RSTB(
        sram_rdata_weight[13]), .CLK(clk), .Q(conv1_weight[13]) );
  DFFSSRX1_HVT weight_reg_13_ ( .D(1'b0), .SETB(n2530), .RSTB(conv1_weight[13]), .CLK(clk), .Q(weight[13]) );
  DFFSSRX1_HVT conv1_weight_reg_12_ ( .D(1'b0), .SETB(n2410), .RSTB(
        sram_rdata_weight[12]), .CLK(clk), .Q(conv1_weight[12]) );
  DFFSSRX1_HVT weight_reg_12_ ( .D(1'b0), .SETB(n2460), .RSTB(conv1_weight[12]), .CLK(clk), .Q(weight[12]) );
  DFFSSRX1_HVT conv1_weight_reg_11_ ( .D(1'b0), .SETB(n12400), .RSTB(
        sram_rdata_weight[11]), .CLK(clk), .Q(conv1_weight[11]) );
  DFFSSRX1_HVT weight_reg_11_ ( .D(1'b0), .SETB(n12200), .RSTB(
        conv1_weight[11]), .CLK(clk), .Q(weight[11]) );
  DFFSSRX1_HVT conv1_weight_reg_10_ ( .D(1'b0), .SETB(n12300), .RSTB(
        sram_rdata_weight[10]), .CLK(clk), .Q(conv1_weight[10]) );
  DFFSSRX1_HVT weight_reg_10_ ( .D(1'b0), .SETB(n2850), .RSTB(conv1_weight[10]), .CLK(clk), .Q(weight[10]) );
  DFFSSRX1_HVT conv1_weight_reg_9_ ( .D(1'b0), .SETB(n2510), .RSTB(
        sram_rdata_weight[9]), .CLK(clk), .Q(conv1_weight[9]) );
  DFFSSRX1_HVT weight_reg_9_ ( .D(1'b0), .SETB(n2560), .RSTB(conv1_weight[9]), 
        .CLK(clk), .Q(weight[9]) );
  DFFSSRX1_HVT conv1_weight_reg_8_ ( .D(1'b0), .SETB(n2440), .RSTB(
        sram_rdata_weight[8]), .CLK(clk), .Q(conv1_weight[8]) );
  DFFSSRX1_HVT weight_reg_8_ ( .D(1'b0), .SETB(n2450), .RSTB(conv1_weight[8]), 
        .CLK(clk), .Q(weight[8]) );
  DFFSSRX1_HVT conv1_weight_reg_7_ ( .D(1'b0), .SETB(n2490), .RSTB(
        sram_rdata_weight[7]), .CLK(clk), .Q(conv1_weight[7]) );
  DFFSSRX1_HVT weight_reg_7_ ( .D(1'b0), .SETB(n2540), .RSTB(conv1_weight[7]), 
        .CLK(clk), .Q(weight[7]) );
  DFFSSRX1_HVT conv1_weight_reg_6_ ( .D(1'b0), .SETB(n2420), .RSTB(
        sram_rdata_weight[6]), .CLK(clk), .Q(conv1_weight[6]) );
  DFFSSRX1_HVT weight_reg_6_ ( .D(1'b0), .SETB(n2830), .RSTB(conv1_weight[6]), 
        .CLK(clk), .Q(weight[6]) );
  DFFSSRX1_HVT conv1_weight_reg_5_ ( .D(1'b0), .SETB(n2510), .RSTB(
        sram_rdata_weight[5]), .CLK(clk), .Q(conv1_weight[5]) );
  DFFSSRX1_HVT weight_reg_5_ ( .D(1'b0), .SETB(n2560), .RSTB(conv1_weight[5]), 
        .CLK(clk), .Q(weight[5]) );
  DFFSSRX1_HVT conv1_weight_reg_4_ ( .D(1'b0), .SETB(n2440), .RSTB(
        sram_rdata_weight[4]), .CLK(clk), .Q(conv1_weight[4]) );
  DFFSSRX1_HVT weight_reg_4_ ( .D(1'b0), .SETB(n12400), .RSTB(conv1_weight[4]), 
        .CLK(clk), .Q(weight[4]) );
  DFFSSRX1_HVT conv1_weight_reg_3_ ( .D(1'b0), .SETB(n13300), .RSTB(
        sram_rdata_weight[3]), .CLK(clk), .Q(conv1_weight[3]) );
  DFFSSRX1_HVT weight_reg_3_ ( .D(1'b0), .SETB(n13400), .RSTB(conv1_weight[3]), 
        .CLK(clk), .Q(weight[3]) );
  DFFSSRX1_HVT conv1_weight_reg_2_ ( .D(1'b0), .SETB(n13200), .RSTB(
        sram_rdata_weight[2]), .CLK(clk), .Q(conv1_weight[2]) );
  DFFSSRX1_HVT weight_reg_2_ ( .D(1'b0), .SETB(n2450), .RSTB(conv1_weight[2]), 
        .CLK(clk), .Q(weight[2]) );
  DFFSSRX1_HVT conv1_weight_reg_1_ ( .D(1'b0), .SETB(n2490), .RSTB(
        sram_rdata_weight[1]), .CLK(clk), .Q(conv1_weight[1]) );
  DFFSSRX1_HVT weight_reg_1_ ( .D(1'b0), .SETB(n2540), .RSTB(conv1_weight[1]), 
        .CLK(clk), .Q(weight[1]) );
  DFFSSRX1_HVT conv1_weight_reg_0_ ( .D(1'b0), .SETB(n2420), .RSTB(
        sram_rdata_weight[0]), .CLK(clk), .Q(conv1_weight[0]) );
  DFFSSRX1_HVT weight_reg_0_ ( .D(1'b0), .SETB(n2850), .RSTB(conv1_weight[0]), 
        .CLK(clk), .Q(weight[0]) );
  DFFSSRX1_HVT sram_rdata_8_reg_31_ ( .D(1'b0), .SETB(n2480), .RSTB(N326), 
        .CLK(clk), .Q(sram_rdata_8[31]), .QN(n3170) );
  DFFSSRX1_HVT sram_rdata_8_reg_30_ ( .D(1'b0), .SETB(n12200), .RSTB(N325), 
        .CLK(clk), .Q(sram_rdata_8[30]), .QN(n3160) );
  DFFSSRX1_HVT sram_rdata_8_reg_29_ ( .D(1'b0), .SETB(n2440), .RSTB(N324), 
        .CLK(clk), .Q(sram_rdata_8[29]), .QN(n3150) );
  DFFSSRX1_HVT sram_rdata_8_reg_28_ ( .D(1'b0), .SETB(n2840), .RSTB(N323), 
        .CLK(clk), .Q(sram_rdata_8[28]), .QN(n3140) );
  DFFSSRX1_HVT sram_rdata_8_reg_27_ ( .D(1'b0), .SETB(n2480), .RSTB(N322), 
        .CLK(clk), .Q(sram_rdata_8[27]), .QN(n3130) );
  DFFSSRX1_HVT sram_rdata_8_reg_26_ ( .D(1'b0), .SETB(n2560), .RSTB(N321), 
        .CLK(clk), .Q(sram_rdata_8[26]), .QN(n3120) );
  DFFSSRX1_HVT sram_rdata_8_reg_25_ ( .D(1'b0), .SETB(n2440), .RSTB(N320), 
        .CLK(clk), .Q(sram_rdata_8[25]), .QN(n3110) );
  DFFSSRX1_HVT sram_rdata_8_reg_24_ ( .D(1'b0), .SETB(n2830), .RSTB(N319), 
        .CLK(clk), .Q(sram_rdata_8[24]), .QN(n3100) );
  DFFSSRX1_HVT sram_rdata_8_reg_23_ ( .D(1'b0), .SETB(n12400), .RSTB(N318), 
        .CLK(clk), .Q(sram_rdata_8[23]), .QN(n3090) );
  DFFSSRX1_HVT sram_rdata_8_reg_22_ ( .D(1'b0), .SETB(n2560), .RSTB(N317), 
        .CLK(clk), .Q(sram_rdata_8[22]), .QN(n3080) );
  DFFSSRX1_HVT sram_rdata_8_reg_21_ ( .D(1'b0), .SETB(n13200), .RSTB(N316), 
        .CLK(clk), .Q(sram_rdata_8[21]), .QN(n3070) );
  DFFSSRX1_HVT sram_rdata_8_reg_20_ ( .D(1'b0), .SETB(n12300), .RSTB(N315), 
        .CLK(clk), .Q(sram_rdata_8[20]), .QN(n3060) );
  DFFSSRX1_HVT sram_rdata_8_reg_19_ ( .D(1'b0), .SETB(n2510), .RSTB(N314), 
        .CLK(clk), .Q(sram_rdata_8[19]), .QN(n3050) );
  DFFSSRX1_HVT sram_rdata_8_reg_18_ ( .D(1'b0), .SETB(n2560), .RSTB(N313), 
        .CLK(clk), .Q(sram_rdata_8[18]), .QN(n3040) );
  DFFSSRX1_HVT sram_rdata_8_reg_17_ ( .D(1'b0), .SETB(n2420), .RSTB(N312), 
        .CLK(clk), .Q(sram_rdata_8[17]), .QN(n3030) );
  DFFSSRX1_HVT sram_rdata_8_reg_16_ ( .D(1'b0), .SETB(n2830), .RSTB(N311), 
        .CLK(clk), .Q(sram_rdata_8[16]), .QN(n3020) );
  DFFSSRX1_HVT sram_rdata_8_reg_15_ ( .D(1'b0), .SETB(n2510), .RSTB(N310), 
        .CLK(clk), .Q(sram_rdata_8[15]), .QN(n3010) );
  DFFSSRX1_HVT sram_rdata_8_reg_14_ ( .D(1'b0), .SETB(n12200), .RSTB(N309), 
        .CLK(clk), .Q(sram_rdata_8[14]), .QN(n3000) );
  DFFSSRX1_HVT sram_rdata_8_reg_13_ ( .D(1'b0), .SETB(n2420), .RSTB(N308), 
        .CLK(clk), .Q(sram_rdata_8[13]), .QN(n2990) );
  DFFSSRX1_HVT sram_rdata_8_reg_12_ ( .D(1'b0), .SETB(n2850), .RSTB(N307), 
        .CLK(clk), .Q(sram_rdata_8[12]), .QN(n2980) );
  DFFSSRX1_HVT sram_rdata_8_reg_11_ ( .D(1'b0), .SETB(n2510), .RSTB(N306), 
        .CLK(clk), .Q(sram_rdata_8[11]), .QN(n2970) );
  DFFSSRX1_HVT sram_rdata_8_reg_10_ ( .D(1'b0), .SETB(n2540), .RSTB(N305), 
        .CLK(clk), .Q(sram_rdata_8[10]), .QN(n2960) );
  DFFSSRX1_HVT sram_rdata_8_reg_9_ ( .D(1'b0), .SETB(n2410), .RSTB(N304), 
        .CLK(clk), .Q(sram_rdata_8[9]), .QN(n2950) );
  DFFSSRX1_HVT sram_rdata_8_reg_8_ ( .D(1'b0), .SETB(n2830), .RSTB(N303), 
        .CLK(clk), .Q(sram_rdata_8[8]), .QN(n2940) );
  DFFSSRX1_HVT sram_rdata_8_reg_7_ ( .D(1'b0), .SETB(n12400), .RSTB(N302), 
        .CLK(clk), .Q(sram_rdata_8[7]), .QN(n2930) );
  DFFSSRX1_HVT sram_rdata_8_reg_6_ ( .D(1'b0), .SETB(n2540), .RSTB(N301), 
        .CLK(clk), .Q(sram_rdata_8[6]), .QN(n2920) );
  DFFSSRX1_HVT sram_rdata_8_reg_5_ ( .D(1'b0), .SETB(n13200), .RSTB(N300), 
        .CLK(clk), .Q(sram_rdata_8[5]), .QN(n2910) );
  DFFSSRX1_HVT sram_rdata_8_reg_4_ ( .D(1'b0), .SETB(n2850), .RSTB(N299), 
        .CLK(clk), .Q(sram_rdata_8[4]), .QN(n2900) );
  DFFSSRX1_HVT sram_rdata_8_reg_3_ ( .D(1'b0), .SETB(n2490), .RSTB(N298), 
        .CLK(clk), .Q(sram_rdata_8[3]), .QN(n2890) );
  DFFSSRX1_HVT sram_rdata_8_reg_2_ ( .D(1'b0), .SETB(n2530), .RSTB(N297), 
        .CLK(clk), .Q(sram_rdata_8[2]), .QN(n2880) );
  DFFSSRX1_HVT sram_rdata_8_reg_1_ ( .D(1'b0), .SETB(n2420), .RSTB(N296), 
        .CLK(clk), .Q(sram_rdata_8[1]), .QN(n2870) );
  DFFSSRX1_HVT sram_rdata_8_reg_0_ ( .D(1'b0), .SETB(n2430), .RSTB(N295), 
        .CLK(clk), .Q(sram_rdata_8[0]), .QN(n573) );
  DFFSSRX1_HVT sram_rdata_0_reg_31_ ( .D(1'b0), .SETB(n12300), .RSTB(N70), 
        .CLK(clk), .Q(sram_rdata_0[31]), .QN(n476) );
  DFFSSRX1_HVT sram_rdata_0_reg_30_ ( .D(1'b0), .SETB(n2490), .RSTB(N69), 
        .CLK(clk), .Q(sram_rdata_0[30]), .QN(n475) );
  DFFSSRX1_HVT sram_rdata_0_reg_29_ ( .D(1'b0), .SETB(n2560), .RSTB(N68), 
        .CLK(clk), .Q(sram_rdata_0[29]), .QN(n474) );
  DFFSSRX1_HVT sram_rdata_0_reg_28_ ( .D(1'b0), .SETB(n2410), .RSTB(N67), 
        .CLK(clk), .Q(sram_rdata_0[28]), .QN(n473) );
  DFFSSRX1_HVT sram_rdata_0_reg_27_ ( .D(1'b0), .SETB(n12200), .RSTB(N66), 
        .CLK(clk), .Q(sram_rdata_0[27]), .QN(n472) );
  DFFSSRX1_HVT sram_rdata_0_reg_26_ ( .D(1'b0), .SETB(n2490), .RSTB(N65), 
        .CLK(clk), .Q(sram_rdata_0[26]), .QN(n471) );
  DFFSSRX1_HVT sram_rdata_0_reg_25_ ( .D(1'b0), .SETB(n12200), .RSTB(N64), 
        .CLK(clk), .Q(sram_rdata_0[25]), .QN(n4701) );
  DFFSSRX1_HVT sram_rdata_0_reg_24_ ( .D(1'b0), .SETB(n2410), .RSTB(N63), 
        .CLK(clk), .Q(sram_rdata_0[24]), .QN(n469) );
  DFFSSRX1_HVT sram_rdata_0_reg_23_ ( .D(1'b0), .SETB(n2450), .RSTB(N62), 
        .CLK(clk), .Q(sram_rdata_0[23]), .QN(n468) );
  DFFSSRX1_HVT sram_rdata_0_reg_22_ ( .D(1'b0), .SETB(n2510), .RSTB(N61), 
        .CLK(clk), .Q(sram_rdata_0[22]), .QN(n467) );
  DFFSSRX1_HVT sram_rdata_0_reg_21_ ( .D(1'b0), .SETB(n2530), .RSTB(N60), 
        .CLK(clk), .Q(sram_rdata_0[21]), .QN(n466) );
  DFFSSRX1_HVT sram_rdata_0_reg_20_ ( .D(1'b0), .SETB(n2410), .RSTB(N59), 
        .CLK(clk), .Q(sram_rdata_0[20]), .QN(n465) );
  DFFSSRX1_HVT sram_rdata_0_reg_19_ ( .D(1'b0), .SETB(n2450), .RSTB(N58), 
        .CLK(clk), .Q(sram_rdata_0[19]), .QN(n464) );
  DFFSSRX1_HVT sram_rdata_0_reg_18_ ( .D(1'b0), .SETB(n12400), .RSTB(N57), 
        .CLK(clk), .Q(sram_rdata_0[18]), .QN(n463) );
  DFFSSRX1_HVT sram_rdata_0_reg_17_ ( .D(1'b0), .SETB(n2530), .RSTB(N56), 
        .CLK(clk), .Q(sram_rdata_0[17]), .QN(n462) );
  DFFSSRX1_HVT sram_rdata_0_reg_16_ ( .D(1'b0), .SETB(n13200), .RSTB(N55), 
        .CLK(clk), .Q(sram_rdata_0[16]), .QN(n461) );
  DFFSSRX1_HVT sram_rdata_0_reg_15_ ( .D(1'b0), .SETB(n2850), .RSTB(N54), 
        .CLK(clk), .Q(sram_rdata_0[15]), .QN(n4601) );
  DFFSSRX1_HVT sram_rdata_0_reg_14_ ( .D(1'b0), .SETB(n2480), .RSTB(N53), 
        .CLK(clk), .Q(sram_rdata_0[14]), .QN(n459) );
  DFFSSRX1_HVT sram_rdata_0_reg_13_ ( .D(1'b0), .SETB(n2530), .RSTB(N52), 
        .CLK(clk), .Q(sram_rdata_0[13]), .QN(n458) );
  DFFSSRX1_HVT sram_rdata_0_reg_12_ ( .D(1'b0), .SETB(n2440), .RSTB(N51), 
        .CLK(clk), .Q(sram_rdata_0[12]), .QN(n457) );
  DFFSSRX1_HVT sram_rdata_0_reg_11_ ( .D(1'b0), .SETB(n2500), .RSTB(N50), 
        .CLK(clk), .Q(sram_rdata_0[11]), .QN(n456) );
  DFFSSRX1_HVT sram_rdata_0_reg_10_ ( .D(1'b0), .SETB(n2480), .RSTB(N49), 
        .CLK(clk), .Q(sram_rdata_0[10]), .QN(n455) );
  DFFSSRX1_HVT sram_rdata_0_reg_9_ ( .D(1'b0), .SETB(n12200), .RSTB(N48), 
        .CLK(clk), .Q(sram_rdata_0[9]), .QN(n454) );
  DFFSSRX1_HVT sram_rdata_0_reg_8_ ( .D(1'b0), .SETB(n2440), .RSTB(N47), .CLK(
        clk), .Q(sram_rdata_0[8]), .QN(n453) );
  DFFSSRX1_HVT sram_rdata_0_reg_7_ ( .D(1'b0), .SETB(n2840), .RSTB(N46), .CLK(
        clk), .Q(sram_rdata_0[7]), .QN(n452) );
  DFFSSRX1_HVT sram_rdata_0_reg_6_ ( .D(1'b0), .SETB(n2480), .RSTB(N45), .CLK(
        clk), .Q(sram_rdata_0[6]), .QN(n451) );
  DFFSSRX1_HVT sram_rdata_0_reg_5_ ( .D(1'b0), .SETB(n2560), .RSTB(N44), .CLK(
        clk), .Q(sram_rdata_0[5]), .QN(n4501) );
  DFFSSRX1_HVT sram_rdata_0_reg_4_ ( .D(1'b0), .SETB(n2440), .RSTB(N43), .CLK(
        clk), .Q(sram_rdata_0[4]), .QN(n449) );
  DFFSSRX1_HVT sram_rdata_0_reg_3_ ( .D(1'b0), .SETB(n2830), .RSTB(N42), .CLK(
        clk), .Q(sram_rdata_0[3]), .QN(n448) );
  DFFSSRX1_HVT sram_rdata_0_reg_2_ ( .D(1'b0), .SETB(n12400), .RSTB(N41), 
        .CLK(clk), .Q(sram_rdata_0[2]), .QN(n447) );
  DFFSSRX1_HVT sram_rdata_0_reg_1_ ( .D(1'b0), .SETB(n2560), .RSTB(N40), .CLK(
        clk), .Q(sram_rdata_0[1]), .QN(n446) );
  DFFSSRX1_HVT sram_rdata_0_reg_0_ ( .D(1'b0), .SETB(n13400), .RSTB(N39), 
        .CLK(clk), .Q(sram_rdata_0[0]), .QN(n445) );
  DFFSSRX1_HVT sram_rdata_1_reg_31_ ( .D(1'b0), .SETB(n2530), .RSTB(N102), 
        .CLK(clk), .Q(sram_rdata_1[31]), .QN(n381) );
  DFFSSRX1_HVT sram_rdata_1_reg_30_ ( .D(1'b0), .SETB(n2420), .RSTB(N101), 
        .CLK(clk), .Q(sram_rdata_1[30]), .QN(n380) );
  DFFSSRX1_HVT sram_rdata_1_reg_29_ ( .D(1'b0), .SETB(n12400), .RSTB(N100), 
        .CLK(clk), .Q(sram_rdata_1[29]), .QN(n379) );
  DFFSSRX1_HVT sram_rdata_1_reg_28_ ( .D(1'b0), .SETB(n2490), .RSTB(N99), 
        .CLK(clk), .Q(sram_rdata_1[28]), .QN(n378) );
  DFFSSRX1_HVT sram_rdata_1_reg_27_ ( .D(1'b0), .SETB(n13400), .RSTB(N98), 
        .CLK(clk), .Q(sram_rdata_1[27]), .QN(n377) );
  DFFSSRX1_HVT sram_rdata_1_reg_26_ ( .D(1'b0), .SETB(n2420), .RSTB(N97), 
        .CLK(clk), .Q(sram_rdata_1[26]), .QN(n376) );
  DFFSSRX1_HVT sram_rdata_1_reg_25_ ( .D(1'b0), .SETB(n2450), .RSTB(N96), 
        .CLK(clk), .Q(sram_rdata_1[25]), .QN(n375) );
  DFFSSRX1_HVT sram_rdata_1_reg_24_ ( .D(1'b0), .SETB(n2480), .RSTB(N95), 
        .CLK(clk), .Q(sram_rdata_1[24]), .QN(n374) );
  DFFSSRX1_HVT sram_rdata_1_reg_23_ ( .D(1'b0), .SETB(n2540), .RSTB(N94), 
        .CLK(clk), .Q(sram_rdata_1[23]), .QN(n373) );
  DFFSSRX1_HVT sram_rdata_1_reg_22_ ( .D(1'b0), .SETB(n2440), .RSTB(N93), 
        .CLK(clk), .Q(sram_rdata_1[22]), .QN(n372) );
  DFFSSRX1_HVT sram_rdata_1_reg_21_ ( .D(1'b0), .SETB(n2450), .RSTB(N92), 
        .CLK(clk), .Q(sram_rdata_1[21]), .QN(n371) );
  DFFSSRX1_HVT sram_rdata_1_reg_20_ ( .D(1'b0), .SETB(n12400), .RSTB(N91), 
        .CLK(clk), .Q(sram_rdata_1[20]), .QN(n370) );
  DFFSSRX1_HVT sram_rdata_1_reg_19_ ( .D(1'b0), .SETB(n2540), .RSTB(N90), 
        .CLK(clk), .Q(sram_rdata_1[19]), .QN(n369) );
  DFFSSRX1_HVT sram_rdata_1_reg_18_ ( .D(1'b0), .SETB(n12300), .RSTB(N89), 
        .CLK(clk), .Q(sram_rdata_1[18]), .QN(n368) );
  DFFSSRX1_HVT sram_rdata_1_reg_17_ ( .D(1'b0), .SETB(n12200), .RSTB(N88), 
        .CLK(clk), .Q(sram_rdata_1[17]), .QN(n367) );
  DFFSSRX1_HVT sram_rdata_1_reg_16_ ( .D(1'b0), .SETB(n2490), .RSTB(N87), 
        .CLK(clk), .Q(sram_rdata_1[16]), .QN(n366) );
  DFFSSRX1_HVT sram_rdata_1_reg_15_ ( .D(1'b0), .SETB(n2560), .RSTB(N86), 
        .CLK(clk), .Q(sram_rdata_1[15]), .QN(n365) );
  DFFSSRX1_HVT sram_rdata_1_reg_14_ ( .D(1'b0), .SETB(n2410), .RSTB(N85), 
        .CLK(clk), .Q(sram_rdata_1[14]), .QN(n364) );
  DFFSSRX1_HVT sram_rdata_1_reg_13_ ( .D(1'b0), .SETB(n12400), .RSTB(N84), 
        .CLK(clk), .Q(sram_rdata_1[13]), .QN(n363) );
  DFFSSRX1_HVT sram_rdata_1_reg_12_ ( .D(1'b0), .SETB(n2490), .RSTB(N83), 
        .CLK(clk), .Q(sram_rdata_1[12]), .QN(n362) );
  DFFSSRX1_HVT sram_rdata_1_reg_11_ ( .D(1'b0), .SETB(n13400), .RSTB(N82), 
        .CLK(clk), .Q(sram_rdata_1[11]), .QN(n361) );
  DFFSSRX1_HVT sram_rdata_1_reg_10_ ( .D(1'b0), .SETB(n2410), .RSTB(N81), 
        .CLK(clk), .Q(sram_rdata_1[10]), .QN(n360) );
  DFFSSRX1_HVT sram_rdata_1_reg_9_ ( .D(1'b0), .SETB(n2450), .RSTB(N80), .CLK(
        clk), .Q(sram_rdata_1[9]), .QN(n359) );
  DFFSSRX1_HVT sram_rdata_1_reg_8_ ( .D(1'b0), .SETB(n2510), .RSTB(N79), .CLK(
        clk), .Q(sram_rdata_1[8]), .QN(n358) );
  DFFSSRX1_HVT sram_rdata_1_reg_7_ ( .D(1'b0), .SETB(n2530), .RSTB(N78), .CLK(
        clk), .Q(sram_rdata_1[7]), .QN(n357) );
  DFFSSRX1_HVT sram_rdata_1_reg_6_ ( .D(1'b0), .SETB(n2410), .RSTB(N77), .CLK(
        clk), .Q(sram_rdata_1[6]), .QN(n356) );
  DFFSSRX1_HVT sram_rdata_1_reg_5_ ( .D(1'b0), .SETB(n2450), .RSTB(N76), .CLK(
        clk), .Q(sram_rdata_1[5]), .QN(n355) );
  DFFSSRX1_HVT sram_rdata_1_reg_4_ ( .D(1'b0), .SETB(n12400), .RSTB(N75), 
        .CLK(clk), .Q(sram_rdata_1[4]), .QN(n354) );
  DFFSSRX1_HVT sram_rdata_1_reg_3_ ( .D(1'b0), .SETB(n2530), .RSTB(N74), .CLK(
        clk), .Q(sram_rdata_1[3]), .QN(n353) );
  DFFSSRX1_HVT sram_rdata_1_reg_2_ ( .D(1'b0), .SETB(n12300), .RSTB(N73), 
        .CLK(clk), .Q(sram_rdata_1[2]), .QN(n352) );
  DFFSSRX1_HVT sram_rdata_1_reg_1_ ( .D(1'b0), .SETB(n2830), .RSTB(N72), .CLK(
        clk), .Q(sram_rdata_1[1]), .QN(n351) );
  DFFSSRX1_HVT sram_rdata_1_reg_0_ ( .D(1'b0), .SETB(n2450), .RSTB(N71), .CLK(
        clk), .Q(sram_rdata_1[0]), .QN(n350) );
  DFFSSRX1_HVT sram_rdata_2_reg_31_ ( .D(1'b0), .SETB(n2480), .RSTB(N134), 
        .CLK(clk), .Q(sram_rdata_2[31]), .QN(n572) );
  DFFSSRX1_HVT sram_rdata_2_reg_30_ ( .D(1'b0), .SETB(n2540), .RSTB(N133), 
        .CLK(clk), .Q(sram_rdata_2[30]), .QN(n571) );
  DFFSSRX1_HVT sram_rdata_2_reg_29_ ( .D(1'b0), .SETB(n2440), .RSTB(N132), 
        .CLK(clk), .Q(sram_rdata_2[29]), .QN(n5701) );
  DFFSSRX1_HVT sram_rdata_2_reg_28_ ( .D(1'b0), .SETB(n2450), .RSTB(N131), 
        .CLK(clk), .Q(sram_rdata_2[28]), .QN(n569) );
  DFFSSRX1_HVT sram_rdata_2_reg_27_ ( .D(1'b0), .SETB(n13300), .RSTB(N130), 
        .CLK(clk), .Q(sram_rdata_2[27]), .QN(n568) );
  DFFSSRX1_HVT sram_rdata_2_reg_26_ ( .D(1'b0), .SETB(n2540), .RSTB(N129), 
        .CLK(clk), .Q(sram_rdata_2[26]), .QN(n567) );
  DFFSSRX1_HVT sram_rdata_2_reg_25_ ( .D(1'b0), .SETB(n12300), .RSTB(N128), 
        .CLK(clk), .Q(sram_rdata_2[25]), .QN(n566) );
  DFFSSRX1_HVT sram_rdata_2_reg_24_ ( .D(1'b0), .SETB(n12400), .RSTB(N127), 
        .CLK(clk), .Q(sram_rdata_2[24]), .QN(n565) );
  DFFSSRX1_HVT sram_rdata_2_reg_23_ ( .D(1'b0), .SETB(n2490), .RSTB(N126), 
        .CLK(clk), .Q(sram_rdata_2[23]), .QN(n564) );
  DFFSSRX1_HVT sram_rdata_2_reg_22_ ( .D(1'b0), .SETB(n2560), .RSTB(N125), 
        .CLK(clk), .Q(sram_rdata_2[22]), .QN(n563) );
  DFFSSRX1_HVT sram_rdata_2_reg_21_ ( .D(1'b0), .SETB(n2410), .RSTB(N124), 
        .CLK(clk), .Q(sram_rdata_2[21]), .QN(n562) );
  DFFSSRX1_HVT sram_rdata_2_reg_20_ ( .D(1'b0), .SETB(n12400), .RSTB(N123), 
        .CLK(clk), .Q(sram_rdata_2[20]), .QN(n561) );
  DFFSSRX1_HVT sram_rdata_2_reg_19_ ( .D(1'b0), .SETB(n2490), .RSTB(N122), 
        .CLK(clk), .Q(sram_rdata_2[19]), .QN(n5601) );
  DFFSSRX1_HVT sram_rdata_2_reg_18_ ( .D(1'b0), .SETB(n12200), .RSTB(N121), 
        .CLK(clk), .Q(sram_rdata_2[18]), .QN(n559) );
  DFFSSRX1_HVT sram_rdata_2_reg_17_ ( .D(1'b0), .SETB(n2410), .RSTB(N120), 
        .CLK(clk), .Q(sram_rdata_2[17]), .QN(n558) );
  DFFSSRX1_HVT sram_rdata_2_reg_16_ ( .D(1'b0), .SETB(n2450), .RSTB(N119), 
        .CLK(clk), .Q(sram_rdata_2[16]), .QN(n557) );
  DFFSSRX1_HVT sram_rdata_2_reg_15_ ( .D(1'b0), .SETB(n2510), .RSTB(N118), 
        .CLK(clk), .Q(sram_rdata_2[15]), .QN(n556) );
  DFFSSRX1_HVT sram_rdata_2_reg_14_ ( .D(1'b0), .SETB(n2530), .RSTB(N117), 
        .CLK(clk), .Q(sram_rdata_2[14]), .QN(n555) );
  DFFSSRX1_HVT sram_rdata_2_reg_13_ ( .D(1'b0), .SETB(n2410), .RSTB(N116), 
        .CLK(clk), .Q(sram_rdata_2[13]), .QN(n554) );
  DFFSSRX1_HVT sram_rdata_2_reg_12_ ( .D(1'b0), .SETB(n2450), .RSTB(N115), 
        .CLK(clk), .Q(sram_rdata_2[12]), .QN(n553) );
  DFFSSRX1_HVT sram_rdata_2_reg_11_ ( .D(1'b0), .SETB(n13300), .RSTB(N114), 
        .CLK(clk), .Q(sram_rdata_2[11]), .QN(n552) );
  DFFSSRX1_HVT sram_rdata_2_reg_10_ ( .D(1'b0), .SETB(n2530), .RSTB(N113), 
        .CLK(clk), .Q(sram_rdata_2[10]), .QN(n551) );
  DFFSSRX1_HVT sram_rdata_2_reg_9_ ( .D(1'b0), .SETB(n12300), .RSTB(N112), 
        .CLK(clk), .Q(sram_rdata_2[9]), .QN(n5501) );
  DFFSSRX1_HVT sram_rdata_2_reg_8_ ( .D(1'b0), .SETB(n2840), .RSTB(N111), 
        .CLK(clk), .Q(sram_rdata_2[8]), .QN(n549) );
  DFFSSRX1_HVT sram_rdata_2_reg_7_ ( .D(1'b0), .SETB(n2480), .RSTB(N110), 
        .CLK(clk), .Q(sram_rdata_2[7]), .QN(n548) );
  DFFSSRX1_HVT sram_rdata_2_reg_6_ ( .D(1'b0), .SETB(n2530), .RSTB(N109), 
        .CLK(clk), .Q(sram_rdata_2[6]), .QN(n547) );
  DFFSSRX1_HVT sram_rdata_2_reg_5_ ( .D(1'b0), .SETB(n2440), .RSTB(N108), 
        .CLK(clk), .Q(sram_rdata_2[5]), .QN(n546) );
  DFFSSRX1_HVT sram_rdata_2_reg_4_ ( .D(1'b0), .SETB(n12200), .RSTB(N107), 
        .CLK(clk), .Q(sram_rdata_2[4]), .QN(n545) );
  DFFSSRX1_HVT sram_rdata_2_reg_3_ ( .D(1'b0), .SETB(n2480), .RSTB(N106), 
        .CLK(clk), .Q(sram_rdata_2[3]), .QN(n544) );
  DFFSSRX1_HVT sram_rdata_2_reg_2_ ( .D(1'b0), .SETB(n12200), .RSTB(N105), 
        .CLK(clk), .Q(sram_rdata_2[2]), .QN(n543) );
  DFFSSRX1_HVT sram_rdata_2_reg_1_ ( .D(1'b0), .SETB(n2440), .RSTB(N104), 
        .CLK(clk), .Q(sram_rdata_2[1]), .QN(n542) );
  DFFSSRX1_HVT sram_rdata_2_reg_0_ ( .D(1'b0), .SETB(n13200), .RSTB(N103), 
        .CLK(clk), .Q(sram_rdata_2[0]), .QN(n541) );
  DFFSSRX1_HVT sram_rdata_3_reg_31_ ( .D(1'b0), .SETB(n2410), .RSTB(N166), 
        .CLK(clk), .Q(sram_rdata_3[31]), .QN(n444) );
  DFFSSRX1_HVT sram_rdata_3_reg_30_ ( .D(1'b0), .SETB(n2500), .RSTB(N165), 
        .CLK(clk), .Q(sram_rdata_3[30]), .QN(n443) );
  DFFSSRX1_HVT sram_rdata_3_reg_29_ ( .D(1'b0), .SETB(n12400), .RSTB(N164), 
        .CLK(clk), .Q(sram_rdata_3[29]), .QN(n442) );
  DFFSSRX1_HVT sram_rdata_3_reg_28_ ( .D(1'b0), .SETB(n2540), .RSTB(N163), 
        .CLK(clk), .Q(sram_rdata_3[28]), .QN(n441) );
  DFFSSRX1_HVT sram_rdata_3_reg_27_ ( .D(1'b0), .SETB(n13200), .RSTB(N162), 
        .CLK(clk), .Q(sram_rdata_3[27]), .QN(n4401) );
  DFFSSRX1_HVT sram_rdata_3_reg_26_ ( .D(1'b0), .SETB(n2850), .RSTB(N161), 
        .CLK(clk), .Q(sram_rdata_3[26]), .QN(n439) );
  DFFSSRX1_HVT sram_rdata_3_reg_25_ ( .D(1'b0), .SETB(n2490), .RSTB(N160), 
        .CLK(clk), .Q(sram_rdata_3[25]), .QN(n438) );
  DFFSSRX1_HVT sram_rdata_3_reg_24_ ( .D(1'b0), .SETB(n2530), .RSTB(N159), 
        .CLK(clk), .Q(sram_rdata_3[24]), .QN(n437) );
  DFFSSRX1_HVT sram_rdata_3_reg_23_ ( .D(1'b0), .SETB(n2420), .RSTB(N158), 
        .CLK(clk), .Q(sram_rdata_3[23]), .QN(n436) );
  DFFSSRX1_HVT sram_rdata_3_reg_22_ ( .D(1'b0), .SETB(n12300), .RSTB(N157), 
        .CLK(clk), .Q(sram_rdata_3[22]), .QN(n435) );
  DFFSSRX1_HVT sram_rdata_3_reg_21_ ( .D(1'b0), .SETB(n2490), .RSTB(N156), 
        .CLK(clk), .Q(sram_rdata_3[21]), .QN(n434) );
  DFFSSRX1_HVT sram_rdata_3_reg_20_ ( .D(1'b0), .SETB(n12200), .RSTB(N155), 
        .CLK(clk), .Q(sram_rdata_3[20]), .QN(n433) );
  DFFSSRX1_HVT sram_rdata_3_reg_19_ ( .D(1'b0), .SETB(n2420), .RSTB(N154), 
        .CLK(clk), .Q(sram_rdata_3[19]), .QN(n432) );
  DFFSSRX1_HVT sram_rdata_3_reg_18_ ( .D(1'b0), .SETB(n2450), .RSTB(N153), 
        .CLK(clk), .Q(sram_rdata_3[18]), .QN(n431) );
  DFFSSRX1_HVT sram_rdata_3_reg_17_ ( .D(1'b0), .SETB(n2480), .RSTB(N152), 
        .CLK(clk), .Q(sram_rdata_3[17]), .QN(n4301) );
  DFFSSRX1_HVT sram_rdata_3_reg_16_ ( .D(1'b0), .SETB(n2540), .RSTB(N151), 
        .CLK(clk), .Q(sram_rdata_3[16]), .QN(n429) );
  DFFSSRX1_HVT sram_rdata_3_reg_15_ ( .D(1'b0), .SETB(n2440), .RSTB(N150), 
        .CLK(clk), .Q(sram_rdata_3[15]), .QN(n428) );
  DFFSSRX1_HVT sram_rdata_3_reg_14_ ( .D(1'b0), .SETB(n2450), .RSTB(N149), 
        .CLK(clk), .Q(sram_rdata_3[14]), .QN(n427) );
  DFFSSRX1_HVT sram_rdata_3_reg_13_ ( .D(1'b0), .SETB(n12400), .RSTB(N148), 
        .CLK(clk), .Q(sram_rdata_3[13]), .QN(n426) );
  DFFSSRX1_HVT sram_rdata_3_reg_12_ ( .D(1'b0), .SETB(n2540), .RSTB(N147), 
        .CLK(clk), .Q(sram_rdata_3[12]), .QN(n425) );
  DFFSSRX1_HVT sram_rdata_3_reg_11_ ( .D(1'b0), .SETB(n13200), .RSTB(N146), 
        .CLK(clk), .Q(sram_rdata_3[11]), .QN(n424) );
  DFFSSRX1_HVT sram_rdata_3_reg_10_ ( .D(1'b0), .SETB(n2500), .RSTB(N145), 
        .CLK(clk), .Q(sram_rdata_3[10]), .QN(n423) );
  DFFSSRX1_HVT sram_rdata_3_reg_9_ ( .D(1'b0), .SETB(n2490), .RSTB(N144), 
        .CLK(clk), .Q(sram_rdata_3[9]), .QN(n422) );
  DFFSSRX1_HVT sram_rdata_3_reg_8_ ( .D(1'b0), .SETB(n2560), .RSTB(N143), 
        .CLK(clk), .Q(sram_rdata_3[8]), .QN(n421) );
  DFFSSRX1_HVT sram_rdata_3_reg_7_ ( .D(1'b0), .SETB(n2410), .RSTB(N142), 
        .CLK(clk), .Q(sram_rdata_3[7]), .QN(n4201) );
  DFFSSRX1_HVT sram_rdata_3_reg_6_ ( .D(1'b0), .SETB(n2550), .RSTB(N141), 
        .CLK(clk), .Q(sram_rdata_3[6]), .QN(n419) );
  DFFSSRX1_HVT sram_rdata_3_reg_5_ ( .D(1'b0), .SETB(n2490), .RSTB(N140), 
        .CLK(clk), .Q(sram_rdata_3[5]), .QN(n418) );
  DFFSSRX1_HVT sram_rdata_3_reg_4_ ( .D(1'b0), .SETB(n12200), .RSTB(N139), 
        .CLK(clk), .Q(sram_rdata_3[4]), .QN(n417) );
  DFFSSRX1_HVT sram_rdata_3_reg_3_ ( .D(1'b0), .SETB(n2410), .RSTB(N138), 
        .CLK(clk), .Q(sram_rdata_3[3]), .QN(n416) );
  DFFSSRX1_HVT sram_rdata_3_reg_2_ ( .D(1'b0), .SETB(n2450), .RSTB(N137), 
        .CLK(clk), .Q(sram_rdata_3[2]), .QN(n415) );
  DFFSSRX1_HVT sram_rdata_3_reg_1_ ( .D(1'b0), .SETB(n2510), .RSTB(N136), 
        .CLK(clk), .Q(sram_rdata_3[1]), .QN(n414) );
  DFFSSRX1_HVT sram_rdata_3_reg_0_ ( .D(1'b0), .SETB(n2490), .RSTB(N135), 
        .CLK(clk), .Q(sram_rdata_3[0]), .QN(n382) );
  DFFSSRX1_HVT sram_rdata_4_reg_31_ ( .D(1'b0), .SETB(n12400), .RSTB(N198), 
        .CLK(clk), .Q(sram_rdata_4[31]), .QN(n349) );
  DFFSSRX1_HVT sram_rdata_4_reg_30_ ( .D(1'b0), .SETB(n2560), .RSTB(N197), 
        .CLK(clk), .Q(sram_rdata_4[30]), .QN(n348) );
  DFFSSRX1_HVT sram_rdata_4_reg_29_ ( .D(1'b0), .SETB(n12300), .RSTB(N196), 
        .CLK(clk), .Q(sram_rdata_4[29]), .QN(n347) );
  DFFSSRX1_HVT sram_rdata_4_reg_28_ ( .D(1'b0), .SETB(n12200), .RSTB(N195), 
        .CLK(clk), .Q(sram_rdata_4[28]), .QN(n3460) );
  DFFSSRX1_HVT sram_rdata_4_reg_27_ ( .D(1'b0), .SETB(n2510), .RSTB(N194), 
        .CLK(clk), .Q(sram_rdata_4[27]), .QN(n345) );
  DFFSSRX1_HVT sram_rdata_4_reg_26_ ( .D(1'b0), .SETB(n2560), .RSTB(N193), 
        .CLK(clk), .Q(sram_rdata_4[26]), .QN(n344) );
  DFFSSRX1_HVT sram_rdata_4_reg_25_ ( .D(1'b0), .SETB(n2420), .RSTB(N192), 
        .CLK(clk), .Q(sram_rdata_4[25]), .QN(n343) );
  DFFSSRX1_HVT sram_rdata_4_reg_24_ ( .D(1'b0), .SETB(n12300), .RSTB(N191), 
        .CLK(clk), .Q(sram_rdata_4[24]), .QN(n342) );
  DFFSSRX1_HVT sram_rdata_4_reg_23_ ( .D(1'b0), .SETB(n2510), .RSTB(N190), 
        .CLK(clk), .Q(sram_rdata_4[23]), .QN(n341) );
  DFFSSRX1_HVT sram_rdata_4_reg_22_ ( .D(1'b0), .SETB(n13400), .RSTB(N189), 
        .CLK(clk), .Q(sram_rdata_4[22]), .QN(n340) );
  DFFSSRX1_HVT sram_rdata_4_reg_21_ ( .D(1'b0), .SETB(n2420), .RSTB(N188), 
        .CLK(clk), .Q(sram_rdata_4[21]), .QN(n339) );
  DFFSSRX1_HVT sram_rdata_4_reg_20_ ( .D(1'b0), .SETB(n2830), .RSTB(N187), 
        .CLK(clk), .Q(sram_rdata_4[20]), .QN(n338) );
  DFFSSRX1_HVT sram_rdata_4_reg_19_ ( .D(1'b0), .SETB(n2510), .RSTB(N186), 
        .CLK(clk), .Q(sram_rdata_4[19]), .QN(n337) );
  DFFSSRX1_HVT sram_rdata_4_reg_18_ ( .D(1'b0), .SETB(n2540), .RSTB(N185), 
        .CLK(clk), .Q(sram_rdata_4[18]), .QN(n336) );
  DFFSSRX1_HVT sram_rdata_4_reg_17_ ( .D(1'b0), .SETB(n2410), .RSTB(N184), 
        .CLK(clk), .Q(sram_rdata_4[17]), .QN(n335) );
  DFFSSRX1_HVT sram_rdata_4_reg_16_ ( .D(1'b0), .SETB(n2430), .RSTB(N183), 
        .CLK(clk), .Q(sram_rdata_4[16]), .QN(n334) );
  DFFSSRX1_HVT sram_rdata_4_reg_15_ ( .D(1'b0), .SETB(n12400), .RSTB(N182), 
        .CLK(clk), .Q(sram_rdata_4[15]), .QN(n333) );
  DFFSSRX1_HVT sram_rdata_4_reg_14_ ( .D(1'b0), .SETB(n2540), .RSTB(N181), 
        .CLK(clk), .Q(sram_rdata_4[14]), .QN(n332) );
  DFFSSRX1_HVT sram_rdata_4_reg_13_ ( .D(1'b0), .SETB(n12300), .RSTB(N180), 
        .CLK(clk), .Q(sram_rdata_4[13]), .QN(n331) );
  DFFSSRX1_HVT sram_rdata_4_reg_12_ ( .D(1'b0), .SETB(n2830), .RSTB(N179), 
        .CLK(clk), .Q(sram_rdata_4[12]), .QN(n330) );
  DFFSSRX1_HVT sram_rdata_4_reg_11_ ( .D(1'b0), .SETB(n2490), .RSTB(N178), 
        .CLK(clk), .Q(sram_rdata_4[11]), .QN(n329) );
  DFFSSRX1_HVT sram_rdata_4_reg_10_ ( .D(1'b0), .SETB(n2530), .RSTB(N177), 
        .CLK(clk), .Q(sram_rdata_4[10]), .QN(n328) );
  DFFSSRX1_HVT sram_rdata_4_reg_9_ ( .D(1'b0), .SETB(n2420), .RSTB(N176), 
        .CLK(clk), .Q(sram_rdata_4[9]), .QN(n327) );
  DFFSSRX1_HVT sram_rdata_4_reg_8_ ( .D(1'b0), .SETB(n2430), .RSTB(N175), 
        .CLK(clk), .Q(sram_rdata_4[8]), .QN(n3260) );
  DFFSSRX1_HVT sram_rdata_4_reg_7_ ( .D(1'b0), .SETB(n2490), .RSTB(N174), 
        .CLK(clk), .Q(sram_rdata_4[7]), .QN(n3250) );
  DFFSSRX1_HVT sram_rdata_4_reg_6_ ( .D(1'b0), .SETB(n13400), .RSTB(N173), 
        .CLK(clk), .Q(sram_rdata_4[6]), .QN(n3240) );
  DFFSSRX1_HVT sram_rdata_4_reg_5_ ( .D(1'b0), .SETB(n2420), .RSTB(N172), 
        .CLK(clk), .Q(sram_rdata_4[5]), .QN(n3230) );
  DFFSSRX1_HVT sram_rdata_4_reg_4_ ( .D(1'b0), .SETB(n2450), .RSTB(N171), 
        .CLK(clk), .Q(sram_rdata_4[4]), .QN(n3220) );
  DFFSSRX1_HVT sram_rdata_4_reg_3_ ( .D(1'b0), .SETB(n2480), .RSTB(N170), 
        .CLK(clk), .Q(sram_rdata_4[3]), .QN(n3210) );
  DFFSSRX1_HVT sram_rdata_4_reg_2_ ( .D(1'b0), .SETB(n2540), .RSTB(N169), 
        .CLK(clk), .Q(sram_rdata_4[2]), .QN(n3200) );
  DFFSSRX1_HVT sram_rdata_4_reg_1_ ( .D(1'b0), .SETB(n2440), .RSTB(N168), 
        .CLK(clk), .Q(sram_rdata_4[1]), .QN(n3190) );
  DFFSSRX1_HVT sram_rdata_4_reg_0_ ( .D(1'b0), .SETB(n2420), .RSTB(N167), 
        .CLK(clk), .Q(sram_rdata_4[0]), .QN(n3180) );
  DFFSSRX1_HVT sram_rdata_5_reg_31_ ( .D(1'b0), .SETB(n12300), .RSTB(N230), 
        .CLK(clk), .Q(sram_rdata_5[31]), .QN(n5401) );
  DFFSSRX1_HVT sram_rdata_5_reg_30_ ( .D(1'b0), .SETB(n2510), .RSTB(N229), 
        .CLK(clk), .Q(sram_rdata_5[30]), .QN(n539) );
  DFFSSRX1_HVT sram_rdata_5_reg_29_ ( .D(1'b0), .SETB(n12200), .RSTB(N228), 
        .CLK(clk), .Q(sram_rdata_5[29]), .QN(n538) );
  DFFSSRX1_HVT sram_rdata_5_reg_28_ ( .D(1'b0), .SETB(n2420), .RSTB(N227), 
        .CLK(clk), .Q(sram_rdata_5[28]), .QN(n537) );
  DFFSSRX1_HVT sram_rdata_5_reg_27_ ( .D(1'b0), .SETB(n2840), .RSTB(N226), 
        .CLK(clk), .Q(sram_rdata_5[27]), .QN(n536) );
  DFFSSRX1_HVT sram_rdata_5_reg_26_ ( .D(1'b0), .SETB(n2510), .RSTB(N225), 
        .CLK(clk), .Q(sram_rdata_5[26]), .QN(n535) );
  DFFSSRX1_HVT sram_rdata_5_reg_25_ ( .D(1'b0), .SETB(n2540), .RSTB(N224), 
        .CLK(clk), .Q(sram_rdata_5[25]), .QN(n534) );
  DFFSSRX1_HVT sram_rdata_5_reg_24_ ( .D(1'b0), .SETB(n2410), .RSTB(N223), 
        .CLK(clk), .Q(sram_rdata_5[24]), .QN(n533) );
  DFFSSRX1_HVT sram_rdata_5_reg_23_ ( .D(1'b0), .SETB(n13200), .RSTB(N222), 
        .CLK(clk), .Q(sram_rdata_5[23]), .QN(n532) );
  DFFSSRX1_HVT sram_rdata_5_reg_22_ ( .D(1'b0), .SETB(n13300), .RSTB(N221), 
        .CLK(clk), .Q(sram_rdata_5[22]), .QN(n531) );
  DFFSSRX1_HVT sram_rdata_5_reg_21_ ( .D(1'b0), .SETB(n2540), .RSTB(N220), 
        .CLK(clk), .Q(sram_rdata_5[21]), .QN(n5301) );
  DFFSSRX1_HVT sram_rdata_5_reg_20_ ( .D(1'b0), .SETB(n12300), .RSTB(N219), 
        .CLK(clk), .Q(sram_rdata_5[20]), .QN(n529) );
  DFFSSRX1_HVT sram_rdata_5_reg_19_ ( .D(1'b0), .SETB(n2840), .RSTB(N218), 
        .CLK(clk), .Q(sram_rdata_5[19]), .QN(n528) );
  DFFSSRX1_HVT sram_rdata_5_reg_18_ ( .D(1'b0), .SETB(n2490), .RSTB(N217), 
        .CLK(clk), .Q(sram_rdata_5[18]), .QN(n527) );
  DFFSSRX1_HVT sram_rdata_5_reg_17_ ( .D(1'b0), .SETB(n2530), .RSTB(N216), 
        .CLK(clk), .Q(sram_rdata_5[17]), .QN(n526) );
  DFFSSRX1_HVT sram_rdata_5_reg_16_ ( .D(1'b0), .SETB(n2420), .RSTB(N215), 
        .CLK(clk), .Q(sram_rdata_5[16]), .QN(n525) );
  DFFSSRX1_HVT sram_rdata_5_reg_15_ ( .D(1'b0), .SETB(n2840), .RSTB(N214), 
        .CLK(clk), .Q(sram_rdata_5[15]), .QN(n524) );
  DFFSSRX1_HVT sram_rdata_5_reg_14_ ( .D(1'b0), .SETB(n2490), .RSTB(N213), 
        .CLK(clk), .Q(sram_rdata_5[14]), .QN(n523) );
  DFFSSRX1_HVT sram_rdata_5_reg_13_ ( .D(1'b0), .SETB(n12200), .RSTB(N212), 
        .CLK(clk), .Q(sram_rdata_5[13]), .QN(n522) );
  DFFSSRX1_HVT sram_rdata_5_reg_12_ ( .D(1'b0), .SETB(n2420), .RSTB(N211), 
        .CLK(clk), .Q(sram_rdata_5[12]), .QN(n521) );
  DFFSSRX1_HVT sram_rdata_5_reg_11_ ( .D(1'b0), .SETB(n2450), .RSTB(N210), 
        .CLK(clk), .Q(sram_rdata_5[11]), .QN(n5201) );
  DFFSSRX1_HVT sram_rdata_5_reg_10_ ( .D(1'b0), .SETB(n2480), .RSTB(N209), 
        .CLK(clk), .Q(sram_rdata_5[10]), .QN(n519) );
  DFFSSRX1_HVT sram_rdata_5_reg_9_ ( .D(1'b0), .SETB(n2540), .RSTB(N208), 
        .CLK(clk), .Q(sram_rdata_5[9]), .QN(n518) );
  DFFSSRX1_HVT sram_rdata_5_reg_8_ ( .D(1'b0), .SETB(n2440), .RSTB(N207), 
        .CLK(clk), .Q(sram_rdata_5[8]), .QN(n517) );
  DFFSSRX1_HVT sram_rdata_5_reg_7_ ( .D(1'b0), .SETB(n2450), .RSTB(N206), 
        .CLK(clk), .Q(sram_rdata_5[7]), .QN(n516) );
  DFFSSRX1_HVT sram_rdata_5_reg_6_ ( .D(1'b0), .SETB(n13300), .RSTB(N205), 
        .CLK(clk), .Q(sram_rdata_5[6]), .QN(n515) );
  DFFSSRX1_HVT sram_rdata_5_reg_5_ ( .D(1'b0), .SETB(n2540), .RSTB(N204), 
        .CLK(clk), .Q(sram_rdata_5[5]), .QN(n514) );
  DFFSSRX1_HVT sram_rdata_5_reg_4_ ( .D(1'b0), .SETB(n12300), .RSTB(N203), 
        .CLK(clk), .Q(sram_rdata_5[4]), .QN(n513) );
  DFFSSRX1_HVT sram_rdata_5_reg_3_ ( .D(1'b0), .SETB(n2430), .RSTB(N202), 
        .CLK(clk), .Q(sram_rdata_5[3]), .QN(n512) );
  DFFSSRX1_HVT sram_rdata_5_reg_2_ ( .D(1'b0), .SETB(n2490), .RSTB(N201), 
        .CLK(clk), .Q(sram_rdata_5[2]), .QN(n511) );
  DFFSSRX1_HVT sram_rdata_5_reg_1_ ( .D(1'b0), .SETB(n2560), .RSTB(N200), 
        .CLK(clk), .Q(sram_rdata_5[1]), .QN(n5101) );
  DFFSSRX1_HVT sram_rdata_5_reg_0_ ( .D(1'b0), .SETB(n2540), .RSTB(N199), 
        .CLK(clk), .Q(sram_rdata_5[0]), .QN(n478) );
  DFFSSRX1_HVT sram_rdata_6_reg_31_ ( .D(1'b0), .SETB(n2410), .RSTB(N262), 
        .CLK(clk), .Q(sram_rdata_6[31]), .QN(n509) );
  DFFSSRX1_HVT sram_rdata_6_reg_30_ ( .D(1'b0), .SETB(n2450), .RSTB(N261), 
        .CLK(clk), .Q(sram_rdata_6[30]), .QN(n508) );
  DFFSSRX1_HVT sram_rdata_6_reg_29_ ( .D(1'b0), .SETB(n2510), .RSTB(N260), 
        .CLK(clk), .Q(sram_rdata_6[29]), .QN(n507) );
  DFFSSRX1_HVT sram_rdata_6_reg_28_ ( .D(1'b0), .SETB(n2530), .RSTB(N259), 
        .CLK(clk), .Q(sram_rdata_6[28]), .QN(n506) );
  DFFSSRX1_HVT sram_rdata_6_reg_27_ ( .D(1'b0), .SETB(n2410), .RSTB(N258), 
        .CLK(clk), .Q(sram_rdata_6[27]), .QN(n505) );
  DFFSSRX1_HVT sram_rdata_6_reg_26_ ( .D(1'b0), .SETB(n2450), .RSTB(N257), 
        .CLK(clk), .Q(sram_rdata_6[26]), .QN(n504) );
  DFFSSRX1_HVT sram_rdata_6_reg_25_ ( .D(1'b0), .SETB(n12400), .RSTB(N256), 
        .CLK(clk), .Q(sram_rdata_6[25]), .QN(n503) );
  DFFSSRX1_HVT sram_rdata_6_reg_24_ ( .D(1'b0), .SETB(n2530), .RSTB(N255), 
        .CLK(clk), .Q(sram_rdata_6[24]), .QN(n502) );
  DFFSSRX1_HVT sram_rdata_6_reg_23_ ( .D(1'b0), .SETB(n12300), .RSTB(N254), 
        .CLK(clk), .Q(sram_rdata_6[23]), .QN(n501) );
  DFFSSRX1_HVT sram_rdata_6_reg_22_ ( .D(1'b0), .SETB(n2830), .RSTB(N253), 
        .CLK(clk), .Q(sram_rdata_6[22]), .QN(n5001) );
  DFFSSRX1_HVT sram_rdata_6_reg_21_ ( .D(1'b0), .SETB(n2480), .RSTB(N252), 
        .CLK(clk), .Q(sram_rdata_6[21]), .QN(n499) );
  DFFSSRX1_HVT sram_rdata_6_reg_20_ ( .D(1'b0), .SETB(n2530), .RSTB(N251), 
        .CLK(clk), .Q(sram_rdata_6[20]), .QN(n498) );
  DFFSSRX1_HVT sram_rdata_6_reg_19_ ( .D(1'b0), .SETB(n2440), .RSTB(N250), 
        .CLK(clk), .Q(sram_rdata_6[19]), .QN(n497) );
  DFFSSRX1_HVT sram_rdata_6_reg_18_ ( .D(1'b0), .SETB(n12200), .RSTB(N249), 
        .CLK(clk), .Q(sram_rdata_6[18]), .QN(n496) );
  DFFSSRX1_HVT sram_rdata_6_reg_17_ ( .D(1'b0), .SETB(n2480), .RSTB(N248), 
        .CLK(clk), .Q(sram_rdata_6[17]), .QN(n495) );
  DFFSSRX1_HVT sram_rdata_6_reg_16_ ( .D(1'b0), .SETB(n13400), .RSTB(N247), 
        .CLK(clk), .Q(sram_rdata_6[16]), .QN(n494) );
  DFFSSRX1_HVT sram_rdata_6_reg_15_ ( .D(1'b0), .SETB(n2440), .RSTB(N246), 
        .CLK(clk), .Q(sram_rdata_6[15]), .QN(n493) );
  DFFSSRX1_HVT sram_rdata_6_reg_14_ ( .D(1'b0), .SETB(n2850), .RSTB(N245), 
        .CLK(clk), .Q(sram_rdata_6[14]), .QN(n492) );
  DFFSSRX1_HVT sram_rdata_6_reg_13_ ( .D(1'b0), .SETB(n2480), .RSTB(N244), 
        .CLK(clk), .Q(sram_rdata_6[13]), .QN(n491) );
  DFFSSRX1_HVT sram_rdata_6_reg_12_ ( .D(1'b0), .SETB(n2560), .RSTB(N243), 
        .CLK(clk), .Q(sram_rdata_6[12]), .QN(n4901) );
  DFFSSRX1_HVT sram_rdata_6_reg_11_ ( .D(1'b0), .SETB(n2440), .RSTB(N242), 
        .CLK(clk), .Q(sram_rdata_6[11]), .QN(n489) );
  DFFSSRX1_HVT sram_rdata_6_reg_10_ ( .D(1'b0), .SETB(n2850), .RSTB(N241), 
        .CLK(clk), .Q(sram_rdata_6[10]), .QN(n488) );
  DFFSSRX1_HVT sram_rdata_6_reg_9_ ( .D(1'b0), .SETB(n12400), .RSTB(N240), 
        .CLK(clk), .Q(sram_rdata_6[9]), .QN(n487) );
  DFFSSRX1_HVT sram_rdata_6_reg_8_ ( .D(1'b0), .SETB(n2560), .RSTB(N239), 
        .CLK(clk), .Q(sram_rdata_6[8]), .QN(n486) );
  DFFSSRX1_HVT sram_rdata_6_reg_7_ ( .D(1'b0), .SETB(n12300), .RSTB(N238), 
        .CLK(clk), .Q(sram_rdata_6[7]), .QN(n485) );
  DFFSSRX1_HVT sram_rdata_6_reg_6_ ( .D(1'b0), .SETB(n13200), .RSTB(N237), 
        .CLK(clk), .Q(sram_rdata_6[6]), .QN(n484) );
  DFFSSRX1_HVT sram_rdata_6_reg_5_ ( .D(1'b0), .SETB(n2510), .RSTB(N236), 
        .CLK(clk), .Q(sram_rdata_6[5]), .QN(n483) );
  DFFSSRX1_HVT sram_rdata_6_reg_4_ ( .D(1'b0), .SETB(n2560), .RSTB(N235), 
        .CLK(clk), .Q(sram_rdata_6[4]), .QN(n482) );
  DFFSSRX1_HVT sram_rdata_6_reg_3_ ( .D(1'b0), .SETB(n2420), .RSTB(N234), 
        .CLK(clk), .Q(sram_rdata_6[3]), .QN(n481) );
  DFFSSRX1_HVT sram_rdata_6_reg_2_ ( .D(1'b0), .SETB(n2550), .RSTB(N233), 
        .CLK(clk), .Q(sram_rdata_6[2]), .QN(n4801) );
  DFFSSRX1_HVT sram_rdata_6_reg_1_ ( .D(1'b0), .SETB(n2510), .RSTB(N232), 
        .CLK(clk), .Q(sram_rdata_6[1]), .QN(n479) );
  DFFSSRX1_HVT sram_rdata_6_reg_0_ ( .D(1'b0), .SETB(n12200), .RSTB(N231), 
        .CLK(clk), .Q(sram_rdata_6[0]), .QN(n477) );
  DFFSSRX1_HVT sram_rdata_7_reg_31_ ( .D(1'b0), .SETB(n2530), .RSTB(N294), 
        .CLK(clk), .Q(sram_rdata_7[31]), .QN(n413) );
  DFFSSRX1_HVT sram_rdata_7_reg_30_ ( .D(1'b0), .SETB(n12300), .RSTB(N293), 
        .CLK(clk), .Q(sram_rdata_7[30]), .QN(n412) );
  DFFSSRX1_HVT sram_rdata_7_reg_29_ ( .D(1'b0), .SETB(n2840), .RSTB(N292), 
        .CLK(clk), .Q(sram_rdata_7[29]), .QN(n411) );
  DFFSSRX1_HVT sram_rdata_7_reg_28_ ( .D(1'b0), .SETB(n2480), .RSTB(N291), 
        .CLK(clk), .Q(sram_rdata_7[28]), .QN(n4101) );
  DFFSSRX1_HVT sram_rdata_7_reg_27_ ( .D(1'b0), .SETB(n2530), .RSTB(N290), 
        .CLK(clk), .Q(sram_rdata_7[27]), .QN(n409) );
  DFFSSRX1_HVT sram_rdata_7_reg_26_ ( .D(1'b0), .SETB(n2440), .RSTB(N289), 
        .CLK(clk), .Q(sram_rdata_7[26]), .QN(n408) );
  DFFSSRX1_HVT sram_rdata_7_reg_25_ ( .D(1'b0), .SETB(n12200), .RSTB(N288), 
        .CLK(clk), .Q(sram_rdata_7[25]), .QN(n407) );
  DFFSSRX1_HVT sram_rdata_7_reg_24_ ( .D(1'b0), .SETB(n2480), .RSTB(N287), 
        .CLK(clk), .Q(sram_rdata_7[24]), .QN(n406) );
  DFFSSRX1_HVT sram_rdata_7_reg_23_ ( .D(1'b0), .SETB(n12200), .RSTB(N286), 
        .CLK(clk), .Q(sram_rdata_7[23]), .QN(n405) );
  DFFSSRX1_HVT sram_rdata_7_reg_22_ ( .D(1'b0), .SETB(n2440), .RSTB(N285), 
        .CLK(clk), .Q(sram_rdata_7[22]), .QN(n404) );
  DFFSSRX1_HVT sram_rdata_7_reg_21_ ( .D(1'b0), .SETB(n2830), .RSTB(N284), 
        .CLK(clk), .Q(sram_rdata_7[21]), .QN(n403) );
  DFFSSRX1_HVT sram_rdata_7_reg_20_ ( .D(1'b0), .SETB(n2480), .RSTB(N283), 
        .CLK(clk), .Q(sram_rdata_7[20]), .QN(n402) );
  DFFSSRX1_HVT sram_rdata_7_reg_19_ ( .D(1'b0), .SETB(n2560), .RSTB(N282), 
        .CLK(clk), .Q(sram_rdata_7[19]), .QN(n401) );
  DFFSSRX1_HVT sram_rdata_7_reg_18_ ( .D(1'b0), .SETB(n2440), .RSTB(N281), 
        .CLK(clk), .Q(sram_rdata_7[18]), .QN(n4001) );
  DFFSSRX1_HVT sram_rdata_7_reg_17_ ( .D(1'b0), .SETB(n2840), .RSTB(N280), 
        .CLK(clk), .Q(sram_rdata_7[17]), .QN(n399) );
  DFFSSRX1_HVT sram_rdata_7_reg_16_ ( .D(1'b0), .SETB(n13300), .RSTB(N279), 
        .CLK(clk), .Q(sram_rdata_7[16]), .QN(n398) );
  DFFSSRX1_HVT sram_rdata_7_reg_15_ ( .D(1'b0), .SETB(n2560), .RSTB(N278), 
        .CLK(clk), .Q(sram_rdata_7[15]), .QN(n397) );
  DFFSSRX1_HVT sram_rdata_7_reg_14_ ( .D(1'b0), .SETB(n12300), .RSTB(N277), 
        .CLK(clk), .Q(sram_rdata_7[14]), .QN(n396) );
  DFFSSRX1_HVT sram_rdata_7_reg_13_ ( .D(1'b0), .SETB(n13300), .RSTB(N276), 
        .CLK(clk), .Q(sram_rdata_7[13]), .QN(n395) );
  DFFSSRX1_HVT sram_rdata_7_reg_12_ ( .D(1'b0), .SETB(n2510), .RSTB(N275), 
        .CLK(clk), .Q(sram_rdata_7[12]), .QN(n394) );
  DFFSSRX1_HVT sram_rdata_7_reg_11_ ( .D(1'b0), .SETB(n2560), .RSTB(N274), 
        .CLK(clk), .Q(sram_rdata_7[11]), .QN(n393) );
  DFFSSRX1_HVT sram_rdata_7_reg_10_ ( .D(1'b0), .SETB(n2420), .RSTB(N273), 
        .CLK(clk), .Q(sram_rdata_7[10]), .QN(n392) );
  DFFSSRX1_HVT sram_rdata_7_reg_9_ ( .D(1'b0), .SETB(n12300), .RSTB(N272), 
        .CLK(clk), .Q(sram_rdata_7[9]), .QN(n391) );
  DFFSSRX1_HVT sram_rdata_7_reg_8_ ( .D(1'b0), .SETB(n2510), .RSTB(N271), 
        .CLK(clk), .Q(sram_rdata_7[8]), .QN(n3901) );
  DFFSSRX1_HVT sram_rdata_7_reg_7_ ( .D(1'b0), .SETB(n12200), .RSTB(N270), 
        .CLK(clk), .Q(sram_rdata_7[7]), .QN(n389) );
  DFFSSRX1_HVT sram_rdata_7_reg_6_ ( .D(1'b0), .SETB(n2420), .RSTB(N269), 
        .CLK(clk), .Q(sram_rdata_7[6]), .QN(n388) );
  DFFSSRX1_HVT sram_rdata_7_reg_5_ ( .D(1'b0), .SETB(n2840), .RSTB(N268), 
        .CLK(clk), .Q(sram_rdata_7[5]), .QN(n387) );
  DFFSSRX1_HVT sram_rdata_7_reg_4_ ( .D(1'b0), .SETB(n2510), .RSTB(N267), 
        .CLK(clk), .Q(sram_rdata_7[4]), .QN(n386) );
  DFFSSRX1_HVT sram_rdata_7_reg_3_ ( .D(1'b0), .SETB(n2540), .RSTB(N266), 
        .CLK(clk), .Q(sram_rdata_7[3]), .QN(n385) );
  DFFSSRX1_HVT sram_rdata_7_reg_2_ ( .D(1'b0), .SETB(n2410), .RSTB(N265), 
        .CLK(clk), .Q(sram_rdata_7[2]), .QN(n384) );
  DFFSSRX1_HVT sram_rdata_7_reg_1_ ( .D(1'b0), .SETB(n2850), .RSTB(N264), 
        .CLK(clk), .Q(sram_rdata_7[1]), .QN(n383) );
  DFFSSRX1_HVT sram_rdata_7_reg_0_ ( .D(1'b0), .SETB(n13300), .RSTB(N263), 
        .CLK(clk), .Q(sram_rdata_7[0]), .QN(n2860) );
  AO221X1_HVT U3 ( .A1(1'b1), .A2(n9600), .A3(sram_rdata_1[27]), .A4(n575), 
        .A5(n9700), .Y(n_src_aox[283]) );
  AO221X1_HVT U4 ( .A1(1'b1), .A2(n9300), .A3(sram_rdata_1[18]), .A4(n2220), 
        .A5(n9400), .Y(n_src_aox[274]) );
  AO221X1_HVT U5 ( .A1(1'b1), .A2(n9000), .A3(sram_rdata_1[26]), .A4(n2210), 
        .A5(n9100), .Y(n_src_aox[282]) );
  AO221X1_HVT U6 ( .A1(1'b1), .A2(n8700), .A3(sram_rdata_1[23]), .A4(n2270), 
        .A5(n8800), .Y(n_src_aox[279]) );
  AO221X1_HVT U7 ( .A1(1'b1), .A2(n8400), .A3(sram_rdata_1[25]), .A4(n1720), 
        .A5(n8500), .Y(n_src_aox[281]) );
  AO221X1_HVT U8 ( .A1(1'b1), .A2(n8100), .A3(sram_rdata_0[27]), .A4(n2280), 
        .A5(n8200), .Y(n_src_aox[251]) );
  AO221X1_HVT U9 ( .A1(1'b1), .A2(n7800), .A3(sram_rdata_1[24]), .A4(n2240), 
        .A5(n7900), .Y(n_src_aox[280]) );
  AO221X1_HVT U10 ( .A1(1'b1), .A2(n7500), .A3(sram_rdata_2[26]), .A4(n1810), 
        .A5(n7600), .Y(n_src_aox[266]) );
  AO221X1_HVT U11 ( .A1(1'b1), .A2(n7200), .A3(sram_rdata_1[20]), .A4(n1750), 
        .A5(n7300), .Y(n_src_aox[276]) );
  AO221X1_HVT U12 ( .A1(1'b1), .A2(n6900), .A3(sram_rdata_1[14]), .A4(n2220), 
        .A5(n7000), .Y(n_src_aox[238]) );
  AO221X1_HVT U13 ( .A1(1'b1), .A2(n6600), .A3(sram_rdata_1[19]), .A4(n576), 
        .A5(n6700), .Y(n_src_aox[275]) );
  AO221X1_HVT U14 ( .A1(1'b1), .A2(n6300), .A3(sram_rdata_2[30]), .A4(n2260), 
        .A5(n6400), .Y(n_src_aox[270]) );
  AO221X1_HVT U15 ( .A1(1'b1), .A2(n6000), .A3(sram_rdata_2[25]), .A4(n2280), 
        .A5(n6100), .Y(n_src_aox[265]) );
  AO221X1_HVT U16 ( .A1(1'b1), .A2(n5700), .A3(sram_rdata_5[30]), .A4(n2210), 
        .A5(n5800), .Y(n_src_aox[174]) );
  AO221X1_HVT U17 ( .A1(1'b1), .A2(n5400), .A3(sram_rdata_2[24]), .A4(n574), 
        .A5(n5500), .Y(n_src_aox[264]) );
  AO221X1_HVT U18 ( .A1(1'b1), .A2(n5100), .A3(sram_rdata_1[6]), .A4(n1750), 
        .A5(n5200), .Y(n_src_aox[230]) );
  AO221X1_HVT U19 ( .A1(1'b1), .A2(n4800), .A3(sram_rdata_2[18]), .A4(n2250), 
        .A5(n4900), .Y(n_src_aox[258]) );
  AO221X1_HVT U20 ( .A1(1'b1), .A2(n4500), .A3(sram_rdata_2[7]), .A4(n2260), 
        .A5(n4600), .Y(n_src_aox[215]) );
  AO221X1_HVT U21 ( .A1(1'b1), .A2(n4200), .A3(sram_rdata_0[31]), .A4(n575), 
        .A5(n4300), .Y(n_src_aox[255]) );
  AO221X1_HVT U22 ( .A1(1'b1), .A2(n3900), .A3(sram_rdata_3[26]), .A4(n1760), 
        .A5(n4000), .Y(n_src_aox[154]) );
  AO221X1_HVT U23 ( .A1(1'b1), .A2(n35), .A3(sram_rdata_0[24]), .A4(n1760), 
        .A5(n36), .Y(n_src_aox[248]) );
  AO221X1_HVT U24 ( .A1(1'b1), .A2(n32), .A3(sram_rdata_4[26]), .A4(n2250), 
        .A5(n33), .Y(n_src_aox[186]) );
  AO221X1_HVT U25 ( .A1(1'b1), .A2(n29), .A3(sram_rdata_1[0]), .A4(n2240), 
        .A5(n30), .Y(n_src_aox[224]) );
  AO221X1_HVT U26 ( .A1(1'b1), .A2(n26), .A3(sram_rdata_5[25]), .A4(n1800), 
        .A5(n27), .Y(n_src_aox[169]) );
  AO221X1_HVT U27 ( .A1(1'b1), .A2(n23), .A3(sram_rdata_2[0]), .A4(n1790), 
        .A5(n24), .Y(n_src_aox[208]) );
  AO221X1_HVT U28 ( .A1(1'b1), .A2(n20), .A3(sram_rdata_4[1]), .A4(n575), .A5(
        n21), .Y(n_src_aox[129]) );
  AO221X1_HVT U29 ( .A1(1'b1), .A2(n17), .A3(sram_rdata_0[12]), .A4(n1820), 
        .A5(n18), .Y(n_src_aox[204]) );
  AO221X1_HVT U30 ( .A1(1'b1), .A2(n14), .A3(sram_rdata_7[30]), .A4(n2220), 
        .A5(n15), .Y(n_src_aox[94]) );
  AO221X1_HVT U31 ( .A1(1'b1), .A2(n11), .A3(sram_rdata_0[11]), .A4(n1720), 
        .A5(n12), .Y(n_src_aox[203]) );
  AO221X1_HVT U32 ( .A1(1'b1), .A2(n8), .A3(sram_rdata_4[29]), .A4(n2210), 
        .A5(n9), .Y(n_src_aox[189]) );
  AO221X1_HVT U33 ( .A1(1'b1), .A2(n5), .A3(sram_rdata_0[5]), .A4(n1820), .A5(
        n6), .Y(n_src_aox[197]) );
  AO221X1_HVT U34 ( .A1(1'b1), .A2(n2), .A3(sram_rdata_6[11]), .A4(n2230), 
        .A5(n3), .Y(n_src_aox[11]) );
  NBUFFX2_HVT U35 ( .A(n1658), .Y(n587) );
  INVX1_HVT U36 ( .A(n584), .Y(n10500) );
  INVX1_HVT U37 ( .A(n583), .Y(n10400) );
  INVX1_HVT U38 ( .A(n584), .Y(n10300) );
  INVX1_HVT U39 ( .A(n583), .Y(n10600) );
  AO22X1_HVT U41 ( .A1(n922), .A2(n12600), .A3(n591), .A4(n1297), .Y(n2) );
  OAI22X1_HVT U42 ( .A1(n11800), .A2(n393), .A3(n2730), .A4(n2970), .Y(n3) );
  AO22X1_HVT U44 ( .A1(n1269), .A2(n1663), .A3(n12600), .A4(n12701), .Y(n5) );
  OAI22X1_HVT U45 ( .A1(n2790), .A2(n355), .A3(n10100), .A4(n546), .Y(n6) );
  AO22X1_HVT U47 ( .A1(n1637), .A2(n15100), .A3(n12700), .A4(n1235), .Y(n8) );
  OAI22X1_HVT U48 ( .A1(n12000), .A2(n538), .A3(n2730), .A4(n442), .Y(n9) );
  AO22X1_HVT U50 ( .A1(n1296), .A2(n14900), .A3(n1648), .A4(n1297), .Y(n11) );
  OAI22X1_HVT U51 ( .A1(n10600), .A2(n361), .A3(n2710), .A4(n552), .Y(n12) );
  AO22X1_HVT U53 ( .A1(n1236), .A2(n10900), .A3(n15000), .A4(n1643), .Y(n14)
         );
  OAI22X1_HVT U54 ( .A1(n2780), .A2(n3160), .A3(n14800), .A4(n508), .Y(n15) );
  AO22X1_HVT U56 ( .A1(n1298), .A2(n14900), .A3(n12900), .A4(n1299), .Y(n17)
         );
  OAI22X1_HVT U57 ( .A1(n11900), .A2(n362), .A3(n2710), .A4(n553), .Y(n18) );
  AO22X1_HVT U59 ( .A1(n1391), .A2(n12900), .A3(n12700), .A4(n10101), .Y(n20)
         );
  OAI22X1_HVT U60 ( .A1(n11900), .A2(n5101), .A3(n2730), .A4(n414), .Y(n21) );
  AO22X1_HVT U62 ( .A1(n1315), .A2(n11000), .A3(n591), .A4(n1316), .Y(n23) );
  OAI22X1_HVT U63 ( .A1(n10400), .A2(n445), .A3(n2690), .A4(n350), .Y(n24) );
  AO22X1_HVT U65 ( .A1(n15701), .A2(n12600), .A3(n12800), .A4(n1164), .Y(n26)
         );
  OAI22X1_HVT U66 ( .A1(n2800), .A2(n438), .A3(n14700), .A4(n343), .Y(n27) );
  AO22X1_HVT U68 ( .A1(n1389), .A2(n10900), .A3(n15000), .A4(n13901), .Y(n29)
         );
  OAI22X1_HVT U69 ( .A1(n10400), .A2(n541), .A3(n14500), .A4(n445), .Y(n30) );
  AO22X1_HVT U71 ( .A1(n1628), .A2(n579), .A3(n588), .A4(n1226), .Y(n32) );
  OAI22X1_HVT U72 ( .A1(n2760), .A2(n535), .A3(n2730), .A4(n439), .Y(n33) );
  AO22X1_HVT U74 ( .A1(n15001), .A2(n1663), .A3(n12600), .A4(n1501), .Y(n35)
         );
  OAI22X1_HVT U75 ( .A1(n13700), .A2(n374), .A3(n14500), .A4(n565), .Y(n36) );
  INVX0_HVT U76 ( .A(mode[0]), .Y(n37) );
  AND2X1_HVT U77 ( .A1(mode[1]), .A2(n37), .Y(n1664) );
  AO22X1_HVT U79 ( .A1(n1507), .A2(n15200), .A3(n15000), .A4(n1107), .Y(n3900)
         );
  OAI22X1_HVT U80 ( .A1(n2760), .A2(n344), .A3(n2720), .A4(n535), .Y(n4000) );
  AO22X1_HVT U82 ( .A1(n1529), .A2(n1663), .A3(n12600), .A4(n15301), .Y(n4200)
         );
  OAI22X1_HVT U83 ( .A1(n12100), .A2(n381), .A3(n2700), .A4(n572), .Y(n4300)
         );
  AO22X1_HVT U85 ( .A1(n1347), .A2(n12700), .A3(n11000), .A4(n1348), .Y(n4500)
         );
  OAI22X1_HVT U86 ( .A1(n2760), .A2(n452), .A3(n14500), .A4(n357), .Y(n4600)
         );
  AO22X1_HVT U88 ( .A1(n1541), .A2(n10800), .A3(n579), .A4(n1542), .Y(n4800)
         );
  OAI22X1_HVT U89 ( .A1(n10300), .A2(n463), .A3(n14700), .A4(n368), .Y(n4900)
         );
  AO22X1_HVT U91 ( .A1(n1416), .A2(n10700), .A3(n581), .A4(n1417), .Y(n5100)
         );
  OAI22X1_HVT U92 ( .A1(n11800), .A2(n547), .A3(n2730), .A4(n451), .Y(n5200)
         );
  AO22X1_HVT U94 ( .A1(n1568), .A2(n12700), .A3(n581), .A4(n1569), .Y(n5400)
         );
  OAI22X1_HVT U95 ( .A1(n13700), .A2(n469), .A3(n10000), .A4(n374), .Y(n5500)
         );
  AO22X1_HVT U97 ( .A1(n1589), .A2(n12600), .A3(n591), .A4(n1181), .Y(n5700)
         );
  OAI22X1_HVT U98 ( .A1(n2780), .A2(n443), .A3(n2730), .A4(n348), .Y(n5800) );
  AO22X1_HVT U100 ( .A1(n15701), .A2(n10700), .A3(n5801), .A4(n1571), .Y(n6000) );
  OAI22X1_HVT U101 ( .A1(n2800), .A2(n4701), .A3(n10100), .A4(n375), .Y(n6100)
         );
  AO22X1_HVT U103 ( .A1(n1589), .A2(n10800), .A3(n12900), .A4(n15901), .Y(
        n6300) );
  OAI22X1_HVT U104 ( .A1(n13800), .A2(n475), .A3(n2750), .A4(n380), .Y(n6400)
         );
  AO22X1_HVT U106 ( .A1(n1608), .A2(n10800), .A3(n12600), .A4(n1609), .Y(n6600) );
  OAI22X1_HVT U107 ( .A1(n2780), .A2(n5601), .A3(n14600), .A4(n464), .Y(n6700)
         );
  AO22X1_HVT U109 ( .A1(n1453), .A2(n12700), .A3(n5801), .A4(n1454), .Y(n6900)
         );
  OAI22X1_HVT U110 ( .A1(n2770), .A2(n555), .A3(n2740), .A4(n459), .Y(n7000)
         );
  AO22X1_HVT U112 ( .A1(n16101), .A2(n10800), .A3(n581), .A4(n1611), .Y(n7200)
         );
  OAI22X1_HVT U113 ( .A1(n2800), .A2(n561), .A3(n2690), .A4(n465), .Y(n7300)
         );
  AO22X1_HVT U115 ( .A1(n1572), .A2(n12800), .A3(n581), .A4(n1573), .Y(n7500)
         );
  OAI22X1_HVT U116 ( .A1(n2760), .A2(n471), .A3(n1661), .A4(n376), .Y(n7600)
         );
  AO22X1_HVT U118 ( .A1(n1624), .A2(n10700), .A3(n12900), .A4(n1625), .Y(n7800) );
  OAI22X1_HVT U119 ( .A1(n2790), .A2(n565), .A3(n2710), .A4(n469), .Y(n7900)
         );
  AO22X1_HVT U121 ( .A1(n1512), .A2(n12800), .A3(n578), .A4(n1513), .Y(n8100)
         );
  OAI22X1_HVT U122 ( .A1(n11800), .A2(n377), .A3(n10000), .A4(n568), .Y(n8200)
         );
  AO22X1_HVT U124 ( .A1(n1626), .A2(n12800), .A3(n581), .A4(n1627), .Y(n8400)
         );
  OAI22X1_HVT U125 ( .A1(n2810), .A2(n566), .A3(n2740), .A4(n4701), .Y(n8500)
         );
  AO22X1_HVT U127 ( .A1(n1622), .A2(n12800), .A3(n582), .A4(n1623), .Y(n8700)
         );
  OAI22X1_HVT U128 ( .A1(n2760), .A2(n564), .A3(n14600), .A4(n468), .Y(n8800)
         );
  AO22X1_HVT U130 ( .A1(n1628), .A2(n12700), .A3(n15200), .A4(n1629), .Y(n9000) );
  OAI22X1_HVT U131 ( .A1(n1662), .A2(n567), .A3(n2740), .A4(n471), .Y(n9100)
         );
  AO22X1_HVT U133 ( .A1(n1606), .A2(n10700), .A3(n15200), .A4(n1607), .Y(n9300) );
  OAI22X1_HVT U134 ( .A1(n12100), .A2(n559), .A3(n2720), .A4(n463), .Y(n9400)
         );
  AO22X1_HVT U136 ( .A1(n16301), .A2(n1663), .A3(n12600), .A4(n1631), .Y(n9600) );
  OAI22X1_HVT U137 ( .A1(n10600), .A2(n568), .A3(n2710), .A4(n472), .Y(n9700)
         );
  NBUFFX2_HVT U138 ( .A(n16501), .Y(n1720) );
  INVX1_HVT U139 ( .A(n1659), .Y(n11100) );
  INVX2_HVT U140 ( .A(n2610), .Y(n9800) );
  INVX2_HVT U141 ( .A(n2610), .Y(n9900) );
  INVX1_HVT U142 ( .A(n2350), .Y(n11700) );
  INVX1_HVT U143 ( .A(n14400), .Y(n11600) );
  INVX1_HVT U144 ( .A(n583), .Y(n11800) );
  INVX1_HVT U145 ( .A(n584), .Y(n11900) );
  INVX2_HVT U146 ( .A(n585), .Y(n10000) );
  INVX1_HVT U147 ( .A(n584), .Y(n12000) );
  INVX2_HVT U148 ( .A(n585), .Y(n10100) );
  INVX1_HVT U149 ( .A(n584), .Y(n12100) );
  INVX0_HVT U150 ( .A(n584), .Y(n13700) );
  INVX0_HVT U151 ( .A(n584), .Y(n13800) );
  INVX2_HVT U152 ( .A(n14400), .Y(n10200) );
  INVX1_HVT U153 ( .A(n586), .Y(n2750) );
  INVX2_HVT U154 ( .A(n1661), .Y(n585) );
  INVX1_HVT U155 ( .A(n1661), .Y(n586) );
  INVX2_HVT U156 ( .A(n16200), .Y(n10700) );
  INVX2_HVT U157 ( .A(n16200), .Y(n10800) );
  INVX2_HVT U158 ( .A(n16300), .Y(n10900) );
  INVX2_HVT U159 ( .A(n16300), .Y(n11000) );
  INVX1_HVT U160 ( .A(srstn), .Y(n2830) );
  INVX1_HVT U161 ( .A(srstn), .Y(n2850) );
  INVX1_HVT U162 ( .A(srstn), .Y(n2840) );
  INVX1_HVT U163 ( .A(n16601), .Y(n11200) );
  INVX1_HVT U164 ( .A(n2610), .Y(n13100) );
  INVX1_HVT U165 ( .A(n2610), .Y(n13000) );
  INVX2_HVT U166 ( .A(n2610), .Y(n11300) );
  INVX2_HVT U167 ( .A(n2570), .Y(n11400) );
  INVX2_HVT U168 ( .A(n585), .Y(n11500) );
  INVX2_HVT U169 ( .A(n586), .Y(n2740) );
  INVX1_HVT U170 ( .A(n2570), .Y(n2600) );
  INVX2_HVT U171 ( .A(n585), .Y(n2710) );
  INVX1_HVT U172 ( .A(n577), .Y(n2570) );
  INVX1_HVT U173 ( .A(N346), .Y(n2610) );
  INVX1_HVT U174 ( .A(n15300), .Y(n15800) );
  INVX1_HVT U175 ( .A(n15300), .Y(n16000) );
  INVX1_HVT U176 ( .A(n15300), .Y(n16100) );
  INVX1_HVT U177 ( .A(n15300), .Y(n15900) );
  INVX1_HVT U178 ( .A(n2520), .Y(n13400) );
  INVX1_HVT U179 ( .A(n2400), .Y(n13200) );
  INVX1_HVT U180 ( .A(n2470), .Y(n13300) );
  INVX1_HVT U181 ( .A(n1870), .Y(n1880) );
  INVX1_HVT U182 ( .A(n1870), .Y(n1900) );
  INVX1_HVT U183 ( .A(n1870), .Y(n1890) );
  INVX1_HVT U184 ( .A(n1662), .Y(n584) );
  INVX1_HVT U185 ( .A(n1662), .Y(n583) );
  INVX1_HVT U186 ( .A(n1870), .Y(n1910) );
  INVX1_HVT U187 ( .A(n2820), .Y(n593) );
  INVX2_HVT U188 ( .A(n2520), .Y(n12200) );
  INVX2_HVT U189 ( .A(n2400), .Y(n12300) );
  INVX2_HVT U190 ( .A(n2470), .Y(n12400) );
  INVX1_HVT U191 ( .A(n15300), .Y(n15500) );
  INVX1_HVT U192 ( .A(n15300), .Y(n15600) );
  INVX1_HVT U193 ( .A(n15300), .Y(n15700) );
  INVX1_HVT U194 ( .A(n13900), .Y(n1870) );
  INVX1_HVT U195 ( .A(n15300), .Y(n15400) );
  NAND3X0_HVT U196 ( .A1(n1655), .A2(n1654), .A3(n2070), .Y(n1661) );
  INVX1_HVT U197 ( .A(n11100), .Y(n2070) );
  INVX1_HVT U198 ( .A(n11100), .Y(n13900) );
  NAND3X0_HVT U199 ( .A1(n1655), .A2(n1654), .A3(n2160), .Y(n1662) );
  INVX1_HVT U200 ( .A(n2200), .Y(n2250) );
  NBUFFX2_HVT U201 ( .A(n1664), .Y(n2820) );
  INVX1_HVT U202 ( .A(n13500), .Y(n15300) );
  INVX1_HVT U203 ( .A(n11200), .Y(n1920) );
  INVX1_HVT U204 ( .A(n1780), .Y(n1740) );
  INVX1_HVT U205 ( .A(n11200), .Y(n16600) );
  INVX1_HVT U206 ( .A(n1780), .Y(n1770) );
  INVX1_HVT U207 ( .A(n11200), .Y(n1700) );
  INVX1_HVT U208 ( .A(n1950), .Y(n2000) );
  INVX1_HVT U209 ( .A(n11200), .Y(n1940) );
  INVX1_HVT U210 ( .A(n11200), .Y(n1710) );
  INVX1_HVT U211 ( .A(n1780), .Y(n1760) );
  INVX1_HVT U212 ( .A(n11200), .Y(n1670) );
  INVX1_HVT U213 ( .A(n11200), .Y(n1930) );
  INVX1_HVT U214 ( .A(n2200), .Y(n2230) );
  INVX1_HVT U215 ( .A(n1950), .Y(n1980) );
  INVX1_HVT U216 ( .A(n2200), .Y(n2220) );
  INVX1_HVT U217 ( .A(n1950), .Y(n2010) );
  INVX1_HVT U218 ( .A(n1780), .Y(n1750) );
  INVX1_HVT U219 ( .A(n1950), .Y(n2020) );
  INVX1_HVT U220 ( .A(n1950), .Y(n1990) );
  INVX1_HVT U221 ( .A(n1780), .Y(n1800) );
  INVX1_HVT U222 ( .A(n11200), .Y(n16500) );
  INVX1_HVT U223 ( .A(n2200), .Y(n2210) );
  INVX1_HVT U224 ( .A(n1780), .Y(n1820) );
  INVX1_HVT U225 ( .A(n1780), .Y(n1790) );
  INVX1_HVT U226 ( .A(n11200), .Y(n16400) );
  INVX1_HVT U227 ( .A(n1950), .Y(n1970) );
  INVX1_HVT U228 ( .A(n1950), .Y(n1960) );
  INVX1_HVT U229 ( .A(n11200), .Y(n1680) );
  INVX1_HVT U230 ( .A(n1780), .Y(n1810) );
  INVX1_HVT U231 ( .A(n11200), .Y(n1690) );
  INVX1_HVT U232 ( .A(n2200), .Y(n2240) );
  INVX1_HVT U233 ( .A(n2830), .Y(n2400) );
  INVX1_HVT U234 ( .A(n2840), .Y(n2470) );
  INVX1_HVT U235 ( .A(n2850), .Y(n2520) );
  INVX1_HVT U236 ( .A(n2150), .Y(n2160) );
  INVX1_HVT U237 ( .A(n575), .Y(n2200) );
  INVX1_HVT U238 ( .A(n11100), .Y(n12500) );
  INVX1_HVT U239 ( .A(n2150), .Y(n13500) );
  INVX1_HVT U240 ( .A(n15300), .Y(n2140) );
  INVX2_HVT U241 ( .A(n16300), .Y(n12600) );
  INVX1_HVT U242 ( .A(n16601), .Y(n1950) );
  INVX1_HVT U243 ( .A(n15300), .Y(n2120) );
  INVX1_HVT U244 ( .A(n576), .Y(n1780) );
  INVX1_HVT U245 ( .A(n15300), .Y(n2110) );
  INVX1_HVT U246 ( .A(n2150), .Y(n2130) );
  INVX2_HVT U247 ( .A(n16200), .Y(n12700) );
  INVX2_HVT U248 ( .A(n16200), .Y(n12800) );
  INVX2_HVT U249 ( .A(n16300), .Y(n12900) );
  DELLN1X2_HVT U250 ( .A(n1663), .Y(n589) );
  DELLN1X2_HVT U251 ( .A(n16501), .Y(n574) );
  DELLN1X2_HVT U252 ( .A(n1648), .Y(n581) );
  INVX1_HVT U253 ( .A(n587), .Y(n2150) );
  DELLN1X2_HVT U254 ( .A(n16501), .Y(n576) );
  INVX2_HVT U255 ( .A(n2400), .Y(n2420) );
  INVX1_HVT U256 ( .A(n2400), .Y(n2430) );
  INVX2_HVT U257 ( .A(srstn), .Y(n2450) );
  INVX1_HVT U258 ( .A(srstn), .Y(n2460) );
  INVX2_HVT U259 ( .A(n2470), .Y(n2490) );
  INVX1_HVT U260 ( .A(n2470), .Y(n2500) );
  INVX2_HVT U261 ( .A(n2520), .Y(n2540) );
  INVX1_HVT U262 ( .A(n2520), .Y(n2550) );
  INVX0_HVT U263 ( .A(n2150), .Y(n13600) );
  DELLN1X2_HVT U264 ( .A(n1648), .Y(n578) );
  DELLN1X2_HVT U265 ( .A(n1648), .Y(n579) );
  DELLN1X2_HVT U266 ( .A(n1648), .Y(n582) );
  DELLN1X2_HVT U267 ( .A(n1648), .Y(n5801) );
  DELLN1X2_HVT U268 ( .A(n1648), .Y(n15200) );
  DELLN1X2_HVT U269 ( .A(n1648), .Y(n15100) );
  DELLN1X2_HVT U270 ( .A(n1663), .Y(n591) );
  NBUFFX2_HVT U271 ( .A(n1663), .Y(n588) );
  DELLN1X2_HVT U272 ( .A(n1663), .Y(n592) );
  DELLN1X2_HVT U273 ( .A(n1663), .Y(n5901) );
  DELLN1X2_HVT U274 ( .A(n1663), .Y(n15000) );
  DELLN1X2_HVT U275 ( .A(n1663), .Y(n14900) );
  INVX2_HVT U276 ( .A(n2570), .Y(n2590) );
  INVX2_HVT U277 ( .A(n2570), .Y(n2580) );
  INVX2_HVT U278 ( .A(n2610), .Y(n2630) );
  INVX2_HVT U279 ( .A(n2610), .Y(n2620) );
  NBUFFX2_HVT U280 ( .A(N346), .Y(n577) );
  INVX2_HVT U281 ( .A(n593), .Y(n14000) );
  INVX2_HVT U282 ( .A(n593), .Y(n14100) );
  INVX2_HVT U283 ( .A(n593), .Y(n2650) );
  INVX2_HVT U284 ( .A(n593), .Y(n2640) );
  INVX2_HVT U285 ( .A(n2340), .Y(n14200) );
  INVX2_HVT U286 ( .A(n14400), .Y(n14300) );
  INVX2_HVT U287 ( .A(n14400), .Y(n2680) );
  INVX2_HVT U288 ( .A(n14400), .Y(n2670) );
  INVX2_HVT U289 ( .A(n14400), .Y(n2660) );
  INVX0_HVT U290 ( .A(n2820), .Y(n14400) );
  DELLN1X2_HVT U291 ( .A(n16501), .Y(n575) );
  DELLN1X2_HVT U292 ( .A(n16501), .Y(n1730) );
  INVX2_HVT U293 ( .A(n585), .Y(n14500) );
  INVX2_HVT U294 ( .A(n585), .Y(n14600) );
  INVX2_HVT U295 ( .A(n585), .Y(n2700) );
  INVX2_HVT U296 ( .A(n585), .Y(n2690) );
  INVX2_HVT U297 ( .A(n586), .Y(n14700) );
  INVX2_HVT U298 ( .A(n586), .Y(n14800) );
  INVX2_HVT U299 ( .A(n586), .Y(n2730) );
  INVX2_HVT U300 ( .A(n586), .Y(n2720) );
  INVX1_HVT U301 ( .A(n583), .Y(n2770) );
  INVX1_HVT U302 ( .A(n583), .Y(n2780) );
  INVX1_HVT U303 ( .A(n583), .Y(n2760) );
  INVX1_HVT U304 ( .A(n584), .Y(n2800) );
  INVX1_HVT U305 ( .A(n584), .Y(n2810) );
  INVX1_HVT U306 ( .A(n584), .Y(n2790) );
  INVX0_HVT U307 ( .A(n588), .Y(n16200) );
  INVX0_HVT U308 ( .A(n15100), .Y(n16300) );
  INVX0_HVT U309 ( .A(n11100), .Y(n1830) );
  INVX0_HVT U310 ( .A(n11100), .Y(n1840) );
  INVX0_HVT U311 ( .A(n11100), .Y(n1850) );
  INVX0_HVT U312 ( .A(n11100), .Y(n1860) );
  INVX0_HVT U313 ( .A(n11100), .Y(n2030) );
  INVX0_HVT U314 ( .A(n11100), .Y(n2040) );
  INVX0_HVT U315 ( .A(n11100), .Y(n2050) );
  INVX0_HVT U316 ( .A(n11100), .Y(n2060) );
  INVX0_HVT U317 ( .A(n1870), .Y(n2080) );
  INVX0_HVT U318 ( .A(n1870), .Y(n2090) );
  INVX0_HVT U319 ( .A(n1870), .Y(n2100) );
  INVX0_HVT U320 ( .A(n2150), .Y(n2170) );
  INVX0_HVT U321 ( .A(n2150), .Y(n2180) );
  INVX0_HVT U322 ( .A(n2150), .Y(n2190) );
  INVX0_HVT U323 ( .A(n1780), .Y(n2260) );
  INVX0_HVT U324 ( .A(n1780), .Y(n2270) );
  INVX0_HVT U325 ( .A(n1780), .Y(n2280) );
  INVX2_HVT U326 ( .A(n1664), .Y(n2290) );
  INVX2_HVT U327 ( .A(n1664), .Y(n2300) );
  INVX2_HVT U328 ( .A(n1664), .Y(n2310) );
  INVX2_HVT U329 ( .A(n1664), .Y(n2320) );
  INVX2_HVT U330 ( .A(n2820), .Y(n2330) );
  INVX2_HVT U331 ( .A(n2820), .Y(n2340) );
  INVX2_HVT U332 ( .A(n2820), .Y(n2350) );
  INVX2_HVT U333 ( .A(n2820), .Y(n2360) );
  INVX2_HVT U334 ( .A(n2820), .Y(n2370) );
  INVX2_HVT U335 ( .A(n2820), .Y(n2380) );
  INVX2_HVT U336 ( .A(n2820), .Y(n2390) );
  INVX2_HVT U337 ( .A(n2400), .Y(n2410) );
  INVX2_HVT U338 ( .A(n2400), .Y(n2440) );
  INVX2_HVT U339 ( .A(n2470), .Y(n2480) );
  INVX2_HVT U340 ( .A(n2470), .Y(n2510) );
  INVX2_HVT U341 ( .A(n2520), .Y(n2530) );
  INVX2_HVT U342 ( .A(n2520), .Y(n2560) );
  INVX1_HVT U343 ( .A(box_sel[1]), .Y(n1656) );
  INVX1_HVT U344 ( .A(box_sel[2]), .Y(n1655) );
  INVX1_HVT U345 ( .A(box_sel[3]), .Y(n1654) );
  INVX1_HVT U346 ( .A(box_sel[0]), .Y(n1657) );
  NAND2X0_HVT U347 ( .A1(n2250), .A2(n1656), .Y(n594) );
  AND3X1_HVT U348 ( .A1(n1657), .A2(n1654), .A3(n1655), .Y(n16501) );
  NAND2X0_HVT U349 ( .A1(srstn), .A2(n594), .Y(N346) );
  AO222X1_HVT U350 ( .A1(n2040), .A2(sram_rdata_5[0]), .A3(n2010), .A4(
        sram_rdata_3[0]), .A5(n15400), .A6(sram_rdata_4[0]), .Y(n1244) );
  AND2X1_HVT U351 ( .A1(n1654), .A2(box_sel[2]), .Y(n1648) );
  AO222X1_HVT U352 ( .A1(n1850), .A2(sram_rdata_2[0]), .A3(n15700), .A4(
        sram_rdata_1[0]), .A5(sram_rdata_0[0]), .A6(n1940), .Y(n878) );
  AOI22X1_HVT U353 ( .A1(n1244), .A2(n10800), .A3(n11000), .A4(n878), .Y(n597)
         );
  OA22X1_HVT U354 ( .A1(n2800), .A2(n2860), .A3(n2720), .A4(n573), .Y(n596) );
  NAND2X0_HVT U355 ( .A1(n1770), .A2(sram_rdata_6[0]), .Y(n595) );
  NAND3X0_HVT U356 ( .A1(n597), .A2(n596), .A3(n595), .Y(n_src_aox[0]) );
  AO222X1_HVT U357 ( .A1(n1659), .A2(sram_rdata_5[1]), .A3(n13500), .A4(
        sram_rdata_4[1]), .A5(sram_rdata_3[1]), .A6(n16400), .Y(n12501) );
  AO222X1_HVT U358 ( .A1(n2030), .A2(sram_rdata_2[1]), .A3(n15900), .A4(
        sram_rdata_1[1]), .A5(sram_rdata_0[1]), .A6(n16400), .Y(n882) );
  AOI22X1_HVT U359 ( .A1(n12501), .A2(n14900), .A3(n579), .A4(n882), .Y(n6001)
         );
  OA22X1_HVT U360 ( .A1(n11900), .A2(n383), .A3(n14500), .A4(n2870), .Y(n599)
         );
  NAND2X0_HVT U361 ( .A1(n2240), .A2(sram_rdata_6[1]), .Y(n598) );
  NAND3X0_HVT U362 ( .A1(n6001), .A2(n599), .A3(n598), .Y(n_src_aox[1]) );
  AO222X1_HVT U363 ( .A1(n2040), .A2(sram_rdata_5[2]), .A3(n2120), .A4(
        sram_rdata_4[2]), .A5(sram_rdata_3[2]), .A6(n1670), .Y(n1255) );
  AO222X1_HVT U364 ( .A1(n2050), .A2(sram_rdata_2[2]), .A3(n15900), .A4(
        sram_rdata_1[2]), .A5(sram_rdata_0[2]), .A6(n1690), .Y(n886) );
  AOI22X1_HVT U365 ( .A1(n1255), .A2(n10700), .A3(n579), .A4(n886), .Y(n603)
         );
  OA22X1_HVT U366 ( .A1(n11800), .A2(n384), .A3(n10000), .A4(n2880), .Y(n602)
         );
  NAND2X0_HVT U367 ( .A1(n1800), .A2(sram_rdata_6[2]), .Y(n601) );
  NAND3X0_HVT U368 ( .A1(n603), .A2(n602), .A3(n601), .Y(n_src_aox[2]) );
  AO222X1_HVT U369 ( .A1(n1860), .A2(sram_rdata_5[3]), .A3(n15700), .A4(
        sram_rdata_4[3]), .A5(sram_rdata_3[3]), .A6(n16400), .Y(n12601) );
  AO222X1_HVT U370 ( .A1(n1659), .A2(sram_rdata_2[3]), .A3(n16000), .A4(
        sram_rdata_1[3]), .A5(sram_rdata_0[3]), .A6(n1700), .Y(n8901) );
  AOI22X1_HVT U371 ( .A1(n12601), .A2(n588), .A3(n582), .A4(n8901), .Y(n606)
         );
  OA22X1_HVT U372 ( .A1(n2770), .A2(n385), .A3(n1661), .A4(n2890), .Y(n605) );
  NAND2X0_HVT U373 ( .A1(n574), .A2(sram_rdata_6[3]), .Y(n604) );
  NAND3X0_HVT U374 ( .A1(n606), .A2(n605), .A3(n604), .Y(n_src_aox[3]) );
  AO222X1_HVT U375 ( .A1(n2080), .A2(sram_rdata_5[4]), .A3(n2130), .A4(
        sram_rdata_4[4]), .A5(sram_rdata_3[4]), .A6(n1940), .Y(n1265) );
  AO222X1_HVT U376 ( .A1(n1910), .A2(sram_rdata_2[4]), .A3(n15500), .A4(
        sram_rdata_1[4]), .A5(sram_rdata_0[4]), .A6(n2010), .Y(n894) );
  AOI22X1_HVT U377 ( .A1(n1265), .A2(n10700), .A3(n15100), .A4(n894), .Y(n609)
         );
  OA22X1_HVT U378 ( .A1(n13800), .A2(n386), .A3(n14700), .A4(n2900), .Y(n608)
         );
  NAND2X0_HVT U379 ( .A1(n1790), .A2(sram_rdata_6[4]), .Y(n607) );
  NAND3X0_HVT U380 ( .A1(n609), .A2(n608), .A3(n607), .Y(n_src_aox[4]) );
  AO222X1_HVT U381 ( .A1(n1860), .A2(sram_rdata_5[5]), .A3(n2160), .A4(
        sram_rdata_4[5]), .A5(sram_rdata_3[5]), .A6(n1990), .Y(n12701) );
  AO222X1_HVT U382 ( .A1(n1850), .A2(sram_rdata_2[5]), .A3(n16100), .A4(
        sram_rdata_1[5]), .A5(sram_rdata_0[5]), .A6(n1920), .Y(n898) );
  AOI22X1_HVT U383 ( .A1(n12701), .A2(n10700), .A3(n582), .A4(n898), .Y(n612)
         );
  OA22X1_HVT U384 ( .A1(n2790), .A2(n387), .A3(n2690), .A4(n2910), .Y(n611) );
  NAND2X0_HVT U385 ( .A1(n574), .A2(sram_rdata_6[5]), .Y(n6101) );
  NAND3X0_HVT U386 ( .A1(n612), .A2(n611), .A3(n6101), .Y(n_src_aox[5]) );
  AO222X1_HVT U387 ( .A1(n2030), .A2(sram_rdata_5[6]), .A3(n15500), .A4(
        sram_rdata_4[6]), .A5(sram_rdata_3[6]), .A6(n2000), .Y(n1272) );
  AO222X1_HVT U388 ( .A1(n1659), .A2(sram_rdata_2[6]), .A3(n2120), .A4(
        sram_rdata_1[6]), .A5(sram_rdata_0[6]), .A6(n1980), .Y(n902) );
  AOI22X1_HVT U389 ( .A1(n1272), .A2(n12700), .A3(n15200), .A4(n902), .Y(n615)
         );
  OA22X1_HVT U390 ( .A1(n13800), .A2(n388), .A3(n2710), .A4(n2920), .Y(n614)
         );
  NAND2X0_HVT U391 ( .A1(n2250), .A2(sram_rdata_6[6]), .Y(n613) );
  NAND3X0_HVT U392 ( .A1(n615), .A2(n614), .A3(n613), .Y(n_src_aox[6]) );
  AO222X1_HVT U393 ( .A1(n1840), .A2(sram_rdata_5[7]), .A3(n2140), .A4(
        sram_rdata_4[7]), .A5(sram_rdata_3[7]), .A6(n1980), .Y(n1277) );
  AO222X1_HVT U394 ( .A1(n1900), .A2(sram_rdata_2[7]), .A3(n15900), .A4(
        sram_rdata_1[7]), .A5(sram_rdata_0[7]), .A6(n1710), .Y(n906) );
  AOI22X1_HVT U395 ( .A1(n1277), .A2(n12800), .A3(n15200), .A4(n906), .Y(n618)
         );
  OA22X1_HVT U396 ( .A1(n13800), .A2(n389), .A3(n2750), .A4(n2930), .Y(n617)
         );
  NAND2X0_HVT U397 ( .A1(n1750), .A2(sram_rdata_6[7]), .Y(n616) );
  NAND3X0_HVT U398 ( .A1(n618), .A2(n617), .A3(n616), .Y(n_src_aox[7]) );
  AO222X1_HVT U399 ( .A1(n1850), .A2(sram_rdata_5[8]), .A3(n2120), .A4(
        sram_rdata_4[8]), .A5(sram_rdata_3[8]), .A6(n1690), .Y(n1282) );
  AO222X1_HVT U400 ( .A1(n1840), .A2(sram_rdata_2[8]), .A3(n2120), .A4(
        sram_rdata_1[8]), .A5(sram_rdata_0[8]), .A6(n1670), .Y(n9101) );
  AOI22X1_HVT U401 ( .A1(n1282), .A2(n591), .A3(n11000), .A4(n9101), .Y(n621)
         );
  OA22X1_HVT U402 ( .A1(n11900), .A2(n3901), .A3(n14800), .A4(n2940), .Y(n6201) );
  NAND2X0_HVT U403 ( .A1(n2240), .A2(sram_rdata_6[8]), .Y(n619) );
  NAND3X0_HVT U404 ( .A1(n621), .A2(n6201), .A3(n619), .Y(n_src_aox[8]) );
  AO222X1_HVT U405 ( .A1(n2060), .A2(sram_rdata_5[9]), .A3(n2130), .A4(
        sram_rdata_4[9]), .A5(sram_rdata_3[9]), .A6(n1960), .Y(n1287) );
  AO222X1_HVT U406 ( .A1(n1900), .A2(sram_rdata_2[9]), .A3(n15900), .A4(
        sram_rdata_1[9]), .A5(sram_rdata_0[9]), .A6(n1940), .Y(n914) );
  AOI22X1_HVT U407 ( .A1(n1287), .A2(n5901), .A3(n582), .A4(n914), .Y(n624) );
  OA22X1_HVT U408 ( .A1(n13700), .A2(n391), .A3(n1661), .A4(n2950), .Y(n623)
         );
  NAND2X0_HVT U409 ( .A1(n1800), .A2(sram_rdata_6[9]), .Y(n622) );
  NAND3X0_HVT U410 ( .A1(n624), .A2(n623), .A3(n622), .Y(n_src_aox[9]) );
  AO222X1_HVT U411 ( .A1(n2090), .A2(sram_rdata_5[10]), .A3(n13600), .A4(
        sram_rdata_4[10]), .A5(sram_rdata_3[10]), .A6(n1710), .Y(n1292) );
  AO222X1_HVT U412 ( .A1(n13900), .A2(sram_rdata_2[10]), .A3(n15500), .A4(
        sram_rdata_1[10]), .A5(sram_rdata_0[10]), .A6(n2020), .Y(n918) );
  AOI22X1_HVT U413 ( .A1(n1292), .A2(n12800), .A3(n12900), .A4(n918), .Y(n627)
         );
  OA22X1_HVT U414 ( .A1(n2780), .A2(n392), .A3(n11500), .A4(n2960), .Y(n626)
         );
  NAND2X0_HVT U415 ( .A1(n1770), .A2(sram_rdata_6[10]), .Y(n625) );
  NAND3X0_HVT U416 ( .A1(n627), .A2(n626), .A3(n625), .Y(n_src_aox[10]) );
  AO222X1_HVT U417 ( .A1(n12500), .A2(sram_rdata_5[11]), .A3(n2180), .A4(
        sram_rdata_4[11]), .A5(sram_rdata_3[11]), .A6(n1970), .Y(n1297) );
  AO222X1_HVT U418 ( .A1(n1659), .A2(sram_rdata_2[11]), .A3(n15400), .A4(
        sram_rdata_1[11]), .A5(sram_rdata_0[11]), .A6(n1930), .Y(n922) );
  AO222X1_HVT U419 ( .A1(n2060), .A2(sram_rdata_5[12]), .A3(n13500), .A4(
        sram_rdata_4[12]), .A5(sram_rdata_3[12]), .A6(n1940), .Y(n1299) );
  AO222X1_HVT U420 ( .A1(n1850), .A2(sram_rdata_2[12]), .A3(n16000), .A4(
        sram_rdata_1[12]), .A5(sram_rdata_0[12]), .A6(n1690), .Y(n926) );
  AOI22X1_HVT U421 ( .A1(n1299), .A2(n10800), .A3(n10900), .A4(n926), .Y(n6301) );
  OA22X1_HVT U422 ( .A1(n12000), .A2(n394), .A3(n2750), .A4(n2980), .Y(n629)
         );
  NAND2X0_HVT U423 ( .A1(n574), .A2(sram_rdata_6[12]), .Y(n628) );
  NAND3X0_HVT U424 ( .A1(n6301), .A2(n629), .A3(n628), .Y(n_src_aox[12]) );
  AO222X1_HVT U425 ( .A1(n1880), .A2(sram_rdata_5[13]), .A3(n15400), .A4(
        sram_rdata_4[13]), .A5(sram_rdata_3[13]), .A6(n1710), .Y(n1301) );
  AO222X1_HVT U426 ( .A1(n1860), .A2(sram_rdata_2[13]), .A3(n15900), .A4(
        sram_rdata_1[13]), .A5(sram_rdata_0[13]), .A6(n16500), .Y(n9301) );
  AOI22X1_HVT U427 ( .A1(n1301), .A2(n14900), .A3(n15100), .A4(n9301), .Y(n633) );
  OA22X1_HVT U428 ( .A1(n10400), .A2(n395), .A3(n11500), .A4(n2990), .Y(n632)
         );
  NAND2X0_HVT U429 ( .A1(n2280), .A2(sram_rdata_6[13]), .Y(n631) );
  NAND3X0_HVT U430 ( .A1(n633), .A2(n632), .A3(n631), .Y(n_src_aox[13]) );
  AO222X1_HVT U431 ( .A1(n1850), .A2(sram_rdata_5[14]), .A3(n2110), .A4(
        sram_rdata_4[14]), .A5(sram_rdata_3[14]), .A6(n16601), .Y(n1306) );
  AO222X1_HVT U432 ( .A1(n1880), .A2(sram_rdata_2[14]), .A3(n16100), .A4(
        sram_rdata_1[14]), .A5(sram_rdata_0[14]), .A6(n16600), .Y(n934) );
  AOI22X1_HVT U433 ( .A1(n1306), .A2(n588), .A3(n5801), .A4(n934), .Y(n636) );
  OA22X1_HVT U434 ( .A1(n10300), .A2(n396), .A3(n2710), .A4(n3000), .Y(n635)
         );
  NAND2X0_HVT U435 ( .A1(n1760), .A2(sram_rdata_6[14]), .Y(n634) );
  NAND3X0_HVT U436 ( .A1(n636), .A2(n635), .A3(n634), .Y(n_src_aox[14]) );
  AO222X1_HVT U437 ( .A1(n1659), .A2(sram_rdata_5[15]), .A3(n15500), .A4(
        sram_rdata_4[15]), .A5(sram_rdata_3[15]), .A6(n16500), .Y(n1311) );
  AO222X1_HVT U438 ( .A1(n2070), .A2(sram_rdata_2[15]), .A3(n2160), .A4(
        sram_rdata_1[15]), .A5(sram_rdata_0[15]), .A6(n2020), .Y(n938) );
  AOI22X1_HVT U439 ( .A1(n1311), .A2(n14900), .A3(n579), .A4(n938), .Y(n639)
         );
  OA22X1_HVT U440 ( .A1(n12100), .A2(n397), .A3(n14700), .A4(n3010), .Y(n638)
         );
  NAND2X0_HVT U441 ( .A1(n2230), .A2(sram_rdata_6[15]), .Y(n637) );
  NAND3X0_HVT U442 ( .A1(n639), .A2(n638), .A3(n637), .Y(n_src_aox[15]) );
  AO222X1_HVT U443 ( .A1(n2080), .A2(sram_rdata_4[0]), .A3(n1960), .A4(
        sram_rdata_5[0]), .A5(n15500), .A6(sram_rdata_3[0]), .Y(n1315) );
  AO222X1_HVT U444 ( .A1(n2100), .A2(sram_rdata_1[0]), .A3(n13500), .A4(
        sram_rdata_0[0]), .A5(sram_rdata_2[0]), .A6(n1970), .Y(n942) );
  AOI22X1_HVT U445 ( .A1(n1315), .A2(n589), .A3(n5801), .A4(n942), .Y(n642) );
  OA22X1_HVT U446 ( .A1(n10400), .A2(n477), .A3(n2860), .A4(n2750), .Y(n641)
         );
  NAND2X0_HVT U447 ( .A1(n575), .A2(sram_rdata_8[0]), .Y(n6401) );
  NAND3X0_HVT U448 ( .A1(n642), .A2(n641), .A3(n6401), .Y(n_src_aox[16]) );
  AO222X1_HVT U449 ( .A1(n2090), .A2(sram_rdata_4[1]), .A3(n2130), .A4(
        sram_rdata_3[1]), .A5(sram_rdata_5[1]), .A6(n2010), .Y(n1318) );
  AO222X1_HVT U450 ( .A1(n2070), .A2(sram_rdata_1[1]), .A3(n2170), .A4(
        sram_rdata_0[1]), .A5(sram_rdata_2[1]), .A6(n1970), .Y(n946) );
  AOI22X1_HVT U451 ( .A1(n1318), .A2(n589), .A3(n5801), .A4(n946), .Y(n645) );
  OA22X1_HVT U452 ( .A1(n10500), .A2(n479), .A3(n2720), .A4(n383), .Y(n644) );
  NAND2X0_HVT U453 ( .A1(n1740), .A2(sram_rdata_8[1]), .Y(n643) );
  NAND3X0_HVT U454 ( .A1(n645), .A2(n644), .A3(n643), .Y(n_src_aox[17]) );
  AO222X1_HVT U455 ( .A1(n2040), .A2(sram_rdata_4[2]), .A3(n2160), .A4(
        sram_rdata_3[2]), .A5(sram_rdata_5[2]), .A6(n1960), .Y(n1323) );
  AO222X1_HVT U456 ( .A1(n1830), .A2(sram_rdata_1[2]), .A3(n2170), .A4(
        sram_rdata_0[2]), .A5(sram_rdata_2[2]), .A6(n1680), .Y(n9501) );
  AOI22X1_HVT U457 ( .A1(n1323), .A2(n12700), .A3(n11000), .A4(n9501), .Y(n648) );
  OA22X1_HVT U458 ( .A1(n2800), .A2(n4801), .A3(n2690), .A4(n384), .Y(n647) );
  NAND2X0_HVT U459 ( .A1(n1720), .A2(sram_rdata_8[2]), .Y(n646) );
  NAND3X0_HVT U460 ( .A1(n648), .A2(n647), .A3(n646), .Y(n_src_aox[18]) );
  AO222X1_HVT U461 ( .A1(n2060), .A2(sram_rdata_4[3]), .A3(n16000), .A4(
        sram_rdata_3[3]), .A5(sram_rdata_5[3]), .A6(n1930), .Y(n1328) );
  AO222X1_HVT U462 ( .A1(n2030), .A2(sram_rdata_1[3]), .A3(n2190), .A4(
        sram_rdata_0[3]), .A5(sram_rdata_2[3]), .A6(n16500), .Y(n954) );
  AOI22X1_HVT U463 ( .A1(n1328), .A2(n588), .A3(n582), .A4(n954), .Y(n651) );
  OA22X1_HVT U464 ( .A1(n2780), .A2(n481), .A3(n14600), .A4(n385), .Y(n6501)
         );
  NAND2X0_HVT U465 ( .A1(n1770), .A2(sram_rdata_8[3]), .Y(n649) );
  NAND3X0_HVT U466 ( .A1(n651), .A2(n6501), .A3(n649), .Y(n_src_aox[19]) );
  AO222X1_HVT U467 ( .A1(n2040), .A2(sram_rdata_4[4]), .A3(n13600), .A4(
        sram_rdata_3[4]), .A5(sram_rdata_5[4]), .A6(n1680), .Y(n1333) );
  AO222X1_HVT U468 ( .A1(n2050), .A2(sram_rdata_1[4]), .A3(n2140), .A4(
        sram_rdata_0[4]), .A5(sram_rdata_2[4]), .A6(n1670), .Y(n958) );
  AOI22X1_HVT U469 ( .A1(n1333), .A2(n15000), .A3(n579), .A4(n958), .Y(n654)
         );
  OA22X1_HVT U470 ( .A1(n10600), .A2(n482), .A3(n2730), .A4(n386), .Y(n653) );
  NAND2X0_HVT U471 ( .A1(n2250), .A2(sram_rdata_8[4]), .Y(n652) );
  NAND3X0_HVT U472 ( .A1(n654), .A2(n653), .A3(n652), .Y(n_src_aox[20]) );
  AO222X1_HVT U473 ( .A1(n1880), .A2(sram_rdata_4[5]), .A3(n2160), .A4(
        sram_rdata_3[5]), .A5(sram_rdata_5[5]), .A6(n1690), .Y(n1338) );
  AO222X1_HVT U474 ( .A1(n2030), .A2(sram_rdata_1[5]), .A3(n2170), .A4(
        sram_rdata_0[5]), .A5(sram_rdata_2[5]), .A6(n1680), .Y(n962) );
  AOI22X1_HVT U475 ( .A1(n1338), .A2(n10700), .A3(n10900), .A4(n962), .Y(n657)
         );
  OA22X1_HVT U476 ( .A1(n2790), .A2(n483), .A3(n14800), .A4(n387), .Y(n656) );
  NAND2X0_HVT U477 ( .A1(n576), .A2(sram_rdata_8[5]), .Y(n655) );
  NAND3X0_HVT U478 ( .A1(n657), .A2(n656), .A3(n655), .Y(n_src_aox[21]) );
  AO222X1_HVT U479 ( .A1(n2080), .A2(sram_rdata_4[6]), .A3(n13500), .A4(
        sram_rdata_3[6]), .A5(sram_rdata_5[6]), .A6(n16500), .Y(n1343) );
  AO222X1_HVT U480 ( .A1(n1850), .A2(sram_rdata_1[6]), .A3(n15400), .A4(
        sram_rdata_0[6]), .A5(sram_rdata_2[6]), .A6(n1700), .Y(n966) );
  AOI22X1_HVT U481 ( .A1(n1343), .A2(n15000), .A3(n582), .A4(n966), .Y(n6601)
         );
  OA22X1_HVT U482 ( .A1(n2790), .A2(n484), .A3(n2710), .A4(n388), .Y(n659) );
  NAND2X0_HVT U483 ( .A1(n2220), .A2(sram_rdata_8[6]), .Y(n658) );
  NAND3X0_HVT U484 ( .A1(n6601), .A2(n659), .A3(n658), .Y(n_src_aox[22]) );
  AO222X1_HVT U485 ( .A1(n1830), .A2(sram_rdata_4[7]), .A3(n15600), .A4(
        sram_rdata_3[7]), .A5(sram_rdata_5[7]), .A6(n2010), .Y(n1348) );
  AO222X1_HVT U486 ( .A1(n1840), .A2(sram_rdata_1[7]), .A3(n2160), .A4(
        sram_rdata_0[7]), .A5(sram_rdata_2[7]), .A6(n1960), .Y(n9701) );
  AOI22X1_HVT U487 ( .A1(n1348), .A2(n15000), .A3(n579), .A4(n9701), .Y(n663)
         );
  OA22X1_HVT U488 ( .A1(n2760), .A2(n485), .A3(n2700), .A4(n389), .Y(n662) );
  NAND2X0_HVT U489 ( .A1(n1770), .A2(sram_rdata_8[7]), .Y(n661) );
  NAND3X0_HVT U490 ( .A1(n663), .A2(n662), .A3(n661), .Y(n_src_aox[23]) );
  AO222X1_HVT U491 ( .A1(n2040), .A2(sram_rdata_4[8]), .A3(n587), .A4(
        sram_rdata_3[8]), .A5(sram_rdata_5[8]), .A6(n1940), .Y(n13501) );
  AO222X1_HVT U492 ( .A1(n1830), .A2(sram_rdata_1[8]), .A3(n2180), .A4(
        sram_rdata_0[8]), .A5(sram_rdata_2[8]), .A6(n2020), .Y(n974) );
  AOI22X1_HVT U493 ( .A1(n13501), .A2(n12700), .A3(n15200), .A4(n974), .Y(n666) );
  OA22X1_HVT U494 ( .A1(n2760), .A2(n486), .A3(n10100), .A4(n3901), .Y(n665)
         );
  NAND2X0_HVT U495 ( .A1(n1820), .A2(sram_rdata_8[8]), .Y(n664) );
  NAND3X0_HVT U496 ( .A1(n666), .A2(n665), .A3(n664), .Y(n_src_aox[24]) );
  AO222X1_HVT U497 ( .A1(n12500), .A2(sram_rdata_4[9]), .A3(n2120), .A4(
        sram_rdata_3[9]), .A5(sram_rdata_5[9]), .A6(n1970), .Y(n1355) );
  AO222X1_HVT U498 ( .A1(n1659), .A2(sram_rdata_1[9]), .A3(n15800), .A4(
        sram_rdata_0[9]), .A5(sram_rdata_2[9]), .A6(n1990), .Y(n978) );
  AOI22X1_HVT U499 ( .A1(n1355), .A2(n589), .A3(n12600), .A4(n978), .Y(n669)
         );
  OA22X1_HVT U500 ( .A1(n2810), .A2(n487), .A3(n2740), .A4(n391), .Y(n668) );
  NAND2X0_HVT U501 ( .A1(n1800), .A2(sram_rdata_8[9]), .Y(n667) );
  NAND3X0_HVT U502 ( .A1(n669), .A2(n668), .A3(n667), .Y(n_src_aox[25]) );
  AO222X1_HVT U503 ( .A1(n1890), .A2(sram_rdata_4[10]), .A3(n2170), .A4(
        sram_rdata_3[10]), .A5(sram_rdata_5[10]), .A6(n1920), .Y(n13601) );
  AO222X1_HVT U504 ( .A1(n1830), .A2(sram_rdata_1[10]), .A3(n2130), .A4(
        sram_rdata_0[10]), .A5(sram_rdata_2[10]), .A6(n1940), .Y(n982) );
  AOI22X1_HVT U505 ( .A1(n13601), .A2(n10700), .A3(n12900), .A4(n982), .Y(n672) );
  OA22X1_HVT U506 ( .A1(n10500), .A2(n488), .A3(n2700), .A4(n392), .Y(n671) );
  NAND2X0_HVT U507 ( .A1(n1790), .A2(sram_rdata_8[10]), .Y(n6701) );
  NAND3X0_HVT U508 ( .A1(n672), .A2(n671), .A3(n6701), .Y(n_src_aox[26]) );
  AO222X1_HVT U509 ( .A1(n1910), .A2(sram_rdata_4[11]), .A3(n2130), .A4(
        sram_rdata_3[11]), .A5(sram_rdata_5[11]), .A6(n1680), .Y(n1365) );
  AO222X1_HVT U510 ( .A1(n12500), .A2(sram_rdata_1[11]), .A3(n2110), .A4(
        sram_rdata_0[11]), .A5(sram_rdata_2[11]), .A6(n1970), .Y(n986) );
  AOI22X1_HVT U511 ( .A1(n1365), .A2(n588), .A3(n15100), .A4(n986), .Y(n675)
         );
  OA22X1_HVT U512 ( .A1(n10600), .A2(n489), .A3(n11500), .A4(n393), .Y(n674)
         );
  NAND2X0_HVT U513 ( .A1(n2270), .A2(sram_rdata_8[11]), .Y(n673) );
  NAND3X0_HVT U514 ( .A1(n675), .A2(n674), .A3(n673), .Y(n_src_aox[27]) );
  AO222X1_HVT U515 ( .A1(n2080), .A2(sram_rdata_4[12]), .A3(n2110), .A4(
        sram_rdata_3[12]), .A5(sram_rdata_5[12]), .A6(n1920), .Y(n13701) );
  AO222X1_HVT U516 ( .A1(n1880), .A2(sram_rdata_1[12]), .A3(n587), .A4(
        sram_rdata_0[12]), .A5(sram_rdata_2[12]), .A6(n1700), .Y(n9901) );
  AOI22X1_HVT U517 ( .A1(n13701), .A2(n10700), .A3(n11000), .A4(n9901), .Y(
        n678) );
  OA22X1_HVT U518 ( .A1(n2770), .A2(n4901), .A3(n14800), .A4(n394), .Y(n677)
         );
  NAND2X0_HVT U519 ( .A1(n1820), .A2(sram_rdata_8[12]), .Y(n676) );
  NAND3X0_HVT U520 ( .A1(n678), .A2(n677), .A3(n676), .Y(n_src_aox[28]) );
  AO222X1_HVT U521 ( .A1(n1830), .A2(sram_rdata_4[13]), .A3(n16100), .A4(
        sram_rdata_3[13]), .A5(sram_rdata_5[13]), .A6(n2000), .Y(n1375) );
  AO222X1_HVT U522 ( .A1(n1840), .A2(sram_rdata_1[13]), .A3(n2180), .A4(
        sram_rdata_0[13]), .A5(sram_rdata_2[13]), .A6(n1980), .Y(n994) );
  AOI22X1_HVT U523 ( .A1(n1375), .A2(n15000), .A3(n582), .A4(n994), .Y(n681)
         );
  OA22X1_HVT U524 ( .A1(n10400), .A2(n491), .A3(n2740), .A4(n395), .Y(n6801)
         );
  NAND2X0_HVT U525 ( .A1(n1730), .A2(sram_rdata_8[13]), .Y(n679) );
  NAND3X0_HVT U526 ( .A1(n681), .A2(n6801), .A3(n679), .Y(n_src_aox[29]) );
  AO222X1_HVT U527 ( .A1(n2030), .A2(sram_rdata_4[14]), .A3(n15600), .A4(
        sram_rdata_3[14]), .A5(sram_rdata_5[14]), .A6(n1990), .Y(n13801) );
  AO222X1_HVT U528 ( .A1(n1860), .A2(sram_rdata_1[14]), .A3(n2190), .A4(
        sram_rdata_0[14]), .A5(sram_rdata_2[14]), .A6(n1930), .Y(n998) );
  AOI22X1_HVT U529 ( .A1(n13801), .A2(n10800), .A3(n15100), .A4(n998), .Y(n684) );
  OA22X1_HVT U530 ( .A1(n12000), .A2(n492), .A3(n2690), .A4(n396), .Y(n683) );
  NAND2X0_HVT U531 ( .A1(n2210), .A2(sram_rdata_8[14]), .Y(n682) );
  NAND3X0_HVT U532 ( .A1(n684), .A2(n683), .A3(n682), .Y(n_src_aox[30]) );
  AO222X1_HVT U533 ( .A1(n1860), .A2(sram_rdata_4[15]), .A3(n15400), .A4(
        sram_rdata_3[15]), .A5(sram_rdata_5[15]), .A6(n16601), .Y(n1385) );
  AO222X1_HVT U534 ( .A1(n1860), .A2(sram_rdata_1[15]), .A3(n15600), .A4(
        sram_rdata_0[15]), .A5(sram_rdata_2[15]), .A6(n16600), .Y(n1002) );
  AOI22X1_HVT U535 ( .A1(n1385), .A2(n10700), .A3(n579), .A4(n1002), .Y(n687)
         );
  OA22X1_HVT U536 ( .A1(n12100), .A2(n493), .A3(n14500), .A4(n397), .Y(n686)
         );
  NAND2X0_HVT U537 ( .A1(n2230), .A2(sram_rdata_8[15]), .Y(n685) );
  NAND3X0_HVT U538 ( .A1(n687), .A2(n686), .A3(n685), .Y(n_src_aox[31]) );
  AO222X1_HVT U539 ( .A1(n1860), .A2(sram_rdata_3[0]), .A3(n1920), .A4(
        sram_rdata_4[0]), .A5(n2160), .A6(sram_rdata_5[0]), .Y(n1389) );
  AO222X1_HVT U540 ( .A1(n1900), .A2(sram_rdata_0[0]), .A3(n15400), .A4(
        sram_rdata_2[0]), .A5(n2000), .A6(sram_rdata_1[0]), .Y(n1006) );
  AOI22X1_HVT U541 ( .A1(n1389), .A2(n591), .A3(n5801), .A4(n1006), .Y(n6901)
         );
  OA22X1_HVT U542 ( .A1(n10300), .A2(n573), .A3(n477), .A4(n10100), .Y(n689)
         );
  NAND2X0_HVT U543 ( .A1(n1810), .A2(sram_rdata_7[0]), .Y(n688) );
  NAND3X0_HVT U544 ( .A1(n6901), .A2(n689), .A3(n688), .Y(n_src_aox[32]) );
  AO222X1_HVT U545 ( .A1(n1910), .A2(sram_rdata_3[1]), .A3(n2140), .A4(
        sram_rdata_5[1]), .A5(n1980), .A6(sram_rdata_4[1]), .Y(n1392) );
  AO222X1_HVT U546 ( .A1(n1900), .A2(sram_rdata_0[1]), .A3(n15600), .A4(
        sram_rdata_2[1]), .A5(n1710), .A6(sram_rdata_1[1]), .Y(n10101) );
  AOI22X1_HVT U547 ( .A1(n1392), .A2(n591), .A3(n1648), .A4(n10101), .Y(n693)
         );
  OA22X1_HVT U548 ( .A1(n10500), .A2(n2870), .A3(n14700), .A4(n479), .Y(n692)
         );
  NAND2X0_HVT U549 ( .A1(n576), .A2(sram_rdata_7[1]), .Y(n691) );
  NAND3X0_HVT U550 ( .A1(n693), .A2(n692), .A3(n691), .Y(n_src_aox[33]) );
  AO222X1_HVT U551 ( .A1(n2080), .A2(sram_rdata_3[2]), .A3(n15700), .A4(
        sram_rdata_5[2]), .A5(n1680), .A6(sram_rdata_4[2]), .Y(n1397) );
  AO222X1_HVT U552 ( .A1(n2090), .A2(sram_rdata_0[2]), .A3(n2180), .A4(
        sram_rdata_2[2]), .A5(n16601), .A6(sram_rdata_1[2]), .Y(n1011) );
  AOI22X1_HVT U553 ( .A1(n1397), .A2(n588), .A3(n5801), .A4(n1011), .Y(n696)
         );
  OA22X1_HVT U554 ( .A1(n10300), .A2(n2880), .A3(n10100), .A4(n4801), .Y(n695)
         );
  NAND2X0_HVT U555 ( .A1(n2260), .A2(sram_rdata_7[2]), .Y(n694) );
  NAND3X0_HVT U556 ( .A1(n696), .A2(n695), .A3(n694), .Y(n_src_aox[34]) );
  AO222X1_HVT U557 ( .A1(n2070), .A2(sram_rdata_3[3]), .A3(n15500), .A4(
        sram_rdata_5[3]), .A5(n1960), .A6(sram_rdata_4[3]), .Y(n1402) );
  AO222X1_HVT U558 ( .A1(n2090), .A2(sram_rdata_0[3]), .A3(n15700), .A4(
        sram_rdata_2[3]), .A5(n1940), .A6(sram_rdata_1[3]), .Y(n1015) );
  AOI22X1_HVT U559 ( .A1(n1402), .A2(n15000), .A3(n15200), .A4(n1015), .Y(n699) );
  OA22X1_HVT U560 ( .A1(n2770), .A2(n2890), .A3(n2700), .A4(n481), .Y(n698) );
  NAND2X0_HVT U561 ( .A1(n2280), .A2(sram_rdata_7[3]), .Y(n697) );
  NAND3X0_HVT U562 ( .A1(n699), .A2(n698), .A3(n697), .Y(n_src_aox[35]) );
  AO222X1_HVT U563 ( .A1(n2050), .A2(sram_rdata_3[4]), .A3(n2190), .A4(
        sram_rdata_5[4]), .A5(n1670), .A6(sram_rdata_4[4]), .Y(n1407) );
  AO222X1_HVT U564 ( .A1(n1910), .A2(sram_rdata_0[4]), .A3(n2190), .A4(
        sram_rdata_2[4]), .A5(n1980), .A6(sram_rdata_1[4]), .Y(n1019) );
  AOI22X1_HVT U565 ( .A1(n1407), .A2(n10800), .A3(n12900), .A4(n1019), .Y(n702) );
  OA22X1_HVT U566 ( .A1(n2810), .A2(n2900), .A3(n14600), .A4(n482), .Y(n701)
         );
  NAND2X0_HVT U567 ( .A1(n1730), .A2(sram_rdata_7[4]), .Y(n7001) );
  NAND3X0_HVT U568 ( .A1(n702), .A2(n701), .A3(n7001), .Y(n_src_aox[36]) );
  AO222X1_HVT U569 ( .A1(n1840), .A2(sram_rdata_3[5]), .A3(n2190), .A4(
        sram_rdata_5[5]), .A5(n1990), .A6(sram_rdata_4[5]), .Y(n1412) );
  AO222X1_HVT U570 ( .A1(n2060), .A2(sram_rdata_0[5]), .A3(n13600), .A4(
        sram_rdata_2[5]), .A5(n1960), .A6(sram_rdata_1[5]), .Y(n1023) );
  AOI22X1_HVT U571 ( .A1(n1412), .A2(n14900), .A3(n582), .A4(n1023), .Y(n705)
         );
  OA22X1_HVT U572 ( .A1(n13800), .A2(n2910), .A3(n2730), .A4(n483), .Y(n704)
         );
  NAND2X0_HVT U573 ( .A1(n2240), .A2(sram_rdata_7[5]), .Y(n703) );
  NAND3X0_HVT U574 ( .A1(n705), .A2(n704), .A3(n703), .Y(n_src_aox[37]) );
  AO222X1_HVT U575 ( .A1(n2030), .A2(sram_rdata_3[6]), .A3(n587), .A4(
        sram_rdata_5[6]), .A5(n1960), .A6(sram_rdata_4[6]), .Y(n1417) );
  AO222X1_HVT U576 ( .A1(n2040), .A2(sram_rdata_0[6]), .A3(n16000), .A4(
        sram_rdata_2[6]), .A5(n16601), .A6(sram_rdata_1[6]), .Y(n1027) );
  AOI22X1_HVT U577 ( .A1(n1417), .A2(n15000), .A3(n582), .A4(n1027), .Y(n708)
         );
  OA22X1_HVT U578 ( .A1(n10600), .A2(n2920), .A3(n2730), .A4(n484), .Y(n707)
         );
  NAND2X0_HVT U579 ( .A1(n1770), .A2(sram_rdata_7[6]), .Y(n706) );
  NAND3X0_HVT U580 ( .A1(n708), .A2(n707), .A3(n706), .Y(n_src_aox[38]) );
  AO222X1_HVT U581 ( .A1(n12500), .A2(sram_rdata_3[7]), .A3(n2110), .A4(
        sram_rdata_5[7]), .A5(n16601), .A6(sram_rdata_4[7]), .Y(n1419) );
  AO222X1_HVT U582 ( .A1(n1659), .A2(sram_rdata_0[7]), .A3(n13600), .A4(
        sram_rdata_2[7]), .A5(n16600), .A6(sram_rdata_1[7]), .Y(n1031) );
  AOI22X1_HVT U583 ( .A1(n1419), .A2(n14900), .A3(n5801), .A4(n1031), .Y(n711)
         );
  OA22X1_HVT U584 ( .A1(n1662), .A2(n2930), .A3(n10000), .A4(n485), .Y(n7101)
         );
  NAND2X0_HVT U585 ( .A1(n1730), .A2(sram_rdata_7[7]), .Y(n709) );
  NAND3X0_HVT U586 ( .A1(n711), .A2(n7101), .A3(n709), .Y(n_src_aox[39]) );
  AO222X1_HVT U587 ( .A1(n2070), .A2(sram_rdata_3[8]), .A3(n16000), .A4(
        sram_rdata_5[8]), .A5(n16600), .A6(sram_rdata_4[8]), .Y(n1424) );
  AO222X1_HVT U588 ( .A1(n1860), .A2(sram_rdata_0[8]), .A3(n13600), .A4(
        sram_rdata_2[8]), .A5(n16500), .A6(sram_rdata_1[8]), .Y(n1035) );
  AOI22X1_HVT U589 ( .A1(n1424), .A2(n588), .A3(n582), .A4(n1035), .Y(n714) );
  OA22X1_HVT U590 ( .A1(n13700), .A2(n2940), .A3(n14500), .A4(n486), .Y(n713)
         );
  NAND2X0_HVT U591 ( .A1(n1800), .A2(sram_rdata_7[8]), .Y(n712) );
  NAND3X0_HVT U592 ( .A1(n714), .A2(n713), .A3(n712), .Y(n_src_aox[40]) );
  AO222X1_HVT U593 ( .A1(n2090), .A2(sram_rdata_3[9]), .A3(n15800), .A4(
        sram_rdata_5[9]), .A5(n1700), .A6(sram_rdata_4[9]), .Y(n1429) );
  AO222X1_HVT U594 ( .A1(n1900), .A2(sram_rdata_0[9]), .A3(n15500), .A4(
        sram_rdata_2[9]), .A5(n2000), .A6(sram_rdata_1[9]), .Y(n1039) );
  AOI22X1_HVT U595 ( .A1(n1429), .A2(n10700), .A3(n581), .A4(n1039), .Y(n717)
         );
  OA22X1_HVT U596 ( .A1(n2800), .A2(n2950), .A3(n14800), .A4(n487), .Y(n716)
         );
  NAND2X0_HVT U597 ( .A1(n576), .A2(sram_rdata_7[9]), .Y(n715) );
  NAND3X0_HVT U598 ( .A1(n717), .A2(n716), .A3(n715), .Y(n_src_aox[41]) );
  AO222X1_HVT U599 ( .A1(n2060), .A2(sram_rdata_3[10]), .A3(n2170), .A4(
        sram_rdata_5[10]), .A5(n1980), .A6(sram_rdata_4[10]), .Y(n1434) );
  AO222X1_HVT U600 ( .A1(n1659), .A2(sram_rdata_0[10]), .A3(n15600), .A4(
        sram_rdata_2[10]), .A5(n2000), .A6(sram_rdata_1[10]), .Y(n1043) );
  AOI22X1_HVT U601 ( .A1(n1434), .A2(n12700), .A3(n15100), .A4(n1043), .Y(
        n7201) );
  OA22X1_HVT U602 ( .A1(n1662), .A2(n2960), .A3(n14700), .A4(n488), .Y(n719)
         );
  NAND2X0_HVT U603 ( .A1(n2250), .A2(sram_rdata_7[10]), .Y(n718) );
  NAND3X0_HVT U604 ( .A1(n7201), .A2(n719), .A3(n718), .Y(n_src_aox[42]) );
  AO222X1_HVT U605 ( .A1(n1880), .A2(sram_rdata_3[11]), .A3(n587), .A4(
        sram_rdata_5[11]), .A5(n1970), .A6(sram_rdata_4[11]), .Y(n1439) );
  AO222X1_HVT U606 ( .A1(n1840), .A2(sram_rdata_0[11]), .A3(n2140), .A4(
        sram_rdata_2[11]), .A5(n1930), .A6(sram_rdata_1[11]), .Y(n1047) );
  AOI22X1_HVT U607 ( .A1(n1439), .A2(n592), .A3(n582), .A4(n1047), .Y(n723) );
  OA22X1_HVT U608 ( .A1(n11800), .A2(n2970), .A3(n2690), .A4(n489), .Y(n722)
         );
  NAND2X0_HVT U609 ( .A1(n1760), .A2(sram_rdata_7[11]), .Y(n721) );
  NAND3X0_HVT U610 ( .A1(n723), .A2(n722), .A3(n721), .Y(n_src_aox[43]) );
  AO222X1_HVT U611 ( .A1(n1850), .A2(sram_rdata_3[12]), .A3(n15900), .A4(
        sram_rdata_5[12]), .A5(n16500), .A6(sram_rdata_4[12]), .Y(n1444) );
  AO222X1_HVT U612 ( .A1(n1880), .A2(sram_rdata_0[12]), .A3(n13600), .A4(
        sram_rdata_2[12]), .A5(n1930), .A6(sram_rdata_1[12]), .Y(n1051) );
  AOI22X1_HVT U613 ( .A1(n1444), .A2(n15000), .A3(n12900), .A4(n1051), .Y(n726) );
  OA22X1_HVT U614 ( .A1(n10500), .A2(n2980), .A3(n10000), .A4(n4901), .Y(n725)
         );
  NAND2X0_HVT U615 ( .A1(n2220), .A2(sram_rdata_7[12]), .Y(n724) );
  NAND3X0_HVT U616 ( .A1(n726), .A2(n725), .A3(n724), .Y(n_src_aox[44]) );
  AO222X1_HVT U617 ( .A1(n1900), .A2(sram_rdata_3[13]), .A3(n2120), .A4(
        sram_rdata_5[13]), .A5(n16400), .A6(sram_rdata_4[13]), .Y(n1449) );
  AO222X1_HVT U618 ( .A1(n1890), .A2(sram_rdata_0[13]), .A3(n2110), .A4(
        sram_rdata_2[13]), .A5(n16601), .A6(sram_rdata_1[13]), .Y(n1055) );
  AOI22X1_HVT U619 ( .A1(n1449), .A2(n15000), .A3(n10900), .A4(n1055), .Y(n729) );
  OA22X1_HVT U620 ( .A1(n12000), .A2(n2990), .A3(n2720), .A4(n491), .Y(n728)
         );
  NAND2X0_HVT U621 ( .A1(n1750), .A2(sram_rdata_7[13]), .Y(n727) );
  NAND3X0_HVT U622 ( .A1(n729), .A2(n728), .A3(n727), .Y(n_src_aox[45]) );
  AO222X1_HVT U623 ( .A1(n2070), .A2(sram_rdata_3[14]), .A3(n2140), .A4(
        sram_rdata_5[14]), .A5(n16400), .A6(sram_rdata_4[14]), .Y(n1454) );
  AO222X1_HVT U624 ( .A1(n13900), .A2(sram_rdata_0[14]), .A3(n15700), .A4(
        sram_rdata_2[14]), .A5(n16500), .A6(sram_rdata_1[14]), .Y(n1059) );
  AOI22X1_HVT U625 ( .A1(n1454), .A2(n589), .A3(n11000), .A4(n1059), .Y(n732)
         );
  OA22X1_HVT U626 ( .A1(n2780), .A2(n3000), .A3(n2720), .A4(n492), .Y(n731) );
  NAND2X0_HVT U627 ( .A1(n1740), .A2(sram_rdata_7[14]), .Y(n7301) );
  NAND3X0_HVT U628 ( .A1(n732), .A2(n731), .A3(n7301), .Y(n_src_aox[46]) );
  AO222X1_HVT U629 ( .A1(n1659), .A2(sram_rdata_3[15]), .A3(n13600), .A4(
        sram_rdata_5[15]), .A5(n16601), .A6(sram_rdata_4[15]), .Y(n1456) );
  AO222X1_HVT U630 ( .A1(n1890), .A2(sram_rdata_0[15]), .A3(n15400), .A4(
        sram_rdata_2[15]), .A5(n1680), .A6(sram_rdata_1[15]), .Y(n1063) );
  AOI22X1_HVT U631 ( .A1(n1456), .A2(n591), .A3(n10900), .A4(n1063), .Y(n735)
         );
  OA22X1_HVT U632 ( .A1(n12100), .A2(n3010), .A3(n14600), .A4(n493), .Y(n734)
         );
  NAND2X0_HVT U633 ( .A1(n2210), .A2(sram_rdata_7[15]), .Y(n733) );
  NAND3X0_HVT U634 ( .A1(n735), .A2(n734), .A3(n733), .Y(n_src_aox[47]) );
  AO222X1_HVT U635 ( .A1(n2040), .A2(sram_rdata_5[16]), .A3(n2180), .A4(
        sram_rdata_4[16]), .A5(sram_rdata_3[16]), .A6(n16601), .Y(n1461) );
  AO222X1_HVT U636 ( .A1(n1910), .A2(sram_rdata_2[16]), .A3(n15400), .A4(
        sram_rdata_1[16]), .A5(sram_rdata_0[16]), .A6(n16500), .Y(n1067) );
  AOI22X1_HVT U637 ( .A1(n1461), .A2(n10800), .A3(n15200), .A4(n1067), .Y(n738) );
  OA22X1_HVT U638 ( .A1(n12000), .A2(n398), .A3(n10000), .A4(n3020), .Y(n737)
         );
  NAND2X0_HVT U639 ( .A1(n1730), .A2(sram_rdata_6[16]), .Y(n736) );
  NAND3X0_HVT U640 ( .A1(n738), .A2(n737), .A3(n736), .Y(n_src_aox[48]) );
  AO222X1_HVT U641 ( .A1(n1659), .A2(sram_rdata_5[17]), .A3(n15600), .A4(
        sram_rdata_4[17]), .A5(sram_rdata_3[17]), .A6(n1670), .Y(n1466) );
  AO222X1_HVT U642 ( .A1(n12500), .A2(sram_rdata_2[17]), .A3(n15500), .A4(
        sram_rdata_1[17]), .A5(sram_rdata_0[17]), .A6(n1690), .Y(n1071) );
  AOI22X1_HVT U643 ( .A1(n1466), .A2(n588), .A3(n15200), .A4(n1071), .Y(n741)
         );
  OA22X1_HVT U644 ( .A1(n11900), .A2(n399), .A3(n10100), .A4(n3030), .Y(n7401)
         );
  NAND2X0_HVT U645 ( .A1(n2280), .A2(sram_rdata_6[17]), .Y(n739) );
  NAND3X0_HVT U646 ( .A1(n741), .A2(n7401), .A3(n739), .Y(n_src_aox[49]) );
  AO222X1_HVT U647 ( .A1(n1890), .A2(sram_rdata_5[18]), .A3(n587), .A4(
        sram_rdata_4[18]), .A5(sram_rdata_3[18]), .A6(n2020), .Y(n1471) );
  AO222X1_HVT U648 ( .A1(n2040), .A2(sram_rdata_2[18]), .A3(n587), .A4(
        sram_rdata_1[18]), .A5(sram_rdata_0[18]), .A6(n1960), .Y(n1075) );
  AOI22X1_HVT U649 ( .A1(n1471), .A2(n589), .A3(n12600), .A4(n1075), .Y(n744)
         );
  OA22X1_HVT U650 ( .A1(n12100), .A2(n4001), .A3(n2730), .A4(n3040), .Y(n743)
         );
  NAND2X0_HVT U651 ( .A1(n1790), .A2(sram_rdata_6[18]), .Y(n742) );
  NAND3X0_HVT U652 ( .A1(n744), .A2(n743), .A3(n742), .Y(n_src_aox[50]) );
  AO222X1_HVT U653 ( .A1(n1910), .A2(sram_rdata_5[19]), .A3(n2140), .A4(
        sram_rdata_4[19]), .A5(sram_rdata_3[19]), .A6(n2020), .Y(n1476) );
  AO222X1_HVT U654 ( .A1(n1890), .A2(sram_rdata_2[19]), .A3(n15400), .A4(
        sram_rdata_1[19]), .A5(sram_rdata_0[19]), .A6(n1980), .Y(n1079) );
  AOI22X1_HVT U655 ( .A1(n1476), .A2(n14900), .A3(n578), .A4(n1079), .Y(n747)
         );
  OA22X1_HVT U656 ( .A1(n2780), .A2(n401), .A3(n11500), .A4(n3050), .Y(n746)
         );
  NAND2X0_HVT U657 ( .A1(n2230), .A2(sram_rdata_6[19]), .Y(n745) );
  NAND3X0_HVT U658 ( .A1(n747), .A2(n746), .A3(n745), .Y(n_src_aox[51]) );
  AO222X1_HVT U659 ( .A1(n2100), .A2(sram_rdata_5[20]), .A3(n16100), .A4(
        sram_rdata_4[20]), .A5(sram_rdata_3[20]), .A6(n1990), .Y(n1481) );
  AO222X1_HVT U660 ( .A1(n2100), .A2(sram_rdata_2[20]), .A3(n2190), .A4(
        sram_rdata_1[20]), .A5(sram_rdata_0[20]), .A6(n1670), .Y(n1083) );
  AOI22X1_HVT U661 ( .A1(n1481), .A2(n15000), .A3(n12600), .A4(n1083), .Y(
        n7501) );
  OA22X1_HVT U662 ( .A1(n2810), .A2(n402), .A3(n2700), .A4(n3060), .Y(n749) );
  NAND2X0_HVT U663 ( .A1(n2250), .A2(sram_rdata_6[20]), .Y(n748) );
  NAND3X0_HVT U664 ( .A1(n7501), .A2(n749), .A3(n748), .Y(n_src_aox[52]) );
  AO222X1_HVT U665 ( .A1(n2100), .A2(sram_rdata_5[21]), .A3(n2170), .A4(
        sram_rdata_4[21]), .A5(sram_rdata_3[21]), .A6(n1930), .Y(n1486) );
  AO222X1_HVT U666 ( .A1(n2080), .A2(sram_rdata_2[21]), .A3(n16000), .A4(
        sram_rdata_1[21]), .A5(sram_rdata_0[21]), .A6(n1920), .Y(n1087) );
  AOI22X1_HVT U667 ( .A1(n1486), .A2(n589), .A3(n12600), .A4(n1087), .Y(n753)
         );
  OA22X1_HVT U668 ( .A1(n2790), .A2(n403), .A3(n2740), .A4(n3070), .Y(n752) );
  NAND2X0_HVT U669 ( .A1(n1770), .A2(sram_rdata_6[21]), .Y(n751) );
  NAND3X0_HVT U670 ( .A1(n753), .A2(n752), .A3(n751), .Y(n_src_aox[53]) );
  AO222X1_HVT U671 ( .A1(n2060), .A2(sram_rdata_5[22]), .A3(n2170), .A4(
        sram_rdata_4[22]), .A5(sram_rdata_3[22]), .A6(n1680), .Y(n1491) );
  AO222X1_HVT U672 ( .A1(n12500), .A2(sram_rdata_2[22]), .A3(n2160), .A4(
        sram_rdata_1[22]), .A5(sram_rdata_0[22]), .A6(n16400), .Y(n1091) );
  AOI22X1_HVT U673 ( .A1(n1491), .A2(n12700), .A3(n12900), .A4(n1091), .Y(n756) );
  OA22X1_HVT U674 ( .A1(n10600), .A2(n404), .A3(n1661), .A4(n3080), .Y(n755)
         );
  NAND2X0_HVT U675 ( .A1(n576), .A2(sram_rdata_6[22]), .Y(n754) );
  NAND3X0_HVT U676 ( .A1(n756), .A2(n755), .A3(n754), .Y(n_src_aox[54]) );
  AO222X1_HVT U677 ( .A1(n1850), .A2(sram_rdata_5[23]), .A3(n2180), .A4(
        sram_rdata_4[23]), .A5(sram_rdata_3[23]), .A6(n1670), .Y(n1496) );
  AO222X1_HVT U678 ( .A1(n2050), .A2(sram_rdata_2[23]), .A3(n15800), .A4(
        sram_rdata_1[23]), .A5(sram_rdata_0[23]), .A6(n1710), .Y(n1095) );
  AOI22X1_HVT U679 ( .A1(n1496), .A2(n588), .A3(n5801), .A4(n1095), .Y(n759)
         );
  OA22X1_HVT U680 ( .A1(n1662), .A2(n405), .A3(n14500), .A4(n3090), .Y(n758)
         );
  NAND2X0_HVT U681 ( .A1(n1760), .A2(sram_rdata_6[23]), .Y(n757) );
  NAND3X0_HVT U682 ( .A1(n759), .A2(n758), .A3(n757), .Y(n_src_aox[55]) );
  AO222X1_HVT U683 ( .A1(n2030), .A2(sram_rdata_5[24]), .A3(n13600), .A4(
        sram_rdata_4[24]), .A5(sram_rdata_3[24]), .A6(n16600), .Y(n1501) );
  AO222X1_HVT U684 ( .A1(n2040), .A2(sram_rdata_2[24]), .A3(n13600), .A4(
        sram_rdata_1[24]), .A5(sram_rdata_0[24]), .A6(n16600), .Y(n1099) );
  AOI22X1_HVT U685 ( .A1(n1501), .A2(n15000), .A3(n582), .A4(n1099), .Y(n762)
         );
  OA22X1_HVT U686 ( .A1(n13800), .A2(n406), .A3(n14600), .A4(n3100), .Y(n761)
         );
  NAND2X0_HVT U687 ( .A1(n2270), .A2(sram_rdata_6[24]), .Y(n7601) );
  NAND3X0_HVT U688 ( .A1(n762), .A2(n761), .A3(n7601), .Y(n_src_aox[56]) );
  AO222X1_HVT U689 ( .A1(n2040), .A2(sram_rdata_5[25]), .A3(n2130), .A4(
        sram_rdata_4[25]), .A5(sram_rdata_3[25]), .A6(n2010), .Y(n1503) );
  AO222X1_HVT U690 ( .A1(n2050), .A2(sram_rdata_2[25]), .A3(n587), .A4(
        sram_rdata_1[25]), .A5(sram_rdata_0[25]), .A6(n1990), .Y(n1103) );
  AOI22X1_HVT U691 ( .A1(n1503), .A2(n12800), .A3(n579), .A4(n1103), .Y(n765)
         );
  OA22X1_HVT U692 ( .A1(n13800), .A2(n407), .A3(n2750), .A4(n3110), .Y(n764)
         );
  NAND2X0_HVT U693 ( .A1(n1810), .A2(sram_rdata_6[25]), .Y(n763) );
  NAND3X0_HVT U694 ( .A1(n765), .A2(n764), .A3(n763), .Y(n_src_aox[57]) );
  AO222X1_HVT U695 ( .A1(n2100), .A2(sram_rdata_5[26]), .A3(n15400), .A4(
        sram_rdata_4[26]), .A5(sram_rdata_3[26]), .A6(n1940), .Y(n1508) );
  AO222X1_HVT U696 ( .A1(n1910), .A2(sram_rdata_2[26]), .A3(n15400), .A4(
        sram_rdata_1[26]), .A5(sram_rdata_0[26]), .A6(n2000), .Y(n1107) );
  AOI22X1_HVT U697 ( .A1(n1508), .A2(n591), .A3(n579), .A4(n1107), .Y(n768) );
  OA22X1_HVT U698 ( .A1(n2760), .A2(n408), .A3(n2740), .A4(n3120), .Y(n767) );
  NAND2X0_HVT U699 ( .A1(n2220), .A2(sram_rdata_6[26]), .Y(n766) );
  NAND3X0_HVT U700 ( .A1(n768), .A2(n767), .A3(n766), .Y(n_src_aox[58]) );
  AO222X1_HVT U701 ( .A1(n1830), .A2(sram_rdata_5[27]), .A3(n16000), .A4(
        sram_rdata_4[27]), .A5(sram_rdata_3[27]), .A6(n1970), .Y(n1513) );
  AO222X1_HVT U702 ( .A1(n1880), .A2(sram_rdata_2[27]), .A3(n13500), .A4(
        sram_rdata_1[27]), .A5(sram_rdata_0[27]), .A6(n1960), .Y(n1108) );
  AOI22X1_HVT U703 ( .A1(n1513), .A2(n591), .A3(n1648), .A4(n1108), .Y(n771)
         );
  OA22X1_HVT U704 ( .A1(n11800), .A2(n409), .A3(n10000), .A4(n3130), .Y(n7701)
         );
  NAND2X0_HVT U705 ( .A1(n576), .A2(sram_rdata_6[27]), .Y(n769) );
  NAND3X0_HVT U706 ( .A1(n771), .A2(n7701), .A3(n769), .Y(n_src_aox[59]) );
  AO222X1_HVT U707 ( .A1(n2030), .A2(sram_rdata_5[28]), .A3(n2160), .A4(
        sram_rdata_4[28]), .A5(sram_rdata_3[28]), .A6(n1710), .Y(n1515) );
  AO222X1_HVT U708 ( .A1(n13900), .A2(sram_rdata_2[28]), .A3(n2190), .A4(
        sram_rdata_1[28]), .A5(sram_rdata_0[28]), .A6(n1680), .Y(n1112) );
  AOI22X1_HVT U709 ( .A1(n1515), .A2(n12700), .A3(n15200), .A4(n1112), .Y(n774) );
  OA22X1_HVT U710 ( .A1(n10500), .A2(n4101), .A3(n2710), .A4(n3140), .Y(n773)
         );
  NAND2X0_HVT U711 ( .A1(n1810), .A2(sram_rdata_6[28]), .Y(n772) );
  NAND3X0_HVT U712 ( .A1(n774), .A2(n773), .A3(n772), .Y(n_src_aox[60]) );
  AO222X1_HVT U713 ( .A1(n13900), .A2(sram_rdata_5[29]), .A3(n13500), .A4(
        sram_rdata_4[29]), .A5(sram_rdata_3[29]), .A6(n1700), .Y(n15201) );
  AO222X1_HVT U714 ( .A1(n1850), .A2(sram_rdata_2[29]), .A3(n2110), .A4(
        sram_rdata_1[29]), .A5(sram_rdata_0[29]), .A6(n1980), .Y(n1116) );
  AOI22X1_HVT U715 ( .A1(n15201), .A2(n14900), .A3(n581), .A4(n1116), .Y(n778)
         );
  OA22X1_HVT U716 ( .A1(n10400), .A2(n411), .A3(n14700), .A4(n3150), .Y(n777)
         );
  NAND2X0_HVT U717 ( .A1(n1790), .A2(sram_rdata_6[29]), .Y(n775) );
  NAND3X0_HVT U718 ( .A1(n778), .A2(n777), .A3(n775), .Y(n_src_aox[61]) );
  AO222X1_HVT U719 ( .A1(n1850), .A2(sram_rdata_5[30]), .A3(n587), .A4(
        sram_rdata_4[30]), .A5(sram_rdata_3[30]), .A6(n1920), .Y(n1525) );
  AO222X1_HVT U720 ( .A1(n1860), .A2(sram_rdata_2[30]), .A3(n15500), .A4(
        sram_rdata_1[30]), .A5(sram_rdata_0[30]), .A6(n1670), .Y(n11201) );
  AOI22X1_HVT U721 ( .A1(n1525), .A2(n15000), .A3(n11000), .A4(n11201), .Y(
        n781) );
  OA22X1_HVT U722 ( .A1(n2770), .A2(n412), .A3(n10100), .A4(n3160), .Y(n7801)
         );
  NAND2X0_HVT U723 ( .A1(n1760), .A2(sram_rdata_6[30]), .Y(n779) );
  NAND3X0_HVT U724 ( .A1(n781), .A2(n7801), .A3(n779), .Y(n_src_aox[62]) );
  AO222X1_HVT U725 ( .A1(n1830), .A2(sram_rdata_5[31]), .A3(n2130), .A4(
        sram_rdata_4[31]), .A5(sram_rdata_3[31]), .A6(n2010), .Y(n15301) );
  AO222X1_HVT U726 ( .A1(n1910), .A2(sram_rdata_2[31]), .A3(n2130), .A4(
        sram_rdata_1[31]), .A5(sram_rdata_0[31]), .A6(n1990), .Y(n1124) );
  AOI22X1_HVT U727 ( .A1(n15301), .A2(n15000), .A3(n5801), .A4(n1124), .Y(n784) );
  OA22X1_HVT U728 ( .A1(n10300), .A2(n413), .A3(n2700), .A4(n3170), .Y(n783)
         );
  NAND2X0_HVT U729 ( .A1(n2270), .A2(sram_rdata_6[31]), .Y(n782) );
  NAND3X0_HVT U730 ( .A1(n784), .A2(n783), .A3(n782), .Y(n_src_aox[63]) );
  AO222X1_HVT U731 ( .A1(n2070), .A2(sram_rdata_4[16]), .A3(n2140), .A4(
        sram_rdata_3[16]), .A5(sram_rdata_5[16]), .A6(n1940), .Y(n1532) );
  AO222X1_HVT U732 ( .A1(n1830), .A2(sram_rdata_1[16]), .A3(n2120), .A4(
        sram_rdata_0[16]), .A5(sram_rdata_2[16]), .A6(n2020), .Y(n1128) );
  AOI22X1_HVT U733 ( .A1(n1532), .A2(n589), .A3(n11000), .A4(n1128), .Y(n787)
         );
  OA22X1_HVT U734 ( .A1(n10400), .A2(n494), .A3(n10100), .A4(n398), .Y(n786)
         );
  NAND2X0_HVT U735 ( .A1(n1820), .A2(sram_rdata_8[16]), .Y(n785) );
  NAND3X0_HVT U736 ( .A1(n787), .A2(n786), .A3(n785), .Y(n_src_aox[64]) );
  AO222X1_HVT U737 ( .A1(n1900), .A2(sram_rdata_4[17]), .A3(n2120), .A4(
        sram_rdata_3[17]), .A5(sram_rdata_5[17]), .A6(n16400), .Y(n1537) );
  AO222X1_HVT U738 ( .A1(n1900), .A2(sram_rdata_1[17]), .A3(n16000), .A4(
        sram_rdata_0[17]), .A5(sram_rdata_2[17]), .A6(n1700), .Y(n1132) );
  AOI22X1_HVT U739 ( .A1(n1537), .A2(n591), .A3(n579), .A4(n1132), .Y(n7901)
         );
  OA22X1_HVT U740 ( .A1(n10500), .A2(n495), .A3(n2730), .A4(n399), .Y(n789) );
  NAND2X0_HVT U741 ( .A1(n575), .A2(sram_rdata_8[17]), .Y(n788) );
  NAND3X0_HVT U742 ( .A1(n7901), .A2(n789), .A3(n788), .Y(n_src_aox[65]) );
  AO222X1_HVT U743 ( .A1(n2060), .A2(sram_rdata_4[18]), .A3(n2190), .A4(
        sram_rdata_3[18]), .A5(sram_rdata_5[18]), .A6(n16500), .Y(n1542) );
  AO222X1_HVT U744 ( .A1(n1850), .A2(sram_rdata_1[18]), .A3(n15900), .A4(
        sram_rdata_0[18]), .A5(sram_rdata_2[18]), .A6(n1690), .Y(n1136) );
  AOI22X1_HVT U745 ( .A1(n1542), .A2(n10800), .A3(n10900), .A4(n1136), .Y(n793) );
  OA22X1_HVT U746 ( .A1(n10300), .A2(n496), .A3(n14800), .A4(n4001), .Y(n792)
         );
  NAND2X0_HVT U747 ( .A1(n2210), .A2(sram_rdata_8[18]), .Y(n791) );
  NAND3X0_HVT U748 ( .A1(n793), .A2(n792), .A3(n791), .Y(n_src_aox[66]) );
  AO222X1_HVT U749 ( .A1(n2100), .A2(sram_rdata_4[19]), .A3(n587), .A4(
        sram_rdata_3[19]), .A5(sram_rdata_5[19]), .A6(n1710), .Y(n1544) );
  AO222X1_HVT U750 ( .A1(n1840), .A2(sram_rdata_1[19]), .A3(n13600), .A4(
        sram_rdata_0[19]), .A5(sram_rdata_2[19]), .A6(n1930), .Y(n11401) );
  AOI22X1_HVT U751 ( .A1(n1544), .A2(n591), .A3(n582), .A4(n11401), .Y(n796)
         );
  OA22X1_HVT U752 ( .A1(n2770), .A2(n497), .A3(n2690), .A4(n401), .Y(n795) );
  NAND2X0_HVT U753 ( .A1(n1810), .A2(sram_rdata_8[19]), .Y(n794) );
  NAND3X0_HVT U754 ( .A1(n796), .A2(n795), .A3(n794), .Y(n_src_aox[67]) );
  AO222X1_HVT U755 ( .A1(n1880), .A2(sram_rdata_4[20]), .A3(n16100), .A4(
        sram_rdata_3[20]), .A5(sram_rdata_5[20]), .A6(n2020), .Y(n1549) );
  AO222X1_HVT U756 ( .A1(n1880), .A2(sram_rdata_1[20]), .A3(n15800), .A4(
        sram_rdata_0[20]), .A5(sram_rdata_2[20]), .A6(n1970), .Y(n1144) );
  AOI22X1_HVT U757 ( .A1(n1549), .A2(n12800), .A3(n15100), .A4(n1144), .Y(n799) );
  OA22X1_HVT U758 ( .A1(n2800), .A2(n498), .A3(n11500), .A4(n402), .Y(n798) );
  NAND2X0_HVT U759 ( .A1(n1800), .A2(sram_rdata_8[20]), .Y(n797) );
  NAND3X0_HVT U760 ( .A1(n799), .A2(n798), .A3(n797), .Y(n_src_aox[68]) );
  AO222X1_HVT U761 ( .A1(n1830), .A2(sram_rdata_4[21]), .A3(n2130), .A4(
        sram_rdata_3[21]), .A5(sram_rdata_5[21]), .A6(n1990), .Y(n1554) );
  AO222X1_HVT U762 ( .A1(n1840), .A2(sram_rdata_1[21]), .A3(n2120), .A4(
        sram_rdata_0[21]), .A5(sram_rdata_2[21]), .A6(n1960), .Y(n1148) );
  AOI22X1_HVT U763 ( .A1(n1554), .A2(n10700), .A3(n578), .A4(n1148), .Y(n802)
         );
  OA22X1_HVT U764 ( .A1(n2790), .A2(n499), .A3(n10100), .A4(n403), .Y(n801) );
  NAND2X0_HVT U765 ( .A1(n1720), .A2(sram_rdata_8[21]), .Y(n8001) );
  NAND3X0_HVT U766 ( .A1(n802), .A2(n801), .A3(n8001), .Y(n_src_aox[69]) );
  AO222X1_HVT U767 ( .A1(n2070), .A2(sram_rdata_4[22]), .A3(n15600), .A4(
        sram_rdata_3[22]), .A5(sram_rdata_5[22]), .A6(n1930), .Y(n1559) );
  AO222X1_HVT U768 ( .A1(n2100), .A2(sram_rdata_1[22]), .A3(n2190), .A4(
        sram_rdata_0[22]), .A5(sram_rdata_2[22]), .A6(n16400), .Y(n1152) );
  AOI22X1_HVT U769 ( .A1(n1559), .A2(n589), .A3(n15200), .A4(n1152), .Y(n805)
         );
  OA22X1_HVT U770 ( .A1(n10600), .A2(n5001), .A3(n2740), .A4(n404), .Y(n804)
         );
  NAND2X0_HVT U771 ( .A1(n2260), .A2(sram_rdata_8[22]), .Y(n803) );
  NAND3X0_HVT U772 ( .A1(n805), .A2(n804), .A3(n803), .Y(n_src_aox[70]) );
  AO222X1_HVT U773 ( .A1(n2100), .A2(sram_rdata_4[23]), .A3(n16100), .A4(
        sram_rdata_3[23]), .A5(sram_rdata_5[23]), .A6(n1920), .Y(n1564) );
  AO222X1_HVT U774 ( .A1(n2100), .A2(sram_rdata_1[23]), .A3(n15800), .A4(
        sram_rdata_0[23]), .A5(sram_rdata_2[23]), .A6(n1930), .Y(n1156) );
  AOI22X1_HVT U775 ( .A1(n1564), .A2(n591), .A3(n582), .A4(n1156), .Y(n808) );
  OA22X1_HVT U776 ( .A1(n13700), .A2(n501), .A3(n2710), .A4(n405), .Y(n807) );
  NAND2X0_HVT U777 ( .A1(n2260), .A2(sram_rdata_8[23]), .Y(n806) );
  NAND3X0_HVT U778 ( .A1(n808), .A2(n807), .A3(n806), .Y(n_src_aox[71]) );
  AO222X1_HVT U779 ( .A1(n2050), .A2(sram_rdata_4[24]), .A3(n2190), .A4(
        sram_rdata_3[24]), .A5(sram_rdata_5[24]), .A6(n1670), .Y(n1569) );
  AO222X1_HVT U780 ( .A1(n1910), .A2(sram_rdata_1[24]), .A3(n2160), .A4(
        sram_rdata_0[24]), .A5(sram_rdata_2[24]), .A6(n16400), .Y(n11601) );
  AOI22X1_HVT U781 ( .A1(n1569), .A2(n10800), .A3(n12900), .A4(n11601), .Y(
        n811) );
  OA22X1_HVT U782 ( .A1(n13700), .A2(n502), .A3(n10000), .A4(n406), .Y(n8101)
         );
  NAND2X0_HVT U783 ( .A1(n574), .A2(sram_rdata_8[24]), .Y(n809) );
  NAND3X0_HVT U784 ( .A1(n811), .A2(n8101), .A3(n809), .Y(n_src_aox[72]) );
  AO222X1_HVT U785 ( .A1(n1659), .A2(sram_rdata_4[25]), .A3(n2170), .A4(
        sram_rdata_3[25]), .A5(sram_rdata_5[25]), .A6(n16600), .Y(n1571) );
  AO222X1_HVT U786 ( .A1(n2060), .A2(sram_rdata_1[25]), .A3(n16100), .A4(
        sram_rdata_0[25]), .A5(sram_rdata_2[25]), .A6(n16400), .Y(n1164) );
  AOI22X1_HVT U787 ( .A1(n1571), .A2(n14900), .A3(n15200), .A4(n1164), .Y(n814) );
  OA22X1_HVT U788 ( .A1(n2810), .A2(n503), .A3(n1661), .A4(n407), .Y(n813) );
  NAND2X0_HVT U789 ( .A1(n2240), .A2(sram_rdata_8[25]), .Y(n812) );
  NAND3X0_HVT U790 ( .A1(n814), .A2(n813), .A3(n812), .Y(n_src_aox[73]) );
  AO222X1_HVT U791 ( .A1(n2060), .A2(sram_rdata_4[26]), .A3(n15700), .A4(
        sram_rdata_3[26]), .A5(sram_rdata_5[26]), .A6(n1920), .Y(n1573) );
  AO222X1_HVT U792 ( .A1(n2050), .A2(sram_rdata_1[26]), .A3(n587), .A4(
        sram_rdata_0[26]), .A5(sram_rdata_2[26]), .A6(n1700), .Y(n1165) );
  AOI22X1_HVT U793 ( .A1(n1573), .A2(n14900), .A3(n579), .A4(n1165), .Y(n817)
         );
  OA22X1_HVT U794 ( .A1(n2760), .A2(n504), .A3(n10100), .A4(n408), .Y(n816) );
  NAND2X0_HVT U795 ( .A1(n1760), .A2(sram_rdata_8[26]), .Y(n815) );
  NAND3X0_HVT U796 ( .A1(n817), .A2(n816), .A3(n815), .Y(n_src_aox[74]) );
  AO222X1_HVT U797 ( .A1(n1860), .A2(sram_rdata_4[27]), .A3(n2110), .A4(
        sram_rdata_3[27]), .A5(sram_rdata_5[27]), .A6(n2000), .Y(n1575) );
  AO222X1_HVT U798 ( .A1(n1890), .A2(sram_rdata_1[27]), .A3(n15600), .A4(
        sram_rdata_0[27]), .A5(sram_rdata_2[27]), .A6(n1980), .Y(n1169) );
  AOI22X1_HVT U799 ( .A1(n1575), .A2(n588), .A3(n15100), .A4(n1169), .Y(n8201)
         );
  OA22X1_HVT U800 ( .A1(n10600), .A2(n505), .A3(n14600), .A4(n409), .Y(n819)
         );
  NAND2X0_HVT U801 ( .A1(n574), .A2(sram_rdata_8[27]), .Y(n818) );
  NAND3X0_HVT U802 ( .A1(n8201), .A2(n819), .A3(n818), .Y(n_src_aox[75]) );
  AO222X1_HVT U803 ( .A1(n2100), .A2(sram_rdata_4[28]), .A3(n15500), .A4(
        sram_rdata_3[28]), .A5(sram_rdata_5[28]), .A6(n1980), .Y(n15801) );
  AO222X1_HVT U804 ( .A1(n2050), .A2(sram_rdata_1[28]), .A3(n16000), .A4(
        sram_rdata_0[28]), .A5(sram_rdata_2[28]), .A6(n2000), .Y(n1173) );
  AOI22X1_HVT U805 ( .A1(n15801), .A2(n12800), .A3(n579), .A4(n1173), .Y(n823)
         );
  OA22X1_HVT U806 ( .A1(n11900), .A2(n506), .A3(n2710), .A4(n4101), .Y(n822)
         );
  NAND2X0_HVT U807 ( .A1(n1810), .A2(sram_rdata_8[28]), .Y(n821) );
  NAND3X0_HVT U808 ( .A1(n823), .A2(n822), .A3(n821), .Y(n_src_aox[76]) );
  AO222X1_HVT U809 ( .A1(n1840), .A2(sram_rdata_4[29]), .A3(n13500), .A4(
        sram_rdata_3[29]), .A5(sram_rdata_5[29]), .A6(n2020), .Y(n1585) );
  AO222X1_HVT U810 ( .A1(n2060), .A2(sram_rdata_1[29]), .A3(n15900), .A4(
        sram_rdata_0[29]), .A5(sram_rdata_2[29]), .A6(n1990), .Y(n1177) );
  AOI22X1_HVT U811 ( .A1(n1585), .A2(n12800), .A3(n1648), .A4(n1177), .Y(n826)
         );
  OA22X1_HVT U812 ( .A1(n12000), .A2(n507), .A3(n14800), .A4(n411), .Y(n825)
         );
  NAND2X0_HVT U813 ( .A1(n1730), .A2(sram_rdata_8[29]), .Y(n824) );
  NAND3X0_HVT U814 ( .A1(n826), .A2(n825), .A3(n824), .Y(n_src_aox[77]) );
  AO222X1_HVT U815 ( .A1(n2050), .A2(sram_rdata_4[30]), .A3(n2180), .A4(
        sram_rdata_3[30]), .A5(sram_rdata_5[30]), .A6(n1690), .Y(n15901) );
  AO222X1_HVT U816 ( .A1(n12500), .A2(sram_rdata_1[30]), .A3(n15400), .A4(
        sram_rdata_0[30]), .A5(sram_rdata_2[30]), .A6(n1710), .Y(n1181) );
  AOI22X1_HVT U817 ( .A1(n15901), .A2(n12700), .A3(n10900), .A4(n1181), .Y(
        n829) );
  OA22X1_HVT U818 ( .A1(n13800), .A2(n508), .A3(n2750), .A4(n412), .Y(n828) );
  NAND2X0_HVT U819 ( .A1(n2250), .A2(sram_rdata_8[30]), .Y(n827) );
  NAND3X0_HVT U820 ( .A1(n829), .A2(n828), .A3(n827), .Y(n_src_aox[78]) );
  AO222X1_HVT U821 ( .A1(n1830), .A2(sram_rdata_4[31]), .A3(n587), .A4(
        sram_rdata_3[31]), .A5(sram_rdata_5[31]), .A6(n1710), .Y(n1592) );
  AO222X1_HVT U822 ( .A1(n2040), .A2(sram_rdata_1[31]), .A3(n2110), .A4(
        sram_rdata_0[31]), .A5(sram_rdata_2[31]), .A6(n1970), .Y(n1182) );
  AOI22X1_HVT U823 ( .A1(n1592), .A2(n589), .A3(n581), .A4(n1182), .Y(n832) );
  OA22X1_HVT U824 ( .A1(n12100), .A2(n509), .A3(n11500), .A4(n413), .Y(n831)
         );
  NAND2X0_HVT U825 ( .A1(n1760), .A2(sram_rdata_8[31]), .Y(n8301) );
  NAND3X0_HVT U826 ( .A1(n832), .A2(n831), .A3(n8301), .Y(n_src_aox[79]) );
  AO222X1_HVT U827 ( .A1(n12500), .A2(sram_rdata_3[16]), .A3(n16000), .A4(
        sram_rdata_5[16]), .A5(n1700), .A6(sram_rdata_4[16]), .Y(n1597) );
  AO222X1_HVT U828 ( .A1(n2060), .A2(sram_rdata_0[16]), .A3(n13600), .A4(
        sram_rdata_2[16]), .A5(n2010), .A6(sram_rdata_1[16]), .Y(n1186) );
  AOI22X1_HVT U829 ( .A1(n1597), .A2(n591), .A3(n11000), .A4(n1186), .Y(n835)
         );
  OA22X1_HVT U830 ( .A1(n10400), .A2(n3020), .A3(n2710), .A4(n494), .Y(n834)
         );
  NAND2X0_HVT U831 ( .A1(n2240), .A2(sram_rdata_7[16]), .Y(n833) );
  NAND3X0_HVT U832 ( .A1(n835), .A2(n834), .A3(n833), .Y(n_src_aox[80]) );
  AO222X1_HVT U833 ( .A1(n1850), .A2(sram_rdata_3[17]), .A3(n2110), .A4(
        sram_rdata_5[17]), .A5(n1990), .A6(sram_rdata_4[17]), .Y(n1602) );
  AO222X1_HVT U834 ( .A1(n1840), .A2(sram_rdata_0[17]), .A3(n2140), .A4(
        sram_rdata_2[17]), .A5(n1920), .A6(sram_rdata_1[17]), .Y(n11901) );
  AOI22X1_HVT U835 ( .A1(n1602), .A2(n589), .A3(n5801), .A4(n11901), .Y(n838)
         );
  OA22X1_HVT U836 ( .A1(n11900), .A2(n3030), .A3(n2740), .A4(n495), .Y(n837)
         );
  NAND2X0_HVT U837 ( .A1(n2270), .A2(sram_rdata_7[17]), .Y(n836) );
  NAND3X0_HVT U838 ( .A1(n838), .A2(n837), .A3(n836), .Y(n_src_aox[81]) );
  AO222X1_HVT U839 ( .A1(n2090), .A2(sram_rdata_3[18]), .A3(n2130), .A4(
        sram_rdata_5[18]), .A5(n2020), .A6(sram_rdata_4[18]), .Y(n1607) );
  AO222X1_HVT U840 ( .A1(n1900), .A2(sram_rdata_0[18]), .A3(n13600), .A4(
        sram_rdata_2[18]), .A5(n2010), .A6(sram_rdata_1[18]), .Y(n1194) );
  AOI22X1_HVT U841 ( .A1(n1607), .A2(n591), .A3(n12900), .A4(n1194), .Y(n841)
         );
  OA22X1_HVT U842 ( .A1(n10300), .A2(n3040), .A3(n2720), .A4(n496), .Y(n8401)
         );
  NAND2X0_HVT U843 ( .A1(n1740), .A2(sram_rdata_7[18]), .Y(n839) );
  NAND3X0_HVT U844 ( .A1(n841), .A2(n8401), .A3(n839), .Y(n_src_aox[82]) );
  AO222X1_HVT U845 ( .A1(n1900), .A2(sram_rdata_3[19]), .A3(n15400), .A4(
        sram_rdata_5[19]), .A5(n1980), .A6(sram_rdata_4[19]), .Y(n1609) );
  AO222X1_HVT U846 ( .A1(n1840), .A2(sram_rdata_0[19]), .A3(n16100), .A4(
        sram_rdata_2[19]), .A5(n16600), .A6(sram_rdata_1[19]), .Y(n1198) );
  AOI22X1_HVT U847 ( .A1(n1609), .A2(n14900), .A3(n5801), .A4(n1198), .Y(n844)
         );
  OA22X1_HVT U848 ( .A1(n2770), .A2(n3050), .A3(n14500), .A4(n497), .Y(n843)
         );
  NAND2X0_HVT U849 ( .A1(n2230), .A2(sram_rdata_7[19]), .Y(n842) );
  NAND3X0_HVT U850 ( .A1(n844), .A2(n843), .A3(n842), .Y(n_src_aox[83]) );
  AO222X1_HVT U851 ( .A1(n2030), .A2(sram_rdata_3[20]), .A3(n2170), .A4(
        sram_rdata_5[20]), .A5(n1680), .A6(sram_rdata_4[20]), .Y(n1611) );
  AO222X1_HVT U852 ( .A1(n1890), .A2(sram_rdata_0[20]), .A3(n2130), .A4(
        sram_rdata_2[20]), .A5(n1690), .A6(sram_rdata_1[20]), .Y(n1202) );
  AOI22X1_HVT U853 ( .A1(n1611), .A2(n12700), .A3(n15100), .A4(n1202), .Y(n847) );
  OA22X1_HVT U854 ( .A1(n2810), .A2(n3060), .A3(n14600), .A4(n498), .Y(n846)
         );
  NAND2X0_HVT U855 ( .A1(n574), .A2(sram_rdata_7[20]), .Y(n845) );
  NAND3X0_HVT U856 ( .A1(n847), .A2(n846), .A3(n845), .Y(n_src_aox[84]) );
  AO222X1_HVT U857 ( .A1(n1890), .A2(sram_rdata_3[21]), .A3(n15900), .A4(
        sram_rdata_5[21]), .A5(n1990), .A6(sram_rdata_4[21]), .Y(n1613) );
  AO222X1_HVT U858 ( .A1(n12500), .A2(sram_rdata_0[21]), .A3(n15500), .A4(
        sram_rdata_2[21]), .A5(n1920), .A6(sram_rdata_1[21]), .Y(n1206) );
  AOI22X1_HVT U859 ( .A1(n1613), .A2(n588), .A3(n579), .A4(n1206), .Y(n8501)
         );
  OA22X1_HVT U860 ( .A1(n2790), .A2(n3070), .A3(n2730), .A4(n499), .Y(n849) );
  NAND2X0_HVT U861 ( .A1(n2280), .A2(sram_rdata_7[21]), .Y(n848) );
  NAND3X0_HVT U862 ( .A1(n8501), .A2(n849), .A3(n848), .Y(n_src_aox[85]) );
  AO222X1_HVT U863 ( .A1(n1910), .A2(sram_rdata_3[22]), .A3(n587), .A4(
        sram_rdata_5[22]), .A5(n1690), .A6(sram_rdata_4[22]), .Y(n1618) );
  AO222X1_HVT U864 ( .A1(n2030), .A2(sram_rdata_0[22]), .A3(n2180), .A4(
        sram_rdata_2[22]), .A5(n2010), .A6(sram_rdata_1[22]), .Y(n12101) );
  AOI22X1_HVT U865 ( .A1(n1618), .A2(n591), .A3(n579), .A4(n12101), .Y(n853)
         );
  OA22X1_HVT U866 ( .A1(n11800), .A2(n3080), .A3(n14700), .A4(n5001), .Y(n852)
         );
  NAND2X0_HVT U867 ( .A1(n1770), .A2(sram_rdata_7[22]), .Y(n851) );
  NAND3X0_HVT U868 ( .A1(n853), .A2(n852), .A3(n851), .Y(n_src_aox[86]) );
  AO222X1_HVT U869 ( .A1(n13900), .A2(sram_rdata_3[23]), .A3(n2120), .A4(
        sram_rdata_5[23]), .A5(n1970), .A6(sram_rdata_4[23]), .Y(n1623) );
  AO222X1_HVT U870 ( .A1(n12500), .A2(sram_rdata_0[23]), .A3(n15800), .A4(
        sram_rdata_2[23]), .A5(n1940), .A6(sram_rdata_1[23]), .Y(n1214) );
  AOI22X1_HVT U871 ( .A1(n1623), .A2(n591), .A3(n582), .A4(n1214), .Y(n856) );
  OA22X1_HVT U872 ( .A1(n2760), .A2(n3090), .A3(n2690), .A4(n501), .Y(n855) );
  NAND2X0_HVT U873 ( .A1(n2230), .A2(sram_rdata_7[23]), .Y(n854) );
  NAND3X0_HVT U874 ( .A1(n856), .A2(n855), .A3(n854), .Y(n_src_aox[87]) );
  AO222X1_HVT U875 ( .A1(n2090), .A2(sram_rdata_3[24]), .A3(n587), .A4(
        sram_rdata_5[24]), .A5(n1940), .A6(sram_rdata_4[24]), .Y(n1625) );
  AO222X1_HVT U876 ( .A1(n2090), .A2(sram_rdata_0[24]), .A3(n2180), .A4(
        sram_rdata_2[24]), .A5(n16600), .A6(sram_rdata_1[24]), .Y(n1218) );
  AOI22X1_HVT U877 ( .A1(n1625), .A2(n589), .A3(n5801), .A4(n1218), .Y(n859)
         );
  OA22X1_HVT U878 ( .A1(n2790), .A2(n3100), .A3(n2690), .A4(n502), .Y(n858) );
  NAND2X0_HVT U879 ( .A1(n2230), .A2(sram_rdata_7[24]), .Y(n857) );
  NAND3X0_HVT U880 ( .A1(n859), .A2(n858), .A3(n857), .Y(n_src_aox[88]) );
  AO222X1_HVT U881 ( .A1(n2090), .A2(sram_rdata_3[25]), .A3(n2140), .A4(
        sram_rdata_5[25]), .A5(n1700), .A6(sram_rdata_4[25]), .Y(n1627) );
  AO222X1_HVT U882 ( .A1(n2070), .A2(sram_rdata_0[25]), .A3(n13500), .A4(
        sram_rdata_2[25]), .A5(n1680), .A6(sram_rdata_1[25]), .Y(n1222) );
  AOI22X1_HVT U883 ( .A1(n1627), .A2(n14900), .A3(n579), .A4(n1222), .Y(n862)
         );
  OA22X1_HVT U884 ( .A1(n2800), .A2(n3110), .A3(n14700), .A4(n503), .Y(n861)
         );
  NAND2X0_HVT U885 ( .A1(n1790), .A2(sram_rdata_7[25]), .Y(n8601) );
  NAND3X0_HVT U886 ( .A1(n862), .A2(n861), .A3(n8601), .Y(n_src_aox[89]) );
  AO222X1_HVT U887 ( .A1(n2050), .A2(sram_rdata_3[26]), .A3(n2160), .A4(
        sram_rdata_5[26]), .A5(n16601), .A6(sram_rdata_4[26]), .Y(n1629) );
  AO222X1_HVT U888 ( .A1(n1659), .A2(sram_rdata_0[26]), .A3(n2190), .A4(
        sram_rdata_2[26]), .A5(n16601), .A6(sram_rdata_1[26]), .Y(n1226) );
  AOI22X1_HVT U889 ( .A1(n1629), .A2(n12700), .A3(n12900), .A4(n1226), .Y(n865) );
  OA22X1_HVT U890 ( .A1(n2760), .A2(n3120), .A3(n14700), .A4(n504), .Y(n864)
         );
  NAND2X0_HVT U891 ( .A1(n1720), .A2(sram_rdata_7[26]), .Y(n863) );
  NAND3X0_HVT U892 ( .A1(n865), .A2(n864), .A3(n863), .Y(n_src_aox[90]) );
  AO222X1_HVT U893 ( .A1(n1900), .A2(sram_rdata_3[27]), .A3(n2170), .A4(
        sram_rdata_5[27]), .A5(n16500), .A6(sram_rdata_4[27]), .Y(n1631) );
  AO222X1_HVT U894 ( .A1(n2060), .A2(sram_rdata_0[27]), .A3(n15800), .A4(
        sram_rdata_2[27]), .A5(n2020), .A6(sram_rdata_1[27]), .Y(n1227) );
  AOI22X1_HVT U895 ( .A1(n1631), .A2(n12800), .A3(n10900), .A4(n1227), .Y(n868) );
  OA22X1_HVT U896 ( .A1(n11800), .A2(n3130), .A3(n14600), .A4(n505), .Y(n867)
         );
  NAND2X0_HVT U897 ( .A1(n1750), .A2(sram_rdata_7[27]), .Y(n866) );
  NAND3X0_HVT U898 ( .A1(n868), .A2(n867), .A3(n866), .Y(n_src_aox[91]) );
  AO222X1_HVT U899 ( .A1(n2040), .A2(sram_rdata_3[28]), .A3(n13500), .A4(
        sram_rdata_5[28]), .A5(n1970), .A6(sram_rdata_4[28]), .Y(n1633) );
  AO222X1_HVT U900 ( .A1(n2030), .A2(sram_rdata_0[28]), .A3(n15600), .A4(
        sram_rdata_2[28]), .A5(n1990), .A6(sram_rdata_1[28]), .Y(n1231) );
  AOI22X1_HVT U901 ( .A1(n1633), .A2(n14900), .A3(n5801), .A4(n1231), .Y(n871)
         );
  OA22X1_HVT U902 ( .A1(n11900), .A2(n3140), .A3(n10000), .A4(n506), .Y(n8701)
         );
  NAND2X0_HVT U903 ( .A1(n2250), .A2(sram_rdata_7[28]), .Y(n869) );
  NAND3X0_HVT U904 ( .A1(n871), .A2(n8701), .A3(n869), .Y(n_src_aox[92]) );
  AO222X1_HVT U905 ( .A1(n1890), .A2(sram_rdata_3[29]), .A3(n2120), .A4(
        sram_rdata_5[29]), .A5(n1960), .A6(sram_rdata_4[29]), .Y(n1638) );
  AO222X1_HVT U906 ( .A1(n1890), .A2(sram_rdata_0[29]), .A3(n587), .A4(
        sram_rdata_2[29]), .A5(n1920), .A6(sram_rdata_1[29]), .Y(n1235) );
  AOI22X1_HVT U907 ( .A1(n1638), .A2(n588), .A3(n15100), .A4(n1235), .Y(n874)
         );
  OA22X1_HVT U908 ( .A1(n12000), .A2(n3150), .A3(n2750), .A4(n507), .Y(n873)
         );
  NAND2X0_HVT U909 ( .A1(n1720), .A2(sram_rdata_7[29]), .Y(n872) );
  NAND3X0_HVT U910 ( .A1(n874), .A2(n873), .A3(n872), .Y(n_src_aox[93]) );
  AO222X1_HVT U911 ( .A1(n2080), .A2(sram_rdata_3[30]), .A3(n15800), .A4(
        sram_rdata_5[30]), .A5(n1710), .A6(sram_rdata_4[30]), .Y(n1643) );
  AO222X1_HVT U912 ( .A1(n1860), .A2(sram_rdata_0[30]), .A3(n15800), .A4(
        sram_rdata_2[30]), .A5(n2010), .A6(sram_rdata_1[30]), .Y(n1236) );
  AO222X1_HVT U913 ( .A1(n1900), .A2(sram_rdata_3[31]), .A3(n15600), .A4(
        sram_rdata_5[31]), .A5(n1670), .A6(sram_rdata_4[31]), .Y(n1649) );
  AO222X1_HVT U914 ( .A1(n1830), .A2(sram_rdata_0[31]), .A3(n13500), .A4(
        sram_rdata_2[31]), .A5(n1700), .A6(sram_rdata_1[31]), .Y(n12401) );
  AOI22X1_HVT U915 ( .A1(n1649), .A2(n589), .A3(n578), .A4(n12401), .Y(n877)
         );
  OA22X1_HVT U916 ( .A1(n10300), .A2(n3170), .A3(n2710), .A4(n509), .Y(n876)
         );
  NAND2X0_HVT U917 ( .A1(n1730), .A2(sram_rdata_7[31]), .Y(n875) );
  NAND3X0_HVT U918 ( .A1(n877), .A2(n876), .A3(n875), .Y(n_src_aox[95]) );
  AO222X1_HVT U919 ( .A1(sram_rdata_6[0]), .A2(n2000), .A3(sram_rdata_8[0]), 
        .A4(n2100), .A5(sram_rdata_7[0]), .A6(n2190), .Y(n1245) );
  AOI22X1_HVT U920 ( .A1(n1245), .A2(n10900), .A3(n12700), .A4(n878), .Y(n881)
         );
  OA22X1_HVT U921 ( .A1(n10400), .A2(n3180), .A3(n14500), .A4(n478), .Y(n8801)
         );
  NAND2X0_HVT U922 ( .A1(n1760), .A2(sram_rdata_3[0]), .Y(n879) );
  NAND3X0_HVT U923 ( .A1(n881), .A2(n8801), .A3(n879), .Y(n_src_aox[96]) );
  AO222X1_HVT U924 ( .A1(n2060), .A2(sram_rdata_8[1]), .A3(n2160), .A4(
        sram_rdata_7[1]), .A5(sram_rdata_6[1]), .A6(n2010), .Y(n1249) );
  AOI22X1_HVT U925 ( .A1(n882), .A2(n10800), .A3(n15100), .A4(n1249), .Y(n885)
         );
  OA22X1_HVT U926 ( .A1(n11900), .A2(n3190), .A3(n2730), .A4(n5101), .Y(n884)
         );
  NAND2X0_HVT U927 ( .A1(n1820), .A2(sram_rdata_3[1]), .Y(n883) );
  NAND3X0_HVT U928 ( .A1(n885), .A2(n884), .A3(n883), .Y(n_src_aox[97]) );
  AO222X1_HVT U929 ( .A1(n1900), .A2(sram_rdata_8[2]), .A3(n15800), .A4(
        sram_rdata_7[2]), .A5(sram_rdata_6[2]), .A6(n16500), .Y(n1254) );
  AOI22X1_HVT U930 ( .A1(n886), .A2(n588), .A3(n1648), .A4(n1254), .Y(n889) );
  OA22X1_HVT U931 ( .A1(n12100), .A2(n3200), .A3(n1661), .A4(n511), .Y(n888)
         );
  NAND2X0_HVT U932 ( .A1(n1800), .A2(sram_rdata_3[2]), .Y(n887) );
  NAND3X0_HVT U933 ( .A1(n889), .A2(n888), .A3(n887), .Y(n_src_aox[98]) );
  AO222X1_HVT U934 ( .A1(n2090), .A2(sram_rdata_8[3]), .A3(n2110), .A4(
        sram_rdata_7[3]), .A5(sram_rdata_6[3]), .A6(n2000), .Y(n1259) );
  AOI22X1_HVT U935 ( .A1(n8901), .A2(n589), .A3(n11000), .A4(n1259), .Y(n893)
         );
  OA22X1_HVT U936 ( .A1(n2780), .A2(n3210), .A3(n2690), .A4(n512), .Y(n892) );
  NAND2X0_HVT U937 ( .A1(n2270), .A2(sram_rdata_3[3]), .Y(n891) );
  NAND3X0_HVT U938 ( .A1(n893), .A2(n892), .A3(n891), .Y(n_src_aox[99]) );
  AO222X1_HVT U939 ( .A1(n12500), .A2(sram_rdata_8[4]), .A3(n2130), .A4(
        sram_rdata_7[4]), .A5(sram_rdata_6[4]), .A6(n1960), .Y(n1264) );
  AOI22X1_HVT U940 ( .A1(n894), .A2(n10700), .A3(n579), .A4(n1264), .Y(n897)
         );
  OA22X1_HVT U941 ( .A1(n2800), .A2(n3220), .A3(n14600), .A4(n513), .Y(n896)
         );
  NAND2X0_HVT U942 ( .A1(n1790), .A2(sram_rdata_3[4]), .Y(n895) );
  NAND3X0_HVT U943 ( .A1(n897), .A2(n896), .A3(n895), .Y(n_src_aox[100]) );
  AO222X1_HVT U944 ( .A1(n1910), .A2(sram_rdata_8[5]), .A3(n15800), .A4(
        sram_rdata_7[5]), .A5(sram_rdata_6[5]), .A6(n1960), .Y(n1269) );
  AOI22X1_HVT U945 ( .A1(n898), .A2(n15000), .A3(n12900), .A4(n1269), .Y(n901)
         );
  OA22X1_HVT U946 ( .A1(n2790), .A2(n3230), .A3(n14800), .A4(n514), .Y(n9001)
         );
  NAND2X0_HVT U947 ( .A1(n574), .A2(sram_rdata_3[5]), .Y(n899) );
  NAND3X0_HVT U948 ( .A1(n901), .A2(n9001), .A3(n899), .Y(n_src_aox[101]) );
  AO222X1_HVT U949 ( .A1(n1910), .A2(sram_rdata_8[6]), .A3(n15800), .A4(
        sram_rdata_7[6]), .A5(sram_rdata_6[6]), .A6(n2010), .Y(n1271) );
  AOI22X1_HVT U950 ( .A1(n902), .A2(n15000), .A3(n5801), .A4(n1271), .Y(n905)
         );
  OA22X1_HVT U951 ( .A1(n11800), .A2(n3240), .A3(n2730), .A4(n515), .Y(n904)
         );
  NAND2X0_HVT U952 ( .A1(n2210), .A2(sram_rdata_3[6]), .Y(n903) );
  NAND3X0_HVT U953 ( .A1(n905), .A2(n904), .A3(n903), .Y(n_src_aox[102]) );
  AO222X1_HVT U954 ( .A1(n2070), .A2(sram_rdata_8[7]), .A3(n2120), .A4(
        sram_rdata_7[7]), .A5(sram_rdata_6[7]), .A6(n1710), .Y(n1276) );
  AOI22X1_HVT U955 ( .A1(n906), .A2(n12700), .A3(n12600), .A4(n1276), .Y(n909)
         );
  OA22X1_HVT U956 ( .A1(n13700), .A2(n3250), .A3(n10000), .A4(n516), .Y(n908)
         );
  NAND2X0_HVT U957 ( .A1(n1800), .A2(sram_rdata_3[7]), .Y(n907) );
  NAND3X0_HVT U958 ( .A1(n909), .A2(n908), .A3(n907), .Y(n_src_aox[103]) );
  AO222X1_HVT U959 ( .A1(n2050), .A2(sram_rdata_8[8]), .A3(n2110), .A4(
        sram_rdata_7[8]), .A5(sram_rdata_6[8]), .A6(n16600), .Y(n1281) );
  AOI22X1_HVT U960 ( .A1(n9101), .A2(n15000), .A3(n12600), .A4(n1281), .Y(n913) );
  OA22X1_HVT U961 ( .A1(n13700), .A2(n3260), .A3(n14500), .A4(n517), .Y(n912)
         );
  NAND2X0_HVT U962 ( .A1(n1740), .A2(sram_rdata_3[8]), .Y(n911) );
  NAND3X0_HVT U963 ( .A1(n913), .A2(n912), .A3(n911), .Y(n_src_aox[104]) );
  AO222X1_HVT U964 ( .A1(n2090), .A2(sram_rdata_8[9]), .A3(n2140), .A4(
        sram_rdata_7[9]), .A5(sram_rdata_6[9]), .A6(n1700), .Y(n1286) );
  AOI22X1_HVT U965 ( .A1(n914), .A2(n591), .A3(n15200), .A4(n1286), .Y(n917)
         );
  OA22X1_HVT U966 ( .A1(n2810), .A2(n327), .A3(n14700), .A4(n518), .Y(n916) );
  NAND2X0_HVT U967 ( .A1(n576), .A2(sram_rdata_3[9]), .Y(n915) );
  NAND3X0_HVT U968 ( .A1(n917), .A2(n916), .A3(n915), .Y(n_src_aox[105]) );
  AO222X1_HVT U969 ( .A1(n1880), .A2(sram_rdata_8[10]), .A3(n13500), .A4(
        sram_rdata_7[10]), .A5(sram_rdata_6[10]), .A6(n16600), .Y(n1291) );
  AOI22X1_HVT U970 ( .A1(n918), .A2(n14900), .A3(n581), .A4(n1291), .Y(n921)
         );
  OA22X1_HVT U971 ( .A1(n13700), .A2(n328), .A3(n2740), .A4(n519), .Y(n9201)
         );
  NAND2X0_HVT U972 ( .A1(n2260), .A2(sram_rdata_3[10]), .Y(n919) );
  NAND3X0_HVT U973 ( .A1(n921), .A2(n9201), .A3(n919), .Y(n_src_aox[106]) );
  AO222X1_HVT U974 ( .A1(n1840), .A2(sram_rdata_8[11]), .A3(n16100), .A4(
        sram_rdata_7[11]), .A5(sram_rdata_6[11]), .A6(n16600), .Y(n1296) );
  AOI22X1_HVT U975 ( .A1(n922), .A2(n591), .A3(n10900), .A4(n1296), .Y(n925)
         );
  OA22X1_HVT U976 ( .A1(n10600), .A2(n329), .A3(n2690), .A4(n5201), .Y(n924)
         );
  NAND2X0_HVT U977 ( .A1(n2280), .A2(sram_rdata_3[11]), .Y(n923) );
  NAND3X0_HVT U978 ( .A1(n925), .A2(n924), .A3(n923), .Y(n_src_aox[107]) );
  AO222X1_HVT U979 ( .A1(n1900), .A2(sram_rdata_8[12]), .A3(n13500), .A4(
        sram_rdata_7[12]), .A5(sram_rdata_6[12]), .A6(n16600), .Y(n1298) );
  AOI22X1_HVT U980 ( .A1(n926), .A2(n589), .A3(n12600), .A4(n1298), .Y(n929)
         );
  OA22X1_HVT U981 ( .A1(n10500), .A2(n330), .A3(n10000), .A4(n521), .Y(n928)
         );
  NAND2X0_HVT U982 ( .A1(n575), .A2(sram_rdata_3[12]), .Y(n927) );
  NAND3X0_HVT U983 ( .A1(n929), .A2(n928), .A3(n927), .Y(n_src_aox[108]) );
  AO222X1_HVT U984 ( .A1(n2050), .A2(sram_rdata_8[13]), .A3(n2190), .A4(
        sram_rdata_7[13]), .A5(sram_rdata_6[13]), .A6(n2020), .Y(n13001) );
  AOI22X1_HVT U985 ( .A1(n9301), .A2(n10800), .A3(n11000), .A4(n13001), .Y(
        n933) );
  OA22X1_HVT U986 ( .A1(n12000), .A2(n331), .A3(n2720), .A4(n522), .Y(n932) );
  NAND2X0_HVT U987 ( .A1(n2240), .A2(sram_rdata_3[13]), .Y(n931) );
  NAND3X0_HVT U988 ( .A1(n933), .A2(n932), .A3(n931), .Y(n_src_aox[109]) );
  AO222X1_HVT U989 ( .A1(n1860), .A2(sram_rdata_8[14]), .A3(n16000), .A4(
        sram_rdata_7[14]), .A5(sram_rdata_6[14]), .A6(n1990), .Y(n1305) );
  AOI22X1_HVT U990 ( .A1(n934), .A2(n591), .A3(n15100), .A4(n1305), .Y(n937)
         );
  OA22X1_HVT U991 ( .A1(n2770), .A2(n332), .A3(n14800), .A4(n523), .Y(n936) );
  NAND2X0_HVT U992 ( .A1(n1800), .A2(sram_rdata_3[14]), .Y(n935) );
  NAND3X0_HVT U993 ( .A1(n937), .A2(n936), .A3(n935), .Y(n_src_aox[110]) );
  AO222X1_HVT U994 ( .A1(n1890), .A2(sram_rdata_8[15]), .A3(n15600), .A4(
        sram_rdata_7[15]), .A5(sram_rdata_6[15]), .A6(n1970), .Y(n13101) );
  AOI22X1_HVT U995 ( .A1(n938), .A2(n14900), .A3(n15100), .A4(n13101), .Y(n941) );
  OA22X1_HVT U996 ( .A1(n10300), .A2(n333), .A3(n2710), .A4(n524), .Y(n9401)
         );
  NAND2X0_HVT U997 ( .A1(n1730), .A2(sram_rdata_3[15]), .Y(n939) );
  NAND3X0_HVT U998 ( .A1(n941), .A2(n9401), .A3(n939), .Y(n_src_aox[111]) );
  AO222X1_HVT U999 ( .A1(sram_rdata_6[0]), .A2(n2170), .A3(sram_rdata_8[0]), 
        .A4(n1920), .A5(n2070), .A6(sram_rdata_7[0]), .Y(n1316) );
  AOI22X1_HVT U1000 ( .A1(n1316), .A2(n578), .A3(n592), .A4(n942), .Y(n945) );
  OA22X1_HVT U1001 ( .A1(n10400), .A2(n382), .A3(n11500), .A4(n3180), .Y(n944)
         );
  NAND2X0_HVT U1002 ( .A1(n1820), .A2(sram_rdata_5[0]), .Y(n943) );
  NAND3X0_HVT U1003 ( .A1(n945), .A2(n944), .A3(n943), .Y(n_src_aox[112]) );
  AO222X1_HVT U1004 ( .A1(n12500), .A2(sram_rdata_7[1]), .A3(n16000), .A4(
        sram_rdata_6[1]), .A5(n1690), .A6(sram_rdata_8[1]), .Y(n1317) );
  AOI22X1_HVT U1005 ( .A1(n946), .A2(n588), .A3(n5801), .A4(n1317), .Y(n949)
         );
  OA22X1_HVT U1006 ( .A1(n10500), .A2(n414), .A3(n10100), .A4(n3190), .Y(n948)
         );
  NAND2X0_HVT U1007 ( .A1(n1720), .A2(sram_rdata_5[1]), .Y(n947) );
  NAND3X0_HVT U1008 ( .A1(n949), .A2(n948), .A3(n947), .Y(n_src_aox[113]) );
  AO222X1_HVT U1009 ( .A1(n2090), .A2(sram_rdata_7[2]), .A3(n15500), .A4(
        sram_rdata_6[2]), .A5(n1680), .A6(sram_rdata_8[2]), .Y(n1322) );
  AOI22X1_HVT U1010 ( .A1(n9501), .A2(n14900), .A3(n5801), .A4(n1322), .Y(n953) );
  OA22X1_HVT U1011 ( .A1(n12100), .A2(n415), .A3(n14700), .A4(n3200), .Y(n952)
         );
  NAND2X0_HVT U1012 ( .A1(n2250), .A2(sram_rdata_5[2]), .Y(n951) );
  NAND3X0_HVT U1013 ( .A1(n953), .A2(n952), .A3(n951), .Y(n_src_aox[114]) );
  AO222X1_HVT U1014 ( .A1(n1880), .A2(sram_rdata_7[3]), .A3(n15900), .A4(
        sram_rdata_6[3]), .A5(n16400), .A6(sram_rdata_8[3]), .Y(n1327) );
  AOI22X1_HVT U1015 ( .A1(n954), .A2(n15000), .A3(n578), .A4(n1327), .Y(n957)
         );
  OA22X1_HVT U1016 ( .A1(n2770), .A2(n416), .A3(n11500), .A4(n3210), .Y(n956)
         );
  NAND2X0_HVT U1017 ( .A1(n1770), .A2(sram_rdata_5[3]), .Y(n955) );
  NAND3X0_HVT U1018 ( .A1(n957), .A2(n956), .A3(n955), .Y(n_src_aox[115]) );
  AO222X1_HVT U1019 ( .A1(n1850), .A2(sram_rdata_7[4]), .A3(n2120), .A4(
        sram_rdata_6[4]), .A5(n16400), .A6(sram_rdata_8[4]), .Y(n1332) );
  AOI22X1_HVT U1020 ( .A1(n958), .A2(n10800), .A3(n15100), .A4(n1332), .Y(n961) );
  OA22X1_HVT U1021 ( .A1(n2800), .A2(n417), .A3(n2690), .A4(n3220), .Y(n9601)
         );
  NAND2X0_HVT U1022 ( .A1(n2220), .A2(sram_rdata_5[4]), .Y(n959) );
  NAND3X0_HVT U1023 ( .A1(n961), .A2(n9601), .A3(n959), .Y(n_src_aox[116]) );
  AO222X1_HVT U1024 ( .A1(n1840), .A2(sram_rdata_7[5]), .A3(n13600), .A4(
        sram_rdata_6[5]), .A5(n1700), .A6(sram_rdata_8[5]), .Y(n1337) );
  AOI22X1_HVT U1025 ( .A1(n962), .A2(n10700), .A3(n1648), .A4(n1337), .Y(n965)
         );
  OA22X1_HVT U1026 ( .A1(n2790), .A2(n418), .A3(n2720), .A4(n3230), .Y(n964)
         );
  NAND2X0_HVT U1027 ( .A1(n1750), .A2(sram_rdata_5[5]), .Y(n963) );
  NAND3X0_HVT U1028 ( .A1(n965), .A2(n964), .A3(n963), .Y(n_src_aox[117]) );
  AO222X1_HVT U1029 ( .A1(n2080), .A2(sram_rdata_7[6]), .A3(n15900), .A4(
        sram_rdata_6[6]), .A5(n2020), .A6(sram_rdata_8[6]), .Y(n1342) );
  AOI22X1_HVT U1030 ( .A1(n966), .A2(n589), .A3(n11000), .A4(n1342), .Y(n969)
         );
  OA22X1_HVT U1031 ( .A1(n10600), .A2(n419), .A3(n1661), .A4(n3240), .Y(n968)
         );
  NAND2X0_HVT U1032 ( .A1(n1750), .A2(sram_rdata_5[6]), .Y(n967) );
  NAND3X0_HVT U1033 ( .A1(n969), .A2(n968), .A3(n967), .Y(n_src_aox[118]) );
  AO222X1_HVT U1034 ( .A1(n2070), .A2(sram_rdata_7[7]), .A3(n2180), .A4(
        sram_rdata_6[7]), .A5(n1970), .A6(sram_rdata_8[7]), .Y(n1347) );
  AOI22X1_HVT U1035 ( .A1(n9701), .A2(n15000), .A3(n579), .A4(n1347), .Y(n973)
         );
  OA22X1_HVT U1036 ( .A1(n13800), .A2(n4201), .A3(n2700), .A4(n3250), .Y(n972)
         );
  NAND2X0_HVT U1037 ( .A1(n2210), .A2(sram_rdata_5[7]), .Y(n971) );
  NAND3X0_HVT U1038 ( .A1(n973), .A2(n972), .A3(n971), .Y(n_src_aox[119]) );
  AO222X1_HVT U1039 ( .A1(n2070), .A2(sram_rdata_7[8]), .A3(n15600), .A4(
        sram_rdata_6[8]), .A5(n1940), .A6(sram_rdata_8[8]), .Y(n1349) );
  AOI22X1_HVT U1040 ( .A1(n974), .A2(n15000), .A3(n12900), .A4(n1349), .Y(n977) );
  OA22X1_HVT U1041 ( .A1(n13800), .A2(n421), .A3(n2700), .A4(n3260), .Y(n976)
         );
  NAND2X0_HVT U1042 ( .A1(n1730), .A2(sram_rdata_5[8]), .Y(n975) );
  NAND3X0_HVT U1043 ( .A1(n977), .A2(n976), .A3(n975), .Y(n_src_aox[120]) );
  AO222X1_HVT U1044 ( .A1(n2070), .A2(sram_rdata_7[9]), .A3(n15800), .A4(
        sram_rdata_6[9]), .A5(n2010), .A6(sram_rdata_8[9]), .Y(n1354) );
  AOI22X1_HVT U1045 ( .A1(n978), .A2(n592), .A3(n582), .A4(n1354), .Y(n981) );
  OA22X1_HVT U1046 ( .A1(n13700), .A2(n422), .A3(n2750), .A4(n327), .Y(n9801)
         );
  NAND2X0_HVT U1047 ( .A1(n2280), .A2(sram_rdata_5[9]), .Y(n979) );
  NAND3X0_HVT U1048 ( .A1(n981), .A2(n9801), .A3(n979), .Y(n_src_aox[121]) );
  AO222X1_HVT U1049 ( .A1(n2040), .A2(sram_rdata_7[10]), .A3(n2190), .A4(
        sram_rdata_6[10]), .A5(n1980), .A6(sram_rdata_8[10]), .Y(n1359) );
  AOI22X1_HVT U1050 ( .A1(n982), .A2(n12700), .A3(n15100), .A4(n1359), .Y(n985) );
  OA22X1_HVT U1051 ( .A1(n2760), .A2(n423), .A3(n2720), .A4(n328), .Y(n984) );
  NAND2X0_HVT U1052 ( .A1(n1810), .A2(sram_rdata_5[10]), .Y(n983) );
  NAND3X0_HVT U1053 ( .A1(n985), .A2(n984), .A3(n983), .Y(n_src_aox[122]) );
  AO222X1_HVT U1054 ( .A1(n2050), .A2(sram_rdata_7[11]), .A3(n2170), .A4(
        sram_rdata_6[11]), .A5(n1960), .A6(sram_rdata_8[11]), .Y(n1364) );
  AOI22X1_HVT U1055 ( .A1(n986), .A2(n588), .A3(n15200), .A4(n1364), .Y(n989)
         );
  OA22X1_HVT U1056 ( .A1(n11800), .A2(n424), .A3(n10000), .A4(n329), .Y(n988)
         );
  NAND2X0_HVT U1057 ( .A1(n2230), .A2(sram_rdata_5[11]), .Y(n987) );
  NAND3X0_HVT U1058 ( .A1(n989), .A2(n988), .A3(n987), .Y(n_src_aox[123]) );
  AO222X1_HVT U1059 ( .A1(n1890), .A2(sram_rdata_7[12]), .A3(n2180), .A4(
        sram_rdata_6[12]), .A5(n1710), .A6(sram_rdata_8[12]), .Y(n1369) );
  AOI22X1_HVT U1060 ( .A1(n9901), .A2(n12800), .A3(n582), .A4(n1369), .Y(n993)
         );
  OA22X1_HVT U1061 ( .A1(n11900), .A2(n425), .A3(n2710), .A4(n330), .Y(n992)
         );
  NAND2X0_HVT U1062 ( .A1(n2280), .A2(sram_rdata_5[12]), .Y(n991) );
  NAND3X0_HVT U1063 ( .A1(n993), .A2(n992), .A3(n991), .Y(n_src_aox[124]) );
  AO222X1_HVT U1064 ( .A1(n2030), .A2(sram_rdata_7[13]), .A3(n2140), .A4(
        sram_rdata_6[13]), .A5(n16500), .A6(sram_rdata_8[13]), .Y(n1374) );
  AOI22X1_HVT U1065 ( .A1(n994), .A2(n14900), .A3(n15200), .A4(n1374), .Y(n997) );
  OA22X1_HVT U1066 ( .A1(n10400), .A2(n426), .A3(n2740), .A4(n331), .Y(n996)
         );
  NAND2X0_HVT U1067 ( .A1(n1800), .A2(sram_rdata_5[13]), .Y(n995) );
  NAND3X0_HVT U1068 ( .A1(n997), .A2(n996), .A3(n995), .Y(n_src_aox[125]) );
  AO222X1_HVT U1069 ( .A1(n2060), .A2(sram_rdata_7[14]), .A3(n1658), .A4(
        sram_rdata_6[14]), .A5(n1710), .A6(sram_rdata_8[14]), .Y(n1379) );
  AOI22X1_HVT U1070 ( .A1(n998), .A2(n14900), .A3(n582), .A4(n1379), .Y(n1001)
         );
  OA22X1_HVT U1071 ( .A1(n2780), .A2(n427), .A3(n10100), .A4(n332), .Y(n10001)
         );
  NAND2X0_HVT U1072 ( .A1(n576), .A2(sram_rdata_5[14]), .Y(n999) );
  NAND3X0_HVT U1073 ( .A1(n1001), .A2(n10001), .A3(n999), .Y(n_src_aox[126])
         );
  AO222X1_HVT U1074 ( .A1(n2060), .A2(sram_rdata_7[15]), .A3(n2180), .A4(
        sram_rdata_6[15]), .A5(n1980), .A6(sram_rdata_8[15]), .Y(n1384) );
  AOI22X1_HVT U1075 ( .A1(n1002), .A2(n589), .A3(n579), .A4(n1384), .Y(n1005)
         );
  OA22X1_HVT U1076 ( .A1(n10300), .A2(n428), .A3(n2700), .A4(n333), .Y(n1004)
         );
  NAND2X0_HVT U1077 ( .A1(n1750), .A2(sram_rdata_5[15]), .Y(n1003) );
  NAND3X0_HVT U1078 ( .A1(n1005), .A2(n1004), .A3(n1003), .Y(n_src_aox[127])
         );
  AO222X1_HVT U1079 ( .A1(sram_rdata_6[0]), .A2(n2080), .A3(sram_rdata_8[0]), 
        .A4(n2180), .A5(n1930), .A6(sram_rdata_7[0]), .Y(n13901) );
  AOI22X1_HVT U1080 ( .A1(n13901), .A2(n11000), .A3(n5901), .A4(n1006), .Y(
        n1009) );
  OA22X1_HVT U1081 ( .A1(n12000), .A2(n478), .A3(n11500), .A4(n382), .Y(n1008)
         );
  NAND2X0_HVT U1082 ( .A1(n2270), .A2(sram_rdata_4[0]), .Y(n1007) );
  NAND3X0_HVT U1083 ( .A1(n1009), .A2(n1008), .A3(n1007), .Y(n_src_aox[128])
         );
  AO222X1_HVT U1084 ( .A1(n1910), .A2(sram_rdata_6[1]), .A3(n2110), .A4(
        sram_rdata_8[1]), .A5(sram_rdata_7[1]), .A6(n1980), .Y(n1391) );
  AO222X1_HVT U1085 ( .A1(n1910), .A2(sram_rdata_6[2]), .A3(n16100), .A4(
        sram_rdata_8[2]), .A5(sram_rdata_7[2]), .A6(n1930), .Y(n1396) );
  AOI22X1_HVT U1086 ( .A1(n1011), .A2(n588), .A3(n579), .A4(n1396), .Y(n1014)
         );
  OA22X1_HVT U1087 ( .A1(n12100), .A2(n511), .A3(n14700), .A4(n415), .Y(n1013)
         );
  NAND2X0_HVT U1088 ( .A1(n2220), .A2(sram_rdata_4[2]), .Y(n1012) );
  NAND3X0_HVT U1089 ( .A1(n1014), .A2(n1013), .A3(n1012), .Y(n_src_aox[130])
         );
  AO222X1_HVT U1090 ( .A1(n2100), .A2(sram_rdata_6[3]), .A3(n15700), .A4(
        sram_rdata_8[3]), .A5(sram_rdata_7[3]), .A6(n16500), .Y(n1401) );
  AOI22X1_HVT U1091 ( .A1(n1015), .A2(n10700), .A3(n5801), .A4(n1401), .Y(
        n1018) );
  OA22X1_HVT U1092 ( .A1(n2780), .A2(n512), .A3(n2700), .A4(n416), .Y(n1017)
         );
  NAND2X0_HVT U1093 ( .A1(n1770), .A2(sram_rdata_4[3]), .Y(n1016) );
  NAND3X0_HVT U1094 ( .A1(n1018), .A2(n1017), .A3(n1016), .Y(n_src_aox[131])
         );
  AO222X1_HVT U1095 ( .A1(n1659), .A2(sram_rdata_6[4]), .A3(n13600), .A4(
        sram_rdata_8[4]), .A5(sram_rdata_7[4]), .A6(n1930), .Y(n1406) );
  AOI22X1_HVT U1096 ( .A1(n1019), .A2(n12800), .A3(n582), .A4(n1406), .Y(n1022) );
  OA22X1_HVT U1097 ( .A1(n2810), .A2(n513), .A3(n10000), .A4(n417), .Y(n1021)
         );
  NAND2X0_HVT U1098 ( .A1(n1740), .A2(sram_rdata_4[4]), .Y(n10201) );
  NAND3X0_HVT U1099 ( .A1(n1022), .A2(n1021), .A3(n10201), .Y(n_src_aox[132])
         );
  AO222X1_HVT U1100 ( .A1(n1890), .A2(sram_rdata_6[5]), .A3(n16000), .A4(
        sram_rdata_8[5]), .A5(sram_rdata_7[5]), .A6(n1700), .Y(n1411) );
  AOI22X1_HVT U1101 ( .A1(n1023), .A2(n15000), .A3(n10900), .A4(n1411), .Y(
        n1026) );
  OA22X1_HVT U1102 ( .A1(n2790), .A2(n514), .A3(n10100), .A4(n418), .Y(n1025)
         );
  NAND2X0_HVT U1103 ( .A1(n1810), .A2(sram_rdata_4[5]), .Y(n1024) );
  NAND3X0_HVT U1104 ( .A1(n1026), .A2(n1025), .A3(n1024), .Y(n_src_aox[133])
         );
  AO222X1_HVT U1105 ( .A1(n2030), .A2(sram_rdata_6[6]), .A3(n15600), .A4(
        sram_rdata_8[6]), .A5(sram_rdata_7[6]), .A6(n1710), .Y(n1416) );
  AOI22X1_HVT U1106 ( .A1(n1027), .A2(n12800), .A3(n15100), .A4(n1416), .Y(
        n10301) );
  OA22X1_HVT U1107 ( .A1(n11800), .A2(n515), .A3(n2740), .A4(n419), .Y(n1029)
         );
  NAND2X0_HVT U1108 ( .A1(n1750), .A2(sram_rdata_4[6]), .Y(n1028) );
  NAND3X0_HVT U1109 ( .A1(n10301), .A2(n1029), .A3(n1028), .Y(n_src_aox[134])
         );
  AO222X1_HVT U1110 ( .A1(n2040), .A2(sram_rdata_6[7]), .A3(n2170), .A4(
        sram_rdata_8[7]), .A5(sram_rdata_7[7]), .A6(n1710), .Y(n1418) );
  AOI22X1_HVT U1111 ( .A1(n1031), .A2(n10800), .A3(n15200), .A4(n1418), .Y(
        n1034) );
  OA22X1_HVT U1112 ( .A1(n13700), .A2(n516), .A3(n14500), .A4(n4201), .Y(n1033) );
  NAND2X0_HVT U1113 ( .A1(n2270), .A2(sram_rdata_4[7]), .Y(n1032) );
  NAND3X0_HVT U1114 ( .A1(n1034), .A2(n1033), .A3(n1032), .Y(n_src_aox[135])
         );
  AO222X1_HVT U1115 ( .A1(n13900), .A2(sram_rdata_6[8]), .A3(n16100), .A4(
        sram_rdata_8[8]), .A5(sram_rdata_7[8]), .A6(n1670), .Y(n1423) );
  AOI22X1_HVT U1116 ( .A1(n1035), .A2(n14900), .A3(n15200), .A4(n1423), .Y(
        n1038) );
  OA22X1_HVT U1117 ( .A1(n13800), .A2(n517), .A3(n11500), .A4(n421), .Y(n1037)
         );
  NAND2X0_HVT U1118 ( .A1(n1800), .A2(sram_rdata_4[8]), .Y(n1036) );
  NAND3X0_HVT U1119 ( .A1(n1038), .A2(n1037), .A3(n1036), .Y(n_src_aox[136])
         );
  AO222X1_HVT U1120 ( .A1(n1850), .A2(sram_rdata_6[9]), .A3(n15500), .A4(
        sram_rdata_8[9]), .A5(sram_rdata_7[9]), .A6(n1680), .Y(n1428) );
  AOI22X1_HVT U1121 ( .A1(n1039), .A2(n589), .A3(n11000), .A4(n1428), .Y(n1042) );
  OA22X1_HVT U1122 ( .A1(n2800), .A2(n518), .A3(n1661), .A4(n422), .Y(n1041)
         );
  NAND2X0_HVT U1123 ( .A1(n1720), .A2(sram_rdata_4[9]), .Y(n10401) );
  NAND3X0_HVT U1124 ( .A1(n1042), .A2(n1041), .A3(n10401), .Y(n_src_aox[137])
         );
  AO222X1_HVT U1125 ( .A1(n2070), .A2(sram_rdata_6[10]), .A3(n2110), .A4(
        sram_rdata_8[10]), .A5(sram_rdata_7[10]), .A6(n1670), .Y(n1433) );
  AOI22X1_HVT U1126 ( .A1(n1043), .A2(n591), .A3(n12600), .A4(n1433), .Y(n1046) );
  OA22X1_HVT U1127 ( .A1(n1662), .A2(n519), .A3(n10100), .A4(n423), .Y(n1045)
         );
  NAND2X0_HVT U1128 ( .A1(n2210), .A2(sram_rdata_4[10]), .Y(n1044) );
  NAND3X0_HVT U1129 ( .A1(n1046), .A2(n1045), .A3(n1044), .Y(n_src_aox[138])
         );
  AO222X1_HVT U1130 ( .A1(n1830), .A2(sram_rdata_6[11]), .A3(n15700), .A4(
        sram_rdata_8[11]), .A5(sram_rdata_7[11]), .A6(n1690), .Y(n1438) );
  AOI22X1_HVT U1131 ( .A1(n1047), .A2(n12800), .A3(n12900), .A4(n1438), .Y(
        n10501) );
  OA22X1_HVT U1132 ( .A1(n10600), .A2(n5201), .A3(n2700), .A4(n424), .Y(n1049)
         );
  NAND2X0_HVT U1133 ( .A1(n1760), .A2(sram_rdata_4[11]), .Y(n1048) );
  NAND3X0_HVT U1134 ( .A1(n10501), .A2(n1049), .A3(n1048), .Y(n_src_aox[139])
         );
  AO222X1_HVT U1135 ( .A1(n1830), .A2(sram_rdata_6[12]), .A3(n15700), .A4(
        sram_rdata_8[12]), .A5(sram_rdata_7[12]), .A6(n2000), .Y(n1443) );
  AOI22X1_HVT U1136 ( .A1(n1051), .A2(n588), .A3(n582), .A4(n1443), .Y(n1054)
         );
  OA22X1_HVT U1137 ( .A1(n10500), .A2(n521), .A3(n2690), .A4(n425), .Y(n1053)
         );
  NAND2X0_HVT U1138 ( .A1(n1790), .A2(sram_rdata_4[12]), .Y(n1052) );
  NAND3X0_HVT U1139 ( .A1(n1054), .A2(n1053), .A3(n1052), .Y(n_src_aox[140])
         );
  AO222X1_HVT U1140 ( .A1(n1830), .A2(sram_rdata_6[13]), .A3(n2140), .A4(
        sram_rdata_8[13]), .A5(sram_rdata_7[13]), .A6(n1970), .Y(n1448) );
  AOI22X1_HVT U1141 ( .A1(n1055), .A2(n12700), .A3(n15200), .A4(n1448), .Y(
        n1058) );
  OA22X1_HVT U1142 ( .A1(n10400), .A2(n522), .A3(n2740), .A4(n426), .Y(n1057)
         );
  NAND2X0_HVT U1143 ( .A1(n1720), .A2(sram_rdata_4[13]), .Y(n1056) );
  NAND3X0_HVT U1144 ( .A1(n1058), .A2(n1057), .A3(n1056), .Y(n_src_aox[141])
         );
  AO222X1_HVT U1145 ( .A1(n1840), .A2(sram_rdata_6[14]), .A3(n2140), .A4(
        sram_rdata_8[14]), .A5(sram_rdata_7[14]), .A6(n1920), .Y(n1453) );
  AOI22X1_HVT U1146 ( .A1(n1059), .A2(n591), .A3(n10900), .A4(n1453), .Y(n1062) );
  OA22X1_HVT U1147 ( .A1(n13700), .A2(n523), .A3(n2750), .A4(n427), .Y(n1061)
         );
  NAND2X0_HVT U1148 ( .A1(n2260), .A2(sram_rdata_4[14]), .Y(n10601) );
  NAND3X0_HVT U1149 ( .A1(n1062), .A2(n1061), .A3(n10601), .Y(n_src_aox[142])
         );
  AO222X1_HVT U1150 ( .A1(n2090), .A2(sram_rdata_6[15]), .A3(n2130), .A4(
        sram_rdata_8[15]), .A5(sram_rdata_7[15]), .A6(n2020), .Y(n1455) );
  AOI22X1_HVT U1151 ( .A1(n1063), .A2(n588), .A3(n15100), .A4(n1455), .Y(n1066) );
  OA22X1_HVT U1152 ( .A1(n10300), .A2(n524), .A3(n11500), .A4(n428), .Y(n1065)
         );
  NAND2X0_HVT U1153 ( .A1(n2260), .A2(sram_rdata_4[15]), .Y(n1064) );
  NAND3X0_HVT U1154 ( .A1(n1066), .A2(n1065), .A3(n1064), .Y(n_src_aox[143])
         );
  AO222X1_HVT U1155 ( .A1(n1890), .A2(sram_rdata_8[16]), .A3(n16100), .A4(
        sram_rdata_7[16]), .A5(sram_rdata_6[16]), .A6(n2000), .Y(n14601) );
  AOI22X1_HVT U1156 ( .A1(n1067), .A2(n591), .A3(n15100), .A4(n14601), .Y(
        n10701) );
  OA22X1_HVT U1157 ( .A1(n12000), .A2(n334), .A3(n14600), .A4(n525), .Y(n1069)
         );
  NAND2X0_HVT U1158 ( .A1(n1730), .A2(sram_rdata_3[16]), .Y(n1068) );
  NAND3X0_HVT U1159 ( .A1(n10701), .A2(n1069), .A3(n1068), .Y(n_src_aox[144])
         );
  AO222X1_HVT U1160 ( .A1(n1900), .A2(sram_rdata_8[17]), .A3(n16100), .A4(
        sram_rdata_7[17]), .A5(sram_rdata_6[17]), .A6(n1980), .Y(n1465) );
  AOI22X1_HVT U1161 ( .A1(n1071), .A2(n14900), .A3(n579), .A4(n1465), .Y(n1074) );
  OA22X1_HVT U1162 ( .A1(n10500), .A2(n335), .A3(n2720), .A4(n526), .Y(n1073)
         );
  NAND2X0_HVT U1163 ( .A1(n2240), .A2(sram_rdata_3[17]), .Y(n1072) );
  NAND3X0_HVT U1164 ( .A1(n1074), .A2(n1073), .A3(n1072), .Y(n_src_aox[145])
         );
  AO222X1_HVT U1165 ( .A1(n1860), .A2(sram_rdata_8[18]), .A3(n15700), .A4(
        sram_rdata_7[18]), .A5(sram_rdata_6[18]), .A6(n16600), .Y(n14701) );
  AOI22X1_HVT U1166 ( .A1(n1075), .A2(n591), .A3(n5801), .A4(n14701), .Y(n1078) );
  OA22X1_HVT U1167 ( .A1(n12100), .A2(n336), .A3(n2720), .A4(n527), .Y(n1077)
         );
  NAND2X0_HVT U1168 ( .A1(n2280), .A2(sram_rdata_3[18]), .Y(n1076) );
  NAND3X0_HVT U1169 ( .A1(n1078), .A2(n1077), .A3(n1076), .Y(n_src_aox[146])
         );
  AO222X1_HVT U1170 ( .A1(n2030), .A2(sram_rdata_8[19]), .A3(n2160), .A4(
        sram_rdata_7[19]), .A5(sram_rdata_6[19]), .A6(n1680), .Y(n1475) );
  AOI22X1_HVT U1171 ( .A1(n1079), .A2(n10800), .A3(n11000), .A4(n1475), .Y(
        n1082) );
  OA22X1_HVT U1172 ( .A1(n2780), .A2(n337), .A3(n14500), .A4(n528), .Y(n1081)
         );
  NAND2X0_HVT U1173 ( .A1(n574), .A2(sram_rdata_3[19]), .Y(n10801) );
  NAND3X0_HVT U1174 ( .A1(n1082), .A2(n1081), .A3(n10801), .Y(n_src_aox[147])
         );
  AO222X1_HVT U1175 ( .A1(n12500), .A2(sram_rdata_8[20]), .A3(n15700), .A4(
        sram_rdata_7[20]), .A5(sram_rdata_6[20]), .A6(n16400), .Y(n14801) );
  AOI22X1_HVT U1176 ( .A1(n1083), .A2(n14900), .A3(n15200), .A4(n14801), .Y(
        n1086) );
  OA22X1_HVT U1177 ( .A1(n2800), .A2(n338), .A3(n2710), .A4(n529), .Y(n1085)
         );
  NAND2X0_HVT U1178 ( .A1(n1790), .A2(sram_rdata_3[20]), .Y(n1084) );
  NAND3X0_HVT U1179 ( .A1(n1086), .A2(n1085), .A3(n1084), .Y(n_src_aox[148])
         );
  AO222X1_HVT U1180 ( .A1(n1880), .A2(sram_rdata_8[21]), .A3(n13500), .A4(
        sram_rdata_7[21]), .A5(sram_rdata_6[21]), .A6(n1990), .Y(n1485) );
  AOI22X1_HVT U1181 ( .A1(n1087), .A2(n589), .A3(n582), .A4(n1485), .Y(n10901)
         );
  OA22X1_HVT U1182 ( .A1(n2790), .A2(n339), .A3(n2720), .A4(n5301), .Y(n1089)
         );
  NAND2X0_HVT U1183 ( .A1(n575), .A2(sram_rdata_3[21]), .Y(n1088) );
  NAND3X0_HVT U1184 ( .A1(n10901), .A2(n1089), .A3(n1088), .Y(n_src_aox[149])
         );
  AO222X1_HVT U1185 ( .A1(n1880), .A2(sram_rdata_8[22]), .A3(n15900), .A4(
        sram_rdata_7[22]), .A5(sram_rdata_6[22]), .A6(n1920), .Y(n14901) );
  AOI22X1_HVT U1186 ( .A1(n1091), .A2(n14900), .A3(n582), .A4(n14901), .Y(
        n1094) );
  OA22X1_HVT U1187 ( .A1(n11800), .A2(n340), .A3(n14800), .A4(n531), .Y(n1093)
         );
  NAND2X0_HVT U1188 ( .A1(n2250), .A2(sram_rdata_3[22]), .Y(n1092) );
  NAND3X0_HVT U1189 ( .A1(n1094), .A2(n1093), .A3(n1092), .Y(n_src_aox[150])
         );
  AO222X1_HVT U1190 ( .A1(n1840), .A2(sram_rdata_8[23]), .A3(n15400), .A4(
        sram_rdata_7[23]), .A5(sram_rdata_6[23]), .A6(n1700), .Y(n1495) );
  AOI22X1_HVT U1191 ( .A1(n1095), .A2(n589), .A3(n12600), .A4(n1495), .Y(n1098) );
  OA22X1_HVT U1192 ( .A1(n2760), .A2(n341), .A3(n2700), .A4(n532), .Y(n1097)
         );
  NAND2X0_HVT U1193 ( .A1(n1770), .A2(sram_rdata_3[23]), .Y(n1096) );
  NAND3X0_HVT U1194 ( .A1(n1098), .A2(n1097), .A3(n1096), .Y(n_src_aox[151])
         );
  AO222X1_HVT U1195 ( .A1(n1830), .A2(sram_rdata_8[24]), .A3(n15700), .A4(
        sram_rdata_7[24]), .A5(sram_rdata_6[24]), .A6(n2010), .Y(n15001) );
  AOI22X1_HVT U1196 ( .A1(n1099), .A2(n15000), .A3(n12600), .A4(n15001), .Y(
        n1102) );
  OA22X1_HVT U1197 ( .A1(n2790), .A2(n342), .A3(n2700), .A4(n533), .Y(n1101)
         );
  NAND2X0_HVT U1198 ( .A1(n2240), .A2(sram_rdata_3[24]), .Y(n11001) );
  NAND3X0_HVT U1199 ( .A1(n1102), .A2(n1101), .A3(n11001), .Y(n_src_aox[152])
         );
  AO222X1_HVT U1200 ( .A1(n13900), .A2(sram_rdata_8[25]), .A3(n2130), .A4(
        sram_rdata_7[25]), .A5(sram_rdata_6[25]), .A6(n1960), .Y(n1502) );
  AOI22X1_HVT U1201 ( .A1(n1103), .A2(n10800), .A3(n15200), .A4(n1502), .Y(
        n1106) );
  OA22X1_HVT U1202 ( .A1(n2810), .A2(n343), .A3(n14800), .A4(n534), .Y(n1105)
         );
  NAND2X0_HVT U1203 ( .A1(n1810), .A2(sram_rdata_3[25]), .Y(n1104) );
  NAND3X0_HVT U1204 ( .A1(n1106), .A2(n1105), .A3(n1104), .Y(n_src_aox[153])
         );
  AO222X1_HVT U1205 ( .A1(n2100), .A2(sram_rdata_8[26]), .A3(n16000), .A4(
        sram_rdata_7[26]), .A5(sram_rdata_6[26]), .A6(n1940), .Y(n1507) );
  AO222X1_HVT U1206 ( .A1(n2080), .A2(sram_rdata_8[27]), .A3(n15400), .A4(
        sram_rdata_7[27]), .A5(sram_rdata_6[27]), .A6(n1930), .Y(n1512) );
  AOI22X1_HVT U1207 ( .A1(n1108), .A2(n589), .A3(n12900), .A4(n1512), .Y(n1111) );
  OA22X1_HVT U1208 ( .A1(n10600), .A2(n345), .A3(n14600), .A4(n536), .Y(n11101) );
  NAND2X0_HVT U1209 ( .A1(n2230), .A2(sram_rdata_3[27]), .Y(n1109) );
  NAND3X0_HVT U1210 ( .A1(n1111), .A2(n11101), .A3(n1109), .Y(n_src_aox[155])
         );
  AO222X1_HVT U1211 ( .A1(n2090), .A2(sram_rdata_8[28]), .A3(n2180), .A4(
        sram_rdata_7[28]), .A5(sram_rdata_6[28]), .A6(n1670), .Y(n1514) );
  AOI22X1_HVT U1212 ( .A1(n1112), .A2(n588), .A3(n582), .A4(n1514), .Y(n1115)
         );
  OA22X1_HVT U1213 ( .A1(n10500), .A2(n3460), .A3(n10000), .A4(n537), .Y(n1114) );
  NAND2X0_HVT U1214 ( .A1(n574), .A2(sram_rdata_3[28]), .Y(n1113) );
  NAND3X0_HVT U1215 ( .A1(n1115), .A2(n1114), .A3(n1113), .Y(n_src_aox[156])
         );
  AO222X1_HVT U1216 ( .A1(n2080), .A2(sram_rdata_8[29]), .A3(n15700), .A4(
        sram_rdata_7[29]), .A5(sram_rdata_6[29]), .A6(n1680), .Y(n1519) );
  AOI22X1_HVT U1217 ( .A1(n1116), .A2(n589), .A3(n11000), .A4(n1519), .Y(n1119) );
  OA22X1_HVT U1218 ( .A1(n10400), .A2(n347), .A3(n10100), .A4(n538), .Y(n1118)
         );
  NAND2X0_HVT U1219 ( .A1(n2280), .A2(sram_rdata_3[29]), .Y(n1117) );
  NAND3X0_HVT U1220 ( .A1(n1119), .A2(n1118), .A3(n1117), .Y(n_src_aox[157])
         );
  AO222X1_HVT U1221 ( .A1(n2080), .A2(sram_rdata_8[30]), .A3(n15900), .A4(
        sram_rdata_7[30]), .A5(sram_rdata_6[30]), .A6(n1680), .Y(n1524) );
  AOI22X1_HVT U1222 ( .A1(n11201), .A2(n15000), .A3(n582), .A4(n1524), .Y(
        n1123) );
  OA22X1_HVT U1223 ( .A1(n2770), .A2(n348), .A3(n2740), .A4(n539), .Y(n1122)
         );
  NAND2X0_HVT U1224 ( .A1(n1740), .A2(sram_rdata_3[30]), .Y(n1121) );
  NAND3X0_HVT U1225 ( .A1(n1123), .A2(n1122), .A3(n1121), .Y(n_src_aox[158])
         );
  AO222X1_HVT U1226 ( .A1(n2060), .A2(sram_rdata_8[31]), .A3(n2190), .A4(
        sram_rdata_7[31]), .A5(sram_rdata_6[31]), .A6(n16400), .Y(n1529) );
  AOI22X1_HVT U1227 ( .A1(n1124), .A2(n12700), .A3(n12600), .A4(n1529), .Y(
        n1127) );
  OA22X1_HVT U1228 ( .A1(n10300), .A2(n349), .A3(n14500), .A4(n5401), .Y(n1126) );
  NAND2X0_HVT U1229 ( .A1(n2230), .A2(sram_rdata_3[31]), .Y(n1125) );
  NAND3X0_HVT U1230 ( .A1(n1127), .A2(n1126), .A3(n1125), .Y(n_src_aox[159])
         );
  AO222X1_HVT U1231 ( .A1(n1910), .A2(sram_rdata_7[16]), .A3(n2160), .A4(
        sram_rdata_6[16]), .A5(n16600), .A6(sram_rdata_8[16]), .Y(n1531) );
  AOI22X1_HVT U1232 ( .A1(n1128), .A2(n10700), .A3(n10900), .A4(n1531), .Y(
        n1131) );
  OA22X1_HVT U1233 ( .A1(n12000), .A2(n429), .A3(n14600), .A4(n334), .Y(n11301) );
  NAND2X0_HVT U1234 ( .A1(n1740), .A2(sram_rdata_5[16]), .Y(n1129) );
  NAND3X0_HVT U1235 ( .A1(n1131), .A2(n11301), .A3(n1129), .Y(n_src_aox[160])
         );
  AO222X1_HVT U1236 ( .A1(n1850), .A2(sram_rdata_7[17]), .A3(n2170), .A4(
        sram_rdata_6[17]), .A5(n2020), .A6(sram_rdata_8[17]), .Y(n1536) );
  AOI22X1_HVT U1237 ( .A1(n1132), .A2(n589), .A3(n5801), .A4(n1536), .Y(n1135)
         );
  OA22X1_HVT U1238 ( .A1(n10500), .A2(n4301), .A3(n14700), .A4(n335), .Y(n1134) );
  NAND2X0_HVT U1239 ( .A1(n1750), .A2(sram_rdata_5[17]), .Y(n1133) );
  NAND3X0_HVT U1240 ( .A1(n1135), .A2(n1134), .A3(n1133), .Y(n_src_aox[161])
         );
  AO222X1_HVT U1241 ( .A1(n2050), .A2(sram_rdata_7[18]), .A3(n15900), .A4(
        sram_rdata_6[18]), .A5(n1980), .A6(sram_rdata_8[18]), .Y(n1541) );
  AOI22X1_HVT U1242 ( .A1(n1136), .A2(n12800), .A3(n15100), .A4(n1541), .Y(
        n1139) );
  OA22X1_HVT U1243 ( .A1(n10300), .A2(n431), .A3(n10100), .A4(n336), .Y(n1138)
         );
  NAND2X0_HVT U1244 ( .A1(n1720), .A2(sram_rdata_5[18]), .Y(n1137) );
  NAND3X0_HVT U1245 ( .A1(n1139), .A2(n1138), .A3(n1137), .Y(n_src_aox[162])
         );
  AO222X1_HVT U1246 ( .A1(n2050), .A2(sram_rdata_7[19]), .A3(n1658), .A4(
        sram_rdata_6[19]), .A5(n2000), .A6(sram_rdata_8[19]), .Y(n1543) );
  AOI22X1_HVT U1247 ( .A1(n11401), .A2(n588), .A3(n15200), .A4(n1543), .Y(
        n1143) );
  OA22X1_HVT U1248 ( .A1(n2770), .A2(n432), .A3(n14500), .A4(n337), .Y(n1142)
         );
  NAND2X0_HVT U1249 ( .A1(n1740), .A2(sram_rdata_5[19]), .Y(n1141) );
  NAND3X0_HVT U1250 ( .A1(n1143), .A2(n1142), .A3(n1141), .Y(n_src_aox[163])
         );
  AO222X1_HVT U1251 ( .A1(n2030), .A2(sram_rdata_7[20]), .A3(n15600), .A4(
        sram_rdata_6[20]), .A5(n1920), .A6(sram_rdata_8[20]), .Y(n1548) );
  AOI22X1_HVT U1252 ( .A1(n1144), .A2(n588), .A3(n579), .A4(n1548), .Y(n1147)
         );
  OA22X1_HVT U1253 ( .A1(n2810), .A2(n433), .A3(n14500), .A4(n338), .Y(n1146)
         );
  NAND2X0_HVT U1254 ( .A1(n2250), .A2(sram_rdata_5[20]), .Y(n1145) );
  NAND3X0_HVT U1255 ( .A1(n1147), .A2(n1146), .A3(n1145), .Y(n_src_aox[164])
         );
  AO222X1_HVT U1256 ( .A1(n1880), .A2(sram_rdata_7[21]), .A3(n2120), .A4(
        sram_rdata_6[21]), .A5(n1680), .A6(sram_rdata_8[21]), .Y(n1553) );
  AOI22X1_HVT U1257 ( .A1(n1148), .A2(n12700), .A3(n12900), .A4(n1553), .Y(
        n1151) );
  OA22X1_HVT U1258 ( .A1(n2790), .A2(n434), .A3(n14800), .A4(n339), .Y(n11501)
         );
  NAND2X0_HVT U1259 ( .A1(n576), .A2(sram_rdata_5[21]), .Y(n1149) );
  NAND3X0_HVT U1260 ( .A1(n1151), .A2(n11501), .A3(n1149), .Y(n_src_aox[165])
         );
  AO222X1_HVT U1261 ( .A1(n1860), .A2(sram_rdata_7[22]), .A3(n1658), .A4(
        sram_rdata_6[22]), .A5(n1700), .A6(sram_rdata_8[22]), .Y(n1558) );
  AOI22X1_HVT U1262 ( .A1(n1152), .A2(n5901), .A3(n582), .A4(n1558), .Y(n1155)
         );
  OA22X1_HVT U1263 ( .A1(n10600), .A2(n435), .A3(n2730), .A4(n340), .Y(n1154)
         );
  NAND2X0_HVT U1264 ( .A1(n2220), .A2(sram_rdata_5[22]), .Y(n1153) );
  NAND3X0_HVT U1265 ( .A1(n1155), .A2(n1154), .A3(n1153), .Y(n_src_aox[166])
         );
  AO222X1_HVT U1266 ( .A1(n2070), .A2(sram_rdata_7[23]), .A3(n15900), .A4(
        sram_rdata_6[23]), .A5(n1690), .A6(sram_rdata_8[23]), .Y(n1563) );
  AOI22X1_HVT U1267 ( .A1(n1156), .A2(n589), .A3(n5801), .A4(n1563), .Y(n1159)
         );
  OA22X1_HVT U1268 ( .A1(n13800), .A2(n436), .A3(n10000), .A4(n341), .Y(n1158)
         );
  NAND2X0_HVT U1269 ( .A1(n574), .A2(sram_rdata_5[23]), .Y(n1157) );
  NAND3X0_HVT U1270 ( .A1(n1159), .A2(n1158), .A3(n1157), .Y(n_src_aox[167])
         );
  AO222X1_HVT U1271 ( .A1(n1880), .A2(sram_rdata_7[24]), .A3(n16100), .A4(
        sram_rdata_6[24]), .A5(n16600), .A6(sram_rdata_8[24]), .Y(n1568) );
  AOI22X1_HVT U1272 ( .A1(n11601), .A2(n588), .A3(n15100), .A4(n1568), .Y(
        n1163) );
  OA22X1_HVT U1273 ( .A1(n13700), .A2(n437), .A3(n2700), .A4(n342), .Y(n1162)
         );
  NAND2X0_HVT U1274 ( .A1(n1760), .A2(sram_rdata_5[24]), .Y(n1161) );
  NAND3X0_HVT U1275 ( .A1(n1163), .A2(n1162), .A3(n1161), .Y(n_src_aox[168])
         );
  AO222X1_HVT U1276 ( .A1(n1890), .A2(sram_rdata_7[25]), .A3(n1658), .A4(
        sram_rdata_6[25]), .A5(n16500), .A6(sram_rdata_8[25]), .Y(n15701) );
  AO222X1_HVT U1277 ( .A1(n1890), .A2(sram_rdata_7[26]), .A3(n2190), .A4(
        sram_rdata_6[26]), .A5(n1670), .A6(sram_rdata_8[26]), .Y(n1572) );
  AOI22X1_HVT U1278 ( .A1(n1165), .A2(n14900), .A3(n15200), .A4(n1572), .Y(
        n1168) );
  OA22X1_HVT U1279 ( .A1(n2760), .A2(n439), .A3(n2720), .A4(n344), .Y(n1167)
         );
  NAND2X0_HVT U1280 ( .A1(n1810), .A2(sram_rdata_5[26]), .Y(n1166) );
  NAND3X0_HVT U1281 ( .A1(n1168), .A2(n1167), .A3(n1166), .Y(n_src_aox[170])
         );
  AO222X1_HVT U1282 ( .A1(n2050), .A2(sram_rdata_7[27]), .A3(n2180), .A4(
        sram_rdata_6[27]), .A5(n2000), .A6(sram_rdata_8[27]), .Y(n1574) );
  AOI22X1_HVT U1283 ( .A1(n1169), .A2(n10800), .A3(n15200), .A4(n1574), .Y(
        n1172) );
  OA22X1_HVT U1284 ( .A1(n11800), .A2(n4401), .A3(n2690), .A4(n345), .Y(n1171)
         );
  NAND2X0_HVT U1285 ( .A1(n2270), .A2(sram_rdata_5[27]), .Y(n11701) );
  NAND3X0_HVT U1286 ( .A1(n1172), .A2(n1171), .A3(n11701), .Y(n_src_aox[171])
         );
  AO222X1_HVT U1287 ( .A1(n1830), .A2(sram_rdata_7[28]), .A3(n15400), .A4(
        sram_rdata_6[28]), .A5(n1990), .A6(sram_rdata_8[28]), .Y(n1579) );
  AOI22X1_HVT U1288 ( .A1(n1173), .A2(n12800), .A3(n5801), .A4(n1579), .Y(
        n1176) );
  OA22X1_HVT U1289 ( .A1(n10500), .A2(n441), .A3(n11500), .A4(n3460), .Y(n1175) );
  NAND2X0_HVT U1290 ( .A1(n1770), .A2(sram_rdata_5[28]), .Y(n1174) );
  NAND3X0_HVT U1291 ( .A1(n1176), .A2(n1175), .A3(n1174), .Y(n_src_aox[172])
         );
  AO222X1_HVT U1292 ( .A1(n1900), .A2(sram_rdata_7[29]), .A3(n2110), .A4(
        sram_rdata_6[29]), .A5(n2010), .A6(sram_rdata_8[29]), .Y(n1584) );
  AOI22X1_HVT U1293 ( .A1(n1177), .A2(n10700), .A3(n11000), .A4(n1584), .Y(
        n11801) );
  OA22X1_HVT U1294 ( .A1(n10400), .A2(n442), .A3(n2720), .A4(n347), .Y(n1179)
         );
  NAND2X0_HVT U1295 ( .A1(n575), .A2(sram_rdata_5[29]), .Y(n1178) );
  NAND3X0_HVT U1296 ( .A1(n11801), .A2(n1179), .A3(n1178), .Y(n_src_aox[173])
         );
  AO222X1_HVT U1297 ( .A1(n2030), .A2(sram_rdata_7[30]), .A3(n2140), .A4(
        sram_rdata_6[30]), .A5(n1990), .A6(sram_rdata_8[30]), .Y(n1589) );
  AO222X1_HVT U1298 ( .A1(n13900), .A2(sram_rdata_7[31]), .A3(n15800), .A4(
        sram_rdata_6[31]), .A5(n1930), .A6(sram_rdata_8[31]), .Y(n1591) );
  AOI22X1_HVT U1299 ( .A1(n1182), .A2(n591), .A3(n11000), .A4(n1591), .Y(n1185) );
  OA22X1_HVT U1300 ( .A1(n12100), .A2(n444), .A3(n14600), .A4(n349), .Y(n1184)
         );
  NAND2X0_HVT U1301 ( .A1(n2270), .A2(sram_rdata_5[31]), .Y(n1183) );
  NAND3X0_HVT U1302 ( .A1(n1185), .A2(n1184), .A3(n1183), .Y(n_src_aox[175])
         );
  AO222X1_HVT U1303 ( .A1(n1860), .A2(sram_rdata_6[16]), .A3(n15500), .A4(
        sram_rdata_8[16]), .A5(sram_rdata_7[16]), .A6(n1940), .Y(n1596) );
  AOI22X1_HVT U1304 ( .A1(n1186), .A2(n10700), .A3(n5801), .A4(n1596), .Y(
        n1189) );
  OA22X1_HVT U1305 ( .A1(n10400), .A2(n525), .A3(n11500), .A4(n429), .Y(n1188)
         );
  NAND2X0_HVT U1306 ( .A1(n1750), .A2(sram_rdata_4[16]), .Y(n1187) );
  NAND3X0_HVT U1307 ( .A1(n1189), .A2(n1188), .A3(n1187), .Y(n_src_aox[176])
         );
  AO222X1_HVT U1308 ( .A1(n1840), .A2(sram_rdata_6[17]), .A3(n2110), .A4(
        sram_rdata_8[17]), .A5(sram_rdata_7[17]), .A6(n16500), .Y(n1601) );
  AOI22X1_HVT U1309 ( .A1(n11901), .A2(n10800), .A3(n15100), .A4(n1601), .Y(
        n1193) );
  OA22X1_HVT U1310 ( .A1(n11900), .A2(n526), .A3(n2750), .A4(n4301), .Y(n1192)
         );
  NAND2X0_HVT U1311 ( .A1(n576), .A2(sram_rdata_4[17]), .Y(n1191) );
  NAND3X0_HVT U1312 ( .A1(n1193), .A2(n1192), .A3(n1191), .Y(n_src_aox[177])
         );
  AO222X1_HVT U1313 ( .A1(n1880), .A2(sram_rdata_6[18]), .A3(n2130), .A4(
        sram_rdata_8[18]), .A5(sram_rdata_7[18]), .A6(n2010), .Y(n1606) );
  AOI22X1_HVT U1314 ( .A1(n1194), .A2(n588), .A3(n5801), .A4(n1606), .Y(n1197)
         );
  OA22X1_HVT U1315 ( .A1(n10300), .A2(n527), .A3(n14800), .A4(n431), .Y(n1196)
         );
  NAND2X0_HVT U1316 ( .A1(n2260), .A2(sram_rdata_4[18]), .Y(n1195) );
  NAND3X0_HVT U1317 ( .A1(n1197), .A2(n1196), .A3(n1195), .Y(n_src_aox[178])
         );
  AO222X1_HVT U1318 ( .A1(n2100), .A2(sram_rdata_6[19]), .A3(n2120), .A4(
        sram_rdata_8[19]), .A5(sram_rdata_7[19]), .A6(n1970), .Y(n1608) );
  AOI22X1_HVT U1319 ( .A1(n1198), .A2(n588), .A3(n579), .A4(n1608), .Y(n1201)
         );
  OA22X1_HVT U1320 ( .A1(n2780), .A2(n528), .A3(n11500), .A4(n432), .Y(n12001)
         );
  NAND2X0_HVT U1321 ( .A1(n2280), .A2(sram_rdata_4[19]), .Y(n1199) );
  NAND3X0_HVT U1322 ( .A1(n1201), .A2(n12001), .A3(n1199), .Y(n_src_aox[179])
         );
  AO222X1_HVT U1323 ( .A1(n12500), .A2(sram_rdata_6[20]), .A3(n15700), .A4(
        sram_rdata_8[20]), .A5(sram_rdata_7[20]), .A6(n2020), .Y(n16101) );
  AOI22X1_HVT U1324 ( .A1(n1202), .A2(n589), .A3(n5801), .A4(n16101), .Y(n1205) );
  OA22X1_HVT U1325 ( .A1(n2810), .A2(n529), .A3(n2700), .A4(n433), .Y(n1204)
         );
  NAND2X0_HVT U1326 ( .A1(n1740), .A2(sram_rdata_4[20]), .Y(n1203) );
  NAND3X0_HVT U1327 ( .A1(n1205), .A2(n1204), .A3(n1203), .Y(n_src_aox[180])
         );
  AO222X1_HVT U1328 ( .A1(n2040), .A2(sram_rdata_6[21]), .A3(n16100), .A4(
        sram_rdata_8[21]), .A5(sram_rdata_7[21]), .A6(n1960), .Y(n1612) );
  AOI22X1_HVT U1329 ( .A1(n1206), .A2(n15000), .A3(n10900), .A4(n1612), .Y(
        n1209) );
  OA22X1_HVT U1330 ( .A1(n13700), .A2(n5301), .A3(n2720), .A4(n434), .Y(n1208)
         );
  NAND2X0_HVT U1331 ( .A1(n2240), .A2(sram_rdata_4[21]), .Y(n1207) );
  NAND3X0_HVT U1332 ( .A1(n1209), .A2(n1208), .A3(n1207), .Y(n_src_aox[181])
         );
  AO222X1_HVT U1333 ( .A1(n12500), .A2(sram_rdata_6[22]), .A3(n15500), .A4(
        sram_rdata_8[22]), .A5(sram_rdata_7[22]), .A6(n1920), .Y(n1617) );
  AOI22X1_HVT U1334 ( .A1(n12101), .A2(n14900), .A3(n5801), .A4(n1617), .Y(
        n1213) );
  OA22X1_HVT U1335 ( .A1(n10600), .A2(n531), .A3(n1661), .A4(n435), .Y(n1212)
         );
  NAND2X0_HVT U1336 ( .A1(n1790), .A2(sram_rdata_4[22]), .Y(n1211) );
  NAND3X0_HVT U1337 ( .A1(n1213), .A2(n1212), .A3(n1211), .Y(n_src_aox[182])
         );
  AO222X1_HVT U1338 ( .A1(n2040), .A2(sram_rdata_6[23]), .A3(n2170), .A4(
        sram_rdata_8[23]), .A5(sram_rdata_7[23]), .A6(n1700), .Y(n1622) );
  AOI22X1_HVT U1339 ( .A1(n1214), .A2(n10800), .A3(n12900), .A4(n1622), .Y(
        n1217) );
  OA22X1_HVT U1340 ( .A1(n1662), .A2(n532), .A3(n14600), .A4(n436), .Y(n1216)
         );
  NAND2X0_HVT U1341 ( .A1(n1730), .A2(sram_rdata_4[23]), .Y(n1215) );
  NAND3X0_HVT U1342 ( .A1(n1217), .A2(n1216), .A3(n1215), .Y(n_src_aox[183])
         );
  AO222X1_HVT U1343 ( .A1(n1659), .A2(sram_rdata_6[24]), .A3(n1658), .A4(
        sram_rdata_8[24]), .A5(sram_rdata_7[24]), .A6(n1940), .Y(n1624) );
  AOI22X1_HVT U1344 ( .A1(n1218), .A2(n14900), .A3(n15100), .A4(n1624), .Y(
        n1221) );
  OA22X1_HVT U1345 ( .A1(n13800), .A2(n533), .A3(n14500), .A4(n437), .Y(n12201) );
  NAND2X0_HVT U1346 ( .A1(n1800), .A2(sram_rdata_4[24]), .Y(n1219) );
  NAND3X0_HVT U1347 ( .A1(n1221), .A2(n12201), .A3(n1219), .Y(n_src_aox[184])
         );
  AO222X1_HVT U1348 ( .A1(n1860), .A2(sram_rdata_6[25]), .A3(n15600), .A4(
        sram_rdata_8[25]), .A5(sram_rdata_7[25]), .A6(n1670), .Y(n1626) );
  AOI22X1_HVT U1349 ( .A1(n1222), .A2(n12800), .A3(n579), .A4(n1626), .Y(n1225) );
  OA22X1_HVT U1350 ( .A1(n13800), .A2(n534), .A3(n2750), .A4(n438), .Y(n1224)
         );
  NAND2X0_HVT U1351 ( .A1(n1820), .A2(sram_rdata_4[25]), .Y(n1223) );
  NAND3X0_HVT U1352 ( .A1(n1225), .A2(n1224), .A3(n1223), .Y(n_src_aox[185])
         );
  AO222X1_HVT U1353 ( .A1(n1910), .A2(sram_rdata_6[26]), .A3(n15800), .A4(
        sram_rdata_8[26]), .A5(sram_rdata_7[26]), .A6(n1930), .Y(n1628) );
  AO222X1_HVT U1354 ( .A1(n12500), .A2(sram_rdata_6[27]), .A3(n15500), .A4(
        sram_rdata_8[27]), .A5(sram_rdata_7[27]), .A6(n1690), .Y(n16301) );
  AOI22X1_HVT U1355 ( .A1(n1227), .A2(n15000), .A3(n15200), .A4(n16301), .Y(
        n12301) );
  OA22X1_HVT U1356 ( .A1(n11800), .A2(n536), .A3(n10000), .A4(n4401), .Y(n1229) );
  NAND2X0_HVT U1357 ( .A1(n2210), .A2(sram_rdata_4[27]), .Y(n1228) );
  NAND3X0_HVT U1358 ( .A1(n12301), .A2(n1229), .A3(n1228), .Y(n_src_aox[187])
         );
  AO222X1_HVT U1359 ( .A1(n2100), .A2(sram_rdata_6[28]), .A3(n16000), .A4(
        sram_rdata_8[28]), .A5(sram_rdata_7[28]), .A6(n1690), .Y(n1632) );
  AOI22X1_HVT U1360 ( .A1(n1231), .A2(n591), .A3(n15100), .A4(n1632), .Y(n1234) );
  OA22X1_HVT U1361 ( .A1(n10500), .A2(n537), .A3(n14600), .A4(n441), .Y(n1233)
         );
  NAND2X0_HVT U1362 ( .A1(n2220), .A2(sram_rdata_4[28]), .Y(n1232) );
  NAND3X0_HVT U1363 ( .A1(n1234), .A2(n1233), .A3(n1232), .Y(n_src_aox[188])
         );
  AO222X1_HVT U1364 ( .A1(n2070), .A2(sram_rdata_6[29]), .A3(n2140), .A4(
        sram_rdata_8[29]), .A5(sram_rdata_7[29]), .A6(n16400), .Y(n1637) );
  AO222X1_HVT U1365 ( .A1(n1850), .A2(sram_rdata_6[30]), .A3(n1658), .A4(
        sram_rdata_8[30]), .A5(sram_rdata_7[30]), .A6(n1690), .Y(n1642) );
  AOI22X1_HVT U1366 ( .A1(n1236), .A2(n589), .A3(n15200), .A4(n1642), .Y(n1239) );
  OA22X1_HVT U1367 ( .A1(n2770), .A2(n539), .A3(n1661), .A4(n443), .Y(n1238)
         );
  NAND2X0_HVT U1368 ( .A1(n1770), .A2(sram_rdata_4[30]), .Y(n1237) );
  NAND3X0_HVT U1369 ( .A1(n1239), .A2(n1238), .A3(n1237), .Y(n_src_aox[190])
         );
  AO222X1_HVT U1370 ( .A1(n2090), .A2(sram_rdata_6[31]), .A3(n13500), .A4(
        sram_rdata_8[31]), .A5(sram_rdata_7[31]), .A6(n16500), .Y(n1647) );
  AOI22X1_HVT U1371 ( .A1(n12401), .A2(n591), .A3(n12900), .A4(n1647), .Y(
        n1243) );
  OA22X1_HVT U1372 ( .A1(n12100), .A2(n5401), .A3(n2700), .A4(n444), .Y(n1242)
         );
  NAND2X0_HVT U1373 ( .A1(n2210), .A2(sram_rdata_4[31]), .Y(n1241) );
  NAND3X0_HVT U1374 ( .A1(n1243), .A2(n1242), .A3(n1241), .Y(n_src_aox[191])
         );
  AOI22X1_HVT U1375 ( .A1(n1245), .A2(n589), .A3(n10900), .A4(n1244), .Y(n1248) );
  OA22X1_HVT U1376 ( .A1(n12000), .A2(n350), .A3(n2750), .A4(n541), .Y(n1247)
         );
  NAND2X0_HVT U1377 ( .A1(n575), .A2(sram_rdata_0[0]), .Y(n1246) );
  NAND3X0_HVT U1378 ( .A1(n1248), .A2(n1247), .A3(n1246), .Y(n_src_aox[192])
         );
  AOI22X1_HVT U1379 ( .A1(n12501), .A2(n581), .A3(n592), .A4(n1249), .Y(n1253)
         );
  OA22X1_HVT U1380 ( .A1(n11900), .A2(n351), .A3(n2730), .A4(n542), .Y(n1252)
         );
  NAND2X0_HVT U1381 ( .A1(n2280), .A2(sram_rdata_0[1]), .Y(n1251) );
  NAND3X0_HVT U1382 ( .A1(n1253), .A2(n1252), .A3(n1251), .Y(n_src_aox[193])
         );
  AOI22X1_HVT U1383 ( .A1(n1255), .A2(n581), .A3(n12800), .A4(n1254), .Y(n1258) );
  OA22X1_HVT U1384 ( .A1(n10300), .A2(n352), .A3(n2730), .A4(n543), .Y(n1257)
         );
  NAND2X0_HVT U1385 ( .A1(n1800), .A2(sram_rdata_0[2]), .Y(n1256) );
  NAND3X0_HVT U1386 ( .A1(n1258), .A2(n1257), .A3(n1256), .Y(n_src_aox[194])
         );
  AOI22X1_HVT U1387 ( .A1(n12601), .A2(n578), .A3(n10800), .A4(n1259), .Y(
        n1263) );
  OA22X1_HVT U1388 ( .A1(n2770), .A2(n353), .A3(n2690), .A4(n544), .Y(n1262)
         );
  NAND2X0_HVT U1389 ( .A1(n2230), .A2(sram_rdata_0[3]), .Y(n1261) );
  NAND3X0_HVT U1390 ( .A1(n1263), .A2(n1262), .A3(n1261), .Y(n_src_aox[195])
         );
  AOI22X1_HVT U1391 ( .A1(n1265), .A2(n11000), .A3(n10800), .A4(n1264), .Y(
        n1268) );
  OA22X1_HVT U1392 ( .A1(n2800), .A2(n354), .A3(n10000), .A4(n545), .Y(n1267)
         );
  NAND2X0_HVT U1393 ( .A1(n1750), .A2(sram_rdata_0[4]), .Y(n1266) );
  NAND3X0_HVT U1394 ( .A1(n1268), .A2(n1267), .A3(n1266), .Y(n_src_aox[196])
         );
  AOI22X1_HVT U1395 ( .A1(n1272), .A2(n578), .A3(n12800), .A4(n1271), .Y(n1275) );
  OA22X1_HVT U1396 ( .A1(n11800), .A2(n356), .A3(n14700), .A4(n547), .Y(n1274)
         );
  NAND2X0_HVT U1397 ( .A1(n576), .A2(sram_rdata_0[6]), .Y(n1273) );
  NAND3X0_HVT U1398 ( .A1(n1275), .A2(n1274), .A3(n1273), .Y(n_src_aox[198])
         );
  AOI22X1_HVT U1399 ( .A1(n1277), .A2(n10900), .A3(n5901), .A4(n1276), .Y(
        n12801) );
  OA22X1_HVT U1400 ( .A1(n1662), .A2(n357), .A3(n2710), .A4(n548), .Y(n1279)
         );
  NAND2X0_HVT U1401 ( .A1(n1770), .A2(sram_rdata_0[7]), .Y(n1278) );
  NAND3X0_HVT U1402 ( .A1(n12801), .A2(n1279), .A3(n1278), .Y(n_src_aox[199])
         );
  AOI22X1_HVT U1403 ( .A1(n1282), .A2(n581), .A3(n592), .A4(n1281), .Y(n1285)
         );
  OA22X1_HVT U1404 ( .A1(n13700), .A2(n358), .A3(n11500), .A4(n549), .Y(n1284)
         );
  NAND2X0_HVT U1405 ( .A1(n2270), .A2(sram_rdata_0[8]), .Y(n1283) );
  NAND3X0_HVT U1406 ( .A1(n1285), .A2(n1284), .A3(n1283), .Y(n_src_aox[200])
         );
  AOI22X1_HVT U1407 ( .A1(n1287), .A2(n1648), .A3(n592), .A4(n1286), .Y(n12901) );
  OA22X1_HVT U1408 ( .A1(n2810), .A2(n359), .A3(n10100), .A4(n5501), .Y(n1289)
         );
  NAND2X0_HVT U1409 ( .A1(n2220), .A2(sram_rdata_0[9]), .Y(n1288) );
  NAND3X0_HVT U1410 ( .A1(n12901), .A2(n1289), .A3(n1288), .Y(n_src_aox[201])
         );
  AOI22X1_HVT U1411 ( .A1(n1292), .A2(n578), .A3(n10800), .A4(n1291), .Y(n1295) );
  OA22X1_HVT U1412 ( .A1(n13700), .A2(n360), .A3(n2750), .A4(n551), .Y(n1294)
         );
  NAND2X0_HVT U1413 ( .A1(n2220), .A2(sram_rdata_0[10]), .Y(n1293) );
  NAND3X0_HVT U1414 ( .A1(n1295), .A2(n1294), .A3(n1293), .Y(n_src_aox[202])
         );
  AOI22X1_HVT U1415 ( .A1(n1301), .A2(n579), .A3(n10700), .A4(n13001), .Y(
        n1304) );
  OA22X1_HVT U1416 ( .A1(n12000), .A2(n363), .A3(n2740), .A4(n554), .Y(n1303)
         );
  NAND2X0_HVT U1417 ( .A1(n1790), .A2(sram_rdata_0[13]), .Y(n1302) );
  NAND3X0_HVT U1418 ( .A1(n1304), .A2(n1303), .A3(n1302), .Y(n_src_aox[205])
         );
  AOI22X1_HVT U1419 ( .A1(n1306), .A2(n12900), .A3(n592), .A4(n1305), .Y(n1309) );
  OA22X1_HVT U1420 ( .A1(n13800), .A2(n364), .A3(n2750), .A4(n555), .Y(n1308)
         );
  NAND2X0_HVT U1421 ( .A1(n1760), .A2(sram_rdata_0[14]), .Y(n1307) );
  NAND3X0_HVT U1422 ( .A1(n1309), .A2(n1308), .A3(n1307), .Y(n_src_aox[206])
         );
  AOI22X1_HVT U1423 ( .A1(n1311), .A2(n10900), .A3(n592), .A4(n13101), .Y(
        n1314) );
  OA22X1_HVT U1424 ( .A1(n12100), .A2(n365), .A3(n10000), .A4(n556), .Y(n1313)
         );
  NAND2X0_HVT U1425 ( .A1(n2270), .A2(sram_rdata_0[15]), .Y(n1312) );
  NAND3X0_HVT U1426 ( .A1(n1314), .A2(n1313), .A3(n1312), .Y(n_src_aox[207])
         );
  AOI22X1_HVT U1427 ( .A1(n1318), .A2(n578), .A3(n12700), .A4(n1317), .Y(n1321) );
  OA22X1_HVT U1428 ( .A1(n11900), .A2(n446), .A3(n2720), .A4(n351), .Y(n13201)
         );
  NAND2X0_HVT U1429 ( .A1(n576), .A2(sram_rdata_2[1]), .Y(n1319) );
  NAND3X0_HVT U1430 ( .A1(n1321), .A2(n13201), .A3(n1319), .Y(n_src_aox[209])
         );
  AOI22X1_HVT U1431 ( .A1(n1323), .A2(n12600), .A3(n5901), .A4(n1322), .Y(
        n1326) );
  OA22X1_HVT U1432 ( .A1(n10300), .A2(n447), .A3(n2720), .A4(n352), .Y(n1325)
         );
  NAND2X0_HVT U1433 ( .A1(n2210), .A2(sram_rdata_2[2]), .Y(n1324) );
  NAND3X0_HVT U1434 ( .A1(n1326), .A2(n1325), .A3(n1324), .Y(n_src_aox[210])
         );
  AOI22X1_HVT U1435 ( .A1(n1328), .A2(n578), .A3(n592), .A4(n1327), .Y(n1331)
         );
  OA22X1_HVT U1436 ( .A1(n2770), .A2(n448), .A3(n2690), .A4(n353), .Y(n13301)
         );
  NAND2X0_HVT U1437 ( .A1(n1820), .A2(sram_rdata_2[3]), .Y(n1329) );
  NAND3X0_HVT U1438 ( .A1(n1331), .A2(n13301), .A3(n1329), .Y(n_src_aox[211])
         );
  AOI22X1_HVT U1439 ( .A1(n1333), .A2(n10900), .A3(n5901), .A4(n1332), .Y(
        n1336) );
  OA22X1_HVT U1440 ( .A1(n2810), .A2(n449), .A3(n14600), .A4(n354), .Y(n1335)
         );
  NAND2X0_HVT U1441 ( .A1(n1820), .A2(sram_rdata_2[4]), .Y(n1334) );
  NAND3X0_HVT U1442 ( .A1(n1336), .A2(n1335), .A3(n1334), .Y(n_src_aox[212])
         );
  AOI22X1_HVT U1443 ( .A1(n1338), .A2(n578), .A3(n592), .A4(n1337), .Y(n1341)
         );
  OA22X1_HVT U1444 ( .A1(n2790), .A2(n4501), .A3(n2740), .A4(n355), .Y(n13401)
         );
  NAND2X0_HVT U1445 ( .A1(n575), .A2(sram_rdata_2[5]), .Y(n1339) );
  NAND3X0_HVT U1446 ( .A1(n1341), .A2(n13401), .A3(n1339), .Y(n_src_aox[213])
         );
  AOI22X1_HVT U1447 ( .A1(n1343), .A2(n579), .A3(n10700), .A4(n1342), .Y(n1346) );
  OA22X1_HVT U1448 ( .A1(n10600), .A2(n451), .A3(n2740), .A4(n356), .Y(n1345)
         );
  NAND2X0_HVT U1449 ( .A1(n2260), .A2(sram_rdata_2[6]), .Y(n1344) );
  NAND3X0_HVT U1450 ( .A1(n1346), .A2(n1345), .A3(n1344), .Y(n_src_aox[214])
         );
  AOI22X1_HVT U1451 ( .A1(n13501), .A2(n581), .A3(n5901), .A4(n1349), .Y(n1353) );
  OA22X1_HVT U1452 ( .A1(n2790), .A2(n453), .A3(n2690), .A4(n358), .Y(n1352)
         );
  NAND2X0_HVT U1453 ( .A1(n1790), .A2(sram_rdata_2[8]), .Y(n1351) );
  NAND3X0_HVT U1454 ( .A1(n1353), .A2(n1352), .A3(n1351), .Y(n_src_aox[216])
         );
  AOI22X1_HVT U1455 ( .A1(n1355), .A2(n12600), .A3(n592), .A4(n1354), .Y(n1358) );
  OA22X1_HVT U1456 ( .A1(n2800), .A2(n454), .A3(n14800), .A4(n359), .Y(n1357)
         );
  NAND2X0_HVT U1457 ( .A1(n2240), .A2(sram_rdata_2[9]), .Y(n1356) );
  NAND3X0_HVT U1458 ( .A1(n1358), .A2(n1357), .A3(n1356), .Y(n_src_aox[217])
         );
  AOI22X1_HVT U1459 ( .A1(n13601), .A2(n581), .A3(n592), .A4(n1359), .Y(n1363)
         );
  OA22X1_HVT U1460 ( .A1(n2760), .A2(n455), .A3(n14800), .A4(n360), .Y(n1362)
         );
  NAND2X0_HVT U1461 ( .A1(n2240), .A2(sram_rdata_2[10]), .Y(n1361) );
  NAND3X0_HVT U1462 ( .A1(n1363), .A2(n1362), .A3(n1361), .Y(n_src_aox[218])
         );
  AOI22X1_HVT U1463 ( .A1(n1365), .A2(n10900), .A3(n5901), .A4(n1364), .Y(
        n1368) );
  OA22X1_HVT U1464 ( .A1(n11800), .A2(n456), .A3(n2700), .A4(n361), .Y(n1367)
         );
  NAND2X0_HVT U1465 ( .A1(n574), .A2(sram_rdata_2[11]), .Y(n1366) );
  NAND3X0_HVT U1466 ( .A1(n1368), .A2(n1367), .A3(n1366), .Y(n_src_aox[219])
         );
  AOI22X1_HVT U1467 ( .A1(n13701), .A2(n12600), .A3(n592), .A4(n1369), .Y(
        n1373) );
  OA22X1_HVT U1468 ( .A1(n11900), .A2(n457), .A3(n11500), .A4(n362), .Y(n1372)
         );
  NAND2X0_HVT U1469 ( .A1(n1810), .A2(sram_rdata_2[12]), .Y(n1371) );
  NAND3X0_HVT U1470 ( .A1(n1373), .A2(n1372), .A3(n1371), .Y(n_src_aox[220])
         );
  AOI22X1_HVT U1471 ( .A1(n1375), .A2(n581), .A3(n10800), .A4(n1374), .Y(n1378) );
  OA22X1_HVT U1472 ( .A1(n10400), .A2(n458), .A3(n1661), .A4(n363), .Y(n1377)
         );
  NAND2X0_HVT U1473 ( .A1(n574), .A2(sram_rdata_2[13]), .Y(n1376) );
  NAND3X0_HVT U1474 ( .A1(n1378), .A2(n1377), .A3(n1376), .Y(n_src_aox[221])
         );
  AOI22X1_HVT U1475 ( .A1(n13801), .A2(n582), .A3(n10700), .A4(n1379), .Y(
        n1383) );
  OA22X1_HVT U1476 ( .A1(n2780), .A2(n459), .A3(n14700), .A4(n364), .Y(n1382)
         );
  NAND2X0_HVT U1477 ( .A1(n2250), .A2(sram_rdata_2[14]), .Y(n1381) );
  NAND3X0_HVT U1478 ( .A1(n1383), .A2(n1382), .A3(n1381), .Y(n_src_aox[222])
         );
  AOI22X1_HVT U1479 ( .A1(n1385), .A2(n11000), .A3(n5901), .A4(n1384), .Y(
        n1388) );
  OA22X1_HVT U1480 ( .A1(n12100), .A2(n4601), .A3(n14500), .A4(n365), .Y(n1387) );
  NAND2X0_HVT U1481 ( .A1(n1760), .A2(sram_rdata_2[15]), .Y(n1386) );
  NAND3X0_HVT U1482 ( .A1(n1388), .A2(n1387), .A3(n1386), .Y(n_src_aox[223])
         );
  AOI22X1_HVT U1483 ( .A1(n1392), .A2(n10900), .A3(n5901), .A4(n1391), .Y(
        n1395) );
  OA22X1_HVT U1484 ( .A1(n10500), .A2(n542), .A3(n14700), .A4(n446), .Y(n1394)
         );
  NAND2X0_HVT U1485 ( .A1(n1810), .A2(sram_rdata_1[1]), .Y(n1393) );
  NAND3X0_HVT U1486 ( .A1(n1395), .A2(n1394), .A3(n1393), .Y(n_src_aox[225])
         );
  AOI22X1_HVT U1487 ( .A1(n1397), .A2(n12900), .A3(n10700), .A4(n1396), .Y(
        n14001) );
  OA22X1_HVT U1488 ( .A1(n12100), .A2(n543), .A3(n10100), .A4(n447), .Y(n1399)
         );
  NAND2X0_HVT U1489 ( .A1(n1740), .A2(sram_rdata_1[2]), .Y(n1398) );
  NAND3X0_HVT U1490 ( .A1(n14001), .A2(n1399), .A3(n1398), .Y(n_src_aox[226])
         );
  AOI22X1_HVT U1491 ( .A1(n1402), .A2(n578), .A3(n12700), .A4(n1401), .Y(n1405) );
  OA22X1_HVT U1492 ( .A1(n2780), .A2(n544), .A3(n14600), .A4(n448), .Y(n1404)
         );
  NAND2X0_HVT U1493 ( .A1(n2230), .A2(sram_rdata_1[3]), .Y(n1403) );
  NAND3X0_HVT U1494 ( .A1(n1405), .A2(n1404), .A3(n1403), .Y(n_src_aox[227])
         );
  AOI22X1_HVT U1495 ( .A1(n1407), .A2(n10900), .A3(n12700), .A4(n1406), .Y(
        n14101) );
  OA22X1_HVT U1496 ( .A1(n2800), .A2(n545), .A3(n2710), .A4(n449), .Y(n1409)
         );
  NAND2X0_HVT U1497 ( .A1(n1730), .A2(sram_rdata_1[4]), .Y(n1408) );
  NAND3X0_HVT U1498 ( .A1(n14101), .A2(n1409), .A3(n1408), .Y(n_src_aox[228])
         );
  AOI22X1_HVT U1499 ( .A1(n1412), .A2(n578), .A3(n10700), .A4(n1411), .Y(n1415) );
  OA22X1_HVT U1500 ( .A1(n13700), .A2(n546), .A3(n2740), .A4(n4501), .Y(n1414)
         );
  NAND2X0_HVT U1501 ( .A1(n2280), .A2(sram_rdata_1[5]), .Y(n1413) );
  NAND3X0_HVT U1502 ( .A1(n1415), .A2(n1414), .A3(n1413), .Y(n_src_aox[229])
         );
  AOI22X1_HVT U1503 ( .A1(n1419), .A2(n578), .A3(n592), .A4(n1418), .Y(n1422)
         );
  OA22X1_HVT U1504 ( .A1(n13700), .A2(n548), .A3(n11500), .A4(n452), .Y(n1421)
         );
  NAND2X0_HVT U1505 ( .A1(n2230), .A2(sram_rdata_1[7]), .Y(n14201) );
  NAND3X0_HVT U1506 ( .A1(n1422), .A2(n1421), .A3(n14201), .Y(n_src_aox[231])
         );
  AOI22X1_HVT U1507 ( .A1(n1424), .A2(n578), .A3(n12800), .A4(n1423), .Y(n1427) );
  OA22X1_HVT U1508 ( .A1(n13800), .A2(n549), .A3(n14600), .A4(n453), .Y(n1426)
         );
  NAND2X0_HVT U1509 ( .A1(n1730), .A2(sram_rdata_1[8]), .Y(n1425) );
  NAND3X0_HVT U1510 ( .A1(n1427), .A2(n1426), .A3(n1425), .Y(n_src_aox[232])
         );
  AOI22X1_HVT U1511 ( .A1(n1429), .A2(n581), .A3(n5901), .A4(n1428), .Y(n1432)
         );
  OA22X1_HVT U1512 ( .A1(n2810), .A2(n5501), .A3(n2740), .A4(n454), .Y(n1431)
         );
  NAND2X0_HVT U1513 ( .A1(n1750), .A2(sram_rdata_1[9]), .Y(n14301) );
  NAND3X0_HVT U1514 ( .A1(n1432), .A2(n1431), .A3(n14301), .Y(n_src_aox[233])
         );
  AOI22X1_HVT U1515 ( .A1(n1434), .A2(n11000), .A3(n12700), .A4(n1433), .Y(
        n1437) );
  OA22X1_HVT U1516 ( .A1(n2760), .A2(n551), .A3(n14800), .A4(n455), .Y(n1436)
         );
  NAND2X0_HVT U1517 ( .A1(n1720), .A2(sram_rdata_1[10]), .Y(n1435) );
  NAND3X0_HVT U1518 ( .A1(n1437), .A2(n1436), .A3(n1435), .Y(n_src_aox[234])
         );
  AOI22X1_HVT U1519 ( .A1(n1439), .A2(n12600), .A3(n5901), .A4(n1438), .Y(
        n1442) );
  OA22X1_HVT U1520 ( .A1(n10600), .A2(n552), .A3(n2690), .A4(n456), .Y(n1441)
         );
  NAND2X0_HVT U1521 ( .A1(n1740), .A2(sram_rdata_1[11]), .Y(n14401) );
  NAND3X0_HVT U1522 ( .A1(n1442), .A2(n1441), .A3(n14401), .Y(n_src_aox[235])
         );
  AOI22X1_HVT U1523 ( .A1(n1444), .A2(n578), .A3(n592), .A4(n1443), .Y(n1447)
         );
  OA22X1_HVT U1524 ( .A1(n11900), .A2(n553), .A3(n2700), .A4(n457), .Y(n1446)
         );
  NAND2X0_HVT U1525 ( .A1(n2250), .A2(sram_rdata_1[12]), .Y(n1445) );
  NAND3X0_HVT U1526 ( .A1(n1447), .A2(n1446), .A3(n1445), .Y(n_src_aox[236])
         );
  AOI22X1_HVT U1527 ( .A1(n1449), .A2(n581), .A3(n5901), .A4(n1448), .Y(n1452)
         );
  OA22X1_HVT U1528 ( .A1(n10400), .A2(n554), .A3(n2720), .A4(n458), .Y(n1451)
         );
  NAND2X0_HVT U1529 ( .A1(n1770), .A2(sram_rdata_1[13]), .Y(n14501) );
  NAND3X0_HVT U1530 ( .A1(n1452), .A2(n1451), .A3(n14501), .Y(n_src_aox[237])
         );
  AOI22X1_HVT U1531 ( .A1(n1456), .A2(n578), .A3(n5901), .A4(n1455), .Y(n1459)
         );
  OA22X1_HVT U1532 ( .A1(n10300), .A2(n556), .A3(n14500), .A4(n4601), .Y(n1458) );
  NAND2X0_HVT U1533 ( .A1(n1730), .A2(sram_rdata_1[15]), .Y(n1457) );
  NAND3X0_HVT U1534 ( .A1(n1459), .A2(n1458), .A3(n1457), .Y(n_src_aox[239])
         );
  AOI22X1_HVT U1535 ( .A1(n1461), .A2(n581), .A3(n10800), .A4(n14601), .Y(
        n1464) );
  OA22X1_HVT U1536 ( .A1(n12000), .A2(n366), .A3(n10000), .A4(n557), .Y(n1463)
         );
  NAND2X0_HVT U1537 ( .A1(n1740), .A2(sram_rdata_0[16]), .Y(n1462) );
  NAND3X0_HVT U1538 ( .A1(n1464), .A2(n1463), .A3(n1462), .Y(n_src_aox[240])
         );
  AOI22X1_HVT U1539 ( .A1(n1466), .A2(n578), .A3(n5901), .A4(n1465), .Y(n1469)
         );
  OA22X1_HVT U1540 ( .A1(n10500), .A2(n367), .A3(n1661), .A4(n558), .Y(n1468)
         );
  NAND2X0_HVT U1541 ( .A1(n1820), .A2(sram_rdata_0[17]), .Y(n1467) );
  NAND3X0_HVT U1542 ( .A1(n1469), .A2(n1468), .A3(n1467), .Y(n_src_aox[241])
         );
  AOI22X1_HVT U1543 ( .A1(n1471), .A2(n12900), .A3(n5901), .A4(n14701), .Y(
        n1474) );
  OA22X1_HVT U1544 ( .A1(n12100), .A2(n368), .A3(n14700), .A4(n559), .Y(n1473)
         );
  NAND2X0_HVT U1545 ( .A1(n1820), .A2(sram_rdata_0[18]), .Y(n1472) );
  NAND3X0_HVT U1546 ( .A1(n1474), .A2(n1473), .A3(n1472), .Y(n_src_aox[242])
         );
  AOI22X1_HVT U1547 ( .A1(n1476), .A2(n578), .A3(n12800), .A4(n1475), .Y(n1479) );
  OA22X1_HVT U1548 ( .A1(n2770), .A2(n369), .A3(n11500), .A4(n5601), .Y(n1478)
         );
  NAND2X0_HVT U1549 ( .A1(n2270), .A2(sram_rdata_0[19]), .Y(n1477) );
  NAND3X0_HVT U1550 ( .A1(n1479), .A2(n1478), .A3(n1477), .Y(n_src_aox[243])
         );
  AOI22X1_HVT U1551 ( .A1(n1481), .A2(n11000), .A3(n5901), .A4(n14801), .Y(
        n1484) );
  OA22X1_HVT U1552 ( .A1(n2800), .A2(n370), .A3(n2690), .A4(n561), .Y(n1483)
         );
  NAND2X0_HVT U1553 ( .A1(n2260), .A2(sram_rdata_0[20]), .Y(n1482) );
  NAND3X0_HVT U1554 ( .A1(n1484), .A2(n1483), .A3(n1482), .Y(n_src_aox[244])
         );
  AOI22X1_HVT U1555 ( .A1(n1486), .A2(n578), .A3(n10700), .A4(n1485), .Y(n1489) );
  OA22X1_HVT U1556 ( .A1(n13800), .A2(n371), .A3(n2730), .A4(n562), .Y(n1488)
         );
  NAND2X0_HVT U1557 ( .A1(n1730), .A2(sram_rdata_0[21]), .Y(n1487) );
  NAND3X0_HVT U1558 ( .A1(n1489), .A2(n1488), .A3(n1487), .Y(n_src_aox[245])
         );
  AOI22X1_HVT U1559 ( .A1(n1491), .A2(n578), .A3(n12700), .A4(n14901), .Y(
        n1494) );
  OA22X1_HVT U1560 ( .A1(n11800), .A2(n372), .A3(n2750), .A4(n563), .Y(n1493)
         );
  NAND2X0_HVT U1561 ( .A1(n2210), .A2(sram_rdata_0[22]), .Y(n1492) );
  NAND3X0_HVT U1562 ( .A1(n1494), .A2(n1493), .A3(n1492), .Y(n_src_aox[246])
         );
  AOI22X1_HVT U1563 ( .A1(n1496), .A2(n12600), .A3(n592), .A4(n1495), .Y(n1499) );
  OA22X1_HVT U1564 ( .A1(n2760), .A2(n373), .A3(n2710), .A4(n564), .Y(n1498)
         );
  NAND2X0_HVT U1565 ( .A1(n575), .A2(sram_rdata_0[23]), .Y(n1497) );
  NAND3X0_HVT U1566 ( .A1(n1499), .A2(n1498), .A3(n1497), .Y(n_src_aox[247])
         );
  AOI22X1_HVT U1567 ( .A1(n1503), .A2(n578), .A3(n592), .A4(n1502), .Y(n1506)
         );
  OA22X1_HVT U1568 ( .A1(n2810), .A2(n375), .A3(n2730), .A4(n566), .Y(n1505)
         );
  NAND2X0_HVT U1569 ( .A1(n1740), .A2(sram_rdata_0[25]), .Y(n1504) );
  NAND3X0_HVT U1570 ( .A1(n1506), .A2(n1505), .A3(n1504), .Y(n_src_aox[249])
         );
  AOI22X1_HVT U1571 ( .A1(n1508), .A2(n15200), .A3(n12800), .A4(n1507), .Y(
        n1511) );
  OA22X1_HVT U1572 ( .A1(n2760), .A2(n376), .A3(n14700), .A4(n567), .Y(n15101)
         );
  NAND2X0_HVT U1573 ( .A1(n2260), .A2(sram_rdata_0[26]), .Y(n1509) );
  NAND3X0_HVT U1574 ( .A1(n1511), .A2(n15101), .A3(n1509), .Y(n_src_aox[250])
         );
  AOI22X1_HVT U1575 ( .A1(n1515), .A2(n11000), .A3(n10800), .A4(n1514), .Y(
        n1518) );
  OA22X1_HVT U1576 ( .A1(n10500), .A2(n378), .A3(n14500), .A4(n569), .Y(n1517)
         );
  NAND2X0_HVT U1577 ( .A1(n1790), .A2(sram_rdata_0[28]), .Y(n1516) );
  NAND3X0_HVT U1578 ( .A1(n1518), .A2(n1517), .A3(n1516), .Y(n_src_aox[252])
         );
  AOI22X1_HVT U1579 ( .A1(n15201), .A2(n578), .A3(n592), .A4(n1519), .Y(n1523)
         );
  OA22X1_HVT U1580 ( .A1(n12000), .A2(n379), .A3(n14800), .A4(n5701), .Y(n1522) );
  NAND2X0_HVT U1581 ( .A1(n2240), .A2(sram_rdata_0[29]), .Y(n1521) );
  NAND3X0_HVT U1582 ( .A1(n1523), .A2(n1522), .A3(n1521), .Y(n_src_aox[253])
         );
  AOI22X1_HVT U1583 ( .A1(n1525), .A2(n581), .A3(n10700), .A4(n1524), .Y(n1528) );
  OA22X1_HVT U1584 ( .A1(n2780), .A2(n380), .A3(n10100), .A4(n571), .Y(n1527)
         );
  NAND2X0_HVT U1585 ( .A1(n16501), .A2(sram_rdata_0[30]), .Y(n1526) );
  NAND3X0_HVT U1586 ( .A1(n1528), .A2(n1527), .A3(n1526), .Y(n_src_aox[254])
         );
  AOI22X1_HVT U1587 ( .A1(n1532), .A2(n578), .A3(n12800), .A4(n1531), .Y(n1535) );
  OA22X1_HVT U1588 ( .A1(n12000), .A2(n461), .A3(n2690), .A4(n366), .Y(n1534)
         );
  NAND2X0_HVT U1589 ( .A1(n1790), .A2(sram_rdata_2[16]), .Y(n1533) );
  NAND3X0_HVT U1590 ( .A1(n1535), .A2(n1534), .A3(n1533), .Y(n_src_aox[256])
         );
  AOI22X1_HVT U1591 ( .A1(n1537), .A2(n581), .A3(n592), .A4(n1536), .Y(n15401)
         );
  OA22X1_HVT U1592 ( .A1(n11900), .A2(n462), .A3(n2730), .A4(n367), .Y(n1539)
         );
  NAND2X0_HVT U1593 ( .A1(n575), .A2(sram_rdata_2[17]), .Y(n1538) );
  NAND3X0_HVT U1594 ( .A1(n15401), .A2(n1539), .A3(n1538), .Y(n_src_aox[257])
         );
  AOI22X1_HVT U1595 ( .A1(n1544), .A2(n581), .A3(n5901), .A4(n1543), .Y(n1547)
         );
  OA22X1_HVT U1596 ( .A1(n2780), .A2(n464), .A3(n2700), .A4(n369), .Y(n1546)
         );
  NAND2X0_HVT U1597 ( .A1(n1820), .A2(sram_rdata_2[19]), .Y(n1545) );
  NAND3X0_HVT U1598 ( .A1(n1547), .A2(n1546), .A3(n1545), .Y(n_src_aox[259])
         );
  AOI22X1_HVT U1599 ( .A1(n1549), .A2(n12900), .A3(n592), .A4(n1548), .Y(n1552) );
  OA22X1_HVT U1600 ( .A1(n2810), .A2(n465), .A3(n11500), .A4(n370), .Y(n1551)
         );
  NAND2X0_HVT U1601 ( .A1(n2220), .A2(sram_rdata_2[20]), .Y(n15501) );
  NAND3X0_HVT U1602 ( .A1(n1552), .A2(n1551), .A3(n15501), .Y(n_src_aox[260])
         );
  AOI22X1_HVT U1603 ( .A1(n1554), .A2(n10900), .A3(n5901), .A4(n1553), .Y(
        n1557) );
  OA22X1_HVT U1604 ( .A1(n13800), .A2(n466), .A3(n10100), .A4(n371), .Y(n1556)
         );
  NAND2X0_HVT U1605 ( .A1(n1820), .A2(sram_rdata_2[21]), .Y(n1555) );
  NAND3X0_HVT U1606 ( .A1(n1557), .A2(n1556), .A3(n1555), .Y(n_src_aox[261])
         );
  AOI22X1_HVT U1607 ( .A1(n1559), .A2(n11000), .A3(n592), .A4(n1558), .Y(n1562) );
  OA22X1_HVT U1608 ( .A1(n10600), .A2(n467), .A3(n14800), .A4(n372), .Y(n1561)
         );
  NAND2X0_HVT U1609 ( .A1(n1750), .A2(sram_rdata_2[22]), .Y(n15601) );
  NAND3X0_HVT U1610 ( .A1(n1562), .A2(n1561), .A3(n15601), .Y(n_src_aox[262])
         );
  AOI22X1_HVT U1611 ( .A1(n1564), .A2(n581), .A3(n5901), .A4(n1563), .Y(n1567)
         );
  OA22X1_HVT U1612 ( .A1(n1662), .A2(n468), .A3(n2710), .A4(n373), .Y(n1566)
         );
  NAND2X0_HVT U1613 ( .A1(n2210), .A2(sram_rdata_2[23]), .Y(n1565) );
  NAND3X0_HVT U1614 ( .A1(n1567), .A2(n1566), .A3(n1565), .Y(n_src_aox[263])
         );
  AOI22X1_HVT U1615 ( .A1(n1575), .A2(n578), .A3(n5901), .A4(n1574), .Y(n1578)
         );
  OA22X1_HVT U1616 ( .A1(n10600), .A2(n472), .A3(n14600), .A4(n377), .Y(n1577)
         );
  NAND2X0_HVT U1617 ( .A1(n2230), .A2(sram_rdata_2[27]), .Y(n1576) );
  NAND3X0_HVT U1618 ( .A1(n1578), .A2(n1577), .A3(n1576), .Y(n_src_aox[267])
         );
  AOI22X1_HVT U1619 ( .A1(n15801), .A2(n12600), .A3(n5901), .A4(n1579), .Y(
        n1583) );
  OA22X1_HVT U1620 ( .A1(n10500), .A2(n473), .A3(n2700), .A4(n378), .Y(n1582)
         );
  NAND2X0_HVT U1621 ( .A1(n574), .A2(sram_rdata_2[28]), .Y(n1581) );
  NAND3X0_HVT U1622 ( .A1(n1583), .A2(n1582), .A3(n1581), .Y(n_src_aox[268])
         );
  AOI22X1_HVT U1623 ( .A1(n1585), .A2(n581), .A3(n592), .A4(n1584), .Y(n1588)
         );
  OA22X1_HVT U1624 ( .A1(n10400), .A2(n474), .A3(n2720), .A4(n379), .Y(n1587)
         );
  NAND2X0_HVT U1625 ( .A1(n1810), .A2(sram_rdata_2[29]), .Y(n1586) );
  NAND3X0_HVT U1626 ( .A1(n1588), .A2(n1587), .A3(n1586), .Y(n_src_aox[269])
         );
  AOI22X1_HVT U1627 ( .A1(n1592), .A2(n581), .A3(n592), .A4(n1591), .Y(n1595)
         );
  OA22X1_HVT U1628 ( .A1(n10300), .A2(n476), .A3(n10000), .A4(n381), .Y(n1594)
         );
  NAND2X0_HVT U1629 ( .A1(n1760), .A2(sram_rdata_2[31]), .Y(n1593) );
  NAND3X0_HVT U1630 ( .A1(n1595), .A2(n1594), .A3(n1593), .Y(n_src_aox[271])
         );
  AOI22X1_HVT U1631 ( .A1(n1597), .A2(n12600), .A3(n5901), .A4(n1596), .Y(
        n16001) );
  OA22X1_HVT U1632 ( .A1(n12000), .A2(n557), .A3(n14500), .A4(n461), .Y(n1599)
         );
  NAND2X0_HVT U1633 ( .A1(n2270), .A2(sram_rdata_1[16]), .Y(n1598) );
  NAND3X0_HVT U1634 ( .A1(n16001), .A2(n1599), .A3(n1598), .Y(n_src_aox[272])
         );
  AOI22X1_HVT U1635 ( .A1(n1602), .A2(n581), .A3(n12800), .A4(n1601), .Y(n1605) );
  OA22X1_HVT U1636 ( .A1(n11900), .A2(n558), .A3(n14800), .A4(n462), .Y(n1604)
         );
  NAND2X0_HVT U1637 ( .A1(n2220), .A2(sram_rdata_1[17]), .Y(n1603) );
  NAND3X0_HVT U1638 ( .A1(n1605), .A2(n1604), .A3(n1603), .Y(n_src_aox[273])
         );
  AOI22X1_HVT U1639 ( .A1(n1613), .A2(n10900), .A3(n592), .A4(n1612), .Y(n1616) );
  OA22X1_HVT U1640 ( .A1(n2790), .A2(n562), .A3(n14800), .A4(n466), .Y(n1615)
         );
  NAND2X0_HVT U1641 ( .A1(n1800), .A2(sram_rdata_1[21]), .Y(n1614) );
  NAND3X0_HVT U1642 ( .A1(n1616), .A2(n1615), .A3(n1614), .Y(n_src_aox[277])
         );
  AOI22X1_HVT U1643 ( .A1(n1618), .A2(n12900), .A3(n5901), .A4(n1617), .Y(
        n1621) );
  OA22X1_HVT U1644 ( .A1(n11800), .A2(n563), .A3(n2740), .A4(n467), .Y(n16201)
         );
  NAND2X0_HVT U1645 ( .A1(n1740), .A2(sram_rdata_1[22]), .Y(n1619) );
  NAND3X0_HVT U1646 ( .A1(n1621), .A2(n16201), .A3(n1619), .Y(n_src_aox[278])
         );
  AOI22X1_HVT U1647 ( .A1(n1633), .A2(n12900), .A3(n5901), .A4(n1632), .Y(
        n1636) );
  OA22X1_HVT U1648 ( .A1(n11900), .A2(n569), .A3(n11500), .A4(n473), .Y(n1635)
         );
  NAND2X0_HVT U1649 ( .A1(n1810), .A2(sram_rdata_1[28]), .Y(n1634) );
  NAND3X0_HVT U1650 ( .A1(n1636), .A2(n1635), .A3(n1634), .Y(n_src_aox[284])
         );
  AOI22X1_HVT U1651 ( .A1(n1638), .A2(n10900), .A3(n592), .A4(n1637), .Y(n1641) );
  OA22X1_HVT U1652 ( .A1(n12000), .A2(n5701), .A3(n2750), .A4(n474), .Y(n16401) );
  NAND2X0_HVT U1653 ( .A1(n1720), .A2(sram_rdata_1[29]), .Y(n1639) );
  NAND3X0_HVT U1654 ( .A1(n1641), .A2(n16401), .A3(n1639), .Y(n_src_aox[285])
         );
  AOI22X1_HVT U1655 ( .A1(n1643), .A2(n10900), .A3(n5901), .A4(n1642), .Y(
        n1646) );
  OA22X1_HVT U1656 ( .A1(n2770), .A2(n571), .A3(n14700), .A4(n475), .Y(n1645)
         );
  NAND2X0_HVT U1657 ( .A1(n2260), .A2(sram_rdata_1[30]), .Y(n1644) );
  NAND3X0_HVT U1658 ( .A1(n1646), .A2(n1645), .A3(n1644), .Y(n_src_aox[286])
         );
  AOI22X1_HVT U1659 ( .A1(n1649), .A2(n581), .A3(n592), .A4(n1647), .Y(n1653)
         );
  OA22X1_HVT U1660 ( .A1(n12100), .A2(n572), .A3(n2710), .A4(n476), .Y(n1652)
         );
  NAND2X0_HVT U1661 ( .A1(n2260), .A2(sram_rdata_1[31]), .Y(n1651) );
  NAND3X0_HVT U1662 ( .A1(n1653), .A2(n1652), .A3(n1651), .Y(n_src_aox[287])
         );
  AND2X1_HVT U1663 ( .A1(box_sel[1]), .A2(box_sel[0]), .Y(n1658) );
  AND2X1_HVT U1664 ( .A1(box_sel[0]), .A2(n1656), .Y(n1659) );
  AND2X1_HVT U1665 ( .A1(box_sel[1]), .A2(n1657), .Y(n16601) );
  AND2X1_HVT U1666 ( .A1(box_sel[3]), .A2(n1655), .Y(n1663) );
  AO22X1_HVT U1667 ( .A1(n14200), .A2(sram_rdata_b1[29]), .A3(n2340), .A4(
        sram_rdata_a1[29]), .Y(N100) );
  AO22X1_HVT U1668 ( .A1(n11600), .A2(sram_rdata_b1[30]), .A3(n2390), .A4(
        sram_rdata_a1[30]), .Y(N101) );
  AO22X1_HVT U1669 ( .A1(n2640), .A2(sram_rdata_b1[31]), .A3(n2300), .A4(
        sram_rdata_a1[31]), .Y(N102) );
  AO22X1_HVT U1670 ( .A1(n14000), .A2(sram_rdata_b2[0]), .A3(n2300), .A4(
        sram_rdata_a2[0]), .Y(N103) );
  AO22X1_HVT U1671 ( .A1(n14300), .A2(sram_rdata_b2[1]), .A3(n2320), .A4(
        sram_rdata_a2[1]), .Y(N104) );
  AO22X1_HVT U1672 ( .A1(n2670), .A2(sram_rdata_b2[2]), .A3(n2320), .A4(
        sram_rdata_a2[2]), .Y(N105) );
  AO22X1_HVT U1673 ( .A1(n14000), .A2(sram_rdata_b2[3]), .A3(n2340), .A4(
        sram_rdata_a2[3]), .Y(N106) );
  AO22X1_HVT U1674 ( .A1(n14100), .A2(sram_rdata_b2[4]), .A3(n2330), .A4(
        sram_rdata_a2[4]), .Y(N107) );
  AO22X1_HVT U1675 ( .A1(n10200), .A2(sram_rdata_b2[5]), .A3(n2290), .A4(
        sram_rdata_a2[5]), .Y(N108) );
  AO22X1_HVT U1676 ( .A1(n14200), .A2(sram_rdata_b2[6]), .A3(n2330), .A4(
        sram_rdata_a2[6]), .Y(N109) );
  AO22X1_HVT U1677 ( .A1(n11700), .A2(sram_rdata_b2[7]), .A3(n2380), .A4(
        sram_rdata_a2[7]), .Y(N110) );
  AO22X1_HVT U1678 ( .A1(n2640), .A2(sram_rdata_b2[8]), .A3(n2390), .A4(
        sram_rdata_a2[8]), .Y(N111) );
  AO22X1_HVT U1679 ( .A1(n2660), .A2(sram_rdata_b2[9]), .A3(n2340), .A4(
        sram_rdata_a2[9]), .Y(N112) );
  AO22X1_HVT U1680 ( .A1(n2660), .A2(sram_rdata_b2[10]), .A3(n2370), .A4(
        sram_rdata_a2[10]), .Y(N113) );
  AO22X1_HVT U1681 ( .A1(n2660), .A2(sram_rdata_b2[11]), .A3(n2320), .A4(
        sram_rdata_a2[11]), .Y(N114) );
  AO22X1_HVT U1682 ( .A1(n10200), .A2(sram_rdata_b2[12]), .A3(n2320), .A4(
        sram_rdata_a2[12]), .Y(N115) );
  AO22X1_HVT U1683 ( .A1(n14300), .A2(sram_rdata_b2[13]), .A3(n2390), .A4(
        sram_rdata_a2[13]), .Y(N116) );
  AO22X1_HVT U1684 ( .A1(n10200), .A2(sram_rdata_b2[14]), .A3(n2290), .A4(
        sram_rdata_a2[14]), .Y(N117) );
  AO22X1_HVT U1685 ( .A1(n2650), .A2(sram_rdata_b2[15]), .A3(n2350), .A4(
        sram_rdata_a2[15]), .Y(N118) );
  AO22X1_HVT U1686 ( .A1(n2650), .A2(sram_rdata_b2[16]), .A3(n2340), .A4(
        sram_rdata_a2[16]), .Y(N119) );
  AO22X1_HVT U1687 ( .A1(n2680), .A2(sram_rdata_b2[17]), .A3(n2290), .A4(
        sram_rdata_a2[17]), .Y(N120) );
  AO22X1_HVT U1688 ( .A1(n2680), .A2(sram_rdata_b2[18]), .A3(n2300), .A4(
        sram_rdata_a2[18]), .Y(N121) );
  AO22X1_HVT U1689 ( .A1(n10200), .A2(sram_rdata_b2[19]), .A3(n2370), .A4(
        sram_rdata_a2[19]), .Y(N122) );
  AO22X1_HVT U1690 ( .A1(n11700), .A2(sram_rdata_b2[20]), .A3(n2330), .A4(
        sram_rdata_a2[20]), .Y(N123) );
  AO22X1_HVT U1691 ( .A1(n14200), .A2(sram_rdata_b2[21]), .A3(n2350), .A4(
        sram_rdata_a2[21]), .Y(N124) );
  AO22X1_HVT U1692 ( .A1(n2660), .A2(sram_rdata_b2[22]), .A3(n2340), .A4(
        sram_rdata_a2[22]), .Y(N125) );
  AO22X1_HVT U1693 ( .A1(n14000), .A2(sram_rdata_b2[23]), .A3(n2370), .A4(
        sram_rdata_a2[23]), .Y(N126) );
  AO22X1_HVT U1694 ( .A1(n14100), .A2(sram_rdata_b2[24]), .A3(n2370), .A4(
        sram_rdata_a2[24]), .Y(N127) );
  AO22X1_HVT U1695 ( .A1(n11600), .A2(sram_rdata_b2[25]), .A3(n2370), .A4(
        sram_rdata_a2[25]), .Y(N128) );
  AO22X1_HVT U1696 ( .A1(n2670), .A2(sram_rdata_b2[26]), .A3(n2300), .A4(
        sram_rdata_a2[26]), .Y(N129) );
  AO22X1_HVT U1697 ( .A1(n2640), .A2(sram_rdata_b2[27]), .A3(n2290), .A4(
        sram_rdata_a2[27]), .Y(N130) );
  AO22X1_HVT U1698 ( .A1(n14000), .A2(sram_rdata_b2[28]), .A3(n2290), .A4(
        sram_rdata_a2[28]), .Y(N131) );
  AO22X1_HVT U1699 ( .A1(n2680), .A2(sram_rdata_b2[29]), .A3(n2340), .A4(
        sram_rdata_a2[29]), .Y(N132) );
  AO22X1_HVT U1700 ( .A1(n11600), .A2(sram_rdata_b2[30]), .A3(n2370), .A4(
        sram_rdata_a2[30]), .Y(N133) );
  AO22X1_HVT U1701 ( .A1(n14100), .A2(sram_rdata_b2[31]), .A3(n2350), .A4(
        sram_rdata_a2[31]), .Y(N134) );
  AO22X1_HVT U1702 ( .A1(n2640), .A2(sram_rdata_b3[0]), .A3(n2380), .A4(
        sram_rdata_a3[0]), .Y(N135) );
  AO22X1_HVT U1703 ( .A1(n2670), .A2(sram_rdata_b3[1]), .A3(n2310), .A4(
        sram_rdata_a3[1]), .Y(N136) );
  AO22X1_HVT U1704 ( .A1(n14300), .A2(sram_rdata_b3[2]), .A3(n2300), .A4(
        sram_rdata_a3[2]), .Y(N137) );
  AO22X1_HVT U1705 ( .A1(n2640), .A2(sram_rdata_b3[3]), .A3(n2300), .A4(
        sram_rdata_a3[3]), .Y(N138) );
  AO22X1_HVT U1706 ( .A1(n14000), .A2(sram_rdata_b3[4]), .A3(n2360), .A4(
        sram_rdata_a3[4]), .Y(N139) );
  AO22X1_HVT U1707 ( .A1(n14300), .A2(sram_rdata_b3[5]), .A3(n2330), .A4(
        sram_rdata_a3[5]), .Y(N140) );
  AO22X1_HVT U1708 ( .A1(n2670), .A2(sram_rdata_b3[6]), .A3(n2350), .A4(
        sram_rdata_a3[6]), .Y(N141) );
  AO22X1_HVT U1709 ( .A1(n11700), .A2(sram_rdata_b3[7]), .A3(n2390), .A4(
        sram_rdata_a3[7]), .Y(N142) );
  AO22X1_HVT U1710 ( .A1(n2650), .A2(sram_rdata_b3[8]), .A3(n2380), .A4(
        sram_rdata_a3[8]), .Y(N143) );
  AO22X1_HVT U1711 ( .A1(n10200), .A2(sram_rdata_b3[9]), .A3(n2330), .A4(
        sram_rdata_a3[9]), .Y(N144) );
  AO22X1_HVT U1712 ( .A1(n2680), .A2(sram_rdata_b3[10]), .A3(n2360), .A4(
        sram_rdata_a3[10]), .Y(N145) );
  AO22X1_HVT U1713 ( .A1(n2650), .A2(sram_rdata_b3[11]), .A3(n2300), .A4(
        sram_rdata_a3[11]), .Y(N146) );
  AO22X1_HVT U1714 ( .A1(n14100), .A2(sram_rdata_b3[12]), .A3(n2310), .A4(
        sram_rdata_a3[12]), .Y(N147) );
  AO22X1_HVT U1715 ( .A1(n2670), .A2(sram_rdata_b3[13]), .A3(n2380), .A4(
        sram_rdata_a3[13]), .Y(N148) );
  AO22X1_HVT U1716 ( .A1(n10200), .A2(sram_rdata_b3[14]), .A3(n2380), .A4(
        sram_rdata_a3[14]), .Y(N149) );
  AO22X1_HVT U1717 ( .A1(n14000), .A2(sram_rdata_b3[15]), .A3(n2360), .A4(
        sram_rdata_a3[15]), .Y(N150) );
  AO22X1_HVT U1718 ( .A1(n2640), .A2(sram_rdata_b3[16]), .A3(n2310), .A4(
        sram_rdata_a3[16]), .Y(N151) );
  AO22X1_HVT U1719 ( .A1(n2660), .A2(sram_rdata_b3[17]), .A3(n2310), .A4(
        sram_rdata_a3[17]), .Y(N152) );
  AO22X1_HVT U1720 ( .A1(n14200), .A2(sram_rdata_b3[18]), .A3(n2390), .A4(
        sram_rdata_a3[18]), .Y(N153) );
  AO22X1_HVT U1721 ( .A1(n2650), .A2(sram_rdata_b3[19]), .A3(n2330), .A4(
        sram_rdata_a3[19]), .Y(N154) );
  AO22X1_HVT U1722 ( .A1(n14300), .A2(sram_rdata_b3[20]), .A3(n2360), .A4(
        sram_rdata_a3[20]), .Y(N155) );
  AO22X1_HVT U1723 ( .A1(n11600), .A2(sram_rdata_b3[21]), .A3(n2310), .A4(
        sram_rdata_a3[21]), .Y(N156) );
  AO22X1_HVT U1724 ( .A1(n2680), .A2(sram_rdata_b3[22]), .A3(n2320), .A4(
        sram_rdata_a3[22]), .Y(N157) );
  AO22X1_HVT U1725 ( .A1(n14100), .A2(sram_rdata_b3[23]), .A3(n2370), .A4(
        sram_rdata_a3[23]), .Y(N158) );
  AO22X1_HVT U1726 ( .A1(n11700), .A2(sram_rdata_b3[24]), .A3(n2330), .A4(
        sram_rdata_a3[24]), .Y(N159) );
  AO22X1_HVT U1727 ( .A1(n2680), .A2(sram_rdata_b3[25]), .A3(n2330), .A4(
        sram_rdata_a3[25]), .Y(N160) );
  AO22X1_HVT U1728 ( .A1(n14300), .A2(sram_rdata_b3[26]), .A3(n2340), .A4(
        sram_rdata_a3[26]), .Y(N161) );
  AO22X1_HVT U1729 ( .A1(n14100), .A2(sram_rdata_b3[27]), .A3(n2370), .A4(
        sram_rdata_a3[27]), .Y(N162) );
  AO22X1_HVT U1730 ( .A1(n2650), .A2(sram_rdata_b3[28]), .A3(n2380), .A4(
        sram_rdata_a3[28]), .Y(N163) );
  AO22X1_HVT U1731 ( .A1(n2660), .A2(sram_rdata_b3[29]), .A3(n2310), .A4(
        sram_rdata_a3[29]), .Y(N164) );
  AO22X1_HVT U1732 ( .A1(n11600), .A2(sram_rdata_b3[30]), .A3(n2320), .A4(
        sram_rdata_a3[30]), .Y(N165) );
  AO22X1_HVT U1733 ( .A1(n14200), .A2(sram_rdata_b3[31]), .A3(n2320), .A4(
        sram_rdata_a3[31]), .Y(N166) );
  AO22X1_HVT U1734 ( .A1(n14300), .A2(sram_rdata_b4[0]), .A3(n2310), .A4(
        sram_rdata_a4[0]), .Y(N167) );
  AO22X1_HVT U1735 ( .A1(n2670), .A2(sram_rdata_b4[1]), .A3(n2330), .A4(
        sram_rdata_a4[1]), .Y(N168) );
  AO22X1_HVT U1736 ( .A1(n2660), .A2(sram_rdata_b4[2]), .A3(n2310), .A4(
        sram_rdata_a4[2]), .Y(N169) );
  AO22X1_HVT U1737 ( .A1(n14100), .A2(sram_rdata_b4[3]), .A3(n2330), .A4(
        sram_rdata_a4[3]), .Y(N170) );
  AO22X1_HVT U1738 ( .A1(n2650), .A2(sram_rdata_b4[4]), .A3(n2380), .A4(
        sram_rdata_a4[4]), .Y(N171) );
  AO22X1_HVT U1739 ( .A1(n2680), .A2(sram_rdata_b4[5]), .A3(n2290), .A4(
        sram_rdata_a4[5]), .Y(N172) );
  AO22X1_HVT U1740 ( .A1(n14300), .A2(sram_rdata_b4[6]), .A3(n2320), .A4(
        sram_rdata_a4[6]), .Y(N173) );
  AO22X1_HVT U1741 ( .A1(n14000), .A2(sram_rdata_b4[7]), .A3(n2320), .A4(
        sram_rdata_a4[7]), .Y(N174) );
  AO22X1_HVT U1742 ( .A1(n2650), .A2(sram_rdata_b4[8]), .A3(n2340), .A4(
        sram_rdata_a4[8]), .Y(N175) );
  AO22X1_HVT U1743 ( .A1(n10200), .A2(sram_rdata_b4[9]), .A3(n2350), .A4(
        sram_rdata_a4[9]), .Y(N176) );
  AO22X1_HVT U1744 ( .A1(n14200), .A2(sram_rdata_b4[10]), .A3(n2340), .A4(
        sram_rdata_a4[10]), .Y(N177) );
  AO22X1_HVT U1745 ( .A1(n11700), .A2(sram_rdata_b4[11]), .A3(n2370), .A4(
        sram_rdata_a4[11]), .Y(N178) );
  AO22X1_HVT U1746 ( .A1(n2640), .A2(sram_rdata_b4[12]), .A3(n2380), .A4(
        sram_rdata_a4[12]), .Y(N179) );
  AO22X1_HVT U1747 ( .A1(n14200), .A2(sram_rdata_b4[13]), .A3(n2360), .A4(
        sram_rdata_a4[13]), .Y(N180) );
  AO22X1_HVT U1748 ( .A1(n10200), .A2(sram_rdata_b4[14]), .A3(n2350), .A4(
        sram_rdata_a4[14]), .Y(N181) );
  AO22X1_HVT U1749 ( .A1(n2640), .A2(sram_rdata_b4[15]), .A3(n2320), .A4(
        sram_rdata_a4[15]), .Y(N182) );
  AO22X1_HVT U1750 ( .A1(n14000), .A2(sram_rdata_b4[16]), .A3(n2290), .A4(
        sram_rdata_a4[16]), .Y(N183) );
  AO22X1_HVT U1751 ( .A1(n2660), .A2(sram_rdata_b4[17]), .A3(n2370), .A4(
        sram_rdata_a4[17]), .Y(N184) );
  AO22X1_HVT U1752 ( .A1(n2670), .A2(sram_rdata_b4[18]), .A3(n2390), .A4(
        sram_rdata_a4[18]), .Y(N185) );
  AO22X1_HVT U1753 ( .A1(n14000), .A2(sram_rdata_b4[19]), .A3(n2340), .A4(
        sram_rdata_a4[19]), .Y(N186) );
  AO22X1_HVT U1754 ( .A1(n2640), .A2(sram_rdata_b4[20]), .A3(n2290), .A4(
        sram_rdata_a4[20]), .Y(N187) );
  AO22X1_HVT U1755 ( .A1(n2670), .A2(sram_rdata_b4[21]), .A3(n2290), .A4(
        sram_rdata_a4[21]), .Y(N188) );
  AO22X1_HVT U1756 ( .A1(n14200), .A2(sram_rdata_b4[22]), .A3(n2390), .A4(
        sram_rdata_a4[22]), .Y(N189) );
  AO22X1_HVT U1757 ( .A1(n2670), .A2(sram_rdata_b4[23]), .A3(n2340), .A4(
        sram_rdata_a4[23]), .Y(N190) );
  AO22X1_HVT U1758 ( .A1(n11700), .A2(sram_rdata_b4[24]), .A3(n2340), .A4(
        sram_rdata_a4[24]), .Y(N191) );
  AO22X1_HVT U1759 ( .A1(n11600), .A2(sram_rdata_b4[25]), .A3(n2300), .A4(
        sram_rdata_a4[25]), .Y(N192) );
  AO22X1_HVT U1760 ( .A1(n2660), .A2(sram_rdata_b4[26]), .A3(n2290), .A4(
        sram_rdata_a4[26]), .Y(N193) );
  AO22X1_HVT U1761 ( .A1(n14100), .A2(sram_rdata_b4[27]), .A3(n593), .A4(
        sram_rdata_a4[27]), .Y(N194) );
  AO22X1_HVT U1762 ( .A1(n2680), .A2(sram_rdata_b4[28]), .A3(n2350), .A4(
        sram_rdata_a4[28]), .Y(N195) );
  AO22X1_HVT U1763 ( .A1(n14300), .A2(sram_rdata_b4[29]), .A3(n2360), .A4(
        sram_rdata_a4[29]), .Y(N196) );
  AO22X1_HVT U1764 ( .A1(n11600), .A2(sram_rdata_b4[30]), .A3(n2360), .A4(
        sram_rdata_a4[30]), .Y(N197) );
  AO22X1_HVT U1765 ( .A1(n2650), .A2(sram_rdata_b4[31]), .A3(n2370), .A4(
        sram_rdata_a4[31]), .Y(N198) );
  AO22X1_HVT U1766 ( .A1(n14200), .A2(sram_rdata_b5[0]), .A3(n2380), .A4(
        sram_rdata_a5[0]), .Y(N199) );
  AO22X1_HVT U1767 ( .A1(n14200), .A2(sram_rdata_b5[1]), .A3(n2380), .A4(
        sram_rdata_a5[1]), .Y(N200) );
  AO22X1_HVT U1768 ( .A1(n2680), .A2(sram_rdata_b5[2]), .A3(n2310), .A4(
        sram_rdata_a5[2]), .Y(N201) );
  AO22X1_HVT U1769 ( .A1(n14300), .A2(sram_rdata_b5[3]), .A3(n2300), .A4(
        sram_rdata_a5[3]), .Y(N202) );
  AO22X1_HVT U1770 ( .A1(n14100), .A2(sram_rdata_b5[4]), .A3(n2290), .A4(
        sram_rdata_a5[4]), .Y(N203) );
  AO22X1_HVT U1771 ( .A1(n2660), .A2(sram_rdata_b5[5]), .A3(n2350), .A4(
        sram_rdata_a5[5]), .Y(N204) );
  AO22X1_HVT U1772 ( .A1(n2660), .A2(sram_rdata_b5[6]), .A3(n2390), .A4(
        sram_rdata_a5[6]), .Y(N205) );
  AO22X1_HVT U1773 ( .A1(n11700), .A2(sram_rdata_b5[7]), .A3(n2350), .A4(
        sram_rdata_a5[7]), .Y(N206) );
  AO22X1_HVT U1774 ( .A1(n10200), .A2(sram_rdata_b5[8]), .A3(n2380), .A4(
        sram_rdata_a5[8]), .Y(N207) );
  AO22X1_HVT U1775 ( .A1(n10200), .A2(sram_rdata_b5[9]), .A3(n2300), .A4(
        sram_rdata_a5[9]), .Y(N208) );
  AO22X1_HVT U1776 ( .A1(n2670), .A2(sram_rdata_b5[10]), .A3(n2310), .A4(
        sram_rdata_a5[10]), .Y(N209) );
  AO22X1_HVT U1777 ( .A1(n2640), .A2(sram_rdata_b5[11]), .A3(n2290), .A4(
        sram_rdata_a5[11]), .Y(N210) );
  AO22X1_HVT U1778 ( .A1(n14000), .A2(sram_rdata_b5[12]), .A3(n2350), .A4(
        sram_rdata_a5[12]), .Y(N211) );
  AO22X1_HVT U1779 ( .A1(n2680), .A2(sram_rdata_b5[13]), .A3(n2330), .A4(
        sram_rdata_a5[13]), .Y(N212) );
  AO22X1_HVT U1780 ( .A1(n10200), .A2(sram_rdata_b5[14]), .A3(n2360), .A4(
        sram_rdata_a5[14]), .Y(N213) );
  AO22X1_HVT U1781 ( .A1(n14100), .A2(sram_rdata_b5[15]), .A3(n2380), .A4(
        sram_rdata_a5[15]), .Y(N214) );
  AO22X1_HVT U1782 ( .A1(n11700), .A2(sram_rdata_b5[16]), .A3(n2390), .A4(
        sram_rdata_a5[16]), .Y(N215) );
  AO22X1_HVT U1783 ( .A1(n14300), .A2(sram_rdata_b5[17]), .A3(n2370), .A4(
        sram_rdata_a5[17]), .Y(N216) );
  AO22X1_HVT U1784 ( .A1(n14300), .A2(sram_rdata_b5[18]), .A3(n2330), .A4(
        sram_rdata_a5[18]), .Y(N217) );
  AO22X1_HVT U1785 ( .A1(n2640), .A2(sram_rdata_b5[19]), .A3(n2300), .A4(
        sram_rdata_a5[19]), .Y(N218) );
  AO22X1_HVT U1786 ( .A1(n2650), .A2(sram_rdata_b5[20]), .A3(n2320), .A4(
        sram_rdata_a5[20]), .Y(N219) );
  AO22X1_HVT U1787 ( .A1(n14200), .A2(sram_rdata_b5[21]), .A3(n2370), .A4(
        sram_rdata_a5[21]), .Y(N220) );
  AO22X1_HVT U1788 ( .A1(n2670), .A2(sram_rdata_b5[22]), .A3(n2370), .A4(
        sram_rdata_a5[22]), .Y(N221) );
  AO22X1_HVT U1789 ( .A1(n2650), .A2(sram_rdata_b5[23]), .A3(n2360), .A4(
        sram_rdata_a5[23]), .Y(N222) );
  AO22X1_HVT U1790 ( .A1(n14000), .A2(sram_rdata_b5[24]), .A3(n2310), .A4(
        sram_rdata_a5[24]), .Y(N223) );
  AO22X1_HVT U1791 ( .A1(n11600), .A2(sram_rdata_b5[25]), .A3(n2300), .A4(
        sram_rdata_a5[25]), .Y(N224) );
  AO22X1_HVT U1792 ( .A1(n2680), .A2(sram_rdata_b5[26]), .A3(n2380), .A4(
        sram_rdata_a5[26]), .Y(N225) );
  AO22X1_HVT U1793 ( .A1(n2650), .A2(sram_rdata_b5[27]), .A3(n2350), .A4(
        sram_rdata_a5[27]), .Y(N226) );
  AO22X1_HVT U1794 ( .A1(n14100), .A2(sram_rdata_b5[28]), .A3(n2360), .A4(
        sram_rdata_a5[28]), .Y(N227) );
  AO22X1_HVT U1795 ( .A1(n2680), .A2(sram_rdata_b5[29]), .A3(n2300), .A4(
        sram_rdata_a5[29]), .Y(N228) );
  AO22X1_HVT U1796 ( .A1(n11600), .A2(sram_rdata_b5[30]), .A3(n2310), .A4(
        sram_rdata_a5[30]), .Y(N229) );
  AO22X1_HVT U1797 ( .A1(n14000), .A2(sram_rdata_b5[31]), .A3(n2370), .A4(
        sram_rdata_a5[31]), .Y(N230) );
  AO22X1_HVT U1798 ( .A1(n14100), .A2(sram_rdata_b6[0]), .A3(n2330), .A4(
        sram_rdata_a6[0]), .Y(N231) );
  AO22X1_HVT U1799 ( .A1(n2670), .A2(sram_rdata_b6[1]), .A3(n2340), .A4(
        sram_rdata_a6[1]), .Y(N232) );
  AO22X1_HVT U1800 ( .A1(n14200), .A2(sram_rdata_b6[2]), .A3(n2340), .A4(
        sram_rdata_a6[2]), .Y(N233) );
  AO22X1_HVT U1801 ( .A1(n2650), .A2(sram_rdata_b6[3]), .A3(n593), .A4(
        sram_rdata_a6[3]), .Y(N234) );
  AO22X1_HVT U1802 ( .A1(n2650), .A2(sram_rdata_b6[4]), .A3(n2390), .A4(
        sram_rdata_a6[4]), .Y(N235) );
  AO22X1_HVT U1803 ( .A1(n14300), .A2(sram_rdata_b6[5]), .A3(n2380), .A4(
        sram_rdata_a6[5]), .Y(N236) );
  AO22X1_HVT U1804 ( .A1(n2680), .A2(sram_rdata_b6[6]), .A3(n2290), .A4(
        sram_rdata_a6[6]), .Y(N237) );
  AO22X1_HVT U1805 ( .A1(n14100), .A2(sram_rdata_b6[7]), .A3(n2300), .A4(
        sram_rdata_a6[7]), .Y(N238) );
  AO22X1_HVT U1806 ( .A1(n2640), .A2(sram_rdata_b6[8]), .A3(n2310), .A4(
        sram_rdata_a6[8]), .Y(N239) );
  AO22X1_HVT U1807 ( .A1(n10200), .A2(sram_rdata_b6[9]), .A3(n2340), .A4(
        sram_rdata_a6[9]), .Y(N240) );
  AO22X1_HVT U1808 ( .A1(n14300), .A2(sram_rdata_b6[10]), .A3(n2380), .A4(
        sram_rdata_a6[10]), .Y(N241) );
  AO22X1_HVT U1809 ( .A1(n11700), .A2(sram_rdata_b6[11]), .A3(n2360), .A4(
        sram_rdata_a6[11]), .Y(N242) );
  AO22X1_HVT U1810 ( .A1(n14100), .A2(sram_rdata_b6[12]), .A3(n2390), .A4(
        sram_rdata_a6[12]), .Y(N243) );
  AO22X1_HVT U1811 ( .A1(n2670), .A2(sram_rdata_b6[13]), .A3(n2300), .A4(
        sram_rdata_a6[13]), .Y(N244) );
  AO22X1_HVT U1812 ( .A1(n10200), .A2(sram_rdata_b6[14]), .A3(n2310), .A4(
        sram_rdata_a6[14]), .Y(N245) );
  AO22X1_HVT U1813 ( .A1(n14200), .A2(sram_rdata_b6[15]), .A3(n2300), .A4(
        sram_rdata_a6[15]), .Y(N246) );
  AO22X1_HVT U1814 ( .A1(n11700), .A2(sram_rdata_b6[16]), .A3(n2360), .A4(
        sram_rdata_a6[16]), .Y(N247) );
  AO22X1_HVT U1815 ( .A1(n2660), .A2(sram_rdata_b6[17]), .A3(n2350), .A4(
        sram_rdata_a6[17]), .Y(N248) );
  AO22X1_HVT U1816 ( .A1(n2660), .A2(sram_rdata_b6[18]), .A3(n2350), .A4(
        sram_rdata_a6[18]), .Y(N249) );
  AO22X1_HVT U1817 ( .A1(n14100), .A2(sram_rdata_b6[19]), .A3(n2390), .A4(
        sram_rdata_a6[19]), .Y(N250) );
  AO22X1_HVT U1818 ( .A1(n2640), .A2(sram_rdata_b6[20]), .A3(n593), .A4(
        sram_rdata_a6[20]), .Y(N251) );
  AO22X1_HVT U1819 ( .A1(n2680), .A2(sram_rdata_b6[21]), .A3(n2370), .A4(
        sram_rdata_a6[21]), .Y(N252) );
  AO22X1_HVT U1820 ( .A1(n14300), .A2(sram_rdata_b6[22]), .A3(n2350), .A4(
        sram_rdata_a6[22]), .Y(N253) );
  AO22X1_HVT U1821 ( .A1(n14000), .A2(sram_rdata_b6[23]), .A3(n2310), .A4(
        sram_rdata_a6[23]), .Y(N254) );
  AO22X1_HVT U1822 ( .A1(n2660), .A2(sram_rdata_b6[24]), .A3(n2310), .A4(
        sram_rdata_a6[24]), .Y(N255) );
  AO22X1_HVT U1823 ( .A1(n11600), .A2(sram_rdata_b6[25]), .A3(n2380), .A4(
        sram_rdata_a6[25]), .Y(N256) );
  AO22X1_HVT U1824 ( .A1(n14200), .A2(sram_rdata_b6[26]), .A3(n2330), .A4(
        sram_rdata_a6[26]), .Y(N257) );
  AO22X1_HVT U1825 ( .A1(n14000), .A2(sram_rdata_b6[27]), .A3(n2360), .A4(
        sram_rdata_a6[27]), .Y(N258) );
  AO22X1_HVT U1826 ( .A1(n2650), .A2(sram_rdata_b6[28]), .A3(n2320), .A4(
        sram_rdata_a6[28]), .Y(N259) );
  AO22X1_HVT U1827 ( .A1(n2660), .A2(sram_rdata_b6[29]), .A3(n2320), .A4(
        sram_rdata_a6[29]), .Y(N260) );
  AO22X1_HVT U1828 ( .A1(n11600), .A2(sram_rdata_b6[30]), .A3(n2380), .A4(
        sram_rdata_a6[30]), .Y(N261) );
  AO22X1_HVT U1829 ( .A1(n2640), .A2(sram_rdata_b6[31]), .A3(n2330), .A4(
        sram_rdata_a6[31]), .Y(N262) );
  AO22X1_HVT U1830 ( .A1(n2820), .A2(sram_rdata_b7[0]), .A3(n2330), .A4(
        sram_rdata_a7[0]), .Y(N263) );
  AO22X1_HVT U1831 ( .A1(n14200), .A2(sram_rdata_b7[1]), .A3(n2320), .A4(
        sram_rdata_a7[1]), .Y(N264) );
  AO22X1_HVT U1832 ( .A1(n2670), .A2(sram_rdata_b7[2]), .A3(n2320), .A4(
        sram_rdata_a7[2]), .Y(N265) );
  AO22X1_HVT U1833 ( .A1(n14000), .A2(sram_rdata_b7[3]), .A3(n2380), .A4(
        sram_rdata_a7[3]), .Y(N266) );
  AO22X1_HVT U1834 ( .A1(n2670), .A2(sram_rdata_b7[4]), .A3(n2330), .A4(
        sram_rdata_a7[4]), .Y(N267) );
  AO22X1_HVT U1835 ( .A1(n2670), .A2(sram_rdata_b7[5]), .A3(n2360), .A4(
        sram_rdata_a7[5]), .Y(N268) );
  AO22X1_HVT U1836 ( .A1(n14200), .A2(sram_rdata_b7[6]), .A3(n2360), .A4(
        sram_rdata_a7[6]), .Y(N269) );
  AO22X1_HVT U1837 ( .A1(n11700), .A2(sram_rdata_b7[7]), .A3(n2380), .A4(
        sram_rdata_a7[7]), .Y(N270) );
  AO22X1_HVT U1838 ( .A1(n14000), .A2(sram_rdata_b7[8]), .A3(n2370), .A4(
        sram_rdata_a7[8]), .Y(N271) );
  AO22X1_HVT U1839 ( .A1(n10200), .A2(sram_rdata_b7[9]), .A3(n2300), .A4(
        sram_rdata_a7[9]), .Y(N272) );
  AO22X1_HVT U1840 ( .A1(n2660), .A2(sram_rdata_b7[10]), .A3(n2310), .A4(
        sram_rdata_a7[10]), .Y(N273) );
  AO22X1_HVT U1841 ( .A1(n2680), .A2(sram_rdata_b7[11]), .A3(n2310), .A4(
        sram_rdata_a7[11]), .Y(N274) );
  AO22X1_HVT U1842 ( .A1(n2640), .A2(sram_rdata_b7[12]), .A3(n2320), .A4(
        sram_rdata_a7[12]), .Y(N275) );
  AO22X1_HVT U1843 ( .A1(n14200), .A2(sram_rdata_b7[13]), .A3(n2340), .A4(
        sram_rdata_a7[13]), .Y(N276) );
  AO22X1_HVT U1844 ( .A1(n10200), .A2(sram_rdata_b7[14]), .A3(n2300), .A4(
        sram_rdata_a7[14]), .Y(N277) );
  AO22X1_HVT U1845 ( .A1(n2650), .A2(sram_rdata_b7[15]), .A3(n2340), .A4(
        sram_rdata_a7[15]), .Y(N278) );
  AO22X1_HVT U1846 ( .A1(n11700), .A2(sram_rdata_b7[16]), .A3(n2390), .A4(
        sram_rdata_a7[16]), .Y(N279) );
  AO22X1_HVT U1847 ( .A1(n14300), .A2(sram_rdata_b7[17]), .A3(n2290), .A4(
        sram_rdata_a7[17]), .Y(N280) );
  AO22X1_HVT U1848 ( .A1(n2680), .A2(sram_rdata_b7[18]), .A3(n2320), .A4(
        sram_rdata_a7[18]), .Y(N281) );
  AO22X1_HVT U1849 ( .A1(n10200), .A2(sram_rdata_b7[19]), .A3(n2290), .A4(
        sram_rdata_a7[19]), .Y(N282) );
  AO22X1_HVT U1850 ( .A1(n14000), .A2(sram_rdata_b7[20]), .A3(n2360), .A4(
        sram_rdata_a7[20]), .Y(N283) );
  AO22X1_HVT U1851 ( .A1(n2660), .A2(sram_rdata_b7[21]), .A3(n2330), .A4(
        sram_rdata_a7[21]), .Y(N284) );
  AO22X1_HVT U1852 ( .A1(n2660), .A2(sram_rdata_b7[22]), .A3(n2330), .A4(
        sram_rdata_a7[22]), .Y(N285) );
  AO22X1_HVT U1853 ( .A1(n2640), .A2(sram_rdata_b7[23]), .A3(n2380), .A4(
        sram_rdata_a7[23]), .Y(N286) );
  AO22X1_HVT U1854 ( .A1(n14100), .A2(sram_rdata_b7[24]), .A3(n593), .A4(
        sram_rdata_a7[24]), .Y(N287) );
  AO22X1_HVT U1855 ( .A1(n11600), .A2(sram_rdata_b7[25]), .A3(n2370), .A4(
        sram_rdata_a7[25]), .Y(N288) );
  AO22X1_HVT U1856 ( .A1(n2670), .A2(sram_rdata_b7[26]), .A3(n2340), .A4(
        sram_rdata_a7[26]), .Y(N289) );
  AO22X1_HVT U1857 ( .A1(n2640), .A2(sram_rdata_b7[27]), .A3(n2320), .A4(
        sram_rdata_a7[27]), .Y(N290) );
  AO22X1_HVT U1858 ( .A1(n10200), .A2(sram_rdata_b7[28]), .A3(n2300), .A4(
        sram_rdata_a7[28]), .Y(N291) );
  AO22X1_HVT U1859 ( .A1(n14300), .A2(sram_rdata_b7[29]), .A3(n2290), .A4(
        sram_rdata_a7[29]), .Y(N292) );
  AO22X1_HVT U1860 ( .A1(n11600), .A2(sram_rdata_b7[30]), .A3(n2390), .A4(
        sram_rdata_a7[30]), .Y(N293) );
  AO22X1_HVT U1861 ( .A1(n14100), .A2(sram_rdata_b7[31]), .A3(n2340), .A4(
        sram_rdata_a7[31]), .Y(N294) );
  AO22X1_HVT U1862 ( .A1(n14100), .A2(sram_rdata_b8[0]), .A3(n2320), .A4(
        sram_rdata_a8[0]), .Y(N295) );
  AO22X1_HVT U1863 ( .A1(n2680), .A2(sram_rdata_b8[1]), .A3(n2290), .A4(
        sram_rdata_a8[1]), .Y(N296) );
  AO22X1_HVT U1864 ( .A1(n14300), .A2(sram_rdata_b8[2]), .A3(n2380), .A4(
        sram_rdata_a8[2]), .Y(N297) );
  AO22X1_HVT U1865 ( .A1(n2640), .A2(sram_rdata_b8[3]), .A3(n2340), .A4(
        sram_rdata_a8[3]), .Y(N298) );
  AO22X1_HVT U1866 ( .A1(n14000), .A2(sram_rdata_b8[4]), .A3(n2350), .A4(
        sram_rdata_a8[4]), .Y(N299) );
  AO22X1_HVT U1867 ( .A1(n14200), .A2(sram_rdata_b8[5]), .A3(n2310), .A4(
        sram_rdata_a8[5]), .Y(N300) );
  AO22X1_HVT U1868 ( .A1(n2670), .A2(sram_rdata_b8[6]), .A3(n2300), .A4(
        sram_rdata_a8[6]), .Y(N301) );
  AO22X1_HVT U1869 ( .A1(n2650), .A2(sram_rdata_b8[7]), .A3(n2390), .A4(
        sram_rdata_a8[7]), .Y(N302) );
  AO22X1_HVT U1870 ( .A1(n2650), .A2(sram_rdata_b8[8]), .A3(n2350), .A4(
        sram_rdata_a8[8]), .Y(N303) );
  AO22X1_HVT U1871 ( .A1(n10200), .A2(sram_rdata_b8[9]), .A3(n2330), .A4(
        sram_rdata_a8[9]), .Y(N304) );
  AO22X1_HVT U1872 ( .A1(n2680), .A2(sram_rdata_b8[10]), .A3(n2350), .A4(
        sram_rdata_a8[10]), .Y(N305) );
  AO22X1_HVT U1873 ( .A1(n11700), .A2(sram_rdata_b8[11]), .A3(n2390), .A4(
        sram_rdata_a8[11]), .Y(N306) );
  AO22X1_HVT U1874 ( .A1(n14000), .A2(sram_rdata_b8[12]), .A3(n593), .A4(
        sram_rdata_a8[12]), .Y(N307) );
  AO22X1_HVT U1875 ( .A1(n2680), .A2(sram_rdata_b8[13]), .A3(n2390), .A4(
        sram_rdata_a8[13]), .Y(N308) );
  AO22X1_HVT U1876 ( .A1(n10200), .A2(sram_rdata_b8[14]), .A3(n2320), .A4(
        sram_rdata_a8[14]), .Y(N309) );
  AO22X1_HVT U1877 ( .A1(n14000), .A2(sram_rdata_b8[15]), .A3(n2290), .A4(
        sram_rdata_a8[15]), .Y(N310) );
  AO22X1_HVT U1878 ( .A1(n2650), .A2(sram_rdata_b8[16]), .A3(n2290), .A4(
        sram_rdata_a8[16]), .Y(N311) );
  AO22X1_HVT U1879 ( .A1(n2670), .A2(sram_rdata_b8[17]), .A3(n2360), .A4(
        sram_rdata_a8[17]), .Y(N312) );
  AO22X1_HVT U1880 ( .A1(n14200), .A2(sram_rdata_b8[18]), .A3(n2390), .A4(
        sram_rdata_a8[18]), .Y(N313) );
  AO22X1_HVT U1881 ( .A1(n2650), .A2(sram_rdata_b8[19]), .A3(n2360), .A4(
        sram_rdata_a8[19]), .Y(N314) );
  AO22X1_HVT U1882 ( .A1(n11700), .A2(sram_rdata_b8[20]), .A3(n2390), .A4(
        sram_rdata_a8[20]), .Y(N315) );
  AO22X1_HVT U1883 ( .A1(n14300), .A2(sram_rdata_b8[21]), .A3(n2310), .A4(
        sram_rdata_a8[21]), .Y(N316) );
  AO22X1_HVT U1884 ( .A1(n2680), .A2(sram_rdata_b8[22]), .A3(n2300), .A4(
        sram_rdata_a8[22]), .Y(N317) );
  AO22X1_HVT U1885 ( .A1(n14100), .A2(sram_rdata_b8[23]), .A3(n2320), .A4(
        sram_rdata_a8[23]), .Y(N318) );
  AO22X1_HVT U1886 ( .A1(n2640), .A2(sram_rdata_b8[24]), .A3(n2350), .A4(
        sram_rdata_a8[24]), .Y(N319) );
  AO22X1_HVT U1887 ( .A1(n11600), .A2(sram_rdata_b8[25]), .A3(n2340), .A4(
        sram_rdata_a8[25]), .Y(N320) );
  AO22X1_HVT U1888 ( .A1(n14300), .A2(sram_rdata_b8[26]), .A3(n2350), .A4(
        sram_rdata_a8[26]), .Y(N321) );
  AO22X1_HVT U1889 ( .A1(n14100), .A2(sram_rdata_b8[27]), .A3(n2390), .A4(
        sram_rdata_a8[27]), .Y(N322) );
  AO22X1_HVT U1890 ( .A1(n14100), .A2(sram_rdata_b8[28]), .A3(n2390), .A4(
        sram_rdata_a8[28]), .Y(N323) );
  AO22X1_HVT U1891 ( .A1(n2670), .A2(sram_rdata_b8[29]), .A3(n2360), .A4(
        sram_rdata_a8[29]), .Y(N324) );
  AO22X1_HVT U1892 ( .A1(n11600), .A2(sram_rdata_b8[30]), .A3(n2340), .A4(
        sram_rdata_a8[30]), .Y(N325) );
  AO22X1_HVT U1893 ( .A1(n10200), .A2(sram_rdata_b8[31]), .A3(n2290), .A4(
        sram_rdata_a8[31]), .Y(N326) );
  AO22X1_HVT U1894 ( .A1(n2640), .A2(sram_rdata_b0[0]), .A3(n2290), .A4(
        sram_rdata_a0[0]), .Y(N39) );
  AO22X1_HVT U1895 ( .A1(n2660), .A2(sram_rdata_b0[1]), .A3(n2370), .A4(
        sram_rdata_a0[1]), .Y(N40) );
  AO22X1_HVT U1896 ( .A1(n2660), .A2(sram_rdata_b0[2]), .A3(n2370), .A4(
        sram_rdata_a0[2]), .Y(N41) );
  AO22X1_HVT U1897 ( .A1(n14100), .A2(sram_rdata_b0[3]), .A3(n2330), .A4(
        sram_rdata_a0[3]), .Y(N42) );
  AO22X1_HVT U1898 ( .A1(n2670), .A2(sram_rdata_b0[4]), .A3(n2300), .A4(
        sram_rdata_a0[4]), .Y(N43) );
  AO22X1_HVT U1899 ( .A1(n2680), .A2(sram_rdata_b0[5]), .A3(n2310), .A4(
        sram_rdata_a0[5]), .Y(N44) );
  AO22X1_HVT U1900 ( .A1(n14300), .A2(sram_rdata_b0[6]), .A3(n2370), .A4(
        sram_rdata_a0[6]), .Y(N45) );
  AO22X1_HVT U1901 ( .A1(n14000), .A2(sram_rdata_b0[7]), .A3(n2330), .A4(
        sram_rdata_a0[7]), .Y(N46) );
  AO22X1_HVT U1902 ( .A1(n2640), .A2(sram_rdata_b0[8]), .A3(n2330), .A4(
        sram_rdata_a0[8]), .Y(N47) );
  AO22X1_HVT U1903 ( .A1(n10200), .A2(sram_rdata_b0[9]), .A3(n2290), .A4(
        sram_rdata_a0[9]), .Y(N48) );
  AO22X1_HVT U1904 ( .A1(n14200), .A2(sram_rdata_b0[10]), .A3(n2310), .A4(
        sram_rdata_a0[10]), .Y(N49) );
  AO22X1_HVT U1905 ( .A1(n11700), .A2(sram_rdata_b0[11]), .A3(n2370), .A4(
        sram_rdata_a0[11]), .Y(N50) );
  AO22X1_HVT U1906 ( .A1(n2650), .A2(sram_rdata_b0[12]), .A3(n2340), .A4(
        sram_rdata_a0[12]), .Y(N51) );
  AO22X1_HVT U1907 ( .A1(n2660), .A2(sram_rdata_b0[13]), .A3(n2350), .A4(
        sram_rdata_a0[13]), .Y(N52) );
  AO22X1_HVT U1908 ( .A1(n10200), .A2(sram_rdata_b0[14]), .A3(n2350), .A4(
        sram_rdata_a0[14]), .Y(N53) );
  AO22X1_HVT U1909 ( .A1(n2640), .A2(sram_rdata_b0[15]), .A3(n2370), .A4(
        sram_rdata_a0[15]), .Y(N54) );
  AO22X1_HVT U1910 ( .A1(n11700), .A2(sram_rdata_b0[16]), .A3(n2370), .A4(
        sram_rdata_a0[16]), .Y(N55) );
  AO22X1_HVT U1911 ( .A1(n14200), .A2(sram_rdata_b0[17]), .A3(n2380), .A4(
        sram_rdata_a0[17]), .Y(N56) );
  AO22X1_HVT U1912 ( .A1(n2670), .A2(sram_rdata_b0[18]), .A3(n2300), .A4(
        sram_rdata_a0[18]), .Y(N57) );
  AO22X1_HVT U1913 ( .A1(n14000), .A2(sram_rdata_b0[19]), .A3(n2310), .A4(
        sram_rdata_a0[19]), .Y(N58) );
  AO22X1_HVT U1914 ( .A1(n2660), .A2(sram_rdata_b0[20]), .A3(n2300), .A4(
        sram_rdata_a0[20]), .Y(N59) );
  AO22X1_HVT U1915 ( .A1(n2670), .A2(sram_rdata_b0[21]), .A3(n2350), .A4(
        sram_rdata_a0[21]), .Y(N60) );
  AO22X1_HVT U1916 ( .A1(n14200), .A2(sram_rdata_b0[22]), .A3(n2380), .A4(
        sram_rdata_a0[22]), .Y(N61) );
  AO22X1_HVT U1917 ( .A1(n2820), .A2(sram_rdata_b0[23]), .A3(n2340), .A4(
        sram_rdata_a0[23]), .Y(N62) );
  AO22X1_HVT U1918 ( .A1(n14000), .A2(sram_rdata_b0[24]), .A3(n2380), .A4(
        sram_rdata_a0[24]), .Y(N63) );
  AO22X1_HVT U1919 ( .A1(n11600), .A2(sram_rdata_b0[25]), .A3(n2320), .A4(
        sram_rdata_a0[25]), .Y(N64) );
  AO22X1_HVT U1920 ( .A1(n2660), .A2(sram_rdata_b0[26]), .A3(n2290), .A4(
        sram_rdata_a0[26]), .Y(N65) );
  AO22X1_HVT U1921 ( .A1(n14300), .A2(sram_rdata_b0[27]), .A3(n2300), .A4(
        sram_rdata_a0[27]), .Y(N66) );
  AO22X1_HVT U1922 ( .A1(n2640), .A2(sram_rdata_b0[28]), .A3(n2360), .A4(
        sram_rdata_a0[28]), .Y(N67) );
  AO22X1_HVT U1923 ( .A1(n14200), .A2(sram_rdata_b0[29]), .A3(n2360), .A4(
        sram_rdata_a0[29]), .Y(N68) );
  AO22X1_HVT U1924 ( .A1(n11600), .A2(sram_rdata_b0[30]), .A3(n2360), .A4(
        sram_rdata_a0[30]), .Y(N69) );
  AO22X1_HVT U1925 ( .A1(n2650), .A2(sram_rdata_b0[31]), .A3(n2380), .A4(
        sram_rdata_a0[31]), .Y(N70) );
  AO22X1_HVT U1926 ( .A1(n14200), .A2(sram_rdata_b1[0]), .A3(n2380), .A4(
        sram_rdata_a1[0]), .Y(N71) );
  AO22X1_HVT U1927 ( .A1(n14300), .A2(sram_rdata_b1[1]), .A3(n2370), .A4(
        sram_rdata_a1[1]), .Y(N72) );
  AO22X1_HVT U1928 ( .A1(n2680), .A2(sram_rdata_b1[2]), .A3(n2350), .A4(
        sram_rdata_a1[2]), .Y(N73) );
  AO22X1_HVT U1929 ( .A1(n2680), .A2(sram_rdata_b1[3]), .A3(n2300), .A4(
        sram_rdata_a1[3]), .Y(N74) );
  AO22X1_HVT U1930 ( .A1(n14000), .A2(sram_rdata_b1[4]), .A3(n2310), .A4(
        sram_rdata_a1[4]), .Y(N75) );
  AO22X1_HVT U1931 ( .A1(n2660), .A2(sram_rdata_b1[5]), .A3(n2320), .A4(
        sram_rdata_a1[5]), .Y(N76) );
  AO22X1_HVT U1932 ( .A1(n2660), .A2(sram_rdata_b1[6]), .A3(n2290), .A4(
        sram_rdata_a1[6]), .Y(N77) );
  AO22X1_HVT U1933 ( .A1(n2640), .A2(sram_rdata_b1[7]), .A3(n2360), .A4(
        sram_rdata_a1[7]), .Y(N78) );
  AO22X1_HVT U1934 ( .A1(n14100), .A2(sram_rdata_b1[8]), .A3(n2320), .A4(
        sram_rdata_a1[8]), .Y(N79) );
  AO22X1_HVT U1935 ( .A1(n10200), .A2(sram_rdata_b1[9]), .A3(n2320), .A4(
        sram_rdata_a1[9]), .Y(N80) );
  AO22X1_HVT U1936 ( .A1(n2670), .A2(sram_rdata_b1[10]), .A3(n2390), .A4(
        sram_rdata_a1[10]), .Y(N81) );
  AO22X1_HVT U1937 ( .A1(n11700), .A2(sram_rdata_b1[11]), .A3(n2330), .A4(
        sram_rdata_a1[11]), .Y(N82) );
  AO22X1_HVT U1938 ( .A1(n10200), .A2(sram_rdata_b1[12]), .A3(n2350), .A4(
        sram_rdata_a1[12]), .Y(N83) );
  AO22X1_HVT U1939 ( .A1(n14300), .A2(sram_rdata_b1[13]), .A3(n2320), .A4(
        sram_rdata_a1[13]), .Y(N84) );
  AO22X1_HVT U1940 ( .A1(n10200), .A2(sram_rdata_b1[14]), .A3(n2290), .A4(
        sram_rdata_a1[14]), .Y(N85) );
  AO22X1_HVT U1941 ( .A1(n14100), .A2(sram_rdata_b1[15]), .A3(n593), .A4(
        sram_rdata_a1[15]), .Y(N86) );
  AO22X1_HVT U1942 ( .A1(n11700), .A2(sram_rdata_b1[16]), .A3(n2330), .A4(
        sram_rdata_a1[16]), .Y(N87) );
  AO22X1_HVT U1943 ( .A1(n2680), .A2(sram_rdata_b1[17]), .A3(n2360), .A4(
        sram_rdata_a1[17]), .Y(N88) );
  AO22X1_HVT U1944 ( .A1(n14300), .A2(sram_rdata_b1[18]), .A3(n2360), .A4(
        sram_rdata_a1[18]), .Y(N89) );
  AO22X1_HVT U1945 ( .A1(n2640), .A2(sram_rdata_b1[19]), .A3(n2390), .A4(
        sram_rdata_a1[19]), .Y(N90) );
  AO22X1_HVT U1946 ( .A1(n14100), .A2(sram_rdata_b1[20]), .A3(n2390), .A4(
        sram_rdata_a1[20]), .Y(N91) );
  AO22X1_HVT U1947 ( .A1(n14200), .A2(sram_rdata_b1[21]), .A3(n2390), .A4(
        sram_rdata_a1[21]), .Y(N92) );
  AO22X1_HVT U1948 ( .A1(n2670), .A2(sram_rdata_b1[22]), .A3(n2310), .A4(
        sram_rdata_a1[22]), .Y(N93) );
  AO22X1_HVT U1949 ( .A1(n2650), .A2(sram_rdata_b1[23]), .A3(n2290), .A4(
        sram_rdata_a1[23]), .Y(N94) );
  AO22X1_HVT U1950 ( .A1(n2650), .A2(sram_rdata_b1[24]), .A3(n2310), .A4(
        sram_rdata_a1[24]), .Y(N95) );
  AO22X1_HVT U1951 ( .A1(n11600), .A2(sram_rdata_b1[25]), .A3(n2330), .A4(
        sram_rdata_a1[25]), .Y(N96) );
  AO22X1_HVT U1952 ( .A1(n2680), .A2(sram_rdata_b1[26]), .A3(n2390), .A4(
        sram_rdata_a1[26]), .Y(N97) );
  AO22X1_HVT U1953 ( .A1(n2650), .A2(sram_rdata_b1[27]), .A3(n2360), .A4(
        sram_rdata_a1[27]), .Y(N98) );
  AO22X1_HVT U1954 ( .A1(n14000), .A2(sram_rdata_b1[28]), .A3(n2370), .A4(
        sram_rdata_a1[28]), .Y(N99) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_0 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22040, n1;

  AND2X1_HVT main_gate ( .A1(net22040), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n1), .D(EN), .Q(net22040) );
  INVX0_HVT U1 ( .A(CLK), .Y(n1) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_20 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22040, n2;

  AND2X1_HVT main_gate ( .A1(net22040), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22040) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_19 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22040, n2;

  AND2X1_HVT main_gate ( .A1(net22040), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22040) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_18 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22040, n2;

  AND2X1_HVT main_gate ( .A1(net22040), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22040) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_17 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22040, n2;

  AND2X1_HVT main_gate ( .A1(net22040), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22040) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_16 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22040, n2;

  AND2X1_HVT main_gate ( .A1(net22040), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22040) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_15 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22040, n2;

  AND2X1_HVT main_gate ( .A1(net22040), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22040) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_14 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22040, n2;

  AND2X1_HVT main_gate ( .A1(net22040), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22040) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_13 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22040, n2;

  AND2X1_HVT main_gate ( .A1(net22040), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22040) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_12 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22040, n2;

  AND2X1_HVT main_gate ( .A1(net22040), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22040) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_11 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22040, n2;

  AND2X1_HVT main_gate ( .A1(net22040), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22040) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_10 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22040, n2;

  AND2X1_HVT main_gate ( .A1(net22040), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22040) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_9 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22040, n2;

  AND2X1_HVT main_gate ( .A1(net22040), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22040) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_8 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22040, n2;

  AND2X1_HVT main_gate ( .A1(net22040), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22040) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_7 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22040, n2;

  AND2X1_HVT main_gate ( .A1(net22040), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22040) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_6 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22040, n2;

  AND2X1_HVT main_gate ( .A1(net22040), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22040) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_5 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22040, n2;

  AND2X1_HVT main_gate ( .A1(net22040), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22040) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_4 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22040, n2;

  AND2X1_HVT main_gate ( .A1(net22040), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22040) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_3 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22040, n2;

  AND2X1_HVT main_gate ( .A1(net22040), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22040) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_2 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22040, n2;

  AND2X1_HVT main_gate ( .A1(net22040), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22040) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_1 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net22040, n2;

  AND2X1_HVT main_gate ( .A1(net22040), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net22040) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module bias_sel ( clk, srstn, mode, load_conv1_bias_enable, 
        load_conv2_bias0_enable, load_conv2_bias1_enable, sram_rdata_weight, 
        bias_data, conv1_bias_set_5_, conv1_bias_set_4_, conv1_bias_set_3_, 
        conv1_bias_set_2_, conv1_bias_set_1_, conv1_bias_set_0_, set_5_, 
        set_4_, set_3_, set_2_, set_1_, set_0_ );
  input [1:0] mode;
  input [99:0] sram_rdata_weight;
  output [3:0] bias_data;
  input clk, srstn, load_conv1_bias_enable, load_conv2_bias0_enable,
         load_conv2_bias1_enable, conv1_bias_set_5_, conv1_bias_set_4_,
         conv1_bias_set_3_, conv1_bias_set_2_, conv1_bias_set_1_,
         conv1_bias_set_0_, set_5_, set_4_, set_3_, set_2_, set_1_, set_0_;
  wire   net22069, net22072, net22073, net22074, net22075, net22076, net22077,
         net22078, net22079, net22080, net22083, net22088, net22089, net22090,
         net22091, net22092, net22093, net22094, net22095, net22096, net22097,
         net22100, net22105, net22106, net22107, net22108, net22109, net22110,
         net22111, net22112, net22113, net22114, net22117, net22122, net22123,
         net22124, net22125, net22126, net22127, net22128, net22129, net22130,
         net22131, net22134, net22139, net22140, net22141, net22142, net22143,
         net22144, net22145, net22146, net22147, net22148, net22151, net22156,
         net22157, net22158, net22159, net22160, net22161, net22162, net22163,
         net22164, net22165, net22168, net22173, net22174, net22175, net22176,
         net22177, net22178, net22179, net22180, net22181, net22182, net22185,
         net22190, net22191, net22192, net22193, net22194, net22195, net22196,
         net22197, net22198, net22199, net22202, net22207, net22208, net22209,
         net22210, net22211, net22212, net22213, net22214, net22215, net22216,
         net22219, net22223, net22224, net22225, net22226, net22227, net22228,
         net22229, net22230, net22231, net22232, net22233, net22236, net22249,
         net22250, net22251, net22252, net22253, net22254, net22255, net22256,
         net22257, net22258, net22261, net22266, net22267, net22268, net22269,
         net22270, net22271, net22272, net22273, net22274, net22275, net22278,
         net22283, net22284, net22285, net22286, net22287, net22288, net22289,
         net22290, net22291, net22292, net22295, net22300, net22301, net22302,
         net22303, net22304, net22305, net22306, net22307, net22308, net22309,
         net22312, net22317, net22318, net22319, net22320, net22321, net22322,
         net22323, net22324, net22325, net22326, net22329, net22334, net22335,
         net22336, net22337, net22338, net22339, net22340, net22341, net22342,
         net22343, net22346, net22351, net22352, net22353, net22354, net22355,
         net22356, net22357, net22358, net22359, net22360, net22363, net22368,
         net22369, net22370, net22371, net22372, net22373, net22374, net22375,
         net22376, net22377, net22380, net22385, net22386, net22387, net22388,
         net22389, net22390, net22391, net22392, net22393, net22394, net22397,
         net22401, net22402, net22403, net22404, net22405, net22406, net22407,
         net22408, net22409, net22410, net22411, net22414, net22425, net22431,
         net22435, net22439, net22443, net22446, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403;
  wire   [199:0] conv_weight_box;
  wire   [99:0] delay_weight;

  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_0 clk_gate_conv_weight_box_reg_0_ ( 
        .CLK(clk), .EN(net22223), .ENCLK(net22083) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_20 clk_gate_conv_weight_box_reg_2_ ( 
        .CLK(clk), .EN(net22223), .ENCLK(net22100) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_19 clk_gate_conv_weight_box_reg_5_ ( 
        .CLK(clk), .EN(net22223), .ENCLK(net22117) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_18 clk_gate_conv_weight_box_reg_7_ ( 
        .CLK(clk), .EN(net22223), .ENCLK(net22134) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_17 clk_gate_conv_weight_box_reg_10_ ( 
        .CLK(clk), .EN(net22223), .ENCLK(net22151) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_16 clk_gate_conv_weight_box_reg_12_ ( 
        .CLK(clk), .EN(net22223), .ENCLK(net22168) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_15 clk_gate_conv_weight_box_reg_15_ ( 
        .CLK(clk), .EN(net22223), .ENCLK(net22185) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_14 clk_gate_conv_weight_box_reg_17_ ( 
        .CLK(clk), .EN(net22223), .ENCLK(net22202) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_13 clk_gate_conv_weight_box_reg_20_ ( 
        .CLK(clk), .EN(net22223), .ENCLK(net22219) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_12 clk_gate_conv_weight_box_reg_22_ ( 
        .CLK(clk), .EN(net22223), .ENCLK(net22236) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_11 clk_gate_conv_weight_box_reg_25_ ( 
        .CLK(clk), .EN(net22401), .ENCLK(net22261) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_10 clk_gate_conv_weight_box_reg_27_ ( 
        .CLK(clk), .EN(net22401), .ENCLK(net22278) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_9 clk_gate_conv_weight_box_reg_30_ ( 
        .CLK(clk), .EN(net22401), .ENCLK(net22295) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_8 clk_gate_conv_weight_box_reg_32_ ( 
        .CLK(clk), .EN(net22401), .ENCLK(net22312) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_7 clk_gate_conv_weight_box_reg_35_ ( 
        .CLK(clk), .EN(net22401), .ENCLK(net22329) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_6 clk_gate_conv_weight_box_reg_37_ ( 
        .CLK(clk), .EN(net22401), .ENCLK(net22346) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_5 clk_gate_conv_weight_box_reg_40_ ( 
        .CLK(clk), .EN(net22401), .ENCLK(net22363) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_4 clk_gate_conv_weight_box_reg_42_ ( 
        .CLK(clk), .EN(net22401), .ENCLK(net22380) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_3 clk_gate_conv_weight_box_reg_45_ ( 
        .CLK(clk), .EN(net22401), .ENCLK(net22397) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_2 clk_gate_conv_weight_box_reg_47_ ( 
        .CLK(clk), .EN(net22401), .ENCLK(net22414) );
  SNPS_CLOCK_GATE_HIGH_bias_sel_mydesign_1 clk_gate_bias_data_reg ( .CLK(clk), 
        .EN(net22425), .ENCLK(net22446) );
  DFFSSRX1_HVT delay_weight_reg_99_ ( .D(1'b0), .SETB(n15), .RSTB(
        sram_rdata_weight[99]), .CLK(clk), .Q(delay_weight[99]) );
  DFFSSRX1_HVT delay_weight_reg_98_ ( .D(1'b0), .SETB(n10), .RSTB(
        sram_rdata_weight[98]), .CLK(clk), .Q(delay_weight[98]) );
  DFFSSRX1_HVT delay_weight_reg_97_ ( .D(1'b0), .SETB(n5), .RSTB(
        sram_rdata_weight[97]), .CLK(clk), .Q(delay_weight[97]) );
  DFFSSRX1_HVT delay_weight_reg_96_ ( .D(1'b0), .SETB(n16), .RSTB(
        sram_rdata_weight[96]), .CLK(clk), .Q(delay_weight[96]) );
  DFFSSRX1_HVT delay_weight_reg_95_ ( .D(1'b0), .SETB(n11), .RSTB(
        sram_rdata_weight[95]), .CLK(clk), .Q(delay_weight[95]) );
  DFFSSRX1_HVT delay_weight_reg_94_ ( .D(1'b0), .SETB(n6), .RSTB(
        sram_rdata_weight[94]), .CLK(clk), .Q(delay_weight[94]) );
  DFFSSRX1_HVT delay_weight_reg_93_ ( .D(1'b0), .SETB(n17), .RSTB(
        sram_rdata_weight[93]), .CLK(clk), .Q(delay_weight[93]) );
  DFFSSRX1_HVT delay_weight_reg_92_ ( .D(1'b0), .SETB(n12), .RSTB(
        sram_rdata_weight[92]), .CLK(clk), .Q(delay_weight[92]) );
  DFFSSRX1_HVT delay_weight_reg_91_ ( .D(1'b0), .SETB(n7), .RSTB(
        sram_rdata_weight[91]), .CLK(clk), .Q(delay_weight[91]) );
  DFFSSRX1_HVT delay_weight_reg_90_ ( .D(1'b0), .SETB(n14), .RSTB(
        sram_rdata_weight[90]), .CLK(clk), .Q(delay_weight[90]) );
  DFFSSRX1_HVT delay_weight_reg_89_ ( .D(1'b0), .SETB(n9), .RSTB(
        sram_rdata_weight[89]), .CLK(clk), .Q(delay_weight[89]) );
  DFFSSRX1_HVT delay_weight_reg_88_ ( .D(1'b0), .SETB(n4), .RSTB(
        sram_rdata_weight[88]), .CLK(clk), .Q(delay_weight[88]) );
  DFFSSRX1_HVT delay_weight_reg_87_ ( .D(1'b0), .SETB(n15), .RSTB(
        sram_rdata_weight[87]), .CLK(clk), .Q(delay_weight[87]) );
  DFFSSRX1_HVT delay_weight_reg_86_ ( .D(1'b0), .SETB(n10), .RSTB(
        sram_rdata_weight[86]), .CLK(clk), .Q(delay_weight[86]) );
  DFFSSRX1_HVT delay_weight_reg_85_ ( .D(1'b0), .SETB(n5), .RSTB(
        sram_rdata_weight[85]), .CLK(clk), .Q(delay_weight[85]) );
  DFFSSRX1_HVT delay_weight_reg_84_ ( .D(1'b0), .SETB(n16), .RSTB(
        sram_rdata_weight[84]), .CLK(clk), .Q(delay_weight[84]) );
  DFFSSRX1_HVT delay_weight_reg_83_ ( .D(1'b0), .SETB(n11), .RSTB(
        sram_rdata_weight[83]), .CLK(clk), .Q(delay_weight[83]) );
  DFFSSRX1_HVT delay_weight_reg_82_ ( .D(1'b0), .SETB(n6), .RSTB(
        sram_rdata_weight[82]), .CLK(clk), .Q(delay_weight[82]) );
  DFFSSRX1_HVT delay_weight_reg_81_ ( .D(1'b0), .SETB(n17), .RSTB(
        sram_rdata_weight[81]), .CLK(clk), .Q(delay_weight[81]) );
  DFFSSRX1_HVT delay_weight_reg_80_ ( .D(1'b0), .SETB(n12), .RSTB(
        sram_rdata_weight[80]), .CLK(clk), .Q(delay_weight[80]) );
  DFFSSRX1_HVT delay_weight_reg_79_ ( .D(1'b0), .SETB(n7), .RSTB(
        sram_rdata_weight[79]), .CLK(clk), .Q(delay_weight[79]) );
  DFFSSRX1_HVT delay_weight_reg_78_ ( .D(1'b0), .SETB(n14), .RSTB(
        sram_rdata_weight[78]), .CLK(clk), .Q(delay_weight[78]) );
  DFFSSRX1_HVT delay_weight_reg_77_ ( .D(1'b0), .SETB(n9), .RSTB(
        sram_rdata_weight[77]), .CLK(clk), .Q(delay_weight[77]) );
  DFFSSRX1_HVT delay_weight_reg_76_ ( .D(1'b0), .SETB(n4), .RSTB(
        sram_rdata_weight[76]), .CLK(clk), .Q(delay_weight[76]) );
  DFFSSRX1_HVT delay_weight_reg_75_ ( .D(1'b0), .SETB(n15), .RSTB(
        sram_rdata_weight[75]), .CLK(clk), .Q(delay_weight[75]) );
  DFFSSRX1_HVT delay_weight_reg_74_ ( .D(1'b0), .SETB(n10), .RSTB(
        sram_rdata_weight[74]), .CLK(clk), .Q(delay_weight[74]) );
  DFFSSRX1_HVT delay_weight_reg_73_ ( .D(1'b0), .SETB(n5), .RSTB(
        sram_rdata_weight[73]), .CLK(clk), .Q(delay_weight[73]) );
  DFFSSRX1_HVT delay_weight_reg_72_ ( .D(1'b0), .SETB(n16), .RSTB(
        sram_rdata_weight[72]), .CLK(clk), .Q(delay_weight[72]) );
  DFFSSRX1_HVT delay_weight_reg_71_ ( .D(1'b0), .SETB(n11), .RSTB(
        sram_rdata_weight[71]), .CLK(clk), .Q(delay_weight[71]) );
  DFFSSRX1_HVT delay_weight_reg_70_ ( .D(1'b0), .SETB(n6), .RSTB(
        sram_rdata_weight[70]), .CLK(clk), .Q(delay_weight[70]) );
  DFFSSRX1_HVT delay_weight_reg_69_ ( .D(1'b0), .SETB(n17), .RSTB(
        sram_rdata_weight[69]), .CLK(clk), .Q(delay_weight[69]) );
  DFFSSRX1_HVT delay_weight_reg_68_ ( .D(1'b0), .SETB(n12), .RSTB(
        sram_rdata_weight[68]), .CLK(clk), .Q(delay_weight[68]) );
  DFFSSRX1_HVT delay_weight_reg_67_ ( .D(1'b0), .SETB(n7), .RSTB(
        sram_rdata_weight[67]), .CLK(clk), .Q(delay_weight[67]) );
  DFFSSRX1_HVT delay_weight_reg_66_ ( .D(1'b0), .SETB(n14), .RSTB(
        sram_rdata_weight[66]), .CLK(clk), .Q(delay_weight[66]) );
  DFFSSRX1_HVT delay_weight_reg_65_ ( .D(1'b0), .SETB(n9), .RSTB(
        sram_rdata_weight[65]), .CLK(clk), .Q(delay_weight[65]) );
  DFFSSRX1_HVT delay_weight_reg_64_ ( .D(1'b0), .SETB(n4), .RSTB(
        sram_rdata_weight[64]), .CLK(clk), .Q(delay_weight[64]) );
  DFFSSRX1_HVT delay_weight_reg_63_ ( .D(1'b0), .SETB(n15), .RSTB(
        sram_rdata_weight[63]), .CLK(clk), .Q(delay_weight[63]) );
  DFFSSRX1_HVT delay_weight_reg_62_ ( .D(1'b0), .SETB(n10), .RSTB(
        sram_rdata_weight[62]), .CLK(clk), .Q(delay_weight[62]) );
  DFFSSRX1_HVT delay_weight_reg_61_ ( .D(1'b0), .SETB(n5), .RSTB(
        sram_rdata_weight[61]), .CLK(clk), .Q(delay_weight[61]) );
  DFFSSRX1_HVT delay_weight_reg_60_ ( .D(1'b0), .SETB(n16), .RSTB(
        sram_rdata_weight[60]), .CLK(clk), .Q(delay_weight[60]) );
  DFFSSRX1_HVT delay_weight_reg_59_ ( .D(1'b0), .SETB(n11), .RSTB(
        sram_rdata_weight[59]), .CLK(clk), .Q(delay_weight[59]) );
  DFFSSRX1_HVT delay_weight_reg_58_ ( .D(1'b0), .SETB(n6), .RSTB(
        sram_rdata_weight[58]), .CLK(clk), .Q(delay_weight[58]) );
  DFFSSRX1_HVT delay_weight_reg_57_ ( .D(1'b0), .SETB(n17), .RSTB(
        sram_rdata_weight[57]), .CLK(clk), .Q(delay_weight[57]) );
  DFFSSRX1_HVT delay_weight_reg_56_ ( .D(1'b0), .SETB(n12), .RSTB(
        sram_rdata_weight[56]), .CLK(clk), .Q(delay_weight[56]) );
  DFFSSRX1_HVT delay_weight_reg_55_ ( .D(1'b0), .SETB(n7), .RSTB(
        sram_rdata_weight[55]), .CLK(clk), .Q(delay_weight[55]) );
  DFFSSRX1_HVT delay_weight_reg_54_ ( .D(1'b0), .SETB(n14), .RSTB(
        sram_rdata_weight[54]), .CLK(clk), .Q(delay_weight[54]) );
  DFFSSRX1_HVT delay_weight_reg_53_ ( .D(1'b0), .SETB(n9), .RSTB(
        sram_rdata_weight[53]), .CLK(clk), .Q(delay_weight[53]) );
  DFFSSRX1_HVT delay_weight_reg_52_ ( .D(1'b0), .SETB(n4), .RSTB(
        sram_rdata_weight[52]), .CLK(clk), .Q(delay_weight[52]) );
  DFFSSRX1_HVT delay_weight_reg_51_ ( .D(1'b0), .SETB(n15), .RSTB(
        sram_rdata_weight[51]), .CLK(clk), .Q(delay_weight[51]) );
  DFFSSRX1_HVT delay_weight_reg_50_ ( .D(1'b0), .SETB(n10), .RSTB(
        sram_rdata_weight[50]), .CLK(clk), .Q(delay_weight[50]) );
  DFFSSRX1_HVT delay_weight_reg_49_ ( .D(1'b0), .SETB(n5), .RSTB(
        sram_rdata_weight[49]), .CLK(clk), .Q(delay_weight[49]) );
  DFFSSRX1_HVT delay_weight_reg_48_ ( .D(1'b0), .SETB(n16), .RSTB(
        sram_rdata_weight[48]), .CLK(clk), .Q(delay_weight[48]) );
  DFFSSRX1_HVT delay_weight_reg_47_ ( .D(1'b0), .SETB(n11), .RSTB(
        sram_rdata_weight[47]), .CLK(clk), .Q(delay_weight[47]) );
  DFFSSRX1_HVT delay_weight_reg_46_ ( .D(1'b0), .SETB(n6), .RSTB(
        sram_rdata_weight[46]), .CLK(clk), .Q(delay_weight[46]) );
  DFFSSRX1_HVT delay_weight_reg_45_ ( .D(1'b0), .SETB(n17), .RSTB(
        sram_rdata_weight[45]), .CLK(clk), .Q(delay_weight[45]) );
  DFFSSRX1_HVT delay_weight_reg_44_ ( .D(1'b0), .SETB(n12), .RSTB(
        sram_rdata_weight[44]), .CLK(clk), .Q(delay_weight[44]) );
  DFFSSRX1_HVT delay_weight_reg_43_ ( .D(1'b0), .SETB(n7), .RSTB(
        sram_rdata_weight[43]), .CLK(clk), .Q(delay_weight[43]) );
  DFFSSRX1_HVT delay_weight_reg_42_ ( .D(1'b0), .SETB(n14), .RSTB(
        sram_rdata_weight[42]), .CLK(clk), .Q(delay_weight[42]) );
  DFFSSRX1_HVT delay_weight_reg_41_ ( .D(1'b0), .SETB(n9), .RSTB(
        sram_rdata_weight[41]), .CLK(clk), .Q(delay_weight[41]) );
  DFFSSRX1_HVT delay_weight_reg_40_ ( .D(1'b0), .SETB(n4), .RSTB(
        sram_rdata_weight[40]), .CLK(clk), .Q(delay_weight[40]) );
  DFFSSRX1_HVT delay_weight_reg_39_ ( .D(1'b0), .SETB(n15), .RSTB(
        sram_rdata_weight[39]), .CLK(clk), .Q(delay_weight[39]) );
  DFFSSRX1_HVT delay_weight_reg_38_ ( .D(1'b0), .SETB(n10), .RSTB(
        sram_rdata_weight[38]), .CLK(clk), .Q(delay_weight[38]) );
  DFFSSRX1_HVT delay_weight_reg_37_ ( .D(1'b0), .SETB(n5), .RSTB(
        sram_rdata_weight[37]), .CLK(clk), .Q(delay_weight[37]) );
  DFFSSRX1_HVT delay_weight_reg_36_ ( .D(1'b0), .SETB(n16), .RSTB(
        sram_rdata_weight[36]), .CLK(clk), .Q(delay_weight[36]) );
  DFFSSRX1_HVT delay_weight_reg_35_ ( .D(1'b0), .SETB(n11), .RSTB(
        sram_rdata_weight[35]), .CLK(clk), .Q(delay_weight[35]) );
  DFFSSRX1_HVT delay_weight_reg_34_ ( .D(1'b0), .SETB(n6), .RSTB(
        sram_rdata_weight[34]), .CLK(clk), .Q(delay_weight[34]) );
  DFFSSRX1_HVT delay_weight_reg_33_ ( .D(1'b0), .SETB(n17), .RSTB(
        sram_rdata_weight[33]), .CLK(clk), .Q(delay_weight[33]) );
  DFFSSRX1_HVT delay_weight_reg_32_ ( .D(1'b0), .SETB(n12), .RSTB(
        sram_rdata_weight[32]), .CLK(clk), .Q(delay_weight[32]) );
  DFFSSRX1_HVT delay_weight_reg_31_ ( .D(1'b0), .SETB(n7), .RSTB(
        sram_rdata_weight[31]), .CLK(clk), .Q(delay_weight[31]) );
  DFFSSRX1_HVT delay_weight_reg_30_ ( .D(1'b0), .SETB(n14), .RSTB(
        sram_rdata_weight[30]), .CLK(clk), .Q(delay_weight[30]) );
  DFFSSRX1_HVT delay_weight_reg_29_ ( .D(1'b0), .SETB(n9), .RSTB(
        sram_rdata_weight[29]), .CLK(clk), .Q(delay_weight[29]) );
  DFFSSRX1_HVT delay_weight_reg_28_ ( .D(1'b0), .SETB(n4), .RSTB(
        sram_rdata_weight[28]), .CLK(clk), .Q(delay_weight[28]) );
  DFFSSRX1_HVT delay_weight_reg_27_ ( .D(1'b0), .SETB(n15), .RSTB(
        sram_rdata_weight[27]), .CLK(clk), .Q(delay_weight[27]) );
  DFFSSRX1_HVT delay_weight_reg_26_ ( .D(1'b0), .SETB(n10), .RSTB(
        sram_rdata_weight[26]), .CLK(clk), .Q(delay_weight[26]) );
  DFFSSRX1_HVT delay_weight_reg_25_ ( .D(1'b0), .SETB(n5), .RSTB(
        sram_rdata_weight[25]), .CLK(clk), .Q(delay_weight[25]) );
  DFFSSRX1_HVT delay_weight_reg_24_ ( .D(1'b0), .SETB(n16), .RSTB(
        sram_rdata_weight[24]), .CLK(clk), .Q(delay_weight[24]) );
  DFFSSRX1_HVT delay_weight_reg_23_ ( .D(1'b0), .SETB(n11), .RSTB(
        sram_rdata_weight[23]), .CLK(clk), .Q(delay_weight[23]) );
  DFFSSRX1_HVT delay_weight_reg_22_ ( .D(1'b0), .SETB(n6), .RSTB(
        sram_rdata_weight[22]), .CLK(clk), .Q(delay_weight[22]) );
  DFFSSRX1_HVT delay_weight_reg_21_ ( .D(1'b0), .SETB(n17), .RSTB(
        sram_rdata_weight[21]), .CLK(clk), .Q(delay_weight[21]) );
  DFFSSRX1_HVT delay_weight_reg_20_ ( .D(1'b0), .SETB(n12), .RSTB(
        sram_rdata_weight[20]), .CLK(clk), .Q(delay_weight[20]) );
  DFFSSRX1_HVT delay_weight_reg_19_ ( .D(1'b0), .SETB(n7), .RSTB(
        sram_rdata_weight[19]), .CLK(clk), .Q(delay_weight[19]) );
  DFFSSRX1_HVT delay_weight_reg_18_ ( .D(1'b0), .SETB(n14), .RSTB(
        sram_rdata_weight[18]), .CLK(clk), .Q(delay_weight[18]) );
  DFFSSRX1_HVT delay_weight_reg_17_ ( .D(1'b0), .SETB(n9), .RSTB(
        sram_rdata_weight[17]), .CLK(clk), .Q(delay_weight[17]) );
  DFFSSRX1_HVT delay_weight_reg_16_ ( .D(1'b0), .SETB(n4), .RSTB(
        sram_rdata_weight[16]), .CLK(clk), .Q(delay_weight[16]) );
  DFFSSRX1_HVT delay_weight_reg_15_ ( .D(1'b0), .SETB(n15), .RSTB(
        sram_rdata_weight[15]), .CLK(clk), .Q(delay_weight[15]) );
  DFFSSRX1_HVT delay_weight_reg_14_ ( .D(1'b0), .SETB(n10), .RSTB(
        sram_rdata_weight[14]), .CLK(clk), .Q(delay_weight[14]) );
  DFFSSRX1_HVT delay_weight_reg_13_ ( .D(1'b0), .SETB(n5), .RSTB(
        sram_rdata_weight[13]), .CLK(clk), .Q(delay_weight[13]) );
  DFFSSRX1_HVT delay_weight_reg_12_ ( .D(1'b0), .SETB(n16), .RSTB(
        sram_rdata_weight[12]), .CLK(clk), .Q(delay_weight[12]) );
  DFFSSRX1_HVT delay_weight_reg_11_ ( .D(1'b0), .SETB(n11), .RSTB(
        sram_rdata_weight[11]), .CLK(clk), .Q(delay_weight[11]) );
  DFFSSRX1_HVT delay_weight_reg_10_ ( .D(1'b0), .SETB(n6), .RSTB(
        sram_rdata_weight[10]), .CLK(clk), .Q(delay_weight[10]) );
  DFFSSRX1_HVT delay_weight_reg_9_ ( .D(1'b0), .SETB(n17), .RSTB(
        sram_rdata_weight[9]), .CLK(clk), .Q(delay_weight[9]) );
  DFFSSRX1_HVT delay_weight_reg_8_ ( .D(1'b0), .SETB(n12), .RSTB(
        sram_rdata_weight[8]), .CLK(clk), .Q(delay_weight[8]) );
  DFFSSRX1_HVT delay_weight_reg_7_ ( .D(1'b0), .SETB(n7), .RSTB(
        sram_rdata_weight[7]), .CLK(clk), .Q(delay_weight[7]) );
  DFFSSRX1_HVT delay_weight_reg_6_ ( .D(1'b0), .SETB(n14), .RSTB(
        sram_rdata_weight[6]), .CLK(clk), .Q(delay_weight[6]) );
  DFFSSRX1_HVT delay_weight_reg_5_ ( .D(1'b0), .SETB(n9), .RSTB(
        sram_rdata_weight[5]), .CLK(clk), .Q(delay_weight[5]) );
  DFFSSRX1_HVT delay_weight_reg_4_ ( .D(1'b0), .SETB(n4), .RSTB(
        sram_rdata_weight[4]), .CLK(clk), .Q(delay_weight[4]) );
  DFFSSRX1_HVT delay_weight_reg_3_ ( .D(1'b0), .SETB(n15), .RSTB(
        sram_rdata_weight[3]), .CLK(clk), .Q(delay_weight[3]) );
  DFFSSRX1_HVT delay_weight_reg_2_ ( .D(1'b0), .SETB(n10), .RSTB(
        sram_rdata_weight[2]), .CLK(clk), .Q(delay_weight[2]) );
  DFFSSRX1_HVT delay_weight_reg_1_ ( .D(1'b0), .SETB(n5), .RSTB(
        sram_rdata_weight[1]), .CLK(clk), .Q(delay_weight[1]) );
  DFFSSRX1_HVT delay_weight_reg_0_ ( .D(1'b0), .SETB(n16), .RSTB(
        sram_rdata_weight[0]), .CLK(clk), .Q(delay_weight[0]) );
  DFFSSRX1_HVT conv_weight_box_reg_0__3_ ( .D(1'b0), .SETB(n11), .RSTB(
        net22069), .CLK(net22083), .Q(conv_weight_box[199]) );
  DFFSSRX1_HVT conv_weight_box_reg_0__2_ ( .D(1'b0), .SETB(n6), .RSTB(net22072), .CLK(net22083), .Q(conv_weight_box[198]) );
  DFFSSRX1_HVT conv_weight_box_reg_0__1_ ( .D(1'b0), .SETB(n17), .RSTB(
        net22073), .CLK(net22083), .Q(conv_weight_box[197]) );
  DFFSSRX1_HVT conv_weight_box_reg_0__0_ ( .D(1'b0), .SETB(n12), .RSTB(
        net22074), .CLK(net22083), .Q(conv_weight_box[196]) );
  DFFSSRX1_HVT conv_weight_box_reg_1__3_ ( .D(1'b0), .SETB(n7), .RSTB(net22075), .CLK(net22083), .Q(conv_weight_box[195]) );
  DFFSSRX1_HVT conv_weight_box_reg_1__2_ ( .D(1'b0), .SETB(n14), .RSTB(
        net22076), .CLK(net22083), .Q(conv_weight_box[194]) );
  DFFSSRX1_HVT conv_weight_box_reg_1__1_ ( .D(1'b0), .SETB(n9), .RSTB(net22077), .CLK(net22083), .Q(conv_weight_box[193]) );
  DFFSSRX1_HVT conv_weight_box_reg_1__0_ ( .D(1'b0), .SETB(n4), .RSTB(net22078), .CLK(net22083), .Q(conv_weight_box[192]) );
  DFFSSRX1_HVT conv_weight_box_reg_2__3_ ( .D(1'b0), .SETB(n15), .RSTB(
        net22079), .CLK(net22083), .Q(conv_weight_box[191]) );
  DFFSSRX1_HVT conv_weight_box_reg_2__2_ ( .D(1'b0), .SETB(n10), .RSTB(
        net22080), .CLK(net22083), .Q(conv_weight_box[190]) );
  DFFSSRX1_HVT conv_weight_box_reg_2__1_ ( .D(1'b0), .SETB(n5), .RSTB(net22088), .CLK(net22100), .Q(conv_weight_box[189]) );
  DFFSSRX1_HVT conv_weight_box_reg_2__0_ ( .D(1'b0), .SETB(n16), .RSTB(
        net22089), .CLK(net22100), .Q(conv_weight_box[188]) );
  DFFSSRX1_HVT conv_weight_box_reg_3__3_ ( .D(1'b0), .SETB(n11), .RSTB(
        net22090), .CLK(net22100), .Q(conv_weight_box[187]) );
  DFFSSRX1_HVT conv_weight_box_reg_3__2_ ( .D(1'b0), .SETB(n6), .RSTB(net22091), .CLK(net22100), .Q(conv_weight_box[186]) );
  DFFSSRX1_HVT conv_weight_box_reg_3__1_ ( .D(1'b0), .SETB(n17), .RSTB(
        net22092), .CLK(net22100), .Q(conv_weight_box[185]) );
  DFFSSRX1_HVT conv_weight_box_reg_3__0_ ( .D(1'b0), .SETB(n12), .RSTB(
        net22093), .CLK(net22100), .Q(conv_weight_box[184]) );
  DFFSSRX1_HVT conv_weight_box_reg_4__3_ ( .D(1'b0), .SETB(n7), .RSTB(net22094), .CLK(net22100), .Q(conv_weight_box[183]) );
  DFFSSRX1_HVT conv_weight_box_reg_4__2_ ( .D(1'b0), .SETB(n14), .RSTB(
        net22095), .CLK(net22100), .Q(conv_weight_box[182]) );
  DFFSSRX1_HVT conv_weight_box_reg_4__1_ ( .D(1'b0), .SETB(n9), .RSTB(net22096), .CLK(net22100), .Q(conv_weight_box[181]) );
  DFFSSRX1_HVT conv_weight_box_reg_4__0_ ( .D(1'b0), .SETB(n4), .RSTB(net22097), .CLK(net22100), .Q(conv_weight_box[180]) );
  DFFSSRX1_HVT conv_weight_box_reg_5__3_ ( .D(1'b0), .SETB(n15), .RSTB(
        net22105), .CLK(net22117), .Q(conv_weight_box[179]) );
  DFFSSRX1_HVT conv_weight_box_reg_5__2_ ( .D(1'b0), .SETB(n10), .RSTB(
        net22106), .CLK(net22117), .Q(conv_weight_box[178]) );
  DFFSSRX1_HVT conv_weight_box_reg_5__1_ ( .D(1'b0), .SETB(n5), .RSTB(net22107), .CLK(net22117), .Q(conv_weight_box[177]) );
  DFFSSRX1_HVT conv_weight_box_reg_5__0_ ( .D(1'b0), .SETB(n16), .RSTB(
        net22108), .CLK(net22117), .Q(conv_weight_box[176]) );
  DFFSSRX1_HVT conv_weight_box_reg_6__3_ ( .D(1'b0), .SETB(n11), .RSTB(
        net22109), .CLK(net22117), .Q(conv_weight_box[175]) );
  DFFSSRX1_HVT conv_weight_box_reg_6__2_ ( .D(1'b0), .SETB(n6), .RSTB(net22110), .CLK(net22117), .Q(conv_weight_box[174]) );
  DFFSSRX1_HVT conv_weight_box_reg_6__1_ ( .D(1'b0), .SETB(n17), .RSTB(
        net22111), .CLK(net22117), .Q(conv_weight_box[173]) );
  DFFSSRX1_HVT conv_weight_box_reg_6__0_ ( .D(1'b0), .SETB(n12), .RSTB(
        net22112), .CLK(net22117), .Q(conv_weight_box[172]) );
  DFFSSRX1_HVT conv_weight_box_reg_7__3_ ( .D(1'b0), .SETB(n7), .RSTB(net22113), .CLK(net22117), .Q(conv_weight_box[171]) );
  DFFSSRX1_HVT conv_weight_box_reg_7__2_ ( .D(1'b0), .SETB(n14), .RSTB(
        net22114), .CLK(net22117), .Q(conv_weight_box[170]) );
  DFFSSRX1_HVT conv_weight_box_reg_7__1_ ( .D(1'b0), .SETB(n9), .RSTB(net22122), .CLK(net22134), .Q(conv_weight_box[169]) );
  DFFSSRX1_HVT conv_weight_box_reg_7__0_ ( .D(1'b0), .SETB(n4), .RSTB(net22123), .CLK(net22134), .Q(conv_weight_box[168]) );
  DFFSSRX1_HVT conv_weight_box_reg_8__3_ ( .D(1'b0), .SETB(n15), .RSTB(
        net22124), .CLK(net22134), .Q(conv_weight_box[167]) );
  DFFSSRX1_HVT conv_weight_box_reg_8__2_ ( .D(1'b0), .SETB(n10), .RSTB(
        net22125), .CLK(net22134), .Q(conv_weight_box[166]) );
  DFFSSRX1_HVT conv_weight_box_reg_8__1_ ( .D(1'b0), .SETB(n5), .RSTB(net22126), .CLK(net22134), .Q(conv_weight_box[165]) );
  DFFSSRX1_HVT conv_weight_box_reg_8__0_ ( .D(1'b0), .SETB(n16), .RSTB(
        net22127), .CLK(net22134), .Q(conv_weight_box[164]) );
  DFFSSRX1_HVT conv_weight_box_reg_9__3_ ( .D(1'b0), .SETB(n11), .RSTB(
        net22128), .CLK(net22134), .Q(conv_weight_box[163]) );
  DFFSSRX1_HVT conv_weight_box_reg_9__2_ ( .D(1'b0), .SETB(n6), .RSTB(net22129), .CLK(net22134), .Q(conv_weight_box[162]) );
  DFFSSRX1_HVT conv_weight_box_reg_9__1_ ( .D(1'b0), .SETB(n17), .RSTB(
        net22130), .CLK(net22134), .Q(conv_weight_box[161]) );
  DFFSSRX1_HVT conv_weight_box_reg_9__0_ ( .D(1'b0), .SETB(n12), .RSTB(
        net22131), .CLK(net22134), .Q(conv_weight_box[160]) );
  DFFSSRX1_HVT conv_weight_box_reg_10__3_ ( .D(1'b0), .SETB(n7), .RSTB(
        net22139), .CLK(net22151), .Q(conv_weight_box[159]) );
  DFFSSRX1_HVT conv_weight_box_reg_10__2_ ( .D(1'b0), .SETB(n14), .RSTB(
        net22140), .CLK(net22151), .Q(conv_weight_box[158]) );
  DFFSSRX1_HVT conv_weight_box_reg_10__1_ ( .D(1'b0), .SETB(n9), .RSTB(
        net22141), .CLK(net22151), .Q(conv_weight_box[157]) );
  DFFSSRX1_HVT conv_weight_box_reg_10__0_ ( .D(1'b0), .SETB(n4), .RSTB(
        net22142), .CLK(net22151), .Q(conv_weight_box[156]) );
  DFFSSRX1_HVT conv_weight_box_reg_11__3_ ( .D(1'b0), .SETB(n15), .RSTB(
        net22143), .CLK(net22151), .Q(conv_weight_box[155]) );
  DFFSSRX1_HVT conv_weight_box_reg_11__2_ ( .D(1'b0), .SETB(n10), .RSTB(
        net22144), .CLK(net22151), .Q(conv_weight_box[154]) );
  DFFSSRX1_HVT conv_weight_box_reg_11__1_ ( .D(1'b0), .SETB(n5), .RSTB(
        net22145), .CLK(net22151), .Q(conv_weight_box[153]) );
  DFFSSRX1_HVT conv_weight_box_reg_11__0_ ( .D(1'b0), .SETB(n16), .RSTB(
        net22146), .CLK(net22151), .Q(conv_weight_box[152]) );
  DFFSSRX1_HVT conv_weight_box_reg_12__3_ ( .D(1'b0), .SETB(n11), .RSTB(
        net22147), .CLK(net22151), .Q(conv_weight_box[151]) );
  DFFSSRX1_HVT conv_weight_box_reg_12__2_ ( .D(1'b0), .SETB(n6), .RSTB(
        net22148), .CLK(net22151), .Q(conv_weight_box[150]) );
  DFFSSRX1_HVT conv_weight_box_reg_12__1_ ( .D(1'b0), .SETB(n17), .RSTB(
        net22156), .CLK(net22168), .Q(conv_weight_box[149]) );
  DFFSSRX1_HVT conv_weight_box_reg_12__0_ ( .D(1'b0), .SETB(n12), .RSTB(
        net22157), .CLK(net22168), .Q(conv_weight_box[148]) );
  DFFSSRX1_HVT conv_weight_box_reg_13__3_ ( .D(1'b0), .SETB(n7), .RSTB(
        net22158), .CLK(net22168), .Q(conv_weight_box[147]) );
  DFFSSRX1_HVT conv_weight_box_reg_13__2_ ( .D(1'b0), .SETB(n14), .RSTB(
        net22159), .CLK(net22168), .Q(conv_weight_box[146]) );
  DFFSSRX1_HVT conv_weight_box_reg_13__1_ ( .D(1'b0), .SETB(n9), .RSTB(
        net22160), .CLK(net22168), .Q(conv_weight_box[145]) );
  DFFSSRX1_HVT conv_weight_box_reg_13__0_ ( .D(1'b0), .SETB(n4), .RSTB(
        net22161), .CLK(net22168), .Q(conv_weight_box[144]) );
  DFFSSRX1_HVT conv_weight_box_reg_14__3_ ( .D(1'b0), .SETB(n15), .RSTB(
        net22162), .CLK(net22168), .Q(conv_weight_box[143]) );
  DFFSSRX1_HVT conv_weight_box_reg_14__2_ ( .D(1'b0), .SETB(n10), .RSTB(
        net22163), .CLK(net22168), .Q(conv_weight_box[142]) );
  DFFSSRX1_HVT conv_weight_box_reg_14__1_ ( .D(1'b0), .SETB(n5), .RSTB(
        net22164), .CLK(net22168), .Q(conv_weight_box[141]) );
  DFFSSRX1_HVT conv_weight_box_reg_14__0_ ( .D(1'b0), .SETB(n16), .RSTB(
        net22165), .CLK(net22168), .Q(conv_weight_box[140]) );
  DFFSSRX1_HVT conv_weight_box_reg_15__3_ ( .D(1'b0), .SETB(n11), .RSTB(
        net22173), .CLK(net22185), .Q(conv_weight_box[139]) );
  DFFSSRX1_HVT conv_weight_box_reg_15__2_ ( .D(1'b0), .SETB(n6), .RSTB(
        net22174), .CLK(net22185), .Q(conv_weight_box[138]) );
  DFFSSRX1_HVT conv_weight_box_reg_15__1_ ( .D(1'b0), .SETB(n17), .RSTB(
        net22175), .CLK(net22185), .Q(conv_weight_box[137]) );
  DFFSSRX1_HVT conv_weight_box_reg_15__0_ ( .D(1'b0), .SETB(n12), .RSTB(
        net22176), .CLK(net22185), .Q(conv_weight_box[136]) );
  DFFSSRX1_HVT conv_weight_box_reg_16__3_ ( .D(1'b0), .SETB(n7), .RSTB(
        net22177), .CLK(net22185), .Q(conv_weight_box[135]) );
  DFFSSRX1_HVT conv_weight_box_reg_16__2_ ( .D(1'b0), .SETB(n14), .RSTB(
        net22178), .CLK(net22185), .Q(conv_weight_box[134]) );
  DFFSSRX1_HVT conv_weight_box_reg_16__1_ ( .D(1'b0), .SETB(n9), .RSTB(
        net22179), .CLK(net22185), .Q(conv_weight_box[133]) );
  DFFSSRX1_HVT conv_weight_box_reg_16__0_ ( .D(1'b0), .SETB(n4), .RSTB(
        net22180), .CLK(net22185), .Q(conv_weight_box[132]) );
  DFFSSRX1_HVT conv_weight_box_reg_17__3_ ( .D(1'b0), .SETB(n15), .RSTB(
        net22181), .CLK(net22185), .Q(conv_weight_box[131]) );
  DFFSSRX1_HVT conv_weight_box_reg_17__2_ ( .D(1'b0), .SETB(n10), .RSTB(
        net22182), .CLK(net22185), .Q(conv_weight_box[130]) );
  DFFSSRX1_HVT conv_weight_box_reg_17__1_ ( .D(1'b0), .SETB(n5), .RSTB(
        net22190), .CLK(net22202), .Q(conv_weight_box[129]) );
  DFFSSRX1_HVT conv_weight_box_reg_17__0_ ( .D(1'b0), .SETB(n16), .RSTB(
        net22191), .CLK(net22202), .Q(conv_weight_box[128]) );
  DFFSSRX1_HVT conv_weight_box_reg_18__3_ ( .D(1'b0), .SETB(n11), .RSTB(
        net22192), .CLK(net22202), .Q(conv_weight_box[127]) );
  DFFSSRX1_HVT conv_weight_box_reg_18__2_ ( .D(1'b0), .SETB(n6), .RSTB(
        net22193), .CLK(net22202), .Q(conv_weight_box[126]) );
  DFFSSRX1_HVT conv_weight_box_reg_18__1_ ( .D(1'b0), .SETB(n17), .RSTB(
        net22194), .CLK(net22202), .Q(conv_weight_box[125]) );
  DFFSSRX1_HVT conv_weight_box_reg_18__0_ ( .D(1'b0), .SETB(n12), .RSTB(
        net22195), .CLK(net22202), .Q(conv_weight_box[124]) );
  DFFSSRX1_HVT conv_weight_box_reg_19__3_ ( .D(1'b0), .SETB(n7), .RSTB(
        net22196), .CLK(net22202), .Q(conv_weight_box[123]) );
  DFFSSRX1_HVT conv_weight_box_reg_19__2_ ( .D(1'b0), .SETB(n14), .RSTB(
        net22197), .CLK(net22202), .Q(conv_weight_box[122]) );
  DFFSSRX1_HVT conv_weight_box_reg_19__1_ ( .D(1'b0), .SETB(n9), .RSTB(
        net22198), .CLK(net22202), .Q(conv_weight_box[121]) );
  DFFSSRX1_HVT conv_weight_box_reg_19__0_ ( .D(1'b0), .SETB(n4), .RSTB(
        net22199), .CLK(net22202), .Q(conv_weight_box[120]) );
  DFFSSRX1_HVT conv_weight_box_reg_20__3_ ( .D(1'b0), .SETB(n15), .RSTB(
        net22207), .CLK(net22219), .Q(conv_weight_box[119]) );
  DFFSSRX1_HVT conv_weight_box_reg_20__2_ ( .D(1'b0), .SETB(n10), .RSTB(
        net22208), .CLK(net22219), .Q(conv_weight_box[118]) );
  DFFSSRX1_HVT conv_weight_box_reg_20__1_ ( .D(1'b0), .SETB(n5), .RSTB(
        net22209), .CLK(net22219), .Q(conv_weight_box[117]) );
  DFFSSRX1_HVT conv_weight_box_reg_20__0_ ( .D(1'b0), .SETB(n16), .RSTB(
        net22210), .CLK(net22219), .Q(conv_weight_box[116]) );
  DFFSSRX1_HVT conv_weight_box_reg_21__3_ ( .D(1'b0), .SETB(n11), .RSTB(
        net22211), .CLK(net22219), .Q(conv_weight_box[115]) );
  DFFSSRX1_HVT conv_weight_box_reg_21__2_ ( .D(1'b0), .SETB(n6), .RSTB(
        net22212), .CLK(net22219), .Q(conv_weight_box[114]) );
  DFFSSRX1_HVT conv_weight_box_reg_21__1_ ( .D(1'b0), .SETB(n17), .RSTB(
        net22213), .CLK(net22219), .Q(conv_weight_box[113]) );
  DFFSSRX1_HVT conv_weight_box_reg_21__0_ ( .D(1'b0), .SETB(n12), .RSTB(
        net22214), .CLK(net22219), .Q(conv_weight_box[112]) );
  DFFSSRX1_HVT conv_weight_box_reg_22__3_ ( .D(1'b0), .SETB(n7), .RSTB(
        net22215), .CLK(net22219), .Q(conv_weight_box[111]) );
  DFFSSRX1_HVT conv_weight_box_reg_22__2_ ( .D(1'b0), .SETB(n14), .RSTB(
        net22216), .CLK(net22219), .Q(conv_weight_box[110]) );
  DFFSSRX1_HVT conv_weight_box_reg_22__1_ ( .D(1'b0), .SETB(n9), .RSTB(
        net22224), .CLK(net22236), .Q(conv_weight_box[109]) );
  DFFSSRX1_HVT conv_weight_box_reg_22__0_ ( .D(1'b0), .SETB(n4), .RSTB(
        net22225), .CLK(net22236), .Q(conv_weight_box[108]) );
  DFFSSRX1_HVT conv_weight_box_reg_23__3_ ( .D(1'b0), .SETB(n15), .RSTB(
        net22226), .CLK(net22236), .Q(conv_weight_box[107]) );
  DFFSSRX1_HVT conv_weight_box_reg_23__2_ ( .D(1'b0), .SETB(n10), .RSTB(
        net22227), .CLK(net22236), .Q(conv_weight_box[106]) );
  DFFSSRX1_HVT conv_weight_box_reg_23__1_ ( .D(1'b0), .SETB(n5), .RSTB(
        net22228), .CLK(net22236), .Q(conv_weight_box[105]) );
  DFFSSRX1_HVT conv_weight_box_reg_23__0_ ( .D(1'b0), .SETB(n16), .RSTB(
        net22229), .CLK(net22236), .Q(conv_weight_box[104]) );
  DFFSSRX1_HVT conv_weight_box_reg_24__3_ ( .D(1'b0), .SETB(n11), .RSTB(
        net22230), .CLK(net22236), .Q(conv_weight_box[103]) );
  DFFSSRX1_HVT conv_weight_box_reg_24__2_ ( .D(1'b0), .SETB(n6), .RSTB(
        net22231), .CLK(net22236), .Q(conv_weight_box[102]) );
  DFFSSRX1_HVT conv_weight_box_reg_24__1_ ( .D(1'b0), .SETB(n17), .RSTB(
        net22232), .CLK(net22236), .Q(conv_weight_box[101]) );
  DFFSSRX1_HVT conv_weight_box_reg_24__0_ ( .D(1'b0), .SETB(n12), .RSTB(
        net22233), .CLK(net22236), .Q(conv_weight_box[100]) );
  DFFSSRX1_HVT conv_weight_box_reg_25__3_ ( .D(1'b0), .SETB(n7), .RSTB(
        net22249), .CLK(net22261), .Q(conv_weight_box[99]) );
  DFFSSRX1_HVT conv_weight_box_reg_25__2_ ( .D(1'b0), .SETB(n14), .RSTB(
        net22250), .CLK(net22261), .Q(conv_weight_box[98]) );
  DFFSSRX1_HVT conv_weight_box_reg_25__1_ ( .D(1'b0), .SETB(n9), .RSTB(
        net22251), .CLK(net22261), .Q(conv_weight_box[97]) );
  DFFSSRX1_HVT conv_weight_box_reg_25__0_ ( .D(1'b0), .SETB(n4), .RSTB(
        net22252), .CLK(net22261), .Q(conv_weight_box[96]) );
  DFFSSRX1_HVT conv_weight_box_reg_26__3_ ( .D(1'b0), .SETB(n15), .RSTB(
        net22253), .CLK(net22261), .Q(conv_weight_box[95]) );
  DFFSSRX1_HVT conv_weight_box_reg_26__2_ ( .D(1'b0), .SETB(n10), .RSTB(
        net22254), .CLK(net22261), .Q(conv_weight_box[94]) );
  DFFSSRX1_HVT conv_weight_box_reg_26__1_ ( .D(1'b0), .SETB(n5), .RSTB(
        net22255), .CLK(net22261), .Q(conv_weight_box[93]) );
  DFFSSRX1_HVT conv_weight_box_reg_26__0_ ( .D(1'b0), .SETB(n16), .RSTB(
        net22256), .CLK(net22261), .Q(conv_weight_box[92]) );
  DFFSSRX1_HVT conv_weight_box_reg_27__3_ ( .D(1'b0), .SETB(n11), .RSTB(
        net22257), .CLK(net22261), .Q(conv_weight_box[91]) );
  DFFSSRX1_HVT conv_weight_box_reg_27__2_ ( .D(1'b0), .SETB(n6), .RSTB(
        net22258), .CLK(net22261), .Q(conv_weight_box[90]) );
  DFFSSRX1_HVT conv_weight_box_reg_27__1_ ( .D(1'b0), .SETB(n17), .RSTB(
        net22266), .CLK(net22278), .Q(conv_weight_box[89]) );
  DFFSSRX1_HVT conv_weight_box_reg_27__0_ ( .D(1'b0), .SETB(n12), .RSTB(
        net22267), .CLK(net22278), .Q(conv_weight_box[88]) );
  DFFSSRX1_HVT conv_weight_box_reg_28__3_ ( .D(1'b0), .SETB(n7), .RSTB(
        net22268), .CLK(net22278), .Q(conv_weight_box[87]) );
  DFFSSRX1_HVT conv_weight_box_reg_28__2_ ( .D(1'b0), .SETB(n14), .RSTB(
        net22269), .CLK(net22278), .Q(conv_weight_box[86]) );
  DFFSSRX1_HVT conv_weight_box_reg_28__1_ ( .D(1'b0), .SETB(n9), .RSTB(
        net22270), .CLK(net22278), .Q(conv_weight_box[85]) );
  DFFSSRX1_HVT conv_weight_box_reg_28__0_ ( .D(1'b0), .SETB(n4), .RSTB(
        net22271), .CLK(net22278), .Q(conv_weight_box[84]) );
  DFFSSRX1_HVT conv_weight_box_reg_29__3_ ( .D(1'b0), .SETB(n15), .RSTB(
        net22272), .CLK(net22278), .Q(conv_weight_box[83]) );
  DFFSSRX1_HVT conv_weight_box_reg_29__2_ ( .D(1'b0), .SETB(n10), .RSTB(
        net22273), .CLK(net22278), .Q(conv_weight_box[82]) );
  DFFSSRX1_HVT conv_weight_box_reg_29__1_ ( .D(1'b0), .SETB(n5), .RSTB(
        net22274), .CLK(net22278), .Q(conv_weight_box[81]) );
  DFFSSRX1_HVT conv_weight_box_reg_29__0_ ( .D(1'b0), .SETB(n16), .RSTB(
        net22275), .CLK(net22278), .Q(conv_weight_box[80]) );
  DFFSSRX1_HVT conv_weight_box_reg_30__3_ ( .D(1'b0), .SETB(n11), .RSTB(
        net22283), .CLK(net22295), .Q(conv_weight_box[79]) );
  DFFSSRX1_HVT conv_weight_box_reg_30__2_ ( .D(1'b0), .SETB(n6), .RSTB(
        net22284), .CLK(net22295), .Q(conv_weight_box[78]) );
  DFFSSRX1_HVT conv_weight_box_reg_30__1_ ( .D(1'b0), .SETB(n17), .RSTB(
        net22285), .CLK(net22295), .Q(conv_weight_box[77]) );
  DFFSSRX1_HVT conv_weight_box_reg_30__0_ ( .D(1'b0), .SETB(n12), .RSTB(
        net22286), .CLK(net22295), .Q(conv_weight_box[76]) );
  DFFSSRX1_HVT conv_weight_box_reg_31__3_ ( .D(1'b0), .SETB(n7), .RSTB(
        net22287), .CLK(net22295), .Q(conv_weight_box[75]) );
  DFFSSRX1_HVT conv_weight_box_reg_31__2_ ( .D(1'b0), .SETB(n14), .RSTB(
        net22288), .CLK(net22295), .Q(conv_weight_box[74]) );
  DFFSSRX1_HVT conv_weight_box_reg_31__1_ ( .D(1'b0), .SETB(n9), .RSTB(
        net22289), .CLK(net22295), .Q(conv_weight_box[73]) );
  DFFSSRX1_HVT conv_weight_box_reg_31__0_ ( .D(1'b0), .SETB(n4), .RSTB(
        net22290), .CLK(net22295), .Q(conv_weight_box[72]) );
  DFFSSRX1_HVT conv_weight_box_reg_32__3_ ( .D(1'b0), .SETB(n15), .RSTB(
        net22291), .CLK(net22295), .Q(conv_weight_box[71]) );
  DFFSSRX1_HVT conv_weight_box_reg_32__2_ ( .D(1'b0), .SETB(n10), .RSTB(
        net22292), .CLK(net22295), .Q(conv_weight_box[70]) );
  DFFSSRX1_HVT conv_weight_box_reg_32__1_ ( .D(1'b0), .SETB(n5), .RSTB(
        net22300), .CLK(net22312), .Q(conv_weight_box[69]) );
  DFFSSRX1_HVT conv_weight_box_reg_32__0_ ( .D(1'b0), .SETB(n16), .RSTB(
        net22301), .CLK(net22312), .Q(conv_weight_box[68]) );
  DFFSSRX1_HVT conv_weight_box_reg_33__3_ ( .D(1'b0), .SETB(n11), .RSTB(
        net22302), .CLK(net22312), .Q(conv_weight_box[67]) );
  DFFSSRX1_HVT conv_weight_box_reg_33__2_ ( .D(1'b0), .SETB(n6), .RSTB(
        net22303), .CLK(net22312), .Q(conv_weight_box[66]) );
  DFFSSRX1_HVT conv_weight_box_reg_33__1_ ( .D(1'b0), .SETB(n17), .RSTB(
        net22304), .CLK(net22312), .Q(conv_weight_box[65]) );
  DFFSSRX1_HVT conv_weight_box_reg_33__0_ ( .D(1'b0), .SETB(n12), .RSTB(
        net22305), .CLK(net22312), .Q(conv_weight_box[64]) );
  DFFSSRX1_HVT conv_weight_box_reg_34__3_ ( .D(1'b0), .SETB(n7), .RSTB(
        net22306), .CLK(net22312), .Q(conv_weight_box[63]) );
  DFFSSRX1_HVT conv_weight_box_reg_34__2_ ( .D(1'b0), .SETB(n14), .RSTB(
        net22307), .CLK(net22312), .Q(conv_weight_box[62]) );
  DFFSSRX1_HVT conv_weight_box_reg_34__1_ ( .D(1'b0), .SETB(n9), .RSTB(
        net22308), .CLK(net22312), .Q(conv_weight_box[61]) );
  DFFSSRX1_HVT conv_weight_box_reg_34__0_ ( .D(1'b0), .SETB(n4), .RSTB(
        net22309), .CLK(net22312), .Q(conv_weight_box[60]) );
  DFFSSRX1_HVT conv_weight_box_reg_35__3_ ( .D(1'b0), .SETB(n15), .RSTB(
        net22317), .CLK(net22329), .Q(conv_weight_box[59]) );
  DFFSSRX1_HVT conv_weight_box_reg_35__2_ ( .D(1'b0), .SETB(n10), .RSTB(
        net22318), .CLK(net22329), .Q(conv_weight_box[58]) );
  DFFSSRX1_HVT conv_weight_box_reg_35__1_ ( .D(1'b0), .SETB(n5), .RSTB(
        net22319), .CLK(net22329), .Q(conv_weight_box[57]) );
  DFFSSRX1_HVT conv_weight_box_reg_35__0_ ( .D(1'b0), .SETB(n16), .RSTB(
        net22320), .CLK(net22329), .Q(conv_weight_box[56]) );
  DFFSSRX1_HVT conv_weight_box_reg_36__3_ ( .D(1'b0), .SETB(n11), .RSTB(
        net22321), .CLK(net22329), .Q(conv_weight_box[55]) );
  DFFSSRX1_HVT conv_weight_box_reg_36__2_ ( .D(1'b0), .SETB(n6), .RSTB(
        net22322), .CLK(net22329), .Q(conv_weight_box[54]) );
  DFFSSRX1_HVT conv_weight_box_reg_36__1_ ( .D(1'b0), .SETB(n17), .RSTB(
        net22323), .CLK(net22329), .Q(conv_weight_box[53]) );
  DFFSSRX1_HVT conv_weight_box_reg_36__0_ ( .D(1'b0), .SETB(n12), .RSTB(
        net22324), .CLK(net22329), .Q(conv_weight_box[52]) );
  DFFSSRX1_HVT conv_weight_box_reg_37__3_ ( .D(1'b0), .SETB(n7), .RSTB(
        net22325), .CLK(net22329), .Q(conv_weight_box[51]) );
  DFFSSRX1_HVT conv_weight_box_reg_37__2_ ( .D(1'b0), .SETB(n14), .RSTB(
        net22326), .CLK(net22329), .Q(conv_weight_box[50]) );
  DFFSSRX1_HVT conv_weight_box_reg_37__1_ ( .D(1'b0), .SETB(n9), .RSTB(
        net22334), .CLK(net22346), .Q(conv_weight_box[49]) );
  DFFSSRX1_HVT conv_weight_box_reg_37__0_ ( .D(1'b0), .SETB(n4), .RSTB(
        net22335), .CLK(net22346), .Q(conv_weight_box[48]) );
  DFFSSRX1_HVT conv_weight_box_reg_38__3_ ( .D(1'b0), .SETB(n15), .RSTB(
        net22336), .CLK(net22346), .Q(conv_weight_box[47]) );
  DFFSSRX1_HVT conv_weight_box_reg_38__2_ ( .D(1'b0), .SETB(n10), .RSTB(
        net22337), .CLK(net22346), .Q(conv_weight_box[46]) );
  DFFSSRX1_HVT conv_weight_box_reg_38__1_ ( .D(1'b0), .SETB(n5), .RSTB(
        net22338), .CLK(net22346), .Q(conv_weight_box[45]) );
  DFFSSRX1_HVT conv_weight_box_reg_38__0_ ( .D(1'b0), .SETB(n16), .RSTB(
        net22339), .CLK(net22346), .Q(conv_weight_box[44]) );
  DFFSSRX1_HVT conv_weight_box_reg_39__3_ ( .D(1'b0), .SETB(n11), .RSTB(
        net22340), .CLK(net22346), .Q(conv_weight_box[43]) );
  DFFSSRX1_HVT conv_weight_box_reg_39__2_ ( .D(1'b0), .SETB(n6), .RSTB(
        net22341), .CLK(net22346), .Q(conv_weight_box[42]) );
  DFFSSRX1_HVT conv_weight_box_reg_39__1_ ( .D(1'b0), .SETB(n17), .RSTB(
        net22342), .CLK(net22346), .Q(conv_weight_box[41]) );
  DFFSSRX1_HVT conv_weight_box_reg_39__0_ ( .D(1'b0), .SETB(n12), .RSTB(
        net22343), .CLK(net22346), .Q(conv_weight_box[40]) );
  DFFSSRX1_HVT conv_weight_box_reg_40__3_ ( .D(1'b0), .SETB(n7), .RSTB(
        net22351), .CLK(net22363), .Q(conv_weight_box[39]) );
  DFFSSRX1_HVT conv_weight_box_reg_40__2_ ( .D(1'b0), .SETB(n14), .RSTB(
        net22352), .CLK(net22363), .Q(conv_weight_box[38]) );
  DFFSSRX1_HVT conv_weight_box_reg_40__1_ ( .D(1'b0), .SETB(n9), .RSTB(
        net22353), .CLK(net22363), .Q(conv_weight_box[37]) );
  DFFSSRX1_HVT conv_weight_box_reg_40__0_ ( .D(1'b0), .SETB(n4), .RSTB(
        net22354), .CLK(net22363), .Q(conv_weight_box[36]) );
  DFFSSRX1_HVT conv_weight_box_reg_41__3_ ( .D(1'b0), .SETB(n15), .RSTB(
        net22355), .CLK(net22363), .Q(conv_weight_box[35]) );
  DFFSSRX1_HVT conv_weight_box_reg_41__2_ ( .D(1'b0), .SETB(n10), .RSTB(
        net22356), .CLK(net22363), .Q(conv_weight_box[34]) );
  DFFSSRX1_HVT conv_weight_box_reg_41__1_ ( .D(1'b0), .SETB(n5), .RSTB(
        net22357), .CLK(net22363), .Q(conv_weight_box[33]) );
  DFFSSRX1_HVT conv_weight_box_reg_41__0_ ( .D(1'b0), .SETB(n16), .RSTB(
        net22358), .CLK(net22363), .Q(conv_weight_box[32]) );
  DFFSSRX1_HVT conv_weight_box_reg_42__3_ ( .D(1'b0), .SETB(n11), .RSTB(
        net22359), .CLK(net22363), .Q(conv_weight_box[31]) );
  DFFSSRX1_HVT conv_weight_box_reg_42__2_ ( .D(1'b0), .SETB(n6), .RSTB(
        net22360), .CLK(net22363), .Q(conv_weight_box[30]) );
  DFFSSRX1_HVT conv_weight_box_reg_42__1_ ( .D(1'b0), .SETB(n17), .RSTB(
        net22368), .CLK(net22380), .Q(conv_weight_box[29]) );
  DFFSSRX1_HVT conv_weight_box_reg_42__0_ ( .D(1'b0), .SETB(n12), .RSTB(
        net22369), .CLK(net22380), .Q(conv_weight_box[28]) );
  DFFSSRX1_HVT conv_weight_box_reg_43__3_ ( .D(1'b0), .SETB(n7), .RSTB(
        net22370), .CLK(net22380), .Q(conv_weight_box[27]) );
  DFFSSRX1_HVT conv_weight_box_reg_43__2_ ( .D(1'b0), .SETB(n14), .RSTB(
        net22371), .CLK(net22380), .Q(conv_weight_box[26]) );
  DFFSSRX1_HVT conv_weight_box_reg_43__1_ ( .D(1'b0), .SETB(n9), .RSTB(
        net22372), .CLK(net22380), .Q(conv_weight_box[25]) );
  DFFSSRX1_HVT conv_weight_box_reg_43__0_ ( .D(1'b0), .SETB(n4), .RSTB(
        net22373), .CLK(net22380), .Q(conv_weight_box[24]) );
  DFFSSRX1_HVT conv_weight_box_reg_44__3_ ( .D(1'b0), .SETB(n15), .RSTB(
        net22374), .CLK(net22380), .Q(conv_weight_box[23]) );
  DFFSSRX1_HVT conv_weight_box_reg_44__2_ ( .D(1'b0), .SETB(n10), .RSTB(
        net22375), .CLK(net22380), .Q(conv_weight_box[22]) );
  DFFSSRX1_HVT conv_weight_box_reg_44__1_ ( .D(1'b0), .SETB(n5), .RSTB(
        net22376), .CLK(net22380), .Q(conv_weight_box[21]) );
  DFFSSRX1_HVT conv_weight_box_reg_44__0_ ( .D(1'b0), .SETB(n16), .RSTB(
        net22377), .CLK(net22380), .Q(conv_weight_box[20]) );
  DFFSSRX1_HVT conv_weight_box_reg_45__3_ ( .D(1'b0), .SETB(n11), .RSTB(
        net22385), .CLK(net22397), .Q(conv_weight_box[19]) );
  DFFSSRX1_HVT conv_weight_box_reg_45__2_ ( .D(1'b0), .SETB(n6), .RSTB(
        net22386), .CLK(net22397), .Q(conv_weight_box[18]) );
  DFFSSRX1_HVT conv_weight_box_reg_45__1_ ( .D(1'b0), .SETB(n17), .RSTB(
        net22387), .CLK(net22397), .Q(conv_weight_box[17]) );
  DFFSSRX1_HVT conv_weight_box_reg_45__0_ ( .D(1'b0), .SETB(n12), .RSTB(
        net22388), .CLK(net22397), .Q(conv_weight_box[16]) );
  DFFSSRX1_HVT conv_weight_box_reg_46__3_ ( .D(1'b0), .SETB(n7), .RSTB(
        net22389), .CLK(net22397), .Q(conv_weight_box[15]) );
  DFFSSRX1_HVT conv_weight_box_reg_46__2_ ( .D(1'b0), .SETB(n14), .RSTB(
        net22390), .CLK(net22397), .Q(conv_weight_box[14]) );
  DFFSSRX1_HVT conv_weight_box_reg_46__1_ ( .D(1'b0), .SETB(n9), .RSTB(
        net22391), .CLK(net22397), .Q(conv_weight_box[13]) );
  DFFSSRX1_HVT conv_weight_box_reg_46__0_ ( .D(1'b0), .SETB(n4), .RSTB(
        net22392), .CLK(net22397), .Q(conv_weight_box[12]) );
  DFFSSRX1_HVT conv_weight_box_reg_47__3_ ( .D(1'b0), .SETB(n15), .RSTB(
        net22393), .CLK(net22397), .Q(conv_weight_box[11]) );
  DFFSSRX1_HVT conv_weight_box_reg_47__2_ ( .D(1'b0), .SETB(n10), .RSTB(
        net22394), .CLK(net22397), .Q(conv_weight_box[10]) );
  DFFSSRX1_HVT conv_weight_box_reg_47__1_ ( .D(1'b0), .SETB(n5), .RSTB(
        net22402), .CLK(net22414), .Q(conv_weight_box[9]) );
  DFFSSRX1_HVT conv_weight_box_reg_47__0_ ( .D(1'b0), .SETB(n16), .RSTB(
        net22403), .CLK(net22414), .Q(conv_weight_box[8]) );
  DFFSSRX1_HVT conv_weight_box_reg_48__3_ ( .D(1'b0), .SETB(n11), .RSTB(
        net22404), .CLK(net22414), .Q(conv_weight_box[7]) );
  DFFSSRX1_HVT conv_weight_box_reg_48__2_ ( .D(1'b0), .SETB(n6), .RSTB(
        net22405), .CLK(net22414), .Q(conv_weight_box[6]) );
  DFFSSRX1_HVT conv_weight_box_reg_48__1_ ( .D(1'b0), .SETB(n17), .RSTB(
        net22406), .CLK(net22414), .Q(conv_weight_box[5]) );
  DFFSSRX1_HVT conv_weight_box_reg_48__0_ ( .D(1'b0), .SETB(n12), .RSTB(
        net22407), .CLK(net22414), .Q(conv_weight_box[4]) );
  DFFSSRX1_HVT conv_weight_box_reg_49__3_ ( .D(1'b0), .SETB(n7), .RSTB(
        net22408), .CLK(net22414), .Q(conv_weight_box[3]) );
  DFFSSRX1_HVT conv_weight_box_reg_49__2_ ( .D(1'b0), .SETB(n14), .RSTB(
        net22409), .CLK(net22414), .Q(conv_weight_box[2]) );
  DFFSSRX1_HVT conv_weight_box_reg_49__1_ ( .D(1'b0), .SETB(n9), .RSTB(
        net22410), .CLK(net22414), .Q(conv_weight_box[1]) );
  DFFSSRX1_HVT conv_weight_box_reg_49__0_ ( .D(1'b0), .SETB(n4), .RSTB(
        net22411), .CLK(net22414), .Q(conv_weight_box[0]) );
  DFFSSRX1_HVT bias_data_reg_3_ ( .D(1'b0), .SETB(n15), .RSTB(net22431), .CLK(
        net22446), .Q(bias_data[3]) );
  DFFSSRX1_HVT bias_data_reg_2_ ( .D(1'b0), .SETB(n10), .RSTB(net22435), .CLK(
        net22446), .Q(bias_data[2]) );
  DFFSSRX1_HVT bias_data_reg_1_ ( .D(1'b0), .SETB(n5), .RSTB(net22439), .CLK(
        net22446), .Q(bias_data[1]) );
  DFFSSRX1_HVT bias_data_reg_0_ ( .D(1'b0), .SETB(n16), .RSTB(net22443), .CLK(
        net22446), .Q(bias_data[0]) );
  NOR3X0_HVT U3 ( .A1(n90), .A2(load_conv2_bias1_enable), .A3(
        load_conv2_bias0_enable), .Y(n28) );
  INVX1_HVT U4 ( .A(srstn), .Y(n26) );
  INVX0_HVT U5 ( .A(n42), .Y(n19) );
  NAND2X0_HVT U6 ( .A1(load_conv2_bias1_enable), .A2(n40), .Y(n42) );
  INVX1_HVT U7 ( .A(mode[1]), .Y(n38) );
  INVX1_HVT U8 ( .A(n349), .Y(n115) );
  INVX1_HVT U9 ( .A(n285), .Y(n68) );
  INVX1_HVT U10 ( .A(set_4_), .Y(n106) );
  INVX1_HVT U11 ( .A(set_2_), .Y(n105) );
  INVX1_HVT U12 ( .A(set_0_), .Y(n113) );
  INVX1_HVT U13 ( .A(n22), .Y(n2) );
  NOR2X1_HVT U14 ( .A1(load_conv1_bias_enable), .A2(n43), .Y(n27) );
  INVX1_HVT U15 ( .A(n26), .Y(n13) );
  INVX1_HVT U16 ( .A(n26), .Y(n8) );
  INVX0_HVT U17 ( .A(n287), .Y(n65) );
  INVX0_HVT U18 ( .A(n351), .Y(n112) );
  INVX0_HVT U19 ( .A(set_1_), .Y(n99) );
  INVX1_HVT U20 ( .A(n42), .Y(n3) );
  INVX2_HVT U21 ( .A(n13), .Y(n4) );
  INVX2_HVT U22 ( .A(n8), .Y(n5) );
  INVX2_HVT U23 ( .A(n8), .Y(n6) );
  INVX2_HVT U24 ( .A(n13), .Y(n7) );
  INVX2_HVT U25 ( .A(n8), .Y(n9) );
  INVX2_HVT U26 ( .A(n8), .Y(n10) );
  INVX2_HVT U27 ( .A(n8), .Y(n11) );
  INVX2_HVT U28 ( .A(n8), .Y(n12) );
  INVX2_HVT U29 ( .A(n13), .Y(n14) );
  INVX2_HVT U30 ( .A(n13), .Y(n15) );
  INVX2_HVT U31 ( .A(n13), .Y(n16) );
  INVX2_HVT U32 ( .A(n13), .Y(n17) );
  INVX2_HVT U33 ( .A(n42), .Y(n18) );
  INVX2_HVT U34 ( .A(n42), .Y(n20) );
  INVX2_HVT U35 ( .A(n42), .Y(n21) );
  INVX1_HVT U36 ( .A(n39), .Y(n22) );
  INVX2_HVT U37 ( .A(n22), .Y(n23) );
  INVX2_HVT U38 ( .A(n22), .Y(n24) );
  INVX2_HVT U39 ( .A(n22), .Y(n25) );
  OR2X4_HVT U40 ( .A1(n38), .A2(mode[0]), .Y(n90) );
  INVX1_HVT U41 ( .A(n90), .Y(n40) );
  AO22X2_HVT U42 ( .A1(n40), .A2(load_conv2_bias0_enable), .A3(mode[0]), .A4(
        n38), .Y(n39) );
  NOR4X1_HVT U43 ( .A1(n255), .A2(n254), .A3(n253), .A4(n252), .Y(n275) );
  NOR4X1_HVT U44 ( .A1(n249), .A2(n248), .A3(n247), .A4(n246), .Y(n250) );
  NOR4X1_HVT U45 ( .A1(n245), .A2(n244), .A3(n243), .A4(n242), .Y(n251) );
  NOR4X1_HVT U46 ( .A1(n220), .A2(n219), .A3(n218), .A4(n217), .Y(n240) );
  NOR4X1_HVT U47 ( .A1(n214), .A2(n213), .A3(n212), .A4(n211), .Y(n215) );
  NOR4X1_HVT U48 ( .A1(n210), .A2(n209), .A3(n208), .A4(n207), .Y(n216) );
  NOR4X1_HVT U49 ( .A1(n185), .A2(n184), .A3(n183), .A4(n182), .Y(n205) );
  NOR4X1_HVT U50 ( .A1(n179), .A2(n178), .A3(n177), .A4(n176), .Y(n180) );
  NOR4X1_HVT U51 ( .A1(n175), .A2(n174), .A3(n173), .A4(n172), .Y(n181) );
  NOR4X1_HVT U52 ( .A1(n150), .A2(n149), .A3(n148), .A4(n147), .Y(n170) );
  NOR4X1_HVT U53 ( .A1(n144), .A2(n143), .A3(n142), .A4(n141), .Y(n145) );
  NOR4X1_HVT U54 ( .A1(n140), .A2(n139), .A3(n138), .A4(n137), .Y(n146) );
  NOR4X1_HVT U55 ( .A1(n364), .A2(n363), .A3(n362), .A4(n361), .Y(n402) );
  NOR4X1_HVT U56 ( .A1(n348), .A2(n347), .A3(n346), .A4(n345), .Y(n350) );
  NOR4X1_HVT U57 ( .A1(n344), .A2(n343), .A3(n342), .A4(n341), .Y(n352) );
  NOR4X1_HVT U58 ( .A1(n300), .A2(n299), .A3(n298), .A4(n297), .Y(n339) );
  NOR4X1_HVT U59 ( .A1(n284), .A2(n283), .A3(n282), .A4(n281), .Y(n286) );
  NOR4X1_HVT U60 ( .A1(n280), .A2(n279), .A3(n278), .A4(n277), .Y(n288) );
  NOR4X1_HVT U61 ( .A1(n110), .A2(n109), .A3(n108), .A4(n107), .Y(n135) );
  NOR4X1_HVT U62 ( .A1(n98), .A2(n97), .A3(n96), .A4(n95), .Y(n100) );
  NOR4X1_HVT U63 ( .A1(n94), .A2(n93), .A3(n92), .A4(n91), .Y(n101) );
  AND2X1_HVT U64 ( .A1(set_4_), .A2(n111), .Y(n388) );
  AND3X1_HVT U65 ( .A1(set_3_), .A2(set_4_), .A3(n105), .Y(n389) );
  AND2X1_HVT U66 ( .A1(set_5_), .A2(n111), .Y(n386) );
  AND3X1_HVT U67 ( .A1(set_2_), .A2(set_4_), .A3(n104), .Y(n387) );
  AND3X1_HVT U68 ( .A1(set_5_), .A2(set_3_), .A3(n105), .Y(n383) );
  INVX1_HVT U69 ( .A(set_5_), .Y(n114) );
  AND3X1_HVT U70 ( .A1(set_2_), .A2(set_5_), .A3(n104), .Y(n381) );
  INVX1_HVT U71 ( .A(set_3_), .Y(n104) );
  NOR4X1_HVT U72 ( .A1(n63), .A2(n62), .A3(n61), .A4(n60), .Y(n88) );
  NOR4X1_HVT U73 ( .A1(n51), .A2(n50), .A3(n49), .A4(n48), .Y(n53) );
  INVX1_HVT U74 ( .A(conv1_bias_set_1_), .Y(n52) );
  NOR4X1_HVT U75 ( .A1(n47), .A2(n46), .A3(n45), .A4(n44), .Y(n54) );
  AND2X1_HVT U76 ( .A1(conv1_bias_set_4_), .A2(n64), .Y(n325) );
  AND3X1_HVT U77 ( .A1(conv1_bias_set_3_), .A2(conv1_bias_set_4_), .A3(n58), 
        .Y(n326) );
  AND2X1_HVT U78 ( .A1(conv1_bias_set_5_), .A2(n64), .Y(n323) );
  AND3X1_HVT U79 ( .A1(conv1_bias_set_2_), .A2(conv1_bias_set_4_), .A3(n57), 
        .Y(n324) );
  AND3X1_HVT U80 ( .A1(conv1_bias_set_5_), .A2(conv1_bias_set_3_), .A3(n58), 
        .Y(n320) );
  INVX1_HVT U81 ( .A(conv1_bias_set_2_), .Y(n58) );
  INVX1_HVT U82 ( .A(conv1_bias_set_4_), .Y(n59) );
  INVX1_HVT U83 ( .A(conv1_bias_set_5_), .Y(n67) );
  AND3X1_HVT U84 ( .A1(conv1_bias_set_2_), .A2(conv1_bias_set_5_), .A3(n57), 
        .Y(n318) );
  INVX1_HVT U85 ( .A(conv1_bias_set_3_), .Y(n57) );
  INVX1_HVT U86 ( .A(conv1_bias_set_0_), .Y(n66) );
  NAND2X0_HVT U87 ( .A1(srstn), .A2(n37), .Y(net22223) );
  INVX1_HVT U88 ( .A(load_conv2_bias0_enable), .Y(n41) );
  NAND4X0_HVT U89 ( .A1(n337), .A2(n340), .A3(n339), .A4(n338), .Y(n30) );
  NAND4X0_HVT U90 ( .A1(n400), .A2(n403), .A3(n402), .A4(n401), .Y(n29) );
  AO22X1_HVT U91 ( .A1(n30), .A2(n27), .A3(n28), .A4(n29), .Y(net22443) );
  NAND4X0_HVT U92 ( .A1(n238), .A2(n241), .A3(n240), .A4(n239), .Y(n32) );
  NAND4X0_HVT U93 ( .A1(n273), .A2(n276), .A3(n275), .A4(n274), .Y(n31) );
  AO22X1_HVT U94 ( .A1(n32), .A2(n27), .A3(n28), .A4(n31), .Y(net22439) );
  NAND4X0_HVT U95 ( .A1(n168), .A2(n171), .A3(n170), .A4(n169), .Y(n34) );
  NAND4X0_HVT U96 ( .A1(n203), .A2(n206), .A3(n205), .A4(n204), .Y(n33) );
  AO22X1_HVT U97 ( .A1(n34), .A2(n27), .A3(n28), .A4(n33), .Y(net22435) );
  NAND4X0_HVT U98 ( .A1(n86), .A2(n89), .A3(n88), .A4(n87), .Y(n36) );
  NAND4X0_HVT U99 ( .A1(n133), .A2(n136), .A3(n135), .A4(n134), .Y(n35) );
  AO22X1_HVT U100 ( .A1(n36), .A2(n27), .A3(n28), .A4(n35), .Y(net22431) );
  NAND2X0_HVT U101 ( .A1(mode[0]), .A2(n38), .Y(n43) );
  AO221X1_HVT U102 ( .A1(n40), .A2(n41), .A3(n90), .A4(n43), .A5(n27), .Y(n37)
         );
  AND2X1_HVT U103 ( .A1(delay_weight[99]), .A2(n25), .Y(net22069) );
  AND2X1_HVT U104 ( .A1(delay_weight[98]), .A2(n39), .Y(net22072) );
  AND2X1_HVT U105 ( .A1(delay_weight[97]), .A2(n25), .Y(net22073) );
  AND2X1_HVT U106 ( .A1(delay_weight[96]), .A2(n24), .Y(net22074) );
  AND2X1_HVT U107 ( .A1(delay_weight[95]), .A2(n23), .Y(net22075) );
  AND2X1_HVT U108 ( .A1(delay_weight[94]), .A2(n24), .Y(net22076) );
  AND2X1_HVT U109 ( .A1(delay_weight[93]), .A2(n2), .Y(net22077) );
  AND2X1_HVT U110 ( .A1(delay_weight[92]), .A2(n24), .Y(net22078) );
  AND2X1_HVT U111 ( .A1(delay_weight[91]), .A2(n23), .Y(net22079) );
  AND2X1_HVT U112 ( .A1(delay_weight[90]), .A2(n23), .Y(net22080) );
  AND2X1_HVT U113 ( .A1(delay_weight[89]), .A2(n24), .Y(net22088) );
  AND2X1_HVT U114 ( .A1(delay_weight[88]), .A2(n25), .Y(net22089) );
  AND2X1_HVT U115 ( .A1(delay_weight[87]), .A2(n24), .Y(net22090) );
  AND2X1_HVT U116 ( .A1(delay_weight[86]), .A2(n25), .Y(net22091) );
  AND2X1_HVT U117 ( .A1(delay_weight[85]), .A2(n39), .Y(net22092) );
  AND2X1_HVT U118 ( .A1(delay_weight[84]), .A2(n23), .Y(net22093) );
  AND2X1_HVT U119 ( .A1(delay_weight[83]), .A2(n23), .Y(net22094) );
  AND2X1_HVT U120 ( .A1(delay_weight[82]), .A2(n23), .Y(net22095) );
  AND2X1_HVT U121 ( .A1(delay_weight[81]), .A2(n2), .Y(net22096) );
  AND2X1_HVT U122 ( .A1(delay_weight[80]), .A2(n24), .Y(net22097) );
  AND2X1_HVT U123 ( .A1(delay_weight[79]), .A2(n25), .Y(net22105) );
  AND2X1_HVT U124 ( .A1(delay_weight[78]), .A2(n25), .Y(net22106) );
  AND2X1_HVT U125 ( .A1(delay_weight[77]), .A2(n39), .Y(net22107) );
  AND2X1_HVT U126 ( .A1(delay_weight[76]), .A2(n24), .Y(net22108) );
  AND2X1_HVT U127 ( .A1(delay_weight[75]), .A2(n23), .Y(net22109) );
  AND2X1_HVT U128 ( .A1(delay_weight[74]), .A2(n2), .Y(net22110) );
  AND2X1_HVT U129 ( .A1(delay_weight[73]), .A2(n2), .Y(net22111) );
  AND2X1_HVT U130 ( .A1(delay_weight[72]), .A2(n25), .Y(net22112) );
  AND2X1_HVT U131 ( .A1(delay_weight[71]), .A2(n25), .Y(net22113) );
  AND2X1_HVT U132 ( .A1(delay_weight[70]), .A2(n25), .Y(net22114) );
  AND2X1_HVT U133 ( .A1(delay_weight[69]), .A2(n39), .Y(net22122) );
  AND2X1_HVT U134 ( .A1(delay_weight[68]), .A2(n23), .Y(net22123) );
  AND2X1_HVT U135 ( .A1(delay_weight[67]), .A2(n39), .Y(net22124) );
  AND2X1_HVT U136 ( .A1(delay_weight[66]), .A2(n24), .Y(net22125) );
  AND2X1_HVT U137 ( .A1(delay_weight[65]), .A2(n23), .Y(net22126) );
  AND2X1_HVT U138 ( .A1(delay_weight[64]), .A2(n23), .Y(net22127) );
  AND2X1_HVT U139 ( .A1(delay_weight[63]), .A2(n25), .Y(net22128) );
  AND2X1_HVT U140 ( .A1(delay_weight[62]), .A2(n24), .Y(net22129) );
  AND2X1_HVT U141 ( .A1(delay_weight[61]), .A2(n2), .Y(net22130) );
  AND2X1_HVT U142 ( .A1(delay_weight[60]), .A2(n24), .Y(net22131) );
  AND2X1_HVT U143 ( .A1(delay_weight[59]), .A2(n25), .Y(net22139) );
  AND2X1_HVT U144 ( .A1(delay_weight[58]), .A2(n24), .Y(net22140) );
  AND2X1_HVT U145 ( .A1(delay_weight[57]), .A2(n2), .Y(net22141) );
  AND2X1_HVT U146 ( .A1(delay_weight[56]), .A2(n23), .Y(net22142) );
  AND2X1_HVT U147 ( .A1(delay_weight[55]), .A2(n39), .Y(net22143) );
  AND2X1_HVT U148 ( .A1(delay_weight[54]), .A2(n23), .Y(net22144) );
  AND2X1_HVT U149 ( .A1(delay_weight[53]), .A2(n39), .Y(net22145) );
  AND2X1_HVT U150 ( .A1(delay_weight[52]), .A2(n25), .Y(net22146) );
  AND2X1_HVT U151 ( .A1(delay_weight[51]), .A2(n24), .Y(net22147) );
  AND2X1_HVT U152 ( .A1(delay_weight[50]), .A2(n39), .Y(net22148) );
  AND2X1_HVT U153 ( .A1(delay_weight[49]), .A2(n39), .Y(net22156) );
  AND2X1_HVT U154 ( .A1(delay_weight[48]), .A2(n23), .Y(net22157) );
  AND2X1_HVT U155 ( .A1(delay_weight[47]), .A2(n24), .Y(net22158) );
  AND2X1_HVT U156 ( .A1(delay_weight[46]), .A2(n23), .Y(net22159) );
  AND2X1_HVT U157 ( .A1(delay_weight[45]), .A2(n2), .Y(net22160) );
  AND2X1_HVT U158 ( .A1(delay_weight[44]), .A2(n25), .Y(net22161) );
  AND2X1_HVT U159 ( .A1(delay_weight[43]), .A2(n39), .Y(net22162) );
  AND2X1_HVT U160 ( .A1(delay_weight[42]), .A2(n25), .Y(net22163) );
  AND2X1_HVT U161 ( .A1(delay_weight[41]), .A2(n25), .Y(net22164) );
  AND2X1_HVT U162 ( .A1(delay_weight[40]), .A2(n24), .Y(net22165) );
  AND2X1_HVT U163 ( .A1(delay_weight[39]), .A2(n23), .Y(net22173) );
  AND2X1_HVT U164 ( .A1(delay_weight[38]), .A2(n23), .Y(net22174) );
  AND2X1_HVT U165 ( .A1(delay_weight[37]), .A2(n2), .Y(net22175) );
  AND2X1_HVT U166 ( .A1(delay_weight[36]), .A2(n25), .Y(net22176) );
  AND2X1_HVT U167 ( .A1(delay_weight[35]), .A2(n24), .Y(net22177) );
  AND2X1_HVT U168 ( .A1(delay_weight[34]), .A2(n25), .Y(net22178) );
  AND2X1_HVT U169 ( .A1(delay_weight[33]), .A2(n39), .Y(net22179) );
  AND2X1_HVT U170 ( .A1(delay_weight[32]), .A2(n25), .Y(net22180) );
  AND2X1_HVT U171 ( .A1(delay_weight[31]), .A2(n39), .Y(net22181) );
  AND2X1_HVT U172 ( .A1(delay_weight[30]), .A2(n24), .Y(net22182) );
  AND2X1_HVT U173 ( .A1(delay_weight[29]), .A2(n2), .Y(net22190) );
  AND2X1_HVT U174 ( .A1(delay_weight[28]), .A2(n23), .Y(net22191) );
  AND2X1_HVT U175 ( .A1(delay_weight[27]), .A2(n25), .Y(net22192) );
  AND2X1_HVT U176 ( .A1(delay_weight[26]), .A2(n39), .Y(net22193) );
  AND2X1_HVT U177 ( .A1(delay_weight[25]), .A2(n39), .Y(net22194) );
  AND2X1_HVT U178 ( .A1(delay_weight[24]), .A2(n24), .Y(net22195) );
  AND2X1_HVT U179 ( .A1(delay_weight[23]), .A2(n23), .Y(net22196) );
  AND2X1_HVT U180 ( .A1(delay_weight[22]), .A2(n24), .Y(net22197) );
  AND2X1_HVT U181 ( .A1(delay_weight[21]), .A2(n2), .Y(net22198) );
  AND2X1_HVT U182 ( .A1(delay_weight[20]), .A2(n24), .Y(net22199) );
  AND2X1_HVT U183 ( .A1(delay_weight[19]), .A2(n39), .Y(net22207) );
  AND2X1_HVT U184 ( .A1(delay_weight[18]), .A2(n23), .Y(net22208) );
  AND2X1_HVT U185 ( .A1(delay_weight[17]), .A2(n24), .Y(net22209) );
  AND2X1_HVT U186 ( .A1(delay_weight[16]), .A2(n25), .Y(net22210) );
  AND2X1_HVT U187 ( .A1(delay_weight[15]), .A2(n24), .Y(net22211) );
  AND2X1_HVT U188 ( .A1(delay_weight[14]), .A2(n25), .Y(net22212) );
  AND2X1_HVT U189 ( .A1(delay_weight[13]), .A2(n39), .Y(net22213) );
  AND2X1_HVT U190 ( .A1(delay_weight[12]), .A2(n23), .Y(net22214) );
  AND2X1_HVT U191 ( .A1(delay_weight[11]), .A2(n23), .Y(net22215) );
  AND2X1_HVT U192 ( .A1(delay_weight[10]), .A2(n23), .Y(net22216) );
  AND2X1_HVT U193 ( .A1(delay_weight[9]), .A2(n39), .Y(net22224) );
  AND2X1_HVT U194 ( .A1(delay_weight[8]), .A2(n24), .Y(net22225) );
  AND2X1_HVT U195 ( .A1(delay_weight[7]), .A2(n39), .Y(net22226) );
  AND2X1_HVT U196 ( .A1(delay_weight[6]), .A2(n25), .Y(net22227) );
  AND2X1_HVT U197 ( .A1(delay_weight[5]), .A2(n39), .Y(net22228) );
  AND2X1_HVT U198 ( .A1(delay_weight[4]), .A2(n24), .Y(net22229) );
  AND2X1_HVT U199 ( .A1(delay_weight[3]), .A2(n23), .Y(net22230) );
  AND2X1_HVT U200 ( .A1(delay_weight[2]), .A2(n2), .Y(net22231) );
  AND2X1_HVT U201 ( .A1(delay_weight[1]), .A2(n2), .Y(net22232) );
  AND2X1_HVT U202 ( .A1(delay_weight[0]), .A2(n25), .Y(net22233) );
  AO21X1_HVT U203 ( .A1(n3), .A2(n41), .A3(n26), .Y(net22401) );
  AND2X1_HVT U204 ( .A1(delay_weight[99]), .A2(n20), .Y(net22249) );
  AND2X1_HVT U205 ( .A1(delay_weight[98]), .A2(n20), .Y(net22250) );
  AND2X1_HVT U206 ( .A1(delay_weight[97]), .A2(n19), .Y(net22251) );
  AND2X1_HVT U207 ( .A1(delay_weight[96]), .A2(n21), .Y(net22252) );
  AND2X1_HVT U208 ( .A1(delay_weight[95]), .A2(n3), .Y(net22253) );
  AND2X1_HVT U209 ( .A1(delay_weight[94]), .A2(n18), .Y(net22254) );
  AND2X1_HVT U210 ( .A1(delay_weight[93]), .A2(n21), .Y(net22255) );
  AND2X1_HVT U211 ( .A1(delay_weight[92]), .A2(n18), .Y(net22256) );
  AND2X1_HVT U212 ( .A1(delay_weight[91]), .A2(n21), .Y(net22257) );
  AND2X1_HVT U213 ( .A1(delay_weight[90]), .A2(n21), .Y(net22258) );
  AND2X1_HVT U214 ( .A1(delay_weight[89]), .A2(n21), .Y(net22266) );
  AND2X1_HVT U215 ( .A1(delay_weight[88]), .A2(n18), .Y(net22267) );
  AND2X1_HVT U216 ( .A1(delay_weight[87]), .A2(n18), .Y(net22268) );
  AND2X1_HVT U217 ( .A1(delay_weight[86]), .A2(n3), .Y(net22269) );
  AND2X1_HVT U218 ( .A1(delay_weight[85]), .A2(n20), .Y(net22270) );
  AND2X1_HVT U219 ( .A1(delay_weight[84]), .A2(n18), .Y(net22271) );
  AND2X1_HVT U220 ( .A1(delay_weight[83]), .A2(n20), .Y(net22272) );
  AND2X1_HVT U221 ( .A1(delay_weight[82]), .A2(n19), .Y(net22273) );
  AND2X1_HVT U222 ( .A1(delay_weight[81]), .A2(n18), .Y(net22274) );
  AND2X1_HVT U223 ( .A1(delay_weight[80]), .A2(n18), .Y(net22275) );
  AND2X1_HVT U224 ( .A1(delay_weight[79]), .A2(n20), .Y(net22283) );
  AND2X1_HVT U225 ( .A1(delay_weight[78]), .A2(n19), .Y(net22284) );
  AND2X1_HVT U226 ( .A1(delay_weight[77]), .A2(n3), .Y(net22285) );
  AND2X1_HVT U227 ( .A1(delay_weight[76]), .A2(n19), .Y(net22286) );
  AND2X1_HVT U228 ( .A1(delay_weight[75]), .A2(n19), .Y(net22287) );
  AND2X1_HVT U229 ( .A1(delay_weight[74]), .A2(n21), .Y(net22288) );
  AND2X1_HVT U230 ( .A1(delay_weight[73]), .A2(n18), .Y(net22289) );
  AND2X1_HVT U231 ( .A1(delay_weight[72]), .A2(n19), .Y(net22290) );
  AND2X1_HVT U232 ( .A1(delay_weight[71]), .A2(n20), .Y(net22291) );
  AND2X1_HVT U233 ( .A1(delay_weight[70]), .A2(n19), .Y(net22292) );
  AND2X1_HVT U234 ( .A1(delay_weight[69]), .A2(n19), .Y(net22300) );
  AND2X1_HVT U235 ( .A1(delay_weight[68]), .A2(n3), .Y(net22301) );
  AND2X1_HVT U236 ( .A1(delay_weight[67]), .A2(n21), .Y(net22302) );
  AND2X1_HVT U237 ( .A1(delay_weight[66]), .A2(n20), .Y(net22303) );
  AND2X1_HVT U238 ( .A1(delay_weight[65]), .A2(n18), .Y(net22304) );
  AND2X1_HVT U239 ( .A1(delay_weight[64]), .A2(n20), .Y(net22305) );
  AND2X1_HVT U240 ( .A1(delay_weight[63]), .A2(n20), .Y(net22306) );
  AND2X1_HVT U241 ( .A1(delay_weight[62]), .A2(n21), .Y(net22307) );
  AND2X1_HVT U242 ( .A1(delay_weight[61]), .A2(n21), .Y(net22308) );
  AND2X1_HVT U243 ( .A1(delay_weight[60]), .A2(n19), .Y(net22309) );
  AND2X1_HVT U244 ( .A1(delay_weight[59]), .A2(n3), .Y(net22317) );
  AND2X1_HVT U245 ( .A1(delay_weight[58]), .A2(n20), .Y(net22318) );
  AND2X1_HVT U246 ( .A1(delay_weight[57]), .A2(n21), .Y(net22319) );
  AND2X1_HVT U247 ( .A1(delay_weight[56]), .A2(n19), .Y(net22320) );
  AND2X1_HVT U248 ( .A1(delay_weight[55]), .A2(n19), .Y(net22321) );
  AND2X1_HVT U249 ( .A1(delay_weight[54]), .A2(n21), .Y(net22322) );
  AND2X1_HVT U250 ( .A1(delay_weight[53]), .A2(n18), .Y(net22323) );
  AND2X1_HVT U251 ( .A1(delay_weight[52]), .A2(n20), .Y(net22324) );
  AND2X1_HVT U252 ( .A1(delay_weight[51]), .A2(n19), .Y(net22325) );
  AND2X1_HVT U253 ( .A1(delay_weight[50]), .A2(n3), .Y(net22326) );
  AND2X1_HVT U254 ( .A1(delay_weight[49]), .A2(n18), .Y(net22334) );
  AND2X1_HVT U255 ( .A1(delay_weight[48]), .A2(n18), .Y(net22335) );
  AND2X1_HVT U256 ( .A1(delay_weight[47]), .A2(n20), .Y(net22336) );
  AND2X1_HVT U257 ( .A1(delay_weight[46]), .A2(n21), .Y(net22337) );
  AND2X1_HVT U258 ( .A1(delay_weight[45]), .A2(n20), .Y(net22338) );
  AND2X1_HVT U259 ( .A1(delay_weight[44]), .A2(n19), .Y(net22339) );
  AND2X1_HVT U260 ( .A1(delay_weight[43]), .A2(n18), .Y(net22340) );
  AND2X1_HVT U261 ( .A1(delay_weight[42]), .A2(n18), .Y(net22341) );
  AND2X1_HVT U262 ( .A1(delay_weight[41]), .A2(n3), .Y(net22342) );
  AND2X1_HVT U263 ( .A1(delay_weight[40]), .A2(n21), .Y(net22343) );
  AND2X1_HVT U264 ( .A1(delay_weight[39]), .A2(n19), .Y(net22351) );
  AND2X1_HVT U265 ( .A1(delay_weight[38]), .A2(n21), .Y(net22352) );
  AND2X1_HVT U266 ( .A1(delay_weight[37]), .A2(n20), .Y(net22353) );
  AND2X1_HVT U267 ( .A1(delay_weight[36]), .A2(n21), .Y(net22354) );
  AND2X1_HVT U268 ( .A1(delay_weight[35]), .A2(n20), .Y(net22355) );
  AND2X1_HVT U269 ( .A1(delay_weight[34]), .A2(n21), .Y(net22356) );
  AND2X1_HVT U270 ( .A1(delay_weight[33]), .A2(n20), .Y(net22357) );
  AND2X1_HVT U271 ( .A1(delay_weight[32]), .A2(n3), .Y(net22358) );
  AND2X1_HVT U272 ( .A1(delay_weight[31]), .A2(n20), .Y(net22359) );
  AND2X1_HVT U273 ( .A1(delay_weight[30]), .A2(n19), .Y(net22360) );
  AND2X1_HVT U274 ( .A1(delay_weight[29]), .A2(n18), .Y(net22368) );
  AND2X1_HVT U275 ( .A1(delay_weight[28]), .A2(n18), .Y(net22369) );
  AND2X1_HVT U276 ( .A1(delay_weight[27]), .A2(n18), .Y(net22370) );
  AND2X1_HVT U277 ( .A1(delay_weight[26]), .A2(n21), .Y(net22371) );
  AND2X1_HVT U278 ( .A1(delay_weight[25]), .A2(n20), .Y(net22372) );
  AND2X1_HVT U279 ( .A1(delay_weight[24]), .A2(n21), .Y(net22373) );
  AND2X1_HVT U280 ( .A1(delay_weight[23]), .A2(n3), .Y(net22374) );
  AND2X1_HVT U281 ( .A1(delay_weight[22]), .A2(n18), .Y(net22375) );
  AND2X1_HVT U282 ( .A1(delay_weight[21]), .A2(n3), .Y(net22376) );
  AND2X1_HVT U283 ( .A1(delay_weight[20]), .A2(n20), .Y(net22377) );
  AND2X1_HVT U284 ( .A1(delay_weight[19]), .A2(n21), .Y(net22385) );
  AND2X1_HVT U285 ( .A1(delay_weight[18]), .A2(n19), .Y(net22386) );
  AND2X1_HVT U286 ( .A1(delay_weight[17]), .A2(n18), .Y(net22387) );
  AND2X1_HVT U287 ( .A1(delay_weight[16]), .A2(n18), .Y(net22388) );
  AND2X1_HVT U288 ( .A1(delay_weight[15]), .A2(n18), .Y(net22389) );
  AND2X1_HVT U289 ( .A1(delay_weight[14]), .A2(n3), .Y(net22390) );
  AND2X1_HVT U290 ( .A1(delay_weight[13]), .A2(n21), .Y(net22391) );
  AND2X1_HVT U291 ( .A1(delay_weight[12]), .A2(n3), .Y(net22392) );
  AND2X1_HVT U292 ( .A1(delay_weight[11]), .A2(n21), .Y(net22393) );
  AND2X1_HVT U293 ( .A1(delay_weight[10]), .A2(n20), .Y(net22394) );
  AND2X1_HVT U294 ( .A1(delay_weight[9]), .A2(n20), .Y(net22402) );
  AND2X1_HVT U295 ( .A1(delay_weight[8]), .A2(n20), .Y(net22403) );
  AND2X1_HVT U296 ( .A1(delay_weight[7]), .A2(n21), .Y(net22404) );
  AND2X1_HVT U297 ( .A1(delay_weight[6]), .A2(n19), .Y(net22405) );
  AND2X1_HVT U298 ( .A1(delay_weight[5]), .A2(n3), .Y(net22406) );
  AND2X1_HVT U299 ( .A1(delay_weight[4]), .A2(n20), .Y(net22407) );
  AND2X1_HVT U300 ( .A1(delay_weight[3]), .A2(n3), .Y(net22408) );
  AND2X1_HVT U301 ( .A1(delay_weight[2]), .A2(n18), .Y(net22409) );
  AND2X1_HVT U302 ( .A1(delay_weight[1]), .A2(n18), .Y(net22410) );
  AND2X1_HVT U303 ( .A1(delay_weight[0]), .A2(n21), .Y(net22411) );
  NAND3X0_HVT U304 ( .A1(srstn), .A2(n43), .A3(n90), .Y(net22425) );
  AO22X1_HVT U305 ( .A1(n326), .A2(conv_weight_box[103]), .A3(n324), .A4(
        conv_weight_box[119]), .Y(n47) );
  AO22X1_HVT U306 ( .A1(n318), .A2(conv_weight_box[55]), .A3(n320), .A4(
        conv_weight_box[39]), .Y(n46) );
  AND4X1_HVT U307 ( .A1(conv1_bias_set_2_), .A2(n67), .A3(n57), .A4(n59), .Y(
        n317) );
  AND4X1_HVT U308 ( .A1(n67), .A2(n58), .A3(n57), .A4(n59), .Y(n319) );
  AO22X1_HVT U309 ( .A1(n317), .A2(conv_weight_box[183]), .A3(n319), .A4(
        conv_weight_box[199]), .Y(n45) );
  AND4X1_HVT U310 ( .A1(conv1_bias_set_2_), .A2(conv1_bias_set_3_), .A3(n67), 
        .A4(n59), .Y(n322) );
  AND4X1_HVT U311 ( .A1(conv1_bias_set_3_), .A2(n67), .A3(n58), .A4(n59), .Y(
        n321) );
  AO22X1_HVT U312 ( .A1(n322), .A2(conv_weight_box[151]), .A3(n321), .A4(
        conv_weight_box[167]), .Y(n44) );
  NAND2X0_HVT U313 ( .A1(n52), .A2(n66), .Y(n287) );
  AO22X1_HVT U314 ( .A1(n326), .A2(conv_weight_box[99]), .A3(n324), .A4(
        conv_weight_box[115]), .Y(n51) );
  AO22X1_HVT U315 ( .A1(n318), .A2(conv_weight_box[51]), .A3(n320), .A4(
        conv_weight_box[35]), .Y(n50) );
  AO22X1_HVT U316 ( .A1(n317), .A2(conv_weight_box[179]), .A3(n319), .A4(
        conv_weight_box[195]), .Y(n49) );
  AO22X1_HVT U317 ( .A1(n322), .A2(conv_weight_box[147]), .A3(n321), .A4(
        conv_weight_box[163]), .Y(n48) );
  NAND2X0_HVT U318 ( .A1(conv1_bias_set_0_), .A2(n52), .Y(n285) );
  OA22X1_HVT U319 ( .A1(n54), .A2(n287), .A3(n53), .A4(n285), .Y(n89) );
  AND2X1_HVT U320 ( .A1(conv1_bias_set_1_), .A2(n66), .Y(n336) );
  AND4X1_HVT U321 ( .A1(n336), .A2(conv1_bias_set_5_), .A3(conv1_bias_set_2_), 
        .A4(conv1_bias_set_3_), .Y(n290) );
  AND3X1_HVT U322 ( .A1(conv1_bias_set_5_), .A2(conv1_bias_set_2_), .A3(
        conv1_bias_set_3_), .Y(n55) );
  AND3X1_HVT U323 ( .A1(conv1_bias_set_1_), .A2(conv1_bias_set_0_), .A3(n55), 
        .Y(n289) );
  AO22X1_HVT U324 ( .A1(n290), .A2(conv_weight_box[15]), .A3(n289), .A4(
        conv_weight_box[11]), .Y(n63) );
  AND4X1_HVT U325 ( .A1(conv1_bias_set_2_), .A2(conv1_bias_set_3_), .A3(
        conv1_bias_set_4_), .A4(n68), .Y(n292) );
  AND4X1_HVT U326 ( .A1(conv1_bias_set_2_), .A2(conv1_bias_set_3_), .A3(
        conv1_bias_set_4_), .A4(n65), .Y(n291) );
  AO22X1_HVT U327 ( .A1(n292), .A2(conv_weight_box[83]), .A3(n291), .A4(
        conv_weight_box[87]), .Y(n62) );
  AND3X1_HVT U328 ( .A1(conv1_bias_set_2_), .A2(conv1_bias_set_3_), .A3(
        conv1_bias_set_4_), .Y(n56) );
  AND3X1_HVT U329 ( .A1(conv1_bias_set_1_), .A2(conv1_bias_set_0_), .A3(n56), 
        .Y(n294) );
  AND4X1_HVT U330 ( .A1(conv1_bias_set_5_), .A2(conv1_bias_set_2_), .A3(
        conv1_bias_set_3_), .A4(n65), .Y(n293) );
  AO22X1_HVT U331 ( .A1(n294), .A2(conv_weight_box[75]), .A3(n293), .A4(
        conv_weight_box[23]), .Y(n61) );
  AND2X1_HVT U332 ( .A1(n58), .A2(n57), .Y(n64) );
  AND3X1_HVT U333 ( .A1(n323), .A2(n68), .A3(n59), .Y(n296) );
  AND3X1_HVT U334 ( .A1(n323), .A2(n65), .A3(n59), .Y(n295) );
  AO22X1_HVT U335 ( .A1(n296), .A2(conv_weight_box[67]), .A3(n295), .A4(
        conv_weight_box[71]), .Y(n60) );
  AND4X1_HVT U336 ( .A1(conv1_bias_set_5_), .A2(conv1_bias_set_2_), .A3(
        conv1_bias_set_3_), .A4(n68), .Y(n302) );
  AND3X1_HVT U337 ( .A1(n325), .A2(n65), .A3(n67), .Y(n301) );
  AO22X1_HVT U338 ( .A1(n302), .A2(conv_weight_box[19]), .A3(n301), .A4(
        conv_weight_box[135]), .Y(n71) );
  AND3X1_HVT U339 ( .A1(conv1_bias_set_0_), .A2(conv1_bias_set_5_), .A3(
        conv1_bias_set_4_), .Y(n305) );
  AND3X1_HVT U340 ( .A1(conv1_bias_set_5_), .A2(conv1_bias_set_4_), .A3(n66), 
        .Y(n303) );
  AO22X1_HVT U341 ( .A1(n305), .A2(conv_weight_box[3]), .A3(n303), .A4(
        conv_weight_box[7]), .Y(n70) );
  AND3X1_HVT U342 ( .A1(n325), .A2(n68), .A3(n67), .Y(n307) );
  AND4X1_HVT U343 ( .A1(n336), .A2(conv1_bias_set_2_), .A3(conv1_bias_set_3_), 
        .A4(conv1_bias_set_4_), .Y(n306) );
  AO22X1_HVT U344 ( .A1(n307), .A2(conv_weight_box[131]), .A3(n306), .A4(
        conv_weight_box[79]), .Y(n69) );
  NOR3X0_HVT U345 ( .A1(n71), .A2(n70), .A3(n69), .Y(n87) );
  AO22X1_HVT U346 ( .A1(n318), .A2(conv_weight_box[47]), .A3(n317), .A4(
        conv_weight_box[175]), .Y(n77) );
  AO22X1_HVT U347 ( .A1(n320), .A2(conv_weight_box[31]), .A3(n319), .A4(
        conv_weight_box[191]), .Y(n76) );
  AO22X1_HVT U348 ( .A1(n322), .A2(conv_weight_box[143]), .A3(n321), .A4(
        conv_weight_box[159]), .Y(n74) );
  AO22X1_HVT U349 ( .A1(n324), .A2(conv_weight_box[111]), .A3(n323), .A4(
        conv_weight_box[63]), .Y(n73) );
  AO22X1_HVT U350 ( .A1(n326), .A2(conv_weight_box[95]), .A3(n325), .A4(
        conv_weight_box[127]), .Y(n72) );
  OR3X1_HVT U351 ( .A1(n74), .A2(n73), .A3(n72), .Y(n75) );
  OR3X1_HVT U352 ( .A1(n77), .A2(n76), .A3(n75), .Y(n85) );
  AND2X1_HVT U353 ( .A1(conv1_bias_set_1_), .A2(conv1_bias_set_0_), .Y(n334)
         );
  AO22X1_HVT U354 ( .A1(n318), .A2(conv_weight_box[43]), .A3(n317), .A4(
        conv_weight_box[171]), .Y(n83) );
  AO22X1_HVT U355 ( .A1(n320), .A2(conv_weight_box[27]), .A3(n319), .A4(
        conv_weight_box[187]), .Y(n82) );
  AO22X1_HVT U356 ( .A1(n322), .A2(conv_weight_box[139]), .A3(n321), .A4(
        conv_weight_box[155]), .Y(n80) );
  AO22X1_HVT U357 ( .A1(n324), .A2(conv_weight_box[107]), .A3(n323), .A4(
        conv_weight_box[59]), .Y(n79) );
  AO22X1_HVT U358 ( .A1(n326), .A2(conv_weight_box[91]), .A3(n325), .A4(
        conv_weight_box[123]), .Y(n78) );
  OR3X1_HVT U359 ( .A1(n80), .A2(n79), .A3(n78), .Y(n81) );
  OR3X1_HVT U360 ( .A1(n83), .A2(n82), .A3(n81), .Y(n84) );
  AOI22X1_HVT U361 ( .A1(n336), .A2(n85), .A3(n334), .A4(n84), .Y(n86) );
  AO22X1_HVT U362 ( .A1(conv_weight_box[119]), .A2(n387), .A3(
        conv_weight_box[103]), .A4(n389), .Y(n94) );
  AO22X1_HVT U363 ( .A1(conv_weight_box[55]), .A2(n381), .A3(
        conv_weight_box[39]), .A4(n383), .Y(n93) );
  AND4X1_HVT U364 ( .A1(n114), .A2(n105), .A3(n104), .A4(n106), .Y(n382) );
  AND4X1_HVT U365 ( .A1(set_2_), .A2(n114), .A3(n104), .A4(n106), .Y(n380) );
  AO22X1_HVT U366 ( .A1(conv_weight_box[199]), .A2(n382), .A3(
        conv_weight_box[183]), .A4(n380), .Y(n92) );
  AND4X1_HVT U367 ( .A1(set_2_), .A2(set_3_), .A3(n114), .A4(n106), .Y(n385)
         );
  AND4X1_HVT U368 ( .A1(set_3_), .A2(n114), .A3(n105), .A4(n106), .Y(n384) );
  AO22X1_HVT U369 ( .A1(conv_weight_box[151]), .A2(n385), .A3(
        conv_weight_box[167]), .A4(n384), .Y(n91) );
  NAND2X0_HVT U370 ( .A1(n99), .A2(n113), .Y(n351) );
  AO22X1_HVT U371 ( .A1(conv_weight_box[115]), .A2(n387), .A3(
        conv_weight_box[99]), .A4(n389), .Y(n98) );
  AO22X1_HVT U372 ( .A1(conv_weight_box[51]), .A2(n381), .A3(
        conv_weight_box[35]), .A4(n383), .Y(n97) );
  AO22X1_HVT U373 ( .A1(conv_weight_box[195]), .A2(n382), .A3(
        conv_weight_box[179]), .A4(n380), .Y(n96) );
  AO22X1_HVT U374 ( .A1(conv_weight_box[147]), .A2(n385), .A3(
        conv_weight_box[163]), .A4(n384), .Y(n95) );
  NAND2X0_HVT U375 ( .A1(set_0_), .A2(n99), .Y(n349) );
  OA22X1_HVT U376 ( .A1(n101), .A2(n351), .A3(n100), .A4(n349), .Y(n136) );
  AND2X1_HVT U377 ( .A1(set_1_), .A2(n113), .Y(n399) );
  AND4X1_HVT U378 ( .A1(n399), .A2(set_5_), .A3(set_2_), .A4(set_3_), .Y(n354)
         );
  AND3X1_HVT U379 ( .A1(set_5_), .A2(set_2_), .A3(set_3_), .Y(n102) );
  AND3X1_HVT U380 ( .A1(set_1_), .A2(set_0_), .A3(n102), .Y(n353) );
  AO22X1_HVT U381 ( .A1(conv_weight_box[15]), .A2(n354), .A3(
        conv_weight_box[11]), .A4(n353), .Y(n110) );
  AND4X1_HVT U382 ( .A1(set_2_), .A2(set_3_), .A3(set_4_), .A4(n115), .Y(n356)
         );
  AND4X1_HVT U383 ( .A1(set_2_), .A2(set_3_), .A3(set_4_), .A4(n112), .Y(n355)
         );
  AO22X1_HVT U384 ( .A1(conv_weight_box[83]), .A2(n356), .A3(
        conv_weight_box[87]), .A4(n355), .Y(n109) );
  AND3X1_HVT U385 ( .A1(set_2_), .A2(set_3_), .A3(set_4_), .Y(n103) );
  AND3X1_HVT U386 ( .A1(set_1_), .A2(set_0_), .A3(n103), .Y(n358) );
  AND4X1_HVT U387 ( .A1(set_5_), .A2(set_2_), .A3(set_3_), .A4(n112), .Y(n357)
         );
  AO22X1_HVT U388 ( .A1(conv_weight_box[75]), .A2(n358), .A3(
        conv_weight_box[23]), .A4(n357), .Y(n108) );
  AND2X1_HVT U389 ( .A1(n105), .A2(n104), .Y(n111) );
  AND3X1_HVT U390 ( .A1(n386), .A2(n115), .A3(n106), .Y(n360) );
  AND3X1_HVT U391 ( .A1(n386), .A2(n112), .A3(n106), .Y(n359) );
  AO22X1_HVT U392 ( .A1(conv_weight_box[67]), .A2(n360), .A3(
        conv_weight_box[71]), .A4(n359), .Y(n107) );
  AND4X1_HVT U393 ( .A1(set_5_), .A2(set_2_), .A3(set_3_), .A4(n115), .Y(n366)
         );
  AND3X1_HVT U394 ( .A1(n388), .A2(n112), .A3(n114), .Y(n365) );
  AO22X1_HVT U395 ( .A1(conv_weight_box[19]), .A2(n366), .A3(
        conv_weight_box[135]), .A4(n365), .Y(n118) );
  AND3X1_HVT U396 ( .A1(set_0_), .A2(set_5_), .A3(set_4_), .Y(n368) );
  AND3X1_HVT U397 ( .A1(set_5_), .A2(set_4_), .A3(n113), .Y(n367) );
  AO22X1_HVT U398 ( .A1(conv_weight_box[3]), .A2(n368), .A3(conv_weight_box[7]), .A4(n367), .Y(n117) );
  AND3X1_HVT U399 ( .A1(n388), .A2(n115), .A3(n114), .Y(n370) );
  AND4X1_HVT U400 ( .A1(n399), .A2(set_2_), .A3(set_3_), .A4(set_4_), .Y(n369)
         );
  AO22X1_HVT U401 ( .A1(conv_weight_box[131]), .A2(n370), .A3(
        conv_weight_box[79]), .A4(n369), .Y(n116) );
  NOR3X0_HVT U402 ( .A1(n118), .A2(n117), .A3(n116), .Y(n134) );
  AO22X1_HVT U403 ( .A1(conv_weight_box[47]), .A2(n381), .A3(
        conv_weight_box[175]), .A4(n380), .Y(n124) );
  AO22X1_HVT U404 ( .A1(conv_weight_box[31]), .A2(n383), .A3(
        conv_weight_box[191]), .A4(n382), .Y(n123) );
  AO22X1_HVT U405 ( .A1(conv_weight_box[143]), .A2(n385), .A3(
        conv_weight_box[159]), .A4(n384), .Y(n121) );
  AO22X1_HVT U406 ( .A1(conv_weight_box[111]), .A2(n387), .A3(
        conv_weight_box[63]), .A4(n386), .Y(n120) );
  AO22X1_HVT U407 ( .A1(conv_weight_box[95]), .A2(n389), .A3(
        conv_weight_box[127]), .A4(n388), .Y(n119) );
  OR3X1_HVT U408 ( .A1(n121), .A2(n120), .A3(n119), .Y(n122) );
  OR3X1_HVT U409 ( .A1(n124), .A2(n123), .A3(n122), .Y(n132) );
  AND2X1_HVT U410 ( .A1(set_1_), .A2(set_0_), .Y(n397) );
  AO22X1_HVT U411 ( .A1(conv_weight_box[43]), .A2(n381), .A3(
        conv_weight_box[171]), .A4(n380), .Y(n130) );
  AO22X1_HVT U412 ( .A1(conv_weight_box[27]), .A2(n383), .A3(
        conv_weight_box[187]), .A4(n382), .Y(n129) );
  AO22X1_HVT U413 ( .A1(conv_weight_box[139]), .A2(n385), .A3(
        conv_weight_box[155]), .A4(n384), .Y(n127) );
  AO22X1_HVT U414 ( .A1(conv_weight_box[107]), .A2(n387), .A3(
        conv_weight_box[59]), .A4(n386), .Y(n126) );
  AO22X1_HVT U415 ( .A1(conv_weight_box[91]), .A2(n389), .A3(
        conv_weight_box[123]), .A4(n388), .Y(n125) );
  OR3X1_HVT U416 ( .A1(n127), .A2(n126), .A3(n125), .Y(n128) );
  OR3X1_HVT U417 ( .A1(n130), .A2(n129), .A3(n128), .Y(n131) );
  AOI22X1_HVT U418 ( .A1(n399), .A2(n132), .A3(n397), .A4(n131), .Y(n133) );
  AO22X1_HVT U419 ( .A1(n326), .A2(conv_weight_box[102]), .A3(n324), .A4(
        conv_weight_box[118]), .Y(n140) );
  AO22X1_HVT U420 ( .A1(n318), .A2(conv_weight_box[54]), .A3(n320), .A4(
        conv_weight_box[38]), .Y(n139) );
  AO22X1_HVT U421 ( .A1(n317), .A2(conv_weight_box[182]), .A3(n319), .A4(
        conv_weight_box[198]), .Y(n138) );
  AO22X1_HVT U422 ( .A1(n322), .A2(conv_weight_box[150]), .A3(n321), .A4(
        conv_weight_box[166]), .Y(n137) );
  AO22X1_HVT U423 ( .A1(n326), .A2(conv_weight_box[98]), .A3(n324), .A4(
        conv_weight_box[114]), .Y(n144) );
  AO22X1_HVT U424 ( .A1(n318), .A2(conv_weight_box[50]), .A3(n320), .A4(
        conv_weight_box[34]), .Y(n143) );
  AO22X1_HVT U425 ( .A1(n317), .A2(conv_weight_box[178]), .A3(n319), .A4(
        conv_weight_box[194]), .Y(n142) );
  AO22X1_HVT U426 ( .A1(n322), .A2(conv_weight_box[146]), .A3(n321), .A4(
        conv_weight_box[162]), .Y(n141) );
  OA22X1_HVT U427 ( .A1(n146), .A2(n287), .A3(n145), .A4(n285), .Y(n171) );
  AO22X1_HVT U428 ( .A1(n290), .A2(conv_weight_box[14]), .A3(n289), .A4(
        conv_weight_box[10]), .Y(n150) );
  AO22X1_HVT U429 ( .A1(n292), .A2(conv_weight_box[82]), .A3(n291), .A4(
        conv_weight_box[86]), .Y(n149) );
  AO22X1_HVT U430 ( .A1(n294), .A2(conv_weight_box[74]), .A3(n293), .A4(
        conv_weight_box[22]), .Y(n148) );
  AO22X1_HVT U431 ( .A1(n296), .A2(conv_weight_box[66]), .A3(n295), .A4(
        conv_weight_box[70]), .Y(n147) );
  AO22X1_HVT U432 ( .A1(n302), .A2(conv_weight_box[18]), .A3(n301), .A4(
        conv_weight_box[134]), .Y(n153) );
  AO22X1_HVT U433 ( .A1(n305), .A2(conv_weight_box[2]), .A3(n303), .A4(
        conv_weight_box[6]), .Y(n152) );
  AO22X1_HVT U434 ( .A1(n307), .A2(conv_weight_box[130]), .A3(n306), .A4(
        conv_weight_box[78]), .Y(n151) );
  NOR3X0_HVT U435 ( .A1(n153), .A2(n152), .A3(n151), .Y(n169) );
  AO22X1_HVT U436 ( .A1(n318), .A2(conv_weight_box[46]), .A3(n317), .A4(
        conv_weight_box[174]), .Y(n159) );
  AO22X1_HVT U437 ( .A1(n320), .A2(conv_weight_box[30]), .A3(n319), .A4(
        conv_weight_box[190]), .Y(n158) );
  AO22X1_HVT U438 ( .A1(n322), .A2(conv_weight_box[142]), .A3(n321), .A4(
        conv_weight_box[158]), .Y(n156) );
  AO22X1_HVT U439 ( .A1(n324), .A2(conv_weight_box[110]), .A3(n323), .A4(
        conv_weight_box[62]), .Y(n155) );
  AO22X1_HVT U440 ( .A1(n326), .A2(conv_weight_box[94]), .A3(n325), .A4(
        conv_weight_box[126]), .Y(n154) );
  OR3X1_HVT U441 ( .A1(n156), .A2(n155), .A3(n154), .Y(n157) );
  OR3X1_HVT U442 ( .A1(n159), .A2(n158), .A3(n157), .Y(n167) );
  AO22X1_HVT U443 ( .A1(n318), .A2(conv_weight_box[42]), .A3(n317), .A4(
        conv_weight_box[170]), .Y(n165) );
  AO22X1_HVT U444 ( .A1(n320), .A2(conv_weight_box[26]), .A3(n319), .A4(
        conv_weight_box[186]), .Y(n164) );
  AO22X1_HVT U445 ( .A1(n322), .A2(conv_weight_box[138]), .A3(n321), .A4(
        conv_weight_box[154]), .Y(n162) );
  AO22X1_HVT U446 ( .A1(n324), .A2(conv_weight_box[106]), .A3(n323), .A4(
        conv_weight_box[58]), .Y(n161) );
  AO22X1_HVT U447 ( .A1(n326), .A2(conv_weight_box[90]), .A3(n325), .A4(
        conv_weight_box[122]), .Y(n160) );
  OR3X1_HVT U448 ( .A1(n162), .A2(n161), .A3(n160), .Y(n163) );
  OR3X1_HVT U449 ( .A1(n165), .A2(n164), .A3(n163), .Y(n166) );
  AOI22X1_HVT U450 ( .A1(n336), .A2(n167), .A3(n334), .A4(n166), .Y(n168) );
  AO22X1_HVT U451 ( .A1(n389), .A2(conv_weight_box[102]), .A3(n387), .A4(
        conv_weight_box[118]), .Y(n175) );
  AO22X1_HVT U452 ( .A1(n381), .A2(conv_weight_box[54]), .A3(n383), .A4(
        conv_weight_box[38]), .Y(n174) );
  AO22X1_HVT U453 ( .A1(n380), .A2(conv_weight_box[182]), .A3(n382), .A4(
        conv_weight_box[198]), .Y(n173) );
  AO22X1_HVT U454 ( .A1(n385), .A2(conv_weight_box[150]), .A3(n384), .A4(
        conv_weight_box[166]), .Y(n172) );
  AO22X1_HVT U455 ( .A1(n389), .A2(conv_weight_box[98]), .A3(n387), .A4(
        conv_weight_box[114]), .Y(n179) );
  AO22X1_HVT U456 ( .A1(n381), .A2(conv_weight_box[50]), .A3(n383), .A4(
        conv_weight_box[34]), .Y(n178) );
  AO22X1_HVT U457 ( .A1(n380), .A2(conv_weight_box[178]), .A3(n382), .A4(
        conv_weight_box[194]), .Y(n177) );
  AO22X1_HVT U458 ( .A1(n385), .A2(conv_weight_box[146]), .A3(n384), .A4(
        conv_weight_box[162]), .Y(n176) );
  OA22X1_HVT U459 ( .A1(n181), .A2(n351), .A3(n180), .A4(n349), .Y(n206) );
  AO22X1_HVT U460 ( .A1(n354), .A2(conv_weight_box[14]), .A3(n353), .A4(
        conv_weight_box[10]), .Y(n185) );
  AO22X1_HVT U461 ( .A1(n356), .A2(conv_weight_box[82]), .A3(n355), .A4(
        conv_weight_box[86]), .Y(n184) );
  AO22X1_HVT U462 ( .A1(n358), .A2(conv_weight_box[74]), .A3(n357), .A4(
        conv_weight_box[22]), .Y(n183) );
  AO22X1_HVT U463 ( .A1(n360), .A2(conv_weight_box[66]), .A3(n359), .A4(
        conv_weight_box[70]), .Y(n182) );
  AO22X1_HVT U464 ( .A1(n366), .A2(conv_weight_box[18]), .A3(n365), .A4(
        conv_weight_box[134]), .Y(n188) );
  AO22X1_HVT U465 ( .A1(n368), .A2(conv_weight_box[2]), .A3(n367), .A4(
        conv_weight_box[6]), .Y(n187) );
  AO22X1_HVT U466 ( .A1(n370), .A2(conv_weight_box[130]), .A3(n369), .A4(
        conv_weight_box[78]), .Y(n186) );
  NOR3X0_HVT U467 ( .A1(n188), .A2(n187), .A3(n186), .Y(n204) );
  AO22X1_HVT U468 ( .A1(n381), .A2(conv_weight_box[46]), .A3(n380), .A4(
        conv_weight_box[174]), .Y(n194) );
  AO22X1_HVT U469 ( .A1(n383), .A2(conv_weight_box[30]), .A3(n382), .A4(
        conv_weight_box[190]), .Y(n193) );
  AO22X1_HVT U470 ( .A1(n385), .A2(conv_weight_box[142]), .A3(n384), .A4(
        conv_weight_box[158]), .Y(n191) );
  AO22X1_HVT U471 ( .A1(n387), .A2(conv_weight_box[110]), .A3(n386), .A4(
        conv_weight_box[62]), .Y(n190) );
  AO22X1_HVT U472 ( .A1(n389), .A2(conv_weight_box[94]), .A3(n388), .A4(
        conv_weight_box[126]), .Y(n189) );
  OR3X1_HVT U473 ( .A1(n191), .A2(n190), .A3(n189), .Y(n192) );
  OR3X1_HVT U474 ( .A1(n194), .A2(n193), .A3(n192), .Y(n202) );
  AO22X1_HVT U475 ( .A1(n381), .A2(conv_weight_box[42]), .A3(n380), .A4(
        conv_weight_box[170]), .Y(n200) );
  AO22X1_HVT U476 ( .A1(n383), .A2(conv_weight_box[26]), .A3(n382), .A4(
        conv_weight_box[186]), .Y(n199) );
  AO22X1_HVT U477 ( .A1(n385), .A2(conv_weight_box[138]), .A3(n384), .A4(
        conv_weight_box[154]), .Y(n197) );
  AO22X1_HVT U478 ( .A1(n387), .A2(conv_weight_box[106]), .A3(n386), .A4(
        conv_weight_box[58]), .Y(n196) );
  AO22X1_HVT U479 ( .A1(n389), .A2(conv_weight_box[90]), .A3(n388), .A4(
        conv_weight_box[122]), .Y(n195) );
  OR3X1_HVT U480 ( .A1(n197), .A2(n196), .A3(n195), .Y(n198) );
  OR3X1_HVT U481 ( .A1(n200), .A2(n199), .A3(n198), .Y(n201) );
  AOI22X1_HVT U482 ( .A1(n399), .A2(n202), .A3(n397), .A4(n201), .Y(n203) );
  AO22X1_HVT U483 ( .A1(n326), .A2(conv_weight_box[101]), .A3(n324), .A4(
        conv_weight_box[117]), .Y(n210) );
  AO22X1_HVT U484 ( .A1(n318), .A2(conv_weight_box[53]), .A3(n320), .A4(
        conv_weight_box[37]), .Y(n209) );
  AO22X1_HVT U485 ( .A1(n317), .A2(conv_weight_box[181]), .A3(n319), .A4(
        conv_weight_box[197]), .Y(n208) );
  AO22X1_HVT U486 ( .A1(n322), .A2(conv_weight_box[149]), .A3(n321), .A4(
        conv_weight_box[165]), .Y(n207) );
  AO22X1_HVT U487 ( .A1(n326), .A2(conv_weight_box[97]), .A3(n324), .A4(
        conv_weight_box[113]), .Y(n214) );
  AO22X1_HVT U488 ( .A1(n318), .A2(conv_weight_box[49]), .A3(n320), .A4(
        conv_weight_box[33]), .Y(n213) );
  AO22X1_HVT U489 ( .A1(n317), .A2(conv_weight_box[177]), .A3(n319), .A4(
        conv_weight_box[193]), .Y(n212) );
  AO22X1_HVT U490 ( .A1(n322), .A2(conv_weight_box[145]), .A3(n321), .A4(
        conv_weight_box[161]), .Y(n211) );
  OA22X1_HVT U491 ( .A1(n216), .A2(n287), .A3(n215), .A4(n285), .Y(n241) );
  AO22X1_HVT U492 ( .A1(n290), .A2(conv_weight_box[13]), .A3(n289), .A4(
        conv_weight_box[9]), .Y(n220) );
  AO22X1_HVT U493 ( .A1(n292), .A2(conv_weight_box[81]), .A3(n291), .A4(
        conv_weight_box[85]), .Y(n219) );
  AO22X1_HVT U494 ( .A1(n294), .A2(conv_weight_box[73]), .A3(n293), .A4(
        conv_weight_box[21]), .Y(n218) );
  AO22X1_HVT U495 ( .A1(n296), .A2(conv_weight_box[65]), .A3(n295), .A4(
        conv_weight_box[69]), .Y(n217) );
  AO22X1_HVT U496 ( .A1(n302), .A2(conv_weight_box[17]), .A3(n301), .A4(
        conv_weight_box[133]), .Y(n223) );
  AO22X1_HVT U497 ( .A1(n305), .A2(conv_weight_box[1]), .A3(n303), .A4(
        conv_weight_box[5]), .Y(n222) );
  AO22X1_HVT U498 ( .A1(n307), .A2(conv_weight_box[129]), .A3(n306), .A4(
        conv_weight_box[77]), .Y(n221) );
  NOR3X0_HVT U499 ( .A1(n223), .A2(n222), .A3(n221), .Y(n239) );
  AO22X1_HVT U500 ( .A1(n318), .A2(conv_weight_box[45]), .A3(n317), .A4(
        conv_weight_box[173]), .Y(n229) );
  AO22X1_HVT U501 ( .A1(n320), .A2(conv_weight_box[29]), .A3(n319), .A4(
        conv_weight_box[189]), .Y(n228) );
  AO22X1_HVT U502 ( .A1(n322), .A2(conv_weight_box[141]), .A3(n321), .A4(
        conv_weight_box[157]), .Y(n226) );
  AO22X1_HVT U503 ( .A1(n324), .A2(conv_weight_box[109]), .A3(n323), .A4(
        conv_weight_box[61]), .Y(n225) );
  AO22X1_HVT U504 ( .A1(n326), .A2(conv_weight_box[93]), .A3(n325), .A4(
        conv_weight_box[125]), .Y(n224) );
  OR3X1_HVT U505 ( .A1(n226), .A2(n225), .A3(n224), .Y(n227) );
  OR3X1_HVT U506 ( .A1(n229), .A2(n228), .A3(n227), .Y(n237) );
  AO22X1_HVT U507 ( .A1(n318), .A2(conv_weight_box[41]), .A3(n317), .A4(
        conv_weight_box[169]), .Y(n235) );
  AO22X1_HVT U508 ( .A1(n320), .A2(conv_weight_box[25]), .A3(n319), .A4(
        conv_weight_box[185]), .Y(n234) );
  AO22X1_HVT U509 ( .A1(n322), .A2(conv_weight_box[137]), .A3(n321), .A4(
        conv_weight_box[153]), .Y(n232) );
  AO22X1_HVT U510 ( .A1(n324), .A2(conv_weight_box[105]), .A3(n323), .A4(
        conv_weight_box[57]), .Y(n231) );
  AO22X1_HVT U511 ( .A1(n326), .A2(conv_weight_box[89]), .A3(n325), .A4(
        conv_weight_box[121]), .Y(n230) );
  OR3X1_HVT U512 ( .A1(n232), .A2(n231), .A3(n230), .Y(n233) );
  OR3X1_HVT U513 ( .A1(n235), .A2(n234), .A3(n233), .Y(n236) );
  AOI22X1_HVT U514 ( .A1(n336), .A2(n237), .A3(n334), .A4(n236), .Y(n238) );
  AO22X1_HVT U515 ( .A1(n389), .A2(conv_weight_box[101]), .A3(n387), .A4(
        conv_weight_box[117]), .Y(n245) );
  AO22X1_HVT U516 ( .A1(n381), .A2(conv_weight_box[53]), .A3(n383), .A4(
        conv_weight_box[37]), .Y(n244) );
  AO22X1_HVT U517 ( .A1(n380), .A2(conv_weight_box[181]), .A3(n382), .A4(
        conv_weight_box[197]), .Y(n243) );
  AO22X1_HVT U518 ( .A1(n385), .A2(conv_weight_box[149]), .A3(n384), .A4(
        conv_weight_box[165]), .Y(n242) );
  AO22X1_HVT U519 ( .A1(n389), .A2(conv_weight_box[97]), .A3(n387), .A4(
        conv_weight_box[113]), .Y(n249) );
  AO22X1_HVT U520 ( .A1(n381), .A2(conv_weight_box[49]), .A3(n383), .A4(
        conv_weight_box[33]), .Y(n248) );
  AO22X1_HVT U521 ( .A1(n380), .A2(conv_weight_box[177]), .A3(n382), .A4(
        conv_weight_box[193]), .Y(n247) );
  AO22X1_HVT U522 ( .A1(n385), .A2(conv_weight_box[145]), .A3(n384), .A4(
        conv_weight_box[161]), .Y(n246) );
  OA22X1_HVT U523 ( .A1(n251), .A2(n351), .A3(n250), .A4(n349), .Y(n276) );
  AO22X1_HVT U524 ( .A1(n354), .A2(conv_weight_box[13]), .A3(n353), .A4(
        conv_weight_box[9]), .Y(n255) );
  AO22X1_HVT U525 ( .A1(n356), .A2(conv_weight_box[81]), .A3(n355), .A4(
        conv_weight_box[85]), .Y(n254) );
  AO22X1_HVT U526 ( .A1(n358), .A2(conv_weight_box[73]), .A3(n357), .A4(
        conv_weight_box[21]), .Y(n253) );
  AO22X1_HVT U527 ( .A1(n360), .A2(conv_weight_box[65]), .A3(n359), .A4(
        conv_weight_box[69]), .Y(n252) );
  AO22X1_HVT U528 ( .A1(n366), .A2(conv_weight_box[17]), .A3(n365), .A4(
        conv_weight_box[133]), .Y(n258) );
  AO22X1_HVT U529 ( .A1(n368), .A2(conv_weight_box[1]), .A3(n367), .A4(
        conv_weight_box[5]), .Y(n257) );
  AO22X1_HVT U530 ( .A1(n370), .A2(conv_weight_box[129]), .A3(n369), .A4(
        conv_weight_box[77]), .Y(n256) );
  NOR3X0_HVT U531 ( .A1(n258), .A2(n257), .A3(n256), .Y(n274) );
  AO22X1_HVT U532 ( .A1(n381), .A2(conv_weight_box[45]), .A3(n380), .A4(
        conv_weight_box[173]), .Y(n264) );
  AO22X1_HVT U533 ( .A1(n383), .A2(conv_weight_box[29]), .A3(n382), .A4(
        conv_weight_box[189]), .Y(n263) );
  AO22X1_HVT U534 ( .A1(n385), .A2(conv_weight_box[141]), .A3(n384), .A4(
        conv_weight_box[157]), .Y(n261) );
  AO22X1_HVT U535 ( .A1(n387), .A2(conv_weight_box[109]), .A3(n386), .A4(
        conv_weight_box[61]), .Y(n260) );
  AO22X1_HVT U536 ( .A1(n389), .A2(conv_weight_box[93]), .A3(n388), .A4(
        conv_weight_box[125]), .Y(n259) );
  OR3X1_HVT U537 ( .A1(n261), .A2(n260), .A3(n259), .Y(n262) );
  OR3X1_HVT U538 ( .A1(n264), .A2(n263), .A3(n262), .Y(n272) );
  AO22X1_HVT U539 ( .A1(n381), .A2(conv_weight_box[41]), .A3(n380), .A4(
        conv_weight_box[169]), .Y(n270) );
  AO22X1_HVT U540 ( .A1(n383), .A2(conv_weight_box[25]), .A3(n382), .A4(
        conv_weight_box[185]), .Y(n269) );
  AO22X1_HVT U541 ( .A1(n385), .A2(conv_weight_box[137]), .A3(n384), .A4(
        conv_weight_box[153]), .Y(n267) );
  AO22X1_HVT U542 ( .A1(n387), .A2(conv_weight_box[105]), .A3(n386), .A4(
        conv_weight_box[57]), .Y(n266) );
  AO22X1_HVT U543 ( .A1(n389), .A2(conv_weight_box[89]), .A3(n388), .A4(
        conv_weight_box[121]), .Y(n265) );
  OR3X1_HVT U544 ( .A1(n267), .A2(n266), .A3(n265), .Y(n268) );
  OR3X1_HVT U545 ( .A1(n270), .A2(n269), .A3(n268), .Y(n271) );
  AOI22X1_HVT U546 ( .A1(n399), .A2(n272), .A3(n397), .A4(n271), .Y(n273) );
  AO22X1_HVT U547 ( .A1(n326), .A2(conv_weight_box[100]), .A3(n324), .A4(
        conv_weight_box[116]), .Y(n280) );
  AO22X1_HVT U548 ( .A1(n318), .A2(conv_weight_box[52]), .A3(n320), .A4(
        conv_weight_box[36]), .Y(n279) );
  AO22X1_HVT U549 ( .A1(n317), .A2(conv_weight_box[180]), .A3(n319), .A4(
        conv_weight_box[196]), .Y(n278) );
  AO22X1_HVT U550 ( .A1(n322), .A2(conv_weight_box[148]), .A3(n321), .A4(
        conv_weight_box[164]), .Y(n277) );
  AO22X1_HVT U551 ( .A1(n326), .A2(conv_weight_box[96]), .A3(n324), .A4(
        conv_weight_box[112]), .Y(n284) );
  AO22X1_HVT U552 ( .A1(n318), .A2(conv_weight_box[48]), .A3(n320), .A4(
        conv_weight_box[32]), .Y(n283) );
  AO22X1_HVT U553 ( .A1(n317), .A2(conv_weight_box[176]), .A3(n319), .A4(
        conv_weight_box[192]), .Y(n282) );
  AO22X1_HVT U554 ( .A1(n322), .A2(conv_weight_box[144]), .A3(n321), .A4(
        conv_weight_box[160]), .Y(n281) );
  OA22X1_HVT U555 ( .A1(n288), .A2(n287), .A3(n286), .A4(n285), .Y(n340) );
  AO22X1_HVT U556 ( .A1(n290), .A2(conv_weight_box[12]), .A3(n289), .A4(
        conv_weight_box[8]), .Y(n300) );
  AO22X1_HVT U557 ( .A1(n292), .A2(conv_weight_box[80]), .A3(n291), .A4(
        conv_weight_box[84]), .Y(n299) );
  AO22X1_HVT U558 ( .A1(n294), .A2(conv_weight_box[72]), .A3(n293), .A4(
        conv_weight_box[20]), .Y(n298) );
  AO22X1_HVT U559 ( .A1(n296), .A2(conv_weight_box[64]), .A3(n295), .A4(
        conv_weight_box[68]), .Y(n297) );
  AO22X1_HVT U560 ( .A1(n302), .A2(conv_weight_box[16]), .A3(n301), .A4(
        conv_weight_box[132]), .Y(n310) );
  AO22X1_HVT U561 ( .A1(n305), .A2(conv_weight_box[0]), .A3(n303), .A4(
        conv_weight_box[4]), .Y(n309) );
  AO22X1_HVT U562 ( .A1(n307), .A2(conv_weight_box[128]), .A3(n306), .A4(
        conv_weight_box[76]), .Y(n308) );
  NOR3X0_HVT U563 ( .A1(n310), .A2(n309), .A3(n308), .Y(n338) );
  AO22X1_HVT U564 ( .A1(n318), .A2(conv_weight_box[44]), .A3(n317), .A4(
        conv_weight_box[172]), .Y(n316) );
  AO22X1_HVT U565 ( .A1(n320), .A2(conv_weight_box[28]), .A3(n319), .A4(
        conv_weight_box[188]), .Y(n315) );
  AO22X1_HVT U566 ( .A1(n322), .A2(conv_weight_box[140]), .A3(n321), .A4(
        conv_weight_box[156]), .Y(n313) );
  AO22X1_HVT U567 ( .A1(n324), .A2(conv_weight_box[108]), .A3(n323), .A4(
        conv_weight_box[60]), .Y(n312) );
  AO22X1_HVT U568 ( .A1(n326), .A2(conv_weight_box[92]), .A3(n325), .A4(
        conv_weight_box[124]), .Y(n311) );
  OR3X1_HVT U569 ( .A1(n313), .A2(n312), .A3(n311), .Y(n314) );
  OR3X1_HVT U570 ( .A1(n316), .A2(n315), .A3(n314), .Y(n335) );
  AO22X1_HVT U571 ( .A1(n318), .A2(conv_weight_box[40]), .A3(n317), .A4(
        conv_weight_box[168]), .Y(n332) );
  AO22X1_HVT U572 ( .A1(n320), .A2(conv_weight_box[24]), .A3(n319), .A4(
        conv_weight_box[184]), .Y(n331) );
  AO22X1_HVT U573 ( .A1(n322), .A2(conv_weight_box[136]), .A3(n321), .A4(
        conv_weight_box[152]), .Y(n329) );
  AO22X1_HVT U574 ( .A1(n324), .A2(conv_weight_box[104]), .A3(n323), .A4(
        conv_weight_box[56]), .Y(n328) );
  AO22X1_HVT U575 ( .A1(n326), .A2(conv_weight_box[88]), .A3(n325), .A4(
        conv_weight_box[120]), .Y(n327) );
  OR3X1_HVT U576 ( .A1(n329), .A2(n328), .A3(n327), .Y(n330) );
  OR3X1_HVT U577 ( .A1(n332), .A2(n331), .A3(n330), .Y(n333) );
  AOI22X1_HVT U578 ( .A1(n336), .A2(n335), .A3(n334), .A4(n333), .Y(n337) );
  AO22X1_HVT U579 ( .A1(n389), .A2(conv_weight_box[100]), .A3(n387), .A4(
        conv_weight_box[116]), .Y(n344) );
  AO22X1_HVT U580 ( .A1(n381), .A2(conv_weight_box[52]), .A3(n383), .A4(
        conv_weight_box[36]), .Y(n343) );
  AO22X1_HVT U581 ( .A1(n380), .A2(conv_weight_box[180]), .A3(n382), .A4(
        conv_weight_box[196]), .Y(n342) );
  AO22X1_HVT U582 ( .A1(n385), .A2(conv_weight_box[148]), .A3(n384), .A4(
        conv_weight_box[164]), .Y(n341) );
  AO22X1_HVT U583 ( .A1(n389), .A2(conv_weight_box[96]), .A3(n387), .A4(
        conv_weight_box[112]), .Y(n348) );
  AO22X1_HVT U584 ( .A1(n381), .A2(conv_weight_box[48]), .A3(n383), .A4(
        conv_weight_box[32]), .Y(n347) );
  AO22X1_HVT U585 ( .A1(n380), .A2(conv_weight_box[176]), .A3(n382), .A4(
        conv_weight_box[192]), .Y(n346) );
  AO22X1_HVT U586 ( .A1(n385), .A2(conv_weight_box[144]), .A3(n384), .A4(
        conv_weight_box[160]), .Y(n345) );
  OA22X1_HVT U587 ( .A1(n352), .A2(n351), .A3(n350), .A4(n349), .Y(n403) );
  AO22X1_HVT U588 ( .A1(n354), .A2(conv_weight_box[12]), .A3(n353), .A4(
        conv_weight_box[8]), .Y(n364) );
  AO22X1_HVT U589 ( .A1(n356), .A2(conv_weight_box[80]), .A3(n355), .A4(
        conv_weight_box[84]), .Y(n363) );
  AO22X1_HVT U590 ( .A1(n358), .A2(conv_weight_box[72]), .A3(n357), .A4(
        conv_weight_box[20]), .Y(n362) );
  AO22X1_HVT U591 ( .A1(n360), .A2(conv_weight_box[64]), .A3(n359), .A4(
        conv_weight_box[68]), .Y(n361) );
  AO22X1_HVT U592 ( .A1(n366), .A2(conv_weight_box[16]), .A3(n365), .A4(
        conv_weight_box[132]), .Y(n373) );
  AO22X1_HVT U593 ( .A1(n368), .A2(conv_weight_box[0]), .A3(n367), .A4(
        conv_weight_box[4]), .Y(n372) );
  AO22X1_HVT U594 ( .A1(n370), .A2(conv_weight_box[128]), .A3(n369), .A4(
        conv_weight_box[76]), .Y(n371) );
  NOR3X0_HVT U595 ( .A1(n373), .A2(n372), .A3(n371), .Y(n401) );
  AO22X1_HVT U596 ( .A1(n381), .A2(conv_weight_box[44]), .A3(n380), .A4(
        conv_weight_box[172]), .Y(n379) );
  AO22X1_HVT U597 ( .A1(n383), .A2(conv_weight_box[28]), .A3(n382), .A4(
        conv_weight_box[188]), .Y(n378) );
  AO22X1_HVT U598 ( .A1(n385), .A2(conv_weight_box[140]), .A3(n384), .A4(
        conv_weight_box[156]), .Y(n376) );
  AO22X1_HVT U599 ( .A1(n387), .A2(conv_weight_box[108]), .A3(n386), .A4(
        conv_weight_box[60]), .Y(n375) );
  AO22X1_HVT U600 ( .A1(n389), .A2(conv_weight_box[92]), .A3(n388), .A4(
        conv_weight_box[124]), .Y(n374) );
  OR3X1_HVT U601 ( .A1(n376), .A2(n375), .A3(n374), .Y(n377) );
  OR3X1_HVT U602 ( .A1(n379), .A2(n378), .A3(n377), .Y(n398) );
  AO22X1_HVT U603 ( .A1(n381), .A2(conv_weight_box[40]), .A3(n380), .A4(
        conv_weight_box[168]), .Y(n395) );
  AO22X1_HVT U604 ( .A1(n383), .A2(conv_weight_box[24]), .A3(n382), .A4(
        conv_weight_box[184]), .Y(n394) );
  AO22X1_HVT U605 ( .A1(n385), .A2(conv_weight_box[136]), .A3(n384), .A4(
        conv_weight_box[152]), .Y(n392) );
  AO22X1_HVT U606 ( .A1(n387), .A2(conv_weight_box[104]), .A3(n386), .A4(
        conv_weight_box[56]), .Y(n391) );
  AO22X1_HVT U607 ( .A1(n389), .A2(conv_weight_box[88]), .A3(n388), .A4(
        conv_weight_box[120]), .Y(n390) );
  OR3X1_HVT U608 ( .A1(n392), .A2(n391), .A3(n390), .Y(n393) );
  OR3X1_HVT U609 ( .A1(n395), .A2(n394), .A3(n393), .Y(n396) );
  AOI22X1_HVT U610 ( .A1(n399), .A2(n398), .A3(n397), .A4(n396), .Y(n400) );
endmodule


module multiply_compare ( clk, srstn, mode, channel, conv1_sram_rdata_weight, 
        conv2_sram_rdata_weight, src_window, data_out );
  input [1:0] mode;
  input [4:0] channel;
  input [99:0] conv1_sram_rdata_weight;
  input [99:0] conv2_sram_rdata_weight;
  input [287:0] src_window;
  output [31:0] data_out;
  input clk, srstn;
  wire   N7, N9, DP_OP_425J2_127_3477_n3066, DP_OP_425J2_127_3477_n3065,
         DP_OP_425J2_127_3477_n3063, DP_OP_425J2_127_3477_n3062,
         DP_OP_425J2_127_3477_n3061, DP_OP_425J2_127_3477_n3060,
         DP_OP_425J2_127_3477_n3059, DP_OP_425J2_127_3477_n3058,
         DP_OP_425J2_127_3477_n3057, DP_OP_425J2_127_3477_n3056,
         DP_OP_425J2_127_3477_n3055, DP_OP_425J2_127_3477_n3054,
         DP_OP_425J2_127_3477_n3053, DP_OP_425J2_127_3477_n3052,
         DP_OP_425J2_127_3477_n3051, DP_OP_425J2_127_3477_n3050,
         DP_OP_425J2_127_3477_n3049, DP_OP_425J2_127_3477_n3048,
         DP_OP_425J2_127_3477_n3047, DP_OP_425J2_127_3477_n3046,
         DP_OP_425J2_127_3477_n3045, DP_OP_425J2_127_3477_n3044,
         DP_OP_425J2_127_3477_n3043, DP_OP_425J2_127_3477_n3042,
         DP_OP_425J2_127_3477_n3041, DP_OP_425J2_127_3477_n3040,
         DP_OP_425J2_127_3477_n3039, DP_OP_425J2_127_3477_n3038,
         DP_OP_425J2_127_3477_n3037, DP_OP_425J2_127_3477_n3036,
         DP_OP_425J2_127_3477_n3035, DP_OP_425J2_127_3477_n3034,
         DP_OP_425J2_127_3477_n3033, DP_OP_425J2_127_3477_n3032,
         DP_OP_425J2_127_3477_n3031, DP_OP_425J2_127_3477_n3030,
         DP_OP_425J2_127_3477_n3029, DP_OP_425J2_127_3477_n3028,
         DP_OP_425J2_127_3477_n3027, DP_OP_425J2_127_3477_n3026,
         DP_OP_425J2_127_3477_n3025, DP_OP_425J2_127_3477_n3024,
         DP_OP_425J2_127_3477_n3023, DP_OP_425J2_127_3477_n3021,
         DP_OP_425J2_127_3477_n3020, DP_OP_425J2_127_3477_n3019,
         DP_OP_425J2_127_3477_n3013, DP_OP_425J2_127_3477_n3012,
         DP_OP_425J2_127_3477_n3011, DP_OP_425J2_127_3477_n3010,
         DP_OP_425J2_127_3477_n3009, DP_OP_425J2_127_3477_n3008,
         DP_OP_425J2_127_3477_n3007, DP_OP_425J2_127_3477_n3006,
         DP_OP_425J2_127_3477_n3005, DP_OP_425J2_127_3477_n3004,
         DP_OP_425J2_127_3477_n3003, DP_OP_425J2_127_3477_n3002,
         DP_OP_425J2_127_3477_n3001, DP_OP_425J2_127_3477_n3000,
         DP_OP_425J2_127_3477_n2999, DP_OP_425J2_127_3477_n2998,
         DP_OP_425J2_127_3477_n2997, DP_OP_425J2_127_3477_n2996,
         DP_OP_425J2_127_3477_n2995, DP_OP_425J2_127_3477_n2994,
         DP_OP_425J2_127_3477_n2993, DP_OP_425J2_127_3477_n2992,
         DP_OP_425J2_127_3477_n2991, DP_OP_425J2_127_3477_n2990,
         DP_OP_425J2_127_3477_n2989, DP_OP_425J2_127_3477_n2988,
         DP_OP_425J2_127_3477_n2987, DP_OP_425J2_127_3477_n2986,
         DP_OP_425J2_127_3477_n2985, DP_OP_425J2_127_3477_n2984,
         DP_OP_425J2_127_3477_n2983, DP_OP_425J2_127_3477_n2982,
         DP_OP_425J2_127_3477_n2981, DP_OP_425J2_127_3477_n2980,
         DP_OP_425J2_127_3477_n2977, DP_OP_425J2_127_3477_n2976,
         DP_OP_425J2_127_3477_n2974, DP_OP_425J2_127_3477_n2973,
         DP_OP_425J2_127_3477_n2972, DP_OP_425J2_127_3477_n2971,
         DP_OP_425J2_127_3477_n2970, DP_OP_425J2_127_3477_n2969,
         DP_OP_425J2_127_3477_n2968, DP_OP_425J2_127_3477_n2967,
         DP_OP_425J2_127_3477_n2966, DP_OP_425J2_127_3477_n2965,
         DP_OP_425J2_127_3477_n2964, DP_OP_425J2_127_3477_n2963,
         DP_OP_425J2_127_3477_n2962, DP_OP_425J2_127_3477_n2961,
         DP_OP_425J2_127_3477_n2960, DP_OP_425J2_127_3477_n2959,
         DP_OP_425J2_127_3477_n2958, DP_OP_425J2_127_3477_n2957,
         DP_OP_425J2_127_3477_n2956, DP_OP_425J2_127_3477_n2955,
         DP_OP_425J2_127_3477_n2954, DP_OP_425J2_127_3477_n2953,
         DP_OP_425J2_127_3477_n2951, DP_OP_425J2_127_3477_n2950,
         DP_OP_425J2_127_3477_n2949, DP_OP_425J2_127_3477_n2948,
         DP_OP_425J2_127_3477_n2947, DP_OP_425J2_127_3477_n2946,
         DP_OP_425J2_127_3477_n2945, DP_OP_425J2_127_3477_n2944,
         DP_OP_425J2_127_3477_n2943, DP_OP_425J2_127_3477_n2942,
         DP_OP_425J2_127_3477_n2941, DP_OP_425J2_127_3477_n2940,
         DP_OP_425J2_127_3477_n2939, DP_OP_425J2_127_3477_n2938,
         DP_OP_425J2_127_3477_n2935, DP_OP_425J2_127_3477_n2933,
         DP_OP_425J2_127_3477_n2925, DP_OP_425J2_127_3477_n2924,
         DP_OP_425J2_127_3477_n2923, DP_OP_425J2_127_3477_n2922,
         DP_OP_425J2_127_3477_n2921, DP_OP_425J2_127_3477_n2920,
         DP_OP_425J2_127_3477_n2919, DP_OP_425J2_127_3477_n2918,
         DP_OP_425J2_127_3477_n2917, DP_OP_425J2_127_3477_n2916,
         DP_OP_425J2_127_3477_n2915, DP_OP_425J2_127_3477_n2914,
         DP_OP_425J2_127_3477_n2913, DP_OP_425J2_127_3477_n2912,
         DP_OP_425J2_127_3477_n2911, DP_OP_425J2_127_3477_n2910,
         DP_OP_425J2_127_3477_n2909, DP_OP_425J2_127_3477_n2908,
         DP_OP_425J2_127_3477_n2907, DP_OP_425J2_127_3477_n2906,
         DP_OP_425J2_127_3477_n2905, DP_OP_425J2_127_3477_n2904,
         DP_OP_425J2_127_3477_n2903, DP_OP_425J2_127_3477_n2902,
         DP_OP_425J2_127_3477_n2901, DP_OP_425J2_127_3477_n2900,
         DP_OP_425J2_127_3477_n2899, DP_OP_425J2_127_3477_n2898,
         DP_OP_425J2_127_3477_n2897, DP_OP_425J2_127_3477_n2896,
         DP_OP_425J2_127_3477_n2895, DP_OP_425J2_127_3477_n2894,
         DP_OP_425J2_127_3477_n2893, DP_OP_425J2_127_3477_n2891,
         DP_OP_425J2_127_3477_n2888, DP_OP_425J2_127_3477_n2886,
         DP_OP_425J2_127_3477_n2885, DP_OP_425J2_127_3477_n2883,
         DP_OP_425J2_127_3477_n2882, DP_OP_425J2_127_3477_n2881,
         DP_OP_425J2_127_3477_n2880, DP_OP_425J2_127_3477_n2879,
         DP_OP_425J2_127_3477_n2878, DP_OP_425J2_127_3477_n2877,
         DP_OP_425J2_127_3477_n2876, DP_OP_425J2_127_3477_n2875,
         DP_OP_425J2_127_3477_n2874, DP_OP_425J2_127_3477_n2873,
         DP_OP_425J2_127_3477_n2872, DP_OP_425J2_127_3477_n2871,
         DP_OP_425J2_127_3477_n2870, DP_OP_425J2_127_3477_n2869,
         DP_OP_425J2_127_3477_n2868, DP_OP_425J2_127_3477_n2867,
         DP_OP_425J2_127_3477_n2866, DP_OP_425J2_127_3477_n2865,
         DP_OP_425J2_127_3477_n2864, DP_OP_425J2_127_3477_n2863,
         DP_OP_425J2_127_3477_n2862, DP_OP_425J2_127_3477_n2861,
         DP_OP_425J2_127_3477_n2860, DP_OP_425J2_127_3477_n2859,
         DP_OP_425J2_127_3477_n2858, DP_OP_425J2_127_3477_n2857,
         DP_OP_425J2_127_3477_n2856, DP_OP_425J2_127_3477_n2855,
         DP_OP_425J2_127_3477_n2854, DP_OP_425J2_127_3477_n2853,
         DP_OP_425J2_127_3477_n2852, DP_OP_425J2_127_3477_n2851,
         DP_OP_425J2_127_3477_n2850, DP_OP_425J2_127_3477_n2848,
         DP_OP_425J2_127_3477_n2847, DP_OP_425J2_127_3477_n2846,
         DP_OP_425J2_127_3477_n2843, DP_OP_425J2_127_3477_n2841,
         DP_OP_425J2_127_3477_n2840, DP_OP_425J2_127_3477_n2839,
         DP_OP_425J2_127_3477_n2837, DP_OP_425J2_127_3477_n2836,
         DP_OP_425J2_127_3477_n2835, DP_OP_425J2_127_3477_n2834,
         DP_OP_425J2_127_3477_n2833, DP_OP_425J2_127_3477_n2832,
         DP_OP_425J2_127_3477_n2831, DP_OP_425J2_127_3477_n2830,
         DP_OP_425J2_127_3477_n2829, DP_OP_425J2_127_3477_n2828,
         DP_OP_425J2_127_3477_n2827, DP_OP_425J2_127_3477_n2826,
         DP_OP_425J2_127_3477_n2825, DP_OP_425J2_127_3477_n2824,
         DP_OP_425J2_127_3477_n2823, DP_OP_425J2_127_3477_n2822,
         DP_OP_425J2_127_3477_n2821, DP_OP_425J2_127_3477_n2820,
         DP_OP_425J2_127_3477_n2819, DP_OP_425J2_127_3477_n2818,
         DP_OP_425J2_127_3477_n2817, DP_OP_425J2_127_3477_n2816,
         DP_OP_425J2_127_3477_n2815, DP_OP_425J2_127_3477_n2814,
         DP_OP_425J2_127_3477_n2813, DP_OP_425J2_127_3477_n2812,
         DP_OP_425J2_127_3477_n2811, DP_OP_425J2_127_3477_n2810,
         DP_OP_425J2_127_3477_n2809, DP_OP_425J2_127_3477_n2808,
         DP_OP_425J2_127_3477_n2807, DP_OP_425J2_127_3477_n2806,
         DP_OP_425J2_127_3477_n2801, DP_OP_425J2_127_3477_n2800,
         DP_OP_425J2_127_3477_n2799, DP_OP_425J2_127_3477_n2798,
         DP_OP_425J2_127_3477_n2797, DP_OP_425J2_127_3477_n2796,
         DP_OP_425J2_127_3477_n2793, DP_OP_425J2_127_3477_n2792,
         DP_OP_425J2_127_3477_n2791, DP_OP_425J2_127_3477_n2790,
         DP_OP_425J2_127_3477_n2789, DP_OP_425J2_127_3477_n2788,
         DP_OP_425J2_127_3477_n2787, DP_OP_425J2_127_3477_n2786,
         DP_OP_425J2_127_3477_n2785, DP_OP_425J2_127_3477_n2784,
         DP_OP_425J2_127_3477_n2783, DP_OP_425J2_127_3477_n2782,
         DP_OP_425J2_127_3477_n2781, DP_OP_425J2_127_3477_n2780,
         DP_OP_425J2_127_3477_n2779, DP_OP_425J2_127_3477_n2778,
         DP_OP_425J2_127_3477_n2777, DP_OP_425J2_127_3477_n2776,
         DP_OP_425J2_127_3477_n2775, DP_OP_425J2_127_3477_n2774,
         DP_OP_425J2_127_3477_n2773, DP_OP_425J2_127_3477_n2772,
         DP_OP_425J2_127_3477_n2771, DP_OP_425J2_127_3477_n2770,
         DP_OP_425J2_127_3477_n2769, DP_OP_425J2_127_3477_n2768,
         DP_OP_425J2_127_3477_n2767, DP_OP_425J2_127_3477_n2766,
         DP_OP_425J2_127_3477_n2765, DP_OP_425J2_127_3477_n2764,
         DP_OP_425J2_127_3477_n2763, DP_OP_425J2_127_3477_n2762,
         DP_OP_425J2_127_3477_n2761, DP_OP_425J2_127_3477_n2760,
         DP_OP_425J2_127_3477_n2756, DP_OP_425J2_127_3477_n2755,
         DP_OP_425J2_127_3477_n2754, DP_OP_425J2_127_3477_n2749,
         DP_OP_425J2_127_3477_n2748, DP_OP_425J2_127_3477_n2747,
         DP_OP_425J2_127_3477_n2746, DP_OP_425J2_127_3477_n2745,
         DP_OP_425J2_127_3477_n2744, DP_OP_425J2_127_3477_n2743,
         DP_OP_425J2_127_3477_n2742, DP_OP_425J2_127_3477_n2741,
         DP_OP_425J2_127_3477_n2740, DP_OP_425J2_127_3477_n2739,
         DP_OP_425J2_127_3477_n2738, DP_OP_425J2_127_3477_n2737,
         DP_OP_425J2_127_3477_n2736, DP_OP_425J2_127_3477_n2735,
         DP_OP_425J2_127_3477_n2734, DP_OP_425J2_127_3477_n2733,
         DP_OP_425J2_127_3477_n2732, DP_OP_425J2_127_3477_n2731,
         DP_OP_425J2_127_3477_n2730, DP_OP_425J2_127_3477_n2729,
         DP_OP_425J2_127_3477_n2728, DP_OP_425J2_127_3477_n2727,
         DP_OP_425J2_127_3477_n2726, DP_OP_425J2_127_3477_n2725,
         DP_OP_425J2_127_3477_n2724, DP_OP_425J2_127_3477_n2723,
         DP_OP_425J2_127_3477_n2722, DP_OP_425J2_127_3477_n2721,
         DP_OP_425J2_127_3477_n2720, DP_OP_425J2_127_3477_n2719,
         DP_OP_425J2_127_3477_n2718, DP_OP_425J2_127_3477_n2714,
         DP_OP_425J2_127_3477_n2712, DP_OP_425J2_127_3477_n2710,
         DP_OP_425J2_127_3477_n2708, DP_OP_425J2_127_3477_n2705,
         DP_OP_425J2_127_3477_n2704, DP_OP_425J2_127_3477_n2703,
         DP_OP_425J2_127_3477_n2702, DP_OP_425J2_127_3477_n2701,
         DP_OP_425J2_127_3477_n2700, DP_OP_425J2_127_3477_n2699,
         DP_OP_425J2_127_3477_n2698, DP_OP_425J2_127_3477_n2697,
         DP_OP_425J2_127_3477_n2696, DP_OP_425J2_127_3477_n2695,
         DP_OP_425J2_127_3477_n2694, DP_OP_425J2_127_3477_n2693,
         DP_OP_425J2_127_3477_n2692, DP_OP_425J2_127_3477_n2691,
         DP_OP_425J2_127_3477_n2690, DP_OP_425J2_127_3477_n2689,
         DP_OP_425J2_127_3477_n2688, DP_OP_425J2_127_3477_n2687,
         DP_OP_425J2_127_3477_n2686, DP_OP_425J2_127_3477_n2685,
         DP_OP_425J2_127_3477_n2684, DP_OP_425J2_127_3477_n2683,
         DP_OP_425J2_127_3477_n2682, DP_OP_425J2_127_3477_n2681,
         DP_OP_425J2_127_3477_n2680, DP_OP_425J2_127_3477_n2679,
         DP_OP_425J2_127_3477_n2678, DP_OP_425J2_127_3477_n2677,
         DP_OP_425J2_127_3477_n2676, DP_OP_425J2_127_3477_n2675,
         DP_OP_425J2_127_3477_n2674, DP_OP_425J2_127_3477_n2673,
         DP_OP_425J2_127_3477_n2671, DP_OP_425J2_127_3477_n2661,
         DP_OP_425J2_127_3477_n2660, DP_OP_425J2_127_3477_n2659,
         DP_OP_425J2_127_3477_n2658, DP_OP_425J2_127_3477_n2657,
         DP_OP_425J2_127_3477_n2656, DP_OP_425J2_127_3477_n2655,
         DP_OP_425J2_127_3477_n2654, DP_OP_425J2_127_3477_n2653,
         DP_OP_425J2_127_3477_n2652, DP_OP_425J2_127_3477_n2651,
         DP_OP_425J2_127_3477_n2650, DP_OP_425J2_127_3477_n2649,
         DP_OP_425J2_127_3477_n2648, DP_OP_425J2_127_3477_n2647,
         DP_OP_425J2_127_3477_n2646, DP_OP_425J2_127_3477_n2645,
         DP_OP_425J2_127_3477_n2644, DP_OP_425J2_127_3477_n2643,
         DP_OP_425J2_127_3477_n2642, DP_OP_425J2_127_3477_n2641,
         DP_OP_425J2_127_3477_n2640, DP_OP_425J2_127_3477_n2639,
         DP_OP_425J2_127_3477_n2638, DP_OP_425J2_127_3477_n2637,
         DP_OP_425J2_127_3477_n2636, DP_OP_425J2_127_3477_n2635,
         DP_OP_425J2_127_3477_n2634, DP_OP_425J2_127_3477_n2633,
         DP_OP_425J2_127_3477_n2632, DP_OP_425J2_127_3477_n2631,
         DP_OP_425J2_127_3477_n2630, DP_OP_425J2_127_3477_n2622,
         DP_OP_425J2_127_3477_n2621, DP_OP_425J2_127_3477_n2620,
         DP_OP_425J2_127_3477_n2617, DP_OP_425J2_127_3477_n2616,
         DP_OP_425J2_127_3477_n2615, DP_OP_425J2_127_3477_n2614,
         DP_OP_425J2_127_3477_n2613, DP_OP_425J2_127_3477_n2612,
         DP_OP_425J2_127_3477_n2611, DP_OP_425J2_127_3477_n2610,
         DP_OP_425J2_127_3477_n2609, DP_OP_425J2_127_3477_n2608,
         DP_OP_425J2_127_3477_n2607, DP_OP_425J2_127_3477_n2606,
         DP_OP_425J2_127_3477_n2605, DP_OP_425J2_127_3477_n2604,
         DP_OP_425J2_127_3477_n2603, DP_OP_425J2_127_3477_n2602,
         DP_OP_425J2_127_3477_n2601, DP_OP_425J2_127_3477_n2600,
         DP_OP_425J2_127_3477_n2599, DP_OP_425J2_127_3477_n2598,
         DP_OP_425J2_127_3477_n2597, DP_OP_425J2_127_3477_n2596,
         DP_OP_425J2_127_3477_n2595, DP_OP_425J2_127_3477_n2594,
         DP_OP_425J2_127_3477_n2593, DP_OP_425J2_127_3477_n2592,
         DP_OP_425J2_127_3477_n2591, DP_OP_425J2_127_3477_n2590,
         DP_OP_425J2_127_3477_n2589, DP_OP_425J2_127_3477_n2588,
         DP_OP_425J2_127_3477_n2587, DP_OP_425J2_127_3477_n2586,
         DP_OP_425J2_127_3477_n2582, DP_OP_425J2_127_3477_n2581,
         DP_OP_425J2_127_3477_n2580, DP_OP_425J2_127_3477_n2579,
         DP_OP_425J2_127_3477_n2578, DP_OP_425J2_127_3477_n2577,
         DP_OP_425J2_127_3477_n2576, DP_OP_425J2_127_3477_n2574,
         DP_OP_425J2_127_3477_n2573, DP_OP_425J2_127_3477_n2572,
         DP_OP_425J2_127_3477_n2571, DP_OP_425J2_127_3477_n2569,
         DP_OP_425J2_127_3477_n2568, DP_OP_425J2_127_3477_n2567,
         DP_OP_425J2_127_3477_n2566, DP_OP_425J2_127_3477_n2565,
         DP_OP_425J2_127_3477_n2564, DP_OP_425J2_127_3477_n2563,
         DP_OP_425J2_127_3477_n2562, DP_OP_425J2_127_3477_n2561,
         DP_OP_425J2_127_3477_n2560, DP_OP_425J2_127_3477_n2559,
         DP_OP_425J2_127_3477_n2558, DP_OP_425J2_127_3477_n2557,
         DP_OP_425J2_127_3477_n2556, DP_OP_425J2_127_3477_n2555,
         DP_OP_425J2_127_3477_n2554, DP_OP_425J2_127_3477_n2553,
         DP_OP_425J2_127_3477_n2552, DP_OP_425J2_127_3477_n2551,
         DP_OP_425J2_127_3477_n2550, DP_OP_425J2_127_3477_n2549,
         DP_OP_425J2_127_3477_n2548, DP_OP_425J2_127_3477_n2547,
         DP_OP_425J2_127_3477_n2546, DP_OP_425J2_127_3477_n2545,
         DP_OP_425J2_127_3477_n2544, DP_OP_425J2_127_3477_n2543,
         DP_OP_425J2_127_3477_n2542, DP_OP_425J2_127_3477_n2541,
         DP_OP_425J2_127_3477_n2539, DP_OP_425J2_127_3477_n2536,
         DP_OP_425J2_127_3477_n2534, DP_OP_425J2_127_3477_n2529,
         DP_OP_425J2_127_3477_n2528, DP_OP_425J2_127_3477_n2527,
         DP_OP_425J2_127_3477_n2526, DP_OP_425J2_127_3477_n2525,
         DP_OP_425J2_127_3477_n2524, DP_OP_425J2_127_3477_n2523,
         DP_OP_425J2_127_3477_n2522, DP_OP_425J2_127_3477_n2521,
         DP_OP_425J2_127_3477_n2520, DP_OP_425J2_127_3477_n2519,
         DP_OP_425J2_127_3477_n2518, DP_OP_425J2_127_3477_n2517,
         DP_OP_425J2_127_3477_n2516, DP_OP_425J2_127_3477_n2515,
         DP_OP_425J2_127_3477_n2514, DP_OP_425J2_127_3477_n2513,
         DP_OP_425J2_127_3477_n2512, DP_OP_425J2_127_3477_n2511,
         DP_OP_425J2_127_3477_n2510, DP_OP_425J2_127_3477_n2509,
         DP_OP_425J2_127_3477_n2508, DP_OP_425J2_127_3477_n2507,
         DP_OP_425J2_127_3477_n2506, DP_OP_425J2_127_3477_n2505,
         DP_OP_425J2_127_3477_n2504, DP_OP_425J2_127_3477_n2503,
         DP_OP_425J2_127_3477_n2502, DP_OP_425J2_127_3477_n2501,
         DP_OP_425J2_127_3477_n2500, DP_OP_425J2_127_3477_n2499,
         DP_OP_425J2_127_3477_n2498, DP_OP_425J2_127_3477_n2497,
         DP_OP_425J2_127_3477_n2495, DP_OP_425J2_127_3477_n2493,
         DP_OP_425J2_127_3477_n2485, DP_OP_425J2_127_3477_n2484,
         DP_OP_425J2_127_3477_n2483, DP_OP_425J2_127_3477_n2482,
         DP_OP_425J2_127_3477_n2481, DP_OP_425J2_127_3477_n2480,
         DP_OP_425J2_127_3477_n2479, DP_OP_425J2_127_3477_n2478,
         DP_OP_425J2_127_3477_n2477, DP_OP_425J2_127_3477_n2476,
         DP_OP_425J2_127_3477_n2475, DP_OP_425J2_127_3477_n2474,
         DP_OP_425J2_127_3477_n2473, DP_OP_425J2_127_3477_n2472,
         DP_OP_425J2_127_3477_n2471, DP_OP_425J2_127_3477_n2470,
         DP_OP_425J2_127_3477_n2469, DP_OP_425J2_127_3477_n2468,
         DP_OP_425J2_127_3477_n2467, DP_OP_425J2_127_3477_n2466,
         DP_OP_425J2_127_3477_n2465, DP_OP_425J2_127_3477_n2464,
         DP_OP_425J2_127_3477_n2463, DP_OP_425J2_127_3477_n2462,
         DP_OP_425J2_127_3477_n2461, DP_OP_425J2_127_3477_n2460,
         DP_OP_425J2_127_3477_n2459, DP_OP_425J2_127_3477_n2458,
         DP_OP_425J2_127_3477_n2457, DP_OP_425J2_127_3477_n2456,
         DP_OP_425J2_127_3477_n2455, DP_OP_425J2_127_3477_n2454,
         DP_OP_425J2_127_3477_n2453, DP_OP_425J2_127_3477_n2449,
         DP_OP_425J2_127_3477_n2448, DP_OP_425J2_127_3477_n2447,
         DP_OP_425J2_127_3477_n2445, DP_OP_425J2_127_3477_n2441,
         DP_OP_425J2_127_3477_n2440, DP_OP_425J2_127_3477_n2439,
         DP_OP_425J2_127_3477_n2438, DP_OP_425J2_127_3477_n2437,
         DP_OP_425J2_127_3477_n2436, DP_OP_425J2_127_3477_n2435,
         DP_OP_425J2_127_3477_n2434, DP_OP_425J2_127_3477_n2433,
         DP_OP_425J2_127_3477_n2432, DP_OP_425J2_127_3477_n2431,
         DP_OP_425J2_127_3477_n2430, DP_OP_425J2_127_3477_n2429,
         DP_OP_425J2_127_3477_n2428, DP_OP_425J2_127_3477_n2427,
         DP_OP_425J2_127_3477_n2426, DP_OP_425J2_127_3477_n2425,
         DP_OP_425J2_127_3477_n2424, DP_OP_425J2_127_3477_n2423,
         DP_OP_425J2_127_3477_n2422, DP_OP_425J2_127_3477_n2421,
         DP_OP_425J2_127_3477_n2420, DP_OP_425J2_127_3477_n2419,
         DP_OP_425J2_127_3477_n2418, DP_OP_425J2_127_3477_n2417,
         DP_OP_425J2_127_3477_n2416, DP_OP_425J2_127_3477_n2415,
         DP_OP_425J2_127_3477_n2414, DP_OP_425J2_127_3477_n2413,
         DP_OP_425J2_127_3477_n2412, DP_OP_425J2_127_3477_n2411,
         DP_OP_425J2_127_3477_n2410, DP_OP_425J2_127_3477_n2409,
         DP_OP_425J2_127_3477_n2404, DP_OP_425J2_127_3477_n2403,
         DP_OP_425J2_127_3477_n2401, DP_OP_425J2_127_3477_n2400,
         DP_OP_425J2_127_3477_n2397, DP_OP_425J2_127_3477_n2396,
         DP_OP_425J2_127_3477_n2395, DP_OP_425J2_127_3477_n2394,
         DP_OP_425J2_127_3477_n2393, DP_OP_425J2_127_3477_n2392,
         DP_OP_425J2_127_3477_n2391, DP_OP_425J2_127_3477_n2390,
         DP_OP_425J2_127_3477_n2389, DP_OP_425J2_127_3477_n2388,
         DP_OP_425J2_127_3477_n2387, DP_OP_425J2_127_3477_n2386,
         DP_OP_425J2_127_3477_n2385, DP_OP_425J2_127_3477_n2384,
         DP_OP_425J2_127_3477_n2383, DP_OP_425J2_127_3477_n2382,
         DP_OP_425J2_127_3477_n2381, DP_OP_425J2_127_3477_n2379,
         DP_OP_425J2_127_3477_n2378, DP_OP_425J2_127_3477_n2377,
         DP_OP_425J2_127_3477_n2376, DP_OP_425J2_127_3477_n2375,
         DP_OP_425J2_127_3477_n2374, DP_OP_425J2_127_3477_n2373,
         DP_OP_425J2_127_3477_n2372, DP_OP_425J2_127_3477_n2371,
         DP_OP_425J2_127_3477_n2370, DP_OP_425J2_127_3477_n2369,
         DP_OP_425J2_127_3477_n2368, DP_OP_425J2_127_3477_n2367,
         DP_OP_425J2_127_3477_n2366, DP_OP_425J2_127_3477_n2365,
         DP_OP_425J2_127_3477_n2359, DP_OP_425J2_127_3477_n2358,
         DP_OP_425J2_127_3477_n2357, DP_OP_425J2_127_3477_n2356,
         DP_OP_425J2_127_3477_n2353, DP_OP_425J2_127_3477_n2352,
         DP_OP_425J2_127_3477_n2351, DP_OP_425J2_127_3477_n2350,
         DP_OP_425J2_127_3477_n2349, DP_OP_425J2_127_3477_n2348,
         DP_OP_425J2_127_3477_n2347, DP_OP_425J2_127_3477_n2346,
         DP_OP_425J2_127_3477_n2345, DP_OP_425J2_127_3477_n2344,
         DP_OP_425J2_127_3477_n2343, DP_OP_425J2_127_3477_n2342,
         DP_OP_425J2_127_3477_n2341, DP_OP_425J2_127_3477_n2340,
         DP_OP_425J2_127_3477_n2339, DP_OP_425J2_127_3477_n2338,
         DP_OP_425J2_127_3477_n2337, DP_OP_425J2_127_3477_n2336,
         DP_OP_425J2_127_3477_n2335, DP_OP_425J2_127_3477_n2334,
         DP_OP_425J2_127_3477_n2333, DP_OP_425J2_127_3477_n2332,
         DP_OP_425J2_127_3477_n2331, DP_OP_425J2_127_3477_n2330,
         DP_OP_425J2_127_3477_n2329, DP_OP_425J2_127_3477_n2328,
         DP_OP_425J2_127_3477_n2327, DP_OP_425J2_127_3477_n2326,
         DP_OP_425J2_127_3477_n2325, DP_OP_425J2_127_3477_n2324,
         DP_OP_425J2_127_3477_n2323, DP_OP_425J2_127_3477_n2322,
         DP_OP_425J2_127_3477_n2321, DP_OP_425J2_127_3477_n2320,
         DP_OP_425J2_127_3477_n2319, DP_OP_425J2_127_3477_n2312,
         DP_OP_425J2_127_3477_n2311, DP_OP_425J2_127_3477_n2310,
         DP_OP_425J2_127_3477_n2309, DP_OP_425J2_127_3477_n2308,
         DP_OP_425J2_127_3477_n2307, DP_OP_425J2_127_3477_n2306,
         DP_OP_425J2_127_3477_n2305, DP_OP_425J2_127_3477_n2304,
         DP_OP_425J2_127_3477_n2303, DP_OP_425J2_127_3477_n2302,
         DP_OP_425J2_127_3477_n2301, DP_OP_425J2_127_3477_n2300,
         DP_OP_425J2_127_3477_n2299, DP_OP_425J2_127_3477_n2298,
         DP_OP_425J2_127_3477_n2297, DP_OP_425J2_127_3477_n2296,
         DP_OP_425J2_127_3477_n2295, DP_OP_425J2_127_3477_n2294,
         DP_OP_425J2_127_3477_n2293, DP_OP_425J2_127_3477_n2292,
         DP_OP_425J2_127_3477_n2291, DP_OP_425J2_127_3477_n2290,
         DP_OP_425J2_127_3477_n2289, DP_OP_425J2_127_3477_n2288,
         DP_OP_425J2_127_3477_n2287, DP_OP_425J2_127_3477_n2286,
         DP_OP_425J2_127_3477_n2285, DP_OP_425J2_127_3477_n2284,
         DP_OP_425J2_127_3477_n2283, DP_OP_425J2_127_3477_n2282,
         DP_OP_425J2_127_3477_n2281, DP_OP_425J2_127_3477_n2280,
         DP_OP_425J2_127_3477_n2279, DP_OP_425J2_127_3477_n2278,
         DP_OP_425J2_127_3477_n2272, DP_OP_425J2_127_3477_n2269,
         DP_OP_425J2_127_3477_n2268, DP_OP_425J2_127_3477_n2265,
         DP_OP_425J2_127_3477_n2264, DP_OP_425J2_127_3477_n2263,
         DP_OP_425J2_127_3477_n2262, DP_OP_425J2_127_3477_n2261,
         DP_OP_425J2_127_3477_n2260, DP_OP_425J2_127_3477_n2259,
         DP_OP_425J2_127_3477_n2258, DP_OP_425J2_127_3477_n2257,
         DP_OP_425J2_127_3477_n2256, DP_OP_425J2_127_3477_n2255,
         DP_OP_425J2_127_3477_n2254, DP_OP_425J2_127_3477_n2253,
         DP_OP_425J2_127_3477_n2252, DP_OP_425J2_127_3477_n2251,
         DP_OP_425J2_127_3477_n2250, DP_OP_425J2_127_3477_n2249,
         DP_OP_425J2_127_3477_n2248, DP_OP_425J2_127_3477_n2247,
         DP_OP_425J2_127_3477_n2246, DP_OP_425J2_127_3477_n2245,
         DP_OP_425J2_127_3477_n2244, DP_OP_425J2_127_3477_n2243,
         DP_OP_425J2_127_3477_n2242, DP_OP_425J2_127_3477_n2241,
         DP_OP_425J2_127_3477_n2240, DP_OP_425J2_127_3477_n2239,
         DP_OP_425J2_127_3477_n2238, DP_OP_425J2_127_3477_n2237,
         DP_OP_425J2_127_3477_n2236, DP_OP_425J2_127_3477_n2235,
         DP_OP_425J2_127_3477_n2234, DP_OP_425J2_127_3477_n2231,
         DP_OP_425J2_127_3477_n2230, DP_OP_425J2_127_3477_n2226,
         DP_OP_425J2_127_3477_n2221, DP_OP_425J2_127_3477_n2220,
         DP_OP_425J2_127_3477_n2219, DP_OP_425J2_127_3477_n2218,
         DP_OP_425J2_127_3477_n2217, DP_OP_425J2_127_3477_n2216,
         DP_OP_425J2_127_3477_n2215, DP_OP_425J2_127_3477_n2214,
         DP_OP_425J2_127_3477_n2213, DP_OP_425J2_127_3477_n2212,
         DP_OP_425J2_127_3477_n2211, DP_OP_425J2_127_3477_n2210,
         DP_OP_425J2_127_3477_n2209, DP_OP_425J2_127_3477_n2208,
         DP_OP_425J2_127_3477_n2207, DP_OP_425J2_127_3477_n2206,
         DP_OP_425J2_127_3477_n2205, DP_OP_425J2_127_3477_n2204,
         DP_OP_425J2_127_3477_n2203, DP_OP_425J2_127_3477_n2202,
         DP_OP_425J2_127_3477_n2201, DP_OP_425J2_127_3477_n2200,
         DP_OP_425J2_127_3477_n2199, DP_OP_425J2_127_3477_n2198,
         DP_OP_425J2_127_3477_n2197, DP_OP_425J2_127_3477_n2196,
         DP_OP_425J2_127_3477_n2195, DP_OP_425J2_127_3477_n2194,
         DP_OP_425J2_127_3477_n2193, DP_OP_425J2_127_3477_n2192,
         DP_OP_425J2_127_3477_n2191, DP_OP_425J2_127_3477_n2190,
         DP_OP_425J2_127_3477_n2189, DP_OP_425J2_127_3477_n2188,
         DP_OP_425J2_127_3477_n2186, DP_OP_425J2_127_3477_n2185,
         DP_OP_425J2_127_3477_n2184, DP_OP_425J2_127_3477_n2182,
         DP_OP_425J2_127_3477_n2180, DP_OP_425J2_127_3477_n2177,
         DP_OP_425J2_127_3477_n2176, DP_OP_425J2_127_3477_n2175,
         DP_OP_425J2_127_3477_n2174, DP_OP_425J2_127_3477_n2173,
         DP_OP_425J2_127_3477_n2172, DP_OP_425J2_127_3477_n2171,
         DP_OP_425J2_127_3477_n2170, DP_OP_425J2_127_3477_n2169,
         DP_OP_425J2_127_3477_n2168, DP_OP_425J2_127_3477_n2167,
         DP_OP_425J2_127_3477_n2166, DP_OP_425J2_127_3477_n2165,
         DP_OP_425J2_127_3477_n2164, DP_OP_425J2_127_3477_n2163,
         DP_OP_425J2_127_3477_n2162, DP_OP_425J2_127_3477_n2161,
         DP_OP_425J2_127_3477_n2160, DP_OP_425J2_127_3477_n2159,
         DP_OP_425J2_127_3477_n2158, DP_OP_425J2_127_3477_n2157,
         DP_OP_425J2_127_3477_n2156, DP_OP_425J2_127_3477_n2155,
         DP_OP_425J2_127_3477_n2154, DP_OP_425J2_127_3477_n2153,
         DP_OP_425J2_127_3477_n2152, DP_OP_425J2_127_3477_n2151,
         DP_OP_425J2_127_3477_n2150, DP_OP_425J2_127_3477_n2149,
         DP_OP_425J2_127_3477_n2148, DP_OP_425J2_127_3477_n2147,
         DP_OP_425J2_127_3477_n2146, DP_OP_425J2_127_3477_n2144,
         DP_OP_425J2_127_3477_n2143, DP_OP_425J2_127_3477_n2138,
         DP_OP_425J2_127_3477_n2133, DP_OP_425J2_127_3477_n2132,
         DP_OP_425J2_127_3477_n2131, DP_OP_425J2_127_3477_n2130,
         DP_OP_425J2_127_3477_n2129, DP_OP_425J2_127_3477_n2128,
         DP_OP_425J2_127_3477_n2127, DP_OP_425J2_127_3477_n2126,
         DP_OP_425J2_127_3477_n2125, DP_OP_425J2_127_3477_n2124,
         DP_OP_425J2_127_3477_n2123, DP_OP_425J2_127_3477_n2122,
         DP_OP_425J2_127_3477_n2121, DP_OP_425J2_127_3477_n2120,
         DP_OP_425J2_127_3477_n2119, DP_OP_425J2_127_3477_n2118,
         DP_OP_425J2_127_3477_n2117, DP_OP_425J2_127_3477_n2116,
         DP_OP_425J2_127_3477_n2115, DP_OP_425J2_127_3477_n2114,
         DP_OP_425J2_127_3477_n2113, DP_OP_425J2_127_3477_n2112,
         DP_OP_425J2_127_3477_n2111, DP_OP_425J2_127_3477_n2110,
         DP_OP_425J2_127_3477_n2109, DP_OP_425J2_127_3477_n2108,
         DP_OP_425J2_127_3477_n2107, DP_OP_425J2_127_3477_n2106,
         DP_OP_425J2_127_3477_n2105, DP_OP_425J2_127_3477_n2104,
         DP_OP_425J2_127_3477_n2103, DP_OP_425J2_127_3477_n2102,
         DP_OP_425J2_127_3477_n2099, DP_OP_425J2_127_3477_n2098,
         DP_OP_425J2_127_3477_n2092, DP_OP_425J2_127_3477_n2089,
         DP_OP_425J2_127_3477_n2088, DP_OP_425J2_127_3477_n2087,
         DP_OP_425J2_127_3477_n2086, DP_OP_425J2_127_3477_n2085,
         DP_OP_425J2_127_3477_n2084, DP_OP_425J2_127_3477_n2083,
         DP_OP_425J2_127_3477_n2082, DP_OP_425J2_127_3477_n2081,
         DP_OP_425J2_127_3477_n2080, DP_OP_425J2_127_3477_n2079,
         DP_OP_425J2_127_3477_n2078, DP_OP_425J2_127_3477_n2077,
         DP_OP_425J2_127_3477_n2076, DP_OP_425J2_127_3477_n2075,
         DP_OP_425J2_127_3477_n2074, DP_OP_425J2_127_3477_n2073,
         DP_OP_425J2_127_3477_n2072, DP_OP_425J2_127_3477_n2071,
         DP_OP_425J2_127_3477_n2070, DP_OP_425J2_127_3477_n2069,
         DP_OP_425J2_127_3477_n2068, DP_OP_425J2_127_3477_n2067,
         DP_OP_425J2_127_3477_n2066, DP_OP_425J2_127_3477_n2065,
         DP_OP_425J2_127_3477_n2064, DP_OP_425J2_127_3477_n2063,
         DP_OP_425J2_127_3477_n2062, DP_OP_425J2_127_3477_n2061,
         DP_OP_425J2_127_3477_n2060, DP_OP_425J2_127_3477_n2059,
         DP_OP_425J2_127_3477_n2058, DP_OP_425J2_127_3477_n2057,
         DP_OP_425J2_127_3477_n2056, DP_OP_425J2_127_3477_n2055,
         DP_OP_425J2_127_3477_n2053, DP_OP_425J2_127_3477_n2050,
         DP_OP_425J2_127_3477_n2049, DP_OP_425J2_127_3477_n2048,
         DP_OP_425J2_127_3477_n2046, DP_OP_425J2_127_3477_n2045,
         DP_OP_425J2_127_3477_n2044, DP_OP_425J2_127_3477_n2043,
         DP_OP_425J2_127_3477_n2042, DP_OP_425J2_127_3477_n2041,
         DP_OP_425J2_127_3477_n2040, DP_OP_425J2_127_3477_n2039,
         DP_OP_425J2_127_3477_n2038, DP_OP_425J2_127_3477_n2037,
         DP_OP_425J2_127_3477_n2036, DP_OP_425J2_127_3477_n2035,
         DP_OP_425J2_127_3477_n2034, DP_OP_425J2_127_3477_n2033,
         DP_OP_425J2_127_3477_n2032, DP_OP_425J2_127_3477_n2031,
         DP_OP_425J2_127_3477_n2030, DP_OP_425J2_127_3477_n2029,
         DP_OP_425J2_127_3477_n2028, DP_OP_425J2_127_3477_n2027,
         DP_OP_425J2_127_3477_n2026, DP_OP_425J2_127_3477_n2025,
         DP_OP_425J2_127_3477_n2024, DP_OP_425J2_127_3477_n2023,
         DP_OP_425J2_127_3477_n2022, DP_OP_425J2_127_3477_n2021,
         DP_OP_425J2_127_3477_n2020, DP_OP_425J2_127_3477_n2019,
         DP_OP_425J2_127_3477_n2018, DP_OP_425J2_127_3477_n2017,
         DP_OP_425J2_127_3477_n2016, DP_OP_425J2_127_3477_n2015,
         DP_OP_425J2_127_3477_n2014, DP_OP_425J2_127_3477_n2011,
         DP_OP_425J2_127_3477_n2010, DP_OP_425J2_127_3477_n2008,
         DP_OP_425J2_127_3477_n2007, DP_OP_425J2_127_3477_n2002,
         DP_OP_425J2_127_3477_n2001, DP_OP_425J2_127_3477_n2000,
         DP_OP_425J2_127_3477_n1999, DP_OP_425J2_127_3477_n1998,
         DP_OP_425J2_127_3477_n1997, DP_OP_425J2_127_3477_n1996,
         DP_OP_425J2_127_3477_n1995, DP_OP_425J2_127_3477_n1994,
         DP_OP_425J2_127_3477_n1993, DP_OP_425J2_127_3477_n1992,
         DP_OP_425J2_127_3477_n1991, DP_OP_425J2_127_3477_n1990,
         DP_OP_425J2_127_3477_n1989, DP_OP_425J2_127_3477_n1988,
         DP_OP_425J2_127_3477_n1987, DP_OP_425J2_127_3477_n1986,
         DP_OP_425J2_127_3477_n1985, DP_OP_425J2_127_3477_n1984,
         DP_OP_425J2_127_3477_n1983, DP_OP_425J2_127_3477_n1982,
         DP_OP_425J2_127_3477_n1981, DP_OP_425J2_127_3477_n1980,
         DP_OP_425J2_127_3477_n1979, DP_OP_425J2_127_3477_n1978,
         DP_OP_425J2_127_3477_n1977, DP_OP_425J2_127_3477_n1976,
         DP_OP_425J2_127_3477_n1975, DP_OP_425J2_127_3477_n1974,
         DP_OP_425J2_127_3477_n1973, DP_OP_425J2_127_3477_n1972,
         DP_OP_425J2_127_3477_n1971, DP_OP_425J2_127_3477_n1970,
         DP_OP_425J2_127_3477_n1968, DP_OP_425J2_127_3477_n1936,
         DP_OP_425J2_127_3477_n1935, DP_OP_425J2_127_3477_n1934,
         DP_OP_425J2_127_3477_n1932, DP_OP_425J2_127_3477_n1931,
         DP_OP_425J2_127_3477_n1930, DP_OP_425J2_127_3477_n1928,
         DP_OP_425J2_127_3477_n1927, DP_OP_425J2_127_3477_n1926,
         DP_OP_425J2_127_3477_n1925, DP_OP_425J2_127_3477_n1924,
         DP_OP_425J2_127_3477_n1923, DP_OP_425J2_127_3477_n1921,
         DP_OP_425J2_127_3477_n1920, DP_OP_425J2_127_3477_n1919,
         DP_OP_425J2_127_3477_n1918, DP_OP_425J2_127_3477_n1917,
         DP_OP_425J2_127_3477_n1916, DP_OP_425J2_127_3477_n1915,
         DP_OP_425J2_127_3477_n1914, DP_OP_425J2_127_3477_n1913,
         DP_OP_425J2_127_3477_n1912, DP_OP_425J2_127_3477_n1911,
         DP_OP_425J2_127_3477_n1910, DP_OP_425J2_127_3477_n1909,
         DP_OP_425J2_127_3477_n1908, DP_OP_425J2_127_3477_n1907,
         DP_OP_425J2_127_3477_n1906, DP_OP_425J2_127_3477_n1905,
         DP_OP_425J2_127_3477_n1904, DP_OP_425J2_127_3477_n1903,
         DP_OP_425J2_127_3477_n1902, DP_OP_425J2_127_3477_n1901,
         DP_OP_425J2_127_3477_n1900, DP_OP_425J2_127_3477_n1899,
         DP_OP_425J2_127_3477_n1898, DP_OP_425J2_127_3477_n1897,
         DP_OP_425J2_127_3477_n1896, DP_OP_425J2_127_3477_n1895,
         DP_OP_425J2_127_3477_n1894, DP_OP_425J2_127_3477_n1893,
         DP_OP_425J2_127_3477_n1892, DP_OP_425J2_127_3477_n1891,
         DP_OP_425J2_127_3477_n1890, DP_OP_425J2_127_3477_n1889,
         DP_OP_425J2_127_3477_n1888, DP_OP_425J2_127_3477_n1887,
         DP_OP_425J2_127_3477_n1886, DP_OP_425J2_127_3477_n1885,
         DP_OP_425J2_127_3477_n1884, DP_OP_425J2_127_3477_n1883,
         DP_OP_425J2_127_3477_n1882, DP_OP_425J2_127_3477_n1881,
         DP_OP_425J2_127_3477_n1880, DP_OP_425J2_127_3477_n1879,
         DP_OP_425J2_127_3477_n1878, DP_OP_425J2_127_3477_n1877,
         DP_OP_425J2_127_3477_n1876, DP_OP_425J2_127_3477_n1875,
         DP_OP_425J2_127_3477_n1874, DP_OP_425J2_127_3477_n1873,
         DP_OP_425J2_127_3477_n1872, DP_OP_425J2_127_3477_n1871,
         DP_OP_425J2_127_3477_n1870, DP_OP_425J2_127_3477_n1869,
         DP_OP_425J2_127_3477_n1868, DP_OP_425J2_127_3477_n1867,
         DP_OP_425J2_127_3477_n1866, DP_OP_425J2_127_3477_n1865,
         DP_OP_425J2_127_3477_n1864, DP_OP_425J2_127_3477_n1863,
         DP_OP_425J2_127_3477_n1862, DP_OP_425J2_127_3477_n1861,
         DP_OP_425J2_127_3477_n1860, DP_OP_425J2_127_3477_n1859,
         DP_OP_425J2_127_3477_n1858, DP_OP_425J2_127_3477_n1857,
         DP_OP_425J2_127_3477_n1856, DP_OP_425J2_127_3477_n1855,
         DP_OP_425J2_127_3477_n1854, DP_OP_425J2_127_3477_n1853,
         DP_OP_425J2_127_3477_n1852, DP_OP_425J2_127_3477_n1851,
         DP_OP_425J2_127_3477_n1850, DP_OP_425J2_127_3477_n1849,
         DP_OP_425J2_127_3477_n1848, DP_OP_425J2_127_3477_n1847,
         DP_OP_425J2_127_3477_n1846, DP_OP_425J2_127_3477_n1845,
         DP_OP_425J2_127_3477_n1844, DP_OP_425J2_127_3477_n1843,
         DP_OP_425J2_127_3477_n1842, DP_OP_425J2_127_3477_n1841,
         DP_OP_425J2_127_3477_n1840, DP_OP_425J2_127_3477_n1839,
         DP_OP_425J2_127_3477_n1838, DP_OP_425J2_127_3477_n1837,
         DP_OP_425J2_127_3477_n1836, DP_OP_425J2_127_3477_n1835,
         DP_OP_425J2_127_3477_n1834, DP_OP_425J2_127_3477_n1833,
         DP_OP_425J2_127_3477_n1832, DP_OP_425J2_127_3477_n1831,
         DP_OP_425J2_127_3477_n1830, DP_OP_425J2_127_3477_n1829,
         DP_OP_425J2_127_3477_n1828, DP_OP_425J2_127_3477_n1827,
         DP_OP_425J2_127_3477_n1826, DP_OP_425J2_127_3477_n1825,
         DP_OP_425J2_127_3477_n1824, DP_OP_425J2_127_3477_n1823,
         DP_OP_425J2_127_3477_n1822, DP_OP_425J2_127_3477_n1821,
         DP_OP_425J2_127_3477_n1820, DP_OP_425J2_127_3477_n1819,
         DP_OP_425J2_127_3477_n1818, DP_OP_425J2_127_3477_n1817,
         DP_OP_425J2_127_3477_n1816, DP_OP_425J2_127_3477_n1815,
         DP_OP_425J2_127_3477_n1814, DP_OP_425J2_127_3477_n1813,
         DP_OP_425J2_127_3477_n1812, DP_OP_425J2_127_3477_n1811,
         DP_OP_425J2_127_3477_n1810, DP_OP_425J2_127_3477_n1809,
         DP_OP_425J2_127_3477_n1808, DP_OP_425J2_127_3477_n1807,
         DP_OP_425J2_127_3477_n1806, DP_OP_425J2_127_3477_n1805,
         DP_OP_425J2_127_3477_n1804, DP_OP_425J2_127_3477_n1803,
         DP_OP_425J2_127_3477_n1802, DP_OP_425J2_127_3477_n1801,
         DP_OP_425J2_127_3477_n1800, DP_OP_425J2_127_3477_n1799,
         DP_OP_425J2_127_3477_n1798, DP_OP_425J2_127_3477_n1797,
         DP_OP_425J2_127_3477_n1796, DP_OP_425J2_127_3477_n1795,
         DP_OP_425J2_127_3477_n1794, DP_OP_425J2_127_3477_n1793,
         DP_OP_425J2_127_3477_n1792, DP_OP_425J2_127_3477_n1791,
         DP_OP_425J2_127_3477_n1790, DP_OP_425J2_127_3477_n1789,
         DP_OP_425J2_127_3477_n1788, DP_OP_425J2_127_3477_n1787,
         DP_OP_425J2_127_3477_n1786, DP_OP_425J2_127_3477_n1785,
         DP_OP_425J2_127_3477_n1784, DP_OP_425J2_127_3477_n1783,
         DP_OP_425J2_127_3477_n1782, DP_OP_425J2_127_3477_n1781,
         DP_OP_425J2_127_3477_n1780, DP_OP_425J2_127_3477_n1779,
         DP_OP_425J2_127_3477_n1778, DP_OP_425J2_127_3477_n1777,
         DP_OP_425J2_127_3477_n1776, DP_OP_425J2_127_3477_n1775,
         DP_OP_425J2_127_3477_n1774, DP_OP_425J2_127_3477_n1773,
         DP_OP_425J2_127_3477_n1772, DP_OP_425J2_127_3477_n1771,
         DP_OP_425J2_127_3477_n1770, DP_OP_425J2_127_3477_n1769,
         DP_OP_425J2_127_3477_n1768, DP_OP_425J2_127_3477_n1767,
         DP_OP_425J2_127_3477_n1766, DP_OP_425J2_127_3477_n1765,
         DP_OP_425J2_127_3477_n1764, DP_OP_425J2_127_3477_n1763,
         DP_OP_425J2_127_3477_n1762, DP_OP_425J2_127_3477_n1761,
         DP_OP_425J2_127_3477_n1760, DP_OP_425J2_127_3477_n1759,
         DP_OP_425J2_127_3477_n1758, DP_OP_425J2_127_3477_n1757,
         DP_OP_425J2_127_3477_n1756, DP_OP_425J2_127_3477_n1755,
         DP_OP_425J2_127_3477_n1754, DP_OP_425J2_127_3477_n1753,
         DP_OP_425J2_127_3477_n1752, DP_OP_425J2_127_3477_n1751,
         DP_OP_425J2_127_3477_n1750, DP_OP_425J2_127_3477_n1749,
         DP_OP_425J2_127_3477_n1748, DP_OP_425J2_127_3477_n1747,
         DP_OP_425J2_127_3477_n1746, DP_OP_425J2_127_3477_n1745,
         DP_OP_425J2_127_3477_n1744, DP_OP_425J2_127_3477_n1743,
         DP_OP_425J2_127_3477_n1742, DP_OP_425J2_127_3477_n1741,
         DP_OP_425J2_127_3477_n1740, DP_OP_425J2_127_3477_n1739,
         DP_OP_425J2_127_3477_n1738, DP_OP_425J2_127_3477_n1737,
         DP_OP_425J2_127_3477_n1736, DP_OP_425J2_127_3477_n1735,
         DP_OP_425J2_127_3477_n1734, DP_OP_425J2_127_3477_n1733,
         DP_OP_425J2_127_3477_n1732, DP_OP_425J2_127_3477_n1731,
         DP_OP_425J2_127_3477_n1730, DP_OP_425J2_127_3477_n1729,
         DP_OP_425J2_127_3477_n1728, DP_OP_425J2_127_3477_n1727,
         DP_OP_425J2_127_3477_n1726, DP_OP_425J2_127_3477_n1725,
         DP_OP_425J2_127_3477_n1724, DP_OP_425J2_127_3477_n1723,
         DP_OP_425J2_127_3477_n1722, DP_OP_425J2_127_3477_n1721,
         DP_OP_425J2_127_3477_n1720, DP_OP_425J2_127_3477_n1719,
         DP_OP_425J2_127_3477_n1718, DP_OP_425J2_127_3477_n1717,
         DP_OP_425J2_127_3477_n1716, DP_OP_425J2_127_3477_n1715,
         DP_OP_425J2_127_3477_n1714, DP_OP_425J2_127_3477_n1713,
         DP_OP_425J2_127_3477_n1712, DP_OP_425J2_127_3477_n1711,
         DP_OP_425J2_127_3477_n1710, DP_OP_425J2_127_3477_n1709,
         DP_OP_425J2_127_3477_n1708, DP_OP_425J2_127_3477_n1707,
         DP_OP_425J2_127_3477_n1706, DP_OP_425J2_127_3477_n1705,
         DP_OP_425J2_127_3477_n1704, DP_OP_425J2_127_3477_n1703,
         DP_OP_425J2_127_3477_n1702, DP_OP_425J2_127_3477_n1701,
         DP_OP_425J2_127_3477_n1700, DP_OP_425J2_127_3477_n1699,
         DP_OP_425J2_127_3477_n1698, DP_OP_425J2_127_3477_n1697,
         DP_OP_425J2_127_3477_n1696, DP_OP_425J2_127_3477_n1695,
         DP_OP_425J2_127_3477_n1694, DP_OP_425J2_127_3477_n1693,
         DP_OP_425J2_127_3477_n1692, DP_OP_425J2_127_3477_n1691,
         DP_OP_425J2_127_3477_n1690, DP_OP_425J2_127_3477_n1689,
         DP_OP_425J2_127_3477_n1688, DP_OP_425J2_127_3477_n1687,
         DP_OP_425J2_127_3477_n1686, DP_OP_425J2_127_3477_n1685,
         DP_OP_425J2_127_3477_n1684, DP_OP_425J2_127_3477_n1683,
         DP_OP_425J2_127_3477_n1682, DP_OP_425J2_127_3477_n1681,
         DP_OP_425J2_127_3477_n1680, DP_OP_425J2_127_3477_n1679,
         DP_OP_425J2_127_3477_n1678, DP_OP_425J2_127_3477_n1676,
         DP_OP_425J2_127_3477_n1675, DP_OP_425J2_127_3477_n1674,
         DP_OP_425J2_127_3477_n1673, DP_OP_425J2_127_3477_n1672,
         DP_OP_425J2_127_3477_n1671, DP_OP_425J2_127_3477_n1670,
         DP_OP_425J2_127_3477_n1669, DP_OP_425J2_127_3477_n1668,
         DP_OP_425J2_127_3477_n1667, DP_OP_425J2_127_3477_n1666,
         DP_OP_425J2_127_3477_n1665, DP_OP_425J2_127_3477_n1664,
         DP_OP_425J2_127_3477_n1663, DP_OP_425J2_127_3477_n1662,
         DP_OP_425J2_127_3477_n1661, DP_OP_425J2_127_3477_n1660,
         DP_OP_425J2_127_3477_n1659, DP_OP_425J2_127_3477_n1658,
         DP_OP_425J2_127_3477_n1657, DP_OP_425J2_127_3477_n1656,
         DP_OP_425J2_127_3477_n1655, DP_OP_425J2_127_3477_n1654,
         DP_OP_425J2_127_3477_n1653, DP_OP_425J2_127_3477_n1652,
         DP_OP_425J2_127_3477_n1651, DP_OP_425J2_127_3477_n1650,
         DP_OP_425J2_127_3477_n1649, DP_OP_425J2_127_3477_n1648,
         DP_OP_425J2_127_3477_n1647, DP_OP_425J2_127_3477_n1646,
         DP_OP_425J2_127_3477_n1645, DP_OP_425J2_127_3477_n1644,
         DP_OP_425J2_127_3477_n1643, DP_OP_425J2_127_3477_n1642,
         DP_OP_425J2_127_3477_n1641, DP_OP_425J2_127_3477_n1640,
         DP_OP_425J2_127_3477_n1639, DP_OP_425J2_127_3477_n1638,
         DP_OP_425J2_127_3477_n1637, DP_OP_425J2_127_3477_n1636,
         DP_OP_425J2_127_3477_n1635, DP_OP_425J2_127_3477_n1634,
         DP_OP_425J2_127_3477_n1633, DP_OP_425J2_127_3477_n1632,
         DP_OP_425J2_127_3477_n1631, DP_OP_425J2_127_3477_n1630,
         DP_OP_425J2_127_3477_n1629, DP_OP_425J2_127_3477_n1628,
         DP_OP_425J2_127_3477_n1627, DP_OP_425J2_127_3477_n1626,
         DP_OP_425J2_127_3477_n1625, DP_OP_425J2_127_3477_n1624,
         DP_OP_425J2_127_3477_n1623, DP_OP_425J2_127_3477_n1622,
         DP_OP_425J2_127_3477_n1621, DP_OP_425J2_127_3477_n1620,
         DP_OP_425J2_127_3477_n1619, DP_OP_425J2_127_3477_n1618,
         DP_OP_425J2_127_3477_n1617, DP_OP_425J2_127_3477_n1616,
         DP_OP_425J2_127_3477_n1615, DP_OP_425J2_127_3477_n1614,
         DP_OP_425J2_127_3477_n1613, DP_OP_425J2_127_3477_n1612,
         DP_OP_425J2_127_3477_n1611, DP_OP_425J2_127_3477_n1610,
         DP_OP_425J2_127_3477_n1609, DP_OP_425J2_127_3477_n1608,
         DP_OP_425J2_127_3477_n1607, DP_OP_425J2_127_3477_n1606,
         DP_OP_425J2_127_3477_n1605, DP_OP_425J2_127_3477_n1604,
         DP_OP_425J2_127_3477_n1603, DP_OP_425J2_127_3477_n1602,
         DP_OP_425J2_127_3477_n1601, DP_OP_425J2_127_3477_n1600,
         DP_OP_425J2_127_3477_n1599, DP_OP_425J2_127_3477_n1598,
         DP_OP_425J2_127_3477_n1597, DP_OP_425J2_127_3477_n1596,
         DP_OP_425J2_127_3477_n1595, DP_OP_425J2_127_3477_n1594,
         DP_OP_425J2_127_3477_n1593, DP_OP_425J2_127_3477_n1592,
         DP_OP_425J2_127_3477_n1591, DP_OP_425J2_127_3477_n1590,
         DP_OP_425J2_127_3477_n1589, DP_OP_425J2_127_3477_n1588,
         DP_OP_425J2_127_3477_n1587, DP_OP_425J2_127_3477_n1586,
         DP_OP_425J2_127_3477_n1585, DP_OP_425J2_127_3477_n1584,
         DP_OP_425J2_127_3477_n1583, DP_OP_425J2_127_3477_n1582,
         DP_OP_425J2_127_3477_n1581, DP_OP_425J2_127_3477_n1580,
         DP_OP_425J2_127_3477_n1579, DP_OP_425J2_127_3477_n1578,
         DP_OP_425J2_127_3477_n1577, DP_OP_425J2_127_3477_n1576,
         DP_OP_425J2_127_3477_n1575, DP_OP_425J2_127_3477_n1574,
         DP_OP_425J2_127_3477_n1573, DP_OP_425J2_127_3477_n1572,
         DP_OP_425J2_127_3477_n1571, DP_OP_425J2_127_3477_n1570,
         DP_OP_425J2_127_3477_n1569, DP_OP_425J2_127_3477_n1568,
         DP_OP_425J2_127_3477_n1567, DP_OP_425J2_127_3477_n1566,
         DP_OP_425J2_127_3477_n1565, DP_OP_425J2_127_3477_n1564,
         DP_OP_425J2_127_3477_n1563, DP_OP_425J2_127_3477_n1562,
         DP_OP_425J2_127_3477_n1561, DP_OP_425J2_127_3477_n1560,
         DP_OP_425J2_127_3477_n1559, DP_OP_425J2_127_3477_n1558,
         DP_OP_425J2_127_3477_n1557, DP_OP_425J2_127_3477_n1556,
         DP_OP_425J2_127_3477_n1555, DP_OP_425J2_127_3477_n1554,
         DP_OP_425J2_127_3477_n1553, DP_OP_425J2_127_3477_n1552,
         DP_OP_425J2_127_3477_n1551, DP_OP_425J2_127_3477_n1550,
         DP_OP_425J2_127_3477_n1549, DP_OP_425J2_127_3477_n1548,
         DP_OP_425J2_127_3477_n1547, DP_OP_425J2_127_3477_n1546,
         DP_OP_425J2_127_3477_n1545, DP_OP_425J2_127_3477_n1544,
         DP_OP_425J2_127_3477_n1543, DP_OP_425J2_127_3477_n1542,
         DP_OP_425J2_127_3477_n1541, DP_OP_425J2_127_3477_n1540,
         DP_OP_425J2_127_3477_n1539, DP_OP_425J2_127_3477_n1538,
         DP_OP_425J2_127_3477_n1537, DP_OP_425J2_127_3477_n1536,
         DP_OP_425J2_127_3477_n1535, DP_OP_425J2_127_3477_n1534,
         DP_OP_425J2_127_3477_n1533, DP_OP_425J2_127_3477_n1532,
         DP_OP_425J2_127_3477_n1531, DP_OP_425J2_127_3477_n1530,
         DP_OP_425J2_127_3477_n1529, DP_OP_425J2_127_3477_n1528,
         DP_OP_425J2_127_3477_n1527, DP_OP_425J2_127_3477_n1526,
         DP_OP_425J2_127_3477_n1525, DP_OP_425J2_127_3477_n1524,
         DP_OP_425J2_127_3477_n1523, DP_OP_425J2_127_3477_n1522,
         DP_OP_425J2_127_3477_n1521, DP_OP_425J2_127_3477_n1520,
         DP_OP_425J2_127_3477_n1519, DP_OP_425J2_127_3477_n1518,
         DP_OP_425J2_127_3477_n1517, DP_OP_425J2_127_3477_n1516,
         DP_OP_425J2_127_3477_n1515, DP_OP_425J2_127_3477_n1514,
         DP_OP_425J2_127_3477_n1513, DP_OP_425J2_127_3477_n1512,
         DP_OP_425J2_127_3477_n1511, DP_OP_425J2_127_3477_n1510,
         DP_OP_425J2_127_3477_n1509, DP_OP_425J2_127_3477_n1508,
         DP_OP_425J2_127_3477_n1507, DP_OP_425J2_127_3477_n1506,
         DP_OP_425J2_127_3477_n1505, DP_OP_425J2_127_3477_n1504,
         DP_OP_425J2_127_3477_n1503, DP_OP_425J2_127_3477_n1502,
         DP_OP_425J2_127_3477_n1501, DP_OP_425J2_127_3477_n1500,
         DP_OP_425J2_127_3477_n1499, DP_OP_425J2_127_3477_n1498,
         DP_OP_425J2_127_3477_n1497, DP_OP_425J2_127_3477_n1496,
         DP_OP_425J2_127_3477_n1495, DP_OP_425J2_127_3477_n1494,
         DP_OP_425J2_127_3477_n1493, DP_OP_425J2_127_3477_n1492,
         DP_OP_425J2_127_3477_n1491, DP_OP_425J2_127_3477_n1490,
         DP_OP_425J2_127_3477_n1489, DP_OP_425J2_127_3477_n1488,
         DP_OP_425J2_127_3477_n1487, DP_OP_425J2_127_3477_n1486,
         DP_OP_425J2_127_3477_n1485, DP_OP_425J2_127_3477_n1484,
         DP_OP_425J2_127_3477_n1483, DP_OP_425J2_127_3477_n1482,
         DP_OP_425J2_127_3477_n1481, DP_OP_425J2_127_3477_n1480,
         DP_OP_425J2_127_3477_n1479, DP_OP_425J2_127_3477_n1478,
         DP_OP_425J2_127_3477_n1477, DP_OP_425J2_127_3477_n1476,
         DP_OP_425J2_127_3477_n1475, DP_OP_425J2_127_3477_n1474,
         DP_OP_425J2_127_3477_n1473, DP_OP_425J2_127_3477_n1472,
         DP_OP_425J2_127_3477_n1471, DP_OP_425J2_127_3477_n1470,
         DP_OP_425J2_127_3477_n1469, DP_OP_425J2_127_3477_n1468,
         DP_OP_425J2_127_3477_n1467, DP_OP_425J2_127_3477_n1466,
         DP_OP_425J2_127_3477_n1465, DP_OP_425J2_127_3477_n1464,
         DP_OP_425J2_127_3477_n1463, DP_OP_425J2_127_3477_n1462,
         DP_OP_425J2_127_3477_n1461, DP_OP_425J2_127_3477_n1460,
         DP_OP_425J2_127_3477_n1459, DP_OP_425J2_127_3477_n1458,
         DP_OP_425J2_127_3477_n1457, DP_OP_425J2_127_3477_n1456,
         DP_OP_425J2_127_3477_n1455, DP_OP_425J2_127_3477_n1454,
         DP_OP_425J2_127_3477_n1453, DP_OP_425J2_127_3477_n1452,
         DP_OP_425J2_127_3477_n1451, DP_OP_425J2_127_3477_n1450,
         DP_OP_425J2_127_3477_n1449, DP_OP_425J2_127_3477_n1448,
         DP_OP_425J2_127_3477_n1447, DP_OP_425J2_127_3477_n1446,
         DP_OP_425J2_127_3477_n1445, DP_OP_425J2_127_3477_n1444,
         DP_OP_425J2_127_3477_n1443, DP_OP_425J2_127_3477_n1442,
         DP_OP_425J2_127_3477_n1441, DP_OP_425J2_127_3477_n1440,
         DP_OP_425J2_127_3477_n1439, DP_OP_425J2_127_3477_n1438,
         DP_OP_425J2_127_3477_n1437, DP_OP_425J2_127_3477_n1436,
         DP_OP_425J2_127_3477_n1435, DP_OP_425J2_127_3477_n1434,
         DP_OP_425J2_127_3477_n1433, DP_OP_425J2_127_3477_n1432,
         DP_OP_425J2_127_3477_n1431, DP_OP_425J2_127_3477_n1430,
         DP_OP_425J2_127_3477_n1429, DP_OP_425J2_127_3477_n1428,
         DP_OP_425J2_127_3477_n1427, DP_OP_425J2_127_3477_n1426,
         DP_OP_425J2_127_3477_n1425, DP_OP_425J2_127_3477_n1424,
         DP_OP_425J2_127_3477_n1423, DP_OP_425J2_127_3477_n1422,
         DP_OP_425J2_127_3477_n1421, DP_OP_425J2_127_3477_n1420,
         DP_OP_425J2_127_3477_n1419, DP_OP_425J2_127_3477_n1418,
         DP_OP_425J2_127_3477_n1417, DP_OP_425J2_127_3477_n1416,
         DP_OP_425J2_127_3477_n1415, DP_OP_425J2_127_3477_n1414,
         DP_OP_425J2_127_3477_n1413, DP_OP_425J2_127_3477_n1412,
         DP_OP_425J2_127_3477_n1411, DP_OP_425J2_127_3477_n1410,
         DP_OP_425J2_127_3477_n1409, DP_OP_425J2_127_3477_n1408,
         DP_OP_425J2_127_3477_n1407, DP_OP_425J2_127_3477_n1406,
         DP_OP_425J2_127_3477_n1405, DP_OP_425J2_127_3477_n1404,
         DP_OP_425J2_127_3477_n1403, DP_OP_425J2_127_3477_n1402,
         DP_OP_425J2_127_3477_n1401, DP_OP_425J2_127_3477_n1400,
         DP_OP_425J2_127_3477_n1399, DP_OP_425J2_127_3477_n1398,
         DP_OP_425J2_127_3477_n1397, DP_OP_425J2_127_3477_n1396,
         DP_OP_425J2_127_3477_n1395, DP_OP_425J2_127_3477_n1394,
         DP_OP_425J2_127_3477_n1393, DP_OP_425J2_127_3477_n1392,
         DP_OP_425J2_127_3477_n1391, DP_OP_425J2_127_3477_n1390,
         DP_OP_425J2_127_3477_n1389, DP_OP_425J2_127_3477_n1388,
         DP_OP_425J2_127_3477_n1387, DP_OP_425J2_127_3477_n1386,
         DP_OP_425J2_127_3477_n1385, DP_OP_425J2_127_3477_n1384,
         DP_OP_425J2_127_3477_n1383, DP_OP_425J2_127_3477_n1382,
         DP_OP_425J2_127_3477_n1381, DP_OP_425J2_127_3477_n1380,
         DP_OP_425J2_127_3477_n1379, DP_OP_425J2_127_3477_n1378,
         DP_OP_425J2_127_3477_n1377, DP_OP_425J2_127_3477_n1376,
         DP_OP_425J2_127_3477_n1375, DP_OP_425J2_127_3477_n1374,
         DP_OP_425J2_127_3477_n1373, DP_OP_425J2_127_3477_n1372,
         DP_OP_425J2_127_3477_n1371, DP_OP_425J2_127_3477_n1370,
         DP_OP_425J2_127_3477_n1369, DP_OP_425J2_127_3477_n1368,
         DP_OP_425J2_127_3477_n1367, DP_OP_425J2_127_3477_n1366,
         DP_OP_425J2_127_3477_n1365, DP_OP_425J2_127_3477_n1364,
         DP_OP_425J2_127_3477_n1363, DP_OP_425J2_127_3477_n1362,
         DP_OP_425J2_127_3477_n1361, DP_OP_425J2_127_3477_n1360,
         DP_OP_425J2_127_3477_n1359, DP_OP_425J2_127_3477_n1358,
         DP_OP_425J2_127_3477_n1357, DP_OP_425J2_127_3477_n1356,
         DP_OP_425J2_127_3477_n1355, DP_OP_425J2_127_3477_n1354,
         DP_OP_425J2_127_3477_n1353, DP_OP_425J2_127_3477_n1352,
         DP_OP_425J2_127_3477_n1351, DP_OP_425J2_127_3477_n1350,
         DP_OP_425J2_127_3477_n1349, DP_OP_425J2_127_3477_n1348,
         DP_OP_425J2_127_3477_n1347, DP_OP_425J2_127_3477_n1346,
         DP_OP_425J2_127_3477_n1345, DP_OP_425J2_127_3477_n1344,
         DP_OP_425J2_127_3477_n1343, DP_OP_425J2_127_3477_n1342,
         DP_OP_425J2_127_3477_n1341, DP_OP_425J2_127_3477_n1340,
         DP_OP_425J2_127_3477_n1339, DP_OP_425J2_127_3477_n1338,
         DP_OP_425J2_127_3477_n1337, DP_OP_425J2_127_3477_n1336,
         DP_OP_425J2_127_3477_n1335, DP_OP_425J2_127_3477_n1334,
         DP_OP_425J2_127_3477_n1333, DP_OP_425J2_127_3477_n1332,
         DP_OP_425J2_127_3477_n1331, DP_OP_425J2_127_3477_n1330,
         DP_OP_425J2_127_3477_n1329, DP_OP_425J2_127_3477_n1328,
         DP_OP_425J2_127_3477_n1327, DP_OP_425J2_127_3477_n1326,
         DP_OP_425J2_127_3477_n1325, DP_OP_425J2_127_3477_n1324,
         DP_OP_425J2_127_3477_n1323, DP_OP_425J2_127_3477_n1322,
         DP_OP_425J2_127_3477_n1321, DP_OP_425J2_127_3477_n1320,
         DP_OP_425J2_127_3477_n1319, DP_OP_425J2_127_3477_n1318,
         DP_OP_425J2_127_3477_n1317, DP_OP_425J2_127_3477_n1316,
         DP_OP_425J2_127_3477_n1315, DP_OP_425J2_127_3477_n1314,
         DP_OP_425J2_127_3477_n1313, DP_OP_425J2_127_3477_n1312,
         DP_OP_425J2_127_3477_n1311, DP_OP_425J2_127_3477_n1310,
         DP_OP_425J2_127_3477_n1309, DP_OP_425J2_127_3477_n1308,
         DP_OP_425J2_127_3477_n1307, DP_OP_425J2_127_3477_n1306,
         DP_OP_425J2_127_3477_n1305, DP_OP_425J2_127_3477_n1304,
         DP_OP_425J2_127_3477_n1303, DP_OP_425J2_127_3477_n1302,
         DP_OP_425J2_127_3477_n1301, DP_OP_425J2_127_3477_n1300,
         DP_OP_425J2_127_3477_n1299, DP_OP_425J2_127_3477_n1298,
         DP_OP_425J2_127_3477_n1297, DP_OP_425J2_127_3477_n1296,
         DP_OP_425J2_127_3477_n1295, DP_OP_425J2_127_3477_n1294,
         DP_OP_425J2_127_3477_n1293, DP_OP_425J2_127_3477_n1292,
         DP_OP_425J2_127_3477_n1291, DP_OP_425J2_127_3477_n1290,
         DP_OP_425J2_127_3477_n1289, DP_OP_425J2_127_3477_n1288,
         DP_OP_425J2_127_3477_n1287, DP_OP_425J2_127_3477_n1286,
         DP_OP_425J2_127_3477_n1285, DP_OP_425J2_127_3477_n1284,
         DP_OP_425J2_127_3477_n1283, DP_OP_425J2_127_3477_n1282,
         DP_OP_425J2_127_3477_n1281, DP_OP_425J2_127_3477_n1280,
         DP_OP_425J2_127_3477_n1279, DP_OP_425J2_127_3477_n1278,
         DP_OP_425J2_127_3477_n1277, DP_OP_425J2_127_3477_n1276,
         DP_OP_425J2_127_3477_n1275, DP_OP_425J2_127_3477_n1274,
         DP_OP_425J2_127_3477_n1273, DP_OP_425J2_127_3477_n1272,
         DP_OP_425J2_127_3477_n1271, DP_OP_425J2_127_3477_n1270,
         DP_OP_425J2_127_3477_n1269, DP_OP_425J2_127_3477_n1268,
         DP_OP_425J2_127_3477_n1267, DP_OP_425J2_127_3477_n1266,
         DP_OP_425J2_127_3477_n1265, DP_OP_425J2_127_3477_n1264,
         DP_OP_425J2_127_3477_n1263, DP_OP_425J2_127_3477_n1262,
         DP_OP_425J2_127_3477_n1261, DP_OP_425J2_127_3477_n1260,
         DP_OP_425J2_127_3477_n1259, DP_OP_425J2_127_3477_n1258,
         DP_OP_425J2_127_3477_n1257, DP_OP_425J2_127_3477_n1256,
         DP_OP_425J2_127_3477_n1255, DP_OP_425J2_127_3477_n1254,
         DP_OP_425J2_127_3477_n1253, DP_OP_425J2_127_3477_n1252,
         DP_OP_425J2_127_3477_n1251, DP_OP_425J2_127_3477_n1250,
         DP_OP_425J2_127_3477_n1249, DP_OP_425J2_127_3477_n1248,
         DP_OP_425J2_127_3477_n1247, DP_OP_425J2_127_3477_n1246,
         DP_OP_425J2_127_3477_n1245, DP_OP_425J2_127_3477_n1244,
         DP_OP_425J2_127_3477_n1243, DP_OP_425J2_127_3477_n1242,
         DP_OP_425J2_127_3477_n1241, DP_OP_425J2_127_3477_n1240,
         DP_OP_425J2_127_3477_n1239, DP_OP_425J2_127_3477_n1238,
         DP_OP_425J2_127_3477_n1237, DP_OP_425J2_127_3477_n1236,
         DP_OP_425J2_127_3477_n1235, DP_OP_425J2_127_3477_n1234,
         DP_OP_425J2_127_3477_n1233, DP_OP_425J2_127_3477_n1232,
         DP_OP_425J2_127_3477_n1231, DP_OP_425J2_127_3477_n1230,
         DP_OP_425J2_127_3477_n1229, DP_OP_425J2_127_3477_n1228,
         DP_OP_425J2_127_3477_n1227, DP_OP_425J2_127_3477_n1226,
         DP_OP_425J2_127_3477_n1225, DP_OP_425J2_127_3477_n1224,
         DP_OP_425J2_127_3477_n1223, DP_OP_425J2_127_3477_n1222,
         DP_OP_425J2_127_3477_n1221, DP_OP_425J2_127_3477_n1220,
         DP_OP_425J2_127_3477_n1219, DP_OP_425J2_127_3477_n1218,
         DP_OP_425J2_127_3477_n1217, DP_OP_425J2_127_3477_n1216,
         DP_OP_425J2_127_3477_n1215, DP_OP_425J2_127_3477_n1214,
         DP_OP_425J2_127_3477_n1213, DP_OP_425J2_127_3477_n1212,
         DP_OP_425J2_127_3477_n1211, DP_OP_425J2_127_3477_n1210,
         DP_OP_425J2_127_3477_n1209, DP_OP_425J2_127_3477_n1208,
         DP_OP_425J2_127_3477_n1207, DP_OP_425J2_127_3477_n1206,
         DP_OP_425J2_127_3477_n1205, DP_OP_425J2_127_3477_n1204,
         DP_OP_425J2_127_3477_n1203, DP_OP_425J2_127_3477_n1202,
         DP_OP_425J2_127_3477_n1201, DP_OP_425J2_127_3477_n1200,
         DP_OP_425J2_127_3477_n1199, DP_OP_425J2_127_3477_n1198,
         DP_OP_425J2_127_3477_n1197, DP_OP_425J2_127_3477_n1196,
         DP_OP_425J2_127_3477_n1195, DP_OP_425J2_127_3477_n1194,
         DP_OP_425J2_127_3477_n1193, DP_OP_425J2_127_3477_n1192,
         DP_OP_425J2_127_3477_n1191, DP_OP_425J2_127_3477_n1190,
         DP_OP_425J2_127_3477_n1189, DP_OP_425J2_127_3477_n1188,
         DP_OP_425J2_127_3477_n1187, DP_OP_425J2_127_3477_n1186,
         DP_OP_425J2_127_3477_n1185, DP_OP_425J2_127_3477_n1184,
         DP_OP_425J2_127_3477_n1183, DP_OP_425J2_127_3477_n1182,
         DP_OP_425J2_127_3477_n1181, DP_OP_425J2_127_3477_n1180,
         DP_OP_425J2_127_3477_n1179, DP_OP_425J2_127_3477_n1178,
         DP_OP_425J2_127_3477_n1177, DP_OP_425J2_127_3477_n1176,
         DP_OP_425J2_127_3477_n1175, DP_OP_425J2_127_3477_n1174,
         DP_OP_425J2_127_3477_n1173, DP_OP_425J2_127_3477_n1172,
         DP_OP_425J2_127_3477_n1171, DP_OP_425J2_127_3477_n1170,
         DP_OP_425J2_127_3477_n1169, DP_OP_425J2_127_3477_n1168,
         DP_OP_425J2_127_3477_n1167, DP_OP_425J2_127_3477_n1166,
         DP_OP_425J2_127_3477_n1165, DP_OP_425J2_127_3477_n1164,
         DP_OP_425J2_127_3477_n1163, DP_OP_425J2_127_3477_n1162,
         DP_OP_425J2_127_3477_n1161, DP_OP_425J2_127_3477_n1160,
         DP_OP_425J2_127_3477_n1159, DP_OP_425J2_127_3477_n1158,
         DP_OP_425J2_127_3477_n1157, DP_OP_425J2_127_3477_n1156,
         DP_OP_425J2_127_3477_n1155, DP_OP_425J2_127_3477_n1154,
         DP_OP_425J2_127_3477_n1153, DP_OP_425J2_127_3477_n1152,
         DP_OP_425J2_127_3477_n1151, DP_OP_425J2_127_3477_n1150,
         DP_OP_425J2_127_3477_n1149, DP_OP_425J2_127_3477_n1148,
         DP_OP_425J2_127_3477_n1147, DP_OP_425J2_127_3477_n1146,
         DP_OP_425J2_127_3477_n1145, DP_OP_425J2_127_3477_n1144,
         DP_OP_425J2_127_3477_n1143, DP_OP_425J2_127_3477_n1142,
         DP_OP_425J2_127_3477_n1141, DP_OP_425J2_127_3477_n1140,
         DP_OP_425J2_127_3477_n1139, DP_OP_425J2_127_3477_n1138,
         DP_OP_425J2_127_3477_n1137, DP_OP_425J2_127_3477_n1136,
         DP_OP_425J2_127_3477_n1135, DP_OP_425J2_127_3477_n1134,
         DP_OP_425J2_127_3477_n1133, DP_OP_425J2_127_3477_n1132,
         DP_OP_425J2_127_3477_n1131, DP_OP_425J2_127_3477_n1130,
         DP_OP_425J2_127_3477_n1129, DP_OP_425J2_127_3477_n1128,
         DP_OP_425J2_127_3477_n1127, DP_OP_425J2_127_3477_n1126,
         DP_OP_425J2_127_3477_n1125, DP_OP_425J2_127_3477_n1124,
         DP_OP_425J2_127_3477_n1123, DP_OP_425J2_127_3477_n1122,
         DP_OP_425J2_127_3477_n1121, DP_OP_425J2_127_3477_n1120,
         DP_OP_425J2_127_3477_n1119, DP_OP_425J2_127_3477_n1118,
         DP_OP_425J2_127_3477_n1117, DP_OP_425J2_127_3477_n1116,
         DP_OP_425J2_127_3477_n1115, DP_OP_425J2_127_3477_n1114,
         DP_OP_425J2_127_3477_n1113, DP_OP_425J2_127_3477_n1112,
         DP_OP_425J2_127_3477_n1111, DP_OP_425J2_127_3477_n1110,
         DP_OP_425J2_127_3477_n1109, DP_OP_425J2_127_3477_n1108,
         DP_OP_425J2_127_3477_n1107, DP_OP_425J2_127_3477_n1106,
         DP_OP_425J2_127_3477_n1105, DP_OP_425J2_127_3477_n1104,
         DP_OP_425J2_127_3477_n1103, DP_OP_425J2_127_3477_n1102,
         DP_OP_425J2_127_3477_n1101, DP_OP_425J2_127_3477_n1100,
         DP_OP_425J2_127_3477_n1099, DP_OP_425J2_127_3477_n1098,
         DP_OP_425J2_127_3477_n1097, DP_OP_425J2_127_3477_n1096,
         DP_OP_425J2_127_3477_n1095, DP_OP_425J2_127_3477_n1094,
         DP_OP_425J2_127_3477_n1093, DP_OP_425J2_127_3477_n1092,
         DP_OP_425J2_127_3477_n1091, DP_OP_425J2_127_3477_n1090,
         DP_OP_425J2_127_3477_n1089, DP_OP_425J2_127_3477_n1088,
         DP_OP_425J2_127_3477_n1087, DP_OP_425J2_127_3477_n1086,
         DP_OP_425J2_127_3477_n1085, DP_OP_425J2_127_3477_n1084,
         DP_OP_425J2_127_3477_n1083, DP_OP_425J2_127_3477_n1082,
         DP_OP_425J2_127_3477_n1081, DP_OP_425J2_127_3477_n1080,
         DP_OP_425J2_127_3477_n1079, DP_OP_425J2_127_3477_n1078,
         DP_OP_425J2_127_3477_n1077, DP_OP_425J2_127_3477_n1076,
         DP_OP_425J2_127_3477_n1075, DP_OP_425J2_127_3477_n1074,
         DP_OP_425J2_127_3477_n1073, DP_OP_425J2_127_3477_n1072,
         DP_OP_425J2_127_3477_n1071, DP_OP_425J2_127_3477_n1070,
         DP_OP_425J2_127_3477_n1069, DP_OP_425J2_127_3477_n1068,
         DP_OP_425J2_127_3477_n1067, DP_OP_425J2_127_3477_n1066,
         DP_OP_425J2_127_3477_n1065, DP_OP_425J2_127_3477_n1064,
         DP_OP_425J2_127_3477_n1063, DP_OP_425J2_127_3477_n1062,
         DP_OP_425J2_127_3477_n1061, DP_OP_425J2_127_3477_n1060,
         DP_OP_425J2_127_3477_n1059, DP_OP_425J2_127_3477_n1058,
         DP_OP_425J2_127_3477_n1057, DP_OP_425J2_127_3477_n1056,
         DP_OP_425J2_127_3477_n1055, DP_OP_425J2_127_3477_n1054,
         DP_OP_425J2_127_3477_n1053, DP_OP_425J2_127_3477_n1052,
         DP_OP_425J2_127_3477_n1051, DP_OP_425J2_127_3477_n1050,
         DP_OP_425J2_127_3477_n1049, DP_OP_425J2_127_3477_n1048,
         DP_OP_425J2_127_3477_n1047, DP_OP_425J2_127_3477_n1046,
         DP_OP_425J2_127_3477_n1045, DP_OP_425J2_127_3477_n1044,
         DP_OP_425J2_127_3477_n1043, DP_OP_425J2_127_3477_n1042,
         DP_OP_425J2_127_3477_n1041, DP_OP_425J2_127_3477_n1040,
         DP_OP_425J2_127_3477_n1039, DP_OP_425J2_127_3477_n1038,
         DP_OP_425J2_127_3477_n1037, DP_OP_425J2_127_3477_n1036,
         DP_OP_425J2_127_3477_n1035, DP_OP_425J2_127_3477_n1034,
         DP_OP_425J2_127_3477_n1033, DP_OP_425J2_127_3477_n1032,
         DP_OP_425J2_127_3477_n1031, DP_OP_425J2_127_3477_n1030,
         DP_OP_425J2_127_3477_n1029, DP_OP_425J2_127_3477_n1028,
         DP_OP_425J2_127_3477_n1027, DP_OP_425J2_127_3477_n1026,
         DP_OP_425J2_127_3477_n1025, DP_OP_425J2_127_3477_n1024,
         DP_OP_425J2_127_3477_n1023, DP_OP_425J2_127_3477_n1022,
         DP_OP_425J2_127_3477_n1021, DP_OP_425J2_127_3477_n1020,
         DP_OP_425J2_127_3477_n1019, DP_OP_425J2_127_3477_n1018,
         DP_OP_425J2_127_3477_n1017, DP_OP_425J2_127_3477_n1016,
         DP_OP_425J2_127_3477_n1015, DP_OP_425J2_127_3477_n1014,
         DP_OP_425J2_127_3477_n1013, DP_OP_425J2_127_3477_n1012,
         DP_OP_425J2_127_3477_n1011, DP_OP_425J2_127_3477_n1010,
         DP_OP_425J2_127_3477_n1009, DP_OP_425J2_127_3477_n1008,
         DP_OP_425J2_127_3477_n1007, DP_OP_425J2_127_3477_n1006,
         DP_OP_425J2_127_3477_n1005, DP_OP_425J2_127_3477_n1004,
         DP_OP_425J2_127_3477_n1003, DP_OP_425J2_127_3477_n1002,
         DP_OP_425J2_127_3477_n1001, DP_OP_425J2_127_3477_n1000,
         DP_OP_425J2_127_3477_n999, DP_OP_425J2_127_3477_n998,
         DP_OP_425J2_127_3477_n997, DP_OP_425J2_127_3477_n996,
         DP_OP_425J2_127_3477_n995, DP_OP_425J2_127_3477_n994,
         DP_OP_425J2_127_3477_n993, DP_OP_425J2_127_3477_n992,
         DP_OP_425J2_127_3477_n991, DP_OP_425J2_127_3477_n990,
         DP_OP_425J2_127_3477_n989, DP_OP_425J2_127_3477_n988,
         DP_OP_425J2_127_3477_n987, DP_OP_425J2_127_3477_n986,
         DP_OP_425J2_127_3477_n985, DP_OP_425J2_127_3477_n984,
         DP_OP_425J2_127_3477_n983, DP_OP_425J2_127_3477_n982,
         DP_OP_425J2_127_3477_n981, DP_OP_425J2_127_3477_n980,
         DP_OP_425J2_127_3477_n979, DP_OP_425J2_127_3477_n978,
         DP_OP_425J2_127_3477_n977, DP_OP_425J2_127_3477_n976,
         DP_OP_425J2_127_3477_n975, DP_OP_425J2_127_3477_n974,
         DP_OP_425J2_127_3477_n973, DP_OP_425J2_127_3477_n972,
         DP_OP_425J2_127_3477_n971, DP_OP_425J2_127_3477_n970,
         DP_OP_425J2_127_3477_n969, DP_OP_425J2_127_3477_n968,
         DP_OP_425J2_127_3477_n967, DP_OP_425J2_127_3477_n966,
         DP_OP_425J2_127_3477_n965, DP_OP_425J2_127_3477_n964,
         DP_OP_425J2_127_3477_n963, DP_OP_425J2_127_3477_n962,
         DP_OP_425J2_127_3477_n961, DP_OP_425J2_127_3477_n960,
         DP_OP_425J2_127_3477_n959, DP_OP_425J2_127_3477_n958,
         DP_OP_425J2_127_3477_n957, DP_OP_425J2_127_3477_n956,
         DP_OP_425J2_127_3477_n955, DP_OP_425J2_127_3477_n954,
         DP_OP_425J2_127_3477_n953, DP_OP_425J2_127_3477_n952,
         DP_OP_425J2_127_3477_n951, DP_OP_425J2_127_3477_n950,
         DP_OP_425J2_127_3477_n949, DP_OP_425J2_127_3477_n948,
         DP_OP_425J2_127_3477_n947, DP_OP_425J2_127_3477_n946,
         DP_OP_425J2_127_3477_n945, DP_OP_425J2_127_3477_n944,
         DP_OP_425J2_127_3477_n943, DP_OP_425J2_127_3477_n942,
         DP_OP_425J2_127_3477_n941, DP_OP_425J2_127_3477_n940,
         DP_OP_425J2_127_3477_n939, DP_OP_425J2_127_3477_n938,
         DP_OP_425J2_127_3477_n937, DP_OP_425J2_127_3477_n936,
         DP_OP_425J2_127_3477_n935, DP_OP_425J2_127_3477_n934,
         DP_OP_425J2_127_3477_n933, DP_OP_425J2_127_3477_n932,
         DP_OP_425J2_127_3477_n931, DP_OP_425J2_127_3477_n930,
         DP_OP_425J2_127_3477_n929, DP_OP_425J2_127_3477_n928,
         DP_OP_425J2_127_3477_n927, DP_OP_425J2_127_3477_n926,
         DP_OP_425J2_127_3477_n925, DP_OP_425J2_127_3477_n924,
         DP_OP_425J2_127_3477_n923, DP_OP_425J2_127_3477_n922,
         DP_OP_425J2_127_3477_n921, DP_OP_425J2_127_3477_n920,
         DP_OP_425J2_127_3477_n919, DP_OP_425J2_127_3477_n918,
         DP_OP_425J2_127_3477_n917, DP_OP_425J2_127_3477_n916,
         DP_OP_425J2_127_3477_n915, DP_OP_425J2_127_3477_n914,
         DP_OP_425J2_127_3477_n913, DP_OP_425J2_127_3477_n912,
         DP_OP_425J2_127_3477_n911, DP_OP_425J2_127_3477_n910,
         DP_OP_425J2_127_3477_n909, DP_OP_425J2_127_3477_n908,
         DP_OP_425J2_127_3477_n907, DP_OP_425J2_127_3477_n906,
         DP_OP_425J2_127_3477_n905, DP_OP_425J2_127_3477_n904,
         DP_OP_425J2_127_3477_n903, DP_OP_425J2_127_3477_n902,
         DP_OP_425J2_127_3477_n901, DP_OP_425J2_127_3477_n900,
         DP_OP_425J2_127_3477_n899, DP_OP_425J2_127_3477_n898,
         DP_OP_425J2_127_3477_n897, DP_OP_425J2_127_3477_n896,
         DP_OP_425J2_127_3477_n895, DP_OP_425J2_127_3477_n894,
         DP_OP_425J2_127_3477_n893, DP_OP_425J2_127_3477_n892,
         DP_OP_425J2_127_3477_n891, DP_OP_425J2_127_3477_n890,
         DP_OP_425J2_127_3477_n889, DP_OP_425J2_127_3477_n888,
         DP_OP_425J2_127_3477_n887, DP_OP_425J2_127_3477_n886,
         DP_OP_425J2_127_3477_n885, DP_OP_425J2_127_3477_n884,
         DP_OP_425J2_127_3477_n883, DP_OP_425J2_127_3477_n882,
         DP_OP_425J2_127_3477_n881, DP_OP_425J2_127_3477_n880,
         DP_OP_425J2_127_3477_n879, DP_OP_425J2_127_3477_n878,
         DP_OP_425J2_127_3477_n877, DP_OP_425J2_127_3477_n876,
         DP_OP_425J2_127_3477_n875, DP_OP_425J2_127_3477_n874,
         DP_OP_425J2_127_3477_n873, DP_OP_425J2_127_3477_n872,
         DP_OP_425J2_127_3477_n871, DP_OP_425J2_127_3477_n870,
         DP_OP_425J2_127_3477_n869, DP_OP_425J2_127_3477_n868,
         DP_OP_425J2_127_3477_n867, DP_OP_425J2_127_3477_n866,
         DP_OP_425J2_127_3477_n865, DP_OP_425J2_127_3477_n864,
         DP_OP_425J2_127_3477_n863, DP_OP_425J2_127_3477_n862,
         DP_OP_425J2_127_3477_n861, DP_OP_425J2_127_3477_n860,
         DP_OP_425J2_127_3477_n859, DP_OP_425J2_127_3477_n858,
         DP_OP_425J2_127_3477_n857, DP_OP_425J2_127_3477_n856,
         DP_OP_425J2_127_3477_n855, DP_OP_425J2_127_3477_n854,
         DP_OP_425J2_127_3477_n853, DP_OP_425J2_127_3477_n852,
         DP_OP_425J2_127_3477_n851, DP_OP_425J2_127_3477_n850,
         DP_OP_425J2_127_3477_n849, DP_OP_425J2_127_3477_n848,
         DP_OP_425J2_127_3477_n847, DP_OP_425J2_127_3477_n846,
         DP_OP_425J2_127_3477_n845, DP_OP_425J2_127_3477_n844,
         DP_OP_425J2_127_3477_n843, DP_OP_425J2_127_3477_n842,
         DP_OP_425J2_127_3477_n841, DP_OP_425J2_127_3477_n840,
         DP_OP_425J2_127_3477_n839, DP_OP_425J2_127_3477_n838,
         DP_OP_425J2_127_3477_n837, DP_OP_425J2_127_3477_n836,
         DP_OP_425J2_127_3477_n835, DP_OP_425J2_127_3477_n834,
         DP_OP_425J2_127_3477_n833, DP_OP_425J2_127_3477_n832,
         DP_OP_425J2_127_3477_n831, DP_OP_425J2_127_3477_n830,
         DP_OP_425J2_127_3477_n829, DP_OP_425J2_127_3477_n828,
         DP_OP_425J2_127_3477_n827, DP_OP_425J2_127_3477_n826,
         DP_OP_425J2_127_3477_n825, DP_OP_425J2_127_3477_n823,
         DP_OP_425J2_127_3477_n822, DP_OP_425J2_127_3477_n821,
         DP_OP_425J2_127_3477_n820, DP_OP_425J2_127_3477_n819,
         DP_OP_425J2_127_3477_n818, DP_OP_425J2_127_3477_n817,
         DP_OP_425J2_127_3477_n816, DP_OP_425J2_127_3477_n815,
         DP_OP_425J2_127_3477_n814, DP_OP_425J2_127_3477_n813,
         DP_OP_425J2_127_3477_n812, DP_OP_425J2_127_3477_n811,
         DP_OP_425J2_127_3477_n810, DP_OP_425J2_127_3477_n809,
         DP_OP_425J2_127_3477_n808, DP_OP_425J2_127_3477_n807,
         DP_OP_425J2_127_3477_n806, DP_OP_425J2_127_3477_n805,
         DP_OP_425J2_127_3477_n804, DP_OP_425J2_127_3477_n803,
         DP_OP_425J2_127_3477_n802, DP_OP_425J2_127_3477_n801,
         DP_OP_425J2_127_3477_n800, DP_OP_425J2_127_3477_n799,
         DP_OP_425J2_127_3477_n798, DP_OP_425J2_127_3477_n797,
         DP_OP_425J2_127_3477_n796, DP_OP_425J2_127_3477_n795,
         DP_OP_425J2_127_3477_n794, DP_OP_425J2_127_3477_n793,
         DP_OP_425J2_127_3477_n792, DP_OP_425J2_127_3477_n791,
         DP_OP_425J2_127_3477_n790, DP_OP_425J2_127_3477_n789,
         DP_OP_425J2_127_3477_n788, DP_OP_425J2_127_3477_n787,
         DP_OP_425J2_127_3477_n786, DP_OP_425J2_127_3477_n785,
         DP_OP_425J2_127_3477_n784, DP_OP_425J2_127_3477_n783,
         DP_OP_425J2_127_3477_n782, DP_OP_425J2_127_3477_n781,
         DP_OP_425J2_127_3477_n780, DP_OP_425J2_127_3477_n779,
         DP_OP_425J2_127_3477_n778, DP_OP_425J2_127_3477_n777,
         DP_OP_425J2_127_3477_n776, DP_OP_425J2_127_3477_n775,
         DP_OP_425J2_127_3477_n774, DP_OP_425J2_127_3477_n773,
         DP_OP_425J2_127_3477_n772, DP_OP_425J2_127_3477_n771,
         DP_OP_425J2_127_3477_n770, DP_OP_425J2_127_3477_n769,
         DP_OP_425J2_127_3477_n768, DP_OP_425J2_127_3477_n767,
         DP_OP_425J2_127_3477_n766, DP_OP_425J2_127_3477_n765,
         DP_OP_425J2_127_3477_n764, DP_OP_425J2_127_3477_n763,
         DP_OP_425J2_127_3477_n762, DP_OP_425J2_127_3477_n761,
         DP_OP_425J2_127_3477_n760, DP_OP_425J2_127_3477_n759,
         DP_OP_425J2_127_3477_n758, DP_OP_425J2_127_3477_n757,
         DP_OP_425J2_127_3477_n756, DP_OP_425J2_127_3477_n755,
         DP_OP_425J2_127_3477_n754, DP_OP_425J2_127_3477_n753,
         DP_OP_425J2_127_3477_n752, DP_OP_425J2_127_3477_n751,
         DP_OP_425J2_127_3477_n750, DP_OP_425J2_127_3477_n749,
         DP_OP_425J2_127_3477_n748, DP_OP_425J2_127_3477_n747,
         DP_OP_425J2_127_3477_n746, DP_OP_425J2_127_3477_n745,
         DP_OP_425J2_127_3477_n744, DP_OP_425J2_127_3477_n743,
         DP_OP_425J2_127_3477_n742, DP_OP_425J2_127_3477_n741,
         DP_OP_425J2_127_3477_n740, DP_OP_425J2_127_3477_n739,
         DP_OP_425J2_127_3477_n738, DP_OP_425J2_127_3477_n737,
         DP_OP_425J2_127_3477_n736, DP_OP_425J2_127_3477_n735,
         DP_OP_425J2_127_3477_n734, DP_OP_425J2_127_3477_n733,
         DP_OP_425J2_127_3477_n732, DP_OP_425J2_127_3477_n731,
         DP_OP_425J2_127_3477_n730, DP_OP_425J2_127_3477_n729,
         DP_OP_425J2_127_3477_n728, DP_OP_425J2_127_3477_n727,
         DP_OP_425J2_127_3477_n726, DP_OP_425J2_127_3477_n725,
         DP_OP_425J2_127_3477_n724, DP_OP_425J2_127_3477_n723,
         DP_OP_425J2_127_3477_n722, DP_OP_425J2_127_3477_n721,
         DP_OP_425J2_127_3477_n720, DP_OP_425J2_127_3477_n719,
         DP_OP_425J2_127_3477_n718, DP_OP_425J2_127_3477_n717,
         DP_OP_425J2_127_3477_n716, DP_OP_425J2_127_3477_n715,
         DP_OP_425J2_127_3477_n714, DP_OP_425J2_127_3477_n713,
         DP_OP_425J2_127_3477_n712, DP_OP_425J2_127_3477_n711,
         DP_OP_425J2_127_3477_n710, DP_OP_425J2_127_3477_n709,
         DP_OP_425J2_127_3477_n708, DP_OP_425J2_127_3477_n707,
         DP_OP_425J2_127_3477_n706, DP_OP_425J2_127_3477_n705,
         DP_OP_425J2_127_3477_n704, DP_OP_425J2_127_3477_n703,
         DP_OP_425J2_127_3477_n702, DP_OP_425J2_127_3477_n701,
         DP_OP_425J2_127_3477_n700, DP_OP_425J2_127_3477_n699,
         DP_OP_425J2_127_3477_n698, DP_OP_425J2_127_3477_n697,
         DP_OP_425J2_127_3477_n696, DP_OP_425J2_127_3477_n695,
         DP_OP_425J2_127_3477_n694, DP_OP_425J2_127_3477_n693,
         DP_OP_425J2_127_3477_n692, DP_OP_425J2_127_3477_n691,
         DP_OP_425J2_127_3477_n690, DP_OP_425J2_127_3477_n689,
         DP_OP_425J2_127_3477_n688, DP_OP_425J2_127_3477_n687,
         DP_OP_425J2_127_3477_n686, DP_OP_425J2_127_3477_n685,
         DP_OP_425J2_127_3477_n684, DP_OP_425J2_127_3477_n683,
         DP_OP_425J2_127_3477_n682, DP_OP_425J2_127_3477_n681,
         DP_OP_425J2_127_3477_n680, DP_OP_425J2_127_3477_n679,
         DP_OP_425J2_127_3477_n678, DP_OP_425J2_127_3477_n677,
         DP_OP_425J2_127_3477_n676, DP_OP_425J2_127_3477_n675,
         DP_OP_425J2_127_3477_n674, DP_OP_425J2_127_3477_n673,
         DP_OP_425J2_127_3477_n672, DP_OP_425J2_127_3477_n671,
         DP_OP_425J2_127_3477_n670, DP_OP_425J2_127_3477_n669,
         DP_OP_425J2_127_3477_n668, DP_OP_425J2_127_3477_n667,
         DP_OP_425J2_127_3477_n666, DP_OP_425J2_127_3477_n665,
         DP_OP_425J2_127_3477_n664, DP_OP_425J2_127_3477_n663,
         DP_OP_425J2_127_3477_n662, DP_OP_425J2_127_3477_n661,
         DP_OP_425J2_127_3477_n660, DP_OP_425J2_127_3477_n659,
         DP_OP_425J2_127_3477_n658, DP_OP_425J2_127_3477_n657,
         DP_OP_425J2_127_3477_n656, DP_OP_425J2_127_3477_n655,
         DP_OP_425J2_127_3477_n654, DP_OP_425J2_127_3477_n653,
         DP_OP_425J2_127_3477_n652, DP_OP_425J2_127_3477_n651,
         DP_OP_425J2_127_3477_n650, DP_OP_425J2_127_3477_n649,
         DP_OP_425J2_127_3477_n648, DP_OP_425J2_127_3477_n647,
         DP_OP_425J2_127_3477_n646, DP_OP_425J2_127_3477_n645,
         DP_OP_425J2_127_3477_n644, DP_OP_425J2_127_3477_n643,
         DP_OP_425J2_127_3477_n642, DP_OP_425J2_127_3477_n641,
         DP_OP_425J2_127_3477_n640, DP_OP_425J2_127_3477_n639,
         DP_OP_425J2_127_3477_n638, DP_OP_425J2_127_3477_n637,
         DP_OP_425J2_127_3477_n636, DP_OP_425J2_127_3477_n635,
         DP_OP_425J2_127_3477_n634, DP_OP_425J2_127_3477_n633,
         DP_OP_425J2_127_3477_n632, DP_OP_425J2_127_3477_n631,
         DP_OP_425J2_127_3477_n630, DP_OP_425J2_127_3477_n629,
         DP_OP_425J2_127_3477_n628, DP_OP_425J2_127_3477_n627,
         DP_OP_425J2_127_3477_n626, DP_OP_425J2_127_3477_n625,
         DP_OP_425J2_127_3477_n624, DP_OP_425J2_127_3477_n623,
         DP_OP_425J2_127_3477_n622, DP_OP_425J2_127_3477_n621,
         DP_OP_425J2_127_3477_n620, DP_OP_425J2_127_3477_n619,
         DP_OP_425J2_127_3477_n618, DP_OP_425J2_127_3477_n617,
         DP_OP_425J2_127_3477_n616, DP_OP_425J2_127_3477_n615,
         DP_OP_425J2_127_3477_n614, DP_OP_425J2_127_3477_n613,
         DP_OP_425J2_127_3477_n612, DP_OP_425J2_127_3477_n611,
         DP_OP_425J2_127_3477_n610, DP_OP_425J2_127_3477_n609,
         DP_OP_425J2_127_3477_n608, DP_OP_425J2_127_3477_n607,
         DP_OP_425J2_127_3477_n606, DP_OP_425J2_127_3477_n605,
         DP_OP_425J2_127_3477_n604, DP_OP_425J2_127_3477_n603,
         DP_OP_425J2_127_3477_n602, DP_OP_425J2_127_3477_n601,
         DP_OP_425J2_127_3477_n600, DP_OP_425J2_127_3477_n599,
         DP_OP_425J2_127_3477_n598, DP_OP_425J2_127_3477_n597,
         DP_OP_425J2_127_3477_n596, DP_OP_425J2_127_3477_n595,
         DP_OP_425J2_127_3477_n594, DP_OP_425J2_127_3477_n593,
         DP_OP_425J2_127_3477_n592, DP_OP_425J2_127_3477_n591,
         DP_OP_425J2_127_3477_n590, DP_OP_425J2_127_3477_n589,
         DP_OP_425J2_127_3477_n588, DP_OP_425J2_127_3477_n587,
         DP_OP_425J2_127_3477_n586, DP_OP_425J2_127_3477_n585,
         DP_OP_425J2_127_3477_n584, DP_OP_425J2_127_3477_n583,
         DP_OP_425J2_127_3477_n582, DP_OP_425J2_127_3477_n581,
         DP_OP_425J2_127_3477_n580, DP_OP_425J2_127_3477_n579,
         DP_OP_425J2_127_3477_n578, DP_OP_425J2_127_3477_n577,
         DP_OP_425J2_127_3477_n576, DP_OP_425J2_127_3477_n575,
         DP_OP_425J2_127_3477_n574, DP_OP_425J2_127_3477_n573,
         DP_OP_425J2_127_3477_n572, DP_OP_425J2_127_3477_n571,
         DP_OP_425J2_127_3477_n570, DP_OP_425J2_127_3477_n569,
         DP_OP_425J2_127_3477_n568, DP_OP_425J2_127_3477_n567,
         DP_OP_425J2_127_3477_n566, DP_OP_425J2_127_3477_n565,
         DP_OP_425J2_127_3477_n564, DP_OP_425J2_127_3477_n563,
         DP_OP_425J2_127_3477_n562, DP_OP_425J2_127_3477_n561,
         DP_OP_425J2_127_3477_n560, DP_OP_425J2_127_3477_n559,
         DP_OP_425J2_127_3477_n558, DP_OP_425J2_127_3477_n557,
         DP_OP_425J2_127_3477_n556, DP_OP_425J2_127_3477_n555,
         DP_OP_425J2_127_3477_n554, DP_OP_425J2_127_3477_n553,
         DP_OP_425J2_127_3477_n552, DP_OP_425J2_127_3477_n551,
         DP_OP_425J2_127_3477_n550, DP_OP_425J2_127_3477_n549,
         DP_OP_425J2_127_3477_n548, DP_OP_425J2_127_3477_n547,
         DP_OP_425J2_127_3477_n546, DP_OP_425J2_127_3477_n545,
         DP_OP_425J2_127_3477_n544, DP_OP_425J2_127_3477_n543,
         DP_OP_425J2_127_3477_n542, DP_OP_425J2_127_3477_n541,
         DP_OP_425J2_127_3477_n540, DP_OP_425J2_127_3477_n539,
         DP_OP_425J2_127_3477_n538, DP_OP_425J2_127_3477_n537,
         DP_OP_425J2_127_3477_n536, DP_OP_425J2_127_3477_n535,
         DP_OP_425J2_127_3477_n534, DP_OP_425J2_127_3477_n533,
         DP_OP_425J2_127_3477_n532, DP_OP_425J2_127_3477_n531,
         DP_OP_425J2_127_3477_n530, DP_OP_425J2_127_3477_n529,
         DP_OP_425J2_127_3477_n528, DP_OP_425J2_127_3477_n527,
         DP_OP_425J2_127_3477_n526, DP_OP_425J2_127_3477_n525,
         DP_OP_425J2_127_3477_n524, DP_OP_425J2_127_3477_n523,
         DP_OP_425J2_127_3477_n522, DP_OP_425J2_127_3477_n521,
         DP_OP_425J2_127_3477_n520, DP_OP_425J2_127_3477_n519,
         DP_OP_425J2_127_3477_n518, DP_OP_425J2_127_3477_n517,
         DP_OP_425J2_127_3477_n516, DP_OP_425J2_127_3477_n515,
         DP_OP_425J2_127_3477_n514, DP_OP_425J2_127_3477_n513,
         DP_OP_425J2_127_3477_n512, DP_OP_425J2_127_3477_n511,
         DP_OP_425J2_127_3477_n510, DP_OP_425J2_127_3477_n509,
         DP_OP_425J2_127_3477_n508, DP_OP_425J2_127_3477_n507,
         DP_OP_425J2_127_3477_n506, DP_OP_425J2_127_3477_n505,
         DP_OP_425J2_127_3477_n504, DP_OP_425J2_127_3477_n503,
         DP_OP_425J2_127_3477_n502, DP_OP_425J2_127_3477_n501,
         DP_OP_425J2_127_3477_n500, DP_OP_425J2_127_3477_n499,
         DP_OP_425J2_127_3477_n498, DP_OP_425J2_127_3477_n497,
         DP_OP_425J2_127_3477_n496, DP_OP_425J2_127_3477_n495,
         DP_OP_425J2_127_3477_n494, DP_OP_425J2_127_3477_n493,
         DP_OP_425J2_127_3477_n492, DP_OP_425J2_127_3477_n491,
         DP_OP_425J2_127_3477_n490, DP_OP_425J2_127_3477_n489,
         DP_OP_425J2_127_3477_n488, DP_OP_425J2_127_3477_n487,
         DP_OP_425J2_127_3477_n486, DP_OP_425J2_127_3477_n485,
         DP_OP_425J2_127_3477_n484, DP_OP_425J2_127_3477_n483,
         DP_OP_425J2_127_3477_n482, DP_OP_425J2_127_3477_n481,
         DP_OP_425J2_127_3477_n480, DP_OP_425J2_127_3477_n479,
         DP_OP_425J2_127_3477_n478, DP_OP_425J2_127_3477_n477,
         DP_OP_425J2_127_3477_n476, DP_OP_425J2_127_3477_n475,
         DP_OP_425J2_127_3477_n474, DP_OP_425J2_127_3477_n473,
         DP_OP_425J2_127_3477_n472, DP_OP_425J2_127_3477_n471,
         DP_OP_425J2_127_3477_n470, DP_OP_425J2_127_3477_n469,
         DP_OP_425J2_127_3477_n468, DP_OP_425J2_127_3477_n467,
         DP_OP_425J2_127_3477_n466, DP_OP_425J2_127_3477_n465,
         DP_OP_425J2_127_3477_n464, DP_OP_425J2_127_3477_n463,
         DP_OP_425J2_127_3477_n462, DP_OP_425J2_127_3477_n461,
         DP_OP_425J2_127_3477_n460, DP_OP_425J2_127_3477_n459,
         DP_OP_425J2_127_3477_n458, DP_OP_425J2_127_3477_n457,
         DP_OP_425J2_127_3477_n456, DP_OP_425J2_127_3477_n455,
         DP_OP_425J2_127_3477_n454, DP_OP_425J2_127_3477_n453,
         DP_OP_425J2_127_3477_n452, DP_OP_425J2_127_3477_n451,
         DP_OP_425J2_127_3477_n450, DP_OP_425J2_127_3477_n449,
         DP_OP_425J2_127_3477_n448, DP_OP_425J2_127_3477_n447,
         DP_OP_425J2_127_3477_n446, DP_OP_425J2_127_3477_n445,
         DP_OP_425J2_127_3477_n444, DP_OP_425J2_127_3477_n443,
         DP_OP_425J2_127_3477_n442, DP_OP_425J2_127_3477_n441,
         DP_OP_425J2_127_3477_n440, DP_OP_425J2_127_3477_n439,
         DP_OP_425J2_127_3477_n438, DP_OP_425J2_127_3477_n437,
         DP_OP_425J2_127_3477_n436, DP_OP_425J2_127_3477_n435,
         DP_OP_425J2_127_3477_n434, DP_OP_425J2_127_3477_n433,
         DP_OP_425J2_127_3477_n432, DP_OP_425J2_127_3477_n431,
         DP_OP_425J2_127_3477_n430, DP_OP_425J2_127_3477_n429,
         DP_OP_425J2_127_3477_n428, DP_OP_425J2_127_3477_n427,
         DP_OP_425J2_127_3477_n426, DP_OP_425J2_127_3477_n425,
         DP_OP_425J2_127_3477_n424, DP_OP_425J2_127_3477_n423,
         DP_OP_425J2_127_3477_n422, DP_OP_425J2_127_3477_n421,
         DP_OP_425J2_127_3477_n420, DP_OP_425J2_127_3477_n419,
         DP_OP_425J2_127_3477_n418, DP_OP_425J2_127_3477_n417,
         DP_OP_425J2_127_3477_n416, DP_OP_425J2_127_3477_n415,
         DP_OP_425J2_127_3477_n414, DP_OP_425J2_127_3477_n413,
         DP_OP_425J2_127_3477_n412, DP_OP_425J2_127_3477_n411,
         DP_OP_425J2_127_3477_n410, DP_OP_425J2_127_3477_n409,
         DP_OP_425J2_127_3477_n408, DP_OP_425J2_127_3477_n407,
         DP_OP_425J2_127_3477_n406, DP_OP_425J2_127_3477_n405,
         DP_OP_425J2_127_3477_n404, DP_OP_425J2_127_3477_n403,
         DP_OP_425J2_127_3477_n402, DP_OP_425J2_127_3477_n401,
         DP_OP_425J2_127_3477_n400, DP_OP_425J2_127_3477_n399,
         DP_OP_425J2_127_3477_n398, DP_OP_425J2_127_3477_n397,
         DP_OP_425J2_127_3477_n396, DP_OP_425J2_127_3477_n395,
         DP_OP_425J2_127_3477_n394, DP_OP_425J2_127_3477_n393,
         DP_OP_425J2_127_3477_n392, DP_OP_425J2_127_3477_n391,
         DP_OP_425J2_127_3477_n390, DP_OP_425J2_127_3477_n389,
         DP_OP_425J2_127_3477_n388, DP_OP_425J2_127_3477_n387,
         DP_OP_425J2_127_3477_n386, DP_OP_425J2_127_3477_n385,
         DP_OP_425J2_127_3477_n384, DP_OP_425J2_127_3477_n383,
         DP_OP_425J2_127_3477_n382, DP_OP_425J2_127_3477_n381,
         DP_OP_425J2_127_3477_n380, DP_OP_425J2_127_3477_n379,
         DP_OP_425J2_127_3477_n378, DP_OP_425J2_127_3477_n377,
         DP_OP_425J2_127_3477_n376, DP_OP_425J2_127_3477_n375,
         DP_OP_425J2_127_3477_n374, DP_OP_425J2_127_3477_n373,
         DP_OP_425J2_127_3477_n372, DP_OP_425J2_127_3477_n371,
         DP_OP_425J2_127_3477_n370, DP_OP_425J2_127_3477_n369,
         DP_OP_425J2_127_3477_n368, DP_OP_425J2_127_3477_n367,
         DP_OP_425J2_127_3477_n366, DP_OP_425J2_127_3477_n365,
         DP_OP_425J2_127_3477_n364, DP_OP_425J2_127_3477_n363,
         DP_OP_425J2_127_3477_n362, DP_OP_425J2_127_3477_n361,
         DP_OP_425J2_127_3477_n360, DP_OP_425J2_127_3477_n359,
         DP_OP_425J2_127_3477_n358, DP_OP_425J2_127_3477_n357,
         DP_OP_425J2_127_3477_n356, DP_OP_425J2_127_3477_n355,
         DP_OP_425J2_127_3477_n354, DP_OP_425J2_127_3477_n353,
         DP_OP_425J2_127_3477_n352, DP_OP_425J2_127_3477_n351,
         DP_OP_425J2_127_3477_n350, DP_OP_425J2_127_3477_n349,
         DP_OP_425J2_127_3477_n348, DP_OP_425J2_127_3477_n347,
         DP_OP_425J2_127_3477_n346, DP_OP_425J2_127_3477_n345,
         DP_OP_425J2_127_3477_n344, DP_OP_425J2_127_3477_n343,
         DP_OP_425J2_127_3477_n342, DP_OP_425J2_127_3477_n341,
         DP_OP_425J2_127_3477_n340, DP_OP_425J2_127_3477_n339,
         DP_OP_425J2_127_3477_n338, DP_OP_425J2_127_3477_n337,
         DP_OP_425J2_127_3477_n336, DP_OP_425J2_127_3477_n335,
         DP_OP_425J2_127_3477_n334, DP_OP_425J2_127_3477_n333,
         DP_OP_425J2_127_3477_n332, DP_OP_425J2_127_3477_n330,
         DP_OP_425J2_127_3477_n329, DP_OP_425J2_127_3477_n328,
         DP_OP_425J2_127_3477_n327, DP_OP_425J2_127_3477_n326,
         DP_OP_425J2_127_3477_n325, DP_OP_425J2_127_3477_n324,
         DP_OP_425J2_127_3477_n323, DP_OP_425J2_127_3477_n322,
         DP_OP_425J2_127_3477_n321, DP_OP_425J2_127_3477_n320,
         DP_OP_425J2_127_3477_n319, DP_OP_425J2_127_3477_n318,
         DP_OP_425J2_127_3477_n317, DP_OP_425J2_127_3477_n316,
         DP_OP_425J2_127_3477_n315, DP_OP_425J2_127_3477_n314,
         DP_OP_425J2_127_3477_n313, DP_OP_425J2_127_3477_n312,
         DP_OP_425J2_127_3477_n311, DP_OP_425J2_127_3477_n310,
         DP_OP_425J2_127_3477_n309, DP_OP_425J2_127_3477_n308,
         DP_OP_425J2_127_3477_n307, DP_OP_425J2_127_3477_n306,
         DP_OP_425J2_127_3477_n305, DP_OP_425J2_127_3477_n304,
         DP_OP_425J2_127_3477_n303, DP_OP_425J2_127_3477_n302,
         DP_OP_425J2_127_3477_n297, DP_OP_425J2_127_3477_n295,
         DP_OP_425J2_127_3477_n287, DP_OP_425J2_127_3477_n286,
         DP_OP_425J2_127_3477_n285, DP_OP_425J2_127_3477_n284,
         DP_OP_425J2_127_3477_n283, DP_OP_425J2_127_3477_n282,
         DP_OP_425J2_127_3477_n281, DP_OP_425J2_127_3477_n280,
         DP_OP_425J2_127_3477_n279, DP_OP_425J2_127_3477_n277,
         DP_OP_425J2_127_3477_n276, DP_OP_425J2_127_3477_n274,
         DP_OP_425J2_127_3477_n272, DP_OP_425J2_127_3477_n269,
         DP_OP_425J2_127_3477_n268, DP_OP_425J2_127_3477_n267,
         DP_OP_425J2_127_3477_n266, DP_OP_425J2_127_3477_n265,
         DP_OP_425J2_127_3477_n261, DP_OP_425J2_127_3477_n260,
         DP_OP_425J2_127_3477_n259, DP_OP_425J2_127_3477_n257,
         DP_OP_425J2_127_3477_n255, DP_OP_425J2_127_3477_n252,
         DP_OP_425J2_127_3477_n250, DP_OP_425J2_127_3477_n249,
         DP_OP_425J2_127_3477_n245, DP_OP_425J2_127_3477_n244,
         DP_OP_425J2_127_3477_n240, DP_OP_425J2_127_3477_n237,
         DP_OP_425J2_127_3477_n236, DP_OP_425J2_127_3477_n233,
         DP_OP_425J2_127_3477_n226, DP_OP_425J2_127_3477_n220,
         DP_OP_425J2_127_3477_n219, DP_OP_425J2_127_3477_n217,
         DP_OP_425J2_127_3477_n214, DP_OP_425J2_127_3477_n213,
         DP_OP_425J2_127_3477_n212, DP_OP_425J2_127_3477_n210,
         DP_OP_425J2_127_3477_n209, DP_OP_425J2_127_3477_n207,
         DP_OP_425J2_127_3477_n203, DP_OP_425J2_127_3477_n202,
         DP_OP_425J2_127_3477_n201, DP_OP_425J2_127_3477_n198,
         DP_OP_425J2_127_3477_n197, DP_OP_425J2_127_3477_n190,
         DP_OP_425J2_127_3477_n189, DP_OP_425J2_127_3477_n187,
         DP_OP_425J2_127_3477_n185, DP_OP_425J2_127_3477_n182,
         DP_OP_425J2_127_3477_n178, DP_OP_425J2_127_3477_n176,
         DP_OP_425J2_127_3477_n174, DP_OP_425J2_127_3477_n171,
         DP_OP_425J2_127_3477_n168, DP_OP_425J2_127_3477_n167,
         DP_OP_425J2_127_3477_n166, DP_OP_425J2_127_3477_n165,
         DP_OP_425J2_127_3477_n162, DP_OP_425J2_127_3477_n160,
         DP_OP_425J2_127_3477_n158, DP_OP_425J2_127_3477_n156,
         DP_OP_425J2_127_3477_n153, DP_OP_425J2_127_3477_n151,
         DP_OP_425J2_127_3477_n149, DP_OP_425J2_127_3477_n148,
         DP_OP_425J2_127_3477_n146, DP_OP_425J2_127_3477_n145,
         DP_OP_425J2_127_3477_n144, DP_OP_425J2_127_3477_n142,
         DP_OP_425J2_127_3477_n141, DP_OP_425J2_127_3477_n140,
         DP_OP_425J2_127_3477_n136, DP_OP_425J2_127_3477_n133,
         DP_OP_425J2_127_3477_n132, DP_OP_425J2_127_3477_n131,
         DP_OP_425J2_127_3477_n129, DP_OP_425J2_127_3477_n128,
         DP_OP_425J2_127_3477_n127, DP_OP_425J2_127_3477_n126,
         DP_OP_425J2_127_3477_n124, DP_OP_425J2_127_3477_n122,
         DP_OP_425J2_127_3477_n120, DP_OP_425J2_127_3477_n115,
         DP_OP_425J2_127_3477_n114, DP_OP_425J2_127_3477_n111,
         DP_OP_425J2_127_3477_n110, DP_OP_425J2_127_3477_n109,
         DP_OP_425J2_127_3477_n107, DP_OP_425J2_127_3477_n105,
         DP_OP_425J2_127_3477_n102, DP_OP_425J2_127_3477_n101,
         DP_OP_425J2_127_3477_n100, DP_OP_425J2_127_3477_n98,
         DP_OP_425J2_127_3477_n97, DP_OP_425J2_127_3477_n96,
         DP_OP_425J2_127_3477_n95, DP_OP_425J2_127_3477_n93,
         DP_OP_425J2_127_3477_n91, DP_OP_425J2_127_3477_n89,
         DP_OP_425J2_127_3477_n85, DP_OP_425J2_127_3477_n82,
         DP_OP_425J2_127_3477_n80, DP_OP_425J2_127_3477_n78,
         DP_OP_425J2_127_3477_n77, DP_OP_425J2_127_3477_n75,
         DP_OP_425J2_127_3477_n73, DP_OP_425J2_127_3477_n72,
         DP_OP_425J2_127_3477_n71, DP_OP_425J2_127_3477_n69,
         DP_OP_425J2_127_3477_n67, DP_OP_425J2_127_3477_n65,
         DP_OP_425J2_127_3477_n60, DP_OP_425J2_127_3477_n58,
         DP_OP_425J2_127_3477_n57, DP_OP_425J2_127_3477_n56,
         DP_OP_425J2_127_3477_n54, DP_OP_425J2_127_3477_n52,
         DP_OP_425J2_127_3477_n51, DP_OP_425J2_127_3477_n50,
         DP_OP_425J2_127_3477_n49, DP_OP_425J2_127_3477_n47,
         DP_OP_425J2_127_3477_n38, DP_OP_425J2_127_3477_n22,
         DP_OP_425J2_127_3477_n19, DP_OP_425J2_127_3477_n17,
         DP_OP_425J2_127_3477_n15, DP_OP_425J2_127_3477_n13,
         DP_OP_425J2_127_3477_n12, DP_OP_425J2_127_3477_n5,
         DP_OP_424J2_126_3477_n3066, DP_OP_424J2_126_3477_n3065,
         DP_OP_424J2_126_3477_n3063, DP_OP_424J2_126_3477_n3060,
         DP_OP_424J2_126_3477_n3059, DP_OP_424J2_126_3477_n3058,
         DP_OP_424J2_126_3477_n3057, DP_OP_424J2_126_3477_n3055,
         DP_OP_424J2_126_3477_n3054, DP_OP_424J2_126_3477_n3053,
         DP_OP_424J2_126_3477_n3052, DP_OP_424J2_126_3477_n3051,
         DP_OP_424J2_126_3477_n3050, DP_OP_424J2_126_3477_n3049,
         DP_OP_424J2_126_3477_n3048, DP_OP_424J2_126_3477_n3047,
         DP_OP_424J2_126_3477_n3046, DP_OP_424J2_126_3477_n3045,
         DP_OP_424J2_126_3477_n3044, DP_OP_424J2_126_3477_n3043,
         DP_OP_424J2_126_3477_n3042, DP_OP_424J2_126_3477_n3041,
         DP_OP_424J2_126_3477_n3040, DP_OP_424J2_126_3477_n3039,
         DP_OP_424J2_126_3477_n3038, DP_OP_424J2_126_3477_n3037,
         DP_OP_424J2_126_3477_n3036, DP_OP_424J2_126_3477_n3035,
         DP_OP_424J2_126_3477_n3034, DP_OP_424J2_126_3477_n3033,
         DP_OP_424J2_126_3477_n3032, DP_OP_424J2_126_3477_n3031,
         DP_OP_424J2_126_3477_n3030, DP_OP_424J2_126_3477_n3029,
         DP_OP_424J2_126_3477_n3028, DP_OP_424J2_126_3477_n3027,
         DP_OP_424J2_126_3477_n3026, DP_OP_424J2_126_3477_n3025,
         DP_OP_424J2_126_3477_n3023, DP_OP_424J2_126_3477_n3020,
         DP_OP_424J2_126_3477_n3019, DP_OP_424J2_126_3477_n3015,
         DP_OP_424J2_126_3477_n3013, DP_OP_424J2_126_3477_n3012,
         DP_OP_424J2_126_3477_n3011, DP_OP_424J2_126_3477_n3010,
         DP_OP_424J2_126_3477_n3009, DP_OP_424J2_126_3477_n3008,
         DP_OP_424J2_126_3477_n3007, DP_OP_424J2_126_3477_n3006,
         DP_OP_424J2_126_3477_n3005, DP_OP_424J2_126_3477_n3004,
         DP_OP_424J2_126_3477_n3003, DP_OP_424J2_126_3477_n3002,
         DP_OP_424J2_126_3477_n3001, DP_OP_424J2_126_3477_n3000,
         DP_OP_424J2_126_3477_n2999, DP_OP_424J2_126_3477_n2998,
         DP_OP_424J2_126_3477_n2997, DP_OP_424J2_126_3477_n2996,
         DP_OP_424J2_126_3477_n2995, DP_OP_424J2_126_3477_n2994,
         DP_OP_424J2_126_3477_n2993, DP_OP_424J2_126_3477_n2992,
         DP_OP_424J2_126_3477_n2991, DP_OP_424J2_126_3477_n2990,
         DP_OP_424J2_126_3477_n2989, DP_OP_424J2_126_3477_n2988,
         DP_OP_424J2_126_3477_n2987, DP_OP_424J2_126_3477_n2986,
         DP_OP_424J2_126_3477_n2985, DP_OP_424J2_126_3477_n2984,
         DP_OP_424J2_126_3477_n2983, DP_OP_424J2_126_3477_n2982,
         DP_OP_424J2_126_3477_n2980, DP_OP_424J2_126_3477_n2979,
         DP_OP_424J2_126_3477_n2977, DP_OP_424J2_126_3477_n2976,
         DP_OP_424J2_126_3477_n2975, DP_OP_424J2_126_3477_n2974,
         DP_OP_424J2_126_3477_n2973, DP_OP_424J2_126_3477_n2972,
         DP_OP_424J2_126_3477_n2971, DP_OP_424J2_126_3477_n2970,
         DP_OP_424J2_126_3477_n2969, DP_OP_424J2_126_3477_n2968,
         DP_OP_424J2_126_3477_n2967, DP_OP_424J2_126_3477_n2966,
         DP_OP_424J2_126_3477_n2965, DP_OP_424J2_126_3477_n2964,
         DP_OP_424J2_126_3477_n2963, DP_OP_424J2_126_3477_n2962,
         DP_OP_424J2_126_3477_n2961, DP_OP_424J2_126_3477_n2960,
         DP_OP_424J2_126_3477_n2959, DP_OP_424J2_126_3477_n2958,
         DP_OP_424J2_126_3477_n2957, DP_OP_424J2_126_3477_n2956,
         DP_OP_424J2_126_3477_n2955, DP_OP_424J2_126_3477_n2954,
         DP_OP_424J2_126_3477_n2953, DP_OP_424J2_126_3477_n2951,
         DP_OP_424J2_126_3477_n2950, DP_OP_424J2_126_3477_n2949,
         DP_OP_424J2_126_3477_n2948, DP_OP_424J2_126_3477_n2947,
         DP_OP_424J2_126_3477_n2946, DP_OP_424J2_126_3477_n2945,
         DP_OP_424J2_126_3477_n2944, DP_OP_424J2_126_3477_n2943,
         DP_OP_424J2_126_3477_n2942, DP_OP_424J2_126_3477_n2941,
         DP_OP_424J2_126_3477_n2940, DP_OP_424J2_126_3477_n2939,
         DP_OP_424J2_126_3477_n2938, DP_OP_424J2_126_3477_n2936,
         DP_OP_424J2_126_3477_n2933, DP_OP_424J2_126_3477_n2932,
         DP_OP_424J2_126_3477_n2929, DP_OP_424J2_126_3477_n2928,
         DP_OP_424J2_126_3477_n2927, DP_OP_424J2_126_3477_n2925,
         DP_OP_424J2_126_3477_n2924, DP_OP_424J2_126_3477_n2923,
         DP_OP_424J2_126_3477_n2922, DP_OP_424J2_126_3477_n2921,
         DP_OP_424J2_126_3477_n2920, DP_OP_424J2_126_3477_n2919,
         DP_OP_424J2_126_3477_n2918, DP_OP_424J2_126_3477_n2917,
         DP_OP_424J2_126_3477_n2916, DP_OP_424J2_126_3477_n2915,
         DP_OP_424J2_126_3477_n2914, DP_OP_424J2_126_3477_n2913,
         DP_OP_424J2_126_3477_n2912, DP_OP_424J2_126_3477_n2911,
         DP_OP_424J2_126_3477_n2910, DP_OP_424J2_126_3477_n2908,
         DP_OP_424J2_126_3477_n2907, DP_OP_424J2_126_3477_n2906,
         DP_OP_424J2_126_3477_n2905, DP_OP_424J2_126_3477_n2904,
         DP_OP_424J2_126_3477_n2903, DP_OP_424J2_126_3477_n2902,
         DP_OP_424J2_126_3477_n2901, DP_OP_424J2_126_3477_n2900,
         DP_OP_424J2_126_3477_n2899, DP_OP_424J2_126_3477_n2898,
         DP_OP_424J2_126_3477_n2897, DP_OP_424J2_126_3477_n2896,
         DP_OP_424J2_126_3477_n2895, DP_OP_424J2_126_3477_n2894,
         DP_OP_424J2_126_3477_n2893, DP_OP_424J2_126_3477_n2891,
         DP_OP_424J2_126_3477_n2890, DP_OP_424J2_126_3477_n2889,
         DP_OP_424J2_126_3477_n2887, DP_OP_424J2_126_3477_n2886,
         DP_OP_424J2_126_3477_n2883, DP_OP_424J2_126_3477_n2882,
         DP_OP_424J2_126_3477_n2881, DP_OP_424J2_126_3477_n2880,
         DP_OP_424J2_126_3477_n2879, DP_OP_424J2_126_3477_n2878,
         DP_OP_424J2_126_3477_n2877, DP_OP_424J2_126_3477_n2876,
         DP_OP_424J2_126_3477_n2875, DP_OP_424J2_126_3477_n2874,
         DP_OP_424J2_126_3477_n2873, DP_OP_424J2_126_3477_n2872,
         DP_OP_424J2_126_3477_n2871, DP_OP_424J2_126_3477_n2870,
         DP_OP_424J2_126_3477_n2869, DP_OP_424J2_126_3477_n2868,
         DP_OP_424J2_126_3477_n2867, DP_OP_424J2_126_3477_n2866,
         DP_OP_424J2_126_3477_n2865, DP_OP_424J2_126_3477_n2864,
         DP_OP_424J2_126_3477_n2863, DP_OP_424J2_126_3477_n2862,
         DP_OP_424J2_126_3477_n2861, DP_OP_424J2_126_3477_n2860,
         DP_OP_424J2_126_3477_n2859, DP_OP_424J2_126_3477_n2858,
         DP_OP_424J2_126_3477_n2857, DP_OP_424J2_126_3477_n2856,
         DP_OP_424J2_126_3477_n2854, DP_OP_424J2_126_3477_n2853,
         DP_OP_424J2_126_3477_n2852, DP_OP_424J2_126_3477_n2851,
         DP_OP_424J2_126_3477_n2850, DP_OP_424J2_126_3477_n2849,
         DP_OP_424J2_126_3477_n2846, DP_OP_424J2_126_3477_n2845,
         DP_OP_424J2_126_3477_n2837, DP_OP_424J2_126_3477_n2836,
         DP_OP_424J2_126_3477_n2835, DP_OP_424J2_126_3477_n2834,
         DP_OP_424J2_126_3477_n2833, DP_OP_424J2_126_3477_n2832,
         DP_OP_424J2_126_3477_n2831, DP_OP_424J2_126_3477_n2830,
         DP_OP_424J2_126_3477_n2829, DP_OP_424J2_126_3477_n2828,
         DP_OP_424J2_126_3477_n2827, DP_OP_424J2_126_3477_n2826,
         DP_OP_424J2_126_3477_n2825, DP_OP_424J2_126_3477_n2824,
         DP_OP_424J2_126_3477_n2823, DP_OP_424J2_126_3477_n2822,
         DP_OP_424J2_126_3477_n2821, DP_OP_424J2_126_3477_n2820,
         DP_OP_424J2_126_3477_n2819, DP_OP_424J2_126_3477_n2818,
         DP_OP_424J2_126_3477_n2817, DP_OP_424J2_126_3477_n2816,
         DP_OP_424J2_126_3477_n2815, DP_OP_424J2_126_3477_n2814,
         DP_OP_424J2_126_3477_n2813, DP_OP_424J2_126_3477_n2812,
         DP_OP_424J2_126_3477_n2811, DP_OP_424J2_126_3477_n2810,
         DP_OP_424J2_126_3477_n2809, DP_OP_424J2_126_3477_n2808,
         DP_OP_424J2_126_3477_n2807, DP_OP_424J2_126_3477_n2806,
         DP_OP_424J2_126_3477_n2805, DP_OP_424J2_126_3477_n2802,
         DP_OP_424J2_126_3477_n2801, DP_OP_424J2_126_3477_n2799,
         DP_OP_424J2_126_3477_n2796, DP_OP_424J2_126_3477_n2795,
         DP_OP_424J2_126_3477_n2794, DP_OP_424J2_126_3477_n2793,
         DP_OP_424J2_126_3477_n2792, DP_OP_424J2_126_3477_n2791,
         DP_OP_424J2_126_3477_n2790, DP_OP_424J2_126_3477_n2789,
         DP_OP_424J2_126_3477_n2788, DP_OP_424J2_126_3477_n2787,
         DP_OP_424J2_126_3477_n2786, DP_OP_424J2_126_3477_n2785,
         DP_OP_424J2_126_3477_n2784, DP_OP_424J2_126_3477_n2783,
         DP_OP_424J2_126_3477_n2782, DP_OP_424J2_126_3477_n2780,
         DP_OP_424J2_126_3477_n2779, DP_OP_424J2_126_3477_n2778,
         DP_OP_424J2_126_3477_n2777, DP_OP_424J2_126_3477_n2776,
         DP_OP_424J2_126_3477_n2775, DP_OP_424J2_126_3477_n2774,
         DP_OP_424J2_126_3477_n2773, DP_OP_424J2_126_3477_n2772,
         DP_OP_424J2_126_3477_n2771, DP_OP_424J2_126_3477_n2770,
         DP_OP_424J2_126_3477_n2769, DP_OP_424J2_126_3477_n2768,
         DP_OP_424J2_126_3477_n2767, DP_OP_424J2_126_3477_n2766,
         DP_OP_424J2_126_3477_n2765, DP_OP_424J2_126_3477_n2764,
         DP_OP_424J2_126_3477_n2763, DP_OP_424J2_126_3477_n2762,
         DP_OP_424J2_126_3477_n2758, DP_OP_424J2_126_3477_n2756,
         DP_OP_424J2_126_3477_n2754, DP_OP_424J2_126_3477_n2752,
         DP_OP_424J2_126_3477_n2749, DP_OP_424J2_126_3477_n2748,
         DP_OP_424J2_126_3477_n2747, DP_OP_424J2_126_3477_n2746,
         DP_OP_424J2_126_3477_n2745, DP_OP_424J2_126_3477_n2744,
         DP_OP_424J2_126_3477_n2743, DP_OP_424J2_126_3477_n2742,
         DP_OP_424J2_126_3477_n2741, DP_OP_424J2_126_3477_n2740,
         DP_OP_424J2_126_3477_n2739, DP_OP_424J2_126_3477_n2738,
         DP_OP_424J2_126_3477_n2737, DP_OP_424J2_126_3477_n2736,
         DP_OP_424J2_126_3477_n2735, DP_OP_424J2_126_3477_n2734,
         DP_OP_424J2_126_3477_n2733, DP_OP_424J2_126_3477_n2732,
         DP_OP_424J2_126_3477_n2731, DP_OP_424J2_126_3477_n2730,
         DP_OP_424J2_126_3477_n2729, DP_OP_424J2_126_3477_n2728,
         DP_OP_424J2_126_3477_n2727, DP_OP_424J2_126_3477_n2726,
         DP_OP_424J2_126_3477_n2725, DP_OP_424J2_126_3477_n2724,
         DP_OP_424J2_126_3477_n2723, DP_OP_424J2_126_3477_n2722,
         DP_OP_424J2_126_3477_n2721, DP_OP_424J2_126_3477_n2720,
         DP_OP_424J2_126_3477_n2719, DP_OP_424J2_126_3477_n2718,
         DP_OP_424J2_126_3477_n2716, DP_OP_424J2_126_3477_n2712,
         DP_OP_424J2_126_3477_n2705, DP_OP_424J2_126_3477_n2704,
         DP_OP_424J2_126_3477_n2703, DP_OP_424J2_126_3477_n2702,
         DP_OP_424J2_126_3477_n2701, DP_OP_424J2_126_3477_n2700,
         DP_OP_424J2_126_3477_n2699, DP_OP_424J2_126_3477_n2698,
         DP_OP_424J2_126_3477_n2697, DP_OP_424J2_126_3477_n2696,
         DP_OP_424J2_126_3477_n2695, DP_OP_424J2_126_3477_n2694,
         DP_OP_424J2_126_3477_n2693, DP_OP_424J2_126_3477_n2692,
         DP_OP_424J2_126_3477_n2691, DP_OP_424J2_126_3477_n2690,
         DP_OP_424J2_126_3477_n2689, DP_OP_424J2_126_3477_n2688,
         DP_OP_424J2_126_3477_n2687, DP_OP_424J2_126_3477_n2686,
         DP_OP_424J2_126_3477_n2685, DP_OP_424J2_126_3477_n2684,
         DP_OP_424J2_126_3477_n2683, DP_OP_424J2_126_3477_n2682,
         DP_OP_424J2_126_3477_n2681, DP_OP_424J2_126_3477_n2680,
         DP_OP_424J2_126_3477_n2679, DP_OP_424J2_126_3477_n2678,
         DP_OP_424J2_126_3477_n2677, DP_OP_424J2_126_3477_n2676,
         DP_OP_424J2_126_3477_n2675, DP_OP_424J2_126_3477_n2674,
         DP_OP_424J2_126_3477_n2673, DP_OP_424J2_126_3477_n2671,
         DP_OP_424J2_126_3477_n2669, DP_OP_424J2_126_3477_n2667,
         DP_OP_424J2_126_3477_n2661, DP_OP_424J2_126_3477_n2660,
         DP_OP_424J2_126_3477_n2659, DP_OP_424J2_126_3477_n2658,
         DP_OP_424J2_126_3477_n2657, DP_OP_424J2_126_3477_n2656,
         DP_OP_424J2_126_3477_n2655, DP_OP_424J2_126_3477_n2654,
         DP_OP_424J2_126_3477_n2653, DP_OP_424J2_126_3477_n2652,
         DP_OP_424J2_126_3477_n2651, DP_OP_424J2_126_3477_n2650,
         DP_OP_424J2_126_3477_n2649, DP_OP_424J2_126_3477_n2648,
         DP_OP_424J2_126_3477_n2647, DP_OP_424J2_126_3477_n2646,
         DP_OP_424J2_126_3477_n2645, DP_OP_424J2_126_3477_n2644,
         DP_OP_424J2_126_3477_n2643, DP_OP_424J2_126_3477_n2642,
         DP_OP_424J2_126_3477_n2641, DP_OP_424J2_126_3477_n2640,
         DP_OP_424J2_126_3477_n2639, DP_OP_424J2_126_3477_n2638,
         DP_OP_424J2_126_3477_n2637, DP_OP_424J2_126_3477_n2636,
         DP_OP_424J2_126_3477_n2635, DP_OP_424J2_126_3477_n2634,
         DP_OP_424J2_126_3477_n2633, DP_OP_424J2_126_3477_n2632,
         DP_OP_424J2_126_3477_n2631, DP_OP_424J2_126_3477_n2630,
         DP_OP_424J2_126_3477_n2629, DP_OP_424J2_126_3477_n2627,
         DP_OP_424J2_126_3477_n2623, DP_OP_424J2_126_3477_n2622,
         DP_OP_424J2_126_3477_n2619, DP_OP_424J2_126_3477_n2617,
         DP_OP_424J2_126_3477_n2616, DP_OP_424J2_126_3477_n2615,
         DP_OP_424J2_126_3477_n2614, DP_OP_424J2_126_3477_n2613,
         DP_OP_424J2_126_3477_n2612, DP_OP_424J2_126_3477_n2611,
         DP_OP_424J2_126_3477_n2610, DP_OP_424J2_126_3477_n2609,
         DP_OP_424J2_126_3477_n2608, DP_OP_424J2_126_3477_n2607,
         DP_OP_424J2_126_3477_n2606, DP_OP_424J2_126_3477_n2605,
         DP_OP_424J2_126_3477_n2604, DP_OP_424J2_126_3477_n2603,
         DP_OP_424J2_126_3477_n2602, DP_OP_424J2_126_3477_n2601,
         DP_OP_424J2_126_3477_n2600, DP_OP_424J2_126_3477_n2599,
         DP_OP_424J2_126_3477_n2598, DP_OP_424J2_126_3477_n2597,
         DP_OP_424J2_126_3477_n2596, DP_OP_424J2_126_3477_n2595,
         DP_OP_424J2_126_3477_n2594, DP_OP_424J2_126_3477_n2593,
         DP_OP_424J2_126_3477_n2592, DP_OP_424J2_126_3477_n2591,
         DP_OP_424J2_126_3477_n2590, DP_OP_424J2_126_3477_n2589,
         DP_OP_424J2_126_3477_n2588, DP_OP_424J2_126_3477_n2587,
         DP_OP_424J2_126_3477_n2586, DP_OP_424J2_126_3477_n2585,
         DP_OP_424J2_126_3477_n2584, DP_OP_424J2_126_3477_n2582,
         DP_OP_424J2_126_3477_n2580, DP_OP_424J2_126_3477_n2579,
         DP_OP_424J2_126_3477_n2576, DP_OP_424J2_126_3477_n2575,
         DP_OP_424J2_126_3477_n2574, DP_OP_424J2_126_3477_n2573,
         DP_OP_424J2_126_3477_n2572, DP_OP_424J2_126_3477_n2571,
         DP_OP_424J2_126_3477_n2569, DP_OP_424J2_126_3477_n2568,
         DP_OP_424J2_126_3477_n2567, DP_OP_424J2_126_3477_n2566,
         DP_OP_424J2_126_3477_n2565, DP_OP_424J2_126_3477_n2564,
         DP_OP_424J2_126_3477_n2563, DP_OP_424J2_126_3477_n2562,
         DP_OP_424J2_126_3477_n2561, DP_OP_424J2_126_3477_n2560,
         DP_OP_424J2_126_3477_n2559, DP_OP_424J2_126_3477_n2558,
         DP_OP_424J2_126_3477_n2557, DP_OP_424J2_126_3477_n2556,
         DP_OP_424J2_126_3477_n2555, DP_OP_424J2_126_3477_n2554,
         DP_OP_424J2_126_3477_n2553, DP_OP_424J2_126_3477_n2552,
         DP_OP_424J2_126_3477_n2551, DP_OP_424J2_126_3477_n2550,
         DP_OP_424J2_126_3477_n2549, DP_OP_424J2_126_3477_n2548,
         DP_OP_424J2_126_3477_n2547, DP_OP_424J2_126_3477_n2546,
         DP_OP_424J2_126_3477_n2545, DP_OP_424J2_126_3477_n2544,
         DP_OP_424J2_126_3477_n2543, DP_OP_424J2_126_3477_n2542,
         DP_OP_424J2_126_3477_n2541, DP_OP_424J2_126_3477_n2540,
         DP_OP_424J2_126_3477_n2535, DP_OP_424J2_126_3477_n2534,
         DP_OP_424J2_126_3477_n2532, DP_OP_424J2_126_3477_n2529,
         DP_OP_424J2_126_3477_n2528, DP_OP_424J2_126_3477_n2527,
         DP_OP_424J2_126_3477_n2526, DP_OP_424J2_126_3477_n2525,
         DP_OP_424J2_126_3477_n2524, DP_OP_424J2_126_3477_n2523,
         DP_OP_424J2_126_3477_n2522, DP_OP_424J2_126_3477_n2521,
         DP_OP_424J2_126_3477_n2520, DP_OP_424J2_126_3477_n2519,
         DP_OP_424J2_126_3477_n2518, DP_OP_424J2_126_3477_n2517,
         DP_OP_424J2_126_3477_n2516, DP_OP_424J2_126_3477_n2515,
         DP_OP_424J2_126_3477_n2514, DP_OP_424J2_126_3477_n2513,
         DP_OP_424J2_126_3477_n2512, DP_OP_424J2_126_3477_n2511,
         DP_OP_424J2_126_3477_n2510, DP_OP_424J2_126_3477_n2509,
         DP_OP_424J2_126_3477_n2508, DP_OP_424J2_126_3477_n2507,
         DP_OP_424J2_126_3477_n2506, DP_OP_424J2_126_3477_n2505,
         DP_OP_424J2_126_3477_n2504, DP_OP_424J2_126_3477_n2503,
         DP_OP_424J2_126_3477_n2502, DP_OP_424J2_126_3477_n2501,
         DP_OP_424J2_126_3477_n2500, DP_OP_424J2_126_3477_n2499,
         DP_OP_424J2_126_3477_n2498, DP_OP_424J2_126_3477_n2497,
         DP_OP_424J2_126_3477_n2491, DP_OP_424J2_126_3477_n2486,
         DP_OP_424J2_126_3477_n2485, DP_OP_424J2_126_3477_n2484,
         DP_OP_424J2_126_3477_n2483, DP_OP_424J2_126_3477_n2482,
         DP_OP_424J2_126_3477_n2481, DP_OP_424J2_126_3477_n2480,
         DP_OP_424J2_126_3477_n2479, DP_OP_424J2_126_3477_n2478,
         DP_OP_424J2_126_3477_n2477, DP_OP_424J2_126_3477_n2476,
         DP_OP_424J2_126_3477_n2475, DP_OP_424J2_126_3477_n2474,
         DP_OP_424J2_126_3477_n2473, DP_OP_424J2_126_3477_n2472,
         DP_OP_424J2_126_3477_n2471, DP_OP_424J2_126_3477_n2470,
         DP_OP_424J2_126_3477_n2469, DP_OP_424J2_126_3477_n2468,
         DP_OP_424J2_126_3477_n2467, DP_OP_424J2_126_3477_n2466,
         DP_OP_424J2_126_3477_n2465, DP_OP_424J2_126_3477_n2464,
         DP_OP_424J2_126_3477_n2463, DP_OP_424J2_126_3477_n2462,
         DP_OP_424J2_126_3477_n2461, DP_OP_424J2_126_3477_n2460,
         DP_OP_424J2_126_3477_n2459, DP_OP_424J2_126_3477_n2458,
         DP_OP_424J2_126_3477_n2457, DP_OP_424J2_126_3477_n2456,
         DP_OP_424J2_126_3477_n2455, DP_OP_424J2_126_3477_n2454,
         DP_OP_424J2_126_3477_n2447, DP_OP_424J2_126_3477_n2443,
         DP_OP_424J2_126_3477_n2441, DP_OP_424J2_126_3477_n2440,
         DP_OP_424J2_126_3477_n2439, DP_OP_424J2_126_3477_n2438,
         DP_OP_424J2_126_3477_n2437, DP_OP_424J2_126_3477_n2436,
         DP_OP_424J2_126_3477_n2435, DP_OP_424J2_126_3477_n2434,
         DP_OP_424J2_126_3477_n2433, DP_OP_424J2_126_3477_n2432,
         DP_OP_424J2_126_3477_n2431, DP_OP_424J2_126_3477_n2430,
         DP_OP_424J2_126_3477_n2429, DP_OP_424J2_126_3477_n2428,
         DP_OP_424J2_126_3477_n2427, DP_OP_424J2_126_3477_n2426,
         DP_OP_424J2_126_3477_n2425, DP_OP_424J2_126_3477_n2424,
         DP_OP_424J2_126_3477_n2423, DP_OP_424J2_126_3477_n2422,
         DP_OP_424J2_126_3477_n2421, DP_OP_424J2_126_3477_n2420,
         DP_OP_424J2_126_3477_n2419, DP_OP_424J2_126_3477_n2418,
         DP_OP_424J2_126_3477_n2417, DP_OP_424J2_126_3477_n2416,
         DP_OP_424J2_126_3477_n2415, DP_OP_424J2_126_3477_n2414,
         DP_OP_424J2_126_3477_n2413, DP_OP_424J2_126_3477_n2412,
         DP_OP_424J2_126_3477_n2411, DP_OP_424J2_126_3477_n2410,
         DP_OP_424J2_126_3477_n2409, DP_OP_424J2_126_3477_n2408,
         DP_OP_424J2_126_3477_n2405, DP_OP_424J2_126_3477_n2403,
         DP_OP_424J2_126_3477_n2400, DP_OP_424J2_126_3477_n2397,
         DP_OP_424J2_126_3477_n2396, DP_OP_424J2_126_3477_n2395,
         DP_OP_424J2_126_3477_n2394, DP_OP_424J2_126_3477_n2393,
         DP_OP_424J2_126_3477_n2392, DP_OP_424J2_126_3477_n2391,
         DP_OP_424J2_126_3477_n2390, DP_OP_424J2_126_3477_n2389,
         DP_OP_424J2_126_3477_n2388, DP_OP_424J2_126_3477_n2387,
         DP_OP_424J2_126_3477_n2386, DP_OP_424J2_126_3477_n2385,
         DP_OP_424J2_126_3477_n2384, DP_OP_424J2_126_3477_n2383,
         DP_OP_424J2_126_3477_n2382, DP_OP_424J2_126_3477_n2381,
         DP_OP_424J2_126_3477_n2380, DP_OP_424J2_126_3477_n2379,
         DP_OP_424J2_126_3477_n2378, DP_OP_424J2_126_3477_n2377,
         DP_OP_424J2_126_3477_n2376, DP_OP_424J2_126_3477_n2375,
         DP_OP_424J2_126_3477_n2374, DP_OP_424J2_126_3477_n2373,
         DP_OP_424J2_126_3477_n2372, DP_OP_424J2_126_3477_n2371,
         DP_OP_424J2_126_3477_n2370, DP_OP_424J2_126_3477_n2369,
         DP_OP_424J2_126_3477_n2368, DP_OP_424J2_126_3477_n2367,
         DP_OP_424J2_126_3477_n2366, DP_OP_424J2_126_3477_n2365,
         DP_OP_424J2_126_3477_n2358, DP_OP_424J2_126_3477_n2354,
         DP_OP_424J2_126_3477_n2353, DP_OP_424J2_126_3477_n2352,
         DP_OP_424J2_126_3477_n2351, DP_OP_424J2_126_3477_n2350,
         DP_OP_424J2_126_3477_n2349, DP_OP_424J2_126_3477_n2348,
         DP_OP_424J2_126_3477_n2347, DP_OP_424J2_126_3477_n2346,
         DP_OP_424J2_126_3477_n2345, DP_OP_424J2_126_3477_n2344,
         DP_OP_424J2_126_3477_n2343, DP_OP_424J2_126_3477_n2342,
         DP_OP_424J2_126_3477_n2340, DP_OP_424J2_126_3477_n2339,
         DP_OP_424J2_126_3477_n2338, DP_OP_424J2_126_3477_n2337,
         DP_OP_424J2_126_3477_n2336, DP_OP_424J2_126_3477_n2335,
         DP_OP_424J2_126_3477_n2334, DP_OP_424J2_126_3477_n2333,
         DP_OP_424J2_126_3477_n2332, DP_OP_424J2_126_3477_n2331,
         DP_OP_424J2_126_3477_n2330, DP_OP_424J2_126_3477_n2329,
         DP_OP_424J2_126_3477_n2328, DP_OP_424J2_126_3477_n2327,
         DP_OP_424J2_126_3477_n2326, DP_OP_424J2_126_3477_n2325,
         DP_OP_424J2_126_3477_n2324, DP_OP_424J2_126_3477_n2323,
         DP_OP_424J2_126_3477_n2322, DP_OP_424J2_126_3477_n2318,
         DP_OP_424J2_126_3477_n2317, DP_OP_424J2_126_3477_n2315,
         DP_OP_424J2_126_3477_n2311, DP_OP_424J2_126_3477_n2309,
         DP_OP_424J2_126_3477_n2308, DP_OP_424J2_126_3477_n2307,
         DP_OP_424J2_126_3477_n2306, DP_OP_424J2_126_3477_n2305,
         DP_OP_424J2_126_3477_n2304, DP_OP_424J2_126_3477_n2303,
         DP_OP_424J2_126_3477_n2302, DP_OP_424J2_126_3477_n2301,
         DP_OP_424J2_126_3477_n2300, DP_OP_424J2_126_3477_n2299,
         DP_OP_424J2_126_3477_n2298, DP_OP_424J2_126_3477_n2297,
         DP_OP_424J2_126_3477_n2296, DP_OP_424J2_126_3477_n2295,
         DP_OP_424J2_126_3477_n2294, DP_OP_424J2_126_3477_n2293,
         DP_OP_424J2_126_3477_n2292, DP_OP_424J2_126_3477_n2291,
         DP_OP_424J2_126_3477_n2289, DP_OP_424J2_126_3477_n2288,
         DP_OP_424J2_126_3477_n2287, DP_OP_424J2_126_3477_n2286,
         DP_OP_424J2_126_3477_n2285, DP_OP_424J2_126_3477_n2284,
         DP_OP_424J2_126_3477_n2283, DP_OP_424J2_126_3477_n2282,
         DP_OP_424J2_126_3477_n2281, DP_OP_424J2_126_3477_n2280,
         DP_OP_424J2_126_3477_n2279, DP_OP_424J2_126_3477_n2278,
         DP_OP_424J2_126_3477_n2277, DP_OP_424J2_126_3477_n2276,
         DP_OP_424J2_126_3477_n2275, DP_OP_424J2_126_3477_n2274,
         DP_OP_424J2_126_3477_n2269, DP_OP_424J2_126_3477_n2268,
         DP_OP_424J2_126_3477_n2267, DP_OP_424J2_126_3477_n2265,
         DP_OP_424J2_126_3477_n2264, DP_OP_424J2_126_3477_n2263,
         DP_OP_424J2_126_3477_n2262, DP_OP_424J2_126_3477_n2261,
         DP_OP_424J2_126_3477_n2259, DP_OP_424J2_126_3477_n2258,
         DP_OP_424J2_126_3477_n2257, DP_OP_424J2_126_3477_n2256,
         DP_OP_424J2_126_3477_n2255, DP_OP_424J2_126_3477_n2254,
         DP_OP_424J2_126_3477_n2253, DP_OP_424J2_126_3477_n2252,
         DP_OP_424J2_126_3477_n2251, DP_OP_424J2_126_3477_n2250,
         DP_OP_424J2_126_3477_n2249, DP_OP_424J2_126_3477_n2248,
         DP_OP_424J2_126_3477_n2247, DP_OP_424J2_126_3477_n2246,
         DP_OP_424J2_126_3477_n2245, DP_OP_424J2_126_3477_n2244,
         DP_OP_424J2_126_3477_n2243, DP_OP_424J2_126_3477_n2242,
         DP_OP_424J2_126_3477_n2241, DP_OP_424J2_126_3477_n2240,
         DP_OP_424J2_126_3477_n2239, DP_OP_424J2_126_3477_n2238,
         DP_OP_424J2_126_3477_n2237, DP_OP_424J2_126_3477_n2236,
         DP_OP_424J2_126_3477_n2235, DP_OP_424J2_126_3477_n2234,
         DP_OP_424J2_126_3477_n2231, DP_OP_424J2_126_3477_n2222,
         DP_OP_424J2_126_3477_n2221, DP_OP_424J2_126_3477_n2220,
         DP_OP_424J2_126_3477_n2219, DP_OP_424J2_126_3477_n2218,
         DP_OP_424J2_126_3477_n2217, DP_OP_424J2_126_3477_n2216,
         DP_OP_424J2_126_3477_n2215, DP_OP_424J2_126_3477_n2214,
         DP_OP_424J2_126_3477_n2213, DP_OP_424J2_126_3477_n2212,
         DP_OP_424J2_126_3477_n2211, DP_OP_424J2_126_3477_n2210,
         DP_OP_424J2_126_3477_n2209, DP_OP_424J2_126_3477_n2208,
         DP_OP_424J2_126_3477_n2207, DP_OP_424J2_126_3477_n2206,
         DP_OP_424J2_126_3477_n2205, DP_OP_424J2_126_3477_n2204,
         DP_OP_424J2_126_3477_n2203, DP_OP_424J2_126_3477_n2202,
         DP_OP_424J2_126_3477_n2201, DP_OP_424J2_126_3477_n2200,
         DP_OP_424J2_126_3477_n2199, DP_OP_424J2_126_3477_n2198,
         DP_OP_424J2_126_3477_n2197, DP_OP_424J2_126_3477_n2196,
         DP_OP_424J2_126_3477_n2195, DP_OP_424J2_126_3477_n2194,
         DP_OP_424J2_126_3477_n2193, DP_OP_424J2_126_3477_n2192,
         DP_OP_424J2_126_3477_n2191, DP_OP_424J2_126_3477_n2190,
         DP_OP_424J2_126_3477_n2189, DP_OP_424J2_126_3477_n2186,
         DP_OP_424J2_126_3477_n2185, DP_OP_424J2_126_3477_n2184,
         DP_OP_424J2_126_3477_n2177, DP_OP_424J2_126_3477_n2176,
         DP_OP_424J2_126_3477_n2175, DP_OP_424J2_126_3477_n2174,
         DP_OP_424J2_126_3477_n2173, DP_OP_424J2_126_3477_n2172,
         DP_OP_424J2_126_3477_n2171, DP_OP_424J2_126_3477_n2170,
         DP_OP_424J2_126_3477_n2169, DP_OP_424J2_126_3477_n2168,
         DP_OP_424J2_126_3477_n2167, DP_OP_424J2_126_3477_n2166,
         DP_OP_424J2_126_3477_n2165, DP_OP_424J2_126_3477_n2164,
         DP_OP_424J2_126_3477_n2163, DP_OP_424J2_126_3477_n2162,
         DP_OP_424J2_126_3477_n2161, DP_OP_424J2_126_3477_n2160,
         DP_OP_424J2_126_3477_n2159, DP_OP_424J2_126_3477_n2158,
         DP_OP_424J2_126_3477_n2157, DP_OP_424J2_126_3477_n2156,
         DP_OP_424J2_126_3477_n2155, DP_OP_424J2_126_3477_n2154,
         DP_OP_424J2_126_3477_n2153, DP_OP_424J2_126_3477_n2152,
         DP_OP_424J2_126_3477_n2151, DP_OP_424J2_126_3477_n2150,
         DP_OP_424J2_126_3477_n2149, DP_OP_424J2_126_3477_n2148,
         DP_OP_424J2_126_3477_n2147, DP_OP_424J2_126_3477_n2146,
         DP_OP_424J2_126_3477_n2144, DP_OP_424J2_126_3477_n2143,
         DP_OP_424J2_126_3477_n2138, DP_OP_424J2_126_3477_n2136,
         DP_OP_424J2_126_3477_n2133, DP_OP_424J2_126_3477_n2132,
         DP_OP_424J2_126_3477_n2131, DP_OP_424J2_126_3477_n2130,
         DP_OP_424J2_126_3477_n2129, DP_OP_424J2_126_3477_n2128,
         DP_OP_424J2_126_3477_n2127, DP_OP_424J2_126_3477_n2126,
         DP_OP_424J2_126_3477_n2125, DP_OP_424J2_126_3477_n2124,
         DP_OP_424J2_126_3477_n2123, DP_OP_424J2_126_3477_n2122,
         DP_OP_424J2_126_3477_n2121, DP_OP_424J2_126_3477_n2120,
         DP_OP_424J2_126_3477_n2119, DP_OP_424J2_126_3477_n2118,
         DP_OP_424J2_126_3477_n2117, DP_OP_424J2_126_3477_n2116,
         DP_OP_424J2_126_3477_n2115, DP_OP_424J2_126_3477_n2114,
         DP_OP_424J2_126_3477_n2113, DP_OP_424J2_126_3477_n2112,
         DP_OP_424J2_126_3477_n2111, DP_OP_424J2_126_3477_n2110,
         DP_OP_424J2_126_3477_n2109, DP_OP_424J2_126_3477_n2108,
         DP_OP_424J2_126_3477_n2106, DP_OP_424J2_126_3477_n2105,
         DP_OP_424J2_126_3477_n2104, DP_OP_424J2_126_3477_n2103,
         DP_OP_424J2_126_3477_n2102, DP_OP_424J2_126_3477_n2100,
         DP_OP_424J2_126_3477_n2099, DP_OP_424J2_126_3477_n2095,
         DP_OP_424J2_126_3477_n2092, DP_OP_424J2_126_3477_n2090,
         DP_OP_424J2_126_3477_n2089, DP_OP_424J2_126_3477_n2088,
         DP_OP_424J2_126_3477_n2087, DP_OP_424J2_126_3477_n2086,
         DP_OP_424J2_126_3477_n2085, DP_OP_424J2_126_3477_n2084,
         DP_OP_424J2_126_3477_n2083, DP_OP_424J2_126_3477_n2082,
         DP_OP_424J2_126_3477_n2081, DP_OP_424J2_126_3477_n2080,
         DP_OP_424J2_126_3477_n2079, DP_OP_424J2_126_3477_n2078,
         DP_OP_424J2_126_3477_n2077, DP_OP_424J2_126_3477_n2076,
         DP_OP_424J2_126_3477_n2075, DP_OP_424J2_126_3477_n2074,
         DP_OP_424J2_126_3477_n2073, DP_OP_424J2_126_3477_n2072,
         DP_OP_424J2_126_3477_n2071, DP_OP_424J2_126_3477_n2070,
         DP_OP_424J2_126_3477_n2069, DP_OP_424J2_126_3477_n2068,
         DP_OP_424J2_126_3477_n2067, DP_OP_424J2_126_3477_n2066,
         DP_OP_424J2_126_3477_n2065, DP_OP_424J2_126_3477_n2064,
         DP_OP_424J2_126_3477_n2063, DP_OP_424J2_126_3477_n2062,
         DP_OP_424J2_126_3477_n2061, DP_OP_424J2_126_3477_n2060,
         DP_OP_424J2_126_3477_n2059, DP_OP_424J2_126_3477_n2058,
         DP_OP_424J2_126_3477_n2057, DP_OP_424J2_126_3477_n2056,
         DP_OP_424J2_126_3477_n2055, DP_OP_424J2_126_3477_n2051,
         DP_OP_424J2_126_3477_n2045, DP_OP_424J2_126_3477_n2044,
         DP_OP_424J2_126_3477_n2043, DP_OP_424J2_126_3477_n2042,
         DP_OP_424J2_126_3477_n2041, DP_OP_424J2_126_3477_n2040,
         DP_OP_424J2_126_3477_n2039, DP_OP_424J2_126_3477_n2038,
         DP_OP_424J2_126_3477_n2037, DP_OP_424J2_126_3477_n2036,
         DP_OP_424J2_126_3477_n2035, DP_OP_424J2_126_3477_n2034,
         DP_OP_424J2_126_3477_n2033, DP_OP_424J2_126_3477_n2032,
         DP_OP_424J2_126_3477_n2031, DP_OP_424J2_126_3477_n2030,
         DP_OP_424J2_126_3477_n2029, DP_OP_424J2_126_3477_n2028,
         DP_OP_424J2_126_3477_n2027, DP_OP_424J2_126_3477_n2026,
         DP_OP_424J2_126_3477_n2025, DP_OP_424J2_126_3477_n2024,
         DP_OP_424J2_126_3477_n2023, DP_OP_424J2_126_3477_n2022,
         DP_OP_424J2_126_3477_n2021, DP_OP_424J2_126_3477_n2020,
         DP_OP_424J2_126_3477_n2019, DP_OP_424J2_126_3477_n2018,
         DP_OP_424J2_126_3477_n2017, DP_OP_424J2_126_3477_n2016,
         DP_OP_424J2_126_3477_n2015, DP_OP_424J2_126_3477_n2014,
         DP_OP_424J2_126_3477_n2011, DP_OP_424J2_126_3477_n2010,
         DP_OP_424J2_126_3477_n2006, DP_OP_424J2_126_3477_n2005,
         DP_OP_424J2_126_3477_n2004, DP_OP_424J2_126_3477_n2003,
         DP_OP_424J2_126_3477_n2002, DP_OP_424J2_126_3477_n2001,
         DP_OP_424J2_126_3477_n2000, DP_OP_424J2_126_3477_n1999,
         DP_OP_424J2_126_3477_n1998, DP_OP_424J2_126_3477_n1997,
         DP_OP_424J2_126_3477_n1996, DP_OP_424J2_126_3477_n1995,
         DP_OP_424J2_126_3477_n1994, DP_OP_424J2_126_3477_n1993,
         DP_OP_424J2_126_3477_n1992, DP_OP_424J2_126_3477_n1991,
         DP_OP_424J2_126_3477_n1990, DP_OP_424J2_126_3477_n1989,
         DP_OP_424J2_126_3477_n1988, DP_OP_424J2_126_3477_n1987,
         DP_OP_424J2_126_3477_n1986, DP_OP_424J2_126_3477_n1985,
         DP_OP_424J2_126_3477_n1984, DP_OP_424J2_126_3477_n1983,
         DP_OP_424J2_126_3477_n1982, DP_OP_424J2_126_3477_n1981,
         DP_OP_424J2_126_3477_n1980, DP_OP_424J2_126_3477_n1979,
         DP_OP_424J2_126_3477_n1978, DP_OP_424J2_126_3477_n1977,
         DP_OP_424J2_126_3477_n1976, DP_OP_424J2_126_3477_n1975,
         DP_OP_424J2_126_3477_n1974, DP_OP_424J2_126_3477_n1973,
         DP_OP_424J2_126_3477_n1972, DP_OP_424J2_126_3477_n1971,
         DP_OP_424J2_126_3477_n1970, DP_OP_424J2_126_3477_n1936,
         DP_OP_424J2_126_3477_n1935, DP_OP_424J2_126_3477_n1934,
         DP_OP_424J2_126_3477_n1933, DP_OP_424J2_126_3477_n1932,
         DP_OP_424J2_126_3477_n1931, DP_OP_424J2_126_3477_n1930,
         DP_OP_424J2_126_3477_n1929, DP_OP_424J2_126_3477_n1928,
         DP_OP_424J2_126_3477_n1927, DP_OP_424J2_126_3477_n1926,
         DP_OP_424J2_126_3477_n1925, DP_OP_424J2_126_3477_n1924,
         DP_OP_424J2_126_3477_n1923, DP_OP_424J2_126_3477_n1921,
         DP_OP_424J2_126_3477_n1920, DP_OP_424J2_126_3477_n1919,
         DP_OP_424J2_126_3477_n1918, DP_OP_424J2_126_3477_n1917,
         DP_OP_424J2_126_3477_n1916, DP_OP_424J2_126_3477_n1915,
         DP_OP_424J2_126_3477_n1914, DP_OP_424J2_126_3477_n1913,
         DP_OP_424J2_126_3477_n1912, DP_OP_424J2_126_3477_n1911,
         DP_OP_424J2_126_3477_n1910, DP_OP_424J2_126_3477_n1909,
         DP_OP_424J2_126_3477_n1908, DP_OP_424J2_126_3477_n1907,
         DP_OP_424J2_126_3477_n1906, DP_OP_424J2_126_3477_n1905,
         DP_OP_424J2_126_3477_n1904, DP_OP_424J2_126_3477_n1903,
         DP_OP_424J2_126_3477_n1902, DP_OP_424J2_126_3477_n1901,
         DP_OP_424J2_126_3477_n1900, DP_OP_424J2_126_3477_n1899,
         DP_OP_424J2_126_3477_n1898, DP_OP_424J2_126_3477_n1897,
         DP_OP_424J2_126_3477_n1896, DP_OP_424J2_126_3477_n1895,
         DP_OP_424J2_126_3477_n1894, DP_OP_424J2_126_3477_n1893,
         DP_OP_424J2_126_3477_n1892, DP_OP_424J2_126_3477_n1891,
         DP_OP_424J2_126_3477_n1890, DP_OP_424J2_126_3477_n1889,
         DP_OP_424J2_126_3477_n1888, DP_OP_424J2_126_3477_n1887,
         DP_OP_424J2_126_3477_n1886, DP_OP_424J2_126_3477_n1885,
         DP_OP_424J2_126_3477_n1884, DP_OP_424J2_126_3477_n1883,
         DP_OP_424J2_126_3477_n1882, DP_OP_424J2_126_3477_n1881,
         DP_OP_424J2_126_3477_n1880, DP_OP_424J2_126_3477_n1879,
         DP_OP_424J2_126_3477_n1878, DP_OP_424J2_126_3477_n1877,
         DP_OP_424J2_126_3477_n1876, DP_OP_424J2_126_3477_n1875,
         DP_OP_424J2_126_3477_n1874, DP_OP_424J2_126_3477_n1873,
         DP_OP_424J2_126_3477_n1872, DP_OP_424J2_126_3477_n1871,
         DP_OP_424J2_126_3477_n1870, DP_OP_424J2_126_3477_n1869,
         DP_OP_424J2_126_3477_n1868, DP_OP_424J2_126_3477_n1867,
         DP_OP_424J2_126_3477_n1866, DP_OP_424J2_126_3477_n1865,
         DP_OP_424J2_126_3477_n1864, DP_OP_424J2_126_3477_n1863,
         DP_OP_424J2_126_3477_n1862, DP_OP_424J2_126_3477_n1861,
         DP_OP_424J2_126_3477_n1860, DP_OP_424J2_126_3477_n1859,
         DP_OP_424J2_126_3477_n1858, DP_OP_424J2_126_3477_n1857,
         DP_OP_424J2_126_3477_n1856, DP_OP_424J2_126_3477_n1855,
         DP_OP_424J2_126_3477_n1854, DP_OP_424J2_126_3477_n1853,
         DP_OP_424J2_126_3477_n1852, DP_OP_424J2_126_3477_n1851,
         DP_OP_424J2_126_3477_n1850, DP_OP_424J2_126_3477_n1849,
         DP_OP_424J2_126_3477_n1848, DP_OP_424J2_126_3477_n1847,
         DP_OP_424J2_126_3477_n1846, DP_OP_424J2_126_3477_n1845,
         DP_OP_424J2_126_3477_n1844, DP_OP_424J2_126_3477_n1843,
         DP_OP_424J2_126_3477_n1842, DP_OP_424J2_126_3477_n1841,
         DP_OP_424J2_126_3477_n1840, DP_OP_424J2_126_3477_n1839,
         DP_OP_424J2_126_3477_n1838, DP_OP_424J2_126_3477_n1837,
         DP_OP_424J2_126_3477_n1836, DP_OP_424J2_126_3477_n1835,
         DP_OP_424J2_126_3477_n1834, DP_OP_424J2_126_3477_n1833,
         DP_OP_424J2_126_3477_n1832, DP_OP_424J2_126_3477_n1831,
         DP_OP_424J2_126_3477_n1830, DP_OP_424J2_126_3477_n1829,
         DP_OP_424J2_126_3477_n1828, DP_OP_424J2_126_3477_n1827,
         DP_OP_424J2_126_3477_n1826, DP_OP_424J2_126_3477_n1825,
         DP_OP_424J2_126_3477_n1824, DP_OP_424J2_126_3477_n1823,
         DP_OP_424J2_126_3477_n1822, DP_OP_424J2_126_3477_n1821,
         DP_OP_424J2_126_3477_n1820, DP_OP_424J2_126_3477_n1819,
         DP_OP_424J2_126_3477_n1818, DP_OP_424J2_126_3477_n1817,
         DP_OP_424J2_126_3477_n1816, DP_OP_424J2_126_3477_n1815,
         DP_OP_424J2_126_3477_n1814, DP_OP_424J2_126_3477_n1813,
         DP_OP_424J2_126_3477_n1812, DP_OP_424J2_126_3477_n1811,
         DP_OP_424J2_126_3477_n1810, DP_OP_424J2_126_3477_n1809,
         DP_OP_424J2_126_3477_n1808, DP_OP_424J2_126_3477_n1807,
         DP_OP_424J2_126_3477_n1806, DP_OP_424J2_126_3477_n1805,
         DP_OP_424J2_126_3477_n1804, DP_OP_424J2_126_3477_n1803,
         DP_OP_424J2_126_3477_n1802, DP_OP_424J2_126_3477_n1801,
         DP_OP_424J2_126_3477_n1800, DP_OP_424J2_126_3477_n1799,
         DP_OP_424J2_126_3477_n1798, DP_OP_424J2_126_3477_n1797,
         DP_OP_424J2_126_3477_n1796, DP_OP_424J2_126_3477_n1795,
         DP_OP_424J2_126_3477_n1794, DP_OP_424J2_126_3477_n1793,
         DP_OP_424J2_126_3477_n1792, DP_OP_424J2_126_3477_n1791,
         DP_OP_424J2_126_3477_n1790, DP_OP_424J2_126_3477_n1789,
         DP_OP_424J2_126_3477_n1788, DP_OP_424J2_126_3477_n1787,
         DP_OP_424J2_126_3477_n1786, DP_OP_424J2_126_3477_n1785,
         DP_OP_424J2_126_3477_n1784, DP_OP_424J2_126_3477_n1783,
         DP_OP_424J2_126_3477_n1782, DP_OP_424J2_126_3477_n1781,
         DP_OP_424J2_126_3477_n1780, DP_OP_424J2_126_3477_n1779,
         DP_OP_424J2_126_3477_n1778, DP_OP_424J2_126_3477_n1777,
         DP_OP_424J2_126_3477_n1776, DP_OP_424J2_126_3477_n1775,
         DP_OP_424J2_126_3477_n1774, DP_OP_424J2_126_3477_n1773,
         DP_OP_424J2_126_3477_n1772, DP_OP_424J2_126_3477_n1771,
         DP_OP_424J2_126_3477_n1770, DP_OP_424J2_126_3477_n1769,
         DP_OP_424J2_126_3477_n1768, DP_OP_424J2_126_3477_n1767,
         DP_OP_424J2_126_3477_n1766, DP_OP_424J2_126_3477_n1765,
         DP_OP_424J2_126_3477_n1764, DP_OP_424J2_126_3477_n1763,
         DP_OP_424J2_126_3477_n1762, DP_OP_424J2_126_3477_n1761,
         DP_OP_424J2_126_3477_n1760, DP_OP_424J2_126_3477_n1759,
         DP_OP_424J2_126_3477_n1758, DP_OP_424J2_126_3477_n1757,
         DP_OP_424J2_126_3477_n1756, DP_OP_424J2_126_3477_n1755,
         DP_OP_424J2_126_3477_n1754, DP_OP_424J2_126_3477_n1753,
         DP_OP_424J2_126_3477_n1752, DP_OP_424J2_126_3477_n1751,
         DP_OP_424J2_126_3477_n1750, DP_OP_424J2_126_3477_n1749,
         DP_OP_424J2_126_3477_n1748, DP_OP_424J2_126_3477_n1747,
         DP_OP_424J2_126_3477_n1746, DP_OP_424J2_126_3477_n1745,
         DP_OP_424J2_126_3477_n1744, DP_OP_424J2_126_3477_n1743,
         DP_OP_424J2_126_3477_n1742, DP_OP_424J2_126_3477_n1741,
         DP_OP_424J2_126_3477_n1740, DP_OP_424J2_126_3477_n1739,
         DP_OP_424J2_126_3477_n1738, DP_OP_424J2_126_3477_n1737,
         DP_OP_424J2_126_3477_n1736, DP_OP_424J2_126_3477_n1735,
         DP_OP_424J2_126_3477_n1734, DP_OP_424J2_126_3477_n1733,
         DP_OP_424J2_126_3477_n1732, DP_OP_424J2_126_3477_n1731,
         DP_OP_424J2_126_3477_n1730, DP_OP_424J2_126_3477_n1729,
         DP_OP_424J2_126_3477_n1728, DP_OP_424J2_126_3477_n1727,
         DP_OP_424J2_126_3477_n1726, DP_OP_424J2_126_3477_n1725,
         DP_OP_424J2_126_3477_n1724, DP_OP_424J2_126_3477_n1723,
         DP_OP_424J2_126_3477_n1722, DP_OP_424J2_126_3477_n1721,
         DP_OP_424J2_126_3477_n1720, DP_OP_424J2_126_3477_n1719,
         DP_OP_424J2_126_3477_n1718, DP_OP_424J2_126_3477_n1717,
         DP_OP_424J2_126_3477_n1716, DP_OP_424J2_126_3477_n1715,
         DP_OP_424J2_126_3477_n1714, DP_OP_424J2_126_3477_n1713,
         DP_OP_424J2_126_3477_n1712, DP_OP_424J2_126_3477_n1711,
         DP_OP_424J2_126_3477_n1710, DP_OP_424J2_126_3477_n1709,
         DP_OP_424J2_126_3477_n1708, DP_OP_424J2_126_3477_n1707,
         DP_OP_424J2_126_3477_n1706, DP_OP_424J2_126_3477_n1705,
         DP_OP_424J2_126_3477_n1704, DP_OP_424J2_126_3477_n1703,
         DP_OP_424J2_126_3477_n1702, DP_OP_424J2_126_3477_n1701,
         DP_OP_424J2_126_3477_n1700, DP_OP_424J2_126_3477_n1699,
         DP_OP_424J2_126_3477_n1698, DP_OP_424J2_126_3477_n1697,
         DP_OP_424J2_126_3477_n1696, DP_OP_424J2_126_3477_n1695,
         DP_OP_424J2_126_3477_n1694, DP_OP_424J2_126_3477_n1693,
         DP_OP_424J2_126_3477_n1692, DP_OP_424J2_126_3477_n1691,
         DP_OP_424J2_126_3477_n1690, DP_OP_424J2_126_3477_n1689,
         DP_OP_424J2_126_3477_n1688, DP_OP_424J2_126_3477_n1687,
         DP_OP_424J2_126_3477_n1686, DP_OP_424J2_126_3477_n1685,
         DP_OP_424J2_126_3477_n1684, DP_OP_424J2_126_3477_n1683,
         DP_OP_424J2_126_3477_n1682, DP_OP_424J2_126_3477_n1681,
         DP_OP_424J2_126_3477_n1680, DP_OP_424J2_126_3477_n1679,
         DP_OP_424J2_126_3477_n1678, DP_OP_424J2_126_3477_n1677,
         DP_OP_424J2_126_3477_n1676, DP_OP_424J2_126_3477_n1675,
         DP_OP_424J2_126_3477_n1674, DP_OP_424J2_126_3477_n1673,
         DP_OP_424J2_126_3477_n1672, DP_OP_424J2_126_3477_n1671,
         DP_OP_424J2_126_3477_n1670, DP_OP_424J2_126_3477_n1669,
         DP_OP_424J2_126_3477_n1668, DP_OP_424J2_126_3477_n1667,
         DP_OP_424J2_126_3477_n1666, DP_OP_424J2_126_3477_n1665,
         DP_OP_424J2_126_3477_n1664, DP_OP_424J2_126_3477_n1663,
         DP_OP_424J2_126_3477_n1662, DP_OP_424J2_126_3477_n1661,
         DP_OP_424J2_126_3477_n1660, DP_OP_424J2_126_3477_n1659,
         DP_OP_424J2_126_3477_n1658, DP_OP_424J2_126_3477_n1657,
         DP_OP_424J2_126_3477_n1656, DP_OP_424J2_126_3477_n1655,
         DP_OP_424J2_126_3477_n1654, DP_OP_424J2_126_3477_n1653,
         DP_OP_424J2_126_3477_n1652, DP_OP_424J2_126_3477_n1651,
         DP_OP_424J2_126_3477_n1650, DP_OP_424J2_126_3477_n1649,
         DP_OP_424J2_126_3477_n1648, DP_OP_424J2_126_3477_n1647,
         DP_OP_424J2_126_3477_n1646, DP_OP_424J2_126_3477_n1645,
         DP_OP_424J2_126_3477_n1644, DP_OP_424J2_126_3477_n1643,
         DP_OP_424J2_126_3477_n1642, DP_OP_424J2_126_3477_n1641,
         DP_OP_424J2_126_3477_n1640, DP_OP_424J2_126_3477_n1639,
         DP_OP_424J2_126_3477_n1638, DP_OP_424J2_126_3477_n1637,
         DP_OP_424J2_126_3477_n1636, DP_OP_424J2_126_3477_n1635,
         DP_OP_424J2_126_3477_n1634, DP_OP_424J2_126_3477_n1633,
         DP_OP_424J2_126_3477_n1632, DP_OP_424J2_126_3477_n1631,
         DP_OP_424J2_126_3477_n1630, DP_OP_424J2_126_3477_n1629,
         DP_OP_424J2_126_3477_n1628, DP_OP_424J2_126_3477_n1627,
         DP_OP_424J2_126_3477_n1626, DP_OP_424J2_126_3477_n1625,
         DP_OP_424J2_126_3477_n1624, DP_OP_424J2_126_3477_n1623,
         DP_OP_424J2_126_3477_n1622, DP_OP_424J2_126_3477_n1621,
         DP_OP_424J2_126_3477_n1620, DP_OP_424J2_126_3477_n1619,
         DP_OP_424J2_126_3477_n1618, DP_OP_424J2_126_3477_n1617,
         DP_OP_424J2_126_3477_n1616, DP_OP_424J2_126_3477_n1615,
         DP_OP_424J2_126_3477_n1614, DP_OP_424J2_126_3477_n1613,
         DP_OP_424J2_126_3477_n1612, DP_OP_424J2_126_3477_n1611,
         DP_OP_424J2_126_3477_n1610, DP_OP_424J2_126_3477_n1609,
         DP_OP_424J2_126_3477_n1608, DP_OP_424J2_126_3477_n1607,
         DP_OP_424J2_126_3477_n1606, DP_OP_424J2_126_3477_n1605,
         DP_OP_424J2_126_3477_n1604, DP_OP_424J2_126_3477_n1603,
         DP_OP_424J2_126_3477_n1602, DP_OP_424J2_126_3477_n1601,
         DP_OP_424J2_126_3477_n1600, DP_OP_424J2_126_3477_n1599,
         DP_OP_424J2_126_3477_n1598, DP_OP_424J2_126_3477_n1597,
         DP_OP_424J2_126_3477_n1596, DP_OP_424J2_126_3477_n1595,
         DP_OP_424J2_126_3477_n1594, DP_OP_424J2_126_3477_n1593,
         DP_OP_424J2_126_3477_n1592, DP_OP_424J2_126_3477_n1591,
         DP_OP_424J2_126_3477_n1590, DP_OP_424J2_126_3477_n1589,
         DP_OP_424J2_126_3477_n1588, DP_OP_424J2_126_3477_n1587,
         DP_OP_424J2_126_3477_n1586, DP_OP_424J2_126_3477_n1585,
         DP_OP_424J2_126_3477_n1584, DP_OP_424J2_126_3477_n1583,
         DP_OP_424J2_126_3477_n1582, DP_OP_424J2_126_3477_n1581,
         DP_OP_424J2_126_3477_n1580, DP_OP_424J2_126_3477_n1579,
         DP_OP_424J2_126_3477_n1578, DP_OP_424J2_126_3477_n1577,
         DP_OP_424J2_126_3477_n1576, DP_OP_424J2_126_3477_n1575,
         DP_OP_424J2_126_3477_n1574, DP_OP_424J2_126_3477_n1573,
         DP_OP_424J2_126_3477_n1572, DP_OP_424J2_126_3477_n1571,
         DP_OP_424J2_126_3477_n1570, DP_OP_424J2_126_3477_n1569,
         DP_OP_424J2_126_3477_n1568, DP_OP_424J2_126_3477_n1567,
         DP_OP_424J2_126_3477_n1566, DP_OP_424J2_126_3477_n1565,
         DP_OP_424J2_126_3477_n1564, DP_OP_424J2_126_3477_n1563,
         DP_OP_424J2_126_3477_n1562, DP_OP_424J2_126_3477_n1561,
         DP_OP_424J2_126_3477_n1560, DP_OP_424J2_126_3477_n1559,
         DP_OP_424J2_126_3477_n1558, DP_OP_424J2_126_3477_n1557,
         DP_OP_424J2_126_3477_n1556, DP_OP_424J2_126_3477_n1555,
         DP_OP_424J2_126_3477_n1554, DP_OP_424J2_126_3477_n1553,
         DP_OP_424J2_126_3477_n1552, DP_OP_424J2_126_3477_n1551,
         DP_OP_424J2_126_3477_n1550, DP_OP_424J2_126_3477_n1549,
         DP_OP_424J2_126_3477_n1548, DP_OP_424J2_126_3477_n1547,
         DP_OP_424J2_126_3477_n1546, DP_OP_424J2_126_3477_n1545,
         DP_OP_424J2_126_3477_n1544, DP_OP_424J2_126_3477_n1543,
         DP_OP_424J2_126_3477_n1542, DP_OP_424J2_126_3477_n1541,
         DP_OP_424J2_126_3477_n1540, DP_OP_424J2_126_3477_n1539,
         DP_OP_424J2_126_3477_n1538, DP_OP_424J2_126_3477_n1537,
         DP_OP_424J2_126_3477_n1536, DP_OP_424J2_126_3477_n1535,
         DP_OP_424J2_126_3477_n1534, DP_OP_424J2_126_3477_n1533,
         DP_OP_424J2_126_3477_n1532, DP_OP_424J2_126_3477_n1531,
         DP_OP_424J2_126_3477_n1530, DP_OP_424J2_126_3477_n1529,
         DP_OP_424J2_126_3477_n1528, DP_OP_424J2_126_3477_n1527,
         DP_OP_424J2_126_3477_n1526, DP_OP_424J2_126_3477_n1525,
         DP_OP_424J2_126_3477_n1524, DP_OP_424J2_126_3477_n1523,
         DP_OP_424J2_126_3477_n1522, DP_OP_424J2_126_3477_n1521,
         DP_OP_424J2_126_3477_n1520, DP_OP_424J2_126_3477_n1519,
         DP_OP_424J2_126_3477_n1518, DP_OP_424J2_126_3477_n1517,
         DP_OP_424J2_126_3477_n1516, DP_OP_424J2_126_3477_n1515,
         DP_OP_424J2_126_3477_n1514, DP_OP_424J2_126_3477_n1513,
         DP_OP_424J2_126_3477_n1512, DP_OP_424J2_126_3477_n1511,
         DP_OP_424J2_126_3477_n1510, DP_OP_424J2_126_3477_n1509,
         DP_OP_424J2_126_3477_n1508, DP_OP_424J2_126_3477_n1507,
         DP_OP_424J2_126_3477_n1506, DP_OP_424J2_126_3477_n1505,
         DP_OP_424J2_126_3477_n1504, DP_OP_424J2_126_3477_n1503,
         DP_OP_424J2_126_3477_n1502, DP_OP_424J2_126_3477_n1501,
         DP_OP_424J2_126_3477_n1500, DP_OP_424J2_126_3477_n1499,
         DP_OP_424J2_126_3477_n1498, DP_OP_424J2_126_3477_n1497,
         DP_OP_424J2_126_3477_n1496, DP_OP_424J2_126_3477_n1495,
         DP_OP_424J2_126_3477_n1494, DP_OP_424J2_126_3477_n1493,
         DP_OP_424J2_126_3477_n1492, DP_OP_424J2_126_3477_n1491,
         DP_OP_424J2_126_3477_n1490, DP_OP_424J2_126_3477_n1489,
         DP_OP_424J2_126_3477_n1488, DP_OP_424J2_126_3477_n1487,
         DP_OP_424J2_126_3477_n1486, DP_OP_424J2_126_3477_n1485,
         DP_OP_424J2_126_3477_n1484, DP_OP_424J2_126_3477_n1483,
         DP_OP_424J2_126_3477_n1482, DP_OP_424J2_126_3477_n1481,
         DP_OP_424J2_126_3477_n1480, DP_OP_424J2_126_3477_n1479,
         DP_OP_424J2_126_3477_n1478, DP_OP_424J2_126_3477_n1477,
         DP_OP_424J2_126_3477_n1476, DP_OP_424J2_126_3477_n1475,
         DP_OP_424J2_126_3477_n1474, DP_OP_424J2_126_3477_n1473,
         DP_OP_424J2_126_3477_n1472, DP_OP_424J2_126_3477_n1471,
         DP_OP_424J2_126_3477_n1470, DP_OP_424J2_126_3477_n1469,
         DP_OP_424J2_126_3477_n1468, DP_OP_424J2_126_3477_n1467,
         DP_OP_424J2_126_3477_n1466, DP_OP_424J2_126_3477_n1465,
         DP_OP_424J2_126_3477_n1464, DP_OP_424J2_126_3477_n1463,
         DP_OP_424J2_126_3477_n1462, DP_OP_424J2_126_3477_n1461,
         DP_OP_424J2_126_3477_n1460, DP_OP_424J2_126_3477_n1459,
         DP_OP_424J2_126_3477_n1458, DP_OP_424J2_126_3477_n1457,
         DP_OP_424J2_126_3477_n1456, DP_OP_424J2_126_3477_n1455,
         DP_OP_424J2_126_3477_n1454, DP_OP_424J2_126_3477_n1453,
         DP_OP_424J2_126_3477_n1452, DP_OP_424J2_126_3477_n1451,
         DP_OP_424J2_126_3477_n1450, DP_OP_424J2_126_3477_n1449,
         DP_OP_424J2_126_3477_n1448, DP_OP_424J2_126_3477_n1447,
         DP_OP_424J2_126_3477_n1446, DP_OP_424J2_126_3477_n1445,
         DP_OP_424J2_126_3477_n1444, DP_OP_424J2_126_3477_n1443,
         DP_OP_424J2_126_3477_n1442, DP_OP_424J2_126_3477_n1441,
         DP_OP_424J2_126_3477_n1440, DP_OP_424J2_126_3477_n1439,
         DP_OP_424J2_126_3477_n1438, DP_OP_424J2_126_3477_n1437,
         DP_OP_424J2_126_3477_n1436, DP_OP_424J2_126_3477_n1435,
         DP_OP_424J2_126_3477_n1434, DP_OP_424J2_126_3477_n1433,
         DP_OP_424J2_126_3477_n1432, DP_OP_424J2_126_3477_n1431,
         DP_OP_424J2_126_3477_n1430, DP_OP_424J2_126_3477_n1429,
         DP_OP_424J2_126_3477_n1428, DP_OP_424J2_126_3477_n1427,
         DP_OP_424J2_126_3477_n1426, DP_OP_424J2_126_3477_n1425,
         DP_OP_424J2_126_3477_n1424, DP_OP_424J2_126_3477_n1423,
         DP_OP_424J2_126_3477_n1422, DP_OP_424J2_126_3477_n1421,
         DP_OP_424J2_126_3477_n1420, DP_OP_424J2_126_3477_n1419,
         DP_OP_424J2_126_3477_n1418, DP_OP_424J2_126_3477_n1417,
         DP_OP_424J2_126_3477_n1416, DP_OP_424J2_126_3477_n1415,
         DP_OP_424J2_126_3477_n1414, DP_OP_424J2_126_3477_n1413,
         DP_OP_424J2_126_3477_n1412, DP_OP_424J2_126_3477_n1411,
         DP_OP_424J2_126_3477_n1410, DP_OP_424J2_126_3477_n1409,
         DP_OP_424J2_126_3477_n1408, DP_OP_424J2_126_3477_n1407,
         DP_OP_424J2_126_3477_n1406, DP_OP_424J2_126_3477_n1405,
         DP_OP_424J2_126_3477_n1404, DP_OP_424J2_126_3477_n1403,
         DP_OP_424J2_126_3477_n1402, DP_OP_424J2_126_3477_n1401,
         DP_OP_424J2_126_3477_n1400, DP_OP_424J2_126_3477_n1399,
         DP_OP_424J2_126_3477_n1398, DP_OP_424J2_126_3477_n1397,
         DP_OP_424J2_126_3477_n1396, DP_OP_424J2_126_3477_n1395,
         DP_OP_424J2_126_3477_n1394, DP_OP_424J2_126_3477_n1393,
         DP_OP_424J2_126_3477_n1392, DP_OP_424J2_126_3477_n1391,
         DP_OP_424J2_126_3477_n1390, DP_OP_424J2_126_3477_n1389,
         DP_OP_424J2_126_3477_n1388, DP_OP_424J2_126_3477_n1387,
         DP_OP_424J2_126_3477_n1386, DP_OP_424J2_126_3477_n1385,
         DP_OP_424J2_126_3477_n1384, DP_OP_424J2_126_3477_n1383,
         DP_OP_424J2_126_3477_n1382, DP_OP_424J2_126_3477_n1381,
         DP_OP_424J2_126_3477_n1380, DP_OP_424J2_126_3477_n1379,
         DP_OP_424J2_126_3477_n1378, DP_OP_424J2_126_3477_n1377,
         DP_OP_424J2_126_3477_n1376, DP_OP_424J2_126_3477_n1375,
         DP_OP_424J2_126_3477_n1374, DP_OP_424J2_126_3477_n1373,
         DP_OP_424J2_126_3477_n1372, DP_OP_424J2_126_3477_n1371,
         DP_OP_424J2_126_3477_n1370, DP_OP_424J2_126_3477_n1369,
         DP_OP_424J2_126_3477_n1368, DP_OP_424J2_126_3477_n1367,
         DP_OP_424J2_126_3477_n1366, DP_OP_424J2_126_3477_n1365,
         DP_OP_424J2_126_3477_n1364, DP_OP_424J2_126_3477_n1363,
         DP_OP_424J2_126_3477_n1362, DP_OP_424J2_126_3477_n1361,
         DP_OP_424J2_126_3477_n1360, DP_OP_424J2_126_3477_n1359,
         DP_OP_424J2_126_3477_n1358, DP_OP_424J2_126_3477_n1357,
         DP_OP_424J2_126_3477_n1356, DP_OP_424J2_126_3477_n1355,
         DP_OP_424J2_126_3477_n1354, DP_OP_424J2_126_3477_n1353,
         DP_OP_424J2_126_3477_n1352, DP_OP_424J2_126_3477_n1351,
         DP_OP_424J2_126_3477_n1350, DP_OP_424J2_126_3477_n1349,
         DP_OP_424J2_126_3477_n1348, DP_OP_424J2_126_3477_n1347,
         DP_OP_424J2_126_3477_n1346, DP_OP_424J2_126_3477_n1345,
         DP_OP_424J2_126_3477_n1344, DP_OP_424J2_126_3477_n1343,
         DP_OP_424J2_126_3477_n1342, DP_OP_424J2_126_3477_n1341,
         DP_OP_424J2_126_3477_n1340, DP_OP_424J2_126_3477_n1339,
         DP_OP_424J2_126_3477_n1338, DP_OP_424J2_126_3477_n1337,
         DP_OP_424J2_126_3477_n1336, DP_OP_424J2_126_3477_n1335,
         DP_OP_424J2_126_3477_n1334, DP_OP_424J2_126_3477_n1333,
         DP_OP_424J2_126_3477_n1332, DP_OP_424J2_126_3477_n1331,
         DP_OP_424J2_126_3477_n1330, DP_OP_424J2_126_3477_n1329,
         DP_OP_424J2_126_3477_n1328, DP_OP_424J2_126_3477_n1327,
         DP_OP_424J2_126_3477_n1326, DP_OP_424J2_126_3477_n1325,
         DP_OP_424J2_126_3477_n1324, DP_OP_424J2_126_3477_n1323,
         DP_OP_424J2_126_3477_n1322, DP_OP_424J2_126_3477_n1321,
         DP_OP_424J2_126_3477_n1320, DP_OP_424J2_126_3477_n1319,
         DP_OP_424J2_126_3477_n1318, DP_OP_424J2_126_3477_n1317,
         DP_OP_424J2_126_3477_n1316, DP_OP_424J2_126_3477_n1315,
         DP_OP_424J2_126_3477_n1314, DP_OP_424J2_126_3477_n1313,
         DP_OP_424J2_126_3477_n1312, DP_OP_424J2_126_3477_n1311,
         DP_OP_424J2_126_3477_n1310, DP_OP_424J2_126_3477_n1309,
         DP_OP_424J2_126_3477_n1308, DP_OP_424J2_126_3477_n1307,
         DP_OP_424J2_126_3477_n1306, DP_OP_424J2_126_3477_n1305,
         DP_OP_424J2_126_3477_n1304, DP_OP_424J2_126_3477_n1303,
         DP_OP_424J2_126_3477_n1302, DP_OP_424J2_126_3477_n1301,
         DP_OP_424J2_126_3477_n1300, DP_OP_424J2_126_3477_n1299,
         DP_OP_424J2_126_3477_n1298, DP_OP_424J2_126_3477_n1297,
         DP_OP_424J2_126_3477_n1296, DP_OP_424J2_126_3477_n1295,
         DP_OP_424J2_126_3477_n1294, DP_OP_424J2_126_3477_n1293,
         DP_OP_424J2_126_3477_n1292, DP_OP_424J2_126_3477_n1291,
         DP_OP_424J2_126_3477_n1290, DP_OP_424J2_126_3477_n1289,
         DP_OP_424J2_126_3477_n1288, DP_OP_424J2_126_3477_n1287,
         DP_OP_424J2_126_3477_n1286, DP_OP_424J2_126_3477_n1285,
         DP_OP_424J2_126_3477_n1284, DP_OP_424J2_126_3477_n1283,
         DP_OP_424J2_126_3477_n1282, DP_OP_424J2_126_3477_n1281,
         DP_OP_424J2_126_3477_n1280, DP_OP_424J2_126_3477_n1279,
         DP_OP_424J2_126_3477_n1278, DP_OP_424J2_126_3477_n1277,
         DP_OP_424J2_126_3477_n1276, DP_OP_424J2_126_3477_n1275,
         DP_OP_424J2_126_3477_n1274, DP_OP_424J2_126_3477_n1273,
         DP_OP_424J2_126_3477_n1272, DP_OP_424J2_126_3477_n1271,
         DP_OP_424J2_126_3477_n1270, DP_OP_424J2_126_3477_n1269,
         DP_OP_424J2_126_3477_n1268, DP_OP_424J2_126_3477_n1267,
         DP_OP_424J2_126_3477_n1266, DP_OP_424J2_126_3477_n1265,
         DP_OP_424J2_126_3477_n1264, DP_OP_424J2_126_3477_n1263,
         DP_OP_424J2_126_3477_n1262, DP_OP_424J2_126_3477_n1261,
         DP_OP_424J2_126_3477_n1260, DP_OP_424J2_126_3477_n1259,
         DP_OP_424J2_126_3477_n1258, DP_OP_424J2_126_3477_n1257,
         DP_OP_424J2_126_3477_n1256, DP_OP_424J2_126_3477_n1255,
         DP_OP_424J2_126_3477_n1254, DP_OP_424J2_126_3477_n1253,
         DP_OP_424J2_126_3477_n1252, DP_OP_424J2_126_3477_n1251,
         DP_OP_424J2_126_3477_n1250, DP_OP_424J2_126_3477_n1249,
         DP_OP_424J2_126_3477_n1248, DP_OP_424J2_126_3477_n1247,
         DP_OP_424J2_126_3477_n1246, DP_OP_424J2_126_3477_n1245,
         DP_OP_424J2_126_3477_n1244, DP_OP_424J2_126_3477_n1243,
         DP_OP_424J2_126_3477_n1242, DP_OP_424J2_126_3477_n1241,
         DP_OP_424J2_126_3477_n1240, DP_OP_424J2_126_3477_n1239,
         DP_OP_424J2_126_3477_n1238, DP_OP_424J2_126_3477_n1237,
         DP_OP_424J2_126_3477_n1236, DP_OP_424J2_126_3477_n1235,
         DP_OP_424J2_126_3477_n1234, DP_OP_424J2_126_3477_n1233,
         DP_OP_424J2_126_3477_n1232, DP_OP_424J2_126_3477_n1231,
         DP_OP_424J2_126_3477_n1230, DP_OP_424J2_126_3477_n1229,
         DP_OP_424J2_126_3477_n1228, DP_OP_424J2_126_3477_n1227,
         DP_OP_424J2_126_3477_n1226, DP_OP_424J2_126_3477_n1225,
         DP_OP_424J2_126_3477_n1224, DP_OP_424J2_126_3477_n1223,
         DP_OP_424J2_126_3477_n1222, DP_OP_424J2_126_3477_n1221,
         DP_OP_424J2_126_3477_n1220, DP_OP_424J2_126_3477_n1219,
         DP_OP_424J2_126_3477_n1218, DP_OP_424J2_126_3477_n1217,
         DP_OP_424J2_126_3477_n1216, DP_OP_424J2_126_3477_n1215,
         DP_OP_424J2_126_3477_n1214, DP_OP_424J2_126_3477_n1213,
         DP_OP_424J2_126_3477_n1212, DP_OP_424J2_126_3477_n1211,
         DP_OP_424J2_126_3477_n1210, DP_OP_424J2_126_3477_n1209,
         DP_OP_424J2_126_3477_n1208, DP_OP_424J2_126_3477_n1207,
         DP_OP_424J2_126_3477_n1206, DP_OP_424J2_126_3477_n1205,
         DP_OP_424J2_126_3477_n1204, DP_OP_424J2_126_3477_n1203,
         DP_OP_424J2_126_3477_n1202, DP_OP_424J2_126_3477_n1201,
         DP_OP_424J2_126_3477_n1200, DP_OP_424J2_126_3477_n1199,
         DP_OP_424J2_126_3477_n1198, DP_OP_424J2_126_3477_n1197,
         DP_OP_424J2_126_3477_n1196, DP_OP_424J2_126_3477_n1195,
         DP_OP_424J2_126_3477_n1194, DP_OP_424J2_126_3477_n1193,
         DP_OP_424J2_126_3477_n1192, DP_OP_424J2_126_3477_n1191,
         DP_OP_424J2_126_3477_n1190, DP_OP_424J2_126_3477_n1189,
         DP_OP_424J2_126_3477_n1188, DP_OP_424J2_126_3477_n1187,
         DP_OP_424J2_126_3477_n1186, DP_OP_424J2_126_3477_n1185,
         DP_OP_424J2_126_3477_n1184, DP_OP_424J2_126_3477_n1183,
         DP_OP_424J2_126_3477_n1182, DP_OP_424J2_126_3477_n1181,
         DP_OP_424J2_126_3477_n1180, DP_OP_424J2_126_3477_n1179,
         DP_OP_424J2_126_3477_n1178, DP_OP_424J2_126_3477_n1177,
         DP_OP_424J2_126_3477_n1176, DP_OP_424J2_126_3477_n1175,
         DP_OP_424J2_126_3477_n1174, DP_OP_424J2_126_3477_n1173,
         DP_OP_424J2_126_3477_n1172, DP_OP_424J2_126_3477_n1171,
         DP_OP_424J2_126_3477_n1170, DP_OP_424J2_126_3477_n1169,
         DP_OP_424J2_126_3477_n1168, DP_OP_424J2_126_3477_n1167,
         DP_OP_424J2_126_3477_n1166, DP_OP_424J2_126_3477_n1165,
         DP_OP_424J2_126_3477_n1164, DP_OP_424J2_126_3477_n1163,
         DP_OP_424J2_126_3477_n1162, DP_OP_424J2_126_3477_n1161,
         DP_OP_424J2_126_3477_n1160, DP_OP_424J2_126_3477_n1159,
         DP_OP_424J2_126_3477_n1158, DP_OP_424J2_126_3477_n1157,
         DP_OP_424J2_126_3477_n1156, DP_OP_424J2_126_3477_n1155,
         DP_OP_424J2_126_3477_n1154, DP_OP_424J2_126_3477_n1153,
         DP_OP_424J2_126_3477_n1152, DP_OP_424J2_126_3477_n1151,
         DP_OP_424J2_126_3477_n1150, DP_OP_424J2_126_3477_n1149,
         DP_OP_424J2_126_3477_n1148, DP_OP_424J2_126_3477_n1147,
         DP_OP_424J2_126_3477_n1146, DP_OP_424J2_126_3477_n1145,
         DP_OP_424J2_126_3477_n1144, DP_OP_424J2_126_3477_n1143,
         DP_OP_424J2_126_3477_n1142, DP_OP_424J2_126_3477_n1141,
         DP_OP_424J2_126_3477_n1140, DP_OP_424J2_126_3477_n1139,
         DP_OP_424J2_126_3477_n1138, DP_OP_424J2_126_3477_n1137,
         DP_OP_424J2_126_3477_n1136, DP_OP_424J2_126_3477_n1135,
         DP_OP_424J2_126_3477_n1134, DP_OP_424J2_126_3477_n1133,
         DP_OP_424J2_126_3477_n1132, DP_OP_424J2_126_3477_n1131,
         DP_OP_424J2_126_3477_n1130, DP_OP_424J2_126_3477_n1129,
         DP_OP_424J2_126_3477_n1128, DP_OP_424J2_126_3477_n1127,
         DP_OP_424J2_126_3477_n1126, DP_OP_424J2_126_3477_n1125,
         DP_OP_424J2_126_3477_n1124, DP_OP_424J2_126_3477_n1123,
         DP_OP_424J2_126_3477_n1122, DP_OP_424J2_126_3477_n1121,
         DP_OP_424J2_126_3477_n1120, DP_OP_424J2_126_3477_n1119,
         DP_OP_424J2_126_3477_n1118, DP_OP_424J2_126_3477_n1117,
         DP_OP_424J2_126_3477_n1116, DP_OP_424J2_126_3477_n1115,
         DP_OP_424J2_126_3477_n1114, DP_OP_424J2_126_3477_n1113,
         DP_OP_424J2_126_3477_n1112, DP_OP_424J2_126_3477_n1111,
         DP_OP_424J2_126_3477_n1110, DP_OP_424J2_126_3477_n1109,
         DP_OP_424J2_126_3477_n1108, DP_OP_424J2_126_3477_n1107,
         DP_OP_424J2_126_3477_n1106, DP_OP_424J2_126_3477_n1105,
         DP_OP_424J2_126_3477_n1104, DP_OP_424J2_126_3477_n1103,
         DP_OP_424J2_126_3477_n1102, DP_OP_424J2_126_3477_n1101,
         DP_OP_424J2_126_3477_n1100, DP_OP_424J2_126_3477_n1099,
         DP_OP_424J2_126_3477_n1098, DP_OP_424J2_126_3477_n1097,
         DP_OP_424J2_126_3477_n1096, DP_OP_424J2_126_3477_n1095,
         DP_OP_424J2_126_3477_n1094, DP_OP_424J2_126_3477_n1093,
         DP_OP_424J2_126_3477_n1092, DP_OP_424J2_126_3477_n1091,
         DP_OP_424J2_126_3477_n1090, DP_OP_424J2_126_3477_n1089,
         DP_OP_424J2_126_3477_n1088, DP_OP_424J2_126_3477_n1087,
         DP_OP_424J2_126_3477_n1086, DP_OP_424J2_126_3477_n1085,
         DP_OP_424J2_126_3477_n1084, DP_OP_424J2_126_3477_n1083,
         DP_OP_424J2_126_3477_n1082, DP_OP_424J2_126_3477_n1081,
         DP_OP_424J2_126_3477_n1080, DP_OP_424J2_126_3477_n1079,
         DP_OP_424J2_126_3477_n1078, DP_OP_424J2_126_3477_n1077,
         DP_OP_424J2_126_3477_n1076, DP_OP_424J2_126_3477_n1075,
         DP_OP_424J2_126_3477_n1074, DP_OP_424J2_126_3477_n1073,
         DP_OP_424J2_126_3477_n1072, DP_OP_424J2_126_3477_n1071,
         DP_OP_424J2_126_3477_n1070, DP_OP_424J2_126_3477_n1069,
         DP_OP_424J2_126_3477_n1068, DP_OP_424J2_126_3477_n1067,
         DP_OP_424J2_126_3477_n1066, DP_OP_424J2_126_3477_n1065,
         DP_OP_424J2_126_3477_n1064, DP_OP_424J2_126_3477_n1063,
         DP_OP_424J2_126_3477_n1062, DP_OP_424J2_126_3477_n1061,
         DP_OP_424J2_126_3477_n1060, DP_OP_424J2_126_3477_n1059,
         DP_OP_424J2_126_3477_n1058, DP_OP_424J2_126_3477_n1057,
         DP_OP_424J2_126_3477_n1056, DP_OP_424J2_126_3477_n1055,
         DP_OP_424J2_126_3477_n1054, DP_OP_424J2_126_3477_n1053,
         DP_OP_424J2_126_3477_n1052, DP_OP_424J2_126_3477_n1051,
         DP_OP_424J2_126_3477_n1050, DP_OP_424J2_126_3477_n1049,
         DP_OP_424J2_126_3477_n1048, DP_OP_424J2_126_3477_n1047,
         DP_OP_424J2_126_3477_n1046, DP_OP_424J2_126_3477_n1045,
         DP_OP_424J2_126_3477_n1044, DP_OP_424J2_126_3477_n1043,
         DP_OP_424J2_126_3477_n1042, DP_OP_424J2_126_3477_n1041,
         DP_OP_424J2_126_3477_n1040, DP_OP_424J2_126_3477_n1039,
         DP_OP_424J2_126_3477_n1038, DP_OP_424J2_126_3477_n1037,
         DP_OP_424J2_126_3477_n1036, DP_OP_424J2_126_3477_n1035,
         DP_OP_424J2_126_3477_n1034, DP_OP_424J2_126_3477_n1033,
         DP_OP_424J2_126_3477_n1032, DP_OP_424J2_126_3477_n1031,
         DP_OP_424J2_126_3477_n1030, DP_OP_424J2_126_3477_n1029,
         DP_OP_424J2_126_3477_n1028, DP_OP_424J2_126_3477_n1027,
         DP_OP_424J2_126_3477_n1026, DP_OP_424J2_126_3477_n1025,
         DP_OP_424J2_126_3477_n1024, DP_OP_424J2_126_3477_n1023,
         DP_OP_424J2_126_3477_n1022, DP_OP_424J2_126_3477_n1021,
         DP_OP_424J2_126_3477_n1020, DP_OP_424J2_126_3477_n1019,
         DP_OP_424J2_126_3477_n1018, DP_OP_424J2_126_3477_n1017,
         DP_OP_424J2_126_3477_n1016, DP_OP_424J2_126_3477_n1015,
         DP_OP_424J2_126_3477_n1014, DP_OP_424J2_126_3477_n1013,
         DP_OP_424J2_126_3477_n1012, DP_OP_424J2_126_3477_n1011,
         DP_OP_424J2_126_3477_n1010, DP_OP_424J2_126_3477_n1009,
         DP_OP_424J2_126_3477_n1008, DP_OP_424J2_126_3477_n1007,
         DP_OP_424J2_126_3477_n1006, DP_OP_424J2_126_3477_n1005,
         DP_OP_424J2_126_3477_n1004, DP_OP_424J2_126_3477_n1003,
         DP_OP_424J2_126_3477_n1002, DP_OP_424J2_126_3477_n1001,
         DP_OP_424J2_126_3477_n1000, DP_OP_424J2_126_3477_n999,
         DP_OP_424J2_126_3477_n998, DP_OP_424J2_126_3477_n997,
         DP_OP_424J2_126_3477_n996, DP_OP_424J2_126_3477_n995,
         DP_OP_424J2_126_3477_n994, DP_OP_424J2_126_3477_n993,
         DP_OP_424J2_126_3477_n992, DP_OP_424J2_126_3477_n991,
         DP_OP_424J2_126_3477_n990, DP_OP_424J2_126_3477_n989,
         DP_OP_424J2_126_3477_n988, DP_OP_424J2_126_3477_n987,
         DP_OP_424J2_126_3477_n986, DP_OP_424J2_126_3477_n985,
         DP_OP_424J2_126_3477_n984, DP_OP_424J2_126_3477_n983,
         DP_OP_424J2_126_3477_n982, DP_OP_424J2_126_3477_n981,
         DP_OP_424J2_126_3477_n980, DP_OP_424J2_126_3477_n979,
         DP_OP_424J2_126_3477_n978, DP_OP_424J2_126_3477_n977,
         DP_OP_424J2_126_3477_n976, DP_OP_424J2_126_3477_n975,
         DP_OP_424J2_126_3477_n974, DP_OP_424J2_126_3477_n973,
         DP_OP_424J2_126_3477_n972, DP_OP_424J2_126_3477_n971,
         DP_OP_424J2_126_3477_n970, DP_OP_424J2_126_3477_n969,
         DP_OP_424J2_126_3477_n968, DP_OP_424J2_126_3477_n967,
         DP_OP_424J2_126_3477_n966, DP_OP_424J2_126_3477_n965,
         DP_OP_424J2_126_3477_n964, DP_OP_424J2_126_3477_n963,
         DP_OP_424J2_126_3477_n962, DP_OP_424J2_126_3477_n961,
         DP_OP_424J2_126_3477_n960, DP_OP_424J2_126_3477_n959,
         DP_OP_424J2_126_3477_n958, DP_OP_424J2_126_3477_n957,
         DP_OP_424J2_126_3477_n956, DP_OP_424J2_126_3477_n955,
         DP_OP_424J2_126_3477_n954, DP_OP_424J2_126_3477_n953,
         DP_OP_424J2_126_3477_n952, DP_OP_424J2_126_3477_n951,
         DP_OP_424J2_126_3477_n950, DP_OP_424J2_126_3477_n949,
         DP_OP_424J2_126_3477_n948, DP_OP_424J2_126_3477_n947,
         DP_OP_424J2_126_3477_n946, DP_OP_424J2_126_3477_n945,
         DP_OP_424J2_126_3477_n944, DP_OP_424J2_126_3477_n943,
         DP_OP_424J2_126_3477_n942, DP_OP_424J2_126_3477_n941,
         DP_OP_424J2_126_3477_n940, DP_OP_424J2_126_3477_n939,
         DP_OP_424J2_126_3477_n938, DP_OP_424J2_126_3477_n937,
         DP_OP_424J2_126_3477_n936, DP_OP_424J2_126_3477_n935,
         DP_OP_424J2_126_3477_n934, DP_OP_424J2_126_3477_n933,
         DP_OP_424J2_126_3477_n932, DP_OP_424J2_126_3477_n931,
         DP_OP_424J2_126_3477_n930, DP_OP_424J2_126_3477_n929,
         DP_OP_424J2_126_3477_n928, DP_OP_424J2_126_3477_n927,
         DP_OP_424J2_126_3477_n926, DP_OP_424J2_126_3477_n925,
         DP_OP_424J2_126_3477_n924, DP_OP_424J2_126_3477_n923,
         DP_OP_424J2_126_3477_n922, DP_OP_424J2_126_3477_n921,
         DP_OP_424J2_126_3477_n920, DP_OP_424J2_126_3477_n919,
         DP_OP_424J2_126_3477_n918, DP_OP_424J2_126_3477_n917,
         DP_OP_424J2_126_3477_n916, DP_OP_424J2_126_3477_n915,
         DP_OP_424J2_126_3477_n914, DP_OP_424J2_126_3477_n913,
         DP_OP_424J2_126_3477_n912, DP_OP_424J2_126_3477_n911,
         DP_OP_424J2_126_3477_n910, DP_OP_424J2_126_3477_n909,
         DP_OP_424J2_126_3477_n908, DP_OP_424J2_126_3477_n907,
         DP_OP_424J2_126_3477_n906, DP_OP_424J2_126_3477_n905,
         DP_OP_424J2_126_3477_n904, DP_OP_424J2_126_3477_n903,
         DP_OP_424J2_126_3477_n902, DP_OP_424J2_126_3477_n901,
         DP_OP_424J2_126_3477_n900, DP_OP_424J2_126_3477_n899,
         DP_OP_424J2_126_3477_n898, DP_OP_424J2_126_3477_n897,
         DP_OP_424J2_126_3477_n896, DP_OP_424J2_126_3477_n895,
         DP_OP_424J2_126_3477_n894, DP_OP_424J2_126_3477_n893,
         DP_OP_424J2_126_3477_n892, DP_OP_424J2_126_3477_n891,
         DP_OP_424J2_126_3477_n890, DP_OP_424J2_126_3477_n889,
         DP_OP_424J2_126_3477_n888, DP_OP_424J2_126_3477_n887,
         DP_OP_424J2_126_3477_n886, DP_OP_424J2_126_3477_n885,
         DP_OP_424J2_126_3477_n884, DP_OP_424J2_126_3477_n883,
         DP_OP_424J2_126_3477_n882, DP_OP_424J2_126_3477_n881,
         DP_OP_424J2_126_3477_n880, DP_OP_424J2_126_3477_n879,
         DP_OP_424J2_126_3477_n878, DP_OP_424J2_126_3477_n877,
         DP_OP_424J2_126_3477_n876, DP_OP_424J2_126_3477_n875,
         DP_OP_424J2_126_3477_n874, DP_OP_424J2_126_3477_n873,
         DP_OP_424J2_126_3477_n872, DP_OP_424J2_126_3477_n871,
         DP_OP_424J2_126_3477_n870, DP_OP_424J2_126_3477_n869,
         DP_OP_424J2_126_3477_n868, DP_OP_424J2_126_3477_n867,
         DP_OP_424J2_126_3477_n866, DP_OP_424J2_126_3477_n865,
         DP_OP_424J2_126_3477_n864, DP_OP_424J2_126_3477_n863,
         DP_OP_424J2_126_3477_n862, DP_OP_424J2_126_3477_n861,
         DP_OP_424J2_126_3477_n860, DP_OP_424J2_126_3477_n859,
         DP_OP_424J2_126_3477_n858, DP_OP_424J2_126_3477_n857,
         DP_OP_424J2_126_3477_n856, DP_OP_424J2_126_3477_n855,
         DP_OP_424J2_126_3477_n854, DP_OP_424J2_126_3477_n853,
         DP_OP_424J2_126_3477_n852, DP_OP_424J2_126_3477_n851,
         DP_OP_424J2_126_3477_n850, DP_OP_424J2_126_3477_n849,
         DP_OP_424J2_126_3477_n848, DP_OP_424J2_126_3477_n847,
         DP_OP_424J2_126_3477_n846, DP_OP_424J2_126_3477_n845,
         DP_OP_424J2_126_3477_n844, DP_OP_424J2_126_3477_n843,
         DP_OP_424J2_126_3477_n842, DP_OP_424J2_126_3477_n841,
         DP_OP_424J2_126_3477_n840, DP_OP_424J2_126_3477_n839,
         DP_OP_424J2_126_3477_n838, DP_OP_424J2_126_3477_n837,
         DP_OP_424J2_126_3477_n836, DP_OP_424J2_126_3477_n835,
         DP_OP_424J2_126_3477_n834, DP_OP_424J2_126_3477_n833,
         DP_OP_424J2_126_3477_n832, DP_OP_424J2_126_3477_n831,
         DP_OP_424J2_126_3477_n830, DP_OP_424J2_126_3477_n829,
         DP_OP_424J2_126_3477_n828, DP_OP_424J2_126_3477_n827,
         DP_OP_424J2_126_3477_n826, DP_OP_424J2_126_3477_n825,
         DP_OP_424J2_126_3477_n824, DP_OP_424J2_126_3477_n823,
         DP_OP_424J2_126_3477_n822, DP_OP_424J2_126_3477_n821,
         DP_OP_424J2_126_3477_n820, DP_OP_424J2_126_3477_n819,
         DP_OP_424J2_126_3477_n818, DP_OP_424J2_126_3477_n817,
         DP_OP_424J2_126_3477_n816, DP_OP_424J2_126_3477_n815,
         DP_OP_424J2_126_3477_n814, DP_OP_424J2_126_3477_n813,
         DP_OP_424J2_126_3477_n812, DP_OP_424J2_126_3477_n811,
         DP_OP_424J2_126_3477_n810, DP_OP_424J2_126_3477_n809,
         DP_OP_424J2_126_3477_n808, DP_OP_424J2_126_3477_n807,
         DP_OP_424J2_126_3477_n806, DP_OP_424J2_126_3477_n805,
         DP_OP_424J2_126_3477_n804, DP_OP_424J2_126_3477_n803,
         DP_OP_424J2_126_3477_n802, DP_OP_424J2_126_3477_n801,
         DP_OP_424J2_126_3477_n800, DP_OP_424J2_126_3477_n799,
         DP_OP_424J2_126_3477_n798, DP_OP_424J2_126_3477_n797,
         DP_OP_424J2_126_3477_n796, DP_OP_424J2_126_3477_n795,
         DP_OP_424J2_126_3477_n794, DP_OP_424J2_126_3477_n793,
         DP_OP_424J2_126_3477_n792, DP_OP_424J2_126_3477_n791,
         DP_OP_424J2_126_3477_n790, DP_OP_424J2_126_3477_n789,
         DP_OP_424J2_126_3477_n788, DP_OP_424J2_126_3477_n787,
         DP_OP_424J2_126_3477_n786, DP_OP_424J2_126_3477_n785,
         DP_OP_424J2_126_3477_n784, DP_OP_424J2_126_3477_n783,
         DP_OP_424J2_126_3477_n782, DP_OP_424J2_126_3477_n781,
         DP_OP_424J2_126_3477_n780, DP_OP_424J2_126_3477_n779,
         DP_OP_424J2_126_3477_n778, DP_OP_424J2_126_3477_n777,
         DP_OP_424J2_126_3477_n776, DP_OP_424J2_126_3477_n775,
         DP_OP_424J2_126_3477_n774, DP_OP_424J2_126_3477_n773,
         DP_OP_424J2_126_3477_n772, DP_OP_424J2_126_3477_n771,
         DP_OP_424J2_126_3477_n770, DP_OP_424J2_126_3477_n769,
         DP_OP_424J2_126_3477_n768, DP_OP_424J2_126_3477_n767,
         DP_OP_424J2_126_3477_n766, DP_OP_424J2_126_3477_n765,
         DP_OP_424J2_126_3477_n764, DP_OP_424J2_126_3477_n763,
         DP_OP_424J2_126_3477_n762, DP_OP_424J2_126_3477_n761,
         DP_OP_424J2_126_3477_n760, DP_OP_424J2_126_3477_n759,
         DP_OP_424J2_126_3477_n758, DP_OP_424J2_126_3477_n757,
         DP_OP_424J2_126_3477_n756, DP_OP_424J2_126_3477_n755,
         DP_OP_424J2_126_3477_n754, DP_OP_424J2_126_3477_n753,
         DP_OP_424J2_126_3477_n752, DP_OP_424J2_126_3477_n751,
         DP_OP_424J2_126_3477_n750, DP_OP_424J2_126_3477_n749,
         DP_OP_424J2_126_3477_n748, DP_OP_424J2_126_3477_n747,
         DP_OP_424J2_126_3477_n746, DP_OP_424J2_126_3477_n745,
         DP_OP_424J2_126_3477_n744, DP_OP_424J2_126_3477_n743,
         DP_OP_424J2_126_3477_n742, DP_OP_424J2_126_3477_n741,
         DP_OP_424J2_126_3477_n740, DP_OP_424J2_126_3477_n739,
         DP_OP_424J2_126_3477_n738, DP_OP_424J2_126_3477_n737,
         DP_OP_424J2_126_3477_n736, DP_OP_424J2_126_3477_n735,
         DP_OP_424J2_126_3477_n734, DP_OP_424J2_126_3477_n733,
         DP_OP_424J2_126_3477_n732, DP_OP_424J2_126_3477_n731,
         DP_OP_424J2_126_3477_n730, DP_OP_424J2_126_3477_n729,
         DP_OP_424J2_126_3477_n728, DP_OP_424J2_126_3477_n727,
         DP_OP_424J2_126_3477_n726, DP_OP_424J2_126_3477_n725,
         DP_OP_424J2_126_3477_n724, DP_OP_424J2_126_3477_n723,
         DP_OP_424J2_126_3477_n722, DP_OP_424J2_126_3477_n721,
         DP_OP_424J2_126_3477_n720, DP_OP_424J2_126_3477_n719,
         DP_OP_424J2_126_3477_n718, DP_OP_424J2_126_3477_n717,
         DP_OP_424J2_126_3477_n716, DP_OP_424J2_126_3477_n715,
         DP_OP_424J2_126_3477_n714, DP_OP_424J2_126_3477_n713,
         DP_OP_424J2_126_3477_n712, DP_OP_424J2_126_3477_n711,
         DP_OP_424J2_126_3477_n710, DP_OP_424J2_126_3477_n709,
         DP_OP_424J2_126_3477_n708, DP_OP_424J2_126_3477_n707,
         DP_OP_424J2_126_3477_n706, DP_OP_424J2_126_3477_n705,
         DP_OP_424J2_126_3477_n704, DP_OP_424J2_126_3477_n703,
         DP_OP_424J2_126_3477_n702, DP_OP_424J2_126_3477_n701,
         DP_OP_424J2_126_3477_n700, DP_OP_424J2_126_3477_n699,
         DP_OP_424J2_126_3477_n698, DP_OP_424J2_126_3477_n697,
         DP_OP_424J2_126_3477_n696, DP_OP_424J2_126_3477_n695,
         DP_OP_424J2_126_3477_n694, DP_OP_424J2_126_3477_n693,
         DP_OP_424J2_126_3477_n692, DP_OP_424J2_126_3477_n691,
         DP_OP_424J2_126_3477_n690, DP_OP_424J2_126_3477_n689,
         DP_OP_424J2_126_3477_n688, DP_OP_424J2_126_3477_n687,
         DP_OP_424J2_126_3477_n686, DP_OP_424J2_126_3477_n685,
         DP_OP_424J2_126_3477_n684, DP_OP_424J2_126_3477_n683,
         DP_OP_424J2_126_3477_n682, DP_OP_424J2_126_3477_n681,
         DP_OP_424J2_126_3477_n680, DP_OP_424J2_126_3477_n679,
         DP_OP_424J2_126_3477_n678, DP_OP_424J2_126_3477_n677,
         DP_OP_424J2_126_3477_n676, DP_OP_424J2_126_3477_n675,
         DP_OP_424J2_126_3477_n674, DP_OP_424J2_126_3477_n673,
         DP_OP_424J2_126_3477_n672, DP_OP_424J2_126_3477_n671,
         DP_OP_424J2_126_3477_n670, DP_OP_424J2_126_3477_n669,
         DP_OP_424J2_126_3477_n668, DP_OP_424J2_126_3477_n667,
         DP_OP_424J2_126_3477_n666, DP_OP_424J2_126_3477_n665,
         DP_OP_424J2_126_3477_n664, DP_OP_424J2_126_3477_n663,
         DP_OP_424J2_126_3477_n662, DP_OP_424J2_126_3477_n661,
         DP_OP_424J2_126_3477_n660, DP_OP_424J2_126_3477_n659,
         DP_OP_424J2_126_3477_n658, DP_OP_424J2_126_3477_n657,
         DP_OP_424J2_126_3477_n656, DP_OP_424J2_126_3477_n655,
         DP_OP_424J2_126_3477_n654, DP_OP_424J2_126_3477_n653,
         DP_OP_424J2_126_3477_n652, DP_OP_424J2_126_3477_n651,
         DP_OP_424J2_126_3477_n650, DP_OP_424J2_126_3477_n649,
         DP_OP_424J2_126_3477_n648, DP_OP_424J2_126_3477_n647,
         DP_OP_424J2_126_3477_n646, DP_OP_424J2_126_3477_n645,
         DP_OP_424J2_126_3477_n644, DP_OP_424J2_126_3477_n643,
         DP_OP_424J2_126_3477_n642, DP_OP_424J2_126_3477_n641,
         DP_OP_424J2_126_3477_n640, DP_OP_424J2_126_3477_n639,
         DP_OP_424J2_126_3477_n638, DP_OP_424J2_126_3477_n637,
         DP_OP_424J2_126_3477_n636, DP_OP_424J2_126_3477_n635,
         DP_OP_424J2_126_3477_n634, DP_OP_424J2_126_3477_n633,
         DP_OP_424J2_126_3477_n632, DP_OP_424J2_126_3477_n631,
         DP_OP_424J2_126_3477_n630, DP_OP_424J2_126_3477_n629,
         DP_OP_424J2_126_3477_n628, DP_OP_424J2_126_3477_n627,
         DP_OP_424J2_126_3477_n626, DP_OP_424J2_126_3477_n625,
         DP_OP_424J2_126_3477_n624, DP_OP_424J2_126_3477_n623,
         DP_OP_424J2_126_3477_n622, DP_OP_424J2_126_3477_n621,
         DP_OP_424J2_126_3477_n620, DP_OP_424J2_126_3477_n619,
         DP_OP_424J2_126_3477_n618, DP_OP_424J2_126_3477_n617,
         DP_OP_424J2_126_3477_n616, DP_OP_424J2_126_3477_n615,
         DP_OP_424J2_126_3477_n614, DP_OP_424J2_126_3477_n613,
         DP_OP_424J2_126_3477_n612, DP_OP_424J2_126_3477_n611,
         DP_OP_424J2_126_3477_n610, DP_OP_424J2_126_3477_n609,
         DP_OP_424J2_126_3477_n608, DP_OP_424J2_126_3477_n607,
         DP_OP_424J2_126_3477_n606, DP_OP_424J2_126_3477_n605,
         DP_OP_424J2_126_3477_n604, DP_OP_424J2_126_3477_n603,
         DP_OP_424J2_126_3477_n602, DP_OP_424J2_126_3477_n601,
         DP_OP_424J2_126_3477_n600, DP_OP_424J2_126_3477_n599,
         DP_OP_424J2_126_3477_n598, DP_OP_424J2_126_3477_n597,
         DP_OP_424J2_126_3477_n596, DP_OP_424J2_126_3477_n595,
         DP_OP_424J2_126_3477_n594, DP_OP_424J2_126_3477_n593,
         DP_OP_424J2_126_3477_n592, DP_OP_424J2_126_3477_n591,
         DP_OP_424J2_126_3477_n590, DP_OP_424J2_126_3477_n589,
         DP_OP_424J2_126_3477_n588, DP_OP_424J2_126_3477_n587,
         DP_OP_424J2_126_3477_n586, DP_OP_424J2_126_3477_n585,
         DP_OP_424J2_126_3477_n584, DP_OP_424J2_126_3477_n583,
         DP_OP_424J2_126_3477_n582, DP_OP_424J2_126_3477_n581,
         DP_OP_424J2_126_3477_n580, DP_OP_424J2_126_3477_n579,
         DP_OP_424J2_126_3477_n578, DP_OP_424J2_126_3477_n577,
         DP_OP_424J2_126_3477_n576, DP_OP_424J2_126_3477_n575,
         DP_OP_424J2_126_3477_n574, DP_OP_424J2_126_3477_n573,
         DP_OP_424J2_126_3477_n572, DP_OP_424J2_126_3477_n571,
         DP_OP_424J2_126_3477_n570, DP_OP_424J2_126_3477_n569,
         DP_OP_424J2_126_3477_n568, DP_OP_424J2_126_3477_n567,
         DP_OP_424J2_126_3477_n566, DP_OP_424J2_126_3477_n565,
         DP_OP_424J2_126_3477_n564, DP_OP_424J2_126_3477_n563,
         DP_OP_424J2_126_3477_n562, DP_OP_424J2_126_3477_n561,
         DP_OP_424J2_126_3477_n560, DP_OP_424J2_126_3477_n559,
         DP_OP_424J2_126_3477_n558, DP_OP_424J2_126_3477_n557,
         DP_OP_424J2_126_3477_n556, DP_OP_424J2_126_3477_n555,
         DP_OP_424J2_126_3477_n554, DP_OP_424J2_126_3477_n553,
         DP_OP_424J2_126_3477_n552, DP_OP_424J2_126_3477_n551,
         DP_OP_424J2_126_3477_n550, DP_OP_424J2_126_3477_n549,
         DP_OP_424J2_126_3477_n548, DP_OP_424J2_126_3477_n547,
         DP_OP_424J2_126_3477_n546, DP_OP_424J2_126_3477_n545,
         DP_OP_424J2_126_3477_n544, DP_OP_424J2_126_3477_n543,
         DP_OP_424J2_126_3477_n542, DP_OP_424J2_126_3477_n541,
         DP_OP_424J2_126_3477_n540, DP_OP_424J2_126_3477_n539,
         DP_OP_424J2_126_3477_n538, DP_OP_424J2_126_3477_n537,
         DP_OP_424J2_126_3477_n536, DP_OP_424J2_126_3477_n535,
         DP_OP_424J2_126_3477_n534, DP_OP_424J2_126_3477_n533,
         DP_OP_424J2_126_3477_n532, DP_OP_424J2_126_3477_n531,
         DP_OP_424J2_126_3477_n530, DP_OP_424J2_126_3477_n529,
         DP_OP_424J2_126_3477_n528, DP_OP_424J2_126_3477_n527,
         DP_OP_424J2_126_3477_n526, DP_OP_424J2_126_3477_n525,
         DP_OP_424J2_126_3477_n524, DP_OP_424J2_126_3477_n523,
         DP_OP_424J2_126_3477_n522, DP_OP_424J2_126_3477_n521,
         DP_OP_424J2_126_3477_n520, DP_OP_424J2_126_3477_n519,
         DP_OP_424J2_126_3477_n518, DP_OP_424J2_126_3477_n517,
         DP_OP_424J2_126_3477_n516, DP_OP_424J2_126_3477_n515,
         DP_OP_424J2_126_3477_n514, DP_OP_424J2_126_3477_n513,
         DP_OP_424J2_126_3477_n512, DP_OP_424J2_126_3477_n510,
         DP_OP_424J2_126_3477_n509, DP_OP_424J2_126_3477_n508,
         DP_OP_424J2_126_3477_n507, DP_OP_424J2_126_3477_n506,
         DP_OP_424J2_126_3477_n505, DP_OP_424J2_126_3477_n504,
         DP_OP_424J2_126_3477_n503, DP_OP_424J2_126_3477_n502,
         DP_OP_424J2_126_3477_n501, DP_OP_424J2_126_3477_n500,
         DP_OP_424J2_126_3477_n499, DP_OP_424J2_126_3477_n498,
         DP_OP_424J2_126_3477_n497, DP_OP_424J2_126_3477_n496,
         DP_OP_424J2_126_3477_n495, DP_OP_424J2_126_3477_n494,
         DP_OP_424J2_126_3477_n493, DP_OP_424J2_126_3477_n492,
         DP_OP_424J2_126_3477_n491, DP_OP_424J2_126_3477_n490,
         DP_OP_424J2_126_3477_n489, DP_OP_424J2_126_3477_n488,
         DP_OP_424J2_126_3477_n487, DP_OP_424J2_126_3477_n486,
         DP_OP_424J2_126_3477_n485, DP_OP_424J2_126_3477_n484,
         DP_OP_424J2_126_3477_n483, DP_OP_424J2_126_3477_n482,
         DP_OP_424J2_126_3477_n481, DP_OP_424J2_126_3477_n480,
         DP_OP_424J2_126_3477_n479, DP_OP_424J2_126_3477_n478,
         DP_OP_424J2_126_3477_n477, DP_OP_424J2_126_3477_n476,
         DP_OP_424J2_126_3477_n475, DP_OP_424J2_126_3477_n474,
         DP_OP_424J2_126_3477_n473, DP_OP_424J2_126_3477_n472,
         DP_OP_424J2_126_3477_n471, DP_OP_424J2_126_3477_n470,
         DP_OP_424J2_126_3477_n469, DP_OP_424J2_126_3477_n468,
         DP_OP_424J2_126_3477_n467, DP_OP_424J2_126_3477_n466,
         DP_OP_424J2_126_3477_n465, DP_OP_424J2_126_3477_n464,
         DP_OP_424J2_126_3477_n463, DP_OP_424J2_126_3477_n462,
         DP_OP_424J2_126_3477_n461, DP_OP_424J2_126_3477_n460,
         DP_OP_424J2_126_3477_n459, DP_OP_424J2_126_3477_n458,
         DP_OP_424J2_126_3477_n457, DP_OP_424J2_126_3477_n456,
         DP_OP_424J2_126_3477_n455, DP_OP_424J2_126_3477_n454,
         DP_OP_424J2_126_3477_n453, DP_OP_424J2_126_3477_n452,
         DP_OP_424J2_126_3477_n451, DP_OP_424J2_126_3477_n450,
         DP_OP_424J2_126_3477_n449, DP_OP_424J2_126_3477_n448,
         DP_OP_424J2_126_3477_n447, DP_OP_424J2_126_3477_n446,
         DP_OP_424J2_126_3477_n445, DP_OP_424J2_126_3477_n444,
         DP_OP_424J2_126_3477_n443, DP_OP_424J2_126_3477_n442,
         DP_OP_424J2_126_3477_n441, DP_OP_424J2_126_3477_n440,
         DP_OP_424J2_126_3477_n439, DP_OP_424J2_126_3477_n438,
         DP_OP_424J2_126_3477_n437, DP_OP_424J2_126_3477_n436,
         DP_OP_424J2_126_3477_n435, DP_OP_424J2_126_3477_n434,
         DP_OP_424J2_126_3477_n433, DP_OP_424J2_126_3477_n432,
         DP_OP_424J2_126_3477_n431, DP_OP_424J2_126_3477_n430,
         DP_OP_424J2_126_3477_n429, DP_OP_424J2_126_3477_n428,
         DP_OP_424J2_126_3477_n427, DP_OP_424J2_126_3477_n426,
         DP_OP_424J2_126_3477_n425, DP_OP_424J2_126_3477_n424,
         DP_OP_424J2_126_3477_n423, DP_OP_424J2_126_3477_n422,
         DP_OP_424J2_126_3477_n421, DP_OP_424J2_126_3477_n420,
         DP_OP_424J2_126_3477_n419, DP_OP_424J2_126_3477_n418,
         DP_OP_424J2_126_3477_n417, DP_OP_424J2_126_3477_n416,
         DP_OP_424J2_126_3477_n415, DP_OP_424J2_126_3477_n414,
         DP_OP_424J2_126_3477_n413, DP_OP_424J2_126_3477_n412,
         DP_OP_424J2_126_3477_n411, DP_OP_424J2_126_3477_n410,
         DP_OP_424J2_126_3477_n409, DP_OP_424J2_126_3477_n408,
         DP_OP_424J2_126_3477_n407, DP_OP_424J2_126_3477_n406,
         DP_OP_424J2_126_3477_n405, DP_OP_424J2_126_3477_n404,
         DP_OP_424J2_126_3477_n403, DP_OP_424J2_126_3477_n402,
         DP_OP_424J2_126_3477_n401, DP_OP_424J2_126_3477_n400,
         DP_OP_424J2_126_3477_n399, DP_OP_424J2_126_3477_n398,
         DP_OP_424J2_126_3477_n397, DP_OP_424J2_126_3477_n396,
         DP_OP_424J2_126_3477_n395, DP_OP_424J2_126_3477_n394,
         DP_OP_424J2_126_3477_n393, DP_OP_424J2_126_3477_n392,
         DP_OP_424J2_126_3477_n391, DP_OP_424J2_126_3477_n390,
         DP_OP_424J2_126_3477_n389, DP_OP_424J2_126_3477_n388,
         DP_OP_424J2_126_3477_n387, DP_OP_424J2_126_3477_n386,
         DP_OP_424J2_126_3477_n385, DP_OP_424J2_126_3477_n384,
         DP_OP_424J2_126_3477_n383, DP_OP_424J2_126_3477_n382,
         DP_OP_424J2_126_3477_n381, DP_OP_424J2_126_3477_n380,
         DP_OP_424J2_126_3477_n379, DP_OP_424J2_126_3477_n378,
         DP_OP_424J2_126_3477_n377, DP_OP_424J2_126_3477_n376,
         DP_OP_424J2_126_3477_n375, DP_OP_424J2_126_3477_n374,
         DP_OP_424J2_126_3477_n373, DP_OP_424J2_126_3477_n372,
         DP_OP_424J2_126_3477_n371, DP_OP_424J2_126_3477_n370,
         DP_OP_424J2_126_3477_n369, DP_OP_424J2_126_3477_n368,
         DP_OP_424J2_126_3477_n367, DP_OP_424J2_126_3477_n366,
         DP_OP_424J2_126_3477_n365, DP_OP_424J2_126_3477_n364,
         DP_OP_424J2_126_3477_n363, DP_OP_424J2_126_3477_n362,
         DP_OP_424J2_126_3477_n361, DP_OP_424J2_126_3477_n360,
         DP_OP_424J2_126_3477_n359, DP_OP_424J2_126_3477_n358,
         DP_OP_424J2_126_3477_n357, DP_OP_424J2_126_3477_n356,
         DP_OP_424J2_126_3477_n355, DP_OP_424J2_126_3477_n354,
         DP_OP_424J2_126_3477_n353, DP_OP_424J2_126_3477_n352,
         DP_OP_424J2_126_3477_n351, DP_OP_424J2_126_3477_n350,
         DP_OP_424J2_126_3477_n349, DP_OP_424J2_126_3477_n348,
         DP_OP_424J2_126_3477_n347, DP_OP_424J2_126_3477_n346,
         DP_OP_424J2_126_3477_n345, DP_OP_424J2_126_3477_n344,
         DP_OP_424J2_126_3477_n343, DP_OP_424J2_126_3477_n342,
         DP_OP_424J2_126_3477_n341, DP_OP_424J2_126_3477_n340,
         DP_OP_424J2_126_3477_n339, DP_OP_424J2_126_3477_n338,
         DP_OP_424J2_126_3477_n337, DP_OP_424J2_126_3477_n336,
         DP_OP_424J2_126_3477_n335, DP_OP_424J2_126_3477_n334,
         DP_OP_424J2_126_3477_n333, DP_OP_424J2_126_3477_n332,
         DP_OP_424J2_126_3477_n331, DP_OP_424J2_126_3477_n330,
         DP_OP_424J2_126_3477_n329, DP_OP_424J2_126_3477_n328,
         DP_OP_424J2_126_3477_n327, DP_OP_424J2_126_3477_n326,
         DP_OP_424J2_126_3477_n325, DP_OP_424J2_126_3477_n324,
         DP_OP_424J2_126_3477_n323, DP_OP_424J2_126_3477_n322,
         DP_OP_424J2_126_3477_n320, DP_OP_424J2_126_3477_n319,
         DP_OP_424J2_126_3477_n318, DP_OP_424J2_126_3477_n317,
         DP_OP_424J2_126_3477_n316, DP_OP_424J2_126_3477_n315,
         DP_OP_424J2_126_3477_n314, DP_OP_424J2_126_3477_n313,
         DP_OP_424J2_126_3477_n312, DP_OP_424J2_126_3477_n311,
         DP_OP_424J2_126_3477_n310, DP_OP_424J2_126_3477_n309,
         DP_OP_424J2_126_3477_n308, DP_OP_424J2_126_3477_n307,
         DP_OP_424J2_126_3477_n306, DP_OP_424J2_126_3477_n305,
         DP_OP_424J2_126_3477_n304, DP_OP_424J2_126_3477_n303,
         DP_OP_424J2_126_3477_n302, DP_OP_424J2_126_3477_n297,
         DP_OP_424J2_126_3477_n295, DP_OP_424J2_126_3477_n287,
         DP_OP_424J2_126_3477_n286, DP_OP_424J2_126_3477_n285,
         DP_OP_424J2_126_3477_n284, DP_OP_424J2_126_3477_n283,
         DP_OP_424J2_126_3477_n282, DP_OP_424J2_126_3477_n281,
         DP_OP_424J2_126_3477_n280, DP_OP_424J2_126_3477_n279,
         DP_OP_424J2_126_3477_n277, DP_OP_424J2_126_3477_n276,
         DP_OP_424J2_126_3477_n274, DP_OP_424J2_126_3477_n272,
         DP_OP_424J2_126_3477_n269, DP_OP_424J2_126_3477_n268,
         DP_OP_424J2_126_3477_n267, DP_OP_424J2_126_3477_n266,
         DP_OP_424J2_126_3477_n265, DP_OP_424J2_126_3477_n261,
         DP_OP_424J2_126_3477_n260, DP_OP_424J2_126_3477_n259,
         DP_OP_424J2_126_3477_n257, DP_OP_424J2_126_3477_n252,
         DP_OP_424J2_126_3477_n250, DP_OP_424J2_126_3477_n249,
         DP_OP_424J2_126_3477_n245, DP_OP_424J2_126_3477_n244,
         DP_OP_424J2_126_3477_n240, DP_OP_424J2_126_3477_n237,
         DP_OP_424J2_126_3477_n236, DP_OP_424J2_126_3477_n233,
         DP_OP_424J2_126_3477_n226, DP_OP_424J2_126_3477_n220,
         DP_OP_424J2_126_3477_n219, DP_OP_424J2_126_3477_n217,
         DP_OP_424J2_126_3477_n214, DP_OP_424J2_126_3477_n213,
         DP_OP_424J2_126_3477_n212, DP_OP_424J2_126_3477_n210,
         DP_OP_424J2_126_3477_n209, DP_OP_424J2_126_3477_n203,
         DP_OP_424J2_126_3477_n202, DP_OP_424J2_126_3477_n201,
         DP_OP_424J2_126_3477_n198, DP_OP_424J2_126_3477_n197,
         DP_OP_424J2_126_3477_n190, DP_OP_424J2_126_3477_n189,
         DP_OP_424J2_126_3477_n187, DP_OP_424J2_126_3477_n185,
         DP_OP_424J2_126_3477_n182, DP_OP_424J2_126_3477_n178,
         DP_OP_424J2_126_3477_n176, DP_OP_424J2_126_3477_n174,
         DP_OP_424J2_126_3477_n171, DP_OP_424J2_126_3477_n167,
         DP_OP_424J2_126_3477_n166, DP_OP_424J2_126_3477_n165,
         DP_OP_424J2_126_3477_n162, DP_OP_424J2_126_3477_n160,
         DP_OP_424J2_126_3477_n156, DP_OP_424J2_126_3477_n153,
         DP_OP_424J2_126_3477_n151, DP_OP_424J2_126_3477_n149,
         DP_OP_424J2_126_3477_n148, DP_OP_424J2_126_3477_n146,
         DP_OP_424J2_126_3477_n145, DP_OP_424J2_126_3477_n144,
         DP_OP_424J2_126_3477_n142, DP_OP_424J2_126_3477_n141,
         DP_OP_424J2_126_3477_n140, DP_OP_424J2_126_3477_n138,
         DP_OP_424J2_126_3477_n136, DP_OP_424J2_126_3477_n133,
         DP_OP_424J2_126_3477_n132, DP_OP_424J2_126_3477_n131,
         DP_OP_424J2_126_3477_n129, DP_OP_424J2_126_3477_n128,
         DP_OP_424J2_126_3477_n127, DP_OP_424J2_126_3477_n126,
         DP_OP_424J2_126_3477_n124, DP_OP_424J2_126_3477_n122,
         DP_OP_424J2_126_3477_n120, DP_OP_424J2_126_3477_n115,
         DP_OP_424J2_126_3477_n114, DP_OP_424J2_126_3477_n111,
         DP_OP_424J2_126_3477_n110, DP_OP_424J2_126_3477_n109,
         DP_OP_424J2_126_3477_n107, DP_OP_424J2_126_3477_n105,
         DP_OP_424J2_126_3477_n102, DP_OP_424J2_126_3477_n100,
         DP_OP_424J2_126_3477_n98, DP_OP_424J2_126_3477_n97,
         DP_OP_424J2_126_3477_n96, DP_OP_424J2_126_3477_n95,
         DP_OP_424J2_126_3477_n93, DP_OP_424J2_126_3477_n91,
         DP_OP_424J2_126_3477_n89, DP_OP_424J2_126_3477_n85,
         DP_OP_424J2_126_3477_n82, DP_OP_424J2_126_3477_n80,
         DP_OP_424J2_126_3477_n78, DP_OP_424J2_126_3477_n77,
         DP_OP_424J2_126_3477_n75, DP_OP_424J2_126_3477_n73,
         DP_OP_424J2_126_3477_n72, DP_OP_424J2_126_3477_n71,
         DP_OP_424J2_126_3477_n69, DP_OP_424J2_126_3477_n67,
         DP_OP_424J2_126_3477_n65, DP_OP_424J2_126_3477_n60,
         DP_OP_424J2_126_3477_n58, DP_OP_424J2_126_3477_n57,
         DP_OP_424J2_126_3477_n56, DP_OP_424J2_126_3477_n54,
         DP_OP_424J2_126_3477_n52, DP_OP_424J2_126_3477_n51,
         DP_OP_424J2_126_3477_n50, DP_OP_424J2_126_3477_n49,
         DP_OP_424J2_126_3477_n47, DP_OP_424J2_126_3477_n38,
         DP_OP_424J2_126_3477_n22, DP_OP_424J2_126_3477_n19,
         DP_OP_424J2_126_3477_n17, DP_OP_424J2_126_3477_n15,
         DP_OP_424J2_126_3477_n13, DP_OP_424J2_126_3477_n5,
         DP_OP_423J2_125_3477_n3066, DP_OP_423J2_125_3477_n3065,
         DP_OP_423J2_125_3477_n3063, DP_OP_423J2_125_3477_n3062,
         DP_OP_423J2_125_3477_n3061, DP_OP_423J2_125_3477_n3060,
         DP_OP_423J2_125_3477_n3059, DP_OP_423J2_125_3477_n3057,
         DP_OP_423J2_125_3477_n3056, DP_OP_423J2_125_3477_n3055,
         DP_OP_423J2_125_3477_n3054, DP_OP_423J2_125_3477_n3053,
         DP_OP_423J2_125_3477_n3052, DP_OP_423J2_125_3477_n3051,
         DP_OP_423J2_125_3477_n3050, DP_OP_423J2_125_3477_n3049,
         DP_OP_423J2_125_3477_n3048, DP_OP_423J2_125_3477_n3047,
         DP_OP_423J2_125_3477_n3046, DP_OP_423J2_125_3477_n3045,
         DP_OP_423J2_125_3477_n3044, DP_OP_423J2_125_3477_n3043,
         DP_OP_423J2_125_3477_n3042, DP_OP_423J2_125_3477_n3041,
         DP_OP_423J2_125_3477_n3040, DP_OP_423J2_125_3477_n3039,
         DP_OP_423J2_125_3477_n3038, DP_OP_423J2_125_3477_n3037,
         DP_OP_423J2_125_3477_n3036, DP_OP_423J2_125_3477_n3035,
         DP_OP_423J2_125_3477_n3034, DP_OP_423J2_125_3477_n3033,
         DP_OP_423J2_125_3477_n3032, DP_OP_423J2_125_3477_n3031,
         DP_OP_423J2_125_3477_n3030, DP_OP_423J2_125_3477_n3029,
         DP_OP_423J2_125_3477_n3028, DP_OP_423J2_125_3477_n3027,
         DP_OP_423J2_125_3477_n3026, DP_OP_423J2_125_3477_n3025,
         DP_OP_423J2_125_3477_n3022, DP_OP_423J2_125_3477_n3021,
         DP_OP_423J2_125_3477_n3019, DP_OP_423J2_125_3477_n3014,
         DP_OP_423J2_125_3477_n3013, DP_OP_423J2_125_3477_n3012,
         DP_OP_423J2_125_3477_n3011, DP_OP_423J2_125_3477_n3010,
         DP_OP_423J2_125_3477_n3009, DP_OP_423J2_125_3477_n3008,
         DP_OP_423J2_125_3477_n3007, DP_OP_423J2_125_3477_n3006,
         DP_OP_423J2_125_3477_n3005, DP_OP_423J2_125_3477_n3003,
         DP_OP_423J2_125_3477_n3002, DP_OP_423J2_125_3477_n3001,
         DP_OP_423J2_125_3477_n3000, DP_OP_423J2_125_3477_n2999,
         DP_OP_423J2_125_3477_n2998, DP_OP_423J2_125_3477_n2997,
         DP_OP_423J2_125_3477_n2996, DP_OP_423J2_125_3477_n2995,
         DP_OP_423J2_125_3477_n2994, DP_OP_423J2_125_3477_n2993,
         DP_OP_423J2_125_3477_n2992, DP_OP_423J2_125_3477_n2991,
         DP_OP_423J2_125_3477_n2990, DP_OP_423J2_125_3477_n2989,
         DP_OP_423J2_125_3477_n2988, DP_OP_423J2_125_3477_n2987,
         DP_OP_423J2_125_3477_n2986, DP_OP_423J2_125_3477_n2985,
         DP_OP_423J2_125_3477_n2984, DP_OP_423J2_125_3477_n2983,
         DP_OP_423J2_125_3477_n2982, DP_OP_423J2_125_3477_n2976,
         DP_OP_423J2_125_3477_n2973, DP_OP_423J2_125_3477_n2969,
         DP_OP_423J2_125_3477_n2968, DP_OP_423J2_125_3477_n2967,
         DP_OP_423J2_125_3477_n2966, DP_OP_423J2_125_3477_n2965,
         DP_OP_423J2_125_3477_n2964, DP_OP_423J2_125_3477_n2963,
         DP_OP_423J2_125_3477_n2962, DP_OP_423J2_125_3477_n2961,
         DP_OP_423J2_125_3477_n2960, DP_OP_423J2_125_3477_n2959,
         DP_OP_423J2_125_3477_n2958, DP_OP_423J2_125_3477_n2957,
         DP_OP_423J2_125_3477_n2956, DP_OP_423J2_125_3477_n2955,
         DP_OP_423J2_125_3477_n2954, DP_OP_423J2_125_3477_n2953,
         DP_OP_423J2_125_3477_n2952, DP_OP_423J2_125_3477_n2951,
         DP_OP_423J2_125_3477_n2950, DP_OP_423J2_125_3477_n2949,
         DP_OP_423J2_125_3477_n2948, DP_OP_423J2_125_3477_n2947,
         DP_OP_423J2_125_3477_n2946, DP_OP_423J2_125_3477_n2945,
         DP_OP_423J2_125_3477_n2944, DP_OP_423J2_125_3477_n2943,
         DP_OP_423J2_125_3477_n2942, DP_OP_423J2_125_3477_n2941,
         DP_OP_423J2_125_3477_n2940, DP_OP_423J2_125_3477_n2939,
         DP_OP_423J2_125_3477_n2938, DP_OP_423J2_125_3477_n2936,
         DP_OP_423J2_125_3477_n2932, DP_OP_423J2_125_3477_n2931,
         DP_OP_423J2_125_3477_n2925, DP_OP_423J2_125_3477_n2924,
         DP_OP_423J2_125_3477_n2923, DP_OP_423J2_125_3477_n2922,
         DP_OP_423J2_125_3477_n2921, DP_OP_423J2_125_3477_n2920,
         DP_OP_423J2_125_3477_n2919, DP_OP_423J2_125_3477_n2918,
         DP_OP_423J2_125_3477_n2917, DP_OP_423J2_125_3477_n2916,
         DP_OP_423J2_125_3477_n2915, DP_OP_423J2_125_3477_n2914,
         DP_OP_423J2_125_3477_n2913, DP_OP_423J2_125_3477_n2912,
         DP_OP_423J2_125_3477_n2911, DP_OP_423J2_125_3477_n2910,
         DP_OP_423J2_125_3477_n2909, DP_OP_423J2_125_3477_n2908,
         DP_OP_423J2_125_3477_n2907, DP_OP_423J2_125_3477_n2906,
         DP_OP_423J2_125_3477_n2905, DP_OP_423J2_125_3477_n2904,
         DP_OP_423J2_125_3477_n2903, DP_OP_423J2_125_3477_n2902,
         DP_OP_423J2_125_3477_n2900, DP_OP_423J2_125_3477_n2899,
         DP_OP_423J2_125_3477_n2898, DP_OP_423J2_125_3477_n2897,
         DP_OP_423J2_125_3477_n2896, DP_OP_423J2_125_3477_n2895,
         DP_OP_423J2_125_3477_n2894, DP_OP_423J2_125_3477_n2892,
         DP_OP_423J2_125_3477_n2891, DP_OP_423J2_125_3477_n2890,
         DP_OP_423J2_125_3477_n2889, DP_OP_423J2_125_3477_n2887,
         DP_OP_423J2_125_3477_n2886, DP_OP_423J2_125_3477_n2881,
         DP_OP_423J2_125_3477_n2880, DP_OP_423J2_125_3477_n2879,
         DP_OP_423J2_125_3477_n2878, DP_OP_423J2_125_3477_n2877,
         DP_OP_423J2_125_3477_n2876, DP_OP_423J2_125_3477_n2875,
         DP_OP_423J2_125_3477_n2874, DP_OP_423J2_125_3477_n2873,
         DP_OP_423J2_125_3477_n2871, DP_OP_423J2_125_3477_n2870,
         DP_OP_423J2_125_3477_n2869, DP_OP_423J2_125_3477_n2868,
         DP_OP_423J2_125_3477_n2867, DP_OP_423J2_125_3477_n2866,
         DP_OP_423J2_125_3477_n2864, DP_OP_423J2_125_3477_n2863,
         DP_OP_423J2_125_3477_n2862, DP_OP_423J2_125_3477_n2861,
         DP_OP_423J2_125_3477_n2860, DP_OP_423J2_125_3477_n2859,
         DP_OP_423J2_125_3477_n2858, DP_OP_423J2_125_3477_n2857,
         DP_OP_423J2_125_3477_n2856, DP_OP_423J2_125_3477_n2855,
         DP_OP_423J2_125_3477_n2854, DP_OP_423J2_125_3477_n2853,
         DP_OP_423J2_125_3477_n2852, DP_OP_423J2_125_3477_n2851,
         DP_OP_423J2_125_3477_n2850, DP_OP_423J2_125_3477_n2849,
         DP_OP_423J2_125_3477_n2845, DP_OP_423J2_125_3477_n2844,
         DP_OP_423J2_125_3477_n2843, DP_OP_423J2_125_3477_n2842,
         DP_OP_423J2_125_3477_n2841, DP_OP_423J2_125_3477_n2837,
         DP_OP_423J2_125_3477_n2836, DP_OP_423J2_125_3477_n2835,
         DP_OP_423J2_125_3477_n2834, DP_OP_423J2_125_3477_n2833,
         DP_OP_423J2_125_3477_n2832, DP_OP_423J2_125_3477_n2831,
         DP_OP_423J2_125_3477_n2830, DP_OP_423J2_125_3477_n2829,
         DP_OP_423J2_125_3477_n2828, DP_OP_423J2_125_3477_n2827,
         DP_OP_423J2_125_3477_n2826, DP_OP_423J2_125_3477_n2825,
         DP_OP_423J2_125_3477_n2824, DP_OP_423J2_125_3477_n2823,
         DP_OP_423J2_125_3477_n2822, DP_OP_423J2_125_3477_n2821,
         DP_OP_423J2_125_3477_n2820, DP_OP_423J2_125_3477_n2819,
         DP_OP_423J2_125_3477_n2818, DP_OP_423J2_125_3477_n2817,
         DP_OP_423J2_125_3477_n2816, DP_OP_423J2_125_3477_n2815,
         DP_OP_423J2_125_3477_n2814, DP_OP_423J2_125_3477_n2813,
         DP_OP_423J2_125_3477_n2812, DP_OP_423J2_125_3477_n2811,
         DP_OP_423J2_125_3477_n2810, DP_OP_423J2_125_3477_n2809,
         DP_OP_423J2_125_3477_n2808, DP_OP_423J2_125_3477_n2807,
         DP_OP_423J2_125_3477_n2806, DP_OP_423J2_125_3477_n2805,
         DP_OP_423J2_125_3477_n2804, DP_OP_423J2_125_3477_n2803,
         DP_OP_423J2_125_3477_n2802, DP_OP_423J2_125_3477_n2801,
         DP_OP_423J2_125_3477_n2800, DP_OP_423J2_125_3477_n2799,
         DP_OP_423J2_125_3477_n2798, DP_OP_423J2_125_3477_n2795,
         DP_OP_423J2_125_3477_n2794, DP_OP_423J2_125_3477_n2793,
         DP_OP_423J2_125_3477_n2792, DP_OP_423J2_125_3477_n2791,
         DP_OP_423J2_125_3477_n2790, DP_OP_423J2_125_3477_n2789,
         DP_OP_423J2_125_3477_n2788, DP_OP_423J2_125_3477_n2787,
         DP_OP_423J2_125_3477_n2786, DP_OP_423J2_125_3477_n2785,
         DP_OP_423J2_125_3477_n2784, DP_OP_423J2_125_3477_n2783,
         DP_OP_423J2_125_3477_n2782, DP_OP_423J2_125_3477_n2781,
         DP_OP_423J2_125_3477_n2780, DP_OP_423J2_125_3477_n2779,
         DP_OP_423J2_125_3477_n2778, DP_OP_423J2_125_3477_n2777,
         DP_OP_423J2_125_3477_n2776, DP_OP_423J2_125_3477_n2775,
         DP_OP_423J2_125_3477_n2774, DP_OP_423J2_125_3477_n2773,
         DP_OP_423J2_125_3477_n2772, DP_OP_423J2_125_3477_n2771,
         DP_OP_423J2_125_3477_n2770, DP_OP_423J2_125_3477_n2768,
         DP_OP_423J2_125_3477_n2767, DP_OP_423J2_125_3477_n2766,
         DP_OP_423J2_125_3477_n2765, DP_OP_423J2_125_3477_n2764,
         DP_OP_423J2_125_3477_n2763, DP_OP_423J2_125_3477_n2762,
         DP_OP_423J2_125_3477_n2758, DP_OP_423J2_125_3477_n2757,
         DP_OP_423J2_125_3477_n2756, DP_OP_423J2_125_3477_n2754,
         DP_OP_423J2_125_3477_n2751, DP_OP_423J2_125_3477_n2750,
         DP_OP_423J2_125_3477_n2749, DP_OP_423J2_125_3477_n2748,
         DP_OP_423J2_125_3477_n2746, DP_OP_423J2_125_3477_n2745,
         DP_OP_423J2_125_3477_n2744, DP_OP_423J2_125_3477_n2743,
         DP_OP_423J2_125_3477_n2742, DP_OP_423J2_125_3477_n2741,
         DP_OP_423J2_125_3477_n2740, DP_OP_423J2_125_3477_n2739,
         DP_OP_423J2_125_3477_n2738, DP_OP_423J2_125_3477_n2737,
         DP_OP_423J2_125_3477_n2736, DP_OP_423J2_125_3477_n2735,
         DP_OP_423J2_125_3477_n2734, DP_OP_423J2_125_3477_n2733,
         DP_OP_423J2_125_3477_n2732, DP_OP_423J2_125_3477_n2731,
         DP_OP_423J2_125_3477_n2730, DP_OP_423J2_125_3477_n2729,
         DP_OP_423J2_125_3477_n2728, DP_OP_423J2_125_3477_n2727,
         DP_OP_423J2_125_3477_n2726, DP_OP_423J2_125_3477_n2725,
         DP_OP_423J2_125_3477_n2724, DP_OP_423J2_125_3477_n2723,
         DP_OP_423J2_125_3477_n2722, DP_OP_423J2_125_3477_n2721,
         DP_OP_423J2_125_3477_n2720, DP_OP_423J2_125_3477_n2719,
         DP_OP_423J2_125_3477_n2718, DP_OP_423J2_125_3477_n2713,
         DP_OP_423J2_125_3477_n2712, DP_OP_423J2_125_3477_n2708,
         DP_OP_423J2_125_3477_n2706, DP_OP_423J2_125_3477_n2705,
         DP_OP_423J2_125_3477_n2704, DP_OP_423J2_125_3477_n2703,
         DP_OP_423J2_125_3477_n2702, DP_OP_423J2_125_3477_n2701,
         DP_OP_423J2_125_3477_n2700, DP_OP_423J2_125_3477_n2699,
         DP_OP_423J2_125_3477_n2698, DP_OP_423J2_125_3477_n2697,
         DP_OP_423J2_125_3477_n2696, DP_OP_423J2_125_3477_n2695,
         DP_OP_423J2_125_3477_n2694, DP_OP_423J2_125_3477_n2693,
         DP_OP_423J2_125_3477_n2692, DP_OP_423J2_125_3477_n2691,
         DP_OP_423J2_125_3477_n2690, DP_OP_423J2_125_3477_n2689,
         DP_OP_423J2_125_3477_n2688, DP_OP_423J2_125_3477_n2687,
         DP_OP_423J2_125_3477_n2686, DP_OP_423J2_125_3477_n2685,
         DP_OP_423J2_125_3477_n2684, DP_OP_423J2_125_3477_n2683,
         DP_OP_423J2_125_3477_n2682, DP_OP_423J2_125_3477_n2681,
         DP_OP_423J2_125_3477_n2680, DP_OP_423J2_125_3477_n2679,
         DP_OP_423J2_125_3477_n2678, DP_OP_423J2_125_3477_n2677,
         DP_OP_423J2_125_3477_n2676, DP_OP_423J2_125_3477_n2675,
         DP_OP_423J2_125_3477_n2674, DP_OP_423J2_125_3477_n2669,
         DP_OP_423J2_125_3477_n2668, DP_OP_423J2_125_3477_n2667,
         DP_OP_423J2_125_3477_n2666, DP_OP_423J2_125_3477_n2665,
         DP_OP_423J2_125_3477_n2661, DP_OP_423J2_125_3477_n2660,
         DP_OP_423J2_125_3477_n2659, DP_OP_423J2_125_3477_n2658,
         DP_OP_423J2_125_3477_n2657, DP_OP_423J2_125_3477_n2656,
         DP_OP_423J2_125_3477_n2655, DP_OP_423J2_125_3477_n2654,
         DP_OP_423J2_125_3477_n2653, DP_OP_423J2_125_3477_n2652,
         DP_OP_423J2_125_3477_n2651, DP_OP_423J2_125_3477_n2650,
         DP_OP_423J2_125_3477_n2649, DP_OP_423J2_125_3477_n2648,
         DP_OP_423J2_125_3477_n2647, DP_OP_423J2_125_3477_n2646,
         DP_OP_423J2_125_3477_n2645, DP_OP_423J2_125_3477_n2644,
         DP_OP_423J2_125_3477_n2643, DP_OP_423J2_125_3477_n2642,
         DP_OP_423J2_125_3477_n2641, DP_OP_423J2_125_3477_n2640,
         DP_OP_423J2_125_3477_n2639, DP_OP_423J2_125_3477_n2638,
         DP_OP_423J2_125_3477_n2637, DP_OP_423J2_125_3477_n2636,
         DP_OP_423J2_125_3477_n2635, DP_OP_423J2_125_3477_n2634,
         DP_OP_423J2_125_3477_n2633, DP_OP_423J2_125_3477_n2632,
         DP_OP_423J2_125_3477_n2631, DP_OP_423J2_125_3477_n2630,
         DP_OP_423J2_125_3477_n2629, DP_OP_423J2_125_3477_n2627,
         DP_OP_423J2_125_3477_n2625, DP_OP_423J2_125_3477_n2624,
         DP_OP_423J2_125_3477_n2623, DP_OP_423J2_125_3477_n2622,
         DP_OP_423J2_125_3477_n2621, DP_OP_423J2_125_3477_n2620,
         DP_OP_423J2_125_3477_n2619, DP_OP_423J2_125_3477_n2618,
         DP_OP_423J2_125_3477_n2617, DP_OP_423J2_125_3477_n2616,
         DP_OP_423J2_125_3477_n2615, DP_OP_423J2_125_3477_n2614,
         DP_OP_423J2_125_3477_n2613, DP_OP_423J2_125_3477_n2612,
         DP_OP_423J2_125_3477_n2611, DP_OP_423J2_125_3477_n2610,
         DP_OP_423J2_125_3477_n2609, DP_OP_423J2_125_3477_n2608,
         DP_OP_423J2_125_3477_n2607, DP_OP_423J2_125_3477_n2606,
         DP_OP_423J2_125_3477_n2605, DP_OP_423J2_125_3477_n2604,
         DP_OP_423J2_125_3477_n2603, DP_OP_423J2_125_3477_n2602,
         DP_OP_423J2_125_3477_n2601, DP_OP_423J2_125_3477_n2600,
         DP_OP_423J2_125_3477_n2599, DP_OP_423J2_125_3477_n2598,
         DP_OP_423J2_125_3477_n2597, DP_OP_423J2_125_3477_n2596,
         DP_OP_423J2_125_3477_n2595, DP_OP_423J2_125_3477_n2594,
         DP_OP_423J2_125_3477_n2593, DP_OP_423J2_125_3477_n2592,
         DP_OP_423J2_125_3477_n2591, DP_OP_423J2_125_3477_n2590,
         DP_OP_423J2_125_3477_n2589, DP_OP_423J2_125_3477_n2588,
         DP_OP_423J2_125_3477_n2587, DP_OP_423J2_125_3477_n2586,
         DP_OP_423J2_125_3477_n2585, DP_OP_423J2_125_3477_n2581,
         DP_OP_423J2_125_3477_n2579, DP_OP_423J2_125_3477_n2573,
         DP_OP_423J2_125_3477_n2572, DP_OP_423J2_125_3477_n2571,
         DP_OP_423J2_125_3477_n2570, DP_OP_423J2_125_3477_n2569,
         DP_OP_423J2_125_3477_n2568, DP_OP_423J2_125_3477_n2567,
         DP_OP_423J2_125_3477_n2566, DP_OP_423J2_125_3477_n2565,
         DP_OP_423J2_125_3477_n2564, DP_OP_423J2_125_3477_n2563,
         DP_OP_423J2_125_3477_n2562, DP_OP_423J2_125_3477_n2561,
         DP_OP_423J2_125_3477_n2560, DP_OP_423J2_125_3477_n2559,
         DP_OP_423J2_125_3477_n2558, DP_OP_423J2_125_3477_n2557,
         DP_OP_423J2_125_3477_n2556, DP_OP_423J2_125_3477_n2555,
         DP_OP_423J2_125_3477_n2554, DP_OP_423J2_125_3477_n2553,
         DP_OP_423J2_125_3477_n2552, DP_OP_423J2_125_3477_n2551,
         DP_OP_423J2_125_3477_n2550, DP_OP_423J2_125_3477_n2549,
         DP_OP_423J2_125_3477_n2548, DP_OP_423J2_125_3477_n2547,
         DP_OP_423J2_125_3477_n2546, DP_OP_423J2_125_3477_n2545,
         DP_OP_423J2_125_3477_n2544, DP_OP_423J2_125_3477_n2543,
         DP_OP_423J2_125_3477_n2542, DP_OP_423J2_125_3477_n2538,
         DP_OP_423J2_125_3477_n2537, DP_OP_423J2_125_3477_n2536,
         DP_OP_423J2_125_3477_n2531, DP_OP_423J2_125_3477_n2529,
         DP_OP_423J2_125_3477_n2528, DP_OP_423J2_125_3477_n2526,
         DP_OP_423J2_125_3477_n2525, DP_OP_423J2_125_3477_n2524,
         DP_OP_423J2_125_3477_n2523, DP_OP_423J2_125_3477_n2522,
         DP_OP_423J2_125_3477_n2521, DP_OP_423J2_125_3477_n2520,
         DP_OP_423J2_125_3477_n2519, DP_OP_423J2_125_3477_n2518,
         DP_OP_423J2_125_3477_n2517, DP_OP_423J2_125_3477_n2516,
         DP_OP_423J2_125_3477_n2515, DP_OP_423J2_125_3477_n2514,
         DP_OP_423J2_125_3477_n2513, DP_OP_423J2_125_3477_n2512,
         DP_OP_423J2_125_3477_n2511, DP_OP_423J2_125_3477_n2510,
         DP_OP_423J2_125_3477_n2509, DP_OP_423J2_125_3477_n2508,
         DP_OP_423J2_125_3477_n2507, DP_OP_423J2_125_3477_n2506,
         DP_OP_423J2_125_3477_n2505, DP_OP_423J2_125_3477_n2504,
         DP_OP_423J2_125_3477_n2503, DP_OP_423J2_125_3477_n2502,
         DP_OP_423J2_125_3477_n2501, DP_OP_423J2_125_3477_n2500,
         DP_OP_423J2_125_3477_n2499, DP_OP_423J2_125_3477_n2498,
         DP_OP_423J2_125_3477_n2496, DP_OP_423J2_125_3477_n2493,
         DP_OP_423J2_125_3477_n2485, DP_OP_423J2_125_3477_n2484,
         DP_OP_423J2_125_3477_n2483, DP_OP_423J2_125_3477_n2482,
         DP_OP_423J2_125_3477_n2481, DP_OP_423J2_125_3477_n2480,
         DP_OP_423J2_125_3477_n2479, DP_OP_423J2_125_3477_n2478,
         DP_OP_423J2_125_3477_n2477, DP_OP_423J2_125_3477_n2476,
         DP_OP_423J2_125_3477_n2475, DP_OP_423J2_125_3477_n2474,
         DP_OP_423J2_125_3477_n2473, DP_OP_423J2_125_3477_n2472,
         DP_OP_423J2_125_3477_n2471, DP_OP_423J2_125_3477_n2470,
         DP_OP_423J2_125_3477_n2469, DP_OP_423J2_125_3477_n2468,
         DP_OP_423J2_125_3477_n2467, DP_OP_423J2_125_3477_n2466,
         DP_OP_423J2_125_3477_n2465, DP_OP_423J2_125_3477_n2464,
         DP_OP_423J2_125_3477_n2463, DP_OP_423J2_125_3477_n2462,
         DP_OP_423J2_125_3477_n2461, DP_OP_423J2_125_3477_n2460,
         DP_OP_423J2_125_3477_n2459, DP_OP_423J2_125_3477_n2458,
         DP_OP_423J2_125_3477_n2457, DP_OP_423J2_125_3477_n2456,
         DP_OP_423J2_125_3477_n2455, DP_OP_423J2_125_3477_n2454,
         DP_OP_423J2_125_3477_n2452, DP_OP_423J2_125_3477_n2448,
         DP_OP_423J2_125_3477_n2447, DP_OP_423J2_125_3477_n2441,
         DP_OP_423J2_125_3477_n2440, DP_OP_423J2_125_3477_n2439,
         DP_OP_423J2_125_3477_n2438, DP_OP_423J2_125_3477_n2437,
         DP_OP_423J2_125_3477_n2436, DP_OP_423J2_125_3477_n2435,
         DP_OP_423J2_125_3477_n2434, DP_OP_423J2_125_3477_n2433,
         DP_OP_423J2_125_3477_n2432, DP_OP_423J2_125_3477_n2431,
         DP_OP_423J2_125_3477_n2430, DP_OP_423J2_125_3477_n2429,
         DP_OP_423J2_125_3477_n2428, DP_OP_423J2_125_3477_n2427,
         DP_OP_423J2_125_3477_n2426, DP_OP_423J2_125_3477_n2425,
         DP_OP_423J2_125_3477_n2424, DP_OP_423J2_125_3477_n2423,
         DP_OP_423J2_125_3477_n2422, DP_OP_423J2_125_3477_n2421,
         DP_OP_423J2_125_3477_n2420, DP_OP_423J2_125_3477_n2419,
         DP_OP_423J2_125_3477_n2418, DP_OP_423J2_125_3477_n2417,
         DP_OP_423J2_125_3477_n2416, DP_OP_423J2_125_3477_n2415,
         DP_OP_423J2_125_3477_n2414, DP_OP_423J2_125_3477_n2413,
         DP_OP_423J2_125_3477_n2412, DP_OP_423J2_125_3477_n2411,
         DP_OP_423J2_125_3477_n2410, DP_OP_423J2_125_3477_n2409,
         DP_OP_423J2_125_3477_n2405, DP_OP_423J2_125_3477_n2404,
         DP_OP_423J2_125_3477_n2401, DP_OP_423J2_125_3477_n2400,
         DP_OP_423J2_125_3477_n2399, DP_OP_423J2_125_3477_n2397,
         DP_OP_423J2_125_3477_n2396, DP_OP_423J2_125_3477_n2395,
         DP_OP_423J2_125_3477_n2394, DP_OP_423J2_125_3477_n2393,
         DP_OP_423J2_125_3477_n2392, DP_OP_423J2_125_3477_n2391,
         DP_OP_423J2_125_3477_n2390, DP_OP_423J2_125_3477_n2389,
         DP_OP_423J2_125_3477_n2388, DP_OP_423J2_125_3477_n2387,
         DP_OP_423J2_125_3477_n2386, DP_OP_423J2_125_3477_n2385,
         DP_OP_423J2_125_3477_n2384, DP_OP_423J2_125_3477_n2383,
         DP_OP_423J2_125_3477_n2382, DP_OP_423J2_125_3477_n2381,
         DP_OP_423J2_125_3477_n2380, DP_OP_423J2_125_3477_n2379,
         DP_OP_423J2_125_3477_n2378, DP_OP_423J2_125_3477_n2377,
         DP_OP_423J2_125_3477_n2376, DP_OP_423J2_125_3477_n2375,
         DP_OP_423J2_125_3477_n2374, DP_OP_423J2_125_3477_n2373,
         DP_OP_423J2_125_3477_n2372, DP_OP_423J2_125_3477_n2371,
         DP_OP_423J2_125_3477_n2370, DP_OP_423J2_125_3477_n2369,
         DP_OP_423J2_125_3477_n2368, DP_OP_423J2_125_3477_n2367,
         DP_OP_423J2_125_3477_n2366, DP_OP_423J2_125_3477_n2364,
         DP_OP_423J2_125_3477_n2363, DP_OP_423J2_125_3477_n2362,
         DP_OP_423J2_125_3477_n2361, DP_OP_423J2_125_3477_n2354,
         DP_OP_423J2_125_3477_n2353, DP_OP_423J2_125_3477_n2352,
         DP_OP_423J2_125_3477_n2351, DP_OP_423J2_125_3477_n2350,
         DP_OP_423J2_125_3477_n2349, DP_OP_423J2_125_3477_n2348,
         DP_OP_423J2_125_3477_n2347, DP_OP_423J2_125_3477_n2346,
         DP_OP_423J2_125_3477_n2345, DP_OP_423J2_125_3477_n2344,
         DP_OP_423J2_125_3477_n2343, DP_OP_423J2_125_3477_n2342,
         DP_OP_423J2_125_3477_n2341, DP_OP_423J2_125_3477_n2340,
         DP_OP_423J2_125_3477_n2339, DP_OP_423J2_125_3477_n2338,
         DP_OP_423J2_125_3477_n2337, DP_OP_423J2_125_3477_n2336,
         DP_OP_423J2_125_3477_n2335, DP_OP_423J2_125_3477_n2334,
         DP_OP_423J2_125_3477_n2333, DP_OP_423J2_125_3477_n2332,
         DP_OP_423J2_125_3477_n2331, DP_OP_423J2_125_3477_n2330,
         DP_OP_423J2_125_3477_n2329, DP_OP_423J2_125_3477_n2328,
         DP_OP_423J2_125_3477_n2327, DP_OP_423J2_125_3477_n2326,
         DP_OP_423J2_125_3477_n2325, DP_OP_423J2_125_3477_n2324,
         DP_OP_423J2_125_3477_n2323, DP_OP_423J2_125_3477_n2322,
         DP_OP_423J2_125_3477_n2321, DP_OP_423J2_125_3477_n2320,
         DP_OP_423J2_125_3477_n2318, DP_OP_423J2_125_3477_n2317,
         DP_OP_423J2_125_3477_n2316, DP_OP_423J2_125_3477_n2315,
         DP_OP_423J2_125_3477_n2311, DP_OP_423J2_125_3477_n2310,
         DP_OP_423J2_125_3477_n2309, DP_OP_423J2_125_3477_n2308,
         DP_OP_423J2_125_3477_n2307, DP_OP_423J2_125_3477_n2306,
         DP_OP_423J2_125_3477_n2305, DP_OP_423J2_125_3477_n2304,
         DP_OP_423J2_125_3477_n2303, DP_OP_423J2_125_3477_n2302,
         DP_OP_423J2_125_3477_n2301, DP_OP_423J2_125_3477_n2300,
         DP_OP_423J2_125_3477_n2299, DP_OP_423J2_125_3477_n2298,
         DP_OP_423J2_125_3477_n2297, DP_OP_423J2_125_3477_n2296,
         DP_OP_423J2_125_3477_n2295, DP_OP_423J2_125_3477_n2294,
         DP_OP_423J2_125_3477_n2293, DP_OP_423J2_125_3477_n2292,
         DP_OP_423J2_125_3477_n2291, DP_OP_423J2_125_3477_n2290,
         DP_OP_423J2_125_3477_n2289, DP_OP_423J2_125_3477_n2288,
         DP_OP_423J2_125_3477_n2287, DP_OP_423J2_125_3477_n2286,
         DP_OP_423J2_125_3477_n2285, DP_OP_423J2_125_3477_n2284,
         DP_OP_423J2_125_3477_n2283, DP_OP_423J2_125_3477_n2282,
         DP_OP_423J2_125_3477_n2281, DP_OP_423J2_125_3477_n2280,
         DP_OP_423J2_125_3477_n2279, DP_OP_423J2_125_3477_n2278,
         DP_OP_423J2_125_3477_n2277, DP_OP_423J2_125_3477_n2276,
         DP_OP_423J2_125_3477_n2273, DP_OP_423J2_125_3477_n2272,
         DP_OP_423J2_125_3477_n2271, DP_OP_423J2_125_3477_n2269,
         DP_OP_423J2_125_3477_n2268, DP_OP_423J2_125_3477_n2267,
         DP_OP_423J2_125_3477_n2265, DP_OP_423J2_125_3477_n2264,
         DP_OP_423J2_125_3477_n2263, DP_OP_423J2_125_3477_n2262,
         DP_OP_423J2_125_3477_n2261, DP_OP_423J2_125_3477_n2260,
         DP_OP_423J2_125_3477_n2259, DP_OP_423J2_125_3477_n2258,
         DP_OP_423J2_125_3477_n2257, DP_OP_423J2_125_3477_n2256,
         DP_OP_423J2_125_3477_n2255, DP_OP_423J2_125_3477_n2254,
         DP_OP_423J2_125_3477_n2253, DP_OP_423J2_125_3477_n2252,
         DP_OP_423J2_125_3477_n2251, DP_OP_423J2_125_3477_n2250,
         DP_OP_423J2_125_3477_n2249, DP_OP_423J2_125_3477_n2248,
         DP_OP_423J2_125_3477_n2247, DP_OP_423J2_125_3477_n2246,
         DP_OP_423J2_125_3477_n2245, DP_OP_423J2_125_3477_n2244,
         DP_OP_423J2_125_3477_n2243, DP_OP_423J2_125_3477_n2242,
         DP_OP_423J2_125_3477_n2241, DP_OP_423J2_125_3477_n2240,
         DP_OP_423J2_125_3477_n2239, DP_OP_423J2_125_3477_n2238,
         DP_OP_423J2_125_3477_n2237, DP_OP_423J2_125_3477_n2236,
         DP_OP_423J2_125_3477_n2235, DP_OP_423J2_125_3477_n2234,
         DP_OP_423J2_125_3477_n2233, DP_OP_423J2_125_3477_n2232,
         DP_OP_423J2_125_3477_n2230, DP_OP_423J2_125_3477_n2229,
         DP_OP_423J2_125_3477_n2228, DP_OP_423J2_125_3477_n2227,
         DP_OP_423J2_125_3477_n2225, DP_OP_423J2_125_3477_n2222,
         DP_OP_423J2_125_3477_n2221, DP_OP_423J2_125_3477_n2220,
         DP_OP_423J2_125_3477_n2219, DP_OP_423J2_125_3477_n2218,
         DP_OP_423J2_125_3477_n2217, DP_OP_423J2_125_3477_n2216,
         DP_OP_423J2_125_3477_n2215, DP_OP_423J2_125_3477_n2214,
         DP_OP_423J2_125_3477_n2213, DP_OP_423J2_125_3477_n2212,
         DP_OP_423J2_125_3477_n2211, DP_OP_423J2_125_3477_n2210,
         DP_OP_423J2_125_3477_n2209, DP_OP_423J2_125_3477_n2208,
         DP_OP_423J2_125_3477_n2207, DP_OP_423J2_125_3477_n2206,
         DP_OP_423J2_125_3477_n2205, DP_OP_423J2_125_3477_n2204,
         DP_OP_423J2_125_3477_n2203, DP_OP_423J2_125_3477_n2202,
         DP_OP_423J2_125_3477_n2201, DP_OP_423J2_125_3477_n2200,
         DP_OP_423J2_125_3477_n2199, DP_OP_423J2_125_3477_n2198,
         DP_OP_423J2_125_3477_n2197, DP_OP_423J2_125_3477_n2196,
         DP_OP_423J2_125_3477_n2195, DP_OP_423J2_125_3477_n2194,
         DP_OP_423J2_125_3477_n2193, DP_OP_423J2_125_3477_n2192,
         DP_OP_423J2_125_3477_n2191, DP_OP_423J2_125_3477_n2190,
         DP_OP_423J2_125_3477_n2185, DP_OP_423J2_125_3477_n2182,
         DP_OP_423J2_125_3477_n2178, DP_OP_423J2_125_3477_n2177,
         DP_OP_423J2_125_3477_n2176, DP_OP_423J2_125_3477_n2175,
         DP_OP_423J2_125_3477_n2174, DP_OP_423J2_125_3477_n2173,
         DP_OP_423J2_125_3477_n2172, DP_OP_423J2_125_3477_n2171,
         DP_OP_423J2_125_3477_n2170, DP_OP_423J2_125_3477_n2169,
         DP_OP_423J2_125_3477_n2168, DP_OP_423J2_125_3477_n2167,
         DP_OP_423J2_125_3477_n2166, DP_OP_423J2_125_3477_n2165,
         DP_OP_423J2_125_3477_n2164, DP_OP_423J2_125_3477_n2163,
         DP_OP_423J2_125_3477_n2162, DP_OP_423J2_125_3477_n2161,
         DP_OP_423J2_125_3477_n2160, DP_OP_423J2_125_3477_n2159,
         DP_OP_423J2_125_3477_n2158, DP_OP_423J2_125_3477_n2157,
         DP_OP_423J2_125_3477_n2156, DP_OP_423J2_125_3477_n2155,
         DP_OP_423J2_125_3477_n2154, DP_OP_423J2_125_3477_n2153,
         DP_OP_423J2_125_3477_n2152, DP_OP_423J2_125_3477_n2151,
         DP_OP_423J2_125_3477_n2150, DP_OP_423J2_125_3477_n2149,
         DP_OP_423J2_125_3477_n2148, DP_OP_423J2_125_3477_n2147,
         DP_OP_423J2_125_3477_n2146, DP_OP_423J2_125_3477_n2140,
         DP_OP_423J2_125_3477_n2135, DP_OP_423J2_125_3477_n2133,
         DP_OP_423J2_125_3477_n2132, DP_OP_423J2_125_3477_n2131,
         DP_OP_423J2_125_3477_n2130, DP_OP_423J2_125_3477_n2129,
         DP_OP_423J2_125_3477_n2128, DP_OP_423J2_125_3477_n2127,
         DP_OP_423J2_125_3477_n2126, DP_OP_423J2_125_3477_n2125,
         DP_OP_423J2_125_3477_n2124, DP_OP_423J2_125_3477_n2123,
         DP_OP_423J2_125_3477_n2122, DP_OP_423J2_125_3477_n2121,
         DP_OP_423J2_125_3477_n2120, DP_OP_423J2_125_3477_n2119,
         DP_OP_423J2_125_3477_n2118, DP_OP_423J2_125_3477_n2117,
         DP_OP_423J2_125_3477_n2116, DP_OP_423J2_125_3477_n2115,
         DP_OP_423J2_125_3477_n2114, DP_OP_423J2_125_3477_n2113,
         DP_OP_423J2_125_3477_n2112, DP_OP_423J2_125_3477_n2111,
         DP_OP_423J2_125_3477_n2110, DP_OP_423J2_125_3477_n2109,
         DP_OP_423J2_125_3477_n2108, DP_OP_423J2_125_3477_n2107,
         DP_OP_423J2_125_3477_n2106, DP_OP_423J2_125_3477_n2105,
         DP_OP_423J2_125_3477_n2104, DP_OP_423J2_125_3477_n2103,
         DP_OP_423J2_125_3477_n2102, DP_OP_423J2_125_3477_n2101,
         DP_OP_423J2_125_3477_n2100, DP_OP_423J2_125_3477_n2099,
         DP_OP_423J2_125_3477_n2098, DP_OP_423J2_125_3477_n2097,
         DP_OP_423J2_125_3477_n2096, DP_OP_423J2_125_3477_n2094,
         DP_OP_423J2_125_3477_n2090, DP_OP_423J2_125_3477_n2089,
         DP_OP_423J2_125_3477_n2088, DP_OP_423J2_125_3477_n2087,
         DP_OP_423J2_125_3477_n2086, DP_OP_423J2_125_3477_n2085,
         DP_OP_423J2_125_3477_n2084, DP_OP_423J2_125_3477_n2083,
         DP_OP_423J2_125_3477_n2082, DP_OP_423J2_125_3477_n2081,
         DP_OP_423J2_125_3477_n2080, DP_OP_423J2_125_3477_n2079,
         DP_OP_423J2_125_3477_n2078, DP_OP_423J2_125_3477_n2077,
         DP_OP_423J2_125_3477_n2076, DP_OP_423J2_125_3477_n2075,
         DP_OP_423J2_125_3477_n2074, DP_OP_423J2_125_3477_n2073,
         DP_OP_423J2_125_3477_n2072, DP_OP_423J2_125_3477_n2071,
         DP_OP_423J2_125_3477_n2070, DP_OP_423J2_125_3477_n2069,
         DP_OP_423J2_125_3477_n2068, DP_OP_423J2_125_3477_n2067,
         DP_OP_423J2_125_3477_n2066, DP_OP_423J2_125_3477_n2064,
         DP_OP_423J2_125_3477_n2063, DP_OP_423J2_125_3477_n2062,
         DP_OP_423J2_125_3477_n2061, DP_OP_423J2_125_3477_n2060,
         DP_OP_423J2_125_3477_n2059, DP_OP_423J2_125_3477_n2058,
         DP_OP_423J2_125_3477_n2053, DP_OP_423J2_125_3477_n2052,
         DP_OP_423J2_125_3477_n2051, DP_OP_423J2_125_3477_n2048,
         DP_OP_423J2_125_3477_n2045, DP_OP_423J2_125_3477_n2044,
         DP_OP_423J2_125_3477_n2043, DP_OP_423J2_125_3477_n2042,
         DP_OP_423J2_125_3477_n2041, DP_OP_423J2_125_3477_n2040,
         DP_OP_423J2_125_3477_n2039, DP_OP_423J2_125_3477_n2038,
         DP_OP_423J2_125_3477_n2037, DP_OP_423J2_125_3477_n2036,
         DP_OP_423J2_125_3477_n2035, DP_OP_423J2_125_3477_n2034,
         DP_OP_423J2_125_3477_n2033, DP_OP_423J2_125_3477_n2032,
         DP_OP_423J2_125_3477_n2031, DP_OP_423J2_125_3477_n2030,
         DP_OP_423J2_125_3477_n2029, DP_OP_423J2_125_3477_n2028,
         DP_OP_423J2_125_3477_n2027, DP_OP_423J2_125_3477_n2026,
         DP_OP_423J2_125_3477_n2025, DP_OP_423J2_125_3477_n2024,
         DP_OP_423J2_125_3477_n2023, DP_OP_423J2_125_3477_n2022,
         DP_OP_423J2_125_3477_n2021, DP_OP_423J2_125_3477_n2020,
         DP_OP_423J2_125_3477_n2019, DP_OP_423J2_125_3477_n2018,
         DP_OP_423J2_125_3477_n2017, DP_OP_423J2_125_3477_n2016,
         DP_OP_423J2_125_3477_n2015, DP_OP_423J2_125_3477_n2014,
         DP_OP_423J2_125_3477_n2013, DP_OP_423J2_125_3477_n2012,
         DP_OP_423J2_125_3477_n2010, DP_OP_423J2_125_3477_n2008,
         DP_OP_423J2_125_3477_n2007, DP_OP_423J2_125_3477_n2006,
         DP_OP_423J2_125_3477_n2005, DP_OP_423J2_125_3477_n2003,
         DP_OP_423J2_125_3477_n2001, DP_OP_423J2_125_3477_n1999,
         DP_OP_423J2_125_3477_n1998, DP_OP_423J2_125_3477_n1997,
         DP_OP_423J2_125_3477_n1996, DP_OP_423J2_125_3477_n1995,
         DP_OP_423J2_125_3477_n1994, DP_OP_423J2_125_3477_n1993,
         DP_OP_423J2_125_3477_n1992, DP_OP_423J2_125_3477_n1991,
         DP_OP_423J2_125_3477_n1990, DP_OP_423J2_125_3477_n1989,
         DP_OP_423J2_125_3477_n1988, DP_OP_423J2_125_3477_n1987,
         DP_OP_423J2_125_3477_n1986, DP_OP_423J2_125_3477_n1985,
         DP_OP_423J2_125_3477_n1984, DP_OP_423J2_125_3477_n1983,
         DP_OP_423J2_125_3477_n1982, DP_OP_423J2_125_3477_n1981,
         DP_OP_423J2_125_3477_n1980, DP_OP_423J2_125_3477_n1979,
         DP_OP_423J2_125_3477_n1978, DP_OP_423J2_125_3477_n1977,
         DP_OP_423J2_125_3477_n1976, DP_OP_423J2_125_3477_n1975,
         DP_OP_423J2_125_3477_n1974, DP_OP_423J2_125_3477_n1973,
         DP_OP_423J2_125_3477_n1972, DP_OP_423J2_125_3477_n1971,
         DP_OP_423J2_125_3477_n1970, DP_OP_423J2_125_3477_n1936,
         DP_OP_423J2_125_3477_n1934, DP_OP_423J2_125_3477_n1933,
         DP_OP_423J2_125_3477_n1932, DP_OP_423J2_125_3477_n1931,
         DP_OP_423J2_125_3477_n1930, DP_OP_423J2_125_3477_n1929,
         DP_OP_423J2_125_3477_n1928, DP_OP_423J2_125_3477_n1927,
         DP_OP_423J2_125_3477_n1926, DP_OP_423J2_125_3477_n1925,
         DP_OP_423J2_125_3477_n1924, DP_OP_423J2_125_3477_n1923,
         DP_OP_423J2_125_3477_n1921, DP_OP_423J2_125_3477_n1920,
         DP_OP_423J2_125_3477_n1919, DP_OP_423J2_125_3477_n1918,
         DP_OP_423J2_125_3477_n1917, DP_OP_423J2_125_3477_n1916,
         DP_OP_423J2_125_3477_n1915, DP_OP_423J2_125_3477_n1914,
         DP_OP_423J2_125_3477_n1913, DP_OP_423J2_125_3477_n1912,
         DP_OP_423J2_125_3477_n1911, DP_OP_423J2_125_3477_n1910,
         DP_OP_423J2_125_3477_n1909, DP_OP_423J2_125_3477_n1908,
         DP_OP_423J2_125_3477_n1907, DP_OP_423J2_125_3477_n1906,
         DP_OP_423J2_125_3477_n1905, DP_OP_423J2_125_3477_n1904,
         DP_OP_423J2_125_3477_n1903, DP_OP_423J2_125_3477_n1902,
         DP_OP_423J2_125_3477_n1901, DP_OP_423J2_125_3477_n1900,
         DP_OP_423J2_125_3477_n1899, DP_OP_423J2_125_3477_n1898,
         DP_OP_423J2_125_3477_n1897, DP_OP_423J2_125_3477_n1895,
         DP_OP_423J2_125_3477_n1894, DP_OP_423J2_125_3477_n1893,
         DP_OP_423J2_125_3477_n1892, DP_OP_423J2_125_3477_n1891,
         DP_OP_423J2_125_3477_n1890, DP_OP_423J2_125_3477_n1889,
         DP_OP_423J2_125_3477_n1888, DP_OP_423J2_125_3477_n1887,
         DP_OP_423J2_125_3477_n1886, DP_OP_423J2_125_3477_n1885,
         DP_OP_423J2_125_3477_n1884, DP_OP_423J2_125_3477_n1883,
         DP_OP_423J2_125_3477_n1882, DP_OP_423J2_125_3477_n1881,
         DP_OP_423J2_125_3477_n1880, DP_OP_423J2_125_3477_n1879,
         DP_OP_423J2_125_3477_n1878, DP_OP_423J2_125_3477_n1877,
         DP_OP_423J2_125_3477_n1876, DP_OP_423J2_125_3477_n1875,
         DP_OP_423J2_125_3477_n1874, DP_OP_423J2_125_3477_n1873,
         DP_OP_423J2_125_3477_n1872, DP_OP_423J2_125_3477_n1871,
         DP_OP_423J2_125_3477_n1870, DP_OP_423J2_125_3477_n1869,
         DP_OP_423J2_125_3477_n1868, DP_OP_423J2_125_3477_n1867,
         DP_OP_423J2_125_3477_n1866, DP_OP_423J2_125_3477_n1865,
         DP_OP_423J2_125_3477_n1864, DP_OP_423J2_125_3477_n1863,
         DP_OP_423J2_125_3477_n1862, DP_OP_423J2_125_3477_n1861,
         DP_OP_423J2_125_3477_n1860, DP_OP_423J2_125_3477_n1859,
         DP_OP_423J2_125_3477_n1858, DP_OP_423J2_125_3477_n1857,
         DP_OP_423J2_125_3477_n1856, DP_OP_423J2_125_3477_n1855,
         DP_OP_423J2_125_3477_n1854, DP_OP_423J2_125_3477_n1853,
         DP_OP_423J2_125_3477_n1852, DP_OP_423J2_125_3477_n1851,
         DP_OP_423J2_125_3477_n1850, DP_OP_423J2_125_3477_n1849,
         DP_OP_423J2_125_3477_n1848, DP_OP_423J2_125_3477_n1847,
         DP_OP_423J2_125_3477_n1846, DP_OP_423J2_125_3477_n1845,
         DP_OP_423J2_125_3477_n1844, DP_OP_423J2_125_3477_n1843,
         DP_OP_423J2_125_3477_n1842, DP_OP_423J2_125_3477_n1841,
         DP_OP_423J2_125_3477_n1840, DP_OP_423J2_125_3477_n1839,
         DP_OP_423J2_125_3477_n1838, DP_OP_423J2_125_3477_n1837,
         DP_OP_423J2_125_3477_n1836, DP_OP_423J2_125_3477_n1835,
         DP_OP_423J2_125_3477_n1834, DP_OP_423J2_125_3477_n1833,
         DP_OP_423J2_125_3477_n1832, DP_OP_423J2_125_3477_n1831,
         DP_OP_423J2_125_3477_n1830, DP_OP_423J2_125_3477_n1829,
         DP_OP_423J2_125_3477_n1828, DP_OP_423J2_125_3477_n1827,
         DP_OP_423J2_125_3477_n1826, DP_OP_423J2_125_3477_n1825,
         DP_OP_423J2_125_3477_n1824, DP_OP_423J2_125_3477_n1823,
         DP_OP_423J2_125_3477_n1822, DP_OP_423J2_125_3477_n1821,
         DP_OP_423J2_125_3477_n1820, DP_OP_423J2_125_3477_n1819,
         DP_OP_423J2_125_3477_n1818, DP_OP_423J2_125_3477_n1817,
         DP_OP_423J2_125_3477_n1816, DP_OP_423J2_125_3477_n1815,
         DP_OP_423J2_125_3477_n1814, DP_OP_423J2_125_3477_n1813,
         DP_OP_423J2_125_3477_n1812, DP_OP_423J2_125_3477_n1811,
         DP_OP_423J2_125_3477_n1810, DP_OP_423J2_125_3477_n1809,
         DP_OP_423J2_125_3477_n1808, DP_OP_423J2_125_3477_n1807,
         DP_OP_423J2_125_3477_n1806, DP_OP_423J2_125_3477_n1805,
         DP_OP_423J2_125_3477_n1804, DP_OP_423J2_125_3477_n1803,
         DP_OP_423J2_125_3477_n1802, DP_OP_423J2_125_3477_n1801,
         DP_OP_423J2_125_3477_n1800, DP_OP_423J2_125_3477_n1799,
         DP_OP_423J2_125_3477_n1798, DP_OP_423J2_125_3477_n1797,
         DP_OP_423J2_125_3477_n1796, DP_OP_423J2_125_3477_n1795,
         DP_OP_423J2_125_3477_n1794, DP_OP_423J2_125_3477_n1793,
         DP_OP_423J2_125_3477_n1792, DP_OP_423J2_125_3477_n1791,
         DP_OP_423J2_125_3477_n1790, DP_OP_423J2_125_3477_n1789,
         DP_OP_423J2_125_3477_n1788, DP_OP_423J2_125_3477_n1787,
         DP_OP_423J2_125_3477_n1786, DP_OP_423J2_125_3477_n1785,
         DP_OP_423J2_125_3477_n1784, DP_OP_423J2_125_3477_n1783,
         DP_OP_423J2_125_3477_n1782, DP_OP_423J2_125_3477_n1781,
         DP_OP_423J2_125_3477_n1780, DP_OP_423J2_125_3477_n1779,
         DP_OP_423J2_125_3477_n1778, DP_OP_423J2_125_3477_n1777,
         DP_OP_423J2_125_3477_n1776, DP_OP_423J2_125_3477_n1775,
         DP_OP_423J2_125_3477_n1774, DP_OP_423J2_125_3477_n1773,
         DP_OP_423J2_125_3477_n1772, DP_OP_423J2_125_3477_n1771,
         DP_OP_423J2_125_3477_n1770, DP_OP_423J2_125_3477_n1769,
         DP_OP_423J2_125_3477_n1768, DP_OP_423J2_125_3477_n1767,
         DP_OP_423J2_125_3477_n1766, DP_OP_423J2_125_3477_n1765,
         DP_OP_423J2_125_3477_n1764, DP_OP_423J2_125_3477_n1763,
         DP_OP_423J2_125_3477_n1762, DP_OP_423J2_125_3477_n1761,
         DP_OP_423J2_125_3477_n1760, DP_OP_423J2_125_3477_n1759,
         DP_OP_423J2_125_3477_n1758, DP_OP_423J2_125_3477_n1757,
         DP_OP_423J2_125_3477_n1756, DP_OP_423J2_125_3477_n1755,
         DP_OP_423J2_125_3477_n1754, DP_OP_423J2_125_3477_n1753,
         DP_OP_423J2_125_3477_n1752, DP_OP_423J2_125_3477_n1751,
         DP_OP_423J2_125_3477_n1750, DP_OP_423J2_125_3477_n1749,
         DP_OP_423J2_125_3477_n1748, DP_OP_423J2_125_3477_n1747,
         DP_OP_423J2_125_3477_n1746, DP_OP_423J2_125_3477_n1745,
         DP_OP_423J2_125_3477_n1744, DP_OP_423J2_125_3477_n1743,
         DP_OP_423J2_125_3477_n1742, DP_OP_423J2_125_3477_n1741,
         DP_OP_423J2_125_3477_n1740, DP_OP_423J2_125_3477_n1739,
         DP_OP_423J2_125_3477_n1738, DP_OP_423J2_125_3477_n1737,
         DP_OP_423J2_125_3477_n1736, DP_OP_423J2_125_3477_n1735,
         DP_OP_423J2_125_3477_n1734, DP_OP_423J2_125_3477_n1733,
         DP_OP_423J2_125_3477_n1732, DP_OP_423J2_125_3477_n1731,
         DP_OP_423J2_125_3477_n1730, DP_OP_423J2_125_3477_n1729,
         DP_OP_423J2_125_3477_n1728, DP_OP_423J2_125_3477_n1727,
         DP_OP_423J2_125_3477_n1726, DP_OP_423J2_125_3477_n1725,
         DP_OP_423J2_125_3477_n1724, DP_OP_423J2_125_3477_n1723,
         DP_OP_423J2_125_3477_n1722, DP_OP_423J2_125_3477_n1721,
         DP_OP_423J2_125_3477_n1720, DP_OP_423J2_125_3477_n1719,
         DP_OP_423J2_125_3477_n1718, DP_OP_423J2_125_3477_n1717,
         DP_OP_423J2_125_3477_n1716, DP_OP_423J2_125_3477_n1715,
         DP_OP_423J2_125_3477_n1714, DP_OP_423J2_125_3477_n1713,
         DP_OP_423J2_125_3477_n1712, DP_OP_423J2_125_3477_n1711,
         DP_OP_423J2_125_3477_n1710, DP_OP_423J2_125_3477_n1709,
         DP_OP_423J2_125_3477_n1708, DP_OP_423J2_125_3477_n1707,
         DP_OP_423J2_125_3477_n1706, DP_OP_423J2_125_3477_n1705,
         DP_OP_423J2_125_3477_n1704, DP_OP_423J2_125_3477_n1703,
         DP_OP_423J2_125_3477_n1702, DP_OP_423J2_125_3477_n1701,
         DP_OP_423J2_125_3477_n1700, DP_OP_423J2_125_3477_n1699,
         DP_OP_423J2_125_3477_n1698, DP_OP_423J2_125_3477_n1697,
         DP_OP_423J2_125_3477_n1696, DP_OP_423J2_125_3477_n1695,
         DP_OP_423J2_125_3477_n1694, DP_OP_423J2_125_3477_n1693,
         DP_OP_423J2_125_3477_n1692, DP_OP_423J2_125_3477_n1691,
         DP_OP_423J2_125_3477_n1690, DP_OP_423J2_125_3477_n1689,
         DP_OP_423J2_125_3477_n1688, DP_OP_423J2_125_3477_n1687,
         DP_OP_423J2_125_3477_n1686, DP_OP_423J2_125_3477_n1685,
         DP_OP_423J2_125_3477_n1684, DP_OP_423J2_125_3477_n1683,
         DP_OP_423J2_125_3477_n1682, DP_OP_423J2_125_3477_n1681,
         DP_OP_423J2_125_3477_n1680, DP_OP_423J2_125_3477_n1679,
         DP_OP_423J2_125_3477_n1678, DP_OP_423J2_125_3477_n1677,
         DP_OP_423J2_125_3477_n1676, DP_OP_423J2_125_3477_n1675,
         DP_OP_423J2_125_3477_n1674, DP_OP_423J2_125_3477_n1673,
         DP_OP_423J2_125_3477_n1672, DP_OP_423J2_125_3477_n1671,
         DP_OP_423J2_125_3477_n1670, DP_OP_423J2_125_3477_n1669,
         DP_OP_423J2_125_3477_n1668, DP_OP_423J2_125_3477_n1667,
         DP_OP_423J2_125_3477_n1666, DP_OP_423J2_125_3477_n1665,
         DP_OP_423J2_125_3477_n1664, DP_OP_423J2_125_3477_n1663,
         DP_OP_423J2_125_3477_n1662, DP_OP_423J2_125_3477_n1661,
         DP_OP_423J2_125_3477_n1660, DP_OP_423J2_125_3477_n1659,
         DP_OP_423J2_125_3477_n1658, DP_OP_423J2_125_3477_n1657,
         DP_OP_423J2_125_3477_n1656, DP_OP_423J2_125_3477_n1655,
         DP_OP_423J2_125_3477_n1654, DP_OP_423J2_125_3477_n1653,
         DP_OP_423J2_125_3477_n1652, DP_OP_423J2_125_3477_n1651,
         DP_OP_423J2_125_3477_n1650, DP_OP_423J2_125_3477_n1649,
         DP_OP_423J2_125_3477_n1648, DP_OP_423J2_125_3477_n1647,
         DP_OP_423J2_125_3477_n1646, DP_OP_423J2_125_3477_n1645,
         DP_OP_423J2_125_3477_n1644, DP_OP_423J2_125_3477_n1643,
         DP_OP_423J2_125_3477_n1642, DP_OP_423J2_125_3477_n1641,
         DP_OP_423J2_125_3477_n1640, DP_OP_423J2_125_3477_n1639,
         DP_OP_423J2_125_3477_n1638, DP_OP_423J2_125_3477_n1637,
         DP_OP_423J2_125_3477_n1636, DP_OP_423J2_125_3477_n1635,
         DP_OP_423J2_125_3477_n1634, DP_OP_423J2_125_3477_n1633,
         DP_OP_423J2_125_3477_n1632, DP_OP_423J2_125_3477_n1631,
         DP_OP_423J2_125_3477_n1630, DP_OP_423J2_125_3477_n1629,
         DP_OP_423J2_125_3477_n1628, DP_OP_423J2_125_3477_n1627,
         DP_OP_423J2_125_3477_n1626, DP_OP_423J2_125_3477_n1625,
         DP_OP_423J2_125_3477_n1624, DP_OP_423J2_125_3477_n1623,
         DP_OP_423J2_125_3477_n1622, DP_OP_423J2_125_3477_n1621,
         DP_OP_423J2_125_3477_n1620, DP_OP_423J2_125_3477_n1619,
         DP_OP_423J2_125_3477_n1618, DP_OP_423J2_125_3477_n1617,
         DP_OP_423J2_125_3477_n1616, DP_OP_423J2_125_3477_n1615,
         DP_OP_423J2_125_3477_n1614, DP_OP_423J2_125_3477_n1613,
         DP_OP_423J2_125_3477_n1612, DP_OP_423J2_125_3477_n1611,
         DP_OP_423J2_125_3477_n1610, DP_OP_423J2_125_3477_n1609,
         DP_OP_423J2_125_3477_n1608, DP_OP_423J2_125_3477_n1607,
         DP_OP_423J2_125_3477_n1606, DP_OP_423J2_125_3477_n1605,
         DP_OP_423J2_125_3477_n1604, DP_OP_423J2_125_3477_n1603,
         DP_OP_423J2_125_3477_n1602, DP_OP_423J2_125_3477_n1601,
         DP_OP_423J2_125_3477_n1600, DP_OP_423J2_125_3477_n1599,
         DP_OP_423J2_125_3477_n1598, DP_OP_423J2_125_3477_n1597,
         DP_OP_423J2_125_3477_n1596, DP_OP_423J2_125_3477_n1595,
         DP_OP_423J2_125_3477_n1594, DP_OP_423J2_125_3477_n1593,
         DP_OP_423J2_125_3477_n1592, DP_OP_423J2_125_3477_n1591,
         DP_OP_423J2_125_3477_n1590, DP_OP_423J2_125_3477_n1589,
         DP_OP_423J2_125_3477_n1588, DP_OP_423J2_125_3477_n1587,
         DP_OP_423J2_125_3477_n1586, DP_OP_423J2_125_3477_n1585,
         DP_OP_423J2_125_3477_n1584, DP_OP_423J2_125_3477_n1583,
         DP_OP_423J2_125_3477_n1582, DP_OP_423J2_125_3477_n1581,
         DP_OP_423J2_125_3477_n1580, DP_OP_423J2_125_3477_n1579,
         DP_OP_423J2_125_3477_n1578, DP_OP_423J2_125_3477_n1577,
         DP_OP_423J2_125_3477_n1576, DP_OP_423J2_125_3477_n1575,
         DP_OP_423J2_125_3477_n1574, DP_OP_423J2_125_3477_n1573,
         DP_OP_423J2_125_3477_n1572, DP_OP_423J2_125_3477_n1571,
         DP_OP_423J2_125_3477_n1570, DP_OP_423J2_125_3477_n1569,
         DP_OP_423J2_125_3477_n1568, DP_OP_423J2_125_3477_n1567,
         DP_OP_423J2_125_3477_n1566, DP_OP_423J2_125_3477_n1565,
         DP_OP_423J2_125_3477_n1564, DP_OP_423J2_125_3477_n1563,
         DP_OP_423J2_125_3477_n1562, DP_OP_423J2_125_3477_n1561,
         DP_OP_423J2_125_3477_n1560, DP_OP_423J2_125_3477_n1559,
         DP_OP_423J2_125_3477_n1558, DP_OP_423J2_125_3477_n1557,
         DP_OP_423J2_125_3477_n1556, DP_OP_423J2_125_3477_n1555,
         DP_OP_423J2_125_3477_n1554, DP_OP_423J2_125_3477_n1553,
         DP_OP_423J2_125_3477_n1552, DP_OP_423J2_125_3477_n1551,
         DP_OP_423J2_125_3477_n1550, DP_OP_423J2_125_3477_n1549,
         DP_OP_423J2_125_3477_n1548, DP_OP_423J2_125_3477_n1547,
         DP_OP_423J2_125_3477_n1546, DP_OP_423J2_125_3477_n1545,
         DP_OP_423J2_125_3477_n1544, DP_OP_423J2_125_3477_n1543,
         DP_OP_423J2_125_3477_n1542, DP_OP_423J2_125_3477_n1541,
         DP_OP_423J2_125_3477_n1540, DP_OP_423J2_125_3477_n1539,
         DP_OP_423J2_125_3477_n1538, DP_OP_423J2_125_3477_n1537,
         DP_OP_423J2_125_3477_n1536, DP_OP_423J2_125_3477_n1535,
         DP_OP_423J2_125_3477_n1534, DP_OP_423J2_125_3477_n1533,
         DP_OP_423J2_125_3477_n1532, DP_OP_423J2_125_3477_n1531,
         DP_OP_423J2_125_3477_n1530, DP_OP_423J2_125_3477_n1529,
         DP_OP_423J2_125_3477_n1528, DP_OP_423J2_125_3477_n1527,
         DP_OP_423J2_125_3477_n1526, DP_OP_423J2_125_3477_n1525,
         DP_OP_423J2_125_3477_n1524, DP_OP_423J2_125_3477_n1523,
         DP_OP_423J2_125_3477_n1522, DP_OP_423J2_125_3477_n1521,
         DP_OP_423J2_125_3477_n1520, DP_OP_423J2_125_3477_n1519,
         DP_OP_423J2_125_3477_n1518, DP_OP_423J2_125_3477_n1517,
         DP_OP_423J2_125_3477_n1516, DP_OP_423J2_125_3477_n1515,
         DP_OP_423J2_125_3477_n1514, DP_OP_423J2_125_3477_n1513,
         DP_OP_423J2_125_3477_n1512, DP_OP_423J2_125_3477_n1511,
         DP_OP_423J2_125_3477_n1510, DP_OP_423J2_125_3477_n1509,
         DP_OP_423J2_125_3477_n1508, DP_OP_423J2_125_3477_n1507,
         DP_OP_423J2_125_3477_n1506, DP_OP_423J2_125_3477_n1505,
         DP_OP_423J2_125_3477_n1504, DP_OP_423J2_125_3477_n1503,
         DP_OP_423J2_125_3477_n1502, DP_OP_423J2_125_3477_n1501,
         DP_OP_423J2_125_3477_n1500, DP_OP_423J2_125_3477_n1499,
         DP_OP_423J2_125_3477_n1498, DP_OP_423J2_125_3477_n1497,
         DP_OP_423J2_125_3477_n1496, DP_OP_423J2_125_3477_n1495,
         DP_OP_423J2_125_3477_n1494, DP_OP_423J2_125_3477_n1493,
         DP_OP_423J2_125_3477_n1492, DP_OP_423J2_125_3477_n1491,
         DP_OP_423J2_125_3477_n1490, DP_OP_423J2_125_3477_n1489,
         DP_OP_423J2_125_3477_n1488, DP_OP_423J2_125_3477_n1487,
         DP_OP_423J2_125_3477_n1486, DP_OP_423J2_125_3477_n1485,
         DP_OP_423J2_125_3477_n1484, DP_OP_423J2_125_3477_n1483,
         DP_OP_423J2_125_3477_n1482, DP_OP_423J2_125_3477_n1481,
         DP_OP_423J2_125_3477_n1480, DP_OP_423J2_125_3477_n1479,
         DP_OP_423J2_125_3477_n1478, DP_OP_423J2_125_3477_n1477,
         DP_OP_423J2_125_3477_n1476, DP_OP_423J2_125_3477_n1475,
         DP_OP_423J2_125_3477_n1474, DP_OP_423J2_125_3477_n1473,
         DP_OP_423J2_125_3477_n1472, DP_OP_423J2_125_3477_n1471,
         DP_OP_423J2_125_3477_n1470, DP_OP_423J2_125_3477_n1469,
         DP_OP_423J2_125_3477_n1468, DP_OP_423J2_125_3477_n1467,
         DP_OP_423J2_125_3477_n1466, DP_OP_423J2_125_3477_n1465,
         DP_OP_423J2_125_3477_n1464, DP_OP_423J2_125_3477_n1463,
         DP_OP_423J2_125_3477_n1462, DP_OP_423J2_125_3477_n1461,
         DP_OP_423J2_125_3477_n1460, DP_OP_423J2_125_3477_n1459,
         DP_OP_423J2_125_3477_n1458, DP_OP_423J2_125_3477_n1457,
         DP_OP_423J2_125_3477_n1456, DP_OP_423J2_125_3477_n1455,
         DP_OP_423J2_125_3477_n1454, DP_OP_423J2_125_3477_n1453,
         DP_OP_423J2_125_3477_n1452, DP_OP_423J2_125_3477_n1451,
         DP_OP_423J2_125_3477_n1450, DP_OP_423J2_125_3477_n1449,
         DP_OP_423J2_125_3477_n1448, DP_OP_423J2_125_3477_n1447,
         DP_OP_423J2_125_3477_n1446, DP_OP_423J2_125_3477_n1445,
         DP_OP_423J2_125_3477_n1444, DP_OP_423J2_125_3477_n1443,
         DP_OP_423J2_125_3477_n1442, DP_OP_423J2_125_3477_n1441,
         DP_OP_423J2_125_3477_n1440, DP_OP_423J2_125_3477_n1439,
         DP_OP_423J2_125_3477_n1438, DP_OP_423J2_125_3477_n1437,
         DP_OP_423J2_125_3477_n1436, DP_OP_423J2_125_3477_n1435,
         DP_OP_423J2_125_3477_n1434, DP_OP_423J2_125_3477_n1433,
         DP_OP_423J2_125_3477_n1432, DP_OP_423J2_125_3477_n1431,
         DP_OP_423J2_125_3477_n1430, DP_OP_423J2_125_3477_n1429,
         DP_OP_423J2_125_3477_n1428, DP_OP_423J2_125_3477_n1427,
         DP_OP_423J2_125_3477_n1426, DP_OP_423J2_125_3477_n1425,
         DP_OP_423J2_125_3477_n1424, DP_OP_423J2_125_3477_n1423,
         DP_OP_423J2_125_3477_n1422, DP_OP_423J2_125_3477_n1421,
         DP_OP_423J2_125_3477_n1420, DP_OP_423J2_125_3477_n1419,
         DP_OP_423J2_125_3477_n1418, DP_OP_423J2_125_3477_n1417,
         DP_OP_423J2_125_3477_n1416, DP_OP_423J2_125_3477_n1415,
         DP_OP_423J2_125_3477_n1414, DP_OP_423J2_125_3477_n1413,
         DP_OP_423J2_125_3477_n1412, DP_OP_423J2_125_3477_n1411,
         DP_OP_423J2_125_3477_n1410, DP_OP_423J2_125_3477_n1409,
         DP_OP_423J2_125_3477_n1408, DP_OP_423J2_125_3477_n1407,
         DP_OP_423J2_125_3477_n1406, DP_OP_423J2_125_3477_n1405,
         DP_OP_423J2_125_3477_n1404, DP_OP_423J2_125_3477_n1403,
         DP_OP_423J2_125_3477_n1402, DP_OP_423J2_125_3477_n1401,
         DP_OP_423J2_125_3477_n1400, DP_OP_423J2_125_3477_n1399,
         DP_OP_423J2_125_3477_n1398, DP_OP_423J2_125_3477_n1397,
         DP_OP_423J2_125_3477_n1396, DP_OP_423J2_125_3477_n1395,
         DP_OP_423J2_125_3477_n1394, DP_OP_423J2_125_3477_n1393,
         DP_OP_423J2_125_3477_n1392, DP_OP_423J2_125_3477_n1391,
         DP_OP_423J2_125_3477_n1390, DP_OP_423J2_125_3477_n1389,
         DP_OP_423J2_125_3477_n1388, DP_OP_423J2_125_3477_n1387,
         DP_OP_423J2_125_3477_n1386, DP_OP_423J2_125_3477_n1385,
         DP_OP_423J2_125_3477_n1384, DP_OP_423J2_125_3477_n1383,
         DP_OP_423J2_125_3477_n1382, DP_OP_423J2_125_3477_n1381,
         DP_OP_423J2_125_3477_n1380, DP_OP_423J2_125_3477_n1379,
         DP_OP_423J2_125_3477_n1378, DP_OP_423J2_125_3477_n1377,
         DP_OP_423J2_125_3477_n1376, DP_OP_423J2_125_3477_n1375,
         DP_OP_423J2_125_3477_n1374, DP_OP_423J2_125_3477_n1373,
         DP_OP_423J2_125_3477_n1372, DP_OP_423J2_125_3477_n1371,
         DP_OP_423J2_125_3477_n1370, DP_OP_423J2_125_3477_n1369,
         DP_OP_423J2_125_3477_n1368, DP_OP_423J2_125_3477_n1367,
         DP_OP_423J2_125_3477_n1366, DP_OP_423J2_125_3477_n1365,
         DP_OP_423J2_125_3477_n1364, DP_OP_423J2_125_3477_n1363,
         DP_OP_423J2_125_3477_n1362, DP_OP_423J2_125_3477_n1361,
         DP_OP_423J2_125_3477_n1360, DP_OP_423J2_125_3477_n1359,
         DP_OP_423J2_125_3477_n1358, DP_OP_423J2_125_3477_n1357,
         DP_OP_423J2_125_3477_n1356, DP_OP_423J2_125_3477_n1355,
         DP_OP_423J2_125_3477_n1354, DP_OP_423J2_125_3477_n1353,
         DP_OP_423J2_125_3477_n1352, DP_OP_423J2_125_3477_n1351,
         DP_OP_423J2_125_3477_n1350, DP_OP_423J2_125_3477_n1349,
         DP_OP_423J2_125_3477_n1348, DP_OP_423J2_125_3477_n1347,
         DP_OP_423J2_125_3477_n1346, DP_OP_423J2_125_3477_n1345,
         DP_OP_423J2_125_3477_n1344, DP_OP_423J2_125_3477_n1343,
         DP_OP_423J2_125_3477_n1342, DP_OP_423J2_125_3477_n1341,
         DP_OP_423J2_125_3477_n1340, DP_OP_423J2_125_3477_n1339,
         DP_OP_423J2_125_3477_n1338, DP_OP_423J2_125_3477_n1337,
         DP_OP_423J2_125_3477_n1336, DP_OP_423J2_125_3477_n1335,
         DP_OP_423J2_125_3477_n1334, DP_OP_423J2_125_3477_n1333,
         DP_OP_423J2_125_3477_n1332, DP_OP_423J2_125_3477_n1331,
         DP_OP_423J2_125_3477_n1330, DP_OP_423J2_125_3477_n1329,
         DP_OP_423J2_125_3477_n1328, DP_OP_423J2_125_3477_n1327,
         DP_OP_423J2_125_3477_n1326, DP_OP_423J2_125_3477_n1325,
         DP_OP_423J2_125_3477_n1324, DP_OP_423J2_125_3477_n1323,
         DP_OP_423J2_125_3477_n1322, DP_OP_423J2_125_3477_n1321,
         DP_OP_423J2_125_3477_n1320, DP_OP_423J2_125_3477_n1319,
         DP_OP_423J2_125_3477_n1318, DP_OP_423J2_125_3477_n1317,
         DP_OP_423J2_125_3477_n1316, DP_OP_423J2_125_3477_n1315,
         DP_OP_423J2_125_3477_n1314, DP_OP_423J2_125_3477_n1313,
         DP_OP_423J2_125_3477_n1312, DP_OP_423J2_125_3477_n1311,
         DP_OP_423J2_125_3477_n1310, DP_OP_423J2_125_3477_n1309,
         DP_OP_423J2_125_3477_n1308, DP_OP_423J2_125_3477_n1307,
         DP_OP_423J2_125_3477_n1306, DP_OP_423J2_125_3477_n1305,
         DP_OP_423J2_125_3477_n1304, DP_OP_423J2_125_3477_n1303,
         DP_OP_423J2_125_3477_n1302, DP_OP_423J2_125_3477_n1301,
         DP_OP_423J2_125_3477_n1300, DP_OP_423J2_125_3477_n1299,
         DP_OP_423J2_125_3477_n1298, DP_OP_423J2_125_3477_n1297,
         DP_OP_423J2_125_3477_n1296, DP_OP_423J2_125_3477_n1295,
         DP_OP_423J2_125_3477_n1294, DP_OP_423J2_125_3477_n1293,
         DP_OP_423J2_125_3477_n1292, DP_OP_423J2_125_3477_n1291,
         DP_OP_423J2_125_3477_n1290, DP_OP_423J2_125_3477_n1289,
         DP_OP_423J2_125_3477_n1288, DP_OP_423J2_125_3477_n1287,
         DP_OP_423J2_125_3477_n1286, DP_OP_423J2_125_3477_n1285,
         DP_OP_423J2_125_3477_n1284, DP_OP_423J2_125_3477_n1283,
         DP_OP_423J2_125_3477_n1282, DP_OP_423J2_125_3477_n1281,
         DP_OP_423J2_125_3477_n1280, DP_OP_423J2_125_3477_n1279,
         DP_OP_423J2_125_3477_n1278, DP_OP_423J2_125_3477_n1277,
         DP_OP_423J2_125_3477_n1276, DP_OP_423J2_125_3477_n1275,
         DP_OP_423J2_125_3477_n1274, DP_OP_423J2_125_3477_n1273,
         DP_OP_423J2_125_3477_n1272, DP_OP_423J2_125_3477_n1271,
         DP_OP_423J2_125_3477_n1270, DP_OP_423J2_125_3477_n1269,
         DP_OP_423J2_125_3477_n1268, DP_OP_423J2_125_3477_n1267,
         DP_OP_423J2_125_3477_n1266, DP_OP_423J2_125_3477_n1265,
         DP_OP_423J2_125_3477_n1264, DP_OP_423J2_125_3477_n1263,
         DP_OP_423J2_125_3477_n1262, DP_OP_423J2_125_3477_n1261,
         DP_OP_423J2_125_3477_n1260, DP_OP_423J2_125_3477_n1259,
         DP_OP_423J2_125_3477_n1258, DP_OP_423J2_125_3477_n1257,
         DP_OP_423J2_125_3477_n1256, DP_OP_423J2_125_3477_n1255,
         DP_OP_423J2_125_3477_n1254, DP_OP_423J2_125_3477_n1253,
         DP_OP_423J2_125_3477_n1252, DP_OP_423J2_125_3477_n1251,
         DP_OP_423J2_125_3477_n1250, DP_OP_423J2_125_3477_n1249,
         DP_OP_423J2_125_3477_n1248, DP_OP_423J2_125_3477_n1247,
         DP_OP_423J2_125_3477_n1246, DP_OP_423J2_125_3477_n1245,
         DP_OP_423J2_125_3477_n1244, DP_OP_423J2_125_3477_n1243,
         DP_OP_423J2_125_3477_n1242, DP_OP_423J2_125_3477_n1241,
         DP_OP_423J2_125_3477_n1240, DP_OP_423J2_125_3477_n1239,
         DP_OP_423J2_125_3477_n1238, DP_OP_423J2_125_3477_n1237,
         DP_OP_423J2_125_3477_n1236, DP_OP_423J2_125_3477_n1235,
         DP_OP_423J2_125_3477_n1234, DP_OP_423J2_125_3477_n1233,
         DP_OP_423J2_125_3477_n1232, DP_OP_423J2_125_3477_n1231,
         DP_OP_423J2_125_3477_n1230, DP_OP_423J2_125_3477_n1229,
         DP_OP_423J2_125_3477_n1228, DP_OP_423J2_125_3477_n1227,
         DP_OP_423J2_125_3477_n1226, DP_OP_423J2_125_3477_n1225,
         DP_OP_423J2_125_3477_n1224, DP_OP_423J2_125_3477_n1223,
         DP_OP_423J2_125_3477_n1222, DP_OP_423J2_125_3477_n1221,
         DP_OP_423J2_125_3477_n1220, DP_OP_423J2_125_3477_n1219,
         DP_OP_423J2_125_3477_n1218, DP_OP_423J2_125_3477_n1217,
         DP_OP_423J2_125_3477_n1216, DP_OP_423J2_125_3477_n1215,
         DP_OP_423J2_125_3477_n1214, DP_OP_423J2_125_3477_n1213,
         DP_OP_423J2_125_3477_n1212, DP_OP_423J2_125_3477_n1211,
         DP_OP_423J2_125_3477_n1210, DP_OP_423J2_125_3477_n1209,
         DP_OP_423J2_125_3477_n1208, DP_OP_423J2_125_3477_n1207,
         DP_OP_423J2_125_3477_n1206, DP_OP_423J2_125_3477_n1205,
         DP_OP_423J2_125_3477_n1204, DP_OP_423J2_125_3477_n1203,
         DP_OP_423J2_125_3477_n1202, DP_OP_423J2_125_3477_n1201,
         DP_OP_423J2_125_3477_n1200, DP_OP_423J2_125_3477_n1199,
         DP_OP_423J2_125_3477_n1198, DP_OP_423J2_125_3477_n1197,
         DP_OP_423J2_125_3477_n1196, DP_OP_423J2_125_3477_n1195,
         DP_OP_423J2_125_3477_n1194, DP_OP_423J2_125_3477_n1193,
         DP_OP_423J2_125_3477_n1192, DP_OP_423J2_125_3477_n1191,
         DP_OP_423J2_125_3477_n1190, DP_OP_423J2_125_3477_n1189,
         DP_OP_423J2_125_3477_n1188, DP_OP_423J2_125_3477_n1187,
         DP_OP_423J2_125_3477_n1186, DP_OP_423J2_125_3477_n1185,
         DP_OP_423J2_125_3477_n1184, DP_OP_423J2_125_3477_n1183,
         DP_OP_423J2_125_3477_n1182, DP_OP_423J2_125_3477_n1181,
         DP_OP_423J2_125_3477_n1180, DP_OP_423J2_125_3477_n1179,
         DP_OP_423J2_125_3477_n1178, DP_OP_423J2_125_3477_n1177,
         DP_OP_423J2_125_3477_n1176, DP_OP_423J2_125_3477_n1175,
         DP_OP_423J2_125_3477_n1174, DP_OP_423J2_125_3477_n1173,
         DP_OP_423J2_125_3477_n1172, DP_OP_423J2_125_3477_n1171,
         DP_OP_423J2_125_3477_n1170, DP_OP_423J2_125_3477_n1169,
         DP_OP_423J2_125_3477_n1168, DP_OP_423J2_125_3477_n1167,
         DP_OP_423J2_125_3477_n1166, DP_OP_423J2_125_3477_n1165,
         DP_OP_423J2_125_3477_n1164, DP_OP_423J2_125_3477_n1163,
         DP_OP_423J2_125_3477_n1162, DP_OP_423J2_125_3477_n1161,
         DP_OP_423J2_125_3477_n1160, DP_OP_423J2_125_3477_n1159,
         DP_OP_423J2_125_3477_n1158, DP_OP_423J2_125_3477_n1157,
         DP_OP_423J2_125_3477_n1156, DP_OP_423J2_125_3477_n1155,
         DP_OP_423J2_125_3477_n1154, DP_OP_423J2_125_3477_n1153,
         DP_OP_423J2_125_3477_n1152, DP_OP_423J2_125_3477_n1151,
         DP_OP_423J2_125_3477_n1150, DP_OP_423J2_125_3477_n1149,
         DP_OP_423J2_125_3477_n1148, DP_OP_423J2_125_3477_n1147,
         DP_OP_423J2_125_3477_n1146, DP_OP_423J2_125_3477_n1145,
         DP_OP_423J2_125_3477_n1144, DP_OP_423J2_125_3477_n1143,
         DP_OP_423J2_125_3477_n1142, DP_OP_423J2_125_3477_n1141,
         DP_OP_423J2_125_3477_n1140, DP_OP_423J2_125_3477_n1139,
         DP_OP_423J2_125_3477_n1138, DP_OP_423J2_125_3477_n1137,
         DP_OP_423J2_125_3477_n1136, DP_OP_423J2_125_3477_n1135,
         DP_OP_423J2_125_3477_n1134, DP_OP_423J2_125_3477_n1133,
         DP_OP_423J2_125_3477_n1132, DP_OP_423J2_125_3477_n1131,
         DP_OP_423J2_125_3477_n1130, DP_OP_423J2_125_3477_n1129,
         DP_OP_423J2_125_3477_n1128, DP_OP_423J2_125_3477_n1127,
         DP_OP_423J2_125_3477_n1126, DP_OP_423J2_125_3477_n1125,
         DP_OP_423J2_125_3477_n1124, DP_OP_423J2_125_3477_n1123,
         DP_OP_423J2_125_3477_n1122, DP_OP_423J2_125_3477_n1121,
         DP_OP_423J2_125_3477_n1120, DP_OP_423J2_125_3477_n1119,
         DP_OP_423J2_125_3477_n1118, DP_OP_423J2_125_3477_n1117,
         DP_OP_423J2_125_3477_n1116, DP_OP_423J2_125_3477_n1115,
         DP_OP_423J2_125_3477_n1114, DP_OP_423J2_125_3477_n1113,
         DP_OP_423J2_125_3477_n1112, DP_OP_423J2_125_3477_n1111,
         DP_OP_423J2_125_3477_n1110, DP_OP_423J2_125_3477_n1109,
         DP_OP_423J2_125_3477_n1108, DP_OP_423J2_125_3477_n1107,
         DP_OP_423J2_125_3477_n1106, DP_OP_423J2_125_3477_n1105,
         DP_OP_423J2_125_3477_n1104, DP_OP_423J2_125_3477_n1103,
         DP_OP_423J2_125_3477_n1102, DP_OP_423J2_125_3477_n1101,
         DP_OP_423J2_125_3477_n1100, DP_OP_423J2_125_3477_n1099,
         DP_OP_423J2_125_3477_n1098, DP_OP_423J2_125_3477_n1097,
         DP_OP_423J2_125_3477_n1096, DP_OP_423J2_125_3477_n1095,
         DP_OP_423J2_125_3477_n1094, DP_OP_423J2_125_3477_n1093,
         DP_OP_423J2_125_3477_n1092, DP_OP_423J2_125_3477_n1091,
         DP_OP_423J2_125_3477_n1090, DP_OP_423J2_125_3477_n1089,
         DP_OP_423J2_125_3477_n1088, DP_OP_423J2_125_3477_n1087,
         DP_OP_423J2_125_3477_n1086, DP_OP_423J2_125_3477_n1085,
         DP_OP_423J2_125_3477_n1084, DP_OP_423J2_125_3477_n1083,
         DP_OP_423J2_125_3477_n1082, DP_OP_423J2_125_3477_n1081,
         DP_OP_423J2_125_3477_n1080, DP_OP_423J2_125_3477_n1079,
         DP_OP_423J2_125_3477_n1078, DP_OP_423J2_125_3477_n1077,
         DP_OP_423J2_125_3477_n1076, DP_OP_423J2_125_3477_n1075,
         DP_OP_423J2_125_3477_n1074, DP_OP_423J2_125_3477_n1073,
         DP_OP_423J2_125_3477_n1072, DP_OP_423J2_125_3477_n1071,
         DP_OP_423J2_125_3477_n1070, DP_OP_423J2_125_3477_n1069,
         DP_OP_423J2_125_3477_n1068, DP_OP_423J2_125_3477_n1067,
         DP_OP_423J2_125_3477_n1066, DP_OP_423J2_125_3477_n1065,
         DP_OP_423J2_125_3477_n1064, DP_OP_423J2_125_3477_n1063,
         DP_OP_423J2_125_3477_n1062, DP_OP_423J2_125_3477_n1061,
         DP_OP_423J2_125_3477_n1060, DP_OP_423J2_125_3477_n1059,
         DP_OP_423J2_125_3477_n1058, DP_OP_423J2_125_3477_n1057,
         DP_OP_423J2_125_3477_n1056, DP_OP_423J2_125_3477_n1055,
         DP_OP_423J2_125_3477_n1054, DP_OP_423J2_125_3477_n1053,
         DP_OP_423J2_125_3477_n1052, DP_OP_423J2_125_3477_n1051,
         DP_OP_423J2_125_3477_n1050, DP_OP_423J2_125_3477_n1049,
         DP_OP_423J2_125_3477_n1048, DP_OP_423J2_125_3477_n1047,
         DP_OP_423J2_125_3477_n1046, DP_OP_423J2_125_3477_n1045,
         DP_OP_423J2_125_3477_n1044, DP_OP_423J2_125_3477_n1043,
         DP_OP_423J2_125_3477_n1042, DP_OP_423J2_125_3477_n1041,
         DP_OP_423J2_125_3477_n1040, DP_OP_423J2_125_3477_n1039,
         DP_OP_423J2_125_3477_n1038, DP_OP_423J2_125_3477_n1037,
         DP_OP_423J2_125_3477_n1036, DP_OP_423J2_125_3477_n1035,
         DP_OP_423J2_125_3477_n1034, DP_OP_423J2_125_3477_n1033,
         DP_OP_423J2_125_3477_n1032, DP_OP_423J2_125_3477_n1031,
         DP_OP_423J2_125_3477_n1030, DP_OP_423J2_125_3477_n1029,
         DP_OP_423J2_125_3477_n1028, DP_OP_423J2_125_3477_n1027,
         DP_OP_423J2_125_3477_n1026, DP_OP_423J2_125_3477_n1025,
         DP_OP_423J2_125_3477_n1024, DP_OP_423J2_125_3477_n1023,
         DP_OP_423J2_125_3477_n1022, DP_OP_423J2_125_3477_n1021,
         DP_OP_423J2_125_3477_n1020, DP_OP_423J2_125_3477_n1019,
         DP_OP_423J2_125_3477_n1018, DP_OP_423J2_125_3477_n1017,
         DP_OP_423J2_125_3477_n1016, DP_OP_423J2_125_3477_n1015,
         DP_OP_423J2_125_3477_n1014, DP_OP_423J2_125_3477_n1013,
         DP_OP_423J2_125_3477_n1012, DP_OP_423J2_125_3477_n1011,
         DP_OP_423J2_125_3477_n1010, DP_OP_423J2_125_3477_n1009,
         DP_OP_423J2_125_3477_n1008, DP_OP_423J2_125_3477_n1007,
         DP_OP_423J2_125_3477_n1006, DP_OP_423J2_125_3477_n1005,
         DP_OP_423J2_125_3477_n1004, DP_OP_423J2_125_3477_n1003,
         DP_OP_423J2_125_3477_n1002, DP_OP_423J2_125_3477_n1001,
         DP_OP_423J2_125_3477_n1000, DP_OP_423J2_125_3477_n999,
         DP_OP_423J2_125_3477_n998, DP_OP_423J2_125_3477_n997,
         DP_OP_423J2_125_3477_n996, DP_OP_423J2_125_3477_n995,
         DP_OP_423J2_125_3477_n994, DP_OP_423J2_125_3477_n993,
         DP_OP_423J2_125_3477_n992, DP_OP_423J2_125_3477_n991,
         DP_OP_423J2_125_3477_n990, DP_OP_423J2_125_3477_n989,
         DP_OP_423J2_125_3477_n988, DP_OP_423J2_125_3477_n987,
         DP_OP_423J2_125_3477_n986, DP_OP_423J2_125_3477_n985,
         DP_OP_423J2_125_3477_n984, DP_OP_423J2_125_3477_n983,
         DP_OP_423J2_125_3477_n982, DP_OP_423J2_125_3477_n981,
         DP_OP_423J2_125_3477_n980, DP_OP_423J2_125_3477_n979,
         DP_OP_423J2_125_3477_n978, DP_OP_423J2_125_3477_n977,
         DP_OP_423J2_125_3477_n976, DP_OP_423J2_125_3477_n975,
         DP_OP_423J2_125_3477_n974, DP_OP_423J2_125_3477_n973,
         DP_OP_423J2_125_3477_n972, DP_OP_423J2_125_3477_n971,
         DP_OP_423J2_125_3477_n970, DP_OP_423J2_125_3477_n969,
         DP_OP_423J2_125_3477_n968, DP_OP_423J2_125_3477_n967,
         DP_OP_423J2_125_3477_n965, DP_OP_423J2_125_3477_n964,
         DP_OP_423J2_125_3477_n963, DP_OP_423J2_125_3477_n962,
         DP_OP_423J2_125_3477_n961, DP_OP_423J2_125_3477_n960,
         DP_OP_423J2_125_3477_n959, DP_OP_423J2_125_3477_n958,
         DP_OP_423J2_125_3477_n957, DP_OP_423J2_125_3477_n956,
         DP_OP_423J2_125_3477_n955, DP_OP_423J2_125_3477_n954,
         DP_OP_423J2_125_3477_n953, DP_OP_423J2_125_3477_n952,
         DP_OP_423J2_125_3477_n951, DP_OP_423J2_125_3477_n950,
         DP_OP_423J2_125_3477_n949, DP_OP_423J2_125_3477_n948,
         DP_OP_423J2_125_3477_n947, DP_OP_423J2_125_3477_n946,
         DP_OP_423J2_125_3477_n945, DP_OP_423J2_125_3477_n944,
         DP_OP_423J2_125_3477_n943, DP_OP_423J2_125_3477_n942,
         DP_OP_423J2_125_3477_n941, DP_OP_423J2_125_3477_n940,
         DP_OP_423J2_125_3477_n939, DP_OP_423J2_125_3477_n938,
         DP_OP_423J2_125_3477_n937, DP_OP_423J2_125_3477_n936,
         DP_OP_423J2_125_3477_n935, DP_OP_423J2_125_3477_n934,
         DP_OP_423J2_125_3477_n933, DP_OP_423J2_125_3477_n932,
         DP_OP_423J2_125_3477_n931, DP_OP_423J2_125_3477_n930,
         DP_OP_423J2_125_3477_n929, DP_OP_423J2_125_3477_n928,
         DP_OP_423J2_125_3477_n927, DP_OP_423J2_125_3477_n926,
         DP_OP_423J2_125_3477_n925, DP_OP_423J2_125_3477_n924,
         DP_OP_423J2_125_3477_n923, DP_OP_423J2_125_3477_n922,
         DP_OP_423J2_125_3477_n921, DP_OP_423J2_125_3477_n920,
         DP_OP_423J2_125_3477_n919, DP_OP_423J2_125_3477_n918,
         DP_OP_423J2_125_3477_n917, DP_OP_423J2_125_3477_n916,
         DP_OP_423J2_125_3477_n915, DP_OP_423J2_125_3477_n914,
         DP_OP_423J2_125_3477_n913, DP_OP_423J2_125_3477_n911,
         DP_OP_423J2_125_3477_n910, DP_OP_423J2_125_3477_n909,
         DP_OP_423J2_125_3477_n908, DP_OP_423J2_125_3477_n907,
         DP_OP_423J2_125_3477_n906, DP_OP_423J2_125_3477_n905,
         DP_OP_423J2_125_3477_n904, DP_OP_423J2_125_3477_n903,
         DP_OP_423J2_125_3477_n902, DP_OP_423J2_125_3477_n901,
         DP_OP_423J2_125_3477_n900, DP_OP_423J2_125_3477_n899,
         DP_OP_423J2_125_3477_n898, DP_OP_423J2_125_3477_n897,
         DP_OP_423J2_125_3477_n896, DP_OP_423J2_125_3477_n895,
         DP_OP_423J2_125_3477_n894, DP_OP_423J2_125_3477_n893,
         DP_OP_423J2_125_3477_n892, DP_OP_423J2_125_3477_n891,
         DP_OP_423J2_125_3477_n890, DP_OP_423J2_125_3477_n889,
         DP_OP_423J2_125_3477_n888, DP_OP_423J2_125_3477_n887,
         DP_OP_423J2_125_3477_n886, DP_OP_423J2_125_3477_n885,
         DP_OP_423J2_125_3477_n884, DP_OP_423J2_125_3477_n883,
         DP_OP_423J2_125_3477_n882, DP_OP_423J2_125_3477_n881,
         DP_OP_423J2_125_3477_n880, DP_OP_423J2_125_3477_n879,
         DP_OP_423J2_125_3477_n878, DP_OP_423J2_125_3477_n877,
         DP_OP_423J2_125_3477_n876, DP_OP_423J2_125_3477_n875,
         DP_OP_423J2_125_3477_n874, DP_OP_423J2_125_3477_n873,
         DP_OP_423J2_125_3477_n872, DP_OP_423J2_125_3477_n871,
         DP_OP_423J2_125_3477_n870, DP_OP_423J2_125_3477_n869,
         DP_OP_423J2_125_3477_n868, DP_OP_423J2_125_3477_n867,
         DP_OP_423J2_125_3477_n866, DP_OP_423J2_125_3477_n865,
         DP_OP_423J2_125_3477_n864, DP_OP_423J2_125_3477_n863,
         DP_OP_423J2_125_3477_n862, DP_OP_423J2_125_3477_n861,
         DP_OP_423J2_125_3477_n860, DP_OP_423J2_125_3477_n859,
         DP_OP_423J2_125_3477_n858, DP_OP_423J2_125_3477_n857,
         DP_OP_423J2_125_3477_n856, DP_OP_423J2_125_3477_n855,
         DP_OP_423J2_125_3477_n854, DP_OP_423J2_125_3477_n853,
         DP_OP_423J2_125_3477_n852, DP_OP_423J2_125_3477_n851,
         DP_OP_423J2_125_3477_n850, DP_OP_423J2_125_3477_n849,
         DP_OP_423J2_125_3477_n848, DP_OP_423J2_125_3477_n847,
         DP_OP_423J2_125_3477_n846, DP_OP_423J2_125_3477_n845,
         DP_OP_423J2_125_3477_n844, DP_OP_423J2_125_3477_n843,
         DP_OP_423J2_125_3477_n842, DP_OP_423J2_125_3477_n841,
         DP_OP_423J2_125_3477_n840, DP_OP_423J2_125_3477_n839,
         DP_OP_423J2_125_3477_n838, DP_OP_423J2_125_3477_n837,
         DP_OP_423J2_125_3477_n836, DP_OP_423J2_125_3477_n835,
         DP_OP_423J2_125_3477_n834, DP_OP_423J2_125_3477_n833,
         DP_OP_423J2_125_3477_n832, DP_OP_423J2_125_3477_n831,
         DP_OP_423J2_125_3477_n830, DP_OP_423J2_125_3477_n829,
         DP_OP_423J2_125_3477_n828, DP_OP_423J2_125_3477_n827,
         DP_OP_423J2_125_3477_n826, DP_OP_423J2_125_3477_n825,
         DP_OP_423J2_125_3477_n824, DP_OP_423J2_125_3477_n823,
         DP_OP_423J2_125_3477_n822, DP_OP_423J2_125_3477_n821,
         DP_OP_423J2_125_3477_n820, DP_OP_423J2_125_3477_n819,
         DP_OP_423J2_125_3477_n818, DP_OP_423J2_125_3477_n817,
         DP_OP_423J2_125_3477_n816, DP_OP_423J2_125_3477_n815,
         DP_OP_423J2_125_3477_n814, DP_OP_423J2_125_3477_n813,
         DP_OP_423J2_125_3477_n812, DP_OP_423J2_125_3477_n811,
         DP_OP_423J2_125_3477_n810, DP_OP_423J2_125_3477_n809,
         DP_OP_423J2_125_3477_n808, DP_OP_423J2_125_3477_n807,
         DP_OP_423J2_125_3477_n806, DP_OP_423J2_125_3477_n805,
         DP_OP_423J2_125_3477_n804, DP_OP_423J2_125_3477_n803,
         DP_OP_423J2_125_3477_n802, DP_OP_423J2_125_3477_n801,
         DP_OP_423J2_125_3477_n800, DP_OP_423J2_125_3477_n799,
         DP_OP_423J2_125_3477_n798, DP_OP_423J2_125_3477_n797,
         DP_OP_423J2_125_3477_n796, DP_OP_423J2_125_3477_n795,
         DP_OP_423J2_125_3477_n794, DP_OP_423J2_125_3477_n793,
         DP_OP_423J2_125_3477_n792, DP_OP_423J2_125_3477_n791,
         DP_OP_423J2_125_3477_n790, DP_OP_423J2_125_3477_n789,
         DP_OP_423J2_125_3477_n788, DP_OP_423J2_125_3477_n787,
         DP_OP_423J2_125_3477_n786, DP_OP_423J2_125_3477_n785,
         DP_OP_423J2_125_3477_n784, DP_OP_423J2_125_3477_n783,
         DP_OP_423J2_125_3477_n782, DP_OP_423J2_125_3477_n781,
         DP_OP_423J2_125_3477_n780, DP_OP_423J2_125_3477_n779,
         DP_OP_423J2_125_3477_n778, DP_OP_423J2_125_3477_n777,
         DP_OP_423J2_125_3477_n776, DP_OP_423J2_125_3477_n775,
         DP_OP_423J2_125_3477_n774, DP_OP_423J2_125_3477_n773,
         DP_OP_423J2_125_3477_n772, DP_OP_423J2_125_3477_n771,
         DP_OP_423J2_125_3477_n770, DP_OP_423J2_125_3477_n769,
         DP_OP_423J2_125_3477_n768, DP_OP_423J2_125_3477_n767,
         DP_OP_423J2_125_3477_n766, DP_OP_423J2_125_3477_n765,
         DP_OP_423J2_125_3477_n764, DP_OP_423J2_125_3477_n763,
         DP_OP_423J2_125_3477_n762, DP_OP_423J2_125_3477_n761,
         DP_OP_423J2_125_3477_n760, DP_OP_423J2_125_3477_n759,
         DP_OP_423J2_125_3477_n758, DP_OP_423J2_125_3477_n757,
         DP_OP_423J2_125_3477_n756, DP_OP_423J2_125_3477_n755,
         DP_OP_423J2_125_3477_n754, DP_OP_423J2_125_3477_n753,
         DP_OP_423J2_125_3477_n752, DP_OP_423J2_125_3477_n751,
         DP_OP_423J2_125_3477_n750, DP_OP_423J2_125_3477_n749,
         DP_OP_423J2_125_3477_n748, DP_OP_423J2_125_3477_n747,
         DP_OP_423J2_125_3477_n746, DP_OP_423J2_125_3477_n745,
         DP_OP_423J2_125_3477_n744, DP_OP_423J2_125_3477_n743,
         DP_OP_423J2_125_3477_n742, DP_OP_423J2_125_3477_n741,
         DP_OP_423J2_125_3477_n740, DP_OP_423J2_125_3477_n739,
         DP_OP_423J2_125_3477_n738, DP_OP_423J2_125_3477_n737,
         DP_OP_423J2_125_3477_n736, DP_OP_423J2_125_3477_n735,
         DP_OP_423J2_125_3477_n734, DP_OP_423J2_125_3477_n733,
         DP_OP_423J2_125_3477_n732, DP_OP_423J2_125_3477_n731,
         DP_OP_423J2_125_3477_n730, DP_OP_423J2_125_3477_n729,
         DP_OP_423J2_125_3477_n728, DP_OP_423J2_125_3477_n727,
         DP_OP_423J2_125_3477_n726, DP_OP_423J2_125_3477_n725,
         DP_OP_423J2_125_3477_n724, DP_OP_423J2_125_3477_n723,
         DP_OP_423J2_125_3477_n722, DP_OP_423J2_125_3477_n721,
         DP_OP_423J2_125_3477_n720, DP_OP_423J2_125_3477_n719,
         DP_OP_423J2_125_3477_n718, DP_OP_423J2_125_3477_n717,
         DP_OP_423J2_125_3477_n716, DP_OP_423J2_125_3477_n715,
         DP_OP_423J2_125_3477_n714, DP_OP_423J2_125_3477_n713,
         DP_OP_423J2_125_3477_n712, DP_OP_423J2_125_3477_n711,
         DP_OP_423J2_125_3477_n710, DP_OP_423J2_125_3477_n709,
         DP_OP_423J2_125_3477_n708, DP_OP_423J2_125_3477_n707,
         DP_OP_423J2_125_3477_n706, DP_OP_423J2_125_3477_n705,
         DP_OP_423J2_125_3477_n704, DP_OP_423J2_125_3477_n703,
         DP_OP_423J2_125_3477_n702, DP_OP_423J2_125_3477_n701,
         DP_OP_423J2_125_3477_n700, DP_OP_423J2_125_3477_n699,
         DP_OP_423J2_125_3477_n698, DP_OP_423J2_125_3477_n697,
         DP_OP_423J2_125_3477_n696, DP_OP_423J2_125_3477_n695,
         DP_OP_423J2_125_3477_n694, DP_OP_423J2_125_3477_n693,
         DP_OP_423J2_125_3477_n692, DP_OP_423J2_125_3477_n691,
         DP_OP_423J2_125_3477_n690, DP_OP_423J2_125_3477_n689,
         DP_OP_423J2_125_3477_n688, DP_OP_423J2_125_3477_n687,
         DP_OP_423J2_125_3477_n686, DP_OP_423J2_125_3477_n685,
         DP_OP_423J2_125_3477_n684, DP_OP_423J2_125_3477_n683,
         DP_OP_423J2_125_3477_n682, DP_OP_423J2_125_3477_n681,
         DP_OP_423J2_125_3477_n680, DP_OP_423J2_125_3477_n679,
         DP_OP_423J2_125_3477_n678, DP_OP_423J2_125_3477_n677,
         DP_OP_423J2_125_3477_n676, DP_OP_423J2_125_3477_n675,
         DP_OP_423J2_125_3477_n674, DP_OP_423J2_125_3477_n673,
         DP_OP_423J2_125_3477_n672, DP_OP_423J2_125_3477_n671,
         DP_OP_423J2_125_3477_n670, DP_OP_423J2_125_3477_n669,
         DP_OP_423J2_125_3477_n668, DP_OP_423J2_125_3477_n667,
         DP_OP_423J2_125_3477_n666, DP_OP_423J2_125_3477_n665,
         DP_OP_423J2_125_3477_n664, DP_OP_423J2_125_3477_n663,
         DP_OP_423J2_125_3477_n662, DP_OP_423J2_125_3477_n661,
         DP_OP_423J2_125_3477_n660, DP_OP_423J2_125_3477_n659,
         DP_OP_423J2_125_3477_n658, DP_OP_423J2_125_3477_n657,
         DP_OP_423J2_125_3477_n656, DP_OP_423J2_125_3477_n655,
         DP_OP_423J2_125_3477_n654, DP_OP_423J2_125_3477_n653,
         DP_OP_423J2_125_3477_n652, DP_OP_423J2_125_3477_n651,
         DP_OP_423J2_125_3477_n650, DP_OP_423J2_125_3477_n649,
         DP_OP_423J2_125_3477_n648, DP_OP_423J2_125_3477_n647,
         DP_OP_423J2_125_3477_n646, DP_OP_423J2_125_3477_n645,
         DP_OP_423J2_125_3477_n644, DP_OP_423J2_125_3477_n643,
         DP_OP_423J2_125_3477_n642, DP_OP_423J2_125_3477_n641,
         DP_OP_423J2_125_3477_n640, DP_OP_423J2_125_3477_n639,
         DP_OP_423J2_125_3477_n638, DP_OP_423J2_125_3477_n637,
         DP_OP_423J2_125_3477_n636, DP_OP_423J2_125_3477_n635,
         DP_OP_423J2_125_3477_n634, DP_OP_423J2_125_3477_n633,
         DP_OP_423J2_125_3477_n632, DP_OP_423J2_125_3477_n631,
         DP_OP_423J2_125_3477_n630, DP_OP_423J2_125_3477_n629,
         DP_OP_423J2_125_3477_n628, DP_OP_423J2_125_3477_n627,
         DP_OP_423J2_125_3477_n626, DP_OP_423J2_125_3477_n625,
         DP_OP_423J2_125_3477_n624, DP_OP_423J2_125_3477_n623,
         DP_OP_423J2_125_3477_n622, DP_OP_423J2_125_3477_n621,
         DP_OP_423J2_125_3477_n620, DP_OP_423J2_125_3477_n619,
         DP_OP_423J2_125_3477_n618, DP_OP_423J2_125_3477_n617,
         DP_OP_423J2_125_3477_n616, DP_OP_423J2_125_3477_n615,
         DP_OP_423J2_125_3477_n614, DP_OP_423J2_125_3477_n613,
         DP_OP_423J2_125_3477_n612, DP_OP_423J2_125_3477_n611,
         DP_OP_423J2_125_3477_n610, DP_OP_423J2_125_3477_n609,
         DP_OP_423J2_125_3477_n608, DP_OP_423J2_125_3477_n607,
         DP_OP_423J2_125_3477_n606, DP_OP_423J2_125_3477_n605,
         DP_OP_423J2_125_3477_n604, DP_OP_423J2_125_3477_n603,
         DP_OP_423J2_125_3477_n602, DP_OP_423J2_125_3477_n601,
         DP_OP_423J2_125_3477_n600, DP_OP_423J2_125_3477_n599,
         DP_OP_423J2_125_3477_n598, DP_OP_423J2_125_3477_n597,
         DP_OP_423J2_125_3477_n596, DP_OP_423J2_125_3477_n595,
         DP_OP_423J2_125_3477_n594, DP_OP_423J2_125_3477_n593,
         DP_OP_423J2_125_3477_n592, DP_OP_423J2_125_3477_n591,
         DP_OP_423J2_125_3477_n590, DP_OP_423J2_125_3477_n589,
         DP_OP_423J2_125_3477_n588, DP_OP_423J2_125_3477_n587,
         DP_OP_423J2_125_3477_n586, DP_OP_423J2_125_3477_n585,
         DP_OP_423J2_125_3477_n584, DP_OP_423J2_125_3477_n583,
         DP_OP_423J2_125_3477_n582, DP_OP_423J2_125_3477_n581,
         DP_OP_423J2_125_3477_n580, DP_OP_423J2_125_3477_n579,
         DP_OP_423J2_125_3477_n578, DP_OP_423J2_125_3477_n577,
         DP_OP_423J2_125_3477_n576, DP_OP_423J2_125_3477_n575,
         DP_OP_423J2_125_3477_n574, DP_OP_423J2_125_3477_n573,
         DP_OP_423J2_125_3477_n572, DP_OP_423J2_125_3477_n571,
         DP_OP_423J2_125_3477_n570, DP_OP_423J2_125_3477_n569,
         DP_OP_423J2_125_3477_n568, DP_OP_423J2_125_3477_n567,
         DP_OP_423J2_125_3477_n566, DP_OP_423J2_125_3477_n565,
         DP_OP_423J2_125_3477_n564, DP_OP_423J2_125_3477_n563,
         DP_OP_423J2_125_3477_n562, DP_OP_423J2_125_3477_n561,
         DP_OP_423J2_125_3477_n560, DP_OP_423J2_125_3477_n559,
         DP_OP_423J2_125_3477_n558, DP_OP_423J2_125_3477_n557,
         DP_OP_423J2_125_3477_n556, DP_OP_423J2_125_3477_n555,
         DP_OP_423J2_125_3477_n554, DP_OP_423J2_125_3477_n553,
         DP_OP_423J2_125_3477_n552, DP_OP_423J2_125_3477_n551,
         DP_OP_423J2_125_3477_n550, DP_OP_423J2_125_3477_n549,
         DP_OP_423J2_125_3477_n548, DP_OP_423J2_125_3477_n547,
         DP_OP_423J2_125_3477_n546, DP_OP_423J2_125_3477_n545,
         DP_OP_423J2_125_3477_n544, DP_OP_423J2_125_3477_n543,
         DP_OP_423J2_125_3477_n542, DP_OP_423J2_125_3477_n541,
         DP_OP_423J2_125_3477_n540, DP_OP_423J2_125_3477_n539,
         DP_OP_423J2_125_3477_n538, DP_OP_423J2_125_3477_n537,
         DP_OP_423J2_125_3477_n536, DP_OP_423J2_125_3477_n535,
         DP_OP_423J2_125_3477_n534, DP_OP_423J2_125_3477_n533,
         DP_OP_423J2_125_3477_n532, DP_OP_423J2_125_3477_n531,
         DP_OP_423J2_125_3477_n530, DP_OP_423J2_125_3477_n529,
         DP_OP_423J2_125_3477_n528, DP_OP_423J2_125_3477_n527,
         DP_OP_423J2_125_3477_n526, DP_OP_423J2_125_3477_n525,
         DP_OP_423J2_125_3477_n524, DP_OP_423J2_125_3477_n523,
         DP_OP_423J2_125_3477_n522, DP_OP_423J2_125_3477_n521,
         DP_OP_423J2_125_3477_n520, DP_OP_423J2_125_3477_n519,
         DP_OP_423J2_125_3477_n518, DP_OP_423J2_125_3477_n517,
         DP_OP_423J2_125_3477_n516, DP_OP_423J2_125_3477_n515,
         DP_OP_423J2_125_3477_n514, DP_OP_423J2_125_3477_n513,
         DP_OP_423J2_125_3477_n512, DP_OP_423J2_125_3477_n511,
         DP_OP_423J2_125_3477_n510, DP_OP_423J2_125_3477_n509,
         DP_OP_423J2_125_3477_n508, DP_OP_423J2_125_3477_n507,
         DP_OP_423J2_125_3477_n506, DP_OP_423J2_125_3477_n505,
         DP_OP_423J2_125_3477_n504, DP_OP_423J2_125_3477_n503,
         DP_OP_423J2_125_3477_n502, DP_OP_423J2_125_3477_n501,
         DP_OP_423J2_125_3477_n500, DP_OP_423J2_125_3477_n499,
         DP_OP_423J2_125_3477_n498, DP_OP_423J2_125_3477_n497,
         DP_OP_423J2_125_3477_n496, DP_OP_423J2_125_3477_n495,
         DP_OP_423J2_125_3477_n494, DP_OP_423J2_125_3477_n493,
         DP_OP_423J2_125_3477_n492, DP_OP_423J2_125_3477_n491,
         DP_OP_423J2_125_3477_n490, DP_OP_423J2_125_3477_n489,
         DP_OP_423J2_125_3477_n488, DP_OP_423J2_125_3477_n487,
         DP_OP_423J2_125_3477_n486, DP_OP_423J2_125_3477_n485,
         DP_OP_423J2_125_3477_n484, DP_OP_423J2_125_3477_n483,
         DP_OP_423J2_125_3477_n482, DP_OP_423J2_125_3477_n481,
         DP_OP_423J2_125_3477_n480, DP_OP_423J2_125_3477_n479,
         DP_OP_423J2_125_3477_n478, DP_OP_423J2_125_3477_n477,
         DP_OP_423J2_125_3477_n476, DP_OP_423J2_125_3477_n475,
         DP_OP_423J2_125_3477_n474, DP_OP_423J2_125_3477_n473,
         DP_OP_423J2_125_3477_n472, DP_OP_423J2_125_3477_n471,
         DP_OP_423J2_125_3477_n470, DP_OP_423J2_125_3477_n469,
         DP_OP_423J2_125_3477_n468, DP_OP_423J2_125_3477_n467,
         DP_OP_423J2_125_3477_n466, DP_OP_423J2_125_3477_n465,
         DP_OP_423J2_125_3477_n464, DP_OP_423J2_125_3477_n463,
         DP_OP_423J2_125_3477_n462, DP_OP_423J2_125_3477_n461,
         DP_OP_423J2_125_3477_n460, DP_OP_423J2_125_3477_n459,
         DP_OP_423J2_125_3477_n458, DP_OP_423J2_125_3477_n457,
         DP_OP_423J2_125_3477_n456, DP_OP_423J2_125_3477_n455,
         DP_OP_423J2_125_3477_n454, DP_OP_423J2_125_3477_n453,
         DP_OP_423J2_125_3477_n452, DP_OP_423J2_125_3477_n451,
         DP_OP_423J2_125_3477_n450, DP_OP_423J2_125_3477_n449,
         DP_OP_423J2_125_3477_n448, DP_OP_423J2_125_3477_n447,
         DP_OP_423J2_125_3477_n446, DP_OP_423J2_125_3477_n445,
         DP_OP_423J2_125_3477_n444, DP_OP_423J2_125_3477_n443,
         DP_OP_423J2_125_3477_n442, DP_OP_423J2_125_3477_n441,
         DP_OP_423J2_125_3477_n440, DP_OP_423J2_125_3477_n439,
         DP_OP_423J2_125_3477_n438, DP_OP_423J2_125_3477_n437,
         DP_OP_423J2_125_3477_n436, DP_OP_423J2_125_3477_n435,
         DP_OP_423J2_125_3477_n434, DP_OP_423J2_125_3477_n433,
         DP_OP_423J2_125_3477_n432, DP_OP_423J2_125_3477_n431,
         DP_OP_423J2_125_3477_n430, DP_OP_423J2_125_3477_n429,
         DP_OP_423J2_125_3477_n428, DP_OP_423J2_125_3477_n427,
         DP_OP_423J2_125_3477_n426, DP_OP_423J2_125_3477_n425,
         DP_OP_423J2_125_3477_n424, DP_OP_423J2_125_3477_n423,
         DP_OP_423J2_125_3477_n422, DP_OP_423J2_125_3477_n421,
         DP_OP_423J2_125_3477_n420, DP_OP_423J2_125_3477_n419,
         DP_OP_423J2_125_3477_n418, DP_OP_423J2_125_3477_n417,
         DP_OP_423J2_125_3477_n416, DP_OP_423J2_125_3477_n415,
         DP_OP_423J2_125_3477_n414, DP_OP_423J2_125_3477_n413,
         DP_OP_423J2_125_3477_n412, DP_OP_423J2_125_3477_n411,
         DP_OP_423J2_125_3477_n410, DP_OP_423J2_125_3477_n409,
         DP_OP_423J2_125_3477_n408, DP_OP_423J2_125_3477_n407,
         DP_OP_423J2_125_3477_n406, DP_OP_423J2_125_3477_n405,
         DP_OP_423J2_125_3477_n404, DP_OP_423J2_125_3477_n403,
         DP_OP_423J2_125_3477_n402, DP_OP_423J2_125_3477_n401,
         DP_OP_423J2_125_3477_n400, DP_OP_423J2_125_3477_n399,
         DP_OP_423J2_125_3477_n398, DP_OP_423J2_125_3477_n397,
         DP_OP_423J2_125_3477_n396, DP_OP_423J2_125_3477_n395,
         DP_OP_423J2_125_3477_n394, DP_OP_423J2_125_3477_n393,
         DP_OP_423J2_125_3477_n392, DP_OP_423J2_125_3477_n391,
         DP_OP_423J2_125_3477_n390, DP_OP_423J2_125_3477_n389,
         DP_OP_423J2_125_3477_n388, DP_OP_423J2_125_3477_n387,
         DP_OP_423J2_125_3477_n386, DP_OP_423J2_125_3477_n385,
         DP_OP_423J2_125_3477_n384, DP_OP_423J2_125_3477_n383,
         DP_OP_423J2_125_3477_n382, DP_OP_423J2_125_3477_n381,
         DP_OP_423J2_125_3477_n380, DP_OP_423J2_125_3477_n379,
         DP_OP_423J2_125_3477_n378, DP_OP_423J2_125_3477_n377,
         DP_OP_423J2_125_3477_n376, DP_OP_423J2_125_3477_n375,
         DP_OP_423J2_125_3477_n374, DP_OP_423J2_125_3477_n373,
         DP_OP_423J2_125_3477_n372, DP_OP_423J2_125_3477_n371,
         DP_OP_423J2_125_3477_n370, DP_OP_423J2_125_3477_n369,
         DP_OP_423J2_125_3477_n368, DP_OP_423J2_125_3477_n367,
         DP_OP_423J2_125_3477_n366, DP_OP_423J2_125_3477_n365,
         DP_OP_423J2_125_3477_n364, DP_OP_423J2_125_3477_n363,
         DP_OP_423J2_125_3477_n362, DP_OP_423J2_125_3477_n361,
         DP_OP_423J2_125_3477_n360, DP_OP_423J2_125_3477_n359,
         DP_OP_423J2_125_3477_n358, DP_OP_423J2_125_3477_n357,
         DP_OP_423J2_125_3477_n356, DP_OP_423J2_125_3477_n355,
         DP_OP_423J2_125_3477_n354, DP_OP_423J2_125_3477_n353,
         DP_OP_423J2_125_3477_n352, DP_OP_423J2_125_3477_n351,
         DP_OP_423J2_125_3477_n350, DP_OP_423J2_125_3477_n349,
         DP_OP_423J2_125_3477_n348, DP_OP_423J2_125_3477_n347,
         DP_OP_423J2_125_3477_n346, DP_OP_423J2_125_3477_n345,
         DP_OP_423J2_125_3477_n344, DP_OP_423J2_125_3477_n343,
         DP_OP_423J2_125_3477_n342, DP_OP_423J2_125_3477_n341,
         DP_OP_423J2_125_3477_n340, DP_OP_423J2_125_3477_n339,
         DP_OP_423J2_125_3477_n338, DP_OP_423J2_125_3477_n337,
         DP_OP_423J2_125_3477_n336, DP_OP_423J2_125_3477_n335,
         DP_OP_423J2_125_3477_n334, DP_OP_423J2_125_3477_n333,
         DP_OP_423J2_125_3477_n332, DP_OP_423J2_125_3477_n331,
         DP_OP_423J2_125_3477_n330, DP_OP_423J2_125_3477_n329,
         DP_OP_423J2_125_3477_n328, DP_OP_423J2_125_3477_n327,
         DP_OP_423J2_125_3477_n326, DP_OP_423J2_125_3477_n325,
         DP_OP_423J2_125_3477_n324, DP_OP_423J2_125_3477_n323,
         DP_OP_423J2_125_3477_n322, DP_OP_423J2_125_3477_n321,
         DP_OP_423J2_125_3477_n320, DP_OP_423J2_125_3477_n319,
         DP_OP_423J2_125_3477_n318, DP_OP_423J2_125_3477_n317,
         DP_OP_423J2_125_3477_n316, DP_OP_423J2_125_3477_n315,
         DP_OP_423J2_125_3477_n314, DP_OP_423J2_125_3477_n312,
         DP_OP_423J2_125_3477_n311, DP_OP_423J2_125_3477_n310,
         DP_OP_423J2_125_3477_n309, DP_OP_423J2_125_3477_n308,
         DP_OP_423J2_125_3477_n307, DP_OP_423J2_125_3477_n306,
         DP_OP_423J2_125_3477_n305, DP_OP_423J2_125_3477_n304,
         DP_OP_423J2_125_3477_n303, DP_OP_423J2_125_3477_n302,
         DP_OP_423J2_125_3477_n295, DP_OP_423J2_125_3477_n286,
         DP_OP_423J2_125_3477_n285, DP_OP_423J2_125_3477_n284,
         DP_OP_423J2_125_3477_n283, DP_OP_423J2_125_3477_n282,
         DP_OP_423J2_125_3477_n281, DP_OP_423J2_125_3477_n280,
         DP_OP_423J2_125_3477_n279, DP_OP_423J2_125_3477_n277,
         DP_OP_423J2_125_3477_n276, DP_OP_423J2_125_3477_n274,
         DP_OP_423J2_125_3477_n272, DP_OP_423J2_125_3477_n269,
         DP_OP_423J2_125_3477_n268, DP_OP_423J2_125_3477_n267,
         DP_OP_423J2_125_3477_n266, DP_OP_423J2_125_3477_n265,
         DP_OP_423J2_125_3477_n261, DP_OP_423J2_125_3477_n260,
         DP_OP_423J2_125_3477_n259, DP_OP_423J2_125_3477_n257,
         DP_OP_423J2_125_3477_n256, DP_OP_423J2_125_3477_n253,
         DP_OP_423J2_125_3477_n252, DP_OP_423J2_125_3477_n250,
         DP_OP_423J2_125_3477_n249, DP_OP_423J2_125_3477_n244,
         DP_OP_423J2_125_3477_n241, DP_OP_423J2_125_3477_n240,
         DP_OP_423J2_125_3477_n237, DP_OP_423J2_125_3477_n226,
         DP_OP_423J2_125_3477_n222, DP_OP_423J2_125_3477_n220,
         DP_OP_423J2_125_3477_n217, DP_OP_423J2_125_3477_n214,
         DP_OP_423J2_125_3477_n213, DP_OP_423J2_125_3477_n212,
         DP_OP_423J2_125_3477_n210, DP_OP_423J2_125_3477_n209,
         DP_OP_423J2_125_3477_n198, DP_OP_423J2_125_3477_n197,
         DP_OP_423J2_125_3477_n190, DP_OP_423J2_125_3477_n189,
         DP_OP_423J2_125_3477_n188, DP_OP_423J2_125_3477_n187,
         DP_OP_423J2_125_3477_n185, DP_OP_423J2_125_3477_n182,
         DP_OP_423J2_125_3477_n179, DP_OP_423J2_125_3477_n178,
         DP_OP_423J2_125_3477_n177, DP_OP_423J2_125_3477_n176,
         DP_OP_423J2_125_3477_n174, DP_OP_423J2_125_3477_n171,
         DP_OP_423J2_125_3477_n167, DP_OP_423J2_125_3477_n166,
         DP_OP_423J2_125_3477_n165, DP_OP_423J2_125_3477_n162,
         DP_OP_423J2_125_3477_n161, DP_OP_423J2_125_3477_n160,
         DP_OP_423J2_125_3477_n159, DP_OP_423J2_125_3477_n158,
         DP_OP_423J2_125_3477_n156, DP_OP_423J2_125_3477_n153,
         DP_OP_423J2_125_3477_n151, DP_OP_423J2_125_3477_n149,
         DP_OP_423J2_125_3477_n148, DP_OP_423J2_125_3477_n146,
         DP_OP_423J2_125_3477_n145, DP_OP_423J2_125_3477_n144,
         DP_OP_423J2_125_3477_n142, DP_OP_423J2_125_3477_n141,
         DP_OP_423J2_125_3477_n140, DP_OP_423J2_125_3477_n138,
         DP_OP_423J2_125_3477_n136, DP_OP_423J2_125_3477_n133,
         DP_OP_423J2_125_3477_n131, DP_OP_423J2_125_3477_n129,
         DP_OP_423J2_125_3477_n128, DP_OP_423J2_125_3477_n127,
         DP_OP_423J2_125_3477_n126, DP_OP_423J2_125_3477_n125,
         DP_OP_423J2_125_3477_n124, DP_OP_423J2_125_3477_n122,
         DP_OP_423J2_125_3477_n120, DP_OP_423J2_125_3477_n115,
         DP_OP_423J2_125_3477_n114, DP_OP_423J2_125_3477_n111,
         DP_OP_423J2_125_3477_n110, DP_OP_423J2_125_3477_n109,
         DP_OP_423J2_125_3477_n108, DP_OP_423J2_125_3477_n107,
         DP_OP_423J2_125_3477_n105, DP_OP_423J2_125_3477_n102,
         DP_OP_423J2_125_3477_n101, DP_OP_423J2_125_3477_n100,
         DP_OP_423J2_125_3477_n98, DP_OP_423J2_125_3477_n97,
         DP_OP_423J2_125_3477_n96, DP_OP_423J2_125_3477_n95,
         DP_OP_423J2_125_3477_n94, DP_OP_423J2_125_3477_n93,
         DP_OP_423J2_125_3477_n92, DP_OP_423J2_125_3477_n91,
         DP_OP_423J2_125_3477_n89, DP_OP_423J2_125_3477_n85,
         DP_OP_423J2_125_3477_n82, DP_OP_423J2_125_3477_n81,
         DP_OP_423J2_125_3477_n80, DP_OP_423J2_125_3477_n78,
         DP_OP_423J2_125_3477_n77, DP_OP_423J2_125_3477_n75,
         DP_OP_423J2_125_3477_n73, DP_OP_423J2_125_3477_n72,
         DP_OP_423J2_125_3477_n71, DP_OP_423J2_125_3477_n69,
         DP_OP_423J2_125_3477_n68, DP_OP_423J2_125_3477_n67,
         DP_OP_423J2_125_3477_n65, DP_OP_423J2_125_3477_n60,
         DP_OP_423J2_125_3477_n58, DP_OP_423J2_125_3477_n57,
         DP_OP_423J2_125_3477_n56, DP_OP_423J2_125_3477_n55,
         DP_OP_423J2_125_3477_n54, DP_OP_423J2_125_3477_n52,
         DP_OP_423J2_125_3477_n51, DP_OP_423J2_125_3477_n50,
         DP_OP_423J2_125_3477_n49, DP_OP_423J2_125_3477_n47,
         DP_OP_423J2_125_3477_n38, DP_OP_423J2_125_3477_n22,
         DP_OP_423J2_125_3477_n21, DP_OP_423J2_125_3477_n20,
         DP_OP_423J2_125_3477_n19, DP_OP_423J2_125_3477_n18,
         DP_OP_423J2_125_3477_n17, DP_OP_423J2_125_3477_n16,
         DP_OP_423J2_125_3477_n14, DP_OP_423J2_125_3477_n13,
         DP_OP_423J2_125_3477_n9, DP_OP_423J2_125_3477_n8,
         DP_OP_423J2_125_3477_n7, DP_OP_423J2_125_3477_n5,
         DP_OP_423J2_125_3477_n4, DP_OP_422J2_124_3477_n3064,
         DP_OP_422J2_124_3477_n3063, DP_OP_422J2_124_3477_n3060,
         DP_OP_422J2_124_3477_n3059, DP_OP_422J2_124_3477_n3058,
         DP_OP_422J2_124_3477_n3057, DP_OP_422J2_124_3477_n3056,
         DP_OP_422J2_124_3477_n3055, DP_OP_422J2_124_3477_n3054,
         DP_OP_422J2_124_3477_n3053, DP_OP_422J2_124_3477_n3052,
         DP_OP_422J2_124_3477_n3051, DP_OP_422J2_124_3477_n3050,
         DP_OP_422J2_124_3477_n3049, DP_OP_422J2_124_3477_n3048,
         DP_OP_422J2_124_3477_n3047, DP_OP_422J2_124_3477_n3046,
         DP_OP_422J2_124_3477_n3045, DP_OP_422J2_124_3477_n3044,
         DP_OP_422J2_124_3477_n3043, DP_OP_422J2_124_3477_n3042,
         DP_OP_422J2_124_3477_n3041, DP_OP_422J2_124_3477_n3040,
         DP_OP_422J2_124_3477_n3039, DP_OP_422J2_124_3477_n3038,
         DP_OP_422J2_124_3477_n3037, DP_OP_422J2_124_3477_n3036,
         DP_OP_422J2_124_3477_n3035, DP_OP_422J2_124_3477_n3034,
         DP_OP_422J2_124_3477_n3033, DP_OP_422J2_124_3477_n3032,
         DP_OP_422J2_124_3477_n3031, DP_OP_422J2_124_3477_n3030,
         DP_OP_422J2_124_3477_n3029, DP_OP_422J2_124_3477_n3028,
         DP_OP_422J2_124_3477_n3027, DP_OP_422J2_124_3477_n3026,
         DP_OP_422J2_124_3477_n3023, DP_OP_422J2_124_3477_n3021,
         DP_OP_422J2_124_3477_n3019, DP_OP_422J2_124_3477_n3017,
         DP_OP_422J2_124_3477_n3015, DP_OP_422J2_124_3477_n3014,
         DP_OP_422J2_124_3477_n3013, DP_OP_422J2_124_3477_n3012,
         DP_OP_422J2_124_3477_n3011, DP_OP_422J2_124_3477_n3010,
         DP_OP_422J2_124_3477_n3009, DP_OP_422J2_124_3477_n3008,
         DP_OP_422J2_124_3477_n3007, DP_OP_422J2_124_3477_n3006,
         DP_OP_422J2_124_3477_n3005, DP_OP_422J2_124_3477_n3004,
         DP_OP_422J2_124_3477_n3003, DP_OP_422J2_124_3477_n3002,
         DP_OP_422J2_124_3477_n3001, DP_OP_422J2_124_3477_n3000,
         DP_OP_422J2_124_3477_n2999, DP_OP_422J2_124_3477_n2998,
         DP_OP_422J2_124_3477_n2997, DP_OP_422J2_124_3477_n2996,
         DP_OP_422J2_124_3477_n2995, DP_OP_422J2_124_3477_n2994,
         DP_OP_422J2_124_3477_n2993, DP_OP_422J2_124_3477_n2992,
         DP_OP_422J2_124_3477_n2991, DP_OP_422J2_124_3477_n2990,
         DP_OP_422J2_124_3477_n2989, DP_OP_422J2_124_3477_n2988,
         DP_OP_422J2_124_3477_n2987, DP_OP_422J2_124_3477_n2986,
         DP_OP_422J2_124_3477_n2985, DP_OP_422J2_124_3477_n2984,
         DP_OP_422J2_124_3477_n2983, DP_OP_422J2_124_3477_n2982,
         DP_OP_422J2_124_3477_n2980, DP_OP_422J2_124_3477_n2975,
         DP_OP_422J2_124_3477_n2974, DP_OP_422J2_124_3477_n2973,
         DP_OP_422J2_124_3477_n2972, DP_OP_422J2_124_3477_n2971,
         DP_OP_422J2_124_3477_n2970, DP_OP_422J2_124_3477_n2969,
         DP_OP_422J2_124_3477_n2968, DP_OP_422J2_124_3477_n2967,
         DP_OP_422J2_124_3477_n2966, DP_OP_422J2_124_3477_n2965,
         DP_OP_422J2_124_3477_n2964, DP_OP_422J2_124_3477_n2963,
         DP_OP_422J2_124_3477_n2962, DP_OP_422J2_124_3477_n2961,
         DP_OP_422J2_124_3477_n2960, DP_OP_422J2_124_3477_n2959,
         DP_OP_422J2_124_3477_n2958, DP_OP_422J2_124_3477_n2957,
         DP_OP_422J2_124_3477_n2956, DP_OP_422J2_124_3477_n2955,
         DP_OP_422J2_124_3477_n2954, DP_OP_422J2_124_3477_n2953,
         DP_OP_422J2_124_3477_n2952, DP_OP_422J2_124_3477_n2951,
         DP_OP_422J2_124_3477_n2950, DP_OP_422J2_124_3477_n2949,
         DP_OP_422J2_124_3477_n2948, DP_OP_422J2_124_3477_n2947,
         DP_OP_422J2_124_3477_n2946, DP_OP_422J2_124_3477_n2945,
         DP_OP_422J2_124_3477_n2944, DP_OP_422J2_124_3477_n2943,
         DP_OP_422J2_124_3477_n2942, DP_OP_422J2_124_3477_n2941,
         DP_OP_422J2_124_3477_n2940, DP_OP_422J2_124_3477_n2939,
         DP_OP_422J2_124_3477_n2938, DP_OP_422J2_124_3477_n2937,
         DP_OP_422J2_124_3477_n2935, DP_OP_422J2_124_3477_n2930,
         DP_OP_422J2_124_3477_n2929, DP_OP_422J2_124_3477_n2928,
         DP_OP_422J2_124_3477_n2927, DP_OP_422J2_124_3477_n2926,
         DP_OP_422J2_124_3477_n2925, DP_OP_422J2_124_3477_n2924,
         DP_OP_422J2_124_3477_n2923, DP_OP_422J2_124_3477_n2922,
         DP_OP_422J2_124_3477_n2921, DP_OP_422J2_124_3477_n2920,
         DP_OP_422J2_124_3477_n2919, DP_OP_422J2_124_3477_n2918,
         DP_OP_422J2_124_3477_n2917, DP_OP_422J2_124_3477_n2916,
         DP_OP_422J2_124_3477_n2915, DP_OP_422J2_124_3477_n2914,
         DP_OP_422J2_124_3477_n2913, DP_OP_422J2_124_3477_n2912,
         DP_OP_422J2_124_3477_n2911, DP_OP_422J2_124_3477_n2910,
         DP_OP_422J2_124_3477_n2909, DP_OP_422J2_124_3477_n2908,
         DP_OP_422J2_124_3477_n2907, DP_OP_422J2_124_3477_n2906,
         DP_OP_422J2_124_3477_n2905, DP_OP_422J2_124_3477_n2904,
         DP_OP_422J2_124_3477_n2903, DP_OP_422J2_124_3477_n2902,
         DP_OP_422J2_124_3477_n2900, DP_OP_422J2_124_3477_n2899,
         DP_OP_422J2_124_3477_n2898, DP_OP_422J2_124_3477_n2897,
         DP_OP_422J2_124_3477_n2896, DP_OP_422J2_124_3477_n2895,
         DP_OP_422J2_124_3477_n2894, DP_OP_422J2_124_3477_n2893,
         DP_OP_422J2_124_3477_n2890, DP_OP_422J2_124_3477_n2889,
         DP_OP_422J2_124_3477_n2888, DP_OP_422J2_124_3477_n2887,
         DP_OP_422J2_124_3477_n2885, DP_OP_422J2_124_3477_n2884,
         DP_OP_422J2_124_3477_n2883, DP_OP_422J2_124_3477_n2882,
         DP_OP_422J2_124_3477_n2881, DP_OP_422J2_124_3477_n2880,
         DP_OP_422J2_124_3477_n2879, DP_OP_422J2_124_3477_n2878,
         DP_OP_422J2_124_3477_n2877, DP_OP_422J2_124_3477_n2876,
         DP_OP_422J2_124_3477_n2875, DP_OP_422J2_124_3477_n2874,
         DP_OP_422J2_124_3477_n2873, DP_OP_422J2_124_3477_n2872,
         DP_OP_422J2_124_3477_n2871, DP_OP_422J2_124_3477_n2870,
         DP_OP_422J2_124_3477_n2869, DP_OP_422J2_124_3477_n2868,
         DP_OP_422J2_124_3477_n2867, DP_OP_422J2_124_3477_n2866,
         DP_OP_422J2_124_3477_n2865, DP_OP_422J2_124_3477_n2864,
         DP_OP_422J2_124_3477_n2863, DP_OP_422J2_124_3477_n2862,
         DP_OP_422J2_124_3477_n2861, DP_OP_422J2_124_3477_n2860,
         DP_OP_422J2_124_3477_n2859, DP_OP_422J2_124_3477_n2858,
         DP_OP_422J2_124_3477_n2857, DP_OP_422J2_124_3477_n2856,
         DP_OP_422J2_124_3477_n2855, DP_OP_422J2_124_3477_n2854,
         DP_OP_422J2_124_3477_n2853, DP_OP_422J2_124_3477_n2852,
         DP_OP_422J2_124_3477_n2851, DP_OP_422J2_124_3477_n2850,
         DP_OP_422J2_124_3477_n2847, DP_OP_422J2_124_3477_n2846,
         DP_OP_422J2_124_3477_n2842, DP_OP_422J2_124_3477_n2841,
         DP_OP_422J2_124_3477_n2840, DP_OP_422J2_124_3477_n2839,
         DP_OP_422J2_124_3477_n2838, DP_OP_422J2_124_3477_n2837,
         DP_OP_422J2_124_3477_n2836, DP_OP_422J2_124_3477_n2835,
         DP_OP_422J2_124_3477_n2834, DP_OP_422J2_124_3477_n2833,
         DP_OP_422J2_124_3477_n2832, DP_OP_422J2_124_3477_n2831,
         DP_OP_422J2_124_3477_n2830, DP_OP_422J2_124_3477_n2829,
         DP_OP_422J2_124_3477_n2828, DP_OP_422J2_124_3477_n2827,
         DP_OP_422J2_124_3477_n2826, DP_OP_422J2_124_3477_n2825,
         DP_OP_422J2_124_3477_n2824, DP_OP_422J2_124_3477_n2823,
         DP_OP_422J2_124_3477_n2822, DP_OP_422J2_124_3477_n2821,
         DP_OP_422J2_124_3477_n2820, DP_OP_422J2_124_3477_n2819,
         DP_OP_422J2_124_3477_n2818, DP_OP_422J2_124_3477_n2817,
         DP_OP_422J2_124_3477_n2816, DP_OP_422J2_124_3477_n2815,
         DP_OP_422J2_124_3477_n2814, DP_OP_422J2_124_3477_n2813,
         DP_OP_422J2_124_3477_n2812, DP_OP_422J2_124_3477_n2811,
         DP_OP_422J2_124_3477_n2810, DP_OP_422J2_124_3477_n2809,
         DP_OP_422J2_124_3477_n2808, DP_OP_422J2_124_3477_n2807,
         DP_OP_422J2_124_3477_n2806, DP_OP_422J2_124_3477_n2805,
         DP_OP_422J2_124_3477_n2803, DP_OP_422J2_124_3477_n2801,
         DP_OP_422J2_124_3477_n2800, DP_OP_422J2_124_3477_n2799,
         DP_OP_422J2_124_3477_n2798, DP_OP_422J2_124_3477_n2797,
         DP_OP_422J2_124_3477_n2796, DP_OP_422J2_124_3477_n2795,
         DP_OP_422J2_124_3477_n2794, DP_OP_422J2_124_3477_n2793,
         DP_OP_422J2_124_3477_n2792, DP_OP_422J2_124_3477_n2791,
         DP_OP_422J2_124_3477_n2790, DP_OP_422J2_124_3477_n2789,
         DP_OP_422J2_124_3477_n2788, DP_OP_422J2_124_3477_n2787,
         DP_OP_422J2_124_3477_n2786, DP_OP_422J2_124_3477_n2785,
         DP_OP_422J2_124_3477_n2784, DP_OP_422J2_124_3477_n2783,
         DP_OP_422J2_124_3477_n2782, DP_OP_422J2_124_3477_n2781,
         DP_OP_422J2_124_3477_n2780, DP_OP_422J2_124_3477_n2779,
         DP_OP_422J2_124_3477_n2778, DP_OP_422J2_124_3477_n2777,
         DP_OP_422J2_124_3477_n2776, DP_OP_422J2_124_3477_n2775,
         DP_OP_422J2_124_3477_n2774, DP_OP_422J2_124_3477_n2773,
         DP_OP_422J2_124_3477_n2772, DP_OP_422J2_124_3477_n2771,
         DP_OP_422J2_124_3477_n2770, DP_OP_422J2_124_3477_n2768,
         DP_OP_422J2_124_3477_n2767, DP_OP_422J2_124_3477_n2766,
         DP_OP_422J2_124_3477_n2765, DP_OP_422J2_124_3477_n2764,
         DP_OP_422J2_124_3477_n2763, DP_OP_422J2_124_3477_n2762,
         DP_OP_422J2_124_3477_n2759, DP_OP_422J2_124_3477_n2758,
         DP_OP_422J2_124_3477_n2756, DP_OP_422J2_124_3477_n2754,
         DP_OP_422J2_124_3477_n2753, DP_OP_422J2_124_3477_n2751,
         DP_OP_422J2_124_3477_n2750, DP_OP_422J2_124_3477_n2749,
         DP_OP_422J2_124_3477_n2748, DP_OP_422J2_124_3477_n2747,
         DP_OP_422J2_124_3477_n2746, DP_OP_422J2_124_3477_n2745,
         DP_OP_422J2_124_3477_n2744, DP_OP_422J2_124_3477_n2743,
         DP_OP_422J2_124_3477_n2742, DP_OP_422J2_124_3477_n2741,
         DP_OP_422J2_124_3477_n2740, DP_OP_422J2_124_3477_n2739,
         DP_OP_422J2_124_3477_n2738, DP_OP_422J2_124_3477_n2737,
         DP_OP_422J2_124_3477_n2736, DP_OP_422J2_124_3477_n2735,
         DP_OP_422J2_124_3477_n2734, DP_OP_422J2_124_3477_n2733,
         DP_OP_422J2_124_3477_n2732, DP_OP_422J2_124_3477_n2731,
         DP_OP_422J2_124_3477_n2730, DP_OP_422J2_124_3477_n2729,
         DP_OP_422J2_124_3477_n2728, DP_OP_422J2_124_3477_n2727,
         DP_OP_422J2_124_3477_n2726, DP_OP_422J2_124_3477_n2725,
         DP_OP_422J2_124_3477_n2724, DP_OP_422J2_124_3477_n2723,
         DP_OP_422J2_124_3477_n2722, DP_OP_422J2_124_3477_n2721,
         DP_OP_422J2_124_3477_n2720, DP_OP_422J2_124_3477_n2719,
         DP_OP_422J2_124_3477_n2718, DP_OP_422J2_124_3477_n2717,
         DP_OP_422J2_124_3477_n2715, DP_OP_422J2_124_3477_n2714,
         DP_OP_422J2_124_3477_n2712, DP_OP_422J2_124_3477_n2710,
         DP_OP_422J2_124_3477_n2709, DP_OP_422J2_124_3477_n2708,
         DP_OP_422J2_124_3477_n2707, DP_OP_422J2_124_3477_n2705,
         DP_OP_422J2_124_3477_n2704, DP_OP_422J2_124_3477_n2703,
         DP_OP_422J2_124_3477_n2702, DP_OP_422J2_124_3477_n2701,
         DP_OP_422J2_124_3477_n2700, DP_OP_422J2_124_3477_n2699,
         DP_OP_422J2_124_3477_n2698, DP_OP_422J2_124_3477_n2697,
         DP_OP_422J2_124_3477_n2696, DP_OP_422J2_124_3477_n2695,
         DP_OP_422J2_124_3477_n2694, DP_OP_422J2_124_3477_n2693,
         DP_OP_422J2_124_3477_n2692, DP_OP_422J2_124_3477_n2691,
         DP_OP_422J2_124_3477_n2690, DP_OP_422J2_124_3477_n2689,
         DP_OP_422J2_124_3477_n2688, DP_OP_422J2_124_3477_n2687,
         DP_OP_422J2_124_3477_n2686, DP_OP_422J2_124_3477_n2685,
         DP_OP_422J2_124_3477_n2684, DP_OP_422J2_124_3477_n2683,
         DP_OP_422J2_124_3477_n2682, DP_OP_422J2_124_3477_n2681,
         DP_OP_422J2_124_3477_n2680, DP_OP_422J2_124_3477_n2679,
         DP_OP_422J2_124_3477_n2678, DP_OP_422J2_124_3477_n2677,
         DP_OP_422J2_124_3477_n2676, DP_OP_422J2_124_3477_n2675,
         DP_OP_422J2_124_3477_n2674, DP_OP_422J2_124_3477_n2673,
         DP_OP_422J2_124_3477_n2670, DP_OP_422J2_124_3477_n2669,
         DP_OP_422J2_124_3477_n2667, DP_OP_422J2_124_3477_n2665,
         DP_OP_422J2_124_3477_n2664, DP_OP_422J2_124_3477_n2663,
         DP_OP_422J2_124_3477_n2662, DP_OP_422J2_124_3477_n2661,
         DP_OP_422J2_124_3477_n2660, DP_OP_422J2_124_3477_n2659,
         DP_OP_422J2_124_3477_n2658, DP_OP_422J2_124_3477_n2657,
         DP_OP_422J2_124_3477_n2656, DP_OP_422J2_124_3477_n2655,
         DP_OP_422J2_124_3477_n2654, DP_OP_422J2_124_3477_n2653,
         DP_OP_422J2_124_3477_n2652, DP_OP_422J2_124_3477_n2651,
         DP_OP_422J2_124_3477_n2650, DP_OP_422J2_124_3477_n2649,
         DP_OP_422J2_124_3477_n2648, DP_OP_422J2_124_3477_n2647,
         DP_OP_422J2_124_3477_n2646, DP_OP_422J2_124_3477_n2645,
         DP_OP_422J2_124_3477_n2644, DP_OP_422J2_124_3477_n2643,
         DP_OP_422J2_124_3477_n2642, DP_OP_422J2_124_3477_n2641,
         DP_OP_422J2_124_3477_n2640, DP_OP_422J2_124_3477_n2639,
         DP_OP_422J2_124_3477_n2638, DP_OP_422J2_124_3477_n2637,
         DP_OP_422J2_124_3477_n2636, DP_OP_422J2_124_3477_n2635,
         DP_OP_422J2_124_3477_n2634, DP_OP_422J2_124_3477_n2633,
         DP_OP_422J2_124_3477_n2632, DP_OP_422J2_124_3477_n2631,
         DP_OP_422J2_124_3477_n2630, DP_OP_422J2_124_3477_n2629,
         DP_OP_422J2_124_3477_n2627, DP_OP_422J2_124_3477_n2626,
         DP_OP_422J2_124_3477_n2625, DP_OP_422J2_124_3477_n2622,
         DP_OP_422J2_124_3477_n2621, DP_OP_422J2_124_3477_n2620,
         DP_OP_422J2_124_3477_n2619, DP_OP_422J2_124_3477_n2618,
         DP_OP_422J2_124_3477_n2617, DP_OP_422J2_124_3477_n2616,
         DP_OP_422J2_124_3477_n2615, DP_OP_422J2_124_3477_n2614,
         DP_OP_422J2_124_3477_n2613, DP_OP_422J2_124_3477_n2612,
         DP_OP_422J2_124_3477_n2611, DP_OP_422J2_124_3477_n2610,
         DP_OP_422J2_124_3477_n2609, DP_OP_422J2_124_3477_n2608,
         DP_OP_422J2_124_3477_n2607, DP_OP_422J2_124_3477_n2606,
         DP_OP_422J2_124_3477_n2605, DP_OP_422J2_124_3477_n2604,
         DP_OP_422J2_124_3477_n2603, DP_OP_422J2_124_3477_n2602,
         DP_OP_422J2_124_3477_n2601, DP_OP_422J2_124_3477_n2600,
         DP_OP_422J2_124_3477_n2599, DP_OP_422J2_124_3477_n2598,
         DP_OP_422J2_124_3477_n2597, DP_OP_422J2_124_3477_n2596,
         DP_OP_422J2_124_3477_n2595, DP_OP_422J2_124_3477_n2594,
         DP_OP_422J2_124_3477_n2593, DP_OP_422J2_124_3477_n2592,
         DP_OP_422J2_124_3477_n2591, DP_OP_422J2_124_3477_n2590,
         DP_OP_422J2_124_3477_n2589, DP_OP_422J2_124_3477_n2588,
         DP_OP_422J2_124_3477_n2587, DP_OP_422J2_124_3477_n2586,
         DP_OP_422J2_124_3477_n2585, DP_OP_422J2_124_3477_n2583,
         DP_OP_422J2_124_3477_n2582, DP_OP_422J2_124_3477_n2580,
         DP_OP_422J2_124_3477_n2579, DP_OP_422J2_124_3477_n2578,
         DP_OP_422J2_124_3477_n2577, DP_OP_422J2_124_3477_n2576,
         DP_OP_422J2_124_3477_n2575, DP_OP_422J2_124_3477_n2574,
         DP_OP_422J2_124_3477_n2573, DP_OP_422J2_124_3477_n2572,
         DP_OP_422J2_124_3477_n2571, DP_OP_422J2_124_3477_n2569,
         DP_OP_422J2_124_3477_n2568, DP_OP_422J2_124_3477_n2567,
         DP_OP_422J2_124_3477_n2566, DP_OP_422J2_124_3477_n2565,
         DP_OP_422J2_124_3477_n2564, DP_OP_422J2_124_3477_n2563,
         DP_OP_422J2_124_3477_n2562, DP_OP_422J2_124_3477_n2561,
         DP_OP_422J2_124_3477_n2560, DP_OP_422J2_124_3477_n2559,
         DP_OP_422J2_124_3477_n2558, DP_OP_422J2_124_3477_n2557,
         DP_OP_422J2_124_3477_n2556, DP_OP_422J2_124_3477_n2555,
         DP_OP_422J2_124_3477_n2554, DP_OP_422J2_124_3477_n2553,
         DP_OP_422J2_124_3477_n2552, DP_OP_422J2_124_3477_n2551,
         DP_OP_422J2_124_3477_n2550, DP_OP_422J2_124_3477_n2549,
         DP_OP_422J2_124_3477_n2548, DP_OP_422J2_124_3477_n2547,
         DP_OP_422J2_124_3477_n2546, DP_OP_422J2_124_3477_n2545,
         DP_OP_422J2_124_3477_n2544, DP_OP_422J2_124_3477_n2543,
         DP_OP_422J2_124_3477_n2542, DP_OP_422J2_124_3477_n2541,
         DP_OP_422J2_124_3477_n2537, DP_OP_422J2_124_3477_n2536,
         DP_OP_422J2_124_3477_n2535, DP_OP_422J2_124_3477_n2534,
         DP_OP_422J2_124_3477_n2533, DP_OP_422J2_124_3477_n2532,
         DP_OP_422J2_124_3477_n2531, DP_OP_422J2_124_3477_n2530,
         DP_OP_422J2_124_3477_n2529, DP_OP_422J2_124_3477_n2528,
         DP_OP_422J2_124_3477_n2527, DP_OP_422J2_124_3477_n2526,
         DP_OP_422J2_124_3477_n2525, DP_OP_422J2_124_3477_n2524,
         DP_OP_422J2_124_3477_n2523, DP_OP_422J2_124_3477_n2522,
         DP_OP_422J2_124_3477_n2521, DP_OP_422J2_124_3477_n2520,
         DP_OP_422J2_124_3477_n2519, DP_OP_422J2_124_3477_n2518,
         DP_OP_422J2_124_3477_n2517, DP_OP_422J2_124_3477_n2516,
         DP_OP_422J2_124_3477_n2515, DP_OP_422J2_124_3477_n2514,
         DP_OP_422J2_124_3477_n2513, DP_OP_422J2_124_3477_n2512,
         DP_OP_422J2_124_3477_n2511, DP_OP_422J2_124_3477_n2510,
         DP_OP_422J2_124_3477_n2509, DP_OP_422J2_124_3477_n2508,
         DP_OP_422J2_124_3477_n2507, DP_OP_422J2_124_3477_n2506,
         DP_OP_422J2_124_3477_n2505, DP_OP_422J2_124_3477_n2504,
         DP_OP_422J2_124_3477_n2503, DP_OP_422J2_124_3477_n2502,
         DP_OP_422J2_124_3477_n2501, DP_OP_422J2_124_3477_n2500,
         DP_OP_422J2_124_3477_n2499, DP_OP_422J2_124_3477_n2498,
         DP_OP_422J2_124_3477_n2497, DP_OP_422J2_124_3477_n2495,
         DP_OP_422J2_124_3477_n2491, DP_OP_422J2_124_3477_n2490,
         DP_OP_422J2_124_3477_n2489, DP_OP_422J2_124_3477_n2488,
         DP_OP_422J2_124_3477_n2486, DP_OP_422J2_124_3477_n2485,
         DP_OP_422J2_124_3477_n2484, DP_OP_422J2_124_3477_n2483,
         DP_OP_422J2_124_3477_n2482, DP_OP_422J2_124_3477_n2481,
         DP_OP_422J2_124_3477_n2480, DP_OP_422J2_124_3477_n2479,
         DP_OP_422J2_124_3477_n2478, DP_OP_422J2_124_3477_n2477,
         DP_OP_422J2_124_3477_n2476, DP_OP_422J2_124_3477_n2475,
         DP_OP_422J2_124_3477_n2474, DP_OP_422J2_124_3477_n2473,
         DP_OP_422J2_124_3477_n2472, DP_OP_422J2_124_3477_n2471,
         DP_OP_422J2_124_3477_n2470, DP_OP_422J2_124_3477_n2469,
         DP_OP_422J2_124_3477_n2468, DP_OP_422J2_124_3477_n2467,
         DP_OP_422J2_124_3477_n2466, DP_OP_422J2_124_3477_n2465,
         DP_OP_422J2_124_3477_n2464, DP_OP_422J2_124_3477_n2463,
         DP_OP_422J2_124_3477_n2462, DP_OP_422J2_124_3477_n2461,
         DP_OP_422J2_124_3477_n2460, DP_OP_422J2_124_3477_n2459,
         DP_OP_422J2_124_3477_n2458, DP_OP_422J2_124_3477_n2457,
         DP_OP_422J2_124_3477_n2456, DP_OP_422J2_124_3477_n2455,
         DP_OP_422J2_124_3477_n2454, DP_OP_422J2_124_3477_n2450,
         DP_OP_422J2_124_3477_n2448, DP_OP_422J2_124_3477_n2446,
         DP_OP_422J2_124_3477_n2445, DP_OP_422J2_124_3477_n2444,
         DP_OP_422J2_124_3477_n2443, DP_OP_422J2_124_3477_n2442,
         DP_OP_422J2_124_3477_n2441, DP_OP_422J2_124_3477_n2440,
         DP_OP_422J2_124_3477_n2439, DP_OP_422J2_124_3477_n2438,
         DP_OP_422J2_124_3477_n2437, DP_OP_422J2_124_3477_n2436,
         DP_OP_422J2_124_3477_n2435, DP_OP_422J2_124_3477_n2434,
         DP_OP_422J2_124_3477_n2433, DP_OP_422J2_124_3477_n2432,
         DP_OP_422J2_124_3477_n2431, DP_OP_422J2_124_3477_n2430,
         DP_OP_422J2_124_3477_n2429, DP_OP_422J2_124_3477_n2428,
         DP_OP_422J2_124_3477_n2427, DP_OP_422J2_124_3477_n2426,
         DP_OP_422J2_124_3477_n2425, DP_OP_422J2_124_3477_n2424,
         DP_OP_422J2_124_3477_n2423, DP_OP_422J2_124_3477_n2422,
         DP_OP_422J2_124_3477_n2421, DP_OP_422J2_124_3477_n2420,
         DP_OP_422J2_124_3477_n2419, DP_OP_422J2_124_3477_n2418,
         DP_OP_422J2_124_3477_n2417, DP_OP_422J2_124_3477_n2416,
         DP_OP_422J2_124_3477_n2415, DP_OP_422J2_124_3477_n2414,
         DP_OP_422J2_124_3477_n2413, DP_OP_422J2_124_3477_n2412,
         DP_OP_422J2_124_3477_n2411, DP_OP_422J2_124_3477_n2410,
         DP_OP_422J2_124_3477_n2409, DP_OP_422J2_124_3477_n2407,
         DP_OP_422J2_124_3477_n2406, DP_OP_422J2_124_3477_n2405,
         DP_OP_422J2_124_3477_n2404, DP_OP_422J2_124_3477_n2401,
         DP_OP_422J2_124_3477_n2399, DP_OP_422J2_124_3477_n2398,
         DP_OP_422J2_124_3477_n2397, DP_OP_422J2_124_3477_n2396,
         DP_OP_422J2_124_3477_n2395, DP_OP_422J2_124_3477_n2394,
         DP_OP_422J2_124_3477_n2393, DP_OP_422J2_124_3477_n2392,
         DP_OP_422J2_124_3477_n2391, DP_OP_422J2_124_3477_n2390,
         DP_OP_422J2_124_3477_n2389, DP_OP_422J2_124_3477_n2388,
         DP_OP_422J2_124_3477_n2387, DP_OP_422J2_124_3477_n2386,
         DP_OP_422J2_124_3477_n2385, DP_OP_422J2_124_3477_n2384,
         DP_OP_422J2_124_3477_n2383, DP_OP_422J2_124_3477_n2382,
         DP_OP_422J2_124_3477_n2381, DP_OP_422J2_124_3477_n2380,
         DP_OP_422J2_124_3477_n2379, DP_OP_422J2_124_3477_n2378,
         DP_OP_422J2_124_3477_n2377, DP_OP_422J2_124_3477_n2376,
         DP_OP_422J2_124_3477_n2375, DP_OP_422J2_124_3477_n2374,
         DP_OP_422J2_124_3477_n2373, DP_OP_422J2_124_3477_n2372,
         DP_OP_422J2_124_3477_n2371, DP_OP_422J2_124_3477_n2370,
         DP_OP_422J2_124_3477_n2369, DP_OP_422J2_124_3477_n2368,
         DP_OP_422J2_124_3477_n2367, DP_OP_422J2_124_3477_n2366,
         DP_OP_422J2_124_3477_n2362, DP_OP_422J2_124_3477_n2358,
         DP_OP_422J2_124_3477_n2357, DP_OP_422J2_124_3477_n2356,
         DP_OP_422J2_124_3477_n2355, DP_OP_422J2_124_3477_n2354,
         DP_OP_422J2_124_3477_n2353, DP_OP_422J2_124_3477_n2352,
         DP_OP_422J2_124_3477_n2351, DP_OP_422J2_124_3477_n2350,
         DP_OP_422J2_124_3477_n2349, DP_OP_422J2_124_3477_n2348,
         DP_OP_422J2_124_3477_n2347, DP_OP_422J2_124_3477_n2346,
         DP_OP_422J2_124_3477_n2345, DP_OP_422J2_124_3477_n2344,
         DP_OP_422J2_124_3477_n2343, DP_OP_422J2_124_3477_n2342,
         DP_OP_422J2_124_3477_n2341, DP_OP_422J2_124_3477_n2340,
         DP_OP_422J2_124_3477_n2339, DP_OP_422J2_124_3477_n2338,
         DP_OP_422J2_124_3477_n2337, DP_OP_422J2_124_3477_n2336,
         DP_OP_422J2_124_3477_n2335, DP_OP_422J2_124_3477_n2334,
         DP_OP_422J2_124_3477_n2333, DP_OP_422J2_124_3477_n2332,
         DP_OP_422J2_124_3477_n2331, DP_OP_422J2_124_3477_n2330,
         DP_OP_422J2_124_3477_n2329, DP_OP_422J2_124_3477_n2328,
         DP_OP_422J2_124_3477_n2327, DP_OP_422J2_124_3477_n2326,
         DP_OP_422J2_124_3477_n2325, DP_OP_422J2_124_3477_n2324,
         DP_OP_422J2_124_3477_n2323, DP_OP_422J2_124_3477_n2322,
         DP_OP_422J2_124_3477_n2321, DP_OP_422J2_124_3477_n2320,
         DP_OP_422J2_124_3477_n2318, DP_OP_422J2_124_3477_n2314,
         DP_OP_422J2_124_3477_n2313, DP_OP_422J2_124_3477_n2312,
         DP_OP_422J2_124_3477_n2311, DP_OP_422J2_124_3477_n2310,
         DP_OP_422J2_124_3477_n2309, DP_OP_422J2_124_3477_n2308,
         DP_OP_422J2_124_3477_n2307, DP_OP_422J2_124_3477_n2306,
         DP_OP_422J2_124_3477_n2305, DP_OP_422J2_124_3477_n2304,
         DP_OP_422J2_124_3477_n2303, DP_OP_422J2_124_3477_n2302,
         DP_OP_422J2_124_3477_n2301, DP_OP_422J2_124_3477_n2300,
         DP_OP_422J2_124_3477_n2299, DP_OP_422J2_124_3477_n2298,
         DP_OP_422J2_124_3477_n2297, DP_OP_422J2_124_3477_n2296,
         DP_OP_422J2_124_3477_n2295, DP_OP_422J2_124_3477_n2294,
         DP_OP_422J2_124_3477_n2293, DP_OP_422J2_124_3477_n2292,
         DP_OP_422J2_124_3477_n2291, DP_OP_422J2_124_3477_n2290,
         DP_OP_422J2_124_3477_n2289, DP_OP_422J2_124_3477_n2288,
         DP_OP_422J2_124_3477_n2287, DP_OP_422J2_124_3477_n2286,
         DP_OP_422J2_124_3477_n2285, DP_OP_422J2_124_3477_n2284,
         DP_OP_422J2_124_3477_n2283, DP_OP_422J2_124_3477_n2282,
         DP_OP_422J2_124_3477_n2281, DP_OP_422J2_124_3477_n2280,
         DP_OP_422J2_124_3477_n2279, DP_OP_422J2_124_3477_n2278,
         DP_OP_422J2_124_3477_n2277, DP_OP_422J2_124_3477_n2276,
         DP_OP_422J2_124_3477_n2275, DP_OP_422J2_124_3477_n2270,
         DP_OP_422J2_124_3477_n2269, DP_OP_422J2_124_3477_n2268,
         DP_OP_422J2_124_3477_n2267, DP_OP_422J2_124_3477_n2266,
         DP_OP_422J2_124_3477_n2265, DP_OP_422J2_124_3477_n2264,
         DP_OP_422J2_124_3477_n2263, DP_OP_422J2_124_3477_n2262,
         DP_OP_422J2_124_3477_n2261, DP_OP_422J2_124_3477_n2260,
         DP_OP_422J2_124_3477_n2259, DP_OP_422J2_124_3477_n2258,
         DP_OP_422J2_124_3477_n2257, DP_OP_422J2_124_3477_n2256,
         DP_OP_422J2_124_3477_n2255, DP_OP_422J2_124_3477_n2254,
         DP_OP_422J2_124_3477_n2253, DP_OP_422J2_124_3477_n2252,
         DP_OP_422J2_124_3477_n2251, DP_OP_422J2_124_3477_n2250,
         DP_OP_422J2_124_3477_n2249, DP_OP_422J2_124_3477_n2248,
         DP_OP_422J2_124_3477_n2247, DP_OP_422J2_124_3477_n2246,
         DP_OP_422J2_124_3477_n2245, DP_OP_422J2_124_3477_n2244,
         DP_OP_422J2_124_3477_n2243, DP_OP_422J2_124_3477_n2242,
         DP_OP_422J2_124_3477_n2241, DP_OP_422J2_124_3477_n2240,
         DP_OP_422J2_124_3477_n2239, DP_OP_422J2_124_3477_n2238,
         DP_OP_422J2_124_3477_n2237, DP_OP_422J2_124_3477_n2236,
         DP_OP_422J2_124_3477_n2235, DP_OP_422J2_124_3477_n2234,
         DP_OP_422J2_124_3477_n2231, DP_OP_422J2_124_3477_n2230,
         DP_OP_422J2_124_3477_n2225, DP_OP_422J2_124_3477_n2224,
         DP_OP_422J2_124_3477_n2223, DP_OP_422J2_124_3477_n2222,
         DP_OP_422J2_124_3477_n2221, DP_OP_422J2_124_3477_n2220,
         DP_OP_422J2_124_3477_n2219, DP_OP_422J2_124_3477_n2218,
         DP_OP_422J2_124_3477_n2217, DP_OP_422J2_124_3477_n2216,
         DP_OP_422J2_124_3477_n2215, DP_OP_422J2_124_3477_n2214,
         DP_OP_422J2_124_3477_n2213, DP_OP_422J2_124_3477_n2212,
         DP_OP_422J2_124_3477_n2211, DP_OP_422J2_124_3477_n2210,
         DP_OP_422J2_124_3477_n2209, DP_OP_422J2_124_3477_n2208,
         DP_OP_422J2_124_3477_n2207, DP_OP_422J2_124_3477_n2206,
         DP_OP_422J2_124_3477_n2205, DP_OP_422J2_124_3477_n2204,
         DP_OP_422J2_124_3477_n2203, DP_OP_422J2_124_3477_n2202,
         DP_OP_422J2_124_3477_n2201, DP_OP_422J2_124_3477_n2200,
         DP_OP_422J2_124_3477_n2199, DP_OP_422J2_124_3477_n2198,
         DP_OP_422J2_124_3477_n2197, DP_OP_422J2_124_3477_n2196,
         DP_OP_422J2_124_3477_n2195, DP_OP_422J2_124_3477_n2194,
         DP_OP_422J2_124_3477_n2193, DP_OP_422J2_124_3477_n2192,
         DP_OP_422J2_124_3477_n2191, DP_OP_422J2_124_3477_n2190,
         DP_OP_422J2_124_3477_n2189, DP_OP_422J2_124_3477_n2186,
         DP_OP_422J2_124_3477_n2185, DP_OP_422J2_124_3477_n2183,
         DP_OP_422J2_124_3477_n2181, DP_OP_422J2_124_3477_n2179,
         DP_OP_422J2_124_3477_n2178, DP_OP_422J2_124_3477_n2177,
         DP_OP_422J2_124_3477_n2176, DP_OP_422J2_124_3477_n2175,
         DP_OP_422J2_124_3477_n2174, DP_OP_422J2_124_3477_n2173,
         DP_OP_422J2_124_3477_n2172, DP_OP_422J2_124_3477_n2171,
         DP_OP_422J2_124_3477_n2170, DP_OP_422J2_124_3477_n2169,
         DP_OP_422J2_124_3477_n2168, DP_OP_422J2_124_3477_n2167,
         DP_OP_422J2_124_3477_n2166, DP_OP_422J2_124_3477_n2165,
         DP_OP_422J2_124_3477_n2164, DP_OP_422J2_124_3477_n2163,
         DP_OP_422J2_124_3477_n2162, DP_OP_422J2_124_3477_n2161,
         DP_OP_422J2_124_3477_n2160, DP_OP_422J2_124_3477_n2159,
         DP_OP_422J2_124_3477_n2158, DP_OP_422J2_124_3477_n2157,
         DP_OP_422J2_124_3477_n2156, DP_OP_422J2_124_3477_n2155,
         DP_OP_422J2_124_3477_n2154, DP_OP_422J2_124_3477_n2153,
         DP_OP_422J2_124_3477_n2152, DP_OP_422J2_124_3477_n2151,
         DP_OP_422J2_124_3477_n2150, DP_OP_422J2_124_3477_n2149,
         DP_OP_422J2_124_3477_n2148, DP_OP_422J2_124_3477_n2147,
         DP_OP_422J2_124_3477_n2146, DP_OP_422J2_124_3477_n2144,
         DP_OP_422J2_124_3477_n2143, DP_OP_422J2_124_3477_n2142,
         DP_OP_422J2_124_3477_n2140, DP_OP_422J2_124_3477_n2138,
         DP_OP_422J2_124_3477_n2137, DP_OP_422J2_124_3477_n2135,
         DP_OP_422J2_124_3477_n2134, DP_OP_422J2_124_3477_n2133,
         DP_OP_422J2_124_3477_n2132, DP_OP_422J2_124_3477_n2131,
         DP_OP_422J2_124_3477_n2130, DP_OP_422J2_124_3477_n2129,
         DP_OP_422J2_124_3477_n2128, DP_OP_422J2_124_3477_n2127,
         DP_OP_422J2_124_3477_n2126, DP_OP_422J2_124_3477_n2125,
         DP_OP_422J2_124_3477_n2124, DP_OP_422J2_124_3477_n2123,
         DP_OP_422J2_124_3477_n2122, DP_OP_422J2_124_3477_n2121,
         DP_OP_422J2_124_3477_n2120, DP_OP_422J2_124_3477_n2119,
         DP_OP_422J2_124_3477_n2118, DP_OP_422J2_124_3477_n2117,
         DP_OP_422J2_124_3477_n2116, DP_OP_422J2_124_3477_n2115,
         DP_OP_422J2_124_3477_n2114, DP_OP_422J2_124_3477_n2113,
         DP_OP_422J2_124_3477_n2112, DP_OP_422J2_124_3477_n2111,
         DP_OP_422J2_124_3477_n2110, DP_OP_422J2_124_3477_n2109,
         DP_OP_422J2_124_3477_n2108, DP_OP_422J2_124_3477_n2107,
         DP_OP_422J2_124_3477_n2106, DP_OP_422J2_124_3477_n2105,
         DP_OP_422J2_124_3477_n2104, DP_OP_422J2_124_3477_n2103,
         DP_OP_422J2_124_3477_n2102, DP_OP_422J2_124_3477_n2100,
         DP_OP_422J2_124_3477_n2093, DP_OP_422J2_124_3477_n2092,
         DP_OP_422J2_124_3477_n2091, DP_OP_422J2_124_3477_n2090,
         DP_OP_422J2_124_3477_n2089, DP_OP_422J2_124_3477_n2088,
         DP_OP_422J2_124_3477_n2087, DP_OP_422J2_124_3477_n2086,
         DP_OP_422J2_124_3477_n2085, DP_OP_422J2_124_3477_n2084,
         DP_OP_422J2_124_3477_n2083, DP_OP_422J2_124_3477_n2082,
         DP_OP_422J2_124_3477_n2081, DP_OP_422J2_124_3477_n2080,
         DP_OP_422J2_124_3477_n2079, DP_OP_422J2_124_3477_n2078,
         DP_OP_422J2_124_3477_n2077, DP_OP_422J2_124_3477_n2076,
         DP_OP_422J2_124_3477_n2075, DP_OP_422J2_124_3477_n2074,
         DP_OP_422J2_124_3477_n2073, DP_OP_422J2_124_3477_n2072,
         DP_OP_422J2_124_3477_n2071, DP_OP_422J2_124_3477_n2070,
         DP_OP_422J2_124_3477_n2069, DP_OP_422J2_124_3477_n2068,
         DP_OP_422J2_124_3477_n2067, DP_OP_422J2_124_3477_n2066,
         DP_OP_422J2_124_3477_n2064, DP_OP_422J2_124_3477_n2063,
         DP_OP_422J2_124_3477_n2062, DP_OP_422J2_124_3477_n2061,
         DP_OP_422J2_124_3477_n2060, DP_OP_422J2_124_3477_n2059,
         DP_OP_422J2_124_3477_n2058, DP_OP_422J2_124_3477_n2056,
         DP_OP_422J2_124_3477_n2055, DP_OP_422J2_124_3477_n2051,
         DP_OP_422J2_124_3477_n2049, DP_OP_422J2_124_3477_n2048,
         DP_OP_422J2_124_3477_n2047, DP_OP_422J2_124_3477_n2046,
         DP_OP_422J2_124_3477_n2045, DP_OP_422J2_124_3477_n2044,
         DP_OP_422J2_124_3477_n2043, DP_OP_422J2_124_3477_n2042,
         DP_OP_422J2_124_3477_n2041, DP_OP_422J2_124_3477_n2040,
         DP_OP_422J2_124_3477_n2039, DP_OP_422J2_124_3477_n2038,
         DP_OP_422J2_124_3477_n2037, DP_OP_422J2_124_3477_n2036,
         DP_OP_422J2_124_3477_n2035, DP_OP_422J2_124_3477_n2034,
         DP_OP_422J2_124_3477_n2033, DP_OP_422J2_124_3477_n2032,
         DP_OP_422J2_124_3477_n2031, DP_OP_422J2_124_3477_n2030,
         DP_OP_422J2_124_3477_n2029, DP_OP_422J2_124_3477_n2028,
         DP_OP_422J2_124_3477_n2027, DP_OP_422J2_124_3477_n2026,
         DP_OP_422J2_124_3477_n2025, DP_OP_422J2_124_3477_n2024,
         DP_OP_422J2_124_3477_n2023, DP_OP_422J2_124_3477_n2022,
         DP_OP_422J2_124_3477_n2021, DP_OP_422J2_124_3477_n2020,
         DP_OP_422J2_124_3477_n2019, DP_OP_422J2_124_3477_n2018,
         DP_OP_422J2_124_3477_n2017, DP_OP_422J2_124_3477_n2016,
         DP_OP_422J2_124_3477_n2015, DP_OP_422J2_124_3477_n2014,
         DP_OP_422J2_124_3477_n2013, DP_OP_422J2_124_3477_n2011,
         DP_OP_422J2_124_3477_n2007, DP_OP_422J2_124_3477_n2006,
         DP_OP_422J2_124_3477_n2005, DP_OP_422J2_124_3477_n2004,
         DP_OP_422J2_124_3477_n2003, DP_OP_422J2_124_3477_n2002,
         DP_OP_422J2_124_3477_n2001, DP_OP_422J2_124_3477_n2000,
         DP_OP_422J2_124_3477_n1999, DP_OP_422J2_124_3477_n1998,
         DP_OP_422J2_124_3477_n1997, DP_OP_422J2_124_3477_n1996,
         DP_OP_422J2_124_3477_n1995, DP_OP_422J2_124_3477_n1994,
         DP_OP_422J2_124_3477_n1993, DP_OP_422J2_124_3477_n1992,
         DP_OP_422J2_124_3477_n1991, DP_OP_422J2_124_3477_n1990,
         DP_OP_422J2_124_3477_n1989, DP_OP_422J2_124_3477_n1988,
         DP_OP_422J2_124_3477_n1987, DP_OP_422J2_124_3477_n1986,
         DP_OP_422J2_124_3477_n1985, DP_OP_422J2_124_3477_n1984,
         DP_OP_422J2_124_3477_n1983, DP_OP_422J2_124_3477_n1982,
         DP_OP_422J2_124_3477_n1981, DP_OP_422J2_124_3477_n1980,
         DP_OP_422J2_124_3477_n1979, DP_OP_422J2_124_3477_n1978,
         DP_OP_422J2_124_3477_n1977, DP_OP_422J2_124_3477_n1976,
         DP_OP_422J2_124_3477_n1975, DP_OP_422J2_124_3477_n1974,
         DP_OP_422J2_124_3477_n1973, DP_OP_422J2_124_3477_n1972,
         DP_OP_422J2_124_3477_n1971, DP_OP_422J2_124_3477_n1970,
         DP_OP_422J2_124_3477_n1936, DP_OP_422J2_124_3477_n1935,
         DP_OP_422J2_124_3477_n1934, DP_OP_422J2_124_3477_n1933,
         DP_OP_422J2_124_3477_n1932, DP_OP_422J2_124_3477_n1931,
         DP_OP_422J2_124_3477_n1930, DP_OP_422J2_124_3477_n1929,
         DP_OP_422J2_124_3477_n1928, DP_OP_422J2_124_3477_n1927,
         DP_OP_422J2_124_3477_n1926, DP_OP_422J2_124_3477_n1925,
         DP_OP_422J2_124_3477_n1924, DP_OP_422J2_124_3477_n1923,
         DP_OP_422J2_124_3477_n1921, DP_OP_422J2_124_3477_n1920,
         DP_OP_422J2_124_3477_n1919, DP_OP_422J2_124_3477_n1918,
         DP_OP_422J2_124_3477_n1917, DP_OP_422J2_124_3477_n1916,
         DP_OP_422J2_124_3477_n1915, DP_OP_422J2_124_3477_n1914,
         DP_OP_422J2_124_3477_n1913, DP_OP_422J2_124_3477_n1912,
         DP_OP_422J2_124_3477_n1911, DP_OP_422J2_124_3477_n1910,
         DP_OP_422J2_124_3477_n1909, DP_OP_422J2_124_3477_n1908,
         DP_OP_422J2_124_3477_n1907, DP_OP_422J2_124_3477_n1906,
         DP_OP_422J2_124_3477_n1905, DP_OP_422J2_124_3477_n1904,
         DP_OP_422J2_124_3477_n1903, DP_OP_422J2_124_3477_n1902,
         DP_OP_422J2_124_3477_n1901, DP_OP_422J2_124_3477_n1900,
         DP_OP_422J2_124_3477_n1899, DP_OP_422J2_124_3477_n1898,
         DP_OP_422J2_124_3477_n1897, DP_OP_422J2_124_3477_n1896,
         DP_OP_422J2_124_3477_n1895, DP_OP_422J2_124_3477_n1894,
         DP_OP_422J2_124_3477_n1893, DP_OP_422J2_124_3477_n1892,
         DP_OP_422J2_124_3477_n1891, DP_OP_422J2_124_3477_n1890,
         DP_OP_422J2_124_3477_n1889, DP_OP_422J2_124_3477_n1888,
         DP_OP_422J2_124_3477_n1887, DP_OP_422J2_124_3477_n1886,
         DP_OP_422J2_124_3477_n1885, DP_OP_422J2_124_3477_n1884,
         DP_OP_422J2_124_3477_n1883, DP_OP_422J2_124_3477_n1882,
         DP_OP_422J2_124_3477_n1881, DP_OP_422J2_124_3477_n1880,
         DP_OP_422J2_124_3477_n1879, DP_OP_422J2_124_3477_n1878,
         DP_OP_422J2_124_3477_n1877, DP_OP_422J2_124_3477_n1876,
         DP_OP_422J2_124_3477_n1875, DP_OP_422J2_124_3477_n1874,
         DP_OP_422J2_124_3477_n1873, DP_OP_422J2_124_3477_n1872,
         DP_OP_422J2_124_3477_n1871, DP_OP_422J2_124_3477_n1870,
         DP_OP_422J2_124_3477_n1869, DP_OP_422J2_124_3477_n1868,
         DP_OP_422J2_124_3477_n1867, DP_OP_422J2_124_3477_n1866,
         DP_OP_422J2_124_3477_n1865, DP_OP_422J2_124_3477_n1864,
         DP_OP_422J2_124_3477_n1863, DP_OP_422J2_124_3477_n1862,
         DP_OP_422J2_124_3477_n1861, DP_OP_422J2_124_3477_n1860,
         DP_OP_422J2_124_3477_n1859, DP_OP_422J2_124_3477_n1858,
         DP_OP_422J2_124_3477_n1857, DP_OP_422J2_124_3477_n1856,
         DP_OP_422J2_124_3477_n1855, DP_OP_422J2_124_3477_n1854,
         DP_OP_422J2_124_3477_n1853, DP_OP_422J2_124_3477_n1852,
         DP_OP_422J2_124_3477_n1851, DP_OP_422J2_124_3477_n1850,
         DP_OP_422J2_124_3477_n1849, DP_OP_422J2_124_3477_n1848,
         DP_OP_422J2_124_3477_n1847, DP_OP_422J2_124_3477_n1846,
         DP_OP_422J2_124_3477_n1845, DP_OP_422J2_124_3477_n1844,
         DP_OP_422J2_124_3477_n1843, DP_OP_422J2_124_3477_n1842,
         DP_OP_422J2_124_3477_n1841, DP_OP_422J2_124_3477_n1840,
         DP_OP_422J2_124_3477_n1839, DP_OP_422J2_124_3477_n1838,
         DP_OP_422J2_124_3477_n1837, DP_OP_422J2_124_3477_n1836,
         DP_OP_422J2_124_3477_n1835, DP_OP_422J2_124_3477_n1834,
         DP_OP_422J2_124_3477_n1833, DP_OP_422J2_124_3477_n1832,
         DP_OP_422J2_124_3477_n1831, DP_OP_422J2_124_3477_n1830,
         DP_OP_422J2_124_3477_n1829, DP_OP_422J2_124_3477_n1828,
         DP_OP_422J2_124_3477_n1827, DP_OP_422J2_124_3477_n1826,
         DP_OP_422J2_124_3477_n1825, DP_OP_422J2_124_3477_n1824,
         DP_OP_422J2_124_3477_n1823, DP_OP_422J2_124_3477_n1822,
         DP_OP_422J2_124_3477_n1821, DP_OP_422J2_124_3477_n1820,
         DP_OP_422J2_124_3477_n1819, DP_OP_422J2_124_3477_n1818,
         DP_OP_422J2_124_3477_n1817, DP_OP_422J2_124_3477_n1816,
         DP_OP_422J2_124_3477_n1815, DP_OP_422J2_124_3477_n1814,
         DP_OP_422J2_124_3477_n1813, DP_OP_422J2_124_3477_n1812,
         DP_OP_422J2_124_3477_n1811, DP_OP_422J2_124_3477_n1810,
         DP_OP_422J2_124_3477_n1809, DP_OP_422J2_124_3477_n1808,
         DP_OP_422J2_124_3477_n1807, DP_OP_422J2_124_3477_n1806,
         DP_OP_422J2_124_3477_n1805, DP_OP_422J2_124_3477_n1804,
         DP_OP_422J2_124_3477_n1803, DP_OP_422J2_124_3477_n1802,
         DP_OP_422J2_124_3477_n1801, DP_OP_422J2_124_3477_n1800,
         DP_OP_422J2_124_3477_n1799, DP_OP_422J2_124_3477_n1798,
         DP_OP_422J2_124_3477_n1797, DP_OP_422J2_124_3477_n1796,
         DP_OP_422J2_124_3477_n1795, DP_OP_422J2_124_3477_n1794,
         DP_OP_422J2_124_3477_n1793, DP_OP_422J2_124_3477_n1792,
         DP_OP_422J2_124_3477_n1791, DP_OP_422J2_124_3477_n1790,
         DP_OP_422J2_124_3477_n1789, DP_OP_422J2_124_3477_n1788,
         DP_OP_422J2_124_3477_n1787, DP_OP_422J2_124_3477_n1786,
         DP_OP_422J2_124_3477_n1785, DP_OP_422J2_124_3477_n1784,
         DP_OP_422J2_124_3477_n1783, DP_OP_422J2_124_3477_n1782,
         DP_OP_422J2_124_3477_n1781, DP_OP_422J2_124_3477_n1780,
         DP_OP_422J2_124_3477_n1779, DP_OP_422J2_124_3477_n1778,
         DP_OP_422J2_124_3477_n1777, DP_OP_422J2_124_3477_n1776,
         DP_OP_422J2_124_3477_n1775, DP_OP_422J2_124_3477_n1774,
         DP_OP_422J2_124_3477_n1773, DP_OP_422J2_124_3477_n1772,
         DP_OP_422J2_124_3477_n1771, DP_OP_422J2_124_3477_n1770,
         DP_OP_422J2_124_3477_n1769, DP_OP_422J2_124_3477_n1768,
         DP_OP_422J2_124_3477_n1767, DP_OP_422J2_124_3477_n1766,
         DP_OP_422J2_124_3477_n1765, DP_OP_422J2_124_3477_n1764,
         DP_OP_422J2_124_3477_n1763, DP_OP_422J2_124_3477_n1762,
         DP_OP_422J2_124_3477_n1761, DP_OP_422J2_124_3477_n1760,
         DP_OP_422J2_124_3477_n1759, DP_OP_422J2_124_3477_n1758,
         DP_OP_422J2_124_3477_n1757, DP_OP_422J2_124_3477_n1756,
         DP_OP_422J2_124_3477_n1755, DP_OP_422J2_124_3477_n1754,
         DP_OP_422J2_124_3477_n1753, DP_OP_422J2_124_3477_n1752,
         DP_OP_422J2_124_3477_n1751, DP_OP_422J2_124_3477_n1750,
         DP_OP_422J2_124_3477_n1749, DP_OP_422J2_124_3477_n1748,
         DP_OP_422J2_124_3477_n1747, DP_OP_422J2_124_3477_n1746,
         DP_OP_422J2_124_3477_n1745, DP_OP_422J2_124_3477_n1744,
         DP_OP_422J2_124_3477_n1743, DP_OP_422J2_124_3477_n1742,
         DP_OP_422J2_124_3477_n1741, DP_OP_422J2_124_3477_n1740,
         DP_OP_422J2_124_3477_n1739, DP_OP_422J2_124_3477_n1738,
         DP_OP_422J2_124_3477_n1737, DP_OP_422J2_124_3477_n1736,
         DP_OP_422J2_124_3477_n1735, DP_OP_422J2_124_3477_n1734,
         DP_OP_422J2_124_3477_n1733, DP_OP_422J2_124_3477_n1732,
         DP_OP_422J2_124_3477_n1731, DP_OP_422J2_124_3477_n1730,
         DP_OP_422J2_124_3477_n1729, DP_OP_422J2_124_3477_n1728,
         DP_OP_422J2_124_3477_n1727, DP_OP_422J2_124_3477_n1726,
         DP_OP_422J2_124_3477_n1725, DP_OP_422J2_124_3477_n1724,
         DP_OP_422J2_124_3477_n1723, DP_OP_422J2_124_3477_n1722,
         DP_OP_422J2_124_3477_n1721, DP_OP_422J2_124_3477_n1720,
         DP_OP_422J2_124_3477_n1719, DP_OP_422J2_124_3477_n1718,
         DP_OP_422J2_124_3477_n1717, DP_OP_422J2_124_3477_n1716,
         DP_OP_422J2_124_3477_n1715, DP_OP_422J2_124_3477_n1714,
         DP_OP_422J2_124_3477_n1713, DP_OP_422J2_124_3477_n1712,
         DP_OP_422J2_124_3477_n1711, DP_OP_422J2_124_3477_n1710,
         DP_OP_422J2_124_3477_n1709, DP_OP_422J2_124_3477_n1708,
         DP_OP_422J2_124_3477_n1707, DP_OP_422J2_124_3477_n1706,
         DP_OP_422J2_124_3477_n1705, DP_OP_422J2_124_3477_n1704,
         DP_OP_422J2_124_3477_n1703, DP_OP_422J2_124_3477_n1702,
         DP_OP_422J2_124_3477_n1701, DP_OP_422J2_124_3477_n1700,
         DP_OP_422J2_124_3477_n1699, DP_OP_422J2_124_3477_n1698,
         DP_OP_422J2_124_3477_n1697, DP_OP_422J2_124_3477_n1696,
         DP_OP_422J2_124_3477_n1695, DP_OP_422J2_124_3477_n1694,
         DP_OP_422J2_124_3477_n1693, DP_OP_422J2_124_3477_n1692,
         DP_OP_422J2_124_3477_n1691, DP_OP_422J2_124_3477_n1690,
         DP_OP_422J2_124_3477_n1689, DP_OP_422J2_124_3477_n1688,
         DP_OP_422J2_124_3477_n1687, DP_OP_422J2_124_3477_n1686,
         DP_OP_422J2_124_3477_n1685, DP_OP_422J2_124_3477_n1684,
         DP_OP_422J2_124_3477_n1683, DP_OP_422J2_124_3477_n1682,
         DP_OP_422J2_124_3477_n1681, DP_OP_422J2_124_3477_n1680,
         DP_OP_422J2_124_3477_n1679, DP_OP_422J2_124_3477_n1678,
         DP_OP_422J2_124_3477_n1677, DP_OP_422J2_124_3477_n1676,
         DP_OP_422J2_124_3477_n1675, DP_OP_422J2_124_3477_n1674,
         DP_OP_422J2_124_3477_n1673, DP_OP_422J2_124_3477_n1672,
         DP_OP_422J2_124_3477_n1671, DP_OP_422J2_124_3477_n1670,
         DP_OP_422J2_124_3477_n1669, DP_OP_422J2_124_3477_n1668,
         DP_OP_422J2_124_3477_n1667, DP_OP_422J2_124_3477_n1666,
         DP_OP_422J2_124_3477_n1665, DP_OP_422J2_124_3477_n1664,
         DP_OP_422J2_124_3477_n1663, DP_OP_422J2_124_3477_n1662,
         DP_OP_422J2_124_3477_n1661, DP_OP_422J2_124_3477_n1660,
         DP_OP_422J2_124_3477_n1659, DP_OP_422J2_124_3477_n1658,
         DP_OP_422J2_124_3477_n1657, DP_OP_422J2_124_3477_n1656,
         DP_OP_422J2_124_3477_n1655, DP_OP_422J2_124_3477_n1654,
         DP_OP_422J2_124_3477_n1653, DP_OP_422J2_124_3477_n1652,
         DP_OP_422J2_124_3477_n1651, DP_OP_422J2_124_3477_n1650,
         DP_OP_422J2_124_3477_n1649, DP_OP_422J2_124_3477_n1648,
         DP_OP_422J2_124_3477_n1647, DP_OP_422J2_124_3477_n1646,
         DP_OP_422J2_124_3477_n1645, DP_OP_422J2_124_3477_n1644,
         DP_OP_422J2_124_3477_n1643, DP_OP_422J2_124_3477_n1642,
         DP_OP_422J2_124_3477_n1641, DP_OP_422J2_124_3477_n1640,
         DP_OP_422J2_124_3477_n1639, DP_OP_422J2_124_3477_n1638,
         DP_OP_422J2_124_3477_n1637, DP_OP_422J2_124_3477_n1636,
         DP_OP_422J2_124_3477_n1635, DP_OP_422J2_124_3477_n1634,
         DP_OP_422J2_124_3477_n1633, DP_OP_422J2_124_3477_n1632,
         DP_OP_422J2_124_3477_n1631, DP_OP_422J2_124_3477_n1630,
         DP_OP_422J2_124_3477_n1629, DP_OP_422J2_124_3477_n1628,
         DP_OP_422J2_124_3477_n1627, DP_OP_422J2_124_3477_n1626,
         DP_OP_422J2_124_3477_n1625, DP_OP_422J2_124_3477_n1624,
         DP_OP_422J2_124_3477_n1623, DP_OP_422J2_124_3477_n1622,
         DP_OP_422J2_124_3477_n1621, DP_OP_422J2_124_3477_n1620,
         DP_OP_422J2_124_3477_n1619, DP_OP_422J2_124_3477_n1618,
         DP_OP_422J2_124_3477_n1617, DP_OP_422J2_124_3477_n1616,
         DP_OP_422J2_124_3477_n1615, DP_OP_422J2_124_3477_n1614,
         DP_OP_422J2_124_3477_n1613, DP_OP_422J2_124_3477_n1612,
         DP_OP_422J2_124_3477_n1611, DP_OP_422J2_124_3477_n1610,
         DP_OP_422J2_124_3477_n1609, DP_OP_422J2_124_3477_n1608,
         DP_OP_422J2_124_3477_n1607, DP_OP_422J2_124_3477_n1606,
         DP_OP_422J2_124_3477_n1605, DP_OP_422J2_124_3477_n1604,
         DP_OP_422J2_124_3477_n1603, DP_OP_422J2_124_3477_n1602,
         DP_OP_422J2_124_3477_n1601, DP_OP_422J2_124_3477_n1600,
         DP_OP_422J2_124_3477_n1599, DP_OP_422J2_124_3477_n1598,
         DP_OP_422J2_124_3477_n1597, DP_OP_422J2_124_3477_n1596,
         DP_OP_422J2_124_3477_n1595, DP_OP_422J2_124_3477_n1594,
         DP_OP_422J2_124_3477_n1593, DP_OP_422J2_124_3477_n1592,
         DP_OP_422J2_124_3477_n1591, DP_OP_422J2_124_3477_n1590,
         DP_OP_422J2_124_3477_n1589, DP_OP_422J2_124_3477_n1588,
         DP_OP_422J2_124_3477_n1587, DP_OP_422J2_124_3477_n1586,
         DP_OP_422J2_124_3477_n1585, DP_OP_422J2_124_3477_n1584,
         DP_OP_422J2_124_3477_n1583, DP_OP_422J2_124_3477_n1582,
         DP_OP_422J2_124_3477_n1581, DP_OP_422J2_124_3477_n1580,
         DP_OP_422J2_124_3477_n1579, DP_OP_422J2_124_3477_n1578,
         DP_OP_422J2_124_3477_n1577, DP_OP_422J2_124_3477_n1576,
         DP_OP_422J2_124_3477_n1575, DP_OP_422J2_124_3477_n1574,
         DP_OP_422J2_124_3477_n1573, DP_OP_422J2_124_3477_n1572,
         DP_OP_422J2_124_3477_n1571, DP_OP_422J2_124_3477_n1570,
         DP_OP_422J2_124_3477_n1569, DP_OP_422J2_124_3477_n1568,
         DP_OP_422J2_124_3477_n1567, DP_OP_422J2_124_3477_n1566,
         DP_OP_422J2_124_3477_n1565, DP_OP_422J2_124_3477_n1564,
         DP_OP_422J2_124_3477_n1563, DP_OP_422J2_124_3477_n1562,
         DP_OP_422J2_124_3477_n1561, DP_OP_422J2_124_3477_n1560,
         DP_OP_422J2_124_3477_n1559, DP_OP_422J2_124_3477_n1558,
         DP_OP_422J2_124_3477_n1557, DP_OP_422J2_124_3477_n1556,
         DP_OP_422J2_124_3477_n1555, DP_OP_422J2_124_3477_n1554,
         DP_OP_422J2_124_3477_n1553, DP_OP_422J2_124_3477_n1552,
         DP_OP_422J2_124_3477_n1551, DP_OP_422J2_124_3477_n1550,
         DP_OP_422J2_124_3477_n1549, DP_OP_422J2_124_3477_n1548,
         DP_OP_422J2_124_3477_n1547, DP_OP_422J2_124_3477_n1546,
         DP_OP_422J2_124_3477_n1545, DP_OP_422J2_124_3477_n1544,
         DP_OP_422J2_124_3477_n1543, DP_OP_422J2_124_3477_n1542,
         DP_OP_422J2_124_3477_n1541, DP_OP_422J2_124_3477_n1540,
         DP_OP_422J2_124_3477_n1539, DP_OP_422J2_124_3477_n1538,
         DP_OP_422J2_124_3477_n1537, DP_OP_422J2_124_3477_n1536,
         DP_OP_422J2_124_3477_n1535, DP_OP_422J2_124_3477_n1534,
         DP_OP_422J2_124_3477_n1533, DP_OP_422J2_124_3477_n1532,
         DP_OP_422J2_124_3477_n1531, DP_OP_422J2_124_3477_n1530,
         DP_OP_422J2_124_3477_n1529, DP_OP_422J2_124_3477_n1528,
         DP_OP_422J2_124_3477_n1527, DP_OP_422J2_124_3477_n1526,
         DP_OP_422J2_124_3477_n1525, DP_OP_422J2_124_3477_n1524,
         DP_OP_422J2_124_3477_n1523, DP_OP_422J2_124_3477_n1522,
         DP_OP_422J2_124_3477_n1521, DP_OP_422J2_124_3477_n1520,
         DP_OP_422J2_124_3477_n1519, DP_OP_422J2_124_3477_n1518,
         DP_OP_422J2_124_3477_n1517, DP_OP_422J2_124_3477_n1516,
         DP_OP_422J2_124_3477_n1515, DP_OP_422J2_124_3477_n1514,
         DP_OP_422J2_124_3477_n1513, DP_OP_422J2_124_3477_n1512,
         DP_OP_422J2_124_3477_n1511, DP_OP_422J2_124_3477_n1510,
         DP_OP_422J2_124_3477_n1509, DP_OP_422J2_124_3477_n1508,
         DP_OP_422J2_124_3477_n1507, DP_OP_422J2_124_3477_n1506,
         DP_OP_422J2_124_3477_n1505, DP_OP_422J2_124_3477_n1504,
         DP_OP_422J2_124_3477_n1503, DP_OP_422J2_124_3477_n1502,
         DP_OP_422J2_124_3477_n1501, DP_OP_422J2_124_3477_n1500,
         DP_OP_422J2_124_3477_n1499, DP_OP_422J2_124_3477_n1498,
         DP_OP_422J2_124_3477_n1497, DP_OP_422J2_124_3477_n1496,
         DP_OP_422J2_124_3477_n1495, DP_OP_422J2_124_3477_n1494,
         DP_OP_422J2_124_3477_n1493, DP_OP_422J2_124_3477_n1492,
         DP_OP_422J2_124_3477_n1491, DP_OP_422J2_124_3477_n1490,
         DP_OP_422J2_124_3477_n1489, DP_OP_422J2_124_3477_n1488,
         DP_OP_422J2_124_3477_n1487, DP_OP_422J2_124_3477_n1486,
         DP_OP_422J2_124_3477_n1485, DP_OP_422J2_124_3477_n1484,
         DP_OP_422J2_124_3477_n1483, DP_OP_422J2_124_3477_n1482,
         DP_OP_422J2_124_3477_n1481, DP_OP_422J2_124_3477_n1480,
         DP_OP_422J2_124_3477_n1479, DP_OP_422J2_124_3477_n1478,
         DP_OP_422J2_124_3477_n1477, DP_OP_422J2_124_3477_n1476,
         DP_OP_422J2_124_3477_n1475, DP_OP_422J2_124_3477_n1474,
         DP_OP_422J2_124_3477_n1473, DP_OP_422J2_124_3477_n1472,
         DP_OP_422J2_124_3477_n1471, DP_OP_422J2_124_3477_n1470,
         DP_OP_422J2_124_3477_n1469, DP_OP_422J2_124_3477_n1468,
         DP_OP_422J2_124_3477_n1467, DP_OP_422J2_124_3477_n1466,
         DP_OP_422J2_124_3477_n1465, DP_OP_422J2_124_3477_n1464,
         DP_OP_422J2_124_3477_n1463, DP_OP_422J2_124_3477_n1462,
         DP_OP_422J2_124_3477_n1461, DP_OP_422J2_124_3477_n1460,
         DP_OP_422J2_124_3477_n1459, DP_OP_422J2_124_3477_n1458,
         DP_OP_422J2_124_3477_n1457, DP_OP_422J2_124_3477_n1456,
         DP_OP_422J2_124_3477_n1455, DP_OP_422J2_124_3477_n1454,
         DP_OP_422J2_124_3477_n1453, DP_OP_422J2_124_3477_n1452,
         DP_OP_422J2_124_3477_n1451, DP_OP_422J2_124_3477_n1450,
         DP_OP_422J2_124_3477_n1449, DP_OP_422J2_124_3477_n1448,
         DP_OP_422J2_124_3477_n1447, DP_OP_422J2_124_3477_n1446,
         DP_OP_422J2_124_3477_n1445, DP_OP_422J2_124_3477_n1444,
         DP_OP_422J2_124_3477_n1443, DP_OP_422J2_124_3477_n1442,
         DP_OP_422J2_124_3477_n1441, DP_OP_422J2_124_3477_n1440,
         DP_OP_422J2_124_3477_n1439, DP_OP_422J2_124_3477_n1438,
         DP_OP_422J2_124_3477_n1437, DP_OP_422J2_124_3477_n1436,
         DP_OP_422J2_124_3477_n1435, DP_OP_422J2_124_3477_n1434,
         DP_OP_422J2_124_3477_n1433, DP_OP_422J2_124_3477_n1432,
         DP_OP_422J2_124_3477_n1431, DP_OP_422J2_124_3477_n1430,
         DP_OP_422J2_124_3477_n1429, DP_OP_422J2_124_3477_n1428,
         DP_OP_422J2_124_3477_n1427, DP_OP_422J2_124_3477_n1426,
         DP_OP_422J2_124_3477_n1425, DP_OP_422J2_124_3477_n1424,
         DP_OP_422J2_124_3477_n1423, DP_OP_422J2_124_3477_n1422,
         DP_OP_422J2_124_3477_n1421, DP_OP_422J2_124_3477_n1420,
         DP_OP_422J2_124_3477_n1419, DP_OP_422J2_124_3477_n1418,
         DP_OP_422J2_124_3477_n1417, DP_OP_422J2_124_3477_n1416,
         DP_OP_422J2_124_3477_n1415, DP_OP_422J2_124_3477_n1414,
         DP_OP_422J2_124_3477_n1413, DP_OP_422J2_124_3477_n1412,
         DP_OP_422J2_124_3477_n1411, DP_OP_422J2_124_3477_n1410,
         DP_OP_422J2_124_3477_n1409, DP_OP_422J2_124_3477_n1408,
         DP_OP_422J2_124_3477_n1407, DP_OP_422J2_124_3477_n1406,
         DP_OP_422J2_124_3477_n1405, DP_OP_422J2_124_3477_n1404,
         DP_OP_422J2_124_3477_n1403, DP_OP_422J2_124_3477_n1402,
         DP_OP_422J2_124_3477_n1401, DP_OP_422J2_124_3477_n1400,
         DP_OP_422J2_124_3477_n1399, DP_OP_422J2_124_3477_n1398,
         DP_OP_422J2_124_3477_n1397, DP_OP_422J2_124_3477_n1396,
         DP_OP_422J2_124_3477_n1395, DP_OP_422J2_124_3477_n1394,
         DP_OP_422J2_124_3477_n1393, DP_OP_422J2_124_3477_n1392,
         DP_OP_422J2_124_3477_n1391, DP_OP_422J2_124_3477_n1390,
         DP_OP_422J2_124_3477_n1389, DP_OP_422J2_124_3477_n1388,
         DP_OP_422J2_124_3477_n1387, DP_OP_422J2_124_3477_n1386,
         DP_OP_422J2_124_3477_n1385, DP_OP_422J2_124_3477_n1384,
         DP_OP_422J2_124_3477_n1383, DP_OP_422J2_124_3477_n1382,
         DP_OP_422J2_124_3477_n1381, DP_OP_422J2_124_3477_n1380,
         DP_OP_422J2_124_3477_n1379, DP_OP_422J2_124_3477_n1378,
         DP_OP_422J2_124_3477_n1377, DP_OP_422J2_124_3477_n1376,
         DP_OP_422J2_124_3477_n1375, DP_OP_422J2_124_3477_n1374,
         DP_OP_422J2_124_3477_n1373, DP_OP_422J2_124_3477_n1372,
         DP_OP_422J2_124_3477_n1371, DP_OP_422J2_124_3477_n1370,
         DP_OP_422J2_124_3477_n1369, DP_OP_422J2_124_3477_n1368,
         DP_OP_422J2_124_3477_n1367, DP_OP_422J2_124_3477_n1366,
         DP_OP_422J2_124_3477_n1365, DP_OP_422J2_124_3477_n1364,
         DP_OP_422J2_124_3477_n1363, DP_OP_422J2_124_3477_n1362,
         DP_OP_422J2_124_3477_n1361, DP_OP_422J2_124_3477_n1360,
         DP_OP_422J2_124_3477_n1359, DP_OP_422J2_124_3477_n1358,
         DP_OP_422J2_124_3477_n1357, DP_OP_422J2_124_3477_n1356,
         DP_OP_422J2_124_3477_n1355, DP_OP_422J2_124_3477_n1354,
         DP_OP_422J2_124_3477_n1353, DP_OP_422J2_124_3477_n1352,
         DP_OP_422J2_124_3477_n1351, DP_OP_422J2_124_3477_n1350,
         DP_OP_422J2_124_3477_n1349, DP_OP_422J2_124_3477_n1348,
         DP_OP_422J2_124_3477_n1347, DP_OP_422J2_124_3477_n1346,
         DP_OP_422J2_124_3477_n1345, DP_OP_422J2_124_3477_n1344,
         DP_OP_422J2_124_3477_n1343, DP_OP_422J2_124_3477_n1342,
         DP_OP_422J2_124_3477_n1341, DP_OP_422J2_124_3477_n1340,
         DP_OP_422J2_124_3477_n1339, DP_OP_422J2_124_3477_n1338,
         DP_OP_422J2_124_3477_n1337, DP_OP_422J2_124_3477_n1336,
         DP_OP_422J2_124_3477_n1335, DP_OP_422J2_124_3477_n1334,
         DP_OP_422J2_124_3477_n1333, DP_OP_422J2_124_3477_n1332,
         DP_OP_422J2_124_3477_n1331, DP_OP_422J2_124_3477_n1330,
         DP_OP_422J2_124_3477_n1329, DP_OP_422J2_124_3477_n1328,
         DP_OP_422J2_124_3477_n1327, DP_OP_422J2_124_3477_n1326,
         DP_OP_422J2_124_3477_n1325, DP_OP_422J2_124_3477_n1324,
         DP_OP_422J2_124_3477_n1323, DP_OP_422J2_124_3477_n1322,
         DP_OP_422J2_124_3477_n1321, DP_OP_422J2_124_3477_n1320,
         DP_OP_422J2_124_3477_n1319, DP_OP_422J2_124_3477_n1318,
         DP_OP_422J2_124_3477_n1317, DP_OP_422J2_124_3477_n1316,
         DP_OP_422J2_124_3477_n1315, DP_OP_422J2_124_3477_n1314,
         DP_OP_422J2_124_3477_n1313, DP_OP_422J2_124_3477_n1312,
         DP_OP_422J2_124_3477_n1311, DP_OP_422J2_124_3477_n1310,
         DP_OP_422J2_124_3477_n1309, DP_OP_422J2_124_3477_n1308,
         DP_OP_422J2_124_3477_n1307, DP_OP_422J2_124_3477_n1306,
         DP_OP_422J2_124_3477_n1305, DP_OP_422J2_124_3477_n1304,
         DP_OP_422J2_124_3477_n1303, DP_OP_422J2_124_3477_n1302,
         DP_OP_422J2_124_3477_n1301, DP_OP_422J2_124_3477_n1300,
         DP_OP_422J2_124_3477_n1299, DP_OP_422J2_124_3477_n1298,
         DP_OP_422J2_124_3477_n1297, DP_OP_422J2_124_3477_n1296,
         DP_OP_422J2_124_3477_n1295, DP_OP_422J2_124_3477_n1294,
         DP_OP_422J2_124_3477_n1293, DP_OP_422J2_124_3477_n1292,
         DP_OP_422J2_124_3477_n1291, DP_OP_422J2_124_3477_n1290,
         DP_OP_422J2_124_3477_n1289, DP_OP_422J2_124_3477_n1288,
         DP_OP_422J2_124_3477_n1287, DP_OP_422J2_124_3477_n1286,
         DP_OP_422J2_124_3477_n1285, DP_OP_422J2_124_3477_n1284,
         DP_OP_422J2_124_3477_n1282, DP_OP_422J2_124_3477_n1281,
         DP_OP_422J2_124_3477_n1280, DP_OP_422J2_124_3477_n1279,
         DP_OP_422J2_124_3477_n1278, DP_OP_422J2_124_3477_n1277,
         DP_OP_422J2_124_3477_n1276, DP_OP_422J2_124_3477_n1275,
         DP_OP_422J2_124_3477_n1274, DP_OP_422J2_124_3477_n1273,
         DP_OP_422J2_124_3477_n1272, DP_OP_422J2_124_3477_n1271,
         DP_OP_422J2_124_3477_n1270, DP_OP_422J2_124_3477_n1269,
         DP_OP_422J2_124_3477_n1268, DP_OP_422J2_124_3477_n1267,
         DP_OP_422J2_124_3477_n1266, DP_OP_422J2_124_3477_n1265,
         DP_OP_422J2_124_3477_n1264, DP_OP_422J2_124_3477_n1263,
         DP_OP_422J2_124_3477_n1262, DP_OP_422J2_124_3477_n1261,
         DP_OP_422J2_124_3477_n1260, DP_OP_422J2_124_3477_n1259,
         DP_OP_422J2_124_3477_n1258, DP_OP_422J2_124_3477_n1257,
         DP_OP_422J2_124_3477_n1256, DP_OP_422J2_124_3477_n1255,
         DP_OP_422J2_124_3477_n1254, DP_OP_422J2_124_3477_n1253,
         DP_OP_422J2_124_3477_n1252, DP_OP_422J2_124_3477_n1251,
         DP_OP_422J2_124_3477_n1250, DP_OP_422J2_124_3477_n1249,
         DP_OP_422J2_124_3477_n1248, DP_OP_422J2_124_3477_n1247,
         DP_OP_422J2_124_3477_n1246, DP_OP_422J2_124_3477_n1245,
         DP_OP_422J2_124_3477_n1244, DP_OP_422J2_124_3477_n1243,
         DP_OP_422J2_124_3477_n1242, DP_OP_422J2_124_3477_n1241,
         DP_OP_422J2_124_3477_n1240, DP_OP_422J2_124_3477_n1239,
         DP_OP_422J2_124_3477_n1238, DP_OP_422J2_124_3477_n1237,
         DP_OP_422J2_124_3477_n1236, DP_OP_422J2_124_3477_n1235,
         DP_OP_422J2_124_3477_n1234, DP_OP_422J2_124_3477_n1233,
         DP_OP_422J2_124_3477_n1232, DP_OP_422J2_124_3477_n1231,
         DP_OP_422J2_124_3477_n1230, DP_OP_422J2_124_3477_n1229,
         DP_OP_422J2_124_3477_n1228, DP_OP_422J2_124_3477_n1227,
         DP_OP_422J2_124_3477_n1226, DP_OP_422J2_124_3477_n1225,
         DP_OP_422J2_124_3477_n1224, DP_OP_422J2_124_3477_n1223,
         DP_OP_422J2_124_3477_n1222, DP_OP_422J2_124_3477_n1221,
         DP_OP_422J2_124_3477_n1220, DP_OP_422J2_124_3477_n1219,
         DP_OP_422J2_124_3477_n1218, DP_OP_422J2_124_3477_n1217,
         DP_OP_422J2_124_3477_n1216, DP_OP_422J2_124_3477_n1215,
         DP_OP_422J2_124_3477_n1214, DP_OP_422J2_124_3477_n1212,
         DP_OP_422J2_124_3477_n1211, DP_OP_422J2_124_3477_n1210,
         DP_OP_422J2_124_3477_n1209, DP_OP_422J2_124_3477_n1208,
         DP_OP_422J2_124_3477_n1207, DP_OP_422J2_124_3477_n1206,
         DP_OP_422J2_124_3477_n1205, DP_OP_422J2_124_3477_n1204,
         DP_OP_422J2_124_3477_n1203, DP_OP_422J2_124_3477_n1202,
         DP_OP_422J2_124_3477_n1201, DP_OP_422J2_124_3477_n1200,
         DP_OP_422J2_124_3477_n1199, DP_OP_422J2_124_3477_n1198,
         DP_OP_422J2_124_3477_n1197, DP_OP_422J2_124_3477_n1196,
         DP_OP_422J2_124_3477_n1195, DP_OP_422J2_124_3477_n1194,
         DP_OP_422J2_124_3477_n1193, DP_OP_422J2_124_3477_n1192,
         DP_OP_422J2_124_3477_n1191, DP_OP_422J2_124_3477_n1190,
         DP_OP_422J2_124_3477_n1189, DP_OP_422J2_124_3477_n1188,
         DP_OP_422J2_124_3477_n1187, DP_OP_422J2_124_3477_n1186,
         DP_OP_422J2_124_3477_n1185, DP_OP_422J2_124_3477_n1184,
         DP_OP_422J2_124_3477_n1183, DP_OP_422J2_124_3477_n1182,
         DP_OP_422J2_124_3477_n1181, DP_OP_422J2_124_3477_n1180,
         DP_OP_422J2_124_3477_n1179, DP_OP_422J2_124_3477_n1178,
         DP_OP_422J2_124_3477_n1177, DP_OP_422J2_124_3477_n1176,
         DP_OP_422J2_124_3477_n1175, DP_OP_422J2_124_3477_n1174,
         DP_OP_422J2_124_3477_n1173, DP_OP_422J2_124_3477_n1172,
         DP_OP_422J2_124_3477_n1171, DP_OP_422J2_124_3477_n1170,
         DP_OP_422J2_124_3477_n1169, DP_OP_422J2_124_3477_n1168,
         DP_OP_422J2_124_3477_n1167, DP_OP_422J2_124_3477_n1166,
         DP_OP_422J2_124_3477_n1165, DP_OP_422J2_124_3477_n1164,
         DP_OP_422J2_124_3477_n1163, DP_OP_422J2_124_3477_n1162,
         DP_OP_422J2_124_3477_n1161, DP_OP_422J2_124_3477_n1160,
         DP_OP_422J2_124_3477_n1159, DP_OP_422J2_124_3477_n1158,
         DP_OP_422J2_124_3477_n1157, DP_OP_422J2_124_3477_n1156,
         DP_OP_422J2_124_3477_n1155, DP_OP_422J2_124_3477_n1154,
         DP_OP_422J2_124_3477_n1153, DP_OP_422J2_124_3477_n1152,
         DP_OP_422J2_124_3477_n1151, DP_OP_422J2_124_3477_n1150,
         DP_OP_422J2_124_3477_n1149, DP_OP_422J2_124_3477_n1148,
         DP_OP_422J2_124_3477_n1147, DP_OP_422J2_124_3477_n1146,
         DP_OP_422J2_124_3477_n1145, DP_OP_422J2_124_3477_n1144,
         DP_OP_422J2_124_3477_n1143, DP_OP_422J2_124_3477_n1142,
         DP_OP_422J2_124_3477_n1141, DP_OP_422J2_124_3477_n1140,
         DP_OP_422J2_124_3477_n1139, DP_OP_422J2_124_3477_n1138,
         DP_OP_422J2_124_3477_n1137, DP_OP_422J2_124_3477_n1136,
         DP_OP_422J2_124_3477_n1135, DP_OP_422J2_124_3477_n1134,
         DP_OP_422J2_124_3477_n1133, DP_OP_422J2_124_3477_n1132,
         DP_OP_422J2_124_3477_n1131, DP_OP_422J2_124_3477_n1130,
         DP_OP_422J2_124_3477_n1129, DP_OP_422J2_124_3477_n1128,
         DP_OP_422J2_124_3477_n1127, DP_OP_422J2_124_3477_n1126,
         DP_OP_422J2_124_3477_n1125, DP_OP_422J2_124_3477_n1124,
         DP_OP_422J2_124_3477_n1123, DP_OP_422J2_124_3477_n1122,
         DP_OP_422J2_124_3477_n1121, DP_OP_422J2_124_3477_n1120,
         DP_OP_422J2_124_3477_n1119, DP_OP_422J2_124_3477_n1118,
         DP_OP_422J2_124_3477_n1117, DP_OP_422J2_124_3477_n1116,
         DP_OP_422J2_124_3477_n1115, DP_OP_422J2_124_3477_n1114,
         DP_OP_422J2_124_3477_n1113, DP_OP_422J2_124_3477_n1112,
         DP_OP_422J2_124_3477_n1111, DP_OP_422J2_124_3477_n1110,
         DP_OP_422J2_124_3477_n1109, DP_OP_422J2_124_3477_n1108,
         DP_OP_422J2_124_3477_n1107, DP_OP_422J2_124_3477_n1106,
         DP_OP_422J2_124_3477_n1105, DP_OP_422J2_124_3477_n1104,
         DP_OP_422J2_124_3477_n1103, DP_OP_422J2_124_3477_n1102,
         DP_OP_422J2_124_3477_n1101, DP_OP_422J2_124_3477_n1100,
         DP_OP_422J2_124_3477_n1099, DP_OP_422J2_124_3477_n1098,
         DP_OP_422J2_124_3477_n1097, DP_OP_422J2_124_3477_n1096,
         DP_OP_422J2_124_3477_n1095, DP_OP_422J2_124_3477_n1094,
         DP_OP_422J2_124_3477_n1093, DP_OP_422J2_124_3477_n1092,
         DP_OP_422J2_124_3477_n1091, DP_OP_422J2_124_3477_n1090,
         DP_OP_422J2_124_3477_n1089, DP_OP_422J2_124_3477_n1088,
         DP_OP_422J2_124_3477_n1087, DP_OP_422J2_124_3477_n1086,
         DP_OP_422J2_124_3477_n1085, DP_OP_422J2_124_3477_n1084,
         DP_OP_422J2_124_3477_n1083, DP_OP_422J2_124_3477_n1082,
         DP_OP_422J2_124_3477_n1081, DP_OP_422J2_124_3477_n1080,
         DP_OP_422J2_124_3477_n1079, DP_OP_422J2_124_3477_n1078,
         DP_OP_422J2_124_3477_n1077, DP_OP_422J2_124_3477_n1076,
         DP_OP_422J2_124_3477_n1075, DP_OP_422J2_124_3477_n1074,
         DP_OP_422J2_124_3477_n1073, DP_OP_422J2_124_3477_n1072,
         DP_OP_422J2_124_3477_n1071, DP_OP_422J2_124_3477_n1070,
         DP_OP_422J2_124_3477_n1069, DP_OP_422J2_124_3477_n1068,
         DP_OP_422J2_124_3477_n1067, DP_OP_422J2_124_3477_n1066,
         DP_OP_422J2_124_3477_n1065, DP_OP_422J2_124_3477_n1064,
         DP_OP_422J2_124_3477_n1063, DP_OP_422J2_124_3477_n1062,
         DP_OP_422J2_124_3477_n1061, DP_OP_422J2_124_3477_n1060,
         DP_OP_422J2_124_3477_n1059, DP_OP_422J2_124_3477_n1058,
         DP_OP_422J2_124_3477_n1057, DP_OP_422J2_124_3477_n1056,
         DP_OP_422J2_124_3477_n1055, DP_OP_422J2_124_3477_n1054,
         DP_OP_422J2_124_3477_n1053, DP_OP_422J2_124_3477_n1052,
         DP_OP_422J2_124_3477_n1051, DP_OP_422J2_124_3477_n1050,
         DP_OP_422J2_124_3477_n1049, DP_OP_422J2_124_3477_n1048,
         DP_OP_422J2_124_3477_n1047, DP_OP_422J2_124_3477_n1046,
         DP_OP_422J2_124_3477_n1045, DP_OP_422J2_124_3477_n1044,
         DP_OP_422J2_124_3477_n1043, DP_OP_422J2_124_3477_n1042,
         DP_OP_422J2_124_3477_n1041, DP_OP_422J2_124_3477_n1040,
         DP_OP_422J2_124_3477_n1039, DP_OP_422J2_124_3477_n1038,
         DP_OP_422J2_124_3477_n1037, DP_OP_422J2_124_3477_n1036,
         DP_OP_422J2_124_3477_n1035, DP_OP_422J2_124_3477_n1034,
         DP_OP_422J2_124_3477_n1033, DP_OP_422J2_124_3477_n1032,
         DP_OP_422J2_124_3477_n1031, DP_OP_422J2_124_3477_n1030,
         DP_OP_422J2_124_3477_n1029, DP_OP_422J2_124_3477_n1028,
         DP_OP_422J2_124_3477_n1027, DP_OP_422J2_124_3477_n1026,
         DP_OP_422J2_124_3477_n1025, DP_OP_422J2_124_3477_n1024,
         DP_OP_422J2_124_3477_n1023, DP_OP_422J2_124_3477_n1022,
         DP_OP_422J2_124_3477_n1021, DP_OP_422J2_124_3477_n1020,
         DP_OP_422J2_124_3477_n1019, DP_OP_422J2_124_3477_n1018,
         DP_OP_422J2_124_3477_n1017, DP_OP_422J2_124_3477_n1016,
         DP_OP_422J2_124_3477_n1015, DP_OP_422J2_124_3477_n1014,
         DP_OP_422J2_124_3477_n1013, DP_OP_422J2_124_3477_n1012,
         DP_OP_422J2_124_3477_n1011, DP_OP_422J2_124_3477_n1010,
         DP_OP_422J2_124_3477_n1009, DP_OP_422J2_124_3477_n1008,
         DP_OP_422J2_124_3477_n1007, DP_OP_422J2_124_3477_n1006,
         DP_OP_422J2_124_3477_n1005, DP_OP_422J2_124_3477_n1004,
         DP_OP_422J2_124_3477_n1003, DP_OP_422J2_124_3477_n1002,
         DP_OP_422J2_124_3477_n1001, DP_OP_422J2_124_3477_n1000,
         DP_OP_422J2_124_3477_n999, DP_OP_422J2_124_3477_n998,
         DP_OP_422J2_124_3477_n997, DP_OP_422J2_124_3477_n996,
         DP_OP_422J2_124_3477_n995, DP_OP_422J2_124_3477_n994,
         DP_OP_422J2_124_3477_n993, DP_OP_422J2_124_3477_n992,
         DP_OP_422J2_124_3477_n991, DP_OP_422J2_124_3477_n990,
         DP_OP_422J2_124_3477_n989, DP_OP_422J2_124_3477_n988,
         DP_OP_422J2_124_3477_n987, DP_OP_422J2_124_3477_n986,
         DP_OP_422J2_124_3477_n985, DP_OP_422J2_124_3477_n984,
         DP_OP_422J2_124_3477_n983, DP_OP_422J2_124_3477_n982,
         DP_OP_422J2_124_3477_n981, DP_OP_422J2_124_3477_n980,
         DP_OP_422J2_124_3477_n979, DP_OP_422J2_124_3477_n978,
         DP_OP_422J2_124_3477_n977, DP_OP_422J2_124_3477_n976,
         DP_OP_422J2_124_3477_n975, DP_OP_422J2_124_3477_n974,
         DP_OP_422J2_124_3477_n973, DP_OP_422J2_124_3477_n972,
         DP_OP_422J2_124_3477_n971, DP_OP_422J2_124_3477_n970,
         DP_OP_422J2_124_3477_n969, DP_OP_422J2_124_3477_n968,
         DP_OP_422J2_124_3477_n967, DP_OP_422J2_124_3477_n966,
         DP_OP_422J2_124_3477_n965, DP_OP_422J2_124_3477_n964,
         DP_OP_422J2_124_3477_n963, DP_OP_422J2_124_3477_n962,
         DP_OP_422J2_124_3477_n961, DP_OP_422J2_124_3477_n960,
         DP_OP_422J2_124_3477_n959, DP_OP_422J2_124_3477_n958,
         DP_OP_422J2_124_3477_n957, DP_OP_422J2_124_3477_n956,
         DP_OP_422J2_124_3477_n955, DP_OP_422J2_124_3477_n954,
         DP_OP_422J2_124_3477_n953, DP_OP_422J2_124_3477_n952,
         DP_OP_422J2_124_3477_n951, DP_OP_422J2_124_3477_n950,
         DP_OP_422J2_124_3477_n949, DP_OP_422J2_124_3477_n948,
         DP_OP_422J2_124_3477_n947, DP_OP_422J2_124_3477_n946,
         DP_OP_422J2_124_3477_n945, DP_OP_422J2_124_3477_n944,
         DP_OP_422J2_124_3477_n943, DP_OP_422J2_124_3477_n942,
         DP_OP_422J2_124_3477_n941, DP_OP_422J2_124_3477_n940,
         DP_OP_422J2_124_3477_n939, DP_OP_422J2_124_3477_n938,
         DP_OP_422J2_124_3477_n937, DP_OP_422J2_124_3477_n936,
         DP_OP_422J2_124_3477_n935, DP_OP_422J2_124_3477_n934,
         DP_OP_422J2_124_3477_n933, DP_OP_422J2_124_3477_n932,
         DP_OP_422J2_124_3477_n931, DP_OP_422J2_124_3477_n930,
         DP_OP_422J2_124_3477_n929, DP_OP_422J2_124_3477_n928,
         DP_OP_422J2_124_3477_n927, DP_OP_422J2_124_3477_n926,
         DP_OP_422J2_124_3477_n925, DP_OP_422J2_124_3477_n924,
         DP_OP_422J2_124_3477_n923, DP_OP_422J2_124_3477_n922,
         DP_OP_422J2_124_3477_n921, DP_OP_422J2_124_3477_n920,
         DP_OP_422J2_124_3477_n919, DP_OP_422J2_124_3477_n918,
         DP_OP_422J2_124_3477_n917, DP_OP_422J2_124_3477_n916,
         DP_OP_422J2_124_3477_n915, DP_OP_422J2_124_3477_n914,
         DP_OP_422J2_124_3477_n913, DP_OP_422J2_124_3477_n912,
         DP_OP_422J2_124_3477_n911, DP_OP_422J2_124_3477_n910,
         DP_OP_422J2_124_3477_n909, DP_OP_422J2_124_3477_n908,
         DP_OP_422J2_124_3477_n907, DP_OP_422J2_124_3477_n906,
         DP_OP_422J2_124_3477_n905, DP_OP_422J2_124_3477_n904,
         DP_OP_422J2_124_3477_n903, DP_OP_422J2_124_3477_n902,
         DP_OP_422J2_124_3477_n901, DP_OP_422J2_124_3477_n900,
         DP_OP_422J2_124_3477_n899, DP_OP_422J2_124_3477_n898,
         DP_OP_422J2_124_3477_n897, DP_OP_422J2_124_3477_n896,
         DP_OP_422J2_124_3477_n895, DP_OP_422J2_124_3477_n894,
         DP_OP_422J2_124_3477_n893, DP_OP_422J2_124_3477_n892,
         DP_OP_422J2_124_3477_n891, DP_OP_422J2_124_3477_n890,
         DP_OP_422J2_124_3477_n889, DP_OP_422J2_124_3477_n888,
         DP_OP_422J2_124_3477_n887, DP_OP_422J2_124_3477_n886,
         DP_OP_422J2_124_3477_n885, DP_OP_422J2_124_3477_n884,
         DP_OP_422J2_124_3477_n883, DP_OP_422J2_124_3477_n882,
         DP_OP_422J2_124_3477_n881, DP_OP_422J2_124_3477_n880,
         DP_OP_422J2_124_3477_n879, DP_OP_422J2_124_3477_n878,
         DP_OP_422J2_124_3477_n877, DP_OP_422J2_124_3477_n876,
         DP_OP_422J2_124_3477_n875, DP_OP_422J2_124_3477_n874,
         DP_OP_422J2_124_3477_n873, DP_OP_422J2_124_3477_n872,
         DP_OP_422J2_124_3477_n871, DP_OP_422J2_124_3477_n870,
         DP_OP_422J2_124_3477_n869, DP_OP_422J2_124_3477_n868,
         DP_OP_422J2_124_3477_n867, DP_OP_422J2_124_3477_n866,
         DP_OP_422J2_124_3477_n865, DP_OP_422J2_124_3477_n864,
         DP_OP_422J2_124_3477_n863, DP_OP_422J2_124_3477_n862,
         DP_OP_422J2_124_3477_n861, DP_OP_422J2_124_3477_n860,
         DP_OP_422J2_124_3477_n859, DP_OP_422J2_124_3477_n858,
         DP_OP_422J2_124_3477_n857, DP_OP_422J2_124_3477_n856,
         DP_OP_422J2_124_3477_n855, DP_OP_422J2_124_3477_n854,
         DP_OP_422J2_124_3477_n853, DP_OP_422J2_124_3477_n852,
         DP_OP_422J2_124_3477_n851, DP_OP_422J2_124_3477_n850,
         DP_OP_422J2_124_3477_n849, DP_OP_422J2_124_3477_n848,
         DP_OP_422J2_124_3477_n847, DP_OP_422J2_124_3477_n846,
         DP_OP_422J2_124_3477_n845, DP_OP_422J2_124_3477_n844,
         DP_OP_422J2_124_3477_n843, DP_OP_422J2_124_3477_n842,
         DP_OP_422J2_124_3477_n841, DP_OP_422J2_124_3477_n840,
         DP_OP_422J2_124_3477_n839, DP_OP_422J2_124_3477_n838,
         DP_OP_422J2_124_3477_n837, DP_OP_422J2_124_3477_n836,
         DP_OP_422J2_124_3477_n835, DP_OP_422J2_124_3477_n834,
         DP_OP_422J2_124_3477_n833, DP_OP_422J2_124_3477_n832,
         DP_OP_422J2_124_3477_n831, DP_OP_422J2_124_3477_n830,
         DP_OP_422J2_124_3477_n829, DP_OP_422J2_124_3477_n828,
         DP_OP_422J2_124_3477_n827, DP_OP_422J2_124_3477_n826,
         DP_OP_422J2_124_3477_n825, DP_OP_422J2_124_3477_n824,
         DP_OP_422J2_124_3477_n823, DP_OP_422J2_124_3477_n822,
         DP_OP_422J2_124_3477_n821, DP_OP_422J2_124_3477_n820,
         DP_OP_422J2_124_3477_n819, DP_OP_422J2_124_3477_n818,
         DP_OP_422J2_124_3477_n817, DP_OP_422J2_124_3477_n816,
         DP_OP_422J2_124_3477_n815, DP_OP_422J2_124_3477_n814,
         DP_OP_422J2_124_3477_n813, DP_OP_422J2_124_3477_n812,
         DP_OP_422J2_124_3477_n811, DP_OP_422J2_124_3477_n810,
         DP_OP_422J2_124_3477_n809, DP_OP_422J2_124_3477_n808,
         DP_OP_422J2_124_3477_n807, DP_OP_422J2_124_3477_n806,
         DP_OP_422J2_124_3477_n805, DP_OP_422J2_124_3477_n804,
         DP_OP_422J2_124_3477_n803, DP_OP_422J2_124_3477_n802,
         DP_OP_422J2_124_3477_n801, DP_OP_422J2_124_3477_n800,
         DP_OP_422J2_124_3477_n799, DP_OP_422J2_124_3477_n798,
         DP_OP_422J2_124_3477_n797, DP_OP_422J2_124_3477_n796,
         DP_OP_422J2_124_3477_n795, DP_OP_422J2_124_3477_n794,
         DP_OP_422J2_124_3477_n793, DP_OP_422J2_124_3477_n792,
         DP_OP_422J2_124_3477_n791, DP_OP_422J2_124_3477_n790,
         DP_OP_422J2_124_3477_n789, DP_OP_422J2_124_3477_n788,
         DP_OP_422J2_124_3477_n787, DP_OP_422J2_124_3477_n786,
         DP_OP_422J2_124_3477_n785, DP_OP_422J2_124_3477_n784,
         DP_OP_422J2_124_3477_n783, DP_OP_422J2_124_3477_n782,
         DP_OP_422J2_124_3477_n781, DP_OP_422J2_124_3477_n780,
         DP_OP_422J2_124_3477_n779, DP_OP_422J2_124_3477_n778,
         DP_OP_422J2_124_3477_n777, DP_OP_422J2_124_3477_n776,
         DP_OP_422J2_124_3477_n775, DP_OP_422J2_124_3477_n774,
         DP_OP_422J2_124_3477_n773, DP_OP_422J2_124_3477_n772,
         DP_OP_422J2_124_3477_n771, DP_OP_422J2_124_3477_n770,
         DP_OP_422J2_124_3477_n769, DP_OP_422J2_124_3477_n768,
         DP_OP_422J2_124_3477_n767, DP_OP_422J2_124_3477_n766,
         DP_OP_422J2_124_3477_n765, DP_OP_422J2_124_3477_n764,
         DP_OP_422J2_124_3477_n763, DP_OP_422J2_124_3477_n762,
         DP_OP_422J2_124_3477_n761, DP_OP_422J2_124_3477_n760,
         DP_OP_422J2_124_3477_n759, DP_OP_422J2_124_3477_n758,
         DP_OP_422J2_124_3477_n757, DP_OP_422J2_124_3477_n756,
         DP_OP_422J2_124_3477_n755, DP_OP_422J2_124_3477_n754,
         DP_OP_422J2_124_3477_n753, DP_OP_422J2_124_3477_n752,
         DP_OP_422J2_124_3477_n751, DP_OP_422J2_124_3477_n750,
         DP_OP_422J2_124_3477_n749, DP_OP_422J2_124_3477_n748,
         DP_OP_422J2_124_3477_n747, DP_OP_422J2_124_3477_n746,
         DP_OP_422J2_124_3477_n745, DP_OP_422J2_124_3477_n744,
         DP_OP_422J2_124_3477_n743, DP_OP_422J2_124_3477_n742,
         DP_OP_422J2_124_3477_n741, DP_OP_422J2_124_3477_n740,
         DP_OP_422J2_124_3477_n739, DP_OP_422J2_124_3477_n738,
         DP_OP_422J2_124_3477_n737, DP_OP_422J2_124_3477_n736,
         DP_OP_422J2_124_3477_n735, DP_OP_422J2_124_3477_n734,
         DP_OP_422J2_124_3477_n733, DP_OP_422J2_124_3477_n732,
         DP_OP_422J2_124_3477_n731, DP_OP_422J2_124_3477_n730,
         DP_OP_422J2_124_3477_n729, DP_OP_422J2_124_3477_n728,
         DP_OP_422J2_124_3477_n727, DP_OP_422J2_124_3477_n726,
         DP_OP_422J2_124_3477_n725, DP_OP_422J2_124_3477_n724,
         DP_OP_422J2_124_3477_n723, DP_OP_422J2_124_3477_n722,
         DP_OP_422J2_124_3477_n721, DP_OP_422J2_124_3477_n720,
         DP_OP_422J2_124_3477_n719, DP_OP_422J2_124_3477_n718,
         DP_OP_422J2_124_3477_n717, DP_OP_422J2_124_3477_n716,
         DP_OP_422J2_124_3477_n715, DP_OP_422J2_124_3477_n714,
         DP_OP_422J2_124_3477_n713, DP_OP_422J2_124_3477_n712,
         DP_OP_422J2_124_3477_n711, DP_OP_422J2_124_3477_n710,
         DP_OP_422J2_124_3477_n709, DP_OP_422J2_124_3477_n708,
         DP_OP_422J2_124_3477_n707, DP_OP_422J2_124_3477_n706,
         DP_OP_422J2_124_3477_n705, DP_OP_422J2_124_3477_n704,
         DP_OP_422J2_124_3477_n703, DP_OP_422J2_124_3477_n702,
         DP_OP_422J2_124_3477_n701, DP_OP_422J2_124_3477_n700,
         DP_OP_422J2_124_3477_n699, DP_OP_422J2_124_3477_n698,
         DP_OP_422J2_124_3477_n697, DP_OP_422J2_124_3477_n696,
         DP_OP_422J2_124_3477_n695, DP_OP_422J2_124_3477_n694,
         DP_OP_422J2_124_3477_n693, DP_OP_422J2_124_3477_n692,
         DP_OP_422J2_124_3477_n691, DP_OP_422J2_124_3477_n690,
         DP_OP_422J2_124_3477_n689, DP_OP_422J2_124_3477_n688,
         DP_OP_422J2_124_3477_n687, DP_OP_422J2_124_3477_n686,
         DP_OP_422J2_124_3477_n685, DP_OP_422J2_124_3477_n684,
         DP_OP_422J2_124_3477_n683, DP_OP_422J2_124_3477_n682,
         DP_OP_422J2_124_3477_n681, DP_OP_422J2_124_3477_n680,
         DP_OP_422J2_124_3477_n679, DP_OP_422J2_124_3477_n678,
         DP_OP_422J2_124_3477_n677, DP_OP_422J2_124_3477_n676,
         DP_OP_422J2_124_3477_n675, DP_OP_422J2_124_3477_n674,
         DP_OP_422J2_124_3477_n673, DP_OP_422J2_124_3477_n672,
         DP_OP_422J2_124_3477_n671, DP_OP_422J2_124_3477_n670,
         DP_OP_422J2_124_3477_n669, DP_OP_422J2_124_3477_n668,
         DP_OP_422J2_124_3477_n667, DP_OP_422J2_124_3477_n666,
         DP_OP_422J2_124_3477_n665, DP_OP_422J2_124_3477_n664,
         DP_OP_422J2_124_3477_n663, DP_OP_422J2_124_3477_n662,
         DP_OP_422J2_124_3477_n661, DP_OP_422J2_124_3477_n660,
         DP_OP_422J2_124_3477_n659, DP_OP_422J2_124_3477_n658,
         DP_OP_422J2_124_3477_n657, DP_OP_422J2_124_3477_n656,
         DP_OP_422J2_124_3477_n655, DP_OP_422J2_124_3477_n654,
         DP_OP_422J2_124_3477_n653, DP_OP_422J2_124_3477_n652,
         DP_OP_422J2_124_3477_n651, DP_OP_422J2_124_3477_n650,
         DP_OP_422J2_124_3477_n649, DP_OP_422J2_124_3477_n648,
         DP_OP_422J2_124_3477_n647, DP_OP_422J2_124_3477_n646,
         DP_OP_422J2_124_3477_n645, DP_OP_422J2_124_3477_n644,
         DP_OP_422J2_124_3477_n643, DP_OP_422J2_124_3477_n642,
         DP_OP_422J2_124_3477_n641, DP_OP_422J2_124_3477_n640,
         DP_OP_422J2_124_3477_n639, DP_OP_422J2_124_3477_n638,
         DP_OP_422J2_124_3477_n637, DP_OP_422J2_124_3477_n636,
         DP_OP_422J2_124_3477_n635, DP_OP_422J2_124_3477_n634,
         DP_OP_422J2_124_3477_n633, DP_OP_422J2_124_3477_n632,
         DP_OP_422J2_124_3477_n631, DP_OP_422J2_124_3477_n630,
         DP_OP_422J2_124_3477_n629, DP_OP_422J2_124_3477_n628,
         DP_OP_422J2_124_3477_n627, DP_OP_422J2_124_3477_n626,
         DP_OP_422J2_124_3477_n625, DP_OP_422J2_124_3477_n624,
         DP_OP_422J2_124_3477_n623, DP_OP_422J2_124_3477_n622,
         DP_OP_422J2_124_3477_n621, DP_OP_422J2_124_3477_n620,
         DP_OP_422J2_124_3477_n619, DP_OP_422J2_124_3477_n618,
         DP_OP_422J2_124_3477_n617, DP_OP_422J2_124_3477_n616,
         DP_OP_422J2_124_3477_n615, DP_OP_422J2_124_3477_n614,
         DP_OP_422J2_124_3477_n613, DP_OP_422J2_124_3477_n612,
         DP_OP_422J2_124_3477_n611, DP_OP_422J2_124_3477_n610,
         DP_OP_422J2_124_3477_n609, DP_OP_422J2_124_3477_n608,
         DP_OP_422J2_124_3477_n607, DP_OP_422J2_124_3477_n606,
         DP_OP_422J2_124_3477_n605, DP_OP_422J2_124_3477_n604,
         DP_OP_422J2_124_3477_n603, DP_OP_422J2_124_3477_n602,
         DP_OP_422J2_124_3477_n601, DP_OP_422J2_124_3477_n600,
         DP_OP_422J2_124_3477_n599, DP_OP_422J2_124_3477_n598,
         DP_OP_422J2_124_3477_n597, DP_OP_422J2_124_3477_n596,
         DP_OP_422J2_124_3477_n595, DP_OP_422J2_124_3477_n594,
         DP_OP_422J2_124_3477_n593, DP_OP_422J2_124_3477_n592,
         DP_OP_422J2_124_3477_n591, DP_OP_422J2_124_3477_n590,
         DP_OP_422J2_124_3477_n589, DP_OP_422J2_124_3477_n588,
         DP_OP_422J2_124_3477_n587, DP_OP_422J2_124_3477_n586,
         DP_OP_422J2_124_3477_n585, DP_OP_422J2_124_3477_n584,
         DP_OP_422J2_124_3477_n583, DP_OP_422J2_124_3477_n582,
         DP_OP_422J2_124_3477_n581, DP_OP_422J2_124_3477_n580,
         DP_OP_422J2_124_3477_n579, DP_OP_422J2_124_3477_n578,
         DP_OP_422J2_124_3477_n577, DP_OP_422J2_124_3477_n576,
         DP_OP_422J2_124_3477_n575, DP_OP_422J2_124_3477_n574,
         DP_OP_422J2_124_3477_n573, DP_OP_422J2_124_3477_n572,
         DP_OP_422J2_124_3477_n571, DP_OP_422J2_124_3477_n570,
         DP_OP_422J2_124_3477_n569, DP_OP_422J2_124_3477_n568,
         DP_OP_422J2_124_3477_n567, DP_OP_422J2_124_3477_n566,
         DP_OP_422J2_124_3477_n565, DP_OP_422J2_124_3477_n564,
         DP_OP_422J2_124_3477_n563, DP_OP_422J2_124_3477_n562,
         DP_OP_422J2_124_3477_n561, DP_OP_422J2_124_3477_n560,
         DP_OP_422J2_124_3477_n559, DP_OP_422J2_124_3477_n558,
         DP_OP_422J2_124_3477_n557, DP_OP_422J2_124_3477_n556,
         DP_OP_422J2_124_3477_n555, DP_OP_422J2_124_3477_n554,
         DP_OP_422J2_124_3477_n553, DP_OP_422J2_124_3477_n552,
         DP_OP_422J2_124_3477_n551, DP_OP_422J2_124_3477_n550,
         DP_OP_422J2_124_3477_n549, DP_OP_422J2_124_3477_n548,
         DP_OP_422J2_124_3477_n547, DP_OP_422J2_124_3477_n546,
         DP_OP_422J2_124_3477_n545, DP_OP_422J2_124_3477_n544,
         DP_OP_422J2_124_3477_n543, DP_OP_422J2_124_3477_n542,
         DP_OP_422J2_124_3477_n541, DP_OP_422J2_124_3477_n540,
         DP_OP_422J2_124_3477_n539, DP_OP_422J2_124_3477_n538,
         DP_OP_422J2_124_3477_n537, DP_OP_422J2_124_3477_n536,
         DP_OP_422J2_124_3477_n535, DP_OP_422J2_124_3477_n534,
         DP_OP_422J2_124_3477_n533, DP_OP_422J2_124_3477_n532,
         DP_OP_422J2_124_3477_n531, DP_OP_422J2_124_3477_n530,
         DP_OP_422J2_124_3477_n529, DP_OP_422J2_124_3477_n528,
         DP_OP_422J2_124_3477_n527, DP_OP_422J2_124_3477_n526,
         DP_OP_422J2_124_3477_n525, DP_OP_422J2_124_3477_n524,
         DP_OP_422J2_124_3477_n523, DP_OP_422J2_124_3477_n522,
         DP_OP_422J2_124_3477_n521, DP_OP_422J2_124_3477_n520,
         DP_OP_422J2_124_3477_n519, DP_OP_422J2_124_3477_n518,
         DP_OP_422J2_124_3477_n517, DP_OP_422J2_124_3477_n515,
         DP_OP_422J2_124_3477_n514, DP_OP_422J2_124_3477_n513,
         DP_OP_422J2_124_3477_n512, DP_OP_422J2_124_3477_n511,
         DP_OP_422J2_124_3477_n510, DP_OP_422J2_124_3477_n509,
         DP_OP_422J2_124_3477_n508, DP_OP_422J2_124_3477_n507,
         DP_OP_422J2_124_3477_n506, DP_OP_422J2_124_3477_n505,
         DP_OP_422J2_124_3477_n504, DP_OP_422J2_124_3477_n503,
         DP_OP_422J2_124_3477_n502, DP_OP_422J2_124_3477_n501,
         DP_OP_422J2_124_3477_n500, DP_OP_422J2_124_3477_n499,
         DP_OP_422J2_124_3477_n498, DP_OP_422J2_124_3477_n497,
         DP_OP_422J2_124_3477_n496, DP_OP_422J2_124_3477_n495,
         DP_OP_422J2_124_3477_n494, DP_OP_422J2_124_3477_n493,
         DP_OP_422J2_124_3477_n492, DP_OP_422J2_124_3477_n491,
         DP_OP_422J2_124_3477_n490, DP_OP_422J2_124_3477_n489,
         DP_OP_422J2_124_3477_n488, DP_OP_422J2_124_3477_n487,
         DP_OP_422J2_124_3477_n486, DP_OP_422J2_124_3477_n485,
         DP_OP_422J2_124_3477_n484, DP_OP_422J2_124_3477_n483,
         DP_OP_422J2_124_3477_n482, DP_OP_422J2_124_3477_n481,
         DP_OP_422J2_124_3477_n480, DP_OP_422J2_124_3477_n479,
         DP_OP_422J2_124_3477_n478, DP_OP_422J2_124_3477_n477,
         DP_OP_422J2_124_3477_n476, DP_OP_422J2_124_3477_n475,
         DP_OP_422J2_124_3477_n474, DP_OP_422J2_124_3477_n473,
         DP_OP_422J2_124_3477_n472, DP_OP_422J2_124_3477_n471,
         DP_OP_422J2_124_3477_n470, DP_OP_422J2_124_3477_n469,
         DP_OP_422J2_124_3477_n468, DP_OP_422J2_124_3477_n467,
         DP_OP_422J2_124_3477_n466, DP_OP_422J2_124_3477_n465,
         DP_OP_422J2_124_3477_n464, DP_OP_422J2_124_3477_n463,
         DP_OP_422J2_124_3477_n462, DP_OP_422J2_124_3477_n461,
         DP_OP_422J2_124_3477_n460, DP_OP_422J2_124_3477_n459,
         DP_OP_422J2_124_3477_n458, DP_OP_422J2_124_3477_n457,
         DP_OP_422J2_124_3477_n456, DP_OP_422J2_124_3477_n455,
         DP_OP_422J2_124_3477_n454, DP_OP_422J2_124_3477_n453,
         DP_OP_422J2_124_3477_n452, DP_OP_422J2_124_3477_n451,
         DP_OP_422J2_124_3477_n450, DP_OP_422J2_124_3477_n449,
         DP_OP_422J2_124_3477_n448, DP_OP_422J2_124_3477_n447,
         DP_OP_422J2_124_3477_n446, DP_OP_422J2_124_3477_n445,
         DP_OP_422J2_124_3477_n444, DP_OP_422J2_124_3477_n443,
         DP_OP_422J2_124_3477_n442, DP_OP_422J2_124_3477_n441,
         DP_OP_422J2_124_3477_n440, DP_OP_422J2_124_3477_n439,
         DP_OP_422J2_124_3477_n438, DP_OP_422J2_124_3477_n437,
         DP_OP_422J2_124_3477_n436, DP_OP_422J2_124_3477_n435,
         DP_OP_422J2_124_3477_n434, DP_OP_422J2_124_3477_n433,
         DP_OP_422J2_124_3477_n432, DP_OP_422J2_124_3477_n431,
         DP_OP_422J2_124_3477_n430, DP_OP_422J2_124_3477_n429,
         DP_OP_422J2_124_3477_n428, DP_OP_422J2_124_3477_n427,
         DP_OP_422J2_124_3477_n426, DP_OP_422J2_124_3477_n425,
         DP_OP_422J2_124_3477_n424, DP_OP_422J2_124_3477_n423,
         DP_OP_422J2_124_3477_n422, DP_OP_422J2_124_3477_n421,
         DP_OP_422J2_124_3477_n420, DP_OP_422J2_124_3477_n419,
         DP_OP_422J2_124_3477_n418, DP_OP_422J2_124_3477_n417,
         DP_OP_422J2_124_3477_n416, DP_OP_422J2_124_3477_n415,
         DP_OP_422J2_124_3477_n414, DP_OP_422J2_124_3477_n413,
         DP_OP_422J2_124_3477_n412, DP_OP_422J2_124_3477_n411,
         DP_OP_422J2_124_3477_n410, DP_OP_422J2_124_3477_n409,
         DP_OP_422J2_124_3477_n408, DP_OP_422J2_124_3477_n407,
         DP_OP_422J2_124_3477_n406, DP_OP_422J2_124_3477_n405,
         DP_OP_422J2_124_3477_n404, DP_OP_422J2_124_3477_n403,
         DP_OP_422J2_124_3477_n402, DP_OP_422J2_124_3477_n401,
         DP_OP_422J2_124_3477_n400, DP_OP_422J2_124_3477_n399,
         DP_OP_422J2_124_3477_n398, DP_OP_422J2_124_3477_n397,
         DP_OP_422J2_124_3477_n396, DP_OP_422J2_124_3477_n395,
         DP_OP_422J2_124_3477_n394, DP_OP_422J2_124_3477_n393,
         DP_OP_422J2_124_3477_n392, DP_OP_422J2_124_3477_n391,
         DP_OP_422J2_124_3477_n390, DP_OP_422J2_124_3477_n389,
         DP_OP_422J2_124_3477_n388, DP_OP_422J2_124_3477_n387,
         DP_OP_422J2_124_3477_n386, DP_OP_422J2_124_3477_n385,
         DP_OP_422J2_124_3477_n384, DP_OP_422J2_124_3477_n383,
         DP_OP_422J2_124_3477_n382, DP_OP_422J2_124_3477_n381,
         DP_OP_422J2_124_3477_n380, DP_OP_422J2_124_3477_n379,
         DP_OP_422J2_124_3477_n378, DP_OP_422J2_124_3477_n377,
         DP_OP_422J2_124_3477_n376, DP_OP_422J2_124_3477_n375,
         DP_OP_422J2_124_3477_n374, DP_OP_422J2_124_3477_n373,
         DP_OP_422J2_124_3477_n371, DP_OP_422J2_124_3477_n370,
         DP_OP_422J2_124_3477_n369, DP_OP_422J2_124_3477_n368,
         DP_OP_422J2_124_3477_n367, DP_OP_422J2_124_3477_n366,
         DP_OP_422J2_124_3477_n365, DP_OP_422J2_124_3477_n364,
         DP_OP_422J2_124_3477_n363, DP_OP_422J2_124_3477_n362,
         DP_OP_422J2_124_3477_n361, DP_OP_422J2_124_3477_n360,
         DP_OP_422J2_124_3477_n359, DP_OP_422J2_124_3477_n358,
         DP_OP_422J2_124_3477_n357, DP_OP_422J2_124_3477_n356,
         DP_OP_422J2_124_3477_n355, DP_OP_422J2_124_3477_n354,
         DP_OP_422J2_124_3477_n353, DP_OP_422J2_124_3477_n352,
         DP_OP_422J2_124_3477_n351, DP_OP_422J2_124_3477_n350,
         DP_OP_422J2_124_3477_n349, DP_OP_422J2_124_3477_n348,
         DP_OP_422J2_124_3477_n347, DP_OP_422J2_124_3477_n346,
         DP_OP_422J2_124_3477_n345, DP_OP_422J2_124_3477_n344,
         DP_OP_422J2_124_3477_n343, DP_OP_422J2_124_3477_n342,
         DP_OP_422J2_124_3477_n341, DP_OP_422J2_124_3477_n340,
         DP_OP_422J2_124_3477_n339, DP_OP_422J2_124_3477_n338,
         DP_OP_422J2_124_3477_n337, DP_OP_422J2_124_3477_n336,
         DP_OP_422J2_124_3477_n335, DP_OP_422J2_124_3477_n334,
         DP_OP_422J2_124_3477_n333, DP_OP_422J2_124_3477_n332,
         DP_OP_422J2_124_3477_n331, DP_OP_422J2_124_3477_n330,
         DP_OP_422J2_124_3477_n329, DP_OP_422J2_124_3477_n328,
         DP_OP_422J2_124_3477_n327, DP_OP_422J2_124_3477_n326,
         DP_OP_422J2_124_3477_n325, DP_OP_422J2_124_3477_n324,
         DP_OP_422J2_124_3477_n323, DP_OP_422J2_124_3477_n322,
         DP_OP_422J2_124_3477_n321, DP_OP_422J2_124_3477_n320,
         DP_OP_422J2_124_3477_n319, DP_OP_422J2_124_3477_n318,
         DP_OP_422J2_124_3477_n317, DP_OP_422J2_124_3477_n316,
         DP_OP_422J2_124_3477_n315, DP_OP_422J2_124_3477_n314,
         DP_OP_422J2_124_3477_n313, DP_OP_422J2_124_3477_n312,
         DP_OP_422J2_124_3477_n311, DP_OP_422J2_124_3477_n310,
         DP_OP_422J2_124_3477_n309, DP_OP_422J2_124_3477_n308,
         DP_OP_422J2_124_3477_n306, DP_OP_422J2_124_3477_n305,
         DP_OP_422J2_124_3477_n304, DP_OP_422J2_124_3477_n303,
         DP_OP_422J2_124_3477_n302, DP_OP_422J2_124_3477_n286,
         DP_OP_422J2_124_3477_n285, DP_OP_422J2_124_3477_n284,
         DP_OP_422J2_124_3477_n283, DP_OP_422J2_124_3477_n282,
         DP_OP_422J2_124_3477_n281, DP_OP_422J2_124_3477_n280,
         DP_OP_422J2_124_3477_n279, DP_OP_422J2_124_3477_n277,
         DP_OP_422J2_124_3477_n276, DP_OP_422J2_124_3477_n274,
         DP_OP_422J2_124_3477_n272, DP_OP_422J2_124_3477_n269,
         DP_OP_422J2_124_3477_n268, DP_OP_422J2_124_3477_n267,
         DP_OP_422J2_124_3477_n266, DP_OP_422J2_124_3477_n265,
         DP_OP_422J2_124_3477_n261, DP_OP_422J2_124_3477_n260,
         DP_OP_422J2_124_3477_n259, DP_OP_422J2_124_3477_n258,
         DP_OP_422J2_124_3477_n257, DP_OP_422J2_124_3477_n253,
         DP_OP_422J2_124_3477_n252, DP_OP_422J2_124_3477_n251,
         DP_OP_422J2_124_3477_n249, DP_OP_422J2_124_3477_n248,
         DP_OP_422J2_124_3477_n245, DP_OP_422J2_124_3477_n244,
         DP_OP_422J2_124_3477_n242, DP_OP_422J2_124_3477_n241,
         DP_OP_422J2_124_3477_n240, DP_OP_422J2_124_3477_n237,
         DP_OP_422J2_124_3477_n236, DP_OP_422J2_124_3477_n233,
         DP_OP_422J2_124_3477_n232, DP_OP_422J2_124_3477_n226,
         DP_OP_422J2_124_3477_n220, DP_OP_422J2_124_3477_n219,
         DP_OP_422J2_124_3477_n217, DP_OP_422J2_124_3477_n214,
         DP_OP_422J2_124_3477_n213, DP_OP_422J2_124_3477_n212,
         DP_OP_422J2_124_3477_n210, DP_OP_422J2_124_3477_n209,
         DP_OP_422J2_124_3477_n198, DP_OP_422J2_124_3477_n197,
         DP_OP_422J2_124_3477_n190, DP_OP_422J2_124_3477_n189,
         DP_OP_422J2_124_3477_n188, DP_OP_422J2_124_3477_n187,
         DP_OP_422J2_124_3477_n185, DP_OP_422J2_124_3477_n182,
         DP_OP_422J2_124_3477_n179, DP_OP_422J2_124_3477_n177,
         DP_OP_422J2_124_3477_n176, DP_OP_422J2_124_3477_n174,
         DP_OP_422J2_124_3477_n171, DP_OP_422J2_124_3477_n170,
         DP_OP_422J2_124_3477_n169, DP_OP_422J2_124_3477_n167,
         DP_OP_422J2_124_3477_n166, DP_OP_422J2_124_3477_n165,
         DP_OP_422J2_124_3477_n162, DP_OP_422J2_124_3477_n161,
         DP_OP_422J2_124_3477_n160, DP_OP_422J2_124_3477_n159,
         DP_OP_422J2_124_3477_n158, DP_OP_422J2_124_3477_n156,
         DP_OP_422J2_124_3477_n153, DP_OP_422J2_124_3477_n152,
         DP_OP_422J2_124_3477_n151, DP_OP_422J2_124_3477_n149,
         DP_OP_422J2_124_3477_n148, DP_OP_422J2_124_3477_n146,
         DP_OP_422J2_124_3477_n145, DP_OP_422J2_124_3477_n144,
         DP_OP_422J2_124_3477_n142, DP_OP_422J2_124_3477_n141,
         DP_OP_422J2_124_3477_n140, DP_OP_422J2_124_3477_n139,
         DP_OP_422J2_124_3477_n138, DP_OP_422J2_124_3477_n136,
         DP_OP_422J2_124_3477_n133, DP_OP_422J2_124_3477_n131,
         DP_OP_422J2_124_3477_n129, DP_OP_422J2_124_3477_n128,
         DP_OP_422J2_124_3477_n127, DP_OP_422J2_124_3477_n126,
         DP_OP_422J2_124_3477_n125, DP_OP_422J2_124_3477_n124,
         DP_OP_422J2_124_3477_n122, DP_OP_422J2_124_3477_n120,
         DP_OP_422J2_124_3477_n115, DP_OP_422J2_124_3477_n114,
         DP_OP_422J2_124_3477_n111, DP_OP_422J2_124_3477_n110,
         DP_OP_422J2_124_3477_n109, DP_OP_422J2_124_3477_n107,
         DP_OP_422J2_124_3477_n105, DP_OP_422J2_124_3477_n102,
         DP_OP_422J2_124_3477_n100, DP_OP_422J2_124_3477_n98,
         DP_OP_422J2_124_3477_n97, DP_OP_422J2_124_3477_n96,
         DP_OP_422J2_124_3477_n95, DP_OP_422J2_124_3477_n94,
         DP_OP_422J2_124_3477_n93, DP_OP_422J2_124_3477_n91,
         DP_OP_422J2_124_3477_n89, DP_OP_422J2_124_3477_n85,
         DP_OP_422J2_124_3477_n82, DP_OP_422J2_124_3477_n80,
         DP_OP_422J2_124_3477_n78, DP_OP_422J2_124_3477_n77,
         DP_OP_422J2_124_3477_n75, DP_OP_422J2_124_3477_n73,
         DP_OP_422J2_124_3477_n72, DP_OP_422J2_124_3477_n71,
         DP_OP_422J2_124_3477_n69, DP_OP_422J2_124_3477_n68,
         DP_OP_422J2_124_3477_n67, DP_OP_422J2_124_3477_n65,
         DP_OP_422J2_124_3477_n60, DP_OP_422J2_124_3477_n58,
         DP_OP_422J2_124_3477_n57, DP_OP_422J2_124_3477_n56,
         DP_OP_422J2_124_3477_n55, DP_OP_422J2_124_3477_n54,
         DP_OP_422J2_124_3477_n52, DP_OP_422J2_124_3477_n51,
         DP_OP_422J2_124_3477_n50, DP_OP_422J2_124_3477_n49,
         DP_OP_422J2_124_3477_n47, DP_OP_422J2_124_3477_n38,
         DP_OP_422J2_124_3477_n22, DP_OP_422J2_124_3477_n5,
         DP_OP_422J2_124_3477_n4, DP_OP_422J2_124_3477_n2, n1, n2, n3, n4, n5,
         n6, n7010, n8, n9010, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n7000, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n9000, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n7001, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n9001, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n977, n978, n979, n980, n981, n982, n983,
         n984, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1011, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1069, n1071,
         n1072, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1120, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178;
  wire   [31:0] conv2_sum_a;
  wire   [31:0] conv2_sum_b;
  wire   [31:0] tmp_big1;
  wire   [31:0] conv2_sum_c;
  wire   [31:0] conv2_sum_d;
  wire   [31:0] tmp_big2;
  wire   [67:0] conv_weight_box;
  wire   [31:0] n_conv2_sum_a;
  wire   [31:0] n_conv2_sum_b;
  wire   [31:0] n_conv2_sum_c;
  wire   [31:0] n_conv2_sum_d;

  DFFSSRX1_HVT conv2_sum_c_reg_31_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_c[31]), .CLK(clk), .Q(conv2_sum_c[31]), .QN(n1324) );
  DFFSSRX1_HVT conv2_sum_c_reg_30_ ( .D(1'b0), .SETB(n1445), .RSTB(
        n_conv2_sum_c[30]), .CLK(clk), .Q(conv2_sum_c[30]), .QN(n1913) );
  DFFSSRX1_HVT conv2_sum_c_reg_29_ ( .D(1'b0), .SETB(n1495), .RSTB(
        n_conv2_sum_c[29]), .CLK(clk), .Q(conv2_sum_c[29]), .QN(n1917) );
  DFFSSRX1_HVT conv2_sum_c_reg_28_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_c[28]), .CLK(clk), .Q(conv2_sum_c[28]), .QN(n1897) );
  DFFSSRX1_HVT conv2_sum_c_reg_27_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_c[27]), .CLK(clk), .Q(conv2_sum_c[27]), .QN(n1911) );
  DFFSSRX1_HVT conv2_sum_c_reg_26_ ( .D(1'b0), .SETB(n1434), .RSTB(
        n_conv2_sum_c[26]), .CLK(clk), .Q(conv2_sum_c[26]), .QN(n1896) );
  DFFSSRX1_HVT conv2_sum_c_reg_25_ ( .D(1'b0), .SETB(n1495), .RSTB(
        n_conv2_sum_c[25]), .CLK(clk), .Q(conv2_sum_c[25]), .QN(n1910) );
  DFFSSRX1_HVT conv2_sum_c_reg_24_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_c[24]), .CLK(clk), .Q(conv2_sum_c[24]), .QN(n1895) );
  DFFSSRX1_HVT conv2_sum_c_reg_23_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_c[23]), .CLK(clk), .Q(conv2_sum_c[23]), .QN(n1909) );
  DFFSSRX1_HVT conv2_sum_c_reg_22_ ( .D(1'b0), .SETB(n1445), .RSTB(
        n_conv2_sum_c[22]), .CLK(clk), .Q(conv2_sum_c[22]), .QN(n1894) );
  DFFSSRX1_HVT conv2_sum_c_reg_21_ ( .D(1'b0), .SETB(n1495), .RSTB(
        n_conv2_sum_c[21]), .CLK(clk), .Q(conv2_sum_c[21]), .QN(n1908) );
  DFFSSRX1_HVT conv2_sum_c_reg_20_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_c[20]), .CLK(clk), .Q(conv2_sum_c[20]), .QN(n1893) );
  DFFSSRX1_HVT conv2_sum_c_reg_19_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_c[19]), .CLK(clk), .Q(conv2_sum_c[19]), .QN(n1907) );
  DFFSSRX1_HVT conv2_sum_c_reg_18_ ( .D(1'b0), .SETB(n1434), .RSTB(
        n_conv2_sum_c[18]), .CLK(clk), .Q(conv2_sum_c[18]), .QN(n1892) );
  DFFSSRX1_HVT conv2_sum_c_reg_17_ ( .D(1'b0), .SETB(n1495), .RSTB(
        n_conv2_sum_c[17]), .CLK(clk), .Q(conv2_sum_c[17]), .QN(n1906) );
  DFFSSRX1_HVT conv2_sum_c_reg_16_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_c[16]), .CLK(clk), .Q(conv2_sum_c[16]), .QN(n1319) );
  DFFSSRX1_HVT conv2_sum_c_reg_15_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_c[15]), .CLK(clk), .Q(conv2_sum_c[15]), .QN(n1905) );
  DFFSSRX1_HVT conv2_sum_c_reg_14_ ( .D(1'b0), .SETB(n1445), .RSTB(
        n_conv2_sum_c[14]), .CLK(clk), .Q(conv2_sum_c[14]), .QN(n1891) );
  DFFSSRX1_HVT conv2_sum_c_reg_13_ ( .D(1'b0), .SETB(n1495), .RSTB(
        n_conv2_sum_c[13]), .CLK(clk), .Q(conv2_sum_c[13]), .QN(n1904) );
  DFFSSRX1_HVT conv2_sum_c_reg_12_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_c[12]), .CLK(clk), .Q(conv2_sum_c[12]), .QN(n1868) );
  DFFSSRX1_HVT conv2_sum_c_reg_11_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_c[11]), .CLK(clk), .Q(conv2_sum_c[11]), .QN(n1982) );
  DFFSSRX1_HVT conv2_sum_c_reg_10_ ( .D(1'b0), .SETB(n1434), .RSTB(
        n_conv2_sum_c[10]), .CLK(clk), .Q(conv2_sum_c[10]), .QN(n1860) );
  DFFSSRX1_HVT conv2_sum_c_reg_9_ ( .D(1'b0), .SETB(n1495), .RSTB(
        n_conv2_sum_c[9]), .CLK(clk), .Q(conv2_sum_c[9]), .QN(n1993) );
  DFFSSRX1_HVT conv2_sum_c_reg_8_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_c[8]), .CLK(clk), .Q(conv2_sum_c[8]), .QN(n1286) );
  DFFSSRX1_HVT conv2_sum_c_reg_7_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_c[7]), .CLK(clk), .Q(conv2_sum_c[7]), .QN(n1855) );
  DFFSSRX1_HVT conv2_sum_c_reg_6_ ( .D(1'b0), .SETB(n1445), .RSTB(
        n_conv2_sum_c[6]), .CLK(clk), .Q(conv2_sum_c[6]), .QN(n1862) );
  DFFSSRX1_HVT conv2_sum_c_reg_5_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_c[5]), .CLK(clk), .Q(conv2_sum_c[5]), .QN(n1854) );
  DFFSSRX1_HVT conv2_sum_c_reg_4_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_c[4]), .CLK(clk), .Q(conv2_sum_c[4]), .QN(n1859) );
  DFFSSRX1_HVT conv2_sum_c_reg_2_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_c[2]), .CLK(clk), .Q(conv2_sum_c[2]), .QN(n1865) );
  DFFSSRX1_HVT conv2_sum_c_reg_1_ ( .D(1'b0), .SETB(n1434), .RSTB(
        n_conv2_sum_c[1]), .CLK(clk), .Q(conv2_sum_c[1]), .QN(n1980) );
  DFFSSRX1_HVT conv2_sum_c_reg_0_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_c[0]), .CLK(clk), .Q(conv2_sum_c[0]), .QN(n1292) );
  DFFSSRX1_HVT conv2_sum_d_reg_31_ ( .D(1'b0), .SETB(n1495), .RSTB(
        n_conv2_sum_d[31]), .CLK(clk), .Q(conv2_sum_d[31]), .QN(n1915) );
  DFFSSRX1_HVT conv2_sum_d_reg_30_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_d[30]), .CLK(clk), .Q(conv2_sum_d[30]), .QN(n1325) );
  DFFSSRX1_HVT conv2_sum_d_reg_29_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_d[29]), .CLK(clk), .Q(conv2_sum_d[29]), .QN(n1330) );
  DFFSSRX1_HVT conv2_sum_d_reg_28_ ( .D(1'b0), .SETB(n1434), .RSTB(
        n_conv2_sum_d[28]), .CLK(clk), .Q(conv2_sum_d[28]), .QN(n1327) );
  DFFSSRX1_HVT conv2_sum_d_reg_27_ ( .D(1'b0), .SETB(n1495), .RSTB(
        n_conv2_sum_d[27]), .CLK(clk), .Q(conv2_sum_d[27]), .QN(n1299) );
  DFFSSRX1_HVT conv2_sum_d_reg_26_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_d[26]), .CLK(clk), .Q(conv2_sum_d[26]), .QN(n1304) );
  DFFSSRX1_HVT conv2_sum_d_reg_25_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_d[25]), .CLK(clk), .Q(conv2_sum_d[25]), .QN(n1314) );
  DFFSSRX1_HVT conv2_sum_d_reg_24_ ( .D(1'b0), .SETB(n1445), .RSTB(
        n_conv2_sum_d[24]), .CLK(clk), .Q(conv2_sum_d[24]), .QN(n1311) );
  DFFSSRX1_HVT conv2_sum_d_reg_23_ ( .D(1'b0), .SETB(n1495), .RSTB(
        n_conv2_sum_d[23]), .CLK(clk), .Q(conv2_sum_d[23]), .QN(n1297) );
  DFFSSRX1_HVT conv2_sum_d_reg_22_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_d[22]), .CLK(clk), .Q(conv2_sum_d[22]), .QN(n1309) );
  DFFSSRX1_HVT conv2_sum_d_reg_21_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_d[21]), .CLK(clk), .Q(conv2_sum_d[21]), .QN(n1313) );
  DFFSSRX1_HVT conv2_sum_d_reg_20_ ( .D(1'b0), .SETB(n1434), .RSTB(
        n_conv2_sum_d[20]), .CLK(clk), .Q(conv2_sum_d[20]), .QN(n1310) );
  DFFSSRX1_HVT conv2_sum_d_reg_19_ ( .D(1'b0), .SETB(n1495), .RSTB(
        n_conv2_sum_d[19]), .CLK(clk), .Q(conv2_sum_d[19]), .QN(n1300) );
  DFFSSRX1_HVT conv2_sum_d_reg_18_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_d[18]), .CLK(clk), .Q(conv2_sum_d[18]), .QN(n1306) );
  DFFSSRX1_HVT conv2_sum_d_reg_17_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_d[17]), .CLK(clk), .Q(conv2_sum_d[17]), .QN(n1321) );
  DFFSSRX1_HVT conv2_sum_d_reg_16_ ( .D(1'b0), .SETB(n1445), .RSTB(
        n_conv2_sum_d[16]), .CLK(clk), .Q(conv2_sum_d[16]), .QN(n1884) );
  DFFSSRX1_HVT conv2_sum_d_reg_15_ ( .D(1'b0), .SETB(n1495), .RSTB(
        n_conv2_sum_d[15]), .CLK(clk), .Q(conv2_sum_d[15]), .QN(n1302) );
  DFFSSRX1_HVT conv2_sum_d_reg_14_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_d[14]), .CLK(clk), .Q(conv2_sum_d[14]), .QN(n1317) );
  DFFSSRX1_HVT conv2_sum_d_reg_13_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_d[13]), .CLK(clk), .Q(conv2_sum_d[13]), .QN(n1320) );
  DFFSSRX1_HVT conv2_sum_d_reg_12_ ( .D(1'b0), .SETB(n1434), .RSTB(
        n_conv2_sum_d[12]), .CLK(clk), .Q(conv2_sum_d[12]), .QN(n1289) );
  DFFSSRX1_HVT conv2_sum_d_reg_11_ ( .D(1'b0), .SETB(n1495), .RSTB(
        n_conv2_sum_d[11]), .CLK(clk), .Q(conv2_sum_d[11]), .QN(n1986) );
  DFFSSRX1_HVT conv2_sum_d_reg_10_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_d[10]), .CLK(clk), .Q(conv2_sum_d[10]), .QN(n1288) );
  DFFSSRX1_HVT conv2_sum_d_reg_8_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_d[8]), .CLK(clk), .Q(conv2_sum_d[8]), .QN(n1856) );
  DFFSSRX1_HVT conv2_sum_d_reg_7_ ( .D(1'b0), .SETB(n1445), .RSTB(
        n_conv2_sum_d[7]), .CLK(clk), .Q(conv2_sum_d[7]), .QN(n1279) );
  DFFSSRX1_HVT conv2_sum_d_reg_6_ ( .D(1'b0), .SETB(n1495), .RSTB(
        n_conv2_sum_d[6]), .CLK(clk), .Q(conv2_sum_d[6]), .QN(n1284) );
  DFFSSRX1_HVT conv2_sum_d_reg_5_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_d[5]), .CLK(clk), .Q(conv2_sum_d[5]), .QN(n1280) );
  DFFSSRX1_HVT conv2_sum_d_reg_4_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_d[4]), .CLK(clk), .Q(conv2_sum_d[4]), .QN(n1283) );
  DFFSSRX1_HVT conv2_sum_d_reg_3_ ( .D(1'b0), .SETB(n1434), .RSTB(
        n_conv2_sum_d[3]), .CLK(clk), .Q(conv2_sum_d[3]), .QN(n1987) );
  DFFSSRX1_HVT conv2_sum_d_reg_2_ ( .D(1'b0), .SETB(n1495), .RSTB(
        n_conv2_sum_d[2]), .CLK(clk), .Q(conv2_sum_d[2]), .QN(n1282) );
  DFFSSRX1_HVT conv2_sum_d_reg_0_ ( .D(1'b0), .SETB(n1445), .RSTB(
        n_conv2_sum_d[0]), .CLK(clk), .Q(conv2_sum_d[0]), .QN(n1294) );
  DFFSSRX1_HVT conv2_sum_a_reg_31_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_a[31]), .CLK(clk), .Q(conv2_sum_a[31]), .QN(n1323) );
  DFFSSRX1_HVT conv2_sum_a_reg_30_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_a[30]), .CLK(clk), .Q(conv2_sum_a[30]), .QN(n1912) );
  DFFSSRX1_HVT conv2_sum_a_reg_29_ ( .D(1'b0), .SETB(n1445), .RSTB(
        n_conv2_sum_a[29]), .CLK(clk), .Q(conv2_sum_a[29]), .QN(n1916) );
  DFFSSRX1_HVT conv2_sum_a_reg_28_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_a[28]), .CLK(clk), .Q(conv2_sum_a[28]), .QN(n1890) );
  DFFSSRX1_HVT conv2_sum_a_reg_27_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_a[27]), .CLK(clk), .QN(n1882) );
  DFFSSRX1_HVT conv2_sum_a_reg_26_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_a[26]), .CLK(clk), .Q(conv2_sum_a[26]), .QN(n1889) );
  DFFSSRX1_HVT conv2_sum_a_reg_25_ ( .D(1'b0), .SETB(n1434), .RSTB(
        n_conv2_sum_a[25]), .CLK(clk), .Q(conv2_sum_a[25]), .QN(n1903) );
  DFFSSRX1_HVT conv2_sum_a_reg_24_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_a[24]), .CLK(clk), .Q(conv2_sum_a[24]), .QN(n1888) );
  DFFSSRX1_HVT conv2_sum_a_reg_23_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_a[23]), .CLK(clk), .Q(conv2_sum_a[23]), .QN(n1902) );
  DFFSSRX1_HVT conv2_sum_a_reg_22_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_a[22]), .CLK(clk), .Q(conv2_sum_a[22]), .QN(n1887) );
  DFFSSRX1_HVT conv2_sum_a_reg_21_ ( .D(1'b0), .SETB(n1445), .RSTB(
        n_conv2_sum_a[21]), .CLK(clk), .Q(conv2_sum_a[21]), .QN(n1901) );
  DFFSSRX1_HVT conv2_sum_a_reg_20_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_a[20]), .CLK(clk), .Q(conv2_sum_a[20]), .QN(n1886) );
  DFFSSRX1_HVT conv2_sum_a_reg_19_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_a[19]), .CLK(clk), .Q(conv2_sum_a[19]), .QN(n1900) );
  DFFSSRX1_HVT conv2_sum_a_reg_18_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_a[18]), .CLK(clk), .Q(conv2_sum_a[18]), .QN(n1885) );
  DFFSSRX1_HVT conv2_sum_a_reg_17_ ( .D(1'b0), .SETB(n1434), .RSTB(
        n_conv2_sum_a[17]), .CLK(clk), .Q(conv2_sum_a[17]), .QN(n1899) );
  DFFSSRX1_HVT conv2_sum_a_reg_16_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_a[16]), .CLK(clk), .Q(conv2_sum_a[16]), .QN(n1318) );
  DFFSSRX1_HVT conv2_sum_a_reg_15_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_a[15]), .CLK(clk), .Q(conv2_sum_a[15]), .QN(n1898) );
  DFFSSRX1_HVT conv2_sum_a_reg_14_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_a[14]), .CLK(clk), .Q(conv2_sum_a[14]), .QN(n1978) );
  DFFSSRX1_HVT conv2_sum_a_reg_13_ ( .D(1'b0), .SETB(n1445), .RSTB(
        n_conv2_sum_a[13]), .CLK(clk), .Q(conv2_sum_a[13]), .QN(n1879) );
  DFFSSRX1_HVT conv2_sum_a_reg_12_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_a[12]), .CLK(clk), .Q(conv2_sum_a[12]), .QN(n1864) );
  DFFSSRX1_HVT conv2_sum_a_reg_11_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_a[11]), .CLK(clk), .Q(conv2_sum_a[11]), .QN(n1973) );
  DFFSSRX1_HVT conv2_sum_a_reg_10_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_a[10]), .CLK(clk), .Q(conv2_sum_a[10]), .QN(n1849) );
  DFFSSRX1_HVT conv2_sum_a_reg_8_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_a[8]), .CLK(clk), .Q(conv2_sum_a[8]), .QN(n1285) );
  DFFSSRX1_HVT conv2_sum_a_reg_7_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_a[7]), .CLK(clk), .Q(conv2_sum_a[7]), .QN(n1853) );
  DFFSSRX1_HVT conv2_sum_a_reg_6_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_a[6]), .CLK(clk), .Q(conv2_sum_a[6]), .QN(n1861) );
  DFFSSRX1_HVT conv2_sum_a_reg_5_ ( .D(1'b0), .SETB(n1445), .RSTB(
        n_conv2_sum_a[5]), .CLK(clk), .QN(n1852) );
  DFFSSRX1_HVT conv2_sum_a_reg_4_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_a[4]), .CLK(clk), .Q(conv2_sum_a[4]), .QN(n1863) );
  DFFSSRX1_HVT conv2_sum_a_reg_3_ ( .D(1'b0), .SETB(n1434), .RSTB(
        n_conv2_sum_a[3]), .CLK(clk), .Q(conv2_sum_a[3]), .QN(n1872) );
  DFFSSRX1_HVT conv2_sum_a_reg_2_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_a[2]), .CLK(clk), .Q(conv2_sum_a[2]), .QN(n1867) );
  DFFSSRX1_HVT conv2_sum_a_reg_1_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_a[1]), .CLK(clk), .Q(conv2_sum_a[1]), .QN(n1975) );
  DFFSSRX1_HVT conv2_sum_a_reg_0_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_a[0]), .CLK(clk), .Q(conv2_sum_a[0]), .QN(n1869) );
  DFFSSRX1_HVT conv2_sum_b_reg_31_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_b[31]), .CLK(clk), .Q(conv2_sum_b[31]), .QN(n1914) );
  DFFSSRX1_HVT conv2_sum_b_reg_30_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_b[30]), .CLK(clk), .Q(conv2_sum_b[30]), .QN(n1326) );
  DFFSSRX1_HVT conv2_sum_b_reg_29_ ( .D(1'b0), .SETB(n1445), .RSTB(
        n_conv2_sum_b[29]), .CLK(clk), .Q(conv2_sum_b[29]), .QN(n1329) );
  DFFSSRX1_HVT conv2_sum_b_reg_28_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_b[28]), .CLK(clk), .Q(conv2_sum_b[28]), .QN(n1328) );
  DFFSSRX1_HVT conv2_sum_b_reg_27_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_b[27]), .CLK(clk), .Q(conv2_sum_b[27]), .QN(n1881) );
  DFFSSRX1_HVT conv2_sum_b_reg_26_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_b[26]), .CLK(clk), .Q(conv2_sum_b[26]), .QN(n1305) );
  DFFSSRX1_HVT conv2_sum_b_reg_25_ ( .D(1'b0), .SETB(n1434), .RSTB(
        n_conv2_sum_b[25]), .CLK(clk), .Q(conv2_sum_b[25]), .QN(n1307) );
  DFFSSRX1_HVT conv2_sum_b_reg_24_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_b[24]), .CLK(clk), .Q(conv2_sum_b[24]), .QN(n1296) );
  DFFSSRX1_HVT conv2_sum_b_reg_23_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_b[23]), .CLK(clk), .Q(conv2_sum_b[23]), .QN(n1298) );
  DFFSSRX1_HVT conv2_sum_b_reg_22_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_b[22]), .CLK(clk), .Q(conv2_sum_b[22]), .QN(n1308) );
  DFFSSRX1_HVT conv2_sum_b_reg_21_ ( .D(1'b0), .SETB(n1445), .RSTB(
        n_conv2_sum_b[21]), .CLK(clk), .Q(conv2_sum_b[21]), .QN(n1315) );
  DFFSSRX1_HVT conv2_sum_b_reg_20_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_b[20]), .CLK(clk), .Q(conv2_sum_b[20]), .QN(n1312) );
  DFFSSRX1_HVT conv2_sum_b_reg_19_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_b[19]), .CLK(clk), .Q(conv2_sum_b[19]), .QN(n1303) );
  DFFSSRX1_HVT conv2_sum_b_reg_18_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_b[18]), .CLK(clk), .Q(conv2_sum_b[18]), .QN(n1316) );
  DFFSSRX1_HVT conv2_sum_b_reg_17_ ( .D(1'b0), .SETB(n1434), .RSTB(
        n_conv2_sum_b[17]), .CLK(clk), .Q(conv2_sum_b[17]), .QN(n1322) );
  DFFSSRX1_HVT conv2_sum_b_reg_16_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_b[16]), .CLK(clk), .Q(conv2_sum_b[16]), .QN(n1883) );
  DFFSSRX1_HVT conv2_sum_b_reg_15_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_b[15]), .CLK(clk), .Q(conv2_sum_b[15]), .QN(n1301) );
  DFFSSRX1_HVT conv2_sum_b_reg_14_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_b[14]), .CLK(clk), .Q(conv2_sum_b[14]), .QN(n1977) );
  DFFSSRX1_HVT conv2_sum_b_reg_13_ ( .D(1'b0), .SETB(n1445), .RSTB(
        n_conv2_sum_b[13]), .CLK(clk), .Q(conv2_sum_b[13]), .QN(n1880) );
  DFFSSRX1_HVT conv2_sum_b_reg_12_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_b[12]), .CLK(clk), .Q(conv2_sum_b[12]), .QN(n1857) );
  DFFSSRX1_HVT conv2_sum_b_reg_11_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_b[11]), .CLK(clk), .Q(conv2_sum_b[11]), .QN(n1524) );
  DFFSSRX1_HVT conv2_sum_b_reg_10_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_b[10]), .CLK(clk), .Q(conv2_sum_b[10]), .QN(n1850) );
  DFFSSRX1_HVT conv2_sum_b_reg_9_ ( .D(1'b0), .SETB(n1434), .RSTB(
        n_conv2_sum_b[9]), .CLK(clk), .Q(conv2_sum_b[9]), .QN(n1984) );
  DFFSSRX1_HVT conv2_sum_b_reg_8_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_b[8]), .CLK(clk), .Q(conv2_sum_b[8]), .QN(n1858) );
  DFFSSRX1_HVT conv2_sum_b_reg_7_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_b[7]), .CLK(clk), .Q(conv2_sum_b[7]), .QN(n1278) );
  DFFSSRX1_HVT conv2_sum_b_reg_6_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_b[6]), .CLK(clk), .Q(conv2_sum_b[6]), .QN(n1281) );
  DFFSSRX1_HVT conv2_sum_b_reg_5_ ( .D(1'b0), .SETB(n1445), .RSTB(
        n_conv2_sum_b[5]), .CLK(clk), .Q(conv2_sum_b[5]), .QN(n1851) );
  DFFSSRX1_HVT conv2_sum_b_reg_4_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_b[4]), .CLK(clk), .Q(conv2_sum_b[4]), .QN(n1287) );
  DFFSSRX1_HVT conv2_sum_b_reg_3_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_b[3]), .CLK(clk), .Q(conv2_sum_b[3]), .QN(n1981) );
  DFFSSRX1_HVT conv2_sum_b_reg_2_ ( .D(1'b0), .SETB(n1494), .RSTB(
        n_conv2_sum_b[2]), .CLK(clk), .Q(conv2_sum_b[2]), .QN(n1866) );
  DFFSSRX1_HVT conv2_sum_b_reg_1_ ( .D(1'b0), .SETB(n1434), .RSTB(
        n_conv2_sum_b[1]), .CLK(clk), .Q(conv2_sum_b[1]), .QN(n1989) );
  DFFSSRX1_HVT conv2_sum_b_reg_0_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_b[0]), .CLK(clk), .Q(conv2_sum_b[0]), .QN(n1293) );
  DFFSSRX1_HVT conv2_sum_d_reg_9_ ( .D(1'b0), .SETB(n1492), .RSTB(
        n_conv2_sum_d[9]), .CLK(clk), .Q(conv2_sum_d[9]), .QN(n1983) );
  DFFSSRX1_HVT conv2_sum_d_reg_1_ ( .D(1'b0), .SETB(n1493), .RSTB(
        n_conv2_sum_d[1]), .CLK(clk), .Q(conv2_sum_d[1]) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U200 ( .A1(n1381), .A2(
        DP_OP_425J2_127_3477_n332), .Y(DP_OP_425J2_127_3477_n182) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U325 ( .A1(DP_OP_425J2_127_3477_n5), .A2(
        DP_OP_425J2_127_3477_n267), .A3(DP_OP_425J2_127_3477_n268), .Y(
        DP_OP_425J2_127_3477_n266) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U173 ( .A1(DP_OP_425J2_127_3477_n174), .A2(
        DP_OP_425J2_127_3477_n166), .A3(DP_OP_425J2_127_3477_n167), .Y(
        DP_OP_425J2_127_3477_n165) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U83 ( .A1(DP_OP_425J2_127_3477_n105), .A2(
        DP_OP_425J2_127_3477_n97), .A3(DP_OP_425J2_127_3477_n98), .Y(
        DP_OP_425J2_127_3477_n96) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U123 ( .A1(DP_OP_425J2_127_3477_n136), .A2(
        DP_OP_425J2_127_3477_n128), .A3(DP_OP_425J2_127_3477_n129), .Y(
        DP_OP_425J2_127_3477_n127) );
  XNOR2X1_HVT DP_OP_425J2_127_3477_U787 ( .A1(DP_OP_425J2_127_3477_n2502), 
        .A2(DP_OP_425J2_127_3477_n3029), .Y(DP_OP_425J2_127_3477_n1211) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2291 ( .A1(DP_OP_425J2_127_3477_n3058), 
        .A2(n690), .Y(DP_OP_425J2_127_3477_n3050) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2290 ( .A1(DP_OP_425J2_127_3477_n3057), 
        .A2(n34), .Y(DP_OP_425J2_127_3477_n3049) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2289 ( .A1(DP_OP_425J2_127_3477_n3056), .A2(
        n34), .Y(DP_OP_425J2_127_3477_n3048) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2282 ( .A1(DP_OP_425J2_127_3477_n3057), 
        .A2(DP_OP_425J2_127_3477_n3066), .Y(DP_OP_425J2_127_3477_n3041) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2273 ( .A1(DP_OP_425J2_127_3477_n3056), .A2(
        DP_OP_425J2_127_3477_n3065), .Y(DP_OP_425J2_127_3477_n3032) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2272 ( .A1(DP_OP_425J2_127_3477_n3063), .A2(
        n215), .Y(DP_OP_425J2_127_3477_n1728) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2271 ( .A1(DP_OP_425J2_127_3477_n3062), .A2(
        n215), .Y(DP_OP_425J2_127_3477_n3031) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2270 ( .A1(DP_OP_425J2_127_3477_n3061), .A2(
        n213), .Y(DP_OP_425J2_127_3477_n3030) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2269 ( .A1(DP_OP_425J2_127_3477_n3060), .A2(
        n215), .Y(DP_OP_425J2_127_3477_n3029) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2268 ( .A1(DP_OP_425J2_127_3477_n3059), .A2(
        n215), .Y(DP_OP_425J2_127_3477_n3028) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2267 ( .A1(DP_OP_425J2_127_3477_n3058), .A2(
        n213), .Y(DP_OP_425J2_127_3477_n820) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2266 ( .A1(DP_OP_425J2_127_3477_n3057), .A2(
        n213), .Y(DP_OP_425J2_127_3477_n3027) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2265 ( .A1(DP_OP_425J2_127_3477_n3056), 
        .A2(n213), .Y(DP_OP_425J2_127_3477_n3026) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2245 ( .A1(DP_OP_424J2_126_3477_n2002), .A2(
        DP_OP_425J2_127_3477_n3025), .Y(DP_OP_425J2_127_3477_n3006) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2238 ( .A1(DP_OP_424J2_126_3477_n2003), 
        .A2(n704), .Y(DP_OP_425J2_127_3477_n2999) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2237 ( .A1(DP_OP_424J2_126_3477_n2002), .A2(
        n698), .Y(DP_OP_425J2_127_3477_n2998) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2226 ( .A1(DP_OP_425J2_127_3477_n3019), .A2(
        DP_OP_423J2_125_3477_n3022), .Y(DP_OP_425J2_127_3477_n2987) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2201 ( .A1(DP_OP_425J2_127_3477_n2970), .A2(
        n677), .Y(DP_OP_425J2_127_3477_n2962) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2193 ( .A1(DP_OP_425J2_127_3477_n2970), .A2(
        DP_OP_424J2_126_3477_n2980), .Y(DP_OP_425J2_127_3477_n2954) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2184 ( .A1(DP_OP_425J2_127_3477_n2977), .A2(
        n663), .Y(DP_OP_425J2_127_3477_n2945) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2157 ( .A1(DP_OP_424J2_126_3477_n2090), .A2(
        n446), .Y(DP_OP_425J2_127_3477_n2918) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2140 ( .A1(DP_OP_425J2_127_3477_n2933), .A2(
        n35), .Y(DP_OP_425J2_127_3477_n2901) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2139 ( .A1(DP_OP_423J2_125_3477_n2008), .A2(
        n35), .Y(DP_OP_425J2_127_3477_n2900) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2138 ( .A1(DP_OP_423J2_125_3477_n2007), .A2(
        n35), .Y(DP_OP_425J2_127_3477_n2899) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2137 ( .A1(DP_OP_422J2_124_3477_n3060), .A2(
        n35), .Y(DP_OP_425J2_127_3477_n2898) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2136 ( .A1(DP_OP_423J2_125_3477_n2005), .A2(
        n35), .Y(DP_OP_425J2_127_3477_n2897) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2135 ( .A1(DP_OP_424J2_126_3477_n2092), .A2(
        n35), .Y(DP_OP_425J2_127_3477_n2896) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2134 ( .A1(DP_OP_423J2_125_3477_n2003), .A2(
        n35), .Y(DP_OP_425J2_127_3477_n2895) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2133 ( .A1(DP_OP_424J2_126_3477_n2090), 
        .A2(n603), .Y(DP_OP_425J2_127_3477_n2894) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2113 ( .A1(DP_OP_425J2_127_3477_n2882), .A2(
        DP_OP_425J2_127_3477_n2893), .Y(DP_OP_425J2_127_3477_n2874) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2098 ( .A1(DP_OP_425J2_127_3477_n2883), 
        .A2(DP_OP_424J2_126_3477_n2891), .Y(DP_OP_425J2_127_3477_n2859) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2097 ( .A1(DP_OP_425J2_127_3477_n2882), .A2(
        DP_OP_425J2_127_3477_n2891), .Y(DP_OP_425J2_127_3477_n2858) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2096 ( .A1(DP_OP_422J2_124_3477_n3021), .A2(
        DP_OP_422J2_124_3477_n2890), .Y(DP_OP_425J2_127_3477_n2857) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2095 ( .A1(DP_OP_425J2_127_3477_n2888), .A2(
        DP_OP_424J2_126_3477_n2890), .Y(DP_OP_425J2_127_3477_n2856) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2094 ( .A1(DP_OP_422J2_124_3477_n3019), .A2(
        DP_OP_422J2_124_3477_n2890), .Y(DP_OP_425J2_127_3477_n2855) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2093 ( .A1(DP_OP_425J2_127_3477_n2886), .A2(
        DP_OP_423J2_125_3477_n2890), .Y(DP_OP_425J2_127_3477_n2854) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2092 ( .A1(DP_OP_425J2_127_3477_n2885), .A2(
        DP_OP_423J2_125_3477_n2890), .Y(DP_OP_425J2_127_3477_n2853) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2091 ( .A1(DP_OP_424J2_126_3477_n2136), .A2(
        DP_OP_424J2_126_3477_n2890), .Y(DP_OP_425J2_127_3477_n2852) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2090 ( .A1(DP_OP_425J2_127_3477_n2883), .A2(
        DP_OP_423J2_125_3477_n2890), .Y(DP_OP_425J2_127_3477_n2851) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2089 ( .A1(DP_OP_425J2_127_3477_n2882), 
        .A2(DP_OP_424J2_126_3477_n2890), .Y(DP_OP_425J2_127_3477_n2850) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2070 ( .A1(DP_OP_425J2_127_3477_n2839), 
        .A2(DP_OP_423J2_125_3477_n2849), .Y(DP_OP_425J2_127_3477_n2831) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2062 ( .A1(DP_OP_425J2_127_3477_n2839), 
        .A2(DP_OP_425J2_127_3477_n2848), .Y(DP_OP_425J2_127_3477_n2823) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2061 ( .A1(DP_OP_423J2_125_3477_n2090), .A2(
        DP_OP_425J2_127_3477_n2848), .Y(DP_OP_425J2_127_3477_n2822) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2054 ( .A1(DP_OP_425J2_127_3477_n2839), 
        .A2(DP_OP_425J2_127_3477_n2847), .Y(DP_OP_425J2_127_3477_n2815) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2052 ( .A1(DP_OP_423J2_125_3477_n2097), .A2(
        DP_OP_425J2_127_3477_n2846), .Y(DP_OP_425J2_127_3477_n2813) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2051 ( .A1(DP_OP_423J2_125_3477_n2096), .A2(
        DP_OP_425J2_127_3477_n2846), .Y(DP_OP_425J2_127_3477_n2812) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2050 ( .A1(DP_OP_425J2_127_3477_n2843), .A2(
        DP_OP_425J2_127_3477_n2846), .Y(DP_OP_425J2_127_3477_n2811) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2049 ( .A1(DP_OP_423J2_125_3477_n2094), .A2(
        DP_OP_425J2_127_3477_n2846), .Y(DP_OP_425J2_127_3477_n2810) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2048 ( .A1(DP_OP_425J2_127_3477_n2841), .A2(
        DP_OP_425J2_127_3477_n2846), .Y(DP_OP_425J2_127_3477_n2809) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2047 ( .A1(DP_OP_425J2_127_3477_n2840), .A2(
        DP_OP_425J2_127_3477_n2846), .Y(DP_OP_425J2_127_3477_n2808) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2046 ( .A1(DP_OP_425J2_127_3477_n2839), .A2(
        DP_OP_425J2_127_3477_n2846), .Y(DP_OP_425J2_127_3477_n2807) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2045 ( .A1(DP_OP_423J2_125_3477_n2090), 
        .A2(DP_OP_425J2_127_3477_n2846), .Y(DP_OP_425J2_127_3477_n2806) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2026 ( .A1(DP_OP_423J2_125_3477_n2135), 
        .A2(DP_OP_423J2_125_3477_n2805), .Y(DP_OP_425J2_127_3477_n2787) );
  OR2X1_HVT DP_OP_425J2_127_3477_U2025 ( .A1(DP_OP_422J2_124_3477_n2926), .A2(
        DP_OP_423J2_125_3477_n2805), .Y(DP_OP_425J2_127_3477_n2786) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2022 ( .A1(DP_OP_425J2_127_3477_n2799), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_425J2_127_3477_n2783) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2021 ( .A1(DP_OP_425J2_127_3477_n2798), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_425J2_127_3477_n2782) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2020 ( .A1(DP_OP_425J2_127_3477_n2797), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_425J2_127_3477_n2781) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2013 ( .A1(DP_OP_425J2_127_3477_n2798), 
        .A2(n1444), .Y(DP_OP_425J2_127_3477_n2774) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2012 ( .A1(DP_OP_425J2_127_3477_n2797), 
        .A2(DP_OP_422J2_124_3477_n2803), .Y(DP_OP_425J2_127_3477_n2773) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1982 ( .A1(DP_OP_424J2_126_3477_n2267), 
        .A2(n66), .Y(DP_OP_425J2_127_3477_n2743) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1981 ( .A1(DP_OP_423J2_125_3477_n2178), .A2(
        n66), .Y(DP_OP_425J2_127_3477_n2742) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1974 ( .A1(DP_OP_422J2_124_3477_n2883), 
        .A2(DP_OP_425J2_127_3477_n2760), .Y(DP_OP_425J2_127_3477_n2735) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1973 ( .A1(DP_OP_423J2_125_3477_n2178), .A2(
        DP_OP_425J2_127_3477_n2760), .Y(DP_OP_425J2_127_3477_n2734) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1964 ( .A1(DP_OP_422J2_124_3477_n2889), .A2(
        DP_OP_422J2_124_3477_n2758), .Y(DP_OP_425J2_127_3477_n2725) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1963 ( .A1(DP_OP_425J2_127_3477_n2756), .A2(
        DP_OP_424J2_126_3477_n2758), .Y(DP_OP_425J2_127_3477_n2724) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1961 ( .A1(DP_OP_425J2_127_3477_n2754), .A2(
        DP_OP_423J2_125_3477_n2758), .Y(DP_OP_425J2_127_3477_n2722) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1937 ( .A1(DP_OP_423J2_125_3477_n2222), .A2(
        n597), .Y(DP_OP_425J2_127_3477_n2698) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1930 ( .A1(DP_OP_424J2_126_3477_n2311), 
        .A2(n1342), .Y(DP_OP_425J2_127_3477_n2691) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1929 ( .A1(DP_OP_423J2_125_3477_n2222), .A2(
        n1342), .Y(DP_OP_425J2_127_3477_n2690) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1923 ( .A1(DP_OP_425J2_127_3477_n2708), 
        .A2(n1440), .Y(DP_OP_425J2_127_3477_n2684) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1920 ( .A1(DP_OP_424J2_126_3477_n2317), .A2(
        DP_OP_425J2_127_3477_n2714), .Y(DP_OP_425J2_127_3477_n2681) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1919 ( .A1(DP_OP_425J2_127_3477_n2712), .A2(
        DP_OP_425J2_127_3477_n2714), .Y(DP_OP_425J2_127_3477_n2680) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1918 ( .A1(DP_OP_423J2_125_3477_n2227), .A2(
        DP_OP_425J2_127_3477_n2714), .Y(DP_OP_425J2_127_3477_n2679) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1916 ( .A1(DP_OP_422J2_124_3477_n2841), .A2(
        DP_OP_425J2_127_3477_n2714), .Y(DP_OP_425J2_127_3477_n2677) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1915 ( .A1(DP_OP_425J2_127_3477_n2708), .A2(
        DP_OP_425J2_127_3477_n2714), .Y(DP_OP_425J2_127_3477_n2676) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1914 ( .A1(DP_OP_424J2_126_3477_n2311), .A2(
        DP_OP_425J2_127_3477_n2714), .Y(DP_OP_425J2_127_3477_n2675) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1913 ( .A1(DP_OP_423J2_125_3477_n2222), 
        .A2(DP_OP_425J2_127_3477_n2714), .Y(DP_OP_425J2_127_3477_n2674) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1893 ( .A1(DP_OP_424J2_126_3477_n2354), .A2(
        DP_OP_425J2_127_3477_n2673), .Y(DP_OP_425J2_127_3477_n2654) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1885 ( .A1(DP_OP_424J2_126_3477_n2354), .A2(
        n279), .Y(DP_OP_425J2_127_3477_n2646) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1884 ( .A1(DP_OP_423J2_125_3477_n2273), 
        .A2(DP_OP_424J2_126_3477_n2671), .Y(DP_OP_425J2_127_3477_n2645) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1882 ( .A1(DP_OP_422J2_124_3477_n2799), 
        .A2(n1400), .Y(DP_OP_425J2_127_3477_n2643) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1873 ( .A1(DP_OP_424J2_126_3477_n2358), .A2(
        DP_OP_422J2_124_3477_n2670), .Y(DP_OP_425J2_127_3477_n2634) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1872 ( .A1(DP_OP_423J2_125_3477_n2269), .A2(
        DP_OP_422J2_124_3477_n2670), .Y(DP_OP_425J2_127_3477_n2633) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1871 ( .A1(DP_OP_422J2_124_3477_n2796), .A2(
        n86), .Y(DP_OP_425J2_127_3477_n2632) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1869 ( .A1(DP_OP_422J2_124_3477_n2794), 
        .A2(n86), .Y(DP_OP_425J2_127_3477_n2630) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1849 ( .A1(DP_OP_423J2_125_3477_n2310), .A2(
        DP_OP_423J2_125_3477_n2629), .Y(DP_OP_425J2_127_3477_n2610) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1833 ( .A1(DP_OP_423J2_125_3477_n2310), .A2(
        DP_OP_424J2_126_3477_n2627), .Y(DP_OP_425J2_127_3477_n2594) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1798 ( .A1(DP_OP_424J2_126_3477_n2443), 
        .A2(n186), .Y(DP_OP_425J2_127_3477_n2559) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1797 ( .A1(DP_OP_425J2_127_3477_n2574), .A2(
        n186), .Y(DP_OP_425J2_127_3477_n2558) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1788 ( .A1(DP_OP_425J2_127_3477_n2581), .A2(
        DP_OP_425J2_127_3477_n2582), .Y(DP_OP_425J2_127_3477_n2549) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1787 ( .A1(DP_OP_425J2_127_3477_n2580), .A2(
        DP_OP_425J2_127_3477_n2582), .Y(DP_OP_425J2_127_3477_n2548) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1786 ( .A1(DP_OP_425J2_127_3477_n2579), .A2(
        DP_OP_425J2_127_3477_n2582), .Y(DP_OP_425J2_127_3477_n2547) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1785 ( .A1(DP_OP_425J2_127_3477_n2578), .A2(
        DP_OP_425J2_127_3477_n2582), .Y(DP_OP_425J2_127_3477_n2546) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1784 ( .A1(DP_OP_425J2_127_3477_n2577), .A2(
        DP_OP_425J2_127_3477_n2582), .Y(DP_OP_425J2_127_3477_n2545) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1783 ( .A1(DP_OP_425J2_127_3477_n2576), .A2(
        DP_OP_425J2_127_3477_n2582), .Y(DP_OP_425J2_127_3477_n2544) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1782 ( .A1(DP_OP_424J2_126_3477_n2443), .A2(
        DP_OP_425J2_127_3477_n2582), .Y(DP_OP_425J2_127_3477_n2543) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1781 ( .A1(DP_OP_425J2_127_3477_n2574), 
        .A2(DP_OP_425J2_127_3477_n2582), .Y(DP_OP_425J2_127_3477_n2542) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1746 ( .A1(DP_OP_423J2_125_3477_n2399), 
        .A2(n772), .Y(DP_OP_425J2_127_3477_n2507) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1745 ( .A1(DP_OP_422J2_124_3477_n2662), .A2(
        n772), .Y(DP_OP_425J2_127_3477_n2506) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1743 ( .A1(DP_OP_425J2_127_3477_n2536), .A2(
        n1336), .Y(DP_OP_425J2_127_3477_n2504) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1742 ( .A1(DP_OP_422J2_124_3477_n2667), .A2(
        n1362), .Y(DP_OP_425J2_127_3477_n2503) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1741 ( .A1(DP_OP_425J2_127_3477_n2534), .A2(
        DP_OP_423J2_125_3477_n2538), .Y(DP_OP_425J2_127_3477_n2502) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1740 ( .A1(DP_OP_423J2_125_3477_n2401), .A2(
        n1336), .Y(DP_OP_425J2_127_3477_n2501) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1739 ( .A1(DP_OP_423J2_125_3477_n2400), .A2(
        n1335), .Y(DP_OP_425J2_127_3477_n2500) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1738 ( .A1(DP_OP_423J2_125_3477_n2399), .A2(
        n1337), .Y(DP_OP_425J2_127_3477_n2499) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1737 ( .A1(DP_OP_424J2_126_3477_n2486), 
        .A2(n1335), .Y(DP_OP_425J2_127_3477_n2498) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1718 ( .A1(DP_OP_424J2_126_3477_n2575), 
        .A2(DP_OP_422J2_124_3477_n2497), .Y(DP_OP_425J2_127_3477_n2479) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1717 ( .A1(DP_OP_424J2_126_3477_n2574), .A2(
        DP_OP_424J2_126_3477_n2497), .Y(DP_OP_425J2_127_3477_n2478) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1709 ( .A1(DP_OP_424J2_126_3477_n2574), .A2(
        n1491), .Y(DP_OP_425J2_127_3477_n2470) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1674 ( .A1(DP_OP_424J2_126_3477_n2619), 
        .A2(DP_OP_425J2_127_3477_n2453), .Y(DP_OP_425J2_127_3477_n2435) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1673 ( .A1(DP_OP_423J2_125_3477_n2706), .A2(
        DP_OP_425J2_127_3477_n2453), .Y(DP_OP_425J2_127_3477_n2434) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1665 ( .A1(DP_OP_423J2_125_3477_n2706), .A2(
        DP_OP_423J2_125_3477_n2452), .Y(DP_OP_425J2_127_3477_n2426) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1657 ( .A1(DP_OP_423J2_125_3477_n2706), .A2(
        n789), .Y(DP_OP_425J2_127_3477_n2418) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1631 ( .A1(DP_OP_425J2_127_3477_n2400), 
        .A2(DP_OP_423J2_125_3477_n2409), .Y(DP_OP_425J2_127_3477_n2392) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1630 ( .A1(DP_OP_423J2_125_3477_n2751), 
        .A2(DP_OP_425J2_127_3477_n2409), .Y(DP_OP_425J2_127_3477_n2391) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1614 ( .A1(DP_OP_422J2_124_3477_n2267), 
        .A2(n793), .Y(DP_OP_425J2_127_3477_n2375) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1613 ( .A1(DP_OP_423J2_125_3477_n2750), .A2(
        n799), .Y(DP_OP_425J2_127_3477_n2374) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1612 ( .A1(DP_OP_424J2_126_3477_n2669), .A2(
        n1426), .Y(DP_OP_425J2_127_3477_n2373) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1610 ( .A1(DP_OP_425J2_127_3477_n2403), .A2(
        n1426), .Y(DP_OP_425J2_127_3477_n2371) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1586 ( .A1(DP_OP_423J2_125_3477_n2795), 
        .A2(DP_OP_425J2_127_3477_n2365), .Y(DP_OP_425J2_127_3477_n2347) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1577 ( .A1(DP_OP_423J2_125_3477_n2794), .A2(
        n1386), .Y(DP_OP_425J2_127_3477_n2338) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1567 ( .A1(DP_OP_424J2_126_3477_n2712), .A2(
        DP_OP_423J2_125_3477_n2362), .Y(DP_OP_425J2_127_3477_n2328) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1565 ( .A1(DP_OP_425J2_127_3477_n2358), .A2(
        DP_OP_423J2_125_3477_n2362), .Y(DP_OP_425J2_127_3477_n2326) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1562 ( .A1(DP_OP_423J2_125_3477_n2795), .A2(
        DP_OP_423J2_125_3477_n2362), .Y(DP_OP_425J2_127_3477_n2323) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1542 ( .A1(DP_OP_425J2_127_3477_n2311), 
        .A2(DP_OP_425J2_127_3477_n2321), .Y(DP_OP_425J2_127_3477_n2303) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1541 ( .A1(DP_OP_425J2_127_3477_n2310), .A2(
        DP_OP_425J2_127_3477_n2321), .Y(DP_OP_425J2_127_3477_n2302) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1533 ( .A1(DP_OP_425J2_127_3477_n2310), .A2(
        DP_OP_425J2_127_3477_n2320), .Y(DP_OP_425J2_127_3477_n2294) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1526 ( .A1(DP_OP_425J2_127_3477_n2311), 
        .A2(DP_OP_425J2_127_3477_n2319), .Y(DP_OP_425J2_127_3477_n2287) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1525 ( .A1(DP_OP_425J2_127_3477_n2310), .A2(
        n317), .Y(DP_OP_425J2_127_3477_n2286) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1524 ( .A1(DP_OP_423J2_125_3477_n2845), .A2(
        DP_OP_424J2_126_3477_n2318), .Y(DP_OP_425J2_127_3477_n2285) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1523 ( .A1(DP_OP_423J2_125_3477_n2844), .A2(
        DP_OP_423J2_125_3477_n2318), .Y(DP_OP_425J2_127_3477_n2284) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1522 ( .A1(DP_OP_423J2_125_3477_n2843), .A2(
        DP_OP_422J2_124_3477_n2318), .Y(DP_OP_425J2_127_3477_n2283) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1521 ( .A1(DP_OP_423J2_125_3477_n2842), .A2(
        DP_OP_422J2_124_3477_n2318), .Y(DP_OP_425J2_127_3477_n2282) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1520 ( .A1(DP_OP_423J2_125_3477_n2841), .A2(
        DP_OP_422J2_124_3477_n2318), .Y(DP_OP_425J2_127_3477_n2281) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1519 ( .A1(DP_OP_425J2_127_3477_n2312), .A2(
        DP_OP_424J2_126_3477_n2318), .Y(DP_OP_425J2_127_3477_n2280) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1518 ( .A1(DP_OP_425J2_127_3477_n2311), .A2(
        DP_OP_423J2_125_3477_n2318), .Y(DP_OP_425J2_127_3477_n2279) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1517 ( .A1(DP_OP_425J2_127_3477_n2310), 
        .A2(DP_OP_424J2_126_3477_n2318), .Y(DP_OP_425J2_127_3477_n2278) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1499 ( .A1(DP_OP_425J2_127_3477_n2268), 
        .A2(DP_OP_423J2_125_3477_n2277), .Y(DP_OP_425J2_127_3477_n2260) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1497 ( .A1(DP_OP_424J2_126_3477_n2794), .A2(
        DP_OP_422J2_124_3477_n2277), .Y(DP_OP_425J2_127_3477_n2258) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1489 ( .A1(DP_OP_422J2_124_3477_n2134), .A2(
        DP_OP_424J2_126_3477_n2276), .Y(DP_OP_425J2_127_3477_n2250) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1481 ( .A1(DP_OP_424J2_126_3477_n2794), .A2(
        DP_OP_422J2_124_3477_n2275), .Y(DP_OP_425J2_127_3477_n2242) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1480 ( .A1(DP_OP_423J2_125_3477_n2889), .A2(
        n1370), .Y(DP_OP_425J2_127_3477_n2241) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1479 ( .A1(DP_OP_425J2_127_3477_n2272), .A2(
        n1338), .Y(DP_OP_425J2_127_3477_n2240) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1478 ( .A1(DP_OP_424J2_126_3477_n2799), .A2(
        n1370), .Y(DP_OP_425J2_127_3477_n2239) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1477 ( .A1(DP_OP_423J2_125_3477_n2886), .A2(
        n1338), .Y(DP_OP_425J2_127_3477_n2238) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1476 ( .A1(DP_OP_425J2_127_3477_n2269), .A2(
        n1370), .Y(DP_OP_425J2_127_3477_n2237) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1475 ( .A1(DP_OP_425J2_127_3477_n2268), .A2(
        n1370), .Y(DP_OP_425J2_127_3477_n2236) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1474 ( .A1(DP_OP_424J2_126_3477_n2795), .A2(
        n1338), .Y(DP_OP_425J2_127_3477_n2235) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1473 ( .A1(DP_OP_424J2_126_3477_n2794), 
        .A2(n1370), .Y(DP_OP_425J2_127_3477_n2234) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1445 ( .A1(DP_OP_422J2_124_3477_n2090), .A2(
        n365), .Y(DP_OP_425J2_127_3477_n2206) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1436 ( .A1(DP_OP_424J2_126_3477_n2845), .A2(
        DP_OP_425J2_127_3477_n2230), .Y(DP_OP_425J2_127_3477_n2197) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1434 ( .A1(DP_OP_423J2_125_3477_n2931), .A2(
        DP_OP_425J2_127_3477_n2230), .Y(DP_OP_425J2_127_3477_n2195) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1433 ( .A1(DP_OP_425J2_127_3477_n2226), .A2(
        DP_OP_425J2_127_3477_n2230), .Y(DP_OP_425J2_127_3477_n2194) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1432 ( .A1(DP_OP_422J2_124_3477_n2093), .A2(
        DP_OP_425J2_127_3477_n2230), .Y(DP_OP_425J2_127_3477_n2193) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1431 ( .A1(DP_OP_422J2_124_3477_n2092), .A2(
        DP_OP_422J2_124_3477_n2230), .Y(DP_OP_425J2_127_3477_n2192) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1430 ( .A1(DP_OP_422J2_124_3477_n2091), .A2(
        DP_OP_423J2_125_3477_n2230), .Y(DP_OP_425J2_127_3477_n2191) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1429 ( .A1(DP_OP_422J2_124_3477_n2090), 
        .A2(DP_OP_425J2_127_3477_n2230), .Y(DP_OP_425J2_127_3477_n2190) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1409 ( .A1(DP_OP_424J2_126_3477_n2882), .A2(
        DP_OP_425J2_127_3477_n2189), .Y(DP_OP_425J2_127_3477_n2170) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1401 ( .A1(DP_OP_424J2_126_3477_n2882), .A2(
        n1345), .Y(DP_OP_425J2_127_3477_n2162) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1394 ( .A1(DP_OP_424J2_126_3477_n2883), 
        .A2(n1339), .Y(DP_OP_425J2_127_3477_n2155) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1393 ( .A1(DP_OP_424J2_126_3477_n2882), .A2(
        n1339), .Y(DP_OP_425J2_127_3477_n2154) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1392 ( .A1(DP_OP_425J2_127_3477_n2185), .A2(
        DP_OP_424J2_126_3477_n2186), .Y(DP_OP_425J2_127_3477_n2153) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1391 ( .A1(DP_OP_425J2_127_3477_n2184), .A2(
        DP_OP_422J2_124_3477_n2186), .Y(DP_OP_425J2_127_3477_n2152) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1389 ( .A1(DP_OP_425J2_127_3477_n2182), .A2(
        DP_OP_425J2_127_3477_n2186), .Y(DP_OP_425J2_127_3477_n2150) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1388 ( .A1(DP_OP_423J2_125_3477_n2973), .A2(
        DP_OP_425J2_127_3477_n2186), .Y(DP_OP_425J2_127_3477_n2149) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1387 ( .A1(DP_OP_425J2_127_3477_n2180), .A2(
        DP_OP_422J2_124_3477_n2186), .Y(DP_OP_425J2_127_3477_n2148) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1386 ( .A1(DP_OP_424J2_126_3477_n2883), .A2(
        DP_OP_425J2_127_3477_n2186), .Y(DP_OP_425J2_127_3477_n2147) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1385 ( .A1(DP_OP_424J2_126_3477_n2882), 
        .A2(DP_OP_422J2_124_3477_n2186), .Y(DP_OP_425J2_127_3477_n2146) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1358 ( .A1(DP_OP_422J2_124_3477_n2003), 
        .A2(DP_OP_422J2_124_3477_n2144), .Y(DP_OP_425J2_127_3477_n2119) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1357 ( .A1(DP_OP_423J2_125_3477_n3014), .A2(
        DP_OP_425J2_127_3477_n2144), .Y(DP_OP_425J2_127_3477_n2118) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1350 ( .A1(DP_OP_424J2_126_3477_n2927), 
        .A2(DP_OP_425J2_127_3477_n2143), .Y(DP_OP_425J2_127_3477_n2111) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1349 ( .A1(DP_OP_423J2_125_3477_n3014), .A2(
        DP_OP_425J2_127_3477_n2143), .Y(DP_OP_425J2_127_3477_n2110) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1348 ( .A1(DP_OP_424J2_126_3477_n2933), .A2(
        DP_OP_422J2_124_3477_n2142), .Y(DP_OP_425J2_127_3477_n2109) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1346 ( .A1(DP_OP_422J2_124_3477_n2007), .A2(
        DP_OP_422J2_124_3477_n2142), .Y(DP_OP_425J2_127_3477_n2107) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1345 ( .A1(DP_OP_425J2_127_3477_n2138), .A2(
        DP_OP_422J2_124_3477_n2142), .Y(DP_OP_425J2_127_3477_n2106) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1344 ( .A1(DP_OP_424J2_126_3477_n2929), .A2(
        DP_OP_422J2_124_3477_n2142), .Y(DP_OP_425J2_127_3477_n2105) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1342 ( .A1(DP_OP_424J2_126_3477_n2927), .A2(
        DP_OP_422J2_124_3477_n2142), .Y(DP_OP_425J2_127_3477_n2103) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1314 ( .A1(DP_OP_423J2_125_3477_n3057), 
        .A2(DP_OP_424J2_126_3477_n2100), .Y(DP_OP_425J2_127_3477_n2075) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1313 ( .A1(DP_OP_423J2_125_3477_n3056), .A2(
        DP_OP_424J2_126_3477_n2100), .Y(DP_OP_425J2_127_3477_n2074) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1306 ( .A1(DP_OP_423J2_125_3477_n3057), 
        .A2(DP_OP_425J2_127_3477_n2099), .Y(DP_OP_425J2_127_3477_n2067) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1305 ( .A1(DP_OP_423J2_125_3477_n3056), .A2(
        DP_OP_425J2_127_3477_n2099), .Y(DP_OP_425J2_127_3477_n2066) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1278 ( .A1(DP_OP_424J2_126_3477_n3015), 
        .A2(DP_OP_425J2_127_3477_n2057), .Y(DP_OP_425J2_127_3477_n2039) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1269 ( .A1(DP_OP_425J2_127_3477_n2046), .A2(
        DP_OP_425J2_127_3477_n2056), .Y(DP_OP_425J2_127_3477_n2030) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1262 ( .A1(DP_OP_424J2_126_3477_n3015), 
        .A2(DP_OP_425J2_127_3477_n2055), .Y(DP_OP_425J2_127_3477_n2023) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1261 ( .A1(DP_OP_425J2_127_3477_n2046), .A2(
        DP_OP_425J2_127_3477_n2055), .Y(DP_OP_425J2_127_3477_n2022) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1260 ( .A1(DP_OP_425J2_127_3477_n2053), .A2(
        n30), .Y(DP_OP_425J2_127_3477_n2021) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1259 ( .A1(DP_OP_424J2_126_3477_n3020), .A2(
        n30), .Y(DP_OP_425J2_127_3477_n2020) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1257 ( .A1(DP_OP_425J2_127_3477_n2050), .A2(
        n30), .Y(DP_OP_425J2_127_3477_n2018) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1256 ( .A1(DP_OP_425J2_127_3477_n2049), .A2(
        n30), .Y(DP_OP_425J2_127_3477_n2017) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1255 ( .A1(DP_OP_425J2_127_3477_n2048), .A2(
        n30), .Y(DP_OP_425J2_127_3477_n2016) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1254 ( .A1(DP_OP_424J2_126_3477_n3015), .A2(
        n777), .Y(DP_OP_425J2_127_3477_n2015) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1225 ( .A1(DP_OP_425J2_127_3477_n2002), .A2(
        n558), .Y(DP_OP_425J2_127_3477_n1986) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1217 ( .A1(DP_OP_425J2_127_3477_n2002), .A2(
        DP_OP_425J2_127_3477_n2011), .Y(DP_OP_425J2_127_3477_n1978) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1216 ( .A1(DP_OP_424J2_126_3477_n3063), .A2(
        DP_OP_425J2_127_3477_n2010), .Y(DP_OP_425J2_127_3477_n1977) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1215 ( .A1(DP_OP_425J2_127_3477_n2008), .A2(
        DP_OP_425J2_127_3477_n2010), .Y(DP_OP_425J2_127_3477_n1976) );
  OR2X1_HVT DP_OP_425J2_127_3477_U1214 ( .A1(DP_OP_425J2_127_3477_n2007), .A2(
        DP_OP_425J2_127_3477_n2010), .Y(DP_OP_425J2_127_3477_n1975) );
  HADDX1_HVT DP_OP_425J2_127_3477_U1143 ( .A0(DP_OP_425J2_127_3477_n1936), 
        .B0(DP_OP_425J2_127_3477_n2045), .C1(DP_OP_425J2_127_3477_n1920), .SO(
        DP_OP_425J2_127_3477_n1921) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1142 ( .A(DP_OP_425J2_127_3477_n2089), .B(
        DP_OP_425J2_127_3477_n2001), .CI(DP_OP_425J2_127_3477_n2133), .CO(
        DP_OP_425J2_127_3477_n1918), .S(DP_OP_425J2_127_3477_n1919) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1141 ( .A(DP_OP_425J2_127_3477_n2221), .B(
        DP_OP_425J2_127_3477_n2177), .CI(DP_OP_425J2_127_3477_n2265), .CO(
        DP_OP_425J2_127_3477_n1916), .S(DP_OP_425J2_127_3477_n1917) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1140 ( .A(DP_OP_425J2_127_3477_n2353), .B(
        DP_OP_425J2_127_3477_n2309), .CI(DP_OP_425J2_127_3477_n2397), .CO(
        DP_OP_425J2_127_3477_n1914), .S(DP_OP_425J2_127_3477_n1915) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1139 ( .A(DP_OP_425J2_127_3477_n2485), .B(
        DP_OP_425J2_127_3477_n2441), .CI(DP_OP_425J2_127_3477_n2529), .CO(
        DP_OP_425J2_127_3477_n1912), .S(DP_OP_425J2_127_3477_n1913) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1138 ( .A(DP_OP_425J2_127_3477_n2617), .B(
        DP_OP_425J2_127_3477_n2573), .CI(DP_OP_425J2_127_3477_n2661), .CO(
        DP_OP_425J2_127_3477_n1910), .S(DP_OP_425J2_127_3477_n1911) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1137 ( .A(DP_OP_425J2_127_3477_n2749), .B(
        DP_OP_425J2_127_3477_n2705), .CI(DP_OP_425J2_127_3477_n2793), .CO(
        DP_OP_425J2_127_3477_n1908), .S(DP_OP_425J2_127_3477_n1909) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1136 ( .A(DP_OP_425J2_127_3477_n3055), .B(
        DP_OP_425J2_127_3477_n2837), .CI(DP_OP_425J2_127_3477_n2881), .CO(
        DP_OP_425J2_127_3477_n1906), .S(DP_OP_425J2_127_3477_n1907) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1135 ( .A(DP_OP_425J2_127_3477_n3013), .B(
        DP_OP_425J2_127_3477_n2925), .CI(DP_OP_425J2_127_3477_n2969), .CO(
        DP_OP_425J2_127_3477_n1904), .S(DP_OP_425J2_127_3477_n1905) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1134 ( .A(DP_OP_425J2_127_3477_n1921), .B(
        DP_OP_425J2_127_3477_n1907), .CI(DP_OP_425J2_127_3477_n1909), .CO(
        DP_OP_425J2_127_3477_n1902), .S(DP_OP_425J2_127_3477_n1903) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1133 ( .A(DP_OP_425J2_127_3477_n1911), .B(
        DP_OP_425J2_127_3477_n1905), .CI(DP_OP_425J2_127_3477_n1913), .CO(
        DP_OP_425J2_127_3477_n1900), .S(DP_OP_425J2_127_3477_n1901) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1132 ( .A(DP_OP_425J2_127_3477_n1919), .B(
        DP_OP_425J2_127_3477_n1915), .CI(DP_OP_425J2_127_3477_n1917), .CO(
        DP_OP_425J2_127_3477_n1898), .S(DP_OP_425J2_127_3477_n1899) );
  HADDX1_HVT DP_OP_425J2_127_3477_U1131 ( .A0(DP_OP_425J2_127_3477_n1935), 
        .B0(DP_OP_425J2_127_3477_n2000), .C1(DP_OP_425J2_127_3477_n1896), .SO(
        DP_OP_425J2_127_3477_n1897) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1130 ( .A(DP_OP_425J2_127_3477_n2037), .B(
        DP_OP_425J2_127_3477_n1993), .CI(DP_OP_425J2_127_3477_n2044), .CO(
        DP_OP_425J2_127_3477_n1894), .S(DP_OP_425J2_127_3477_n1895) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1129 ( .A(DP_OP_425J2_127_3477_n2088), .B(
        DP_OP_425J2_127_3477_n2081), .CI(DP_OP_425J2_127_3477_n2125), .CO(
        DP_OP_425J2_127_3477_n1892), .S(DP_OP_425J2_127_3477_n1893) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1128 ( .A(DP_OP_425J2_127_3477_n2169), .B(
        DP_OP_425J2_127_3477_n2132), .CI(DP_OP_425J2_127_3477_n2176), .CO(
        DP_OP_425J2_127_3477_n1890), .S(DP_OP_425J2_127_3477_n1891) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1127 ( .A(DP_OP_425J2_127_3477_n2220), .B(
        DP_OP_425J2_127_3477_n2213), .CI(DP_OP_425J2_127_3477_n2257), .CO(
        DP_OP_425J2_127_3477_n1888), .S(DP_OP_425J2_127_3477_n1889) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1126 ( .A(DP_OP_425J2_127_3477_n2301), .B(
        DP_OP_425J2_127_3477_n2264), .CI(DP_OP_425J2_127_3477_n2308), .CO(
        DP_OP_425J2_127_3477_n1886), .S(DP_OP_425J2_127_3477_n1887) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1125 ( .A(DP_OP_425J2_127_3477_n2352), .B(
        DP_OP_425J2_127_3477_n2345), .CI(DP_OP_425J2_127_3477_n2389), .CO(
        DP_OP_425J2_127_3477_n1884), .S(DP_OP_425J2_127_3477_n1885) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1124 ( .A(DP_OP_425J2_127_3477_n2433), .B(
        DP_OP_425J2_127_3477_n2396), .CI(DP_OP_425J2_127_3477_n2440), .CO(
        DP_OP_425J2_127_3477_n1882), .S(DP_OP_425J2_127_3477_n1883) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1123 ( .A(DP_OP_425J2_127_3477_n2484), .B(
        DP_OP_425J2_127_3477_n2477), .CI(DP_OP_425J2_127_3477_n2521), .CO(
        DP_OP_425J2_127_3477_n1880), .S(DP_OP_425J2_127_3477_n1881) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1122 ( .A(DP_OP_425J2_127_3477_n2565), .B(
        DP_OP_425J2_127_3477_n2528), .CI(DP_OP_425J2_127_3477_n2572), .CO(
        DP_OP_425J2_127_3477_n1878), .S(DP_OP_425J2_127_3477_n1879) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1121 ( .A(DP_OP_425J2_127_3477_n3054), .B(
        DP_OP_425J2_127_3477_n2609), .CI(DP_OP_425J2_127_3477_n3047), .CO(
        DP_OP_425J2_127_3477_n1876), .S(DP_OP_425J2_127_3477_n1877) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1120 ( .A(DP_OP_425J2_127_3477_n2792), .B(
        DP_OP_425J2_127_3477_n2616), .CI(DP_OP_425J2_127_3477_n2653), .CO(
        DP_OP_425J2_127_3477_n1874), .S(DP_OP_425J2_127_3477_n1875) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1119 ( .A(DP_OP_425J2_127_3477_n2829), .B(
        DP_OP_425J2_127_3477_n3012), .CI(DP_OP_425J2_127_3477_n3005), .CO(
        DP_OP_425J2_127_3477_n1872), .S(DP_OP_425J2_127_3477_n1873) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1118 ( .A(DP_OP_425J2_127_3477_n2748), .B(
        DP_OP_425J2_127_3477_n2968), .CI(DP_OP_425J2_127_3477_n2961), .CO(
        DP_OP_425J2_127_3477_n1870), .S(DP_OP_425J2_127_3477_n1871) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1117 ( .A(DP_OP_425J2_127_3477_n2741), .B(
        DP_OP_425J2_127_3477_n2924), .CI(DP_OP_425J2_127_3477_n2660), .CO(
        DP_OP_425J2_127_3477_n1868), .S(DP_OP_425J2_127_3477_n1869) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1116 ( .A(DP_OP_425J2_127_3477_n2917), .B(
        DP_OP_425J2_127_3477_n2697), .CI(DP_OP_425J2_127_3477_n2704), .CO(
        DP_OP_425J2_127_3477_n1866), .S(DP_OP_425J2_127_3477_n1867) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1115 ( .A(DP_OP_425J2_127_3477_n2873), .B(
        DP_OP_425J2_127_3477_n2785), .CI(DP_OP_425J2_127_3477_n2836), .CO(
        DP_OP_425J2_127_3477_n1864), .S(DP_OP_425J2_127_3477_n1865) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1114 ( .A(DP_OP_425J2_127_3477_n2880), .B(
        DP_OP_425J2_127_3477_n1920), .CI(DP_OP_425J2_127_3477_n1897), .CO(
        DP_OP_425J2_127_3477_n1862), .S(DP_OP_425J2_127_3477_n1863) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1113 ( .A(DP_OP_425J2_127_3477_n1904), .B(
        DP_OP_425J2_127_3477_n1918), .CI(DP_OP_425J2_127_3477_n1916), .CO(
        DP_OP_425J2_127_3477_n1860), .S(DP_OP_425J2_127_3477_n1861) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1112 ( .A(DP_OP_425J2_127_3477_n1910), .B(
        DP_OP_425J2_127_3477_n1906), .CI(DP_OP_425J2_127_3477_n1914), .CO(
        DP_OP_425J2_127_3477_n1858), .S(DP_OP_425J2_127_3477_n1859) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1111 ( .A(DP_OP_425J2_127_3477_n1912), .B(
        DP_OP_425J2_127_3477_n1908), .CI(DP_OP_425J2_127_3477_n1865), .CO(
        DP_OP_425J2_127_3477_n1856), .S(DP_OP_425J2_127_3477_n1857) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1110 ( .A(DP_OP_425J2_127_3477_n1887), .B(
        DP_OP_425J2_127_3477_n1873), .CI(DP_OP_425J2_127_3477_n1871), .CO(
        DP_OP_425J2_127_3477_n1854), .S(DP_OP_425J2_127_3477_n1855) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1109 ( .A(DP_OP_425J2_127_3477_n1891), .B(
        DP_OP_425J2_127_3477_n1875), .CI(DP_OP_425J2_127_3477_n1879), .CO(
        DP_OP_425J2_127_3477_n1852), .S(DP_OP_425J2_127_3477_n1853) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1108 ( .A(DP_OP_425J2_127_3477_n1893), .B(
        DP_OP_425J2_127_3477_n1881), .CI(DP_OP_425J2_127_3477_n1877), .CO(
        DP_OP_425J2_127_3477_n1850), .S(DP_OP_425J2_127_3477_n1851) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1107 ( .A(DP_OP_425J2_127_3477_n1895), .B(
        DP_OP_425J2_127_3477_n1885), .CI(DP_OP_425J2_127_3477_n1869), .CO(
        DP_OP_425J2_127_3477_n1848), .S(DP_OP_425J2_127_3477_n1849) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1106 ( .A(DP_OP_425J2_127_3477_n1889), .B(
        DP_OP_425J2_127_3477_n1883), .CI(DP_OP_425J2_127_3477_n1867), .CO(
        DP_OP_425J2_127_3477_n1846), .S(DP_OP_425J2_127_3477_n1847) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1105 ( .A(DP_OP_425J2_127_3477_n1863), .B(
        DP_OP_425J2_127_3477_n1902), .CI(DP_OP_425J2_127_3477_n1900), .CO(
        DP_OP_425J2_127_3477_n1844), .S(DP_OP_425J2_127_3477_n1845) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1104 ( .A(DP_OP_425J2_127_3477_n1898), .B(
        DP_OP_425J2_127_3477_n1859), .CI(DP_OP_425J2_127_3477_n1861), .CO(
        DP_OP_425J2_127_3477_n1842), .S(DP_OP_425J2_127_3477_n1843) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1103 ( .A(DP_OP_425J2_127_3477_n1857), .B(
        DP_OP_425J2_127_3477_n1849), .CI(DP_OP_425J2_127_3477_n1851), .CO(
        DP_OP_425J2_127_3477_n1840), .S(DP_OP_425J2_127_3477_n1841) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1102 ( .A(DP_OP_425J2_127_3477_n1855), .B(
        DP_OP_425J2_127_3477_n1847), .CI(DP_OP_425J2_127_3477_n1853), .CO(
        DP_OP_425J2_127_3477_n1838), .S(DP_OP_425J2_127_3477_n1839) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1101 ( .A(DP_OP_425J2_127_3477_n1845), .B(
        DP_OP_425J2_127_3477_n1843), .CI(DP_OP_425J2_127_3477_n1841), .CO(
        DP_OP_425J2_127_3477_n1836), .S(DP_OP_425J2_127_3477_n1837) );
  HADDX1_HVT DP_OP_425J2_127_3477_U1100 ( .A0(DP_OP_425J2_127_3477_n1934), 
        .B0(DP_OP_425J2_127_3477_n1999), .C1(DP_OP_425J2_127_3477_n1834), .SO(
        DP_OP_425J2_127_3477_n1835) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1099 ( .A(DP_OP_425J2_127_3477_n2029), .B(
        DP_OP_425J2_127_3477_n1992), .CI(DP_OP_425J2_127_3477_n1985), .CO(
        DP_OP_425J2_127_3477_n1832), .S(DP_OP_425J2_127_3477_n1833) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1098 ( .A(DP_OP_425J2_127_3477_n2043), .B(
        DP_OP_425J2_127_3477_n2036), .CI(DP_OP_425J2_127_3477_n2073), .CO(
        DP_OP_425J2_127_3477_n1830), .S(DP_OP_425J2_127_3477_n1831) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1097 ( .A(DP_OP_425J2_127_3477_n2087), .B(
        DP_OP_425J2_127_3477_n2080), .CI(DP_OP_425J2_127_3477_n2117), .CO(
        DP_OP_425J2_127_3477_n1828), .S(DP_OP_425J2_127_3477_n1829) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1096 ( .A(DP_OP_425J2_127_3477_n2131), .B(
        DP_OP_425J2_127_3477_n2124), .CI(DP_OP_425J2_127_3477_n2161), .CO(
        DP_OP_425J2_127_3477_n1826), .S(DP_OP_425J2_127_3477_n1827) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1095 ( .A(DP_OP_425J2_127_3477_n2175), .B(
        DP_OP_425J2_127_3477_n2168), .CI(DP_OP_425J2_127_3477_n2205), .CO(
        DP_OP_425J2_127_3477_n1824), .S(DP_OP_425J2_127_3477_n1825) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1094 ( .A(DP_OP_425J2_127_3477_n2219), .B(
        DP_OP_425J2_127_3477_n2212), .CI(DP_OP_425J2_127_3477_n2249), .CO(
        DP_OP_425J2_127_3477_n1822), .S(DP_OP_425J2_127_3477_n1823) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1093 ( .A(DP_OP_425J2_127_3477_n2263), .B(
        DP_OP_425J2_127_3477_n2256), .CI(DP_OP_425J2_127_3477_n2293), .CO(
        DP_OP_425J2_127_3477_n1820), .S(DP_OP_425J2_127_3477_n1821) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1092 ( .A(DP_OP_425J2_127_3477_n2307), .B(
        DP_OP_425J2_127_3477_n2300), .CI(DP_OP_425J2_127_3477_n2337), .CO(
        DP_OP_425J2_127_3477_n1818), .S(DP_OP_425J2_127_3477_n1819) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1091 ( .A(DP_OP_425J2_127_3477_n2351), .B(
        DP_OP_425J2_127_3477_n2344), .CI(DP_OP_425J2_127_3477_n2381), .CO(
        DP_OP_425J2_127_3477_n1816), .S(DP_OP_425J2_127_3477_n1817) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1090 ( .A(DP_OP_425J2_127_3477_n2395), .B(
        DP_OP_425J2_127_3477_n2388), .CI(DP_OP_425J2_127_3477_n2425), .CO(
        DP_OP_425J2_127_3477_n1814), .S(DP_OP_425J2_127_3477_n1815) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1089 ( .A(DP_OP_425J2_127_3477_n2439), .B(
        DP_OP_425J2_127_3477_n2432), .CI(DP_OP_425J2_127_3477_n2469), .CO(
        DP_OP_425J2_127_3477_n1812), .S(DP_OP_425J2_127_3477_n1813) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1088 ( .A(DP_OP_425J2_127_3477_n2740), .B(
        DP_OP_425J2_127_3477_n3053), .CI(DP_OP_425J2_127_3477_n3046), .CO(
        DP_OP_425J2_127_3477_n1810), .S(DP_OP_425J2_127_3477_n1811) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1087 ( .A(DP_OP_425J2_127_3477_n2703), .B(
        DP_OP_425J2_127_3477_n2476), .CI(DP_OP_425J2_127_3477_n3039), .CO(
        DP_OP_425J2_127_3477_n1808), .S(DP_OP_425J2_127_3477_n1809) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1086 ( .A(DP_OP_425J2_127_3477_n2696), .B(
        DP_OP_425J2_127_3477_n3011), .CI(DP_OP_425J2_127_3477_n2483), .CO(
        DP_OP_425J2_127_3477_n1806), .S(DP_OP_425J2_127_3477_n1807) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1085 ( .A(DP_OP_425J2_127_3477_n2733), .B(
        DP_OP_425J2_127_3477_n2513), .CI(DP_OP_425J2_127_3477_n2520), .CO(
        DP_OP_425J2_127_3477_n1804), .S(DP_OP_425J2_127_3477_n1805) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1084 ( .A(DP_OP_425J2_127_3477_n2747), .B(
        DP_OP_425J2_127_3477_n2527), .CI(DP_OP_425J2_127_3477_n3004), .CO(
        DP_OP_425J2_127_3477_n1802), .S(DP_OP_425J2_127_3477_n1803) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1083 ( .A(DP_OP_425J2_127_3477_n2777), .B(
        DP_OP_425J2_127_3477_n2557), .CI(DP_OP_425J2_127_3477_n2997), .CO(
        DP_OP_425J2_127_3477_n1800), .S(DP_OP_425J2_127_3477_n1801) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1082 ( .A(DP_OP_425J2_127_3477_n2689), .B(
        DP_OP_425J2_127_3477_n2564), .CI(DP_OP_425J2_127_3477_n2967), .CO(
        DP_OP_425J2_127_3477_n1798), .S(DP_OP_425J2_127_3477_n1799) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1081 ( .A(DP_OP_425J2_127_3477_n2659), .B(
        DP_OP_425J2_127_3477_n2571), .CI(DP_OP_425J2_127_3477_n2960), .CO(
        DP_OP_425J2_127_3477_n1796), .S(DP_OP_425J2_127_3477_n1797) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1080 ( .A(DP_OP_425J2_127_3477_n2953), .B(
        DP_OP_425J2_127_3477_n2601), .CI(DP_OP_425J2_127_3477_n2608), .CO(
        DP_OP_425J2_127_3477_n1794), .S(DP_OP_425J2_127_3477_n1795) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1079 ( .A(DP_OP_425J2_127_3477_n2923), .B(
        DP_OP_425J2_127_3477_n2615), .CI(DP_OP_425J2_127_3477_n2645), .CO(
        DP_OP_425J2_127_3477_n1792), .S(DP_OP_425J2_127_3477_n1793) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1078 ( .A(DP_OP_425J2_127_3477_n2916), .B(
        DP_OP_425J2_127_3477_n2652), .CI(DP_OP_425J2_127_3477_n2784), .CO(
        DP_OP_425J2_127_3477_n1790), .S(DP_OP_425J2_127_3477_n1791) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1077 ( .A(DP_OP_425J2_127_3477_n2909), .B(
        DP_OP_425J2_127_3477_n2791), .CI(DP_OP_425J2_127_3477_n2821), .CO(
        DP_OP_425J2_127_3477_n1788), .S(DP_OP_425J2_127_3477_n1789) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1076 ( .A(DP_OP_425J2_127_3477_n2879), .B(
        DP_OP_425J2_127_3477_n2828), .CI(DP_OP_425J2_127_3477_n2835), .CO(
        DP_OP_425J2_127_3477_n1786), .S(DP_OP_425J2_127_3477_n1787) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1075 ( .A(DP_OP_425J2_127_3477_n2872), .B(
        DP_OP_425J2_127_3477_n2865), .CI(DP_OP_425J2_127_3477_n1896), .CO(
        DP_OP_425J2_127_3477_n1784), .S(DP_OP_425J2_127_3477_n1785) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1074 ( .A(DP_OP_425J2_127_3477_n1835), .B(
        DP_OP_425J2_127_3477_n1864), .CI(DP_OP_425J2_127_3477_n1866), .CO(
        DP_OP_425J2_127_3477_n1782), .S(DP_OP_425J2_127_3477_n1783) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1073 ( .A(DP_OP_425J2_127_3477_n1882), .B(
        DP_OP_425J2_127_3477_n1894), .CI(DP_OP_425J2_127_3477_n1868), .CO(
        DP_OP_425J2_127_3477_n1780), .S(DP_OP_425J2_127_3477_n1781) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1072 ( .A(DP_OP_425J2_127_3477_n1880), .B(
        DP_OP_425J2_127_3477_n1892), .CI(DP_OP_425J2_127_3477_n1870), .CO(
        DP_OP_425J2_127_3477_n1778), .S(DP_OP_425J2_127_3477_n1779) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1071 ( .A(DP_OP_425J2_127_3477_n1876), .B(
        DP_OP_425J2_127_3477_n1890), .CI(DP_OP_425J2_127_3477_n1872), .CO(
        DP_OP_425J2_127_3477_n1776), .S(DP_OP_425J2_127_3477_n1777) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1070 ( .A(DP_OP_425J2_127_3477_n1888), .B(
        DP_OP_425J2_127_3477_n1886), .CI(DP_OP_425J2_127_3477_n1884), .CO(
        DP_OP_425J2_127_3477_n1774), .S(DP_OP_425J2_127_3477_n1775) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1069 ( .A(DP_OP_425J2_127_3477_n1878), .B(
        DP_OP_425J2_127_3477_n1874), .CI(DP_OP_425J2_127_3477_n1807), .CO(
        DP_OP_425J2_127_3477_n1772), .S(DP_OP_425J2_127_3477_n1773) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1068 ( .A(DP_OP_425J2_127_3477_n1801), .B(
        DP_OP_425J2_127_3477_n1815), .CI(DP_OP_425J2_127_3477_n1819), .CO(
        DP_OP_425J2_127_3477_n1770), .S(DP_OP_425J2_127_3477_n1771) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1067 ( .A(DP_OP_425J2_127_3477_n1797), .B(
        DP_OP_425J2_127_3477_n1825), .CI(DP_OP_425J2_127_3477_n1827), .CO(
        DP_OP_425J2_127_3477_n1768), .S(DP_OP_425J2_127_3477_n1769) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1066 ( .A(DP_OP_425J2_127_3477_n1795), .B(
        DP_OP_425J2_127_3477_n1817), .CI(DP_OP_425J2_127_3477_n1831), .CO(
        DP_OP_425J2_127_3477_n1766), .S(DP_OP_425J2_127_3477_n1767) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1065 ( .A(DP_OP_425J2_127_3477_n1793), .B(
        DP_OP_425J2_127_3477_n1811), .CI(DP_OP_425J2_127_3477_n1829), .CO(
        DP_OP_425J2_127_3477_n1764), .S(DP_OP_425J2_127_3477_n1765) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1064 ( .A(DP_OP_425J2_127_3477_n1791), .B(
        DP_OP_425J2_127_3477_n1821), .CI(DP_OP_425J2_127_3477_n1809), .CO(
        DP_OP_425J2_127_3477_n1762), .S(DP_OP_425J2_127_3477_n1763) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1063 ( .A(DP_OP_425J2_127_3477_n1789), .B(
        DP_OP_425J2_127_3477_n1823), .CI(DP_OP_425J2_127_3477_n1833), .CO(
        DP_OP_425J2_127_3477_n1760), .S(DP_OP_425J2_127_3477_n1761) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1062 ( .A(DP_OP_425J2_127_3477_n1787), .B(
        DP_OP_425J2_127_3477_n1813), .CI(DP_OP_425J2_127_3477_n1799), .CO(
        DP_OP_425J2_127_3477_n1758), .S(DP_OP_425J2_127_3477_n1759) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1061 ( .A(DP_OP_425J2_127_3477_n1805), .B(
        DP_OP_425J2_127_3477_n1803), .CI(DP_OP_425J2_127_3477_n1862), .CO(
        DP_OP_425J2_127_3477_n1756), .S(DP_OP_425J2_127_3477_n1757) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1060 ( .A(DP_OP_425J2_127_3477_n1785), .B(
        DP_OP_425J2_127_3477_n1860), .CI(DP_OP_425J2_127_3477_n1858), .CO(
        DP_OP_425J2_127_3477_n1754), .S(DP_OP_425J2_127_3477_n1755) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1059 ( .A(DP_OP_425J2_127_3477_n1856), .B(
        DP_OP_425J2_127_3477_n1783), .CI(DP_OP_425J2_127_3477_n1850), .CO(
        DP_OP_425J2_127_3477_n1752), .S(DP_OP_425J2_127_3477_n1753) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1058 ( .A(DP_OP_425J2_127_3477_n1854), .B(
        DP_OP_425J2_127_3477_n1775), .CI(DP_OP_425J2_127_3477_n1781), .CO(
        DP_OP_425J2_127_3477_n1750), .S(DP_OP_425J2_127_3477_n1751) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1057 ( .A(DP_OP_425J2_127_3477_n1852), .B(
        DP_OP_425J2_127_3477_n1779), .CI(DP_OP_425J2_127_3477_n1777), .CO(
        DP_OP_425J2_127_3477_n1748), .S(DP_OP_425J2_127_3477_n1749) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1056 ( .A(DP_OP_425J2_127_3477_n1848), .B(
        DP_OP_425J2_127_3477_n1846), .CI(DP_OP_425J2_127_3477_n1773), .CO(
        DP_OP_425J2_127_3477_n1746), .S(DP_OP_425J2_127_3477_n1747) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1055 ( .A(DP_OP_425J2_127_3477_n1757), .B(
        DP_OP_425J2_127_3477_n1759), .CI(DP_OP_425J2_127_3477_n1771), .CO(
        DP_OP_425J2_127_3477_n1744), .S(DP_OP_425J2_127_3477_n1745) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1054 ( .A(DP_OP_425J2_127_3477_n1761), .B(
        DP_OP_425J2_127_3477_n1769), .CI(DP_OP_425J2_127_3477_n1767), .CO(
        DP_OP_425J2_127_3477_n1742), .S(DP_OP_425J2_127_3477_n1743) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1053 ( .A(DP_OP_425J2_127_3477_n1763), .B(
        DP_OP_425J2_127_3477_n1765), .CI(DP_OP_425J2_127_3477_n1844), .CO(
        DP_OP_425J2_127_3477_n1740), .S(DP_OP_425J2_127_3477_n1741) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1052 ( .A(DP_OP_425J2_127_3477_n1755), .B(
        DP_OP_425J2_127_3477_n1842), .CI(DP_OP_425J2_127_3477_n1753), .CO(
        DP_OP_425J2_127_3477_n1738), .S(DP_OP_425J2_127_3477_n1739) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1051 ( .A(DP_OP_425J2_127_3477_n1840), .B(
        DP_OP_425J2_127_3477_n1838), .CI(DP_OP_425J2_127_3477_n1749), .CO(
        DP_OP_425J2_127_3477_n1736), .S(DP_OP_425J2_127_3477_n1737) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1050 ( .A(DP_OP_425J2_127_3477_n1751), .B(
        DP_OP_425J2_127_3477_n1747), .CI(DP_OP_425J2_127_3477_n1745), .CO(
        DP_OP_425J2_127_3477_n1734), .S(DP_OP_425J2_127_3477_n1735) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1049 ( .A(DP_OP_425J2_127_3477_n1743), .B(
        DP_OP_425J2_127_3477_n1741), .CI(DP_OP_425J2_127_3477_n1739), .CO(
        DP_OP_425J2_127_3477_n1732), .S(DP_OP_425J2_127_3477_n1733) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1048 ( .A(DP_OP_425J2_127_3477_n1836), .B(
        DP_OP_425J2_127_3477_n1737), .CI(DP_OP_425J2_127_3477_n1735), .CO(
        DP_OP_425J2_127_3477_n1730), .S(DP_OP_425J2_127_3477_n1731) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1045 ( .A(DP_OP_425J2_127_3477_n2197), .B(
        DP_OP_425J2_127_3477_n2637), .CI(DP_OP_425J2_127_3477_n2417), .CO(
        DP_OP_425J2_127_3477_n1724), .S(DP_OP_425J2_127_3477_n1725) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1044 ( .A(DP_OP_425J2_127_3477_n2945), .B(
        DP_OP_425J2_127_3477_n2153), .CI(DP_OP_425J2_127_3477_n2373), .CO(
        DP_OP_425J2_127_3477_n1722), .S(DP_OP_425J2_127_3477_n1723) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1043 ( .A(DP_OP_425J2_127_3477_n2549), .B(
        DP_OP_425J2_127_3477_n2857), .CI(DP_OP_425J2_127_3477_n2461), .CO(
        DP_OP_425J2_127_3477_n1720), .S(DP_OP_425J2_127_3477_n1721) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1042 ( .A(DP_OP_425J2_127_3477_n2285), .B(
        DP_OP_425J2_127_3477_n2329), .CI(DP_OP_425J2_127_3477_n2109), .CO(
        DP_OP_425J2_127_3477_n1718), .S(DP_OP_425J2_127_3477_n1719) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1041 ( .A(DP_OP_425J2_127_3477_n2813), .B(
        DP_OP_425J2_127_3477_n2681), .CI(DP_OP_425J2_127_3477_n2725), .CO(
        DP_OP_425J2_127_3477_n1716), .S(DP_OP_425J2_127_3477_n1717) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1040 ( .A(DP_OP_425J2_127_3477_n2065), .B(
        DP_OP_425J2_127_3477_n2901), .CI(DP_OP_425J2_127_3477_n2769), .CO(
        DP_OP_425J2_127_3477_n1714), .S(DP_OP_425J2_127_3477_n1715) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1039 ( .A(DP_OP_425J2_127_3477_n2989), .B(
        DP_OP_425J2_127_3477_n2593), .CI(DP_OP_425J2_127_3477_n2241), .CO(
        DP_OP_425J2_127_3477_n1712), .S(DP_OP_425J2_127_3477_n1713) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1038 ( .A(DP_OP_425J2_127_3477_n2021), .B(
        DP_OP_425J2_127_3477_n1729), .CI(DP_OP_425J2_127_3477_n1998), .CO(
        DP_OP_425J2_127_3477_n1710), .S(DP_OP_425J2_127_3477_n1711) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1037 ( .A(DP_OP_425J2_127_3477_n2028), .B(
        DP_OP_425J2_127_3477_n1991), .CI(DP_OP_425J2_127_3477_n1984), .CO(
        DP_OP_425J2_127_3477_n1708), .S(DP_OP_425J2_127_3477_n1709) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1036 ( .A(DP_OP_425J2_127_3477_n2042), .B(
        DP_OP_425J2_127_3477_n2035), .CI(DP_OP_425J2_127_3477_n2072), .CO(
        DP_OP_425J2_127_3477_n1706), .S(DP_OP_425J2_127_3477_n1707) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1035 ( .A(DP_OP_425J2_127_3477_n2086), .B(
        DP_OP_425J2_127_3477_n2079), .CI(DP_OP_425J2_127_3477_n2116), .CO(
        DP_OP_425J2_127_3477_n1704), .S(DP_OP_425J2_127_3477_n1705) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1034 ( .A(DP_OP_425J2_127_3477_n3052), .B(
        DP_OP_425J2_127_3477_n2123), .CI(DP_OP_425J2_127_3477_n2130), .CO(
        DP_OP_425J2_127_3477_n1702), .S(DP_OP_425J2_127_3477_n1703) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1033 ( .A(DP_OP_425J2_127_3477_n2563), .B(
        DP_OP_425J2_127_3477_n3045), .CI(DP_OP_425J2_127_3477_n3038), .CO(
        DP_OP_425J2_127_3477_n1700), .S(DP_OP_425J2_127_3477_n1701) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1032 ( .A(DP_OP_425J2_127_3477_n2526), .B(
        DP_OP_425J2_127_3477_n2160), .CI(DP_OP_425J2_127_3477_n3010), .CO(
        DP_OP_425J2_127_3477_n1698), .S(DP_OP_425J2_127_3477_n1699) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1031 ( .A(DP_OP_425J2_127_3477_n2556), .B(
        DP_OP_425J2_127_3477_n2167), .CI(DP_OP_425J2_127_3477_n3003), .CO(
        DP_OP_425J2_127_3477_n1696), .S(DP_OP_425J2_127_3477_n1697) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1030 ( .A(DP_OP_425J2_127_3477_n2996), .B(
        DP_OP_425J2_127_3477_n2174), .CI(DP_OP_425J2_127_3477_n2204), .CO(
        DP_OP_425J2_127_3477_n1694), .S(DP_OP_425J2_127_3477_n1695) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1029 ( .A(DP_OP_425J2_127_3477_n2519), .B(
        DP_OP_425J2_127_3477_n2211), .CI(DP_OP_425J2_127_3477_n2218), .CO(
        DP_OP_425J2_127_3477_n1692), .S(DP_OP_425J2_127_3477_n1693) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1028 ( .A(DP_OP_425J2_127_3477_n2600), .B(
        DP_OP_425J2_127_3477_n2248), .CI(DP_OP_425J2_127_3477_n2255), .CO(
        DP_OP_425J2_127_3477_n1690), .S(DP_OP_425J2_127_3477_n1691) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1027 ( .A(DP_OP_425J2_127_3477_n2607), .B(
        DP_OP_425J2_127_3477_n2262), .CI(DP_OP_425J2_127_3477_n2292), .CO(
        DP_OP_425J2_127_3477_n1688), .S(DP_OP_425J2_127_3477_n1689) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1026 ( .A(DP_OP_425J2_127_3477_n2614), .B(
        DP_OP_425J2_127_3477_n2966), .CI(DP_OP_425J2_127_3477_n2299), .CO(
        DP_OP_425J2_127_3477_n1686), .S(DP_OP_425J2_127_3477_n1687) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1025 ( .A(DP_OP_425J2_127_3477_n2644), .B(
        DP_OP_425J2_127_3477_n2306), .CI(DP_OP_425J2_127_3477_n2959), .CO(
        DP_OP_425J2_127_3477_n1684), .S(DP_OP_425J2_127_3477_n1685) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1023 ( .A(DP_OP_425J2_127_3477_n2482), .B(
        DP_OP_425J2_127_3477_n2915), .CI(DP_OP_425J2_127_3477_n2336), .CO(
        DP_OP_425J2_127_3477_n1680), .S(DP_OP_425J2_127_3477_n1681) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1022 ( .A(DP_OP_425J2_127_3477_n2908), .B(
        DP_OP_425J2_127_3477_n2343), .CI(DP_OP_425J2_127_3477_n2878), .CO(
        DP_OP_425J2_127_3477_n1678), .S(DP_OP_425J2_127_3477_n1679) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1019 ( .A(DP_OP_425J2_127_3477_n2468), .B(
        DP_OP_425J2_127_3477_n2827), .CI(DP_OP_425J2_127_3477_n2820), .CO(
        DP_OP_425J2_127_3477_n1672), .S(DP_OP_425J2_127_3477_n1673) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1018 ( .A(DP_OP_425J2_127_3477_n2424), .B(
        DP_OP_425J2_127_3477_n2790), .CI(DP_OP_425J2_127_3477_n2783), .CO(
        DP_OP_425J2_127_3477_n1670), .S(DP_OP_425J2_127_3477_n1671) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1017 ( .A(DP_OP_425J2_127_3477_n2387), .B(
        DP_OP_425J2_127_3477_n2776), .CI(DP_OP_425J2_127_3477_n2746), .CO(
        DP_OP_425J2_127_3477_n1668), .S(DP_OP_425J2_127_3477_n1669) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1016 ( .A(DP_OP_425J2_127_3477_n2658), .B(
        DP_OP_425J2_127_3477_n2739), .CI(DP_OP_425J2_127_3477_n2394), .CO(
        DP_OP_425J2_127_3477_n1666), .S(DP_OP_425J2_127_3477_n1667) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1015 ( .A(DP_OP_425J2_127_3477_n2512), .B(
        DP_OP_425J2_127_3477_n2431), .CI(DP_OP_425J2_127_3477_n2732), .CO(
        DP_OP_425J2_127_3477_n1664), .S(DP_OP_425J2_127_3477_n1665) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1014 ( .A(DP_OP_425J2_127_3477_n2702), .B(
        DP_OP_425J2_127_3477_n2438), .CI(DP_OP_425J2_127_3477_n2651), .CO(
        DP_OP_425J2_127_3477_n1662), .S(DP_OP_425J2_127_3477_n1663) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1013 ( .A(DP_OP_425J2_127_3477_n2695), .B(
        DP_OP_425J2_127_3477_n2688), .CI(DP_OP_425J2_127_3477_n1834), .CO(
        DP_OP_425J2_127_3477_n1660), .S(DP_OP_425J2_127_3477_n1661) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1012 ( .A(DP_OP_425J2_127_3477_n1810), .B(
        DP_OP_425J2_127_3477_n1832), .CI(DP_OP_425J2_127_3477_n1786), .CO(
        DP_OP_425J2_127_3477_n1658), .S(DP_OP_425J2_127_3477_n1659) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1011 ( .A(DP_OP_425J2_127_3477_n1808), .B(
        DP_OP_425J2_127_3477_n1830), .CI(DP_OP_425J2_127_3477_n1828), .CO(
        DP_OP_425J2_127_3477_n1656), .S(DP_OP_425J2_127_3477_n1657) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1010 ( .A(DP_OP_425J2_127_3477_n1802), .B(
        DP_OP_425J2_127_3477_n1826), .CI(DP_OP_425J2_127_3477_n1824), .CO(
        DP_OP_425J2_127_3477_n1654), .S(DP_OP_425J2_127_3477_n1655) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1009 ( .A(DP_OP_425J2_127_3477_n1798), .B(
        DP_OP_425J2_127_3477_n1788), .CI(DP_OP_425J2_127_3477_n1790), .CO(
        DP_OP_425J2_127_3477_n1652), .S(DP_OP_425J2_127_3477_n1653) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1008 ( .A(DP_OP_425J2_127_3477_n1796), .B(
        DP_OP_425J2_127_3477_n1822), .CI(DP_OP_425J2_127_3477_n1792), .CO(
        DP_OP_425J2_127_3477_n1650), .S(DP_OP_425J2_127_3477_n1651) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1007 ( .A(DP_OP_425J2_127_3477_n1794), .B(
        DP_OP_425J2_127_3477_n1820), .CI(DP_OP_425J2_127_3477_n1818), .CO(
        DP_OP_425J2_127_3477_n1648), .S(DP_OP_425J2_127_3477_n1649) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1006 ( .A(DP_OP_425J2_127_3477_n1806), .B(
        DP_OP_425J2_127_3477_n1816), .CI(DP_OP_425J2_127_3477_n1800), .CO(
        DP_OP_425J2_127_3477_n1646), .S(DP_OP_425J2_127_3477_n1647) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1005 ( .A(DP_OP_425J2_127_3477_n1814), .B(
        DP_OP_425J2_127_3477_n1804), .CI(DP_OP_425J2_127_3477_n1812), .CO(
        DP_OP_425J2_127_3477_n1644), .S(DP_OP_425J2_127_3477_n1645) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1004 ( .A(DP_OP_425J2_127_3477_n1723), .B(
        DP_OP_425J2_127_3477_n1725), .CI(DP_OP_425J2_127_3477_n1711), .CO(
        DP_OP_425J2_127_3477_n1642), .S(DP_OP_425J2_127_3477_n1643) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1003 ( .A(DP_OP_425J2_127_3477_n1717), .B(
        DP_OP_425J2_127_3477_n1719), .CI(DP_OP_425J2_127_3477_n1784), .CO(
        DP_OP_425J2_127_3477_n1640), .S(DP_OP_425J2_127_3477_n1641) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1002 ( .A(DP_OP_425J2_127_3477_n1713), .B(
        DP_OP_425J2_127_3477_n1715), .CI(DP_OP_425J2_127_3477_n1721), .CO(
        DP_OP_425J2_127_3477_n1638), .S(DP_OP_425J2_127_3477_n1639) );
  FADDX1_HVT DP_OP_425J2_127_3477_U1000 ( .A(DP_OP_425J2_127_3477_n1679), .B(
        DP_OP_425J2_127_3477_n1695), .CI(DP_OP_425J2_127_3477_n1703), .CO(
        DP_OP_425J2_127_3477_n1634), .S(DP_OP_425J2_127_3477_n1635) );
  FADDX1_HVT DP_OP_425J2_127_3477_U999 ( .A(DP_OP_425J2_127_3477_n1671), .B(
        DP_OP_425J2_127_3477_n1691), .CI(DP_OP_425J2_127_3477_n1689), .CO(
        DP_OP_425J2_127_3477_n1632), .S(DP_OP_425J2_127_3477_n1633) );
  FADDX1_HVT DP_OP_425J2_127_3477_U998 ( .A(DP_OP_425J2_127_3477_n1669), .B(
        DP_OP_425J2_127_3477_n1705), .CI(DP_OP_425J2_127_3477_n1693), .CO(
        DP_OP_425J2_127_3477_n1630), .S(DP_OP_425J2_127_3477_n1631) );
  FADDX1_HVT DP_OP_425J2_127_3477_U997 ( .A(DP_OP_425J2_127_3477_n1667), .B(
        DP_OP_425J2_127_3477_n1699), .CI(DP_OP_425J2_127_3477_n1701), .CO(
        DP_OP_425J2_127_3477_n1628), .S(DP_OP_425J2_127_3477_n1629) );
  FADDX1_HVT DP_OP_425J2_127_3477_U996 ( .A(DP_OP_425J2_127_3477_n1665), .B(
        DP_OP_425J2_127_3477_n1697), .CI(DP_OP_425J2_127_3477_n1709), .CO(
        DP_OP_425J2_127_3477_n1626), .S(DP_OP_425J2_127_3477_n1627) );
  FADDX1_HVT DP_OP_425J2_127_3477_U995 ( .A(DP_OP_425J2_127_3477_n1687), .B(
        DP_OP_425J2_127_3477_n1707), .CI(DP_OP_425J2_127_3477_n1663), .CO(
        DP_OP_425J2_127_3477_n1624), .S(DP_OP_425J2_127_3477_n1625) );
  FADDX1_HVT DP_OP_425J2_127_3477_U994 ( .A(DP_OP_425J2_127_3477_n1673), .B(
        DP_OP_425J2_127_3477_n1683), .CI(DP_OP_425J2_127_3477_n1685), .CO(
        DP_OP_425J2_127_3477_n1622), .S(DP_OP_425J2_127_3477_n1623) );
  FADDX1_HVT DP_OP_425J2_127_3477_U993 ( .A(DP_OP_425J2_127_3477_n1681), .B(
        DP_OP_425J2_127_3477_n1661), .CI(DP_OP_425J2_127_3477_n1782), .CO(
        DP_OP_425J2_127_3477_n1620), .S(DP_OP_425J2_127_3477_n1621) );
  FADDX1_HVT DP_OP_425J2_127_3477_U992 ( .A(DP_OP_425J2_127_3477_n1780), .B(
        DP_OP_425J2_127_3477_n1778), .CI(DP_OP_425J2_127_3477_n1776), .CO(
        DP_OP_425J2_127_3477_n1618), .S(DP_OP_425J2_127_3477_n1619) );
  FADDX1_HVT DP_OP_425J2_127_3477_U991 ( .A(DP_OP_425J2_127_3477_n1774), .B(
        DP_OP_425J2_127_3477_n1772), .CI(DP_OP_425J2_127_3477_n1760), .CO(
        DP_OP_425J2_127_3477_n1616), .S(DP_OP_425J2_127_3477_n1617) );
  FADDX1_HVT DP_OP_425J2_127_3477_U990 ( .A(DP_OP_425J2_127_3477_n1758), .B(
        DP_OP_425J2_127_3477_n1659), .CI(DP_OP_425J2_127_3477_n1756), .CO(
        DP_OP_425J2_127_3477_n1614), .S(DP_OP_425J2_127_3477_n1615) );
  FADDX1_HVT DP_OP_425J2_127_3477_U989 ( .A(DP_OP_425J2_127_3477_n1657), .B(
        DP_OP_425J2_127_3477_n1649), .CI(DP_OP_425J2_127_3477_n1770), .CO(
        DP_OP_425J2_127_3477_n1612), .S(DP_OP_425J2_127_3477_n1613) );
  FADDX1_HVT DP_OP_425J2_127_3477_U988 ( .A(DP_OP_425J2_127_3477_n1768), .B(
        DP_OP_425J2_127_3477_n1647), .CI(DP_OP_425J2_127_3477_n1651), .CO(
        DP_OP_425J2_127_3477_n1610), .S(DP_OP_425J2_127_3477_n1611) );
  FADDX1_HVT DP_OP_425J2_127_3477_U987 ( .A(DP_OP_425J2_127_3477_n1764), .B(
        DP_OP_425J2_127_3477_n1655), .CI(DP_OP_425J2_127_3477_n1653), .CO(
        DP_OP_425J2_127_3477_n1608), .S(DP_OP_425J2_127_3477_n1609) );
  FADDX1_HVT DP_OP_425J2_127_3477_U986 ( .A(DP_OP_425J2_127_3477_n1762), .B(
        DP_OP_425J2_127_3477_n1766), .CI(DP_OP_425J2_127_3477_n1645), .CO(
        DP_OP_425J2_127_3477_n1606), .S(DP_OP_425J2_127_3477_n1607) );
  FADDX1_HVT DP_OP_425J2_127_3477_U985 ( .A(DP_OP_425J2_127_3477_n1641), .B(
        DP_OP_425J2_127_3477_n1643), .CI(DP_OP_425J2_127_3477_n1637), .CO(
        DP_OP_425J2_127_3477_n1604), .S(DP_OP_425J2_127_3477_n1605) );
  FADDX1_HVT DP_OP_425J2_127_3477_U984 ( .A(DP_OP_425J2_127_3477_n1639), .B(
        DP_OP_425J2_127_3477_n1625), .CI(DP_OP_425J2_127_3477_n1627), .CO(
        DP_OP_425J2_127_3477_n1602), .S(DP_OP_425J2_127_3477_n1603) );
  FADDX1_HVT DP_OP_425J2_127_3477_U983 ( .A(DP_OP_425J2_127_3477_n1633), .B(
        DP_OP_425J2_127_3477_n1631), .CI(DP_OP_425J2_127_3477_n1754), .CO(
        DP_OP_425J2_127_3477_n1600), .S(DP_OP_425J2_127_3477_n1601) );
  FADDX1_HVT DP_OP_425J2_127_3477_U982 ( .A(DP_OP_425J2_127_3477_n1629), .B(
        DP_OP_425J2_127_3477_n1623), .CI(DP_OP_425J2_127_3477_n1635), .CO(
        DP_OP_425J2_127_3477_n1598), .S(DP_OP_425J2_127_3477_n1599) );
  FADDX1_HVT DP_OP_425J2_127_3477_U981 ( .A(DP_OP_425J2_127_3477_n1621), .B(
        DP_OP_425J2_127_3477_n1752), .CI(DP_OP_425J2_127_3477_n1748), .CO(
        DP_OP_425J2_127_3477_n1596), .S(DP_OP_425J2_127_3477_n1597) );
  FADDX1_HVT DP_OP_425J2_127_3477_U980 ( .A(DP_OP_425J2_127_3477_n1750), .B(
        DP_OP_425J2_127_3477_n1619), .CI(DP_OP_425J2_127_3477_n1746), .CO(
        DP_OP_425J2_127_3477_n1594), .S(DP_OP_425J2_127_3477_n1595) );
  FADDX1_HVT DP_OP_425J2_127_3477_U979 ( .A(DP_OP_425J2_127_3477_n1617), .B(
        DP_OP_425J2_127_3477_n1607), .CI(DP_OP_425J2_127_3477_n1609), .CO(
        DP_OP_425J2_127_3477_n1592), .S(DP_OP_425J2_127_3477_n1593) );
  FADDX1_HVT DP_OP_425J2_127_3477_U977 ( .A(DP_OP_425J2_127_3477_n1615), .B(
        DP_OP_425J2_127_3477_n1613), .CI(DP_OP_425J2_127_3477_n1605), .CO(
        DP_OP_425J2_127_3477_n1588), .S(DP_OP_425J2_127_3477_n1589) );
  FADDX1_HVT DP_OP_425J2_127_3477_U976 ( .A(DP_OP_425J2_127_3477_n1740), .B(
        DP_OP_425J2_127_3477_n1603), .CI(DP_OP_425J2_127_3477_n1599), .CO(
        DP_OP_425J2_127_3477_n1586), .S(DP_OP_425J2_127_3477_n1587) );
  FADDX1_HVT DP_OP_425J2_127_3477_U975 ( .A(DP_OP_425J2_127_3477_n1601), .B(
        DP_OP_425J2_127_3477_n1738), .CI(DP_OP_425J2_127_3477_n1597), .CO(
        DP_OP_425J2_127_3477_n1584), .S(DP_OP_425J2_127_3477_n1585) );
  FADDX1_HVT DP_OP_425J2_127_3477_U974 ( .A(DP_OP_425J2_127_3477_n1736), .B(
        DP_OP_425J2_127_3477_n1595), .CI(DP_OP_425J2_127_3477_n1734), .CO(
        DP_OP_425J2_127_3477_n1582), .S(DP_OP_425J2_127_3477_n1583) );
  FADDX1_HVT DP_OP_425J2_127_3477_U973 ( .A(DP_OP_425J2_127_3477_n1593), .B(
        DP_OP_425J2_127_3477_n1591), .CI(DP_OP_425J2_127_3477_n1589), .CO(
        DP_OP_425J2_127_3477_n1580), .S(DP_OP_425J2_127_3477_n1581) );
  FADDX1_HVT DP_OP_425J2_127_3477_U972 ( .A(DP_OP_425J2_127_3477_n1587), .B(
        DP_OP_425J2_127_3477_n1732), .CI(DP_OP_425J2_127_3477_n1585), .CO(
        DP_OP_425J2_127_3477_n1578), .S(DP_OP_425J2_127_3477_n1579) );
  FADDX1_HVT DP_OP_425J2_127_3477_U970 ( .A(DP_OP_425J2_127_3477_n1728), .B(
        DP_OP_425J2_127_3477_n1976), .CI(DP_OP_425J2_127_3477_n1932), .CO(
        DP_OP_425J2_127_3477_n1574), .S(DP_OP_425J2_127_3477_n1575) );
  FADDX1_HVT DP_OP_425J2_127_3477_U969 ( .A(DP_OP_425J2_127_3477_n3031), .B(
        DP_OP_425J2_127_3477_n2548), .CI(DP_OP_425J2_127_3477_n2416), .CO(
        DP_OP_425J2_127_3477_n1572), .S(DP_OP_425J2_127_3477_n1573) );
  FADDX1_HVT DP_OP_425J2_127_3477_U968 ( .A(DP_OP_425J2_127_3477_n2944), .B(
        DP_OP_425J2_127_3477_n2680), .CI(DP_OP_425J2_127_3477_n2328), .CO(
        DP_OP_425J2_127_3477_n1570), .S(DP_OP_425J2_127_3477_n1571) );
  FADDX1_HVT DP_OP_425J2_127_3477_U967 ( .A(DP_OP_425J2_127_3477_n2108), .B(
        DP_OP_425J2_127_3477_n2636), .CI(DP_OP_425J2_127_3477_n2856), .CO(
        DP_OP_425J2_127_3477_n1568), .S(DP_OP_425J2_127_3477_n1569) );
  FADDX1_HVT DP_OP_425J2_127_3477_U966 ( .A(DP_OP_425J2_127_3477_n2196), .B(
        DP_OP_425J2_127_3477_n2372), .CI(DP_OP_425J2_127_3477_n2460), .CO(
        DP_OP_425J2_127_3477_n1566), .S(DP_OP_425J2_127_3477_n1567) );
  FADDX1_HVT DP_OP_425J2_127_3477_U965 ( .A(DP_OP_425J2_127_3477_n2812), .B(
        DP_OP_425J2_127_3477_n2284), .CI(DP_OP_425J2_127_3477_n2900), .CO(
        DP_OP_425J2_127_3477_n1564), .S(DP_OP_425J2_127_3477_n1565) );
  FADDX1_HVT DP_OP_425J2_127_3477_U964 ( .A(DP_OP_425J2_127_3477_n2152), .B(
        DP_OP_425J2_127_3477_n2504), .CI(DP_OP_425J2_127_3477_n2592), .CO(
        DP_OP_425J2_127_3477_n1562), .S(DP_OP_425J2_127_3477_n1563) );
  FADDX1_HVT DP_OP_425J2_127_3477_U963 ( .A(DP_OP_425J2_127_3477_n2988), .B(
        DP_OP_425J2_127_3477_n2724), .CI(DP_OP_425J2_127_3477_n2768), .CO(
        DP_OP_425J2_127_3477_n1560), .S(DP_OP_425J2_127_3477_n1561) );
  FADDX1_HVT DP_OP_425J2_127_3477_U962 ( .A(DP_OP_425J2_127_3477_n2064), .B(
        DP_OP_425J2_127_3477_n2240), .CI(DP_OP_425J2_127_3477_n2020), .CO(
        DP_OP_425J2_127_3477_n1558), .S(DP_OP_425J2_127_3477_n1559) );
  FADDX1_HVT DP_OP_425J2_127_3477_U961 ( .A(DP_OP_425J2_127_3477_n2555), .B(
        DP_OP_425J2_127_3477_n1990), .CI(DP_OP_425J2_127_3477_n1983), .CO(
        DP_OP_425J2_127_3477_n1556), .S(DP_OP_425J2_127_3477_n1557) );
  FADDX1_HVT DP_OP_425J2_127_3477_U960 ( .A(DP_OP_425J2_127_3477_n3051), .B(
        DP_OP_425J2_127_3477_n1997), .CI(DP_OP_425J2_127_3477_n2027), .CO(
        DP_OP_425J2_127_3477_n1554), .S(DP_OP_425J2_127_3477_n1555) );
  FADDX1_HVT DP_OP_425J2_127_3477_U959 ( .A(DP_OP_425J2_127_3477_n2437), .B(
        DP_OP_425J2_127_3477_n3044), .CI(DP_OP_425J2_127_3477_n2034), .CO(
        DP_OP_425J2_127_3477_n1552), .S(DP_OP_425J2_127_3477_n1553) );
  FADDX1_HVT DP_OP_425J2_127_3477_U958 ( .A(DP_OP_425J2_127_3477_n2430), .B(
        DP_OP_425J2_127_3477_n3037), .CI(DP_OP_425J2_127_3477_n2041), .CO(
        DP_OP_425J2_127_3477_n1550), .S(DP_OP_425J2_127_3477_n1551) );
  FADDX1_HVT DP_OP_425J2_127_3477_U957 ( .A(DP_OP_425J2_127_3477_n3009), .B(
        DP_OP_425J2_127_3477_n2071), .CI(DP_OP_425J2_127_3477_n2078), .CO(
        DP_OP_425J2_127_3477_n1548), .S(DP_OP_425J2_127_3477_n1549) );
  FADDX1_HVT DP_OP_425J2_127_3477_U956 ( .A(DP_OP_425J2_127_3477_n2467), .B(
        DP_OP_425J2_127_3477_n3002), .CI(DP_OP_425J2_127_3477_n2995), .CO(
        DP_OP_425J2_127_3477_n1546), .S(DP_OP_425J2_127_3477_n1547) );
  FADDX1_HVT DP_OP_425J2_127_3477_U955 ( .A(DP_OP_425J2_127_3477_n2393), .B(
        DP_OP_425J2_127_3477_n2965), .CI(DP_OP_425J2_127_3477_n2958), .CO(
        DP_OP_425J2_127_3477_n1544), .S(DP_OP_425J2_127_3477_n1545) );
  FADDX1_HVT DP_OP_425J2_127_3477_U954 ( .A(DP_OP_425J2_127_3477_n2386), .B(
        DP_OP_425J2_127_3477_n2951), .CI(DP_OP_425J2_127_3477_n2085), .CO(
        DP_OP_425J2_127_3477_n1542), .S(DP_OP_425J2_127_3477_n1543) );
  FADDX1_HVT DP_OP_425J2_127_3477_U953 ( .A(DP_OP_425J2_127_3477_n2379), .B(
        DP_OP_425J2_127_3477_n2921), .CI(DP_OP_425J2_127_3477_n2914), .CO(
        DP_OP_425J2_127_3477_n1540), .S(DP_OP_425J2_127_3477_n1541) );
  FADDX1_HVT DP_OP_425J2_127_3477_U952 ( .A(DP_OP_425J2_127_3477_n2349), .B(
        DP_OP_425J2_127_3477_n2907), .CI(DP_OP_425J2_127_3477_n2115), .CO(
        DP_OP_425J2_127_3477_n1538), .S(DP_OP_425J2_127_3477_n1539) );
  FADDX1_HVT DP_OP_425J2_127_3477_U951 ( .A(DP_OP_425J2_127_3477_n2342), .B(
        DP_OP_425J2_127_3477_n2122), .CI(DP_OP_425J2_127_3477_n2129), .CO(
        DP_OP_425J2_127_3477_n1536), .S(DP_OP_425J2_127_3477_n1537) );
  FADDX1_HVT DP_OP_425J2_127_3477_U950 ( .A(DP_OP_425J2_127_3477_n2423), .B(
        DP_OP_425J2_127_3477_n2159), .CI(DP_OP_425J2_127_3477_n2877), .CO(
        DP_OP_425J2_127_3477_n1534), .S(DP_OP_425J2_127_3477_n1535) );
  FADDX1_HVT DP_OP_425J2_127_3477_U949 ( .A(DP_OP_425J2_127_3477_n2474), .B(
        DP_OP_425J2_127_3477_n2870), .CI(DP_OP_425J2_127_3477_n2863), .CO(
        DP_OP_425J2_127_3477_n1532), .S(DP_OP_425J2_127_3477_n1533) );
  FADDX1_HVT DP_OP_425J2_127_3477_U948 ( .A(DP_OP_425J2_127_3477_n2833), .B(
        DP_OP_425J2_127_3477_n2166), .CI(DP_OP_425J2_127_3477_n2173), .CO(
        DP_OP_425J2_127_3477_n1530), .S(DP_OP_425J2_127_3477_n1531) );
  FADDX1_HVT DP_OP_425J2_127_3477_U947 ( .A(DP_OP_425J2_127_3477_n2606), .B(
        DP_OP_425J2_127_3477_n2203), .CI(DP_OP_425J2_127_3477_n2210), .CO(
        DP_OP_425J2_127_3477_n1528), .S(DP_OP_425J2_127_3477_n1529) );
  FADDX1_HVT DP_OP_425J2_127_3477_U946 ( .A(DP_OP_425J2_127_3477_n2826), .B(
        DP_OP_425J2_127_3477_n2217), .CI(DP_OP_425J2_127_3477_n2247), .CO(
        DP_OP_425J2_127_3477_n1526), .S(DP_OP_425J2_127_3477_n1527) );
  FADDX1_HVT DP_OP_425J2_127_3477_U945 ( .A(DP_OP_425J2_127_3477_n2819), .B(
        DP_OP_425J2_127_3477_n2254), .CI(DP_OP_425J2_127_3477_n2261), .CO(
        DP_OP_425J2_127_3477_n1524), .S(DP_OP_425J2_127_3477_n1525) );
  FADDX1_HVT DP_OP_425J2_127_3477_U944 ( .A(DP_OP_425J2_127_3477_n2789), .B(
        DP_OP_425J2_127_3477_n2291), .CI(DP_OP_425J2_127_3477_n2298), .CO(
        DP_OP_425J2_127_3477_n1522), .S(DP_OP_425J2_127_3477_n1523) );
  FADDX1_HVT DP_OP_425J2_127_3477_U943 ( .A(DP_OP_425J2_127_3477_n2782), .B(
        DP_OP_425J2_127_3477_n2305), .CI(DP_OP_425J2_127_3477_n2335), .CO(
        DP_OP_425J2_127_3477_n1520), .S(DP_OP_425J2_127_3477_n1521) );
  FADDX1_HVT DP_OP_425J2_127_3477_U942 ( .A(DP_OP_425J2_127_3477_n2775), .B(
        DP_OP_425J2_127_3477_n2481), .CI(DP_OP_425J2_127_3477_n2511), .CO(
        DP_OP_425J2_127_3477_n1518), .S(DP_OP_425J2_127_3477_n1519) );
  FADDX1_HVT DP_OP_425J2_127_3477_U941 ( .A(DP_OP_425J2_127_3477_n2745), .B(
        DP_OP_425J2_127_3477_n2518), .CI(DP_OP_425J2_127_3477_n2738), .CO(
        DP_OP_425J2_127_3477_n1516), .S(DP_OP_425J2_127_3477_n1517) );
  FADDX1_HVT DP_OP_425J2_127_3477_U940 ( .A(DP_OP_425J2_127_3477_n2643), .B(
        DP_OP_425J2_127_3477_n2525), .CI(DP_OP_425J2_127_3477_n2562), .CO(
        DP_OP_425J2_127_3477_n1514), .S(DP_OP_425J2_127_3477_n1515) );
  FADDX1_HVT DP_OP_425J2_127_3477_U939 ( .A(DP_OP_425J2_127_3477_n2613), .B(
        DP_OP_425J2_127_3477_n2569), .CI(DP_OP_425J2_127_3477_n2731), .CO(
        DP_OP_425J2_127_3477_n1512), .S(DP_OP_425J2_127_3477_n1513) );
  FADDX1_HVT DP_OP_425J2_127_3477_U938 ( .A(DP_OP_425J2_127_3477_n2687), .B(
        DP_OP_425J2_127_3477_n2599), .CI(DP_OP_425J2_127_3477_n2701), .CO(
        DP_OP_425J2_127_3477_n1510), .S(DP_OP_425J2_127_3477_n1511) );
  FADDX1_HVT DP_OP_425J2_127_3477_U937 ( .A(DP_OP_425J2_127_3477_n2650), .B(
        DP_OP_425J2_127_3477_n2657), .CI(DP_OP_425J2_127_3477_n2694), .CO(
        DP_OP_425J2_127_3477_n1508), .S(DP_OP_425J2_127_3477_n1509) );
  FADDX1_HVT DP_OP_425J2_127_3477_U936 ( .A(DP_OP_425J2_127_3477_n1716), .B(
        DP_OP_425J2_127_3477_n1712), .CI(DP_OP_425J2_127_3477_n1710), .CO(
        DP_OP_425J2_127_3477_n1506), .S(DP_OP_425J2_127_3477_n1507) );
  FADDX1_HVT DP_OP_425J2_127_3477_U935 ( .A(DP_OP_425J2_127_3477_n1714), .B(
        DP_OP_425J2_127_3477_n1718), .CI(DP_OP_425J2_127_3477_n1720), .CO(
        DP_OP_425J2_127_3477_n1504), .S(DP_OP_425J2_127_3477_n1505) );
  FADDX1_HVT DP_OP_425J2_127_3477_U934 ( .A(DP_OP_425J2_127_3477_n1722), .B(
        DP_OP_425J2_127_3477_n1724), .CI(DP_OP_425J2_127_3477_n1726), .CO(
        DP_OP_425J2_127_3477_n1502), .S(DP_OP_425J2_127_3477_n1503) );
  FADDX1_HVT DP_OP_425J2_127_3477_U933 ( .A(DP_OP_425J2_127_3477_n1686), .B(
        DP_OP_425J2_127_3477_n1708), .CI(DP_OP_425J2_127_3477_n1706), .CO(
        DP_OP_425J2_127_3477_n1500), .S(DP_OP_425J2_127_3477_n1501) );
  FADDX1_HVT DP_OP_425J2_127_3477_U932 ( .A(DP_OP_425J2_127_3477_n1682), .B(
        DP_OP_425J2_127_3477_n1704), .CI(DP_OP_425J2_127_3477_n1702), .CO(
        DP_OP_425J2_127_3477_n1498), .S(DP_OP_425J2_127_3477_n1499) );
  FADDX1_HVT DP_OP_425J2_127_3477_U931 ( .A(DP_OP_425J2_127_3477_n1676), .B(
        DP_OP_425J2_127_3477_n1700), .CI(DP_OP_425J2_127_3477_n1698), .CO(
        DP_OP_425J2_127_3477_n1496), .S(DP_OP_425J2_127_3477_n1497) );
  FADDX1_HVT DP_OP_425J2_127_3477_U930 ( .A(DP_OP_425J2_127_3477_n1672), .B(
        DP_OP_425J2_127_3477_n1696), .CI(DP_OP_425J2_127_3477_n1662), .CO(
        DP_OP_425J2_127_3477_n1494), .S(DP_OP_425J2_127_3477_n1495) );
  FADDX1_HVT DP_OP_425J2_127_3477_U929 ( .A(DP_OP_425J2_127_3477_n1668), .B(
        DP_OP_425J2_127_3477_n1694), .CI(DP_OP_425J2_127_3477_n1692), .CO(
        DP_OP_425J2_127_3477_n1492), .S(DP_OP_425J2_127_3477_n1493) );
  FADDX1_HVT DP_OP_425J2_127_3477_U928 ( .A(DP_OP_425J2_127_3477_n1678), .B(
        DP_OP_425J2_127_3477_n1690), .CI(DP_OP_425J2_127_3477_n1688), .CO(
        DP_OP_425J2_127_3477_n1490), .S(DP_OP_425J2_127_3477_n1491) );
  FADDX1_HVT DP_OP_425J2_127_3477_U927 ( .A(DP_OP_425J2_127_3477_n1670), .B(
        DP_OP_425J2_127_3477_n1684), .CI(DP_OP_425J2_127_3477_n1680), .CO(
        DP_OP_425J2_127_3477_n1488), .S(DP_OP_425J2_127_3477_n1489) );
  FADDX1_HVT DP_OP_425J2_127_3477_U926 ( .A(DP_OP_425J2_127_3477_n1666), .B(
        DP_OP_425J2_127_3477_n1674), .CI(DP_OP_425J2_127_3477_n1664), .CO(
        DP_OP_425J2_127_3477_n1486), .S(DP_OP_425J2_127_3477_n1487) );
  FADDX1_HVT DP_OP_425J2_127_3477_U925 ( .A(DP_OP_425J2_127_3477_n1575), .B(
        DP_OP_425J2_127_3477_n1559), .CI(DP_OP_425J2_127_3477_n1660), .CO(
        DP_OP_425J2_127_3477_n1484), .S(DP_OP_425J2_127_3477_n1485) );
  FADDX1_HVT DP_OP_425J2_127_3477_U924 ( .A(DP_OP_425J2_127_3477_n1573), .B(
        DP_OP_425J2_127_3477_n1561), .CI(DP_OP_425J2_127_3477_n1563), .CO(
        DP_OP_425J2_127_3477_n1482), .S(DP_OP_425J2_127_3477_n1483) );
  FADDX1_HVT DP_OP_425J2_127_3477_U923 ( .A(DP_OP_425J2_127_3477_n1569), .B(
        DP_OP_425J2_127_3477_n1567), .CI(DP_OP_425J2_127_3477_n1571), .CO(
        DP_OP_425J2_127_3477_n1480), .S(DP_OP_425J2_127_3477_n1481) );
  FADDX1_HVT DP_OP_425J2_127_3477_U922 ( .A(DP_OP_425J2_127_3477_n1565), .B(
        DP_OP_425J2_127_3477_n1545), .CI(DP_OP_425J2_127_3477_n1549), .CO(
        DP_OP_425J2_127_3477_n1478), .S(DP_OP_425J2_127_3477_n1479) );
  FADDX1_HVT DP_OP_425J2_127_3477_U921 ( .A(DP_OP_425J2_127_3477_n1547), .B(
        DP_OP_425J2_127_3477_n1555), .CI(DP_OP_425J2_127_3477_n1553), .CO(
        DP_OP_425J2_127_3477_n1476), .S(DP_OP_425J2_127_3477_n1477) );
  FADDX1_HVT DP_OP_425J2_127_3477_U920 ( .A(DP_OP_425J2_127_3477_n1557), .B(
        DP_OP_425J2_127_3477_n1535), .CI(DP_OP_425J2_127_3477_n1529), .CO(
        DP_OP_425J2_127_3477_n1474), .S(DP_OP_425J2_127_3477_n1475) );
  FADDX1_HVT DP_OP_425J2_127_3477_U919 ( .A(DP_OP_425J2_127_3477_n1537), .B(
        DP_OP_425J2_127_3477_n1533), .CI(DP_OP_425J2_127_3477_n1527), .CO(
        DP_OP_425J2_127_3477_n1472), .S(DP_OP_425J2_127_3477_n1473) );
  FADDX1_HVT DP_OP_425J2_127_3477_U918 ( .A(DP_OP_425J2_127_3477_n1539), .B(
        DP_OP_425J2_127_3477_n1513), .CI(DP_OP_425J2_127_3477_n1511), .CO(
        DP_OP_425J2_127_3477_n1470), .S(DP_OP_425J2_127_3477_n1471) );
  FADDX1_HVT DP_OP_425J2_127_3477_U917 ( .A(DP_OP_425J2_127_3477_n1525), .B(
        DP_OP_425J2_127_3477_n1521), .CI(DP_OP_425J2_127_3477_n1523), .CO(
        DP_OP_425J2_127_3477_n1468), .S(DP_OP_425J2_127_3477_n1469) );
  FADDX1_HVT DP_OP_425J2_127_3477_U916 ( .A(DP_OP_425J2_127_3477_n1531), .B(
        DP_OP_425J2_127_3477_n1509), .CI(DP_OP_425J2_127_3477_n1517), .CO(
        DP_OP_425J2_127_3477_n1466), .S(DP_OP_425J2_127_3477_n1467) );
  FADDX1_HVT DP_OP_425J2_127_3477_U915 ( .A(DP_OP_425J2_127_3477_n1519), .B(
        DP_OP_425J2_127_3477_n1543), .CI(DP_OP_425J2_127_3477_n1551), .CO(
        DP_OP_425J2_127_3477_n1464), .S(DP_OP_425J2_127_3477_n1465) );
  FADDX1_HVT DP_OP_425J2_127_3477_U914 ( .A(DP_OP_425J2_127_3477_n1515), .B(
        DP_OP_425J2_127_3477_n1541), .CI(DP_OP_425J2_127_3477_n1658), .CO(
        DP_OP_425J2_127_3477_n1462), .S(DP_OP_425J2_127_3477_n1463) );
  FADDX1_HVT DP_OP_425J2_127_3477_U913 ( .A(DP_OP_425J2_127_3477_n1652), .B(
        DP_OP_425J2_127_3477_n1654), .CI(DP_OP_425J2_127_3477_n1656), .CO(
        DP_OP_425J2_127_3477_n1460), .S(DP_OP_425J2_127_3477_n1461) );
  FADDX1_HVT DP_OP_425J2_127_3477_U912 ( .A(DP_OP_425J2_127_3477_n1646), .B(
        DP_OP_425J2_127_3477_n1650), .CI(DP_OP_425J2_127_3477_n1644), .CO(
        DP_OP_425J2_127_3477_n1458), .S(DP_OP_425J2_127_3477_n1459) );
  FADDX1_HVT DP_OP_425J2_127_3477_U911 ( .A(DP_OP_425J2_127_3477_n1648), .B(
        DP_OP_425J2_127_3477_n1642), .CI(DP_OP_425J2_127_3477_n1503), .CO(
        DP_OP_425J2_127_3477_n1456), .S(DP_OP_425J2_127_3477_n1457) );
  FADDX1_HVT DP_OP_425J2_127_3477_U910 ( .A(DP_OP_425J2_127_3477_n1505), .B(
        DP_OP_425J2_127_3477_n1640), .CI(DP_OP_425J2_127_3477_n1636), .CO(
        DP_OP_425J2_127_3477_n1454), .S(DP_OP_425J2_127_3477_n1455) );
  FADDX1_HVT DP_OP_425J2_127_3477_U909 ( .A(DP_OP_425J2_127_3477_n1507), .B(
        DP_OP_425J2_127_3477_n1638), .CI(DP_OP_425J2_127_3477_n1634), .CO(
        DP_OP_425J2_127_3477_n1452), .S(DP_OP_425J2_127_3477_n1453) );
  FADDX1_HVT DP_OP_425J2_127_3477_U908 ( .A(DP_OP_425J2_127_3477_n1624), .B(
        DP_OP_425J2_127_3477_n1487), .CI(DP_OP_425J2_127_3477_n1499), .CO(
        DP_OP_425J2_127_3477_n1450), .S(DP_OP_425J2_127_3477_n1451) );
  FADDX1_HVT DP_OP_425J2_127_3477_U907 ( .A(DP_OP_425J2_127_3477_n1632), .B(
        DP_OP_425J2_127_3477_n1501), .CI(DP_OP_425J2_127_3477_n1497), .CO(
        DP_OP_425J2_127_3477_n1448), .S(DP_OP_425J2_127_3477_n1449) );
  FADDX1_HVT DP_OP_425J2_127_3477_U906 ( .A(DP_OP_425J2_127_3477_n1630), .B(
        DP_OP_425J2_127_3477_n1489), .CI(DP_OP_425J2_127_3477_n1491), .CO(
        DP_OP_425J2_127_3477_n1446), .S(DP_OP_425J2_127_3477_n1447) );
  FADDX1_HVT DP_OP_425J2_127_3477_U905 ( .A(DP_OP_425J2_127_3477_n1628), .B(
        DP_OP_425J2_127_3477_n1495), .CI(DP_OP_425J2_127_3477_n1493), .CO(
        DP_OP_425J2_127_3477_n1444), .S(DP_OP_425J2_127_3477_n1445) );
  FADDX1_HVT DP_OP_425J2_127_3477_U904 ( .A(DP_OP_425J2_127_3477_n1626), .B(
        DP_OP_425J2_127_3477_n1622), .CI(DP_OP_425J2_127_3477_n1483), .CO(
        DP_OP_425J2_127_3477_n1442), .S(DP_OP_425J2_127_3477_n1443) );
  FADDX1_HVT DP_OP_425J2_127_3477_U903 ( .A(DP_OP_425J2_127_3477_n1485), .B(
        DP_OP_425J2_127_3477_n1481), .CI(DP_OP_425J2_127_3477_n1479), .CO(
        DP_OP_425J2_127_3477_n1440), .S(DP_OP_425J2_127_3477_n1441) );
  FADDX1_HVT DP_OP_425J2_127_3477_U902 ( .A(DP_OP_425J2_127_3477_n1620), .B(
        DP_OP_425J2_127_3477_n1471), .CI(DP_OP_425J2_127_3477_n1469), .CO(
        DP_OP_425J2_127_3477_n1438), .S(DP_OP_425J2_127_3477_n1439) );
  FADDX1_HVT DP_OP_425J2_127_3477_U901 ( .A(DP_OP_425J2_127_3477_n1475), .B(
        DP_OP_425J2_127_3477_n1465), .CI(DP_OP_425J2_127_3477_n1467), .CO(
        DP_OP_425J2_127_3477_n1436), .S(DP_OP_425J2_127_3477_n1437) );
  FADDX1_HVT DP_OP_425J2_127_3477_U900 ( .A(DP_OP_425J2_127_3477_n1473), .B(
        DP_OP_425J2_127_3477_n1477), .CI(DP_OP_425J2_127_3477_n1618), .CO(
        DP_OP_425J2_127_3477_n1434), .S(DP_OP_425J2_127_3477_n1435) );
  FADDX1_HVT DP_OP_425J2_127_3477_U899 ( .A(DP_OP_425J2_127_3477_n1616), .B(
        DP_OP_425J2_127_3477_n1463), .CI(DP_OP_425J2_127_3477_n1614), .CO(
        DP_OP_425J2_127_3477_n1432), .S(DP_OP_425J2_127_3477_n1433) );
  FADDX1_HVT DP_OP_425J2_127_3477_U898 ( .A(DP_OP_425J2_127_3477_n1461), .B(
        DP_OP_425J2_127_3477_n1459), .CI(DP_OP_425J2_127_3477_n1612), .CO(
        DP_OP_425J2_127_3477_n1430), .S(DP_OP_425J2_127_3477_n1431) );
  FADDX1_HVT DP_OP_425J2_127_3477_U897 ( .A(DP_OP_425J2_127_3477_n1610), .B(
        DP_OP_425J2_127_3477_n1606), .CI(DP_OP_425J2_127_3477_n1608), .CO(
        DP_OP_425J2_127_3477_n1428), .S(DP_OP_425J2_127_3477_n1429) );
  FADDX1_HVT DP_OP_425J2_127_3477_U896 ( .A(DP_OP_425J2_127_3477_n1457), .B(
        DP_OP_425J2_127_3477_n1604), .CI(DP_OP_425J2_127_3477_n1602), .CO(
        DP_OP_425J2_127_3477_n1426), .S(DP_OP_425J2_127_3477_n1427) );
  FADDX1_HVT DP_OP_425J2_127_3477_U894 ( .A(DP_OP_425J2_127_3477_n1451), .B(
        DP_OP_425J2_127_3477_n1447), .CI(DP_OP_425J2_127_3477_n1443), .CO(
        DP_OP_425J2_127_3477_n1422), .S(DP_OP_425J2_127_3477_n1423) );
  FADDX1_HVT DP_OP_425J2_127_3477_U893 ( .A(DP_OP_425J2_127_3477_n1600), .B(
        DP_OP_425J2_127_3477_n1445), .CI(DP_OP_425J2_127_3477_n1598), .CO(
        DP_OP_425J2_127_3477_n1420), .S(DP_OP_425J2_127_3477_n1421) );
  FADDX1_HVT DP_OP_425J2_127_3477_U892 ( .A(DP_OP_425J2_127_3477_n1441), .B(
        DP_OP_425J2_127_3477_n1439), .CI(DP_OP_425J2_127_3477_n1437), .CO(
        DP_OP_425J2_127_3477_n1418), .S(DP_OP_425J2_127_3477_n1419) );
  FADDX1_HVT DP_OP_425J2_127_3477_U891 ( .A(DP_OP_425J2_127_3477_n1596), .B(
        DP_OP_425J2_127_3477_n1435), .CI(DP_OP_425J2_127_3477_n1594), .CO(
        DP_OP_425J2_127_3477_n1416), .S(DP_OP_425J2_127_3477_n1417) );
  FADDX1_HVT DP_OP_425J2_127_3477_U890 ( .A(DP_OP_425J2_127_3477_n1433), .B(
        DP_OP_425J2_127_3477_n1592), .CI(DP_OP_425J2_127_3477_n1590), .CO(
        DP_OP_425J2_127_3477_n1414), .S(DP_OP_425J2_127_3477_n1415) );
  FADDX1_HVT DP_OP_425J2_127_3477_U889 ( .A(DP_OP_425J2_127_3477_n1429), .B(
        DP_OP_425J2_127_3477_n1431), .CI(DP_OP_425J2_127_3477_n1588), .CO(
        DP_OP_425J2_127_3477_n1412), .S(DP_OP_425J2_127_3477_n1413) );
  FADDX1_HVT DP_OP_425J2_127_3477_U888 ( .A(DP_OP_425J2_127_3477_n1427), .B(
        DP_OP_425J2_127_3477_n1425), .CI(DP_OP_425J2_127_3477_n1586), .CO(
        DP_OP_425J2_127_3477_n1410), .S(DP_OP_425J2_127_3477_n1411) );
  FADDX1_HVT DP_OP_425J2_127_3477_U887 ( .A(DP_OP_425J2_127_3477_n1421), .B(
        DP_OP_425J2_127_3477_n1423), .CI(DP_OP_425J2_127_3477_n1584), .CO(
        DP_OP_425J2_127_3477_n1408), .S(DP_OP_425J2_127_3477_n1409) );
  FADDX1_HVT DP_OP_425J2_127_3477_U886 ( .A(DP_OP_425J2_127_3477_n1419), .B(
        DP_OP_425J2_127_3477_n1417), .CI(DP_OP_425J2_127_3477_n1582), .CO(
        DP_OP_425J2_127_3477_n1406), .S(DP_OP_425J2_127_3477_n1407) );
  FADDX1_HVT DP_OP_425J2_127_3477_U885 ( .A(DP_OP_425J2_127_3477_n1415), .B(
        DP_OP_425J2_127_3477_n1580), .CI(DP_OP_425J2_127_3477_n1413), .CO(
        DP_OP_425J2_127_3477_n1404), .S(DP_OP_425J2_127_3477_n1405) );
  FADDX1_HVT DP_OP_425J2_127_3477_U884 ( .A(DP_OP_425J2_127_3477_n1411), .B(
        DP_OP_425J2_127_3477_n1578), .CI(DP_OP_425J2_127_3477_n1409), .CO(
        DP_OP_425J2_127_3477_n1402), .S(DP_OP_425J2_127_3477_n1403) );
  FADDX1_HVT DP_OP_425J2_127_3477_U883 ( .A(DP_OP_425J2_127_3477_n1407), .B(
        DP_OP_425J2_127_3477_n1576), .CI(DP_OP_425J2_127_3477_n1405), .CO(
        DP_OP_425J2_127_3477_n1400), .S(DP_OP_425J2_127_3477_n1401) );
  HADDX1_HVT DP_OP_425J2_127_3477_U882 ( .A0(DP_OP_425J2_127_3477_n3030), .B0(
        DP_OP_425J2_127_3477_n1975), .C1(DP_OP_425J2_127_3477_n1398), .SO(
        DP_OP_425J2_127_3477_n1399) );
  FADDX1_HVT DP_OP_425J2_127_3477_U881 ( .A(DP_OP_425J2_127_3477_n2503), .B(
        DP_OP_425J2_127_3477_n2415), .CI(DP_OP_425J2_127_3477_n1931), .CO(
        DP_OP_425J2_127_3477_n1396), .S(DP_OP_425J2_127_3477_n1397) );
  FADDX1_HVT DP_OP_425J2_127_3477_U880 ( .A(DP_OP_425J2_127_3477_n2547), .B(
        DP_OP_425J2_127_3477_n2327), .CI(DP_OP_425J2_127_3477_n2371), .CO(
        DP_OP_425J2_127_3477_n1394), .S(DP_OP_425J2_127_3477_n1395) );
  FADDX1_HVT DP_OP_425J2_127_3477_U879 ( .A(DP_OP_425J2_127_3477_n2855), .B(
        DP_OP_425J2_127_3477_n2019), .CI(DP_OP_425J2_127_3477_n2107), .CO(
        DP_OP_425J2_127_3477_n1392), .S(DP_OP_425J2_127_3477_n1393) );
  FADDX1_HVT DP_OP_425J2_127_3477_U878 ( .A(DP_OP_425J2_127_3477_n2591), .B(
        DP_OP_425J2_127_3477_n2151), .CI(DP_OP_425J2_127_3477_n2679), .CO(
        DP_OP_425J2_127_3477_n1390), .S(DP_OP_425J2_127_3477_n1391) );
  FADDX1_HVT DP_OP_425J2_127_3477_U877 ( .A(DP_OP_425J2_127_3477_n2063), .B(
        DP_OP_425J2_127_3477_n2899), .CI(DP_OP_425J2_127_3477_n2195), .CO(
        DP_OP_425J2_127_3477_n1388), .S(DP_OP_425J2_127_3477_n1389) );
  FADDX1_HVT DP_OP_425J2_127_3477_U876 ( .A(DP_OP_425J2_127_3477_n2459), .B(
        DP_OP_425J2_127_3477_n2943), .CI(DP_OP_425J2_127_3477_n2767), .CO(
        DP_OP_425J2_127_3477_n1386), .S(DP_OP_425J2_127_3477_n1387) );
  FADDX1_HVT DP_OP_425J2_127_3477_U875 ( .A(DP_OP_425J2_127_3477_n2283), .B(
        DP_OP_425J2_127_3477_n2239), .CI(DP_OP_425J2_127_3477_n2723), .CO(
        DP_OP_425J2_127_3477_n1384), .S(DP_OP_425J2_127_3477_n1385) );
  FADDX1_HVT DP_OP_425J2_127_3477_U874 ( .A(DP_OP_425J2_127_3477_n2987), .B(
        DP_OP_425J2_127_3477_n2635), .CI(DP_OP_425J2_127_3477_n2811), .CO(
        DP_OP_425J2_127_3477_n1382), .S(DP_OP_425J2_127_3477_n1383) );
  FADDX1_HVT DP_OP_425J2_127_3477_U873 ( .A(DP_OP_425J2_127_3477_n2429), .B(
        DP_OP_425J2_127_3477_n3050), .CI(DP_OP_425J2_127_3477_n1982), .CO(
        DP_OP_425J2_127_3477_n1380), .S(DP_OP_425J2_127_3477_n1381) );
  FADDX1_HVT DP_OP_425J2_127_3477_U872 ( .A(DP_OP_425J2_127_3477_n2422), .B(
        DP_OP_425J2_127_3477_n1989), .CI(DP_OP_425J2_127_3477_n1996), .CO(
        DP_OP_425J2_127_3477_n1378), .S(DP_OP_425J2_127_3477_n1379) );
  FADDX1_HVT DP_OP_425J2_127_3477_U871 ( .A(DP_OP_425J2_127_3477_n2436), .B(
        DP_OP_425J2_127_3477_n2026), .CI(DP_OP_425J2_127_3477_n3043), .CO(
        DP_OP_425J2_127_3477_n1376), .S(DP_OP_425J2_127_3477_n1377) );
  FADDX1_HVT DP_OP_425J2_127_3477_U870 ( .A(DP_OP_425J2_127_3477_n2392), .B(
        DP_OP_425J2_127_3477_n3036), .CI(DP_OP_425J2_127_3477_n3008), .CO(
        DP_OP_425J2_127_3477_n1374), .S(DP_OP_425J2_127_3477_n1375) );
  FADDX1_HVT DP_OP_425J2_127_3477_U869 ( .A(DP_OP_425J2_127_3477_n2385), .B(
        DP_OP_425J2_127_3477_n3001), .CI(DP_OP_425J2_127_3477_n2994), .CO(
        DP_OP_425J2_127_3477_n1372), .S(DP_OP_425J2_127_3477_n1373) );
  FADDX1_HVT DP_OP_425J2_127_3477_U868 ( .A(DP_OP_425J2_127_3477_n2348), .B(
        DP_OP_425J2_127_3477_n2964), .CI(DP_OP_425J2_127_3477_n2957), .CO(
        DP_OP_425J2_127_3477_n1370), .S(DP_OP_425J2_127_3477_n1371) );
  FADDX1_HVT DP_OP_425J2_127_3477_U867 ( .A(DP_OP_425J2_127_3477_n2341), .B(
        DP_OP_425J2_127_3477_n2033), .CI(DP_OP_425J2_127_3477_n2950), .CO(
        DP_OP_425J2_127_3477_n1368), .S(DP_OP_425J2_127_3477_n1369) );
  FADDX1_HVT DP_OP_425J2_127_3477_U866 ( .A(DP_OP_425J2_127_3477_n2334), .B(
        DP_OP_425J2_127_3477_n2920), .CI(DP_OP_425J2_127_3477_n2913), .CO(
        DP_OP_425J2_127_3477_n1366), .S(DP_OP_425J2_127_3477_n1367) );
  FADDX1_HVT DP_OP_425J2_127_3477_U865 ( .A(DP_OP_425J2_127_3477_n2304), .B(
        DP_OP_425J2_127_3477_n2906), .CI(DP_OP_425J2_127_3477_n2040), .CO(
        DP_OP_425J2_127_3477_n1364), .S(DP_OP_425J2_127_3477_n1365) );
  FADDX1_HVT DP_OP_425J2_127_3477_U864 ( .A(DP_OP_425J2_127_3477_n2297), .B(
        DP_OP_425J2_127_3477_n2070), .CI(DP_OP_425J2_127_3477_n2077), .CO(
        DP_OP_425J2_127_3477_n1362), .S(DP_OP_425J2_127_3477_n1363) );
  FADDX1_HVT DP_OP_425J2_127_3477_U863 ( .A(DP_OP_425J2_127_3477_n2378), .B(
        DP_OP_425J2_127_3477_n2084), .CI(DP_OP_425J2_127_3477_n2876), .CO(
        DP_OP_425J2_127_3477_n1360), .S(DP_OP_425J2_127_3477_n1361) );
  FADDX1_HVT DP_OP_425J2_127_3477_U862 ( .A(DP_OP_425J2_127_3477_n2466), .B(
        DP_OP_425J2_127_3477_n2869), .CI(DP_OP_425J2_127_3477_n2114), .CO(
        DP_OP_425J2_127_3477_n1358), .S(DP_OP_425J2_127_3477_n1359) );
  FADDX1_HVT DP_OP_425J2_127_3477_U861 ( .A(DP_OP_425J2_127_3477_n2862), .B(
        DP_OP_425J2_127_3477_n2121), .CI(DP_OP_425J2_127_3477_n2128), .CO(
        DP_OP_425J2_127_3477_n1356), .S(DP_OP_425J2_127_3477_n1357) );
  FADDX1_HVT DP_OP_425J2_127_3477_U860 ( .A(DP_OP_425J2_127_3477_n2832), .B(
        DP_OP_425J2_127_3477_n2158), .CI(DP_OP_425J2_127_3477_n2165), .CO(
        DP_OP_425J2_127_3477_n1354), .S(DP_OP_425J2_127_3477_n1355) );
  FADDX1_HVT DP_OP_425J2_127_3477_U859 ( .A(DP_OP_425J2_127_3477_n2825), .B(
        DP_OP_425J2_127_3477_n2172), .CI(DP_OP_425J2_127_3477_n2202), .CO(
        DP_OP_425J2_127_3477_n1352), .S(DP_OP_425J2_127_3477_n1353) );
  FADDX1_HVT DP_OP_425J2_127_3477_U858 ( .A(DP_OP_425J2_127_3477_n2818), .B(
        DP_OP_425J2_127_3477_n2209), .CI(DP_OP_425J2_127_3477_n2216), .CO(
        DP_OP_425J2_127_3477_n1350), .S(DP_OP_425J2_127_3477_n1351) );
  FADDX1_HVT DP_OP_425J2_127_3477_U857 ( .A(DP_OP_425J2_127_3477_n2788), .B(
        DP_OP_425J2_127_3477_n2246), .CI(DP_OP_425J2_127_3477_n2253), .CO(
        DP_OP_425J2_127_3477_n1348), .S(DP_OP_425J2_127_3477_n1349) );
  FADDX1_HVT DP_OP_425J2_127_3477_U856 ( .A(DP_OP_425J2_127_3477_n2781), .B(
        DP_OP_425J2_127_3477_n2260), .CI(DP_OP_425J2_127_3477_n2290), .CO(
        DP_OP_425J2_127_3477_n1346), .S(DP_OP_425J2_127_3477_n1347) );
  FADDX1_HVT DP_OP_425J2_127_3477_U855 ( .A(DP_OP_425J2_127_3477_n2774), .B(
        DP_OP_425J2_127_3477_n2473), .CI(DP_OP_425J2_127_3477_n2480), .CO(
        DP_OP_425J2_127_3477_n1344), .S(DP_OP_425J2_127_3477_n1345) );
  FADDX1_HVT DP_OP_425J2_127_3477_U854 ( .A(DP_OP_425J2_127_3477_n2744), .B(
        DP_OP_425J2_127_3477_n2510), .CI(DP_OP_425J2_127_3477_n2517), .CO(
        DP_OP_425J2_127_3477_n1342), .S(DP_OP_425J2_127_3477_n1343) );
  FADDX1_HVT DP_OP_425J2_127_3477_U853 ( .A(DP_OP_425J2_127_3477_n2737), .B(
        DP_OP_425J2_127_3477_n2524), .CI(DP_OP_425J2_127_3477_n2554), .CO(
        DP_OP_425J2_127_3477_n1340), .S(DP_OP_425J2_127_3477_n1341) );
  FADDX1_HVT DP_OP_425J2_127_3477_U852 ( .A(DP_OP_425J2_127_3477_n2730), .B(
        DP_OP_425J2_127_3477_n2561), .CI(DP_OP_425J2_127_3477_n2568), .CO(
        DP_OP_425J2_127_3477_n1338), .S(DP_OP_425J2_127_3477_n1339) );
  FADDX1_HVT DP_OP_425J2_127_3477_U851 ( .A(DP_OP_425J2_127_3477_n2700), .B(
        DP_OP_425J2_127_3477_n2693), .CI(DP_OP_425J2_127_3477_n2686), .CO(
        DP_OP_425J2_127_3477_n1336), .S(DP_OP_425J2_127_3477_n1337) );
  FADDX1_HVT DP_OP_425J2_127_3477_U850 ( .A(DP_OP_425J2_127_3477_n2642), .B(
        DP_OP_425J2_127_3477_n2656), .CI(DP_OP_425J2_127_3477_n2598), .CO(
        DP_OP_425J2_127_3477_n1334), .S(DP_OP_425J2_127_3477_n1335) );
  FADDX1_HVT DP_OP_425J2_127_3477_U849 ( .A(DP_OP_425J2_127_3477_n2605), .B(
        DP_OP_425J2_127_3477_n2612), .CI(DP_OP_425J2_127_3477_n2649), .CO(
        DP_OP_425J2_127_3477_n1332), .S(DP_OP_425J2_127_3477_n1333) );
  FADDX1_HVT DP_OP_425J2_127_3477_U848 ( .A(DP_OP_425J2_127_3477_n1399), .B(
        DP_OP_425J2_127_3477_n1574), .CI(DP_OP_425J2_127_3477_n1564), .CO(
        DP_OP_425J2_127_3477_n1330), .S(DP_OP_425J2_127_3477_n1331) );
  FADDX1_HVT DP_OP_425J2_127_3477_U847 ( .A(DP_OP_425J2_127_3477_n1572), .B(
        DP_OP_425J2_127_3477_n1570), .CI(DP_OP_425J2_127_3477_n1568), .CO(
        DP_OP_425J2_127_3477_n1328), .S(DP_OP_425J2_127_3477_n1329) );
  FADDX1_HVT DP_OP_425J2_127_3477_U846 ( .A(DP_OP_425J2_127_3477_n1566), .B(
        DP_OP_425J2_127_3477_n1562), .CI(DP_OP_425J2_127_3477_n1558), .CO(
        DP_OP_425J2_127_3477_n1326), .S(DP_OP_425J2_127_3477_n1327) );
  FADDX1_HVT DP_OP_425J2_127_3477_U845 ( .A(DP_OP_425J2_127_3477_n1560), .B(
        DP_OP_425J2_127_3477_n1534), .CI(DP_OP_425J2_127_3477_n1532), .CO(
        DP_OP_425J2_127_3477_n1324), .S(DP_OP_425J2_127_3477_n1325) );
  FADDX1_HVT DP_OP_425J2_127_3477_U844 ( .A(DP_OP_425J2_127_3477_n1536), .B(
        DP_OP_425J2_127_3477_n1508), .CI(DP_OP_425J2_127_3477_n1556), .CO(
        DP_OP_425J2_127_3477_n1322), .S(DP_OP_425J2_127_3477_n1323) );
  FADDX1_HVT DP_OP_425J2_127_3477_U843 ( .A(DP_OP_425J2_127_3477_n1528), .B(
        DP_OP_425J2_127_3477_n1554), .CI(DP_OP_425J2_127_3477_n1552), .CO(
        DP_OP_425J2_127_3477_n1320), .S(DP_OP_425J2_127_3477_n1321) );
  FADDX1_HVT DP_OP_425J2_127_3477_U842 ( .A(DP_OP_425J2_127_3477_n1524), .B(
        DP_OP_425J2_127_3477_n1550), .CI(DP_OP_425J2_127_3477_n1548), .CO(
        DP_OP_425J2_127_3477_n1318), .S(DP_OP_425J2_127_3477_n1319) );
  FADDX1_HVT DP_OP_425J2_127_3477_U841 ( .A(DP_OP_425J2_127_3477_n1518), .B(
        DP_OP_425J2_127_3477_n1510), .CI(DP_OP_425J2_127_3477_n1512), .CO(
        DP_OP_425J2_127_3477_n1316), .S(DP_OP_425J2_127_3477_n1317) );
  FADDX1_HVT DP_OP_425J2_127_3477_U840 ( .A(DP_OP_425J2_127_3477_n1516), .B(
        DP_OP_425J2_127_3477_n1546), .CI(DP_OP_425J2_127_3477_n1544), .CO(
        DP_OP_425J2_127_3477_n1314), .S(DP_OP_425J2_127_3477_n1315) );
  FADDX1_HVT DP_OP_425J2_127_3477_U839 ( .A(DP_OP_425J2_127_3477_n1526), .B(
        DP_OP_425J2_127_3477_n1542), .CI(DP_OP_425J2_127_3477_n1514), .CO(
        DP_OP_425J2_127_3477_n1312), .S(DP_OP_425J2_127_3477_n1313) );
  FADDX1_HVT DP_OP_425J2_127_3477_U838 ( .A(DP_OP_425J2_127_3477_n1522), .B(
        DP_OP_425J2_127_3477_n1540), .CI(DP_OP_425J2_127_3477_n1538), .CO(
        DP_OP_425J2_127_3477_n1310), .S(DP_OP_425J2_127_3477_n1311) );
  FADDX1_HVT DP_OP_425J2_127_3477_U837 ( .A(DP_OP_425J2_127_3477_n1520), .B(
        DP_OP_425J2_127_3477_n1530), .CI(DP_OP_425J2_127_3477_n1389), .CO(
        DP_OP_425J2_127_3477_n1308), .S(DP_OP_425J2_127_3477_n1309) );
  FADDX1_HVT DP_OP_425J2_127_3477_U836 ( .A(DP_OP_425J2_127_3477_n1391), .B(
        DP_OP_425J2_127_3477_n1383), .CI(DP_OP_425J2_127_3477_n1385), .CO(
        DP_OP_425J2_127_3477_n1306), .S(DP_OP_425J2_127_3477_n1307) );
  FADDX1_HVT DP_OP_425J2_127_3477_U835 ( .A(DP_OP_425J2_127_3477_n1395), .B(
        DP_OP_425J2_127_3477_n1393), .CI(DP_OP_425J2_127_3477_n1397), .CO(
        DP_OP_425J2_127_3477_n1304), .S(DP_OP_425J2_127_3477_n1305) );
  FADDX1_HVT DP_OP_425J2_127_3477_U834 ( .A(DP_OP_425J2_127_3477_n1387), .B(
        DP_OP_425J2_127_3477_n1339), .CI(DP_OP_425J2_127_3477_n1337), .CO(
        DP_OP_425J2_127_3477_n1302), .S(DP_OP_425J2_127_3477_n1303) );
  FADDX1_HVT DP_OP_425J2_127_3477_U833 ( .A(DP_OP_425J2_127_3477_n1333), .B(
        DP_OP_425J2_127_3477_n1381), .CI(DP_OP_425J2_127_3477_n1379), .CO(
        DP_OP_425J2_127_3477_n1300), .S(DP_OP_425J2_127_3477_n1301) );
  FADDX1_HVT DP_OP_425J2_127_3477_U832 ( .A(DP_OP_425J2_127_3477_n1369), .B(
        DP_OP_425J2_127_3477_n1359), .CI(DP_OP_425J2_127_3477_n1365), .CO(
        DP_OP_425J2_127_3477_n1298), .S(DP_OP_425J2_127_3477_n1299) );
  FADDX1_HVT DP_OP_425J2_127_3477_U831 ( .A(DP_OP_425J2_127_3477_n1363), .B(
        DP_OP_425J2_127_3477_n1361), .CI(DP_OP_425J2_127_3477_n1345), .CO(
        DP_OP_425J2_127_3477_n1296), .S(DP_OP_425J2_127_3477_n1297) );
  FADDX1_HVT DP_OP_425J2_127_3477_U830 ( .A(DP_OP_425J2_127_3477_n1367), .B(
        DP_OP_425J2_127_3477_n1341), .CI(DP_OP_425J2_127_3477_n1335), .CO(
        DP_OP_425J2_127_3477_n1294), .S(DP_OP_425J2_127_3477_n1295) );
  FADDX1_HVT DP_OP_425J2_127_3477_U829 ( .A(DP_OP_425J2_127_3477_n1371), .B(
        DP_OP_425J2_127_3477_n1353), .CI(DP_OP_425J2_127_3477_n1355), .CO(
        DP_OP_425J2_127_3477_n1292), .S(DP_OP_425J2_127_3477_n1293) );
  FADDX1_HVT DP_OP_425J2_127_3477_U828 ( .A(DP_OP_425J2_127_3477_n1351), .B(
        DP_OP_425J2_127_3477_n1349), .CI(DP_OP_425J2_127_3477_n1343), .CO(
        DP_OP_425J2_127_3477_n1290), .S(DP_OP_425J2_127_3477_n1291) );
  FADDX1_HVT DP_OP_425J2_127_3477_U827 ( .A(DP_OP_425J2_127_3477_n1347), .B(
        DP_OP_425J2_127_3477_n1377), .CI(DP_OP_425J2_127_3477_n1373), .CO(
        DP_OP_425J2_127_3477_n1288), .S(DP_OP_425J2_127_3477_n1289) );
  FADDX1_HVT DP_OP_425J2_127_3477_U826 ( .A(DP_OP_425J2_127_3477_n1375), .B(
        DP_OP_425J2_127_3477_n1357), .CI(DP_OP_425J2_127_3477_n1506), .CO(
        DP_OP_425J2_127_3477_n1286), .S(DP_OP_425J2_127_3477_n1287) );
  FADDX1_HVT DP_OP_425J2_127_3477_U825 ( .A(DP_OP_425J2_127_3477_n1504), .B(
        DP_OP_425J2_127_3477_n1502), .CI(DP_OP_425J2_127_3477_n1500), .CO(
        DP_OP_425J2_127_3477_n1284), .S(DP_OP_425J2_127_3477_n1285) );
  FADDX1_HVT DP_OP_425J2_127_3477_U824 ( .A(DP_OP_425J2_127_3477_n1498), .B(
        DP_OP_425J2_127_3477_n1486), .CI(DP_OP_425J2_127_3477_n1488), .CO(
        DP_OP_425J2_127_3477_n1282), .S(DP_OP_425J2_127_3477_n1283) );
  FADDX1_HVT DP_OP_425J2_127_3477_U823 ( .A(DP_OP_425J2_127_3477_n1492), .B(
        DP_OP_425J2_127_3477_n1496), .CI(DP_OP_425J2_127_3477_n1490), .CO(
        DP_OP_425J2_127_3477_n1280), .S(DP_OP_425J2_127_3477_n1281) );
  FADDX1_HVT DP_OP_425J2_127_3477_U822 ( .A(DP_OP_425J2_127_3477_n1494), .B(
        DP_OP_425J2_127_3477_n1331), .CI(DP_OP_425J2_127_3477_n1484), .CO(
        DP_OP_425J2_127_3477_n1278), .S(DP_OP_425J2_127_3477_n1279) );
  FADDX1_HVT DP_OP_425J2_127_3477_U821 ( .A(DP_OP_425J2_127_3477_n1329), .B(
        DP_OP_425J2_127_3477_n1327), .CI(DP_OP_425J2_127_3477_n1325), .CO(
        DP_OP_425J2_127_3477_n1276), .S(DP_OP_425J2_127_3477_n1277) );
  FADDX1_HVT DP_OP_425J2_127_3477_U820 ( .A(DP_OP_425J2_127_3477_n1482), .B(
        DP_OP_425J2_127_3477_n1480), .CI(DP_OP_425J2_127_3477_n1478), .CO(
        DP_OP_425J2_127_3477_n1274), .S(DP_OP_425J2_127_3477_n1275) );
  FADDX1_HVT DP_OP_425J2_127_3477_U819 ( .A(DP_OP_425J2_127_3477_n1466), .B(
        DP_OP_425J2_127_3477_n1311), .CI(DP_OP_425J2_127_3477_n1309), .CO(
        DP_OP_425J2_127_3477_n1272), .S(DP_OP_425J2_127_3477_n1273) );
  FADDX1_HVT DP_OP_425J2_127_3477_U818 ( .A(DP_OP_425J2_127_3477_n1476), .B(
        DP_OP_425J2_127_3477_n1321), .CI(DP_OP_425J2_127_3477_n1323), .CO(
        DP_OP_425J2_127_3477_n1270), .S(DP_OP_425J2_127_3477_n1271) );
  FADDX1_HVT DP_OP_425J2_127_3477_U817 ( .A(DP_OP_425J2_127_3477_n1474), .B(
        DP_OP_425J2_127_3477_n1317), .CI(DP_OP_425J2_127_3477_n1313), .CO(
        DP_OP_425J2_127_3477_n1268), .S(DP_OP_425J2_127_3477_n1269) );
  FADDX1_HVT DP_OP_425J2_127_3477_U816 ( .A(DP_OP_425J2_127_3477_n1472), .B(
        DP_OP_425J2_127_3477_n1319), .CI(DP_OP_425J2_127_3477_n1315), .CO(
        DP_OP_425J2_127_3477_n1266), .S(DP_OP_425J2_127_3477_n1267) );
  FADDX1_HVT DP_OP_425J2_127_3477_U815 ( .A(DP_OP_425J2_127_3477_n1470), .B(
        DP_OP_425J2_127_3477_n1464), .CI(DP_OP_425J2_127_3477_n1468), .CO(
        DP_OP_425J2_127_3477_n1264), .S(DP_OP_425J2_127_3477_n1265) );
  FADDX1_HVT DP_OP_425J2_127_3477_U814 ( .A(DP_OP_425J2_127_3477_n1305), .B(
        DP_OP_425J2_127_3477_n1307), .CI(DP_OP_425J2_127_3477_n1303), .CO(
        DP_OP_425J2_127_3477_n1262), .S(DP_OP_425J2_127_3477_n1263) );
  FADDX1_HVT DP_OP_425J2_127_3477_U813 ( .A(DP_OP_425J2_127_3477_n1295), .B(
        DP_OP_425J2_127_3477_n1297), .CI(DP_OP_425J2_127_3477_n1462), .CO(
        DP_OP_425J2_127_3477_n1260), .S(DP_OP_425J2_127_3477_n1261) );
  FADDX1_HVT DP_OP_425J2_127_3477_U812 ( .A(DP_OP_425J2_127_3477_n1293), .B(
        DP_OP_425J2_127_3477_n1301), .CI(DP_OP_425J2_127_3477_n1299), .CO(
        DP_OP_425J2_127_3477_n1258), .S(DP_OP_425J2_127_3477_n1259) );
  FADDX1_HVT DP_OP_425J2_127_3477_U811 ( .A(DP_OP_425J2_127_3477_n1289), .B(
        DP_OP_425J2_127_3477_n1291), .CI(DP_OP_425J2_127_3477_n1458), .CO(
        DP_OP_425J2_127_3477_n1256), .S(DP_OP_425J2_127_3477_n1257) );
  FADDX1_HVT DP_OP_425J2_127_3477_U810 ( .A(DP_OP_425J2_127_3477_n1287), .B(
        DP_OP_425J2_127_3477_n1460), .CI(DP_OP_425J2_127_3477_n1456), .CO(
        DP_OP_425J2_127_3477_n1254), .S(DP_OP_425J2_127_3477_n1255) );
  FADDX1_HVT DP_OP_425J2_127_3477_U809 ( .A(DP_OP_425J2_127_3477_n1454), .B(
        DP_OP_425J2_127_3477_n1452), .CI(DP_OP_425J2_127_3477_n1285), .CO(
        DP_OP_425J2_127_3477_n1252), .S(DP_OP_425J2_127_3477_n1253) );
  FADDX1_HVT DP_OP_425J2_127_3477_U808 ( .A(DP_OP_425J2_127_3477_n1450), .B(
        DP_OP_425J2_127_3477_n1442), .CI(DP_OP_425J2_127_3477_n1279), .CO(
        DP_OP_425J2_127_3477_n1250), .S(DP_OP_425J2_127_3477_n1251) );
  FADDX1_HVT DP_OP_425J2_127_3477_U807 ( .A(DP_OP_425J2_127_3477_n1448), .B(
        DP_OP_425J2_127_3477_n1281), .CI(DP_OP_425J2_127_3477_n1283), .CO(
        DP_OP_425J2_127_3477_n1248), .S(DP_OP_425J2_127_3477_n1249) );
  FADDX1_HVT DP_OP_425J2_127_3477_U806 ( .A(DP_OP_425J2_127_3477_n1446), .B(
        DP_OP_425J2_127_3477_n1444), .CI(DP_OP_425J2_127_3477_n1440), .CO(
        DP_OP_425J2_127_3477_n1246), .S(DP_OP_425J2_127_3477_n1247) );
  FADDX1_HVT DP_OP_425J2_127_3477_U805 ( .A(DP_OP_425J2_127_3477_n1275), .B(
        DP_OP_425J2_127_3477_n1277), .CI(DP_OP_425J2_127_3477_n1438), .CO(
        DP_OP_425J2_127_3477_n1244), .S(DP_OP_425J2_127_3477_n1245) );
  FADDX1_HVT DP_OP_425J2_127_3477_U804 ( .A(DP_OP_425J2_127_3477_n1436), .B(
        DP_OP_425J2_127_3477_n1269), .CI(DP_OP_425J2_127_3477_n1434), .CO(
        DP_OP_425J2_127_3477_n1242), .S(DP_OP_425J2_127_3477_n1243) );
  FADDX1_HVT DP_OP_425J2_127_3477_U803 ( .A(DP_OP_425J2_127_3477_n1267), .B(
        DP_OP_425J2_127_3477_n1273), .CI(DP_OP_425J2_127_3477_n1271), .CO(
        DP_OP_425J2_127_3477_n1240), .S(DP_OP_425J2_127_3477_n1241) );
  FADDX1_HVT DP_OP_425J2_127_3477_U802 ( .A(DP_OP_425J2_127_3477_n1265), .B(
        DP_OP_425J2_127_3477_n1263), .CI(DP_OP_425J2_127_3477_n1259), .CO(
        DP_OP_425J2_127_3477_n1238), .S(DP_OP_425J2_127_3477_n1239) );
  FADDX1_HVT DP_OP_425J2_127_3477_U801 ( .A(DP_OP_425J2_127_3477_n1261), .B(
        DP_OP_425J2_127_3477_n1432), .CI(DP_OP_425J2_127_3477_n1257), .CO(
        DP_OP_425J2_127_3477_n1236), .S(DP_OP_425J2_127_3477_n1237) );
  FADDX1_HVT DP_OP_425J2_127_3477_U800 ( .A(DP_OP_425J2_127_3477_n1430), .B(
        DP_OP_425J2_127_3477_n1428), .CI(DP_OP_425J2_127_3477_n1255), .CO(
        DP_OP_425J2_127_3477_n1234), .S(DP_OP_425J2_127_3477_n1235) );
  FADDX1_HVT DP_OP_425J2_127_3477_U799 ( .A(DP_OP_425J2_127_3477_n1426), .B(
        DP_OP_425J2_127_3477_n1253), .CI(DP_OP_425J2_127_3477_n1424), .CO(
        DP_OP_425J2_127_3477_n1232), .S(DP_OP_425J2_127_3477_n1233) );
  FADDX1_HVT DP_OP_425J2_127_3477_U798 ( .A(DP_OP_425J2_127_3477_n1422), .B(
        DP_OP_425J2_127_3477_n1249), .CI(DP_OP_425J2_127_3477_n1247), .CO(
        DP_OP_425J2_127_3477_n1230), .S(DP_OP_425J2_127_3477_n1231) );
  FADDX1_HVT DP_OP_425J2_127_3477_U797 ( .A(DP_OP_425J2_127_3477_n1420), .B(
        DP_OP_425J2_127_3477_n1251), .CI(DP_OP_425J2_127_3477_n1245), .CO(
        DP_OP_425J2_127_3477_n1228), .S(DP_OP_425J2_127_3477_n1229) );
  FADDX1_HVT DP_OP_425J2_127_3477_U796 ( .A(DP_OP_425J2_127_3477_n1418), .B(
        DP_OP_425J2_127_3477_n1241), .CI(DP_OP_425J2_127_3477_n1416), .CO(
        DP_OP_425J2_127_3477_n1226), .S(DP_OP_425J2_127_3477_n1227) );
  FADDX1_HVT DP_OP_425J2_127_3477_U795 ( .A(DP_OP_425J2_127_3477_n1243), .B(
        DP_OP_425J2_127_3477_n1239), .CI(DP_OP_425J2_127_3477_n1237), .CO(
        DP_OP_425J2_127_3477_n1224), .S(DP_OP_425J2_127_3477_n1225) );
  FADDX1_HVT DP_OP_425J2_127_3477_U794 ( .A(DP_OP_425J2_127_3477_n1414), .B(
        DP_OP_425J2_127_3477_n1235), .CI(DP_OP_425J2_127_3477_n1412), .CO(
        DP_OP_425J2_127_3477_n1222), .S(DP_OP_425J2_127_3477_n1223) );
  FADDX1_HVT DP_OP_425J2_127_3477_U793 ( .A(DP_OP_425J2_127_3477_n1233), .B(
        DP_OP_425J2_127_3477_n1410), .CI(DP_OP_425J2_127_3477_n1231), .CO(
        DP_OP_425J2_127_3477_n1220), .S(DP_OP_425J2_127_3477_n1221) );
  FADDX1_HVT DP_OP_425J2_127_3477_U792 ( .A(DP_OP_425J2_127_3477_n1229), .B(
        DP_OP_425J2_127_3477_n1408), .CI(DP_OP_425J2_127_3477_n1227), .CO(
        DP_OP_425J2_127_3477_n1218), .S(DP_OP_425J2_127_3477_n1219) );
  FADDX1_HVT DP_OP_425J2_127_3477_U791 ( .A(DP_OP_425J2_127_3477_n1406), .B(
        DP_OP_425J2_127_3477_n1225), .CI(DP_OP_425J2_127_3477_n1404), .CO(
        DP_OP_425J2_127_3477_n1216), .S(DP_OP_425J2_127_3477_n1217) );
  FADDX1_HVT DP_OP_425J2_127_3477_U790 ( .A(DP_OP_425J2_127_3477_n1223), .B(
        DP_OP_425J2_127_3477_n1221), .CI(DP_OP_425J2_127_3477_n1402), .CO(
        DP_OP_425J2_127_3477_n1214), .S(DP_OP_425J2_127_3477_n1215) );
  FADDX1_HVT DP_OP_425J2_127_3477_U789 ( .A(DP_OP_425J2_127_3477_n1219), .B(
        DP_OP_425J2_127_3477_n1217), .CI(DP_OP_425J2_127_3477_n1400), .CO(
        DP_OP_425J2_127_3477_n1212), .S(DP_OP_425J2_127_3477_n1213) );
  OR2X1_HVT DP_OP_425J2_127_3477_U788 ( .A1(DP_OP_425J2_127_3477_n3029), .A2(
        DP_OP_425J2_127_3477_n2502), .Y(DP_OP_425J2_127_3477_n1210) );
  FADDX1_HVT DP_OP_425J2_127_3477_U786 ( .A(DP_OP_425J2_127_3477_n2194), .B(
        DP_OP_425J2_127_3477_n1974), .CI(DP_OP_425J2_127_3477_n1930), .CO(
        DP_OP_425J2_127_3477_n1208), .S(DP_OP_425J2_127_3477_n1209) );
  FADDX1_HVT DP_OP_425J2_127_3477_U785 ( .A(DP_OP_425J2_127_3477_n2634), .B(
        DP_OP_425J2_127_3477_n2062), .CI(DP_OP_425J2_127_3477_n2414), .CO(
        DP_OP_425J2_127_3477_n1206), .S(DP_OP_425J2_127_3477_n1207) );
  FADDX1_HVT DP_OP_425J2_127_3477_U784 ( .A(DP_OP_425J2_127_3477_n2854), .B(
        DP_OP_425J2_127_3477_n2678), .CI(DP_OP_425J2_127_3477_n2238), .CO(
        DP_OP_425J2_127_3477_n1204), .S(DP_OP_425J2_127_3477_n1205) );
  FADDX1_HVT DP_OP_425J2_127_3477_U783 ( .A(DP_OP_425J2_127_3477_n2326), .B(
        DP_OP_425J2_127_3477_n2150), .CI(DP_OP_425J2_127_3477_n2898), .CO(
        DP_OP_425J2_127_3477_n1202), .S(DP_OP_425J2_127_3477_n1203) );
  FADDX1_HVT DP_OP_425J2_127_3477_U782 ( .A(DP_OP_425J2_127_3477_n2458), .B(
        DP_OP_425J2_127_3477_n2942), .CI(DP_OP_425J2_127_3477_n2722), .CO(
        DP_OP_425J2_127_3477_n1200), .S(DP_OP_425J2_127_3477_n1201) );
  FADDX1_HVT DP_OP_425J2_127_3477_U781 ( .A(DP_OP_425J2_127_3477_n2546), .B(
        DP_OP_425J2_127_3477_n2766), .CI(DP_OP_425J2_127_3477_n2590), .CO(
        DP_OP_425J2_127_3477_n1198), .S(DP_OP_425J2_127_3477_n1199) );
  FADDX1_HVT DP_OP_425J2_127_3477_U780 ( .A(DP_OP_425J2_127_3477_n2282), .B(
        DP_OP_425J2_127_3477_n2106), .CI(DP_OP_425J2_127_3477_n2986), .CO(
        DP_OP_425J2_127_3477_n1196), .S(DP_OP_425J2_127_3477_n1197) );
  FADDX1_HVT DP_OP_425J2_127_3477_U779 ( .A(DP_OP_425J2_127_3477_n2810), .B(
        DP_OP_425J2_127_3477_n2018), .CI(DP_OP_425J2_127_3477_n2370), .CO(
        DP_OP_425J2_127_3477_n1194), .S(DP_OP_425J2_127_3477_n1195) );
  FADDX1_HVT DP_OP_425J2_127_3477_U778 ( .A(DP_OP_425J2_127_3477_n2421), .B(
        DP_OP_425J2_127_3477_n3049), .CI(DP_OP_425J2_127_3477_n1981), .CO(
        DP_OP_425J2_127_3477_n1192), .S(DP_OP_425J2_127_3477_n1193) );
  FADDX1_HVT DP_OP_425J2_127_3477_U777 ( .A(DP_OP_425J2_127_3477_n2428), .B(
        DP_OP_425J2_127_3477_n3042), .CI(DP_OP_425J2_127_3477_n3035), .CO(
        DP_OP_425J2_127_3477_n1190), .S(DP_OP_425J2_127_3477_n1191) );
  FADDX1_HVT DP_OP_425J2_127_3477_U776 ( .A(DP_OP_425J2_127_3477_n2384), .B(
        DP_OP_425J2_127_3477_n3007), .CI(DP_OP_425J2_127_3477_n3000), .CO(
        DP_OP_425J2_127_3477_n1188), .S(DP_OP_425J2_127_3477_n1189) );
  FADDX1_HVT DP_OP_425J2_127_3477_U775 ( .A(DP_OP_425J2_127_3477_n2347), .B(
        DP_OP_425J2_127_3477_n2993), .CI(DP_OP_425J2_127_3477_n2963), .CO(
        DP_OP_425J2_127_3477_n1186), .S(DP_OP_425J2_127_3477_n1187) );
  FADDX1_HVT DP_OP_425J2_127_3477_U774 ( .A(DP_OP_425J2_127_3477_n2340), .B(
        DP_OP_425J2_127_3477_n1988), .CI(DP_OP_425J2_127_3477_n2956), .CO(
        DP_OP_425J2_127_3477_n1184), .S(DP_OP_425J2_127_3477_n1185) );
  FADDX1_HVT DP_OP_425J2_127_3477_U773 ( .A(DP_OP_425J2_127_3477_n2377), .B(
        DP_OP_425J2_127_3477_n2949), .CI(DP_OP_425J2_127_3477_n1995), .CO(
        DP_OP_425J2_127_3477_n1182), .S(DP_OP_425J2_127_3477_n1183) );
  FADDX1_HVT DP_OP_425J2_127_3477_U771 ( .A(DP_OP_425J2_127_3477_n2303), .B(
        DP_OP_425J2_127_3477_n2912), .CI(DP_OP_425J2_127_3477_n2905), .CO(
        DP_OP_425J2_127_3477_n1178), .S(DP_OP_425J2_127_3477_n1179) );
  FADDX1_HVT DP_OP_425J2_127_3477_U770 ( .A(DP_OP_425J2_127_3477_n2296), .B(
        DP_OP_425J2_127_3477_n2032), .CI(DP_OP_425J2_127_3477_n2875), .CO(
        DP_OP_425J2_127_3477_n1176), .S(DP_OP_425J2_127_3477_n1177) );
  FADDX1_HVT DP_OP_425J2_127_3477_U769 ( .A(DP_OP_425J2_127_3477_n2289), .B(
        DP_OP_425J2_127_3477_n2039), .CI(DP_OP_425J2_127_3477_n2868), .CO(
        DP_OP_425J2_127_3477_n1174), .S(DP_OP_425J2_127_3477_n1175) );
  FADDX1_HVT DP_OP_425J2_127_3477_U768 ( .A(DP_OP_425J2_127_3477_n2069), .B(
        DP_OP_425J2_127_3477_n2076), .CI(DP_OP_425J2_127_3477_n2083), .CO(
        DP_OP_425J2_127_3477_n1172), .S(DP_OP_425J2_127_3477_n1173) );
  FADDX1_HVT DP_OP_425J2_127_3477_U767 ( .A(DP_OP_425J2_127_3477_n2861), .B(
        DP_OP_425J2_127_3477_n2113), .CI(DP_OP_425J2_127_3477_n2120), .CO(
        DP_OP_425J2_127_3477_n1170), .S(DP_OP_425J2_127_3477_n1171) );
  FADDX1_HVT DP_OP_425J2_127_3477_U766 ( .A(DP_OP_425J2_127_3477_n2831), .B(
        DP_OP_425J2_127_3477_n2127), .CI(DP_OP_425J2_127_3477_n2157), .CO(
        DP_OP_425J2_127_3477_n1168), .S(DP_OP_425J2_127_3477_n1169) );
  FADDX1_HVT DP_OP_425J2_127_3477_U765 ( .A(DP_OP_425J2_127_3477_n2824), .B(
        DP_OP_425J2_127_3477_n2164), .CI(DP_OP_425J2_127_3477_n2171), .CO(
        DP_OP_425J2_127_3477_n1166), .S(DP_OP_425J2_127_3477_n1167) );
  FADDX1_HVT DP_OP_425J2_127_3477_U764 ( .A(DP_OP_425J2_127_3477_n2817), .B(
        DP_OP_425J2_127_3477_n2201), .CI(DP_OP_425J2_127_3477_n2208), .CO(
        DP_OP_425J2_127_3477_n1164), .S(DP_OP_425J2_127_3477_n1165) );
  FADDX1_HVT DP_OP_425J2_127_3477_U763 ( .A(DP_OP_425J2_127_3477_n2787), .B(
        DP_OP_425J2_127_3477_n2215), .CI(DP_OP_425J2_127_3477_n2245), .CO(
        DP_OP_425J2_127_3477_n1162), .S(DP_OP_425J2_127_3477_n1163) );
  FADDX1_HVT DP_OP_425J2_127_3477_U762 ( .A(DP_OP_425J2_127_3477_n2780), .B(
        DP_OP_425J2_127_3477_n2252), .CI(DP_OP_425J2_127_3477_n2259), .CO(
        DP_OP_425J2_127_3477_n1160), .S(DP_OP_425J2_127_3477_n1161) );
  FADDX1_HVT DP_OP_425J2_127_3477_U761 ( .A(DP_OP_425J2_127_3477_n2773), .B(
        DP_OP_425J2_127_3477_n2391), .CI(DP_OP_425J2_127_3477_n2435), .CO(
        DP_OP_425J2_127_3477_n1158), .S(DP_OP_425J2_127_3477_n1159) );
  FADDX1_HVT DP_OP_425J2_127_3477_U760 ( .A(DP_OP_425J2_127_3477_n2743), .B(
        DP_OP_425J2_127_3477_n2465), .CI(DP_OP_425J2_127_3477_n2472), .CO(
        DP_OP_425J2_127_3477_n1156), .S(DP_OP_425J2_127_3477_n1157) );
  FADDX1_HVT DP_OP_425J2_127_3477_U759 ( .A(DP_OP_425J2_127_3477_n2736), .B(
        DP_OP_425J2_127_3477_n2479), .CI(DP_OP_425J2_127_3477_n2509), .CO(
        DP_OP_425J2_127_3477_n1154), .S(DP_OP_425J2_127_3477_n1155) );
  FADDX1_HVT DP_OP_425J2_127_3477_U758 ( .A(DP_OP_425J2_127_3477_n2729), .B(
        DP_OP_425J2_127_3477_n2516), .CI(DP_OP_425J2_127_3477_n2523), .CO(
        DP_OP_425J2_127_3477_n1152), .S(DP_OP_425J2_127_3477_n1153) );
  FADDX1_HVT DP_OP_425J2_127_3477_U757 ( .A(DP_OP_425J2_127_3477_n2699), .B(
        DP_OP_425J2_127_3477_n2553), .CI(DP_OP_425J2_127_3477_n2560), .CO(
        DP_OP_425J2_127_3477_n1150), .S(DP_OP_425J2_127_3477_n1151) );
  FADDX1_HVT DP_OP_425J2_127_3477_U756 ( .A(DP_OP_425J2_127_3477_n2692), .B(
        DP_OP_425J2_127_3477_n2567), .CI(DP_OP_425J2_127_3477_n2597), .CO(
        DP_OP_425J2_127_3477_n1148), .S(DP_OP_425J2_127_3477_n1149) );
  FADDX1_HVT DP_OP_425J2_127_3477_U755 ( .A(DP_OP_425J2_127_3477_n2685), .B(
        DP_OP_425J2_127_3477_n2604), .CI(DP_OP_425J2_127_3477_n2611), .CO(
        DP_OP_425J2_127_3477_n1146), .S(DP_OP_425J2_127_3477_n1147) );
  FADDX1_HVT DP_OP_425J2_127_3477_U754 ( .A(DP_OP_425J2_127_3477_n2641), .B(
        DP_OP_425J2_127_3477_n2648), .CI(DP_OP_425J2_127_3477_n2655), .CO(
        DP_OP_425J2_127_3477_n1144), .S(DP_OP_425J2_127_3477_n1145) );
  FADDX1_HVT DP_OP_425J2_127_3477_U753 ( .A(DP_OP_425J2_127_3477_n1398), .B(
        DP_OP_425J2_127_3477_n1386), .CI(DP_OP_425J2_127_3477_n1384), .CO(
        DP_OP_425J2_127_3477_n1142), .S(DP_OP_425J2_127_3477_n1143) );
  FADDX1_HVT DP_OP_425J2_127_3477_U752 ( .A(DP_OP_425J2_127_3477_n1382), .B(
        DP_OP_425J2_127_3477_n1211), .CI(DP_OP_425J2_127_3477_n1388), .CO(
        DP_OP_425J2_127_3477_n1140), .S(DP_OP_425J2_127_3477_n1141) );
  FADDX1_HVT DP_OP_425J2_127_3477_U751 ( .A(DP_OP_425J2_127_3477_n1392), .B(
        DP_OP_425J2_127_3477_n1396), .CI(DP_OP_425J2_127_3477_n1390), .CO(
        DP_OP_425J2_127_3477_n1138), .S(DP_OP_425J2_127_3477_n1139) );
  FADDX1_HVT DP_OP_425J2_127_3477_U750 ( .A(DP_OP_425J2_127_3477_n1394), .B(
        DP_OP_425J2_127_3477_n1358), .CI(DP_OP_425J2_127_3477_n1356), .CO(
        DP_OP_425J2_127_3477_n1136), .S(DP_OP_425J2_127_3477_n1137) );
  FADDX1_HVT DP_OP_425J2_127_3477_U749 ( .A(DP_OP_425J2_127_3477_n1360), .B(
        DP_OP_425J2_127_3477_n1332), .CI(DP_OP_425J2_127_3477_n1380), .CO(
        DP_OP_425J2_127_3477_n1134), .S(DP_OP_425J2_127_3477_n1135) );
  FADDX1_HVT DP_OP_425J2_127_3477_U748 ( .A(DP_OP_425J2_127_3477_n1352), .B(
        DP_OP_425J2_127_3477_n1334), .CI(DP_OP_425J2_127_3477_n1378), .CO(
        DP_OP_425J2_127_3477_n1132), .S(DP_OP_425J2_127_3477_n1133) );
  FADDX1_HVT DP_OP_425J2_127_3477_U747 ( .A(DP_OP_425J2_127_3477_n1350), .B(
        DP_OP_425J2_127_3477_n1336), .CI(DP_OP_425J2_127_3477_n1376), .CO(
        DP_OP_425J2_127_3477_n1130), .S(DP_OP_425J2_127_3477_n1131) );
  FADDX1_HVT DP_OP_425J2_127_3477_U746 ( .A(DP_OP_425J2_127_3477_n1346), .B(
        DP_OP_425J2_127_3477_n1374), .CI(DP_OP_425J2_127_3477_n1372), .CO(
        DP_OP_425J2_127_3477_n1128), .S(DP_OP_425J2_127_3477_n1129) );
  FADDX1_HVT DP_OP_425J2_127_3477_U745 ( .A(DP_OP_425J2_127_3477_n1340), .B(
        DP_OP_425J2_127_3477_n1370), .CI(DP_OP_425J2_127_3477_n1368), .CO(
        DP_OP_425J2_127_3477_n1126), .S(DP_OP_425J2_127_3477_n1127) );
  FADDX1_HVT DP_OP_425J2_127_3477_U744 ( .A(DP_OP_425J2_127_3477_n1348), .B(
        DP_OP_425J2_127_3477_n1366), .CI(DP_OP_425J2_127_3477_n1364), .CO(
        DP_OP_425J2_127_3477_n1124), .S(DP_OP_425J2_127_3477_n1125) );
  FADDX1_HVT DP_OP_425J2_127_3477_U743 ( .A(DP_OP_425J2_127_3477_n1342), .B(
        DP_OP_425J2_127_3477_n1362), .CI(DP_OP_425J2_127_3477_n1354), .CO(
        DP_OP_425J2_127_3477_n1122), .S(DP_OP_425J2_127_3477_n1123) );
  FADDX1_HVT DP_OP_425J2_127_3477_U742 ( .A(DP_OP_425J2_127_3477_n1338), .B(
        DP_OP_425J2_127_3477_n1344), .CI(DP_OP_425J2_127_3477_n1201), .CO(
        DP_OP_425J2_127_3477_n1120), .S(DP_OP_425J2_127_3477_n1121) );
  FADDX1_HVT DP_OP_425J2_127_3477_U741 ( .A(DP_OP_425J2_127_3477_n1197), .B(
        DP_OP_425J2_127_3477_n1195), .CI(DP_OP_425J2_127_3477_n1199), .CO(
        DP_OP_425J2_127_3477_n1118), .S(DP_OP_425J2_127_3477_n1119) );
  FADDX1_HVT DP_OP_425J2_127_3477_U740 ( .A(DP_OP_425J2_127_3477_n1207), .B(
        DP_OP_425J2_127_3477_n1205), .CI(DP_OP_425J2_127_3477_n1209), .CO(
        DP_OP_425J2_127_3477_n1116), .S(DP_OP_425J2_127_3477_n1117) );
  FADDX1_HVT DP_OP_425J2_127_3477_U739 ( .A(DP_OP_425J2_127_3477_n1203), .B(
        DP_OP_425J2_127_3477_n1151), .CI(DP_OP_425J2_127_3477_n1153), .CO(
        DP_OP_425J2_127_3477_n1114), .S(DP_OP_425J2_127_3477_n1115) );
  FADDX1_HVT DP_OP_425J2_127_3477_U738 ( .A(DP_OP_425J2_127_3477_n1149), .B(
        DP_OP_425J2_127_3477_n1185), .CI(DP_OP_425J2_127_3477_n1181), .CO(
        DP_OP_425J2_127_3477_n1112), .S(DP_OP_425J2_127_3477_n1113) );
  FADDX1_HVT DP_OP_425J2_127_3477_U737 ( .A(DP_OP_425J2_127_3477_n1187), .B(
        DP_OP_425J2_127_3477_n1171), .CI(DP_OP_425J2_127_3477_n1177), .CO(
        DP_OP_425J2_127_3477_n1110), .S(DP_OP_425J2_127_3477_n1111) );
  FADDX1_HVT DP_OP_425J2_127_3477_U736 ( .A(DP_OP_425J2_127_3477_n1175), .B(
        DP_OP_425J2_127_3477_n1173), .CI(DP_OP_425J2_127_3477_n1157), .CO(
        DP_OP_425J2_127_3477_n1108), .S(DP_OP_425J2_127_3477_n1109) );
  FADDX1_HVT DP_OP_425J2_127_3477_U735 ( .A(DP_OP_425J2_127_3477_n1179), .B(
        DP_OP_425J2_127_3477_n1147), .CI(DP_OP_425J2_127_3477_n1145), .CO(
        DP_OP_425J2_127_3477_n1106), .S(DP_OP_425J2_127_3477_n1107) );
  FADDX1_HVT DP_OP_425J2_127_3477_U734 ( .A(DP_OP_425J2_127_3477_n1183), .B(
        DP_OP_425J2_127_3477_n1165), .CI(DP_OP_425J2_127_3477_n1167), .CO(
        DP_OP_425J2_127_3477_n1104), .S(DP_OP_425J2_127_3477_n1105) );
  FADDX1_HVT DP_OP_425J2_127_3477_U733 ( .A(DP_OP_425J2_127_3477_n1163), .B(
        DP_OP_425J2_127_3477_n1161), .CI(DP_OP_425J2_127_3477_n1155), .CO(
        DP_OP_425J2_127_3477_n1102), .S(DP_OP_425J2_127_3477_n1103) );
  FADDX1_HVT DP_OP_425J2_127_3477_U732 ( .A(DP_OP_425J2_127_3477_n1193), .B(
        DP_OP_425J2_127_3477_n1159), .CI(DP_OP_425J2_127_3477_n1191), .CO(
        DP_OP_425J2_127_3477_n1100), .S(DP_OP_425J2_127_3477_n1101) );
  FADDX1_HVT DP_OP_425J2_127_3477_U731 ( .A(DP_OP_425J2_127_3477_n1189), .B(
        DP_OP_425J2_127_3477_n1169), .CI(DP_OP_425J2_127_3477_n1330), .CO(
        DP_OP_425J2_127_3477_n1098), .S(DP_OP_425J2_127_3477_n1099) );
  FADDX1_HVT DP_OP_425J2_127_3477_U730 ( .A(DP_OP_425J2_127_3477_n1328), .B(
        DP_OP_425J2_127_3477_n1326), .CI(DP_OP_425J2_127_3477_n1324), .CO(
        DP_OP_425J2_127_3477_n1096), .S(DP_OP_425J2_127_3477_n1097) );
  FADDX1_HVT DP_OP_425J2_127_3477_U729 ( .A(DP_OP_425J2_127_3477_n1322), .B(
        DP_OP_425J2_127_3477_n1310), .CI(DP_OP_425J2_127_3477_n1308), .CO(
        DP_OP_425J2_127_3477_n1094), .S(DP_OP_425J2_127_3477_n1095) );
  FADDX1_HVT DP_OP_425J2_127_3477_U728 ( .A(DP_OP_425J2_127_3477_n1314), .B(
        DP_OP_425J2_127_3477_n1312), .CI(DP_OP_425J2_127_3477_n1320), .CO(
        DP_OP_425J2_127_3477_n1092), .S(DP_OP_425J2_127_3477_n1093) );
  FADDX1_HVT DP_OP_425J2_127_3477_U727 ( .A(DP_OP_425J2_127_3477_n1318), .B(
        DP_OP_425J2_127_3477_n1316), .CI(DP_OP_425J2_127_3477_n1143), .CO(
        DP_OP_425J2_127_3477_n1090), .S(DP_OP_425J2_127_3477_n1091) );
  FADDX1_HVT DP_OP_425J2_127_3477_U726 ( .A(DP_OP_425J2_127_3477_n1306), .B(
        DP_OP_425J2_127_3477_n1304), .CI(DP_OP_425J2_127_3477_n1137), .CO(
        DP_OP_425J2_127_3477_n1088), .S(DP_OP_425J2_127_3477_n1089) );
  FADDX1_HVT DP_OP_425J2_127_3477_U725 ( .A(DP_OP_425J2_127_3477_n1141), .B(
        DP_OP_425J2_127_3477_n1139), .CI(DP_OP_425J2_127_3477_n1302), .CO(
        DP_OP_425J2_127_3477_n1086), .S(DP_OP_425J2_127_3477_n1087) );
  FADDX1_HVT DP_OP_425J2_127_3477_U724 ( .A(DP_OP_425J2_127_3477_n1290), .B(
        DP_OP_425J2_127_3477_n1135), .CI(DP_OP_425J2_127_3477_n1121), .CO(
        DP_OP_425J2_127_3477_n1084), .S(DP_OP_425J2_127_3477_n1085) );
  FADDX1_HVT DP_OP_425J2_127_3477_U723 ( .A(DP_OP_425J2_127_3477_n1288), .B(
        DP_OP_425J2_127_3477_n1131), .CI(DP_OP_425J2_127_3477_n1133), .CO(
        DP_OP_425J2_127_3477_n1082), .S(DP_OP_425J2_127_3477_n1083) );
  FADDX1_HVT DP_OP_425J2_127_3477_U722 ( .A(DP_OP_425J2_127_3477_n1292), .B(
        DP_OP_425J2_127_3477_n1129), .CI(DP_OP_425J2_127_3477_n1127), .CO(
        DP_OP_425J2_127_3477_n1080), .S(DP_OP_425J2_127_3477_n1081) );
  FADDX1_HVT DP_OP_425J2_127_3477_U721 ( .A(DP_OP_425J2_127_3477_n1300), .B(
        DP_OP_425J2_127_3477_n1123), .CI(DP_OP_425J2_127_3477_n1125), .CO(
        DP_OP_425J2_127_3477_n1078), .S(DP_OP_425J2_127_3477_n1079) );
  FADDX1_HVT DP_OP_425J2_127_3477_U720 ( .A(DP_OP_425J2_127_3477_n1298), .B(
        DP_OP_425J2_127_3477_n1294), .CI(DP_OP_425J2_127_3477_n1296), .CO(
        DP_OP_425J2_127_3477_n1076), .S(DP_OP_425J2_127_3477_n1077) );
  FADDX1_HVT DP_OP_425J2_127_3477_U719 ( .A(DP_OP_425J2_127_3477_n1117), .B(
        DP_OP_425J2_127_3477_n1286), .CI(DP_OP_425J2_127_3477_n1115), .CO(
        DP_OP_425J2_127_3477_n1074), .S(DP_OP_425J2_127_3477_n1075) );
  FADDX1_HVT DP_OP_425J2_127_3477_U717 ( .A(DP_OP_425J2_127_3477_n1107), .B(
        DP_OP_425J2_127_3477_n1101), .CI(DP_OP_425J2_127_3477_n1284), .CO(
        DP_OP_425J2_127_3477_n1070), .S(DP_OP_425J2_127_3477_n1071) );
  FADDX1_HVT DP_OP_425J2_127_3477_U716 ( .A(DP_OP_425J2_127_3477_n1103), .B(
        DP_OP_425J2_127_3477_n1113), .CI(DP_OP_425J2_127_3477_n1105), .CO(
        DP_OP_425J2_127_3477_n1068), .S(DP_OP_425J2_127_3477_n1069) );
  FADDX1_HVT DP_OP_425J2_127_3477_U715 ( .A(DP_OP_425J2_127_3477_n1099), .B(
        DP_OP_425J2_127_3477_n1282), .CI(DP_OP_425J2_127_3477_n1278), .CO(
        DP_OP_425J2_127_3477_n1066), .S(DP_OP_425J2_127_3477_n1067) );
  FADDX1_HVT DP_OP_425J2_127_3477_U714 ( .A(DP_OP_425J2_127_3477_n1280), .B(
        DP_OP_425J2_127_3477_n1276), .CI(DP_OP_425J2_127_3477_n1274), .CO(
        DP_OP_425J2_127_3477_n1064), .S(DP_OP_425J2_127_3477_n1065) );
  FADDX1_HVT DP_OP_425J2_127_3477_U713 ( .A(DP_OP_425J2_127_3477_n1097), .B(
        DP_OP_425J2_127_3477_n1272), .CI(DP_OP_425J2_127_3477_n1270), .CO(
        DP_OP_425J2_127_3477_n1062), .S(DP_OP_425J2_127_3477_n1063) );
  FADDX1_HVT DP_OP_425J2_127_3477_U712 ( .A(DP_OP_425J2_127_3477_n1268), .B(
        DP_OP_425J2_127_3477_n1093), .CI(DP_OP_425J2_127_3477_n1091), .CO(
        DP_OP_425J2_127_3477_n1060), .S(DP_OP_425J2_127_3477_n1061) );
  FADDX1_HVT DP_OP_425J2_127_3477_U711 ( .A(DP_OP_425J2_127_3477_n1266), .B(
        DP_OP_425J2_127_3477_n1264), .CI(DP_OP_425J2_127_3477_n1095), .CO(
        DP_OP_425J2_127_3477_n1058), .S(DP_OP_425J2_127_3477_n1059) );
  FADDX1_HVT DP_OP_425J2_127_3477_U710 ( .A(DP_OP_425J2_127_3477_n1087), .B(
        DP_OP_425J2_127_3477_n1262), .CI(DP_OP_425J2_127_3477_n1089), .CO(
        DP_OP_425J2_127_3477_n1056), .S(DP_OP_425J2_127_3477_n1057) );
  FADDX1_HVT DP_OP_425J2_127_3477_U709 ( .A(DP_OP_425J2_127_3477_n1081), .B(
        DP_OP_425J2_127_3477_n1085), .CI(DP_OP_425J2_127_3477_n1256), .CO(
        DP_OP_425J2_127_3477_n1054), .S(DP_OP_425J2_127_3477_n1055) );
  FADDX1_HVT DP_OP_425J2_127_3477_U708 ( .A(DP_OP_425J2_127_3477_n1260), .B(
        DP_OP_425J2_127_3477_n1079), .CI(DP_OP_425J2_127_3477_n1083), .CO(
        DP_OP_425J2_127_3477_n1052), .S(DP_OP_425J2_127_3477_n1053) );
  FADDX1_HVT DP_OP_425J2_127_3477_U707 ( .A(DP_OP_425J2_127_3477_n1258), .B(
        DP_OP_425J2_127_3477_n1077), .CI(DP_OP_425J2_127_3477_n1254), .CO(
        DP_OP_425J2_127_3477_n1050), .S(DP_OP_425J2_127_3477_n1051) );
  FADDX1_HVT DP_OP_425J2_127_3477_U706 ( .A(DP_OP_425J2_127_3477_n1075), .B(
        DP_OP_425J2_127_3477_n1073), .CI(DP_OP_425J2_127_3477_n1071), .CO(
        DP_OP_425J2_127_3477_n1048), .S(DP_OP_425J2_127_3477_n1049) );
  FADDX1_HVT DP_OP_425J2_127_3477_U705 ( .A(DP_OP_425J2_127_3477_n1069), .B(
        DP_OP_425J2_127_3477_n1252), .CI(DP_OP_425J2_127_3477_n1067), .CO(
        DP_OP_425J2_127_3477_n1046), .S(DP_OP_425J2_127_3477_n1047) );
  FADDX1_HVT DP_OP_425J2_127_3477_U704 ( .A(DP_OP_425J2_127_3477_n1250), .B(
        DP_OP_425J2_127_3477_n1248), .CI(DP_OP_425J2_127_3477_n1246), .CO(
        DP_OP_425J2_127_3477_n1044), .S(DP_OP_425J2_127_3477_n1045) );
  FADDX1_HVT DP_OP_425J2_127_3477_U703 ( .A(DP_OP_425J2_127_3477_n1065), .B(
        DP_OP_425J2_127_3477_n1244), .CI(DP_OP_425J2_127_3477_n1063), .CO(
        DP_OP_425J2_127_3477_n1042), .S(DP_OP_425J2_127_3477_n1043) );
  FADDX1_HVT DP_OP_425J2_127_3477_U702 ( .A(DP_OP_425J2_127_3477_n1061), .B(
        DP_OP_425J2_127_3477_n1059), .CI(DP_OP_425J2_127_3477_n1242), .CO(
        DP_OP_425J2_127_3477_n1040), .S(DP_OP_425J2_127_3477_n1041) );
  FADDX1_HVT DP_OP_425J2_127_3477_U701 ( .A(DP_OP_425J2_127_3477_n1240), .B(
        DP_OP_425J2_127_3477_n1238), .CI(DP_OP_425J2_127_3477_n1057), .CO(
        DP_OP_425J2_127_3477_n1038), .S(DP_OP_425J2_127_3477_n1039) );
  FADDX1_HVT DP_OP_425J2_127_3477_U700 ( .A(DP_OP_425J2_127_3477_n1236), .B(
        DP_OP_425J2_127_3477_n1053), .CI(DP_OP_425J2_127_3477_n1051), .CO(
        DP_OP_425J2_127_3477_n1036), .S(DP_OP_425J2_127_3477_n1037) );
  FADDX1_HVT DP_OP_425J2_127_3477_U699 ( .A(DP_OP_425J2_127_3477_n1055), .B(
        DP_OP_425J2_127_3477_n1234), .CI(DP_OP_425J2_127_3477_n1049), .CO(
        DP_OP_425J2_127_3477_n1034), .S(DP_OP_425J2_127_3477_n1035) );
  FADDX1_HVT DP_OP_425J2_127_3477_U698 ( .A(DP_OP_425J2_127_3477_n1232), .B(
        DP_OP_425J2_127_3477_n1047), .CI(DP_OP_425J2_127_3477_n1230), .CO(
        DP_OP_425J2_127_3477_n1032), .S(DP_OP_425J2_127_3477_n1033) );
  FADDX1_HVT DP_OP_425J2_127_3477_U697 ( .A(DP_OP_425J2_127_3477_n1045), .B(
        DP_OP_425J2_127_3477_n1228), .CI(DP_OP_425J2_127_3477_n1043), .CO(
        DP_OP_425J2_127_3477_n1030), .S(DP_OP_425J2_127_3477_n1031) );
  FADDX1_HVT DP_OP_425J2_127_3477_U696 ( .A(DP_OP_425J2_127_3477_n1226), .B(
        DP_OP_425J2_127_3477_n1041), .CI(DP_OP_425J2_127_3477_n1039), .CO(
        DP_OP_425J2_127_3477_n1028), .S(DP_OP_425J2_127_3477_n1029) );
  FADDX1_HVT DP_OP_425J2_127_3477_U695 ( .A(DP_OP_425J2_127_3477_n1224), .B(
        DP_OP_425J2_127_3477_n1037), .CI(DP_OP_425J2_127_3477_n1222), .CO(
        DP_OP_425J2_127_3477_n1026), .S(DP_OP_425J2_127_3477_n1027) );
  FADDX1_HVT DP_OP_425J2_127_3477_U694 ( .A(DP_OP_425J2_127_3477_n1035), .B(
        DP_OP_425J2_127_3477_n1220), .CI(DP_OP_425J2_127_3477_n1033), .CO(
        DP_OP_425J2_127_3477_n1024), .S(DP_OP_425J2_127_3477_n1025) );
  FADDX1_HVT DP_OP_425J2_127_3477_U693 ( .A(DP_OP_425J2_127_3477_n1031), .B(
        DP_OP_425J2_127_3477_n1218), .CI(DP_OP_425J2_127_3477_n1029), .CO(
        DP_OP_425J2_127_3477_n1022), .S(DP_OP_425J2_127_3477_n1023) );
  FADDX1_HVT DP_OP_425J2_127_3477_U692 ( .A(DP_OP_425J2_127_3477_n1216), .B(
        DP_OP_425J2_127_3477_n1027), .CI(DP_OP_425J2_127_3477_n1025), .CO(
        DP_OP_425J2_127_3477_n1020), .S(DP_OP_425J2_127_3477_n1021) );
  FADDX1_HVT DP_OP_425J2_127_3477_U691 ( .A(DP_OP_425J2_127_3477_n1214), .B(
        DP_OP_425J2_127_3477_n1023), .CI(DP_OP_425J2_127_3477_n1212), .CO(
        DP_OP_425J2_127_3477_n1018), .S(DP_OP_425J2_127_3477_n1019) );
  FADDX1_HVT DP_OP_425J2_127_3477_U690 ( .A(DP_OP_425J2_127_3477_n3028), .B(
        DP_OP_425J2_127_3477_n1973), .CI(n1295), .CO(
        DP_OP_425J2_127_3477_n1016), .S(DP_OP_425J2_127_3477_n1017) );
  FADDX1_HVT DP_OP_425J2_127_3477_U689 ( .A(DP_OP_425J2_127_3477_n2853), .B(
        DP_OP_425J2_127_3477_n2170), .CI(DP_OP_425J2_127_3477_n2434), .CO(
        DP_OP_425J2_127_3477_n1014), .S(DP_OP_425J2_127_3477_n1015) );
  FADDX1_HVT DP_OP_425J2_127_3477_U688 ( .A(DP_OP_425J2_127_3477_n2061), .B(
        DP_OP_425J2_127_3477_n2478), .CI(DP_OP_425J2_127_3477_n2038), .CO(
        DP_OP_425J2_127_3477_n1012), .S(DP_OP_425J2_127_3477_n1013) );
  FADDX1_HVT DP_OP_425J2_127_3477_U687 ( .A(DP_OP_425J2_127_3477_n2369), .B(
        DP_OP_425J2_127_3477_n1994), .CI(DP_OP_425J2_127_3477_n2962), .CO(
        DP_OP_425J2_127_3477_n1010), .S(DP_OP_425J2_127_3477_n1011) );
  FADDX1_HVT DP_OP_425J2_127_3477_U686 ( .A(DP_OP_425J2_127_3477_n2325), .B(
        DP_OP_425J2_127_3477_n2302), .CI(DP_OP_425J2_127_3477_n2654), .CO(
        DP_OP_425J2_127_3477_n1008), .S(DP_OP_425J2_127_3477_n1009) );
  FADDX1_HVT DP_OP_425J2_127_3477_U685 ( .A(DP_OP_425J2_127_3477_n2237), .B(
        DP_OP_425J2_127_3477_n2346), .CI(DP_OP_425J2_127_3477_n3006), .CO(
        DP_OP_425J2_127_3477_n1006), .S(DP_OP_425J2_127_3477_n1007) );
  FADDX1_HVT DP_OP_425J2_127_3477_U684 ( .A(DP_OP_425J2_127_3477_n2017), .B(
        DP_OP_425J2_127_3477_n2082), .CI(DP_OP_425J2_127_3477_n2522), .CO(
        DP_OP_425J2_127_3477_n1004), .S(DP_OP_425J2_127_3477_n1005) );
  FADDX1_HVT DP_OP_425J2_127_3477_U683 ( .A(DP_OP_425J2_127_3477_n2105), .B(
        DP_OP_425J2_127_3477_n2786), .CI(DP_OP_425J2_127_3477_n2830), .CO(
        DP_OP_425J2_127_3477_n1002), .S(DP_OP_425J2_127_3477_n1003) );
  FADDX1_HVT DP_OP_425J2_127_3477_U682 ( .A(DP_OP_425J2_127_3477_n2193), .B(
        DP_OP_425J2_127_3477_n2742), .CI(DP_OP_425J2_127_3477_n2610), .CO(
        DP_OP_425J2_127_3477_n1000), .S(DP_OP_425J2_127_3477_n1001) );
  FADDX1_HVT DP_OP_425J2_127_3477_U681 ( .A(DP_OP_425J2_127_3477_n2545), .B(
        DP_OP_425J2_127_3477_n2390), .CI(DP_OP_425J2_127_3477_n2874), .CO(
        DP_OP_425J2_127_3477_n998), .S(DP_OP_425J2_127_3477_n999) );
  FADDX1_HVT DP_OP_425J2_127_3477_U680 ( .A(DP_OP_425J2_127_3477_n2941), .B(
        DP_OP_425J2_127_3477_n2214), .CI(DP_OP_425J2_127_3477_n2126), .CO(
        DP_OP_425J2_127_3477_n996), .S(DP_OP_425J2_127_3477_n997) );
  FADDX1_HVT DP_OP_425J2_127_3477_U679 ( .A(DP_OP_425J2_127_3477_n2677), .B(
        DP_OP_425J2_127_3477_n2918), .CI(DP_OP_425J2_127_3477_n2566), .CO(
        DP_OP_425J2_127_3477_n994), .S(DP_OP_425J2_127_3477_n995) );
  FADDX1_HVT DP_OP_425J2_127_3477_U678 ( .A(DP_OP_425J2_127_3477_n2457), .B(
        DP_OP_425J2_127_3477_n3048), .CI(DP_OP_425J2_127_3477_n2258), .CO(
        DP_OP_425J2_127_3477_n992), .S(DP_OP_425J2_127_3477_n993) );
  FADDX1_HVT DP_OP_425J2_127_3477_U677 ( .A(DP_OP_425J2_127_3477_n2149), .B(
        DP_OP_425J2_127_3477_n2413), .CI(DP_OP_425J2_127_3477_n2698), .CO(
        DP_OP_425J2_127_3477_n990), .S(DP_OP_425J2_127_3477_n991) );
  FADDX1_HVT DP_OP_425J2_127_3477_U676 ( .A(DP_OP_425J2_127_3477_n2765), .B(
        DP_OP_425J2_127_3477_n2809), .CI(DP_OP_425J2_127_3477_n2897), .CO(
        DP_OP_425J2_127_3477_n988), .S(DP_OP_425J2_127_3477_n989) );
  FADDX1_HVT DP_OP_425J2_127_3477_U675 ( .A(DP_OP_425J2_127_3477_n2501), .B(
        DP_OP_425J2_127_3477_n2589), .CI(DP_OP_425J2_127_3477_n2985), .CO(
        DP_OP_425J2_127_3477_n986), .S(DP_OP_425J2_127_3477_n987) );
  FADDX1_HVT DP_OP_425J2_127_3477_U674 ( .A(DP_OP_425J2_127_3477_n2633), .B(
        DP_OP_425J2_127_3477_n2281), .CI(DP_OP_425J2_127_3477_n2721), .CO(
        DP_OP_425J2_127_3477_n984), .S(DP_OP_425J2_127_3477_n985) );
  FADDX1_HVT DP_OP_425J2_127_3477_U673 ( .A(DP_OP_425J2_127_3477_n3041), .B(
        DP_OP_425J2_127_3477_n1987), .CI(DP_OP_425J2_127_3477_n1980), .CO(
        DP_OP_425J2_127_3477_n982), .S(DP_OP_425J2_127_3477_n983) );
  FADDX1_HVT DP_OP_425J2_127_3477_U672 ( .A(DP_OP_425J2_127_3477_n3034), .B(
        DP_OP_425J2_127_3477_n2999), .CI(DP_OP_425J2_127_3477_n2992), .CO(
        DP_OP_425J2_127_3477_n980), .S(DP_OP_425J2_127_3477_n981) );
  FADDX1_HVT DP_OP_425J2_127_3477_U671 ( .A(DP_OP_425J2_127_3477_n2515), .B(
        DP_OP_425J2_127_3477_n2955), .CI(DP_OP_425J2_127_3477_n2948), .CO(
        DP_OP_425J2_127_3477_n978), .S(DP_OP_425J2_127_3477_n979) );
  FADDX1_HVT DP_OP_425J2_127_3477_U670 ( .A(DP_OP_425J2_127_3477_n2911), .B(
        DP_OP_425J2_127_3477_n2024), .CI(DP_OP_425J2_127_3477_n2031), .CO(
        DP_OP_425J2_127_3477_n976), .S(DP_OP_425J2_127_3477_n977) );
  FADDX1_HVT DP_OP_425J2_127_3477_U669 ( .A(DP_OP_425J2_127_3477_n2904), .B(
        DP_OP_425J2_127_3477_n2068), .CI(DP_OP_425J2_127_3477_n2075), .CO(
        DP_OP_425J2_127_3477_n974), .S(DP_OP_425J2_127_3477_n975) );
  FADDX1_HVT DP_OP_425J2_127_3477_U668 ( .A(DP_OP_425J2_127_3477_n2867), .B(
        DP_OP_425J2_127_3477_n2112), .CI(DP_OP_425J2_127_3477_n2119), .CO(
        DP_OP_425J2_127_3477_n972), .S(DP_OP_425J2_127_3477_n973) );
  FADDX1_HVT DP_OP_425J2_127_3477_U667 ( .A(DP_OP_425J2_127_3477_n2860), .B(
        DP_OP_425J2_127_3477_n2156), .CI(DP_OP_425J2_127_3477_n2163), .CO(
        DP_OP_425J2_127_3477_n970), .S(DP_OP_425J2_127_3477_n971) );
  FADDX1_HVT DP_OP_425J2_127_3477_U666 ( .A(DP_OP_425J2_127_3477_n2823), .B(
        DP_OP_425J2_127_3477_n2200), .CI(DP_OP_425J2_127_3477_n2207), .CO(
        DP_OP_425J2_127_3477_n968), .S(DP_OP_425J2_127_3477_n969) );
  FADDX1_HVT DP_OP_425J2_127_3477_U665 ( .A(DP_OP_425J2_127_3477_n2816), .B(
        DP_OP_425J2_127_3477_n2244), .CI(DP_OP_425J2_127_3477_n2251), .CO(
        DP_OP_425J2_127_3477_n966), .S(DP_OP_425J2_127_3477_n967) );
  FADDX1_HVT DP_OP_425J2_127_3477_U664 ( .A(DP_OP_425J2_127_3477_n2779), .B(
        DP_OP_425J2_127_3477_n2288), .CI(DP_OP_425J2_127_3477_n2295), .CO(
        DP_OP_425J2_127_3477_n964), .S(DP_OP_425J2_127_3477_n965) );
  FADDX1_HVT DP_OP_425J2_127_3477_U663 ( .A(DP_OP_425J2_127_3477_n2772), .B(
        DP_OP_425J2_127_3477_n2332), .CI(DP_OP_425J2_127_3477_n2339), .CO(
        DP_OP_425J2_127_3477_n962), .S(DP_OP_425J2_127_3477_n963) );
  FADDX1_HVT DP_OP_425J2_127_3477_U662 ( .A(DP_OP_425J2_127_3477_n2735), .B(
        DP_OP_425J2_127_3477_n2376), .CI(DP_OP_425J2_127_3477_n2383), .CO(
        DP_OP_425J2_127_3477_n960), .S(DP_OP_425J2_127_3477_n961) );
  FADDX1_HVT DP_OP_425J2_127_3477_U661 ( .A(DP_OP_425J2_127_3477_n2728), .B(
        DP_OP_425J2_127_3477_n2420), .CI(DP_OP_425J2_127_3477_n2427), .CO(
        DP_OP_425J2_127_3477_n958), .S(DP_OP_425J2_127_3477_n959) );
  FADDX1_HVT DP_OP_425J2_127_3477_U660 ( .A(DP_OP_425J2_127_3477_n2691), .B(
        DP_OP_425J2_127_3477_n2464), .CI(DP_OP_425J2_127_3477_n2471), .CO(
        DP_OP_425J2_127_3477_n956), .S(DP_OP_425J2_127_3477_n957) );
  FADDX1_HVT DP_OP_425J2_127_3477_U659 ( .A(DP_OP_425J2_127_3477_n2684), .B(
        DP_OP_425J2_127_3477_n2508), .CI(DP_OP_425J2_127_3477_n2552), .CO(
        DP_OP_425J2_127_3477_n954), .S(DP_OP_425J2_127_3477_n955) );
  FADDX1_HVT DP_OP_425J2_127_3477_U658 ( .A(DP_OP_425J2_127_3477_n2647), .B(
        DP_OP_425J2_127_3477_n2559), .CI(DP_OP_425J2_127_3477_n2596), .CO(
        DP_OP_425J2_127_3477_n952), .S(DP_OP_425J2_127_3477_n953) );
  FADDX1_HVT DP_OP_425J2_127_3477_U657 ( .A(DP_OP_425J2_127_3477_n2640), .B(
        DP_OP_425J2_127_3477_n2603), .CI(DP_OP_425J2_127_3477_n1210), .CO(
        DP_OP_425J2_127_3477_n950), .S(DP_OP_425J2_127_3477_n951) );
  FADDX1_HVT DP_OP_425J2_127_3477_U656 ( .A(DP_OP_425J2_127_3477_n1198), .B(
        DP_OP_425J2_127_3477_n1194), .CI(DP_OP_425J2_127_3477_n1208), .CO(
        DP_OP_425J2_127_3477_n948), .S(DP_OP_425J2_127_3477_n949) );
  FADDX1_HVT DP_OP_425J2_127_3477_U655 ( .A(DP_OP_425J2_127_3477_n1206), .B(
        DP_OP_425J2_127_3477_n1196), .CI(DP_OP_425J2_127_3477_n1204), .CO(
        DP_OP_425J2_127_3477_n946), .S(DP_OP_425J2_127_3477_n947) );
  FADDX1_HVT DP_OP_425J2_127_3477_U654 ( .A(DP_OP_425J2_127_3477_n1202), .B(
        DP_OP_425J2_127_3477_n1200), .CI(DP_OP_425J2_127_3477_n1170), .CO(
        DP_OP_425J2_127_3477_n944), .S(DP_OP_425J2_127_3477_n945) );
  FADDX1_HVT DP_OP_425J2_127_3477_U653 ( .A(DP_OP_425J2_127_3477_n1168), .B(
        DP_OP_425J2_127_3477_n1144), .CI(DP_OP_425J2_127_3477_n1192), .CO(
        DP_OP_425J2_127_3477_n942), .S(DP_OP_425J2_127_3477_n943) );
  FADDX1_HVT DP_OP_425J2_127_3477_U652 ( .A(DP_OP_425J2_127_3477_n1166), .B(
        DP_OP_425J2_127_3477_n1190), .CI(DP_OP_425J2_127_3477_n1188), .CO(
        DP_OP_425J2_127_3477_n940), .S(DP_OP_425J2_127_3477_n941) );
  FADDX1_HVT DP_OP_425J2_127_3477_U651 ( .A(DP_OP_425J2_127_3477_n1160), .B(
        DP_OP_425J2_127_3477_n1186), .CI(DP_OP_425J2_127_3477_n1184), .CO(
        DP_OP_425J2_127_3477_n938), .S(DP_OP_425J2_127_3477_n939) );
  FADDX1_HVT DP_OP_425J2_127_3477_U650 ( .A(DP_OP_425J2_127_3477_n1182), .B(
        DP_OP_425J2_127_3477_n1180), .CI(DP_OP_425J2_127_3477_n1178), .CO(
        DP_OP_425J2_127_3477_n936), .S(DP_OP_425J2_127_3477_n937) );
  FADDX1_HVT DP_OP_425J2_127_3477_U649 ( .A(DP_OP_425J2_127_3477_n1150), .B(
        DP_OP_425J2_127_3477_n1176), .CI(DP_OP_425J2_127_3477_n1174), .CO(
        DP_OP_425J2_127_3477_n934), .S(DP_OP_425J2_127_3477_n935) );
  FADDX1_HVT DP_OP_425J2_127_3477_U648 ( .A(DP_OP_425J2_127_3477_n1156), .B(
        DP_OP_425J2_127_3477_n1172), .CI(DP_OP_425J2_127_3477_n1164), .CO(
        DP_OP_425J2_127_3477_n932), .S(DP_OP_425J2_127_3477_n933) );
  FADDX1_HVT DP_OP_425J2_127_3477_U647 ( .A(DP_OP_425J2_127_3477_n1148), .B(
        DP_OP_425J2_127_3477_n1162), .CI(DP_OP_425J2_127_3477_n1158), .CO(
        DP_OP_425J2_127_3477_n930), .S(DP_OP_425J2_127_3477_n931) );
  FADDX1_HVT DP_OP_425J2_127_3477_U646 ( .A(DP_OP_425J2_127_3477_n1152), .B(
        DP_OP_425J2_127_3477_n1146), .CI(DP_OP_425J2_127_3477_n1154), .CO(
        DP_OP_425J2_127_3477_n928), .S(DP_OP_425J2_127_3477_n929) );
  FADDX1_HVT DP_OP_425J2_127_3477_U645 ( .A(DP_OP_425J2_127_3477_n1017), .B(
        DP_OP_425J2_127_3477_n1003), .CI(DP_OP_425J2_127_3477_n1005), .CO(
        DP_OP_425J2_127_3477_n926), .S(DP_OP_425J2_127_3477_n927) );
  FADDX1_HVT DP_OP_425J2_127_3477_U644 ( .A(DP_OP_425J2_127_3477_n1009), .B(
        DP_OP_425J2_127_3477_n987), .CI(DP_OP_425J2_127_3477_n985), .CO(
        DP_OP_425J2_127_3477_n924), .S(DP_OP_425J2_127_3477_n925) );
  FADDX1_HVT DP_OP_425J2_127_3477_U643 ( .A(DP_OP_425J2_127_3477_n1001), .B(
        DP_OP_425J2_127_3477_n999), .CI(DP_OP_425J2_127_3477_n995), .CO(
        DP_OP_425J2_127_3477_n922), .S(DP_OP_425J2_127_3477_n923) );
  FADDX1_HVT DP_OP_425J2_127_3477_U642 ( .A(DP_OP_425J2_127_3477_n1007), .B(
        DP_OP_425J2_127_3477_n989), .CI(DP_OP_425J2_127_3477_n993), .CO(
        DP_OP_425J2_127_3477_n920), .S(DP_OP_425J2_127_3477_n921) );
  FADDX1_HVT DP_OP_425J2_127_3477_U641 ( .A(DP_OP_425J2_127_3477_n997), .B(
        DP_OP_425J2_127_3477_n1015), .CI(DP_OP_425J2_127_3477_n1011), .CO(
        DP_OP_425J2_127_3477_n918), .S(DP_OP_425J2_127_3477_n919) );
  FADDX1_HVT DP_OP_425J2_127_3477_U640 ( .A(DP_OP_425J2_127_3477_n991), .B(
        DP_OP_425J2_127_3477_n1013), .CI(DP_OP_425J2_127_3477_n973), .CO(
        DP_OP_425J2_127_3477_n916), .S(DP_OP_425J2_127_3477_n917) );
  FADDX1_HVT DP_OP_425J2_127_3477_U639 ( .A(DP_OP_425J2_127_3477_n975), .B(
        DP_OP_425J2_127_3477_n957), .CI(DP_OP_425J2_127_3477_n951), .CO(
        DP_OP_425J2_127_3477_n914), .S(DP_OP_425J2_127_3477_n915) );
  FADDX1_HVT DP_OP_425J2_127_3477_U638 ( .A(DP_OP_425J2_127_3477_n977), .B(
        DP_OP_425J2_127_3477_n953), .CI(DP_OP_425J2_127_3477_n969), .CO(
        DP_OP_425J2_127_3477_n912), .S(DP_OP_425J2_127_3477_n913) );
  FADDX1_HVT DP_OP_425J2_127_3477_U637 ( .A(DP_OP_425J2_127_3477_n967), .B(
        DP_OP_425J2_127_3477_n965), .CI(DP_OP_425J2_127_3477_n955), .CO(
        DP_OP_425J2_127_3477_n910), .S(DP_OP_425J2_127_3477_n911) );
  FADDX1_HVT DP_OP_425J2_127_3477_U636 ( .A(DP_OP_425J2_127_3477_n971), .B(
        DP_OP_425J2_127_3477_n959), .CI(DP_OP_425J2_127_3477_n961), .CO(
        DP_OP_425J2_127_3477_n908), .S(DP_OP_425J2_127_3477_n909) );
  FADDX1_HVT DP_OP_425J2_127_3477_U635 ( .A(DP_OP_425J2_127_3477_n983), .B(
        DP_OP_425J2_127_3477_n979), .CI(DP_OP_425J2_127_3477_n981), .CO(
        DP_OP_425J2_127_3477_n906), .S(DP_OP_425J2_127_3477_n907) );
  FADDX1_HVT DP_OP_425J2_127_3477_U634 ( .A(DP_OP_425J2_127_3477_n963), .B(
        DP_OP_425J2_127_3477_n1142), .CI(DP_OP_425J2_127_3477_n1140), .CO(
        DP_OP_425J2_127_3477_n904), .S(DP_OP_425J2_127_3477_n905) );
  FADDX1_HVT DP_OP_425J2_127_3477_U633 ( .A(DP_OP_425J2_127_3477_n1138), .B(
        DP_OP_425J2_127_3477_n1136), .CI(DP_OP_425J2_127_3477_n1122), .CO(
        DP_OP_425J2_127_3477_n902), .S(DP_OP_425J2_127_3477_n903) );
  FADDX1_HVT DP_OP_425J2_127_3477_U632 ( .A(DP_OP_425J2_127_3477_n1134), .B(
        DP_OP_425J2_127_3477_n1132), .CI(DP_OP_425J2_127_3477_n1120), .CO(
        DP_OP_425J2_127_3477_n900), .S(DP_OP_425J2_127_3477_n901) );
  FADDX1_HVT DP_OP_425J2_127_3477_U631 ( .A(DP_OP_425J2_127_3477_n1130), .B(
        DP_OP_425J2_127_3477_n1124), .CI(DP_OP_425J2_127_3477_n1126), .CO(
        DP_OP_425J2_127_3477_n898), .S(DP_OP_425J2_127_3477_n899) );
  FADDX1_HVT DP_OP_425J2_127_3477_U630 ( .A(DP_OP_425J2_127_3477_n1128), .B(
        DP_OP_425J2_127_3477_n1118), .CI(DP_OP_425J2_127_3477_n1116), .CO(
        DP_OP_425J2_127_3477_n896), .S(DP_OP_425J2_127_3477_n897) );
  FADDX1_HVT DP_OP_425J2_127_3477_U629 ( .A(DP_OP_425J2_127_3477_n949), .B(
        DP_OP_425J2_127_3477_n945), .CI(DP_OP_425J2_127_3477_n1114), .CO(
        DP_OP_425J2_127_3477_n894), .S(DP_OP_425J2_127_3477_n895) );
  FADDX1_HVT DP_OP_425J2_127_3477_U628 ( .A(DP_OP_425J2_127_3477_n947), .B(
        DP_OP_425J2_127_3477_n1102), .CI(DP_OP_425J2_127_3477_n1100), .CO(
        DP_OP_425J2_127_3477_n892), .S(DP_OP_425J2_127_3477_n893) );
  FADDX1_HVT DP_OP_425J2_127_3477_U627 ( .A(DP_OP_425J2_127_3477_n1108), .B(
        DP_OP_425J2_127_3477_n943), .CI(DP_OP_425J2_127_3477_n1098), .CO(
        DP_OP_425J2_127_3477_n890), .S(DP_OP_425J2_127_3477_n891) );
  FADDX1_HVT DP_OP_425J2_127_3477_U626 ( .A(DP_OP_425J2_127_3477_n1106), .B(
        DP_OP_425J2_127_3477_n939), .CI(DP_OP_425J2_127_3477_n929), .CO(
        DP_OP_425J2_127_3477_n888), .S(DP_OP_425J2_127_3477_n889) );
  FADDX1_HVT DP_OP_425J2_127_3477_U625 ( .A(DP_OP_425J2_127_3477_n1112), .B(
        DP_OP_425J2_127_3477_n935), .CI(DP_OP_425J2_127_3477_n937), .CO(
        DP_OP_425J2_127_3477_n886), .S(DP_OP_425J2_127_3477_n887) );
  FADDX1_HVT DP_OP_425J2_127_3477_U624 ( .A(DP_OP_425J2_127_3477_n1110), .B(
        DP_OP_425J2_127_3477_n931), .CI(DP_OP_425J2_127_3477_n933), .CO(
        DP_OP_425J2_127_3477_n884), .S(DP_OP_425J2_127_3477_n885) );
  FADDX1_HVT DP_OP_425J2_127_3477_U623 ( .A(DP_OP_425J2_127_3477_n1104), .B(
        DP_OP_425J2_127_3477_n941), .CI(DP_OP_425J2_127_3477_n927), .CO(
        DP_OP_425J2_127_3477_n882), .S(DP_OP_425J2_127_3477_n883) );
  FADDX1_HVT DP_OP_425J2_127_3477_U622 ( .A(DP_OP_425J2_127_3477_n921), .B(
        DP_OP_425J2_127_3477_n925), .CI(DP_OP_425J2_127_3477_n917), .CO(
        DP_OP_425J2_127_3477_n880), .S(DP_OP_425J2_127_3477_n881) );
  FADDX1_HVT DP_OP_425J2_127_3477_U621 ( .A(DP_OP_425J2_127_3477_n919), .B(
        DP_OP_425J2_127_3477_n923), .CI(DP_OP_425J2_127_3477_n911), .CO(
        DP_OP_425J2_127_3477_n878), .S(DP_OP_425J2_127_3477_n879) );
  FADDX1_HVT DP_OP_425J2_127_3477_U620 ( .A(DP_OP_425J2_127_3477_n909), .B(
        DP_OP_425J2_127_3477_n915), .CI(DP_OP_425J2_127_3477_n1096), .CO(
        DP_OP_425J2_127_3477_n876), .S(DP_OP_425J2_127_3477_n877) );
  FADDX1_HVT DP_OP_425J2_127_3477_U619 ( .A(DP_OP_425J2_127_3477_n907), .B(
        DP_OP_425J2_127_3477_n913), .CI(DP_OP_425J2_127_3477_n1092), .CO(
        DP_OP_425J2_127_3477_n874), .S(DP_OP_425J2_127_3477_n875) );
  FADDX1_HVT DP_OP_425J2_127_3477_U618 ( .A(DP_OP_425J2_127_3477_n905), .B(
        DP_OP_425J2_127_3477_n1090), .CI(DP_OP_425J2_127_3477_n1094), .CO(
        DP_OP_425J2_127_3477_n872), .S(DP_OP_425J2_127_3477_n873) );
  FADDX1_HVT DP_OP_425J2_127_3477_U617 ( .A(DP_OP_425J2_127_3477_n1086), .B(
        DP_OP_425J2_127_3477_n1088), .CI(DP_OP_425J2_127_3477_n903), .CO(
        DP_OP_425J2_127_3477_n870), .S(DP_OP_425J2_127_3477_n871) );
  FADDX1_HVT DP_OP_425J2_127_3477_U616 ( .A(DP_OP_425J2_127_3477_n1084), .B(
        DP_OP_425J2_127_3477_n901), .CI(DP_OP_425J2_127_3477_n899), .CO(
        DP_OP_425J2_127_3477_n868), .S(DP_OP_425J2_127_3477_n869) );
  FADDX1_HVT DP_OP_425J2_127_3477_U615 ( .A(DP_OP_425J2_127_3477_n1082), .B(
        DP_OP_425J2_127_3477_n1076), .CI(DP_OP_425J2_127_3477_n1078), .CO(
        DP_OP_425J2_127_3477_n866), .S(DP_OP_425J2_127_3477_n867) );
  FADDX1_HVT DP_OP_425J2_127_3477_U614 ( .A(DP_OP_425J2_127_3477_n1080), .B(
        DP_OP_425J2_127_3477_n897), .CI(DP_OP_425J2_127_3477_n1074), .CO(
        DP_OP_425J2_127_3477_n864), .S(DP_OP_425J2_127_3477_n865) );
  FADDX1_HVT DP_OP_425J2_127_3477_U613 ( .A(DP_OP_425J2_127_3477_n895), .B(
        DP_OP_425J2_127_3477_n1072), .CI(DP_OP_425J2_127_3477_n893), .CO(
        DP_OP_425J2_127_3477_n862), .S(DP_OP_425J2_127_3477_n863) );
  FADDX1_HVT DP_OP_425J2_127_3477_U612 ( .A(DP_OP_425J2_127_3477_n1070), .B(
        DP_OP_425J2_127_3477_n887), .CI(DP_OP_425J2_127_3477_n883), .CO(
        DP_OP_425J2_127_3477_n860), .S(DP_OP_425J2_127_3477_n861) );
  FADDX1_HVT DP_OP_425J2_127_3477_U611 ( .A(DP_OP_425J2_127_3477_n1068), .B(
        DP_OP_425J2_127_3477_n891), .CI(DP_OP_425J2_127_3477_n889), .CO(
        DP_OP_425J2_127_3477_n858), .S(DP_OP_425J2_127_3477_n859) );
  FADDX1_HVT DP_OP_425J2_127_3477_U610 ( .A(DP_OP_425J2_127_3477_n885), .B(
        DP_OP_425J2_127_3477_n881), .CI(DP_OP_425J2_127_3477_n1066), .CO(
        DP_OP_425J2_127_3477_n856), .S(DP_OP_425J2_127_3477_n857) );
  FADDX1_HVT DP_OP_425J2_127_3477_U609 ( .A(DP_OP_425J2_127_3477_n879), .B(
        DP_OP_425J2_127_3477_n877), .CI(DP_OP_425J2_127_3477_n1064), .CO(
        DP_OP_425J2_127_3477_n854), .S(DP_OP_425J2_127_3477_n855) );
  FADDX1_HVT DP_OP_425J2_127_3477_U608 ( .A(DP_OP_425J2_127_3477_n875), .B(
        DP_OP_425J2_127_3477_n1062), .CI(DP_OP_425J2_127_3477_n1058), .CO(
        DP_OP_425J2_127_3477_n852), .S(DP_OP_425J2_127_3477_n853) );
  FADDX1_HVT DP_OP_425J2_127_3477_U607 ( .A(DP_OP_425J2_127_3477_n1060), .B(
        DP_OP_425J2_127_3477_n873), .CI(DP_OP_425J2_127_3477_n1056), .CO(
        DP_OP_425J2_127_3477_n850), .S(DP_OP_425J2_127_3477_n851) );
  FADDX1_HVT DP_OP_425J2_127_3477_U606 ( .A(DP_OP_425J2_127_3477_n871), .B(
        DP_OP_425J2_127_3477_n1054), .CI(DP_OP_425J2_127_3477_n1052), .CO(
        DP_OP_425J2_127_3477_n848), .S(DP_OP_425J2_127_3477_n849) );
  FADDX1_HVT DP_OP_425J2_127_3477_U605 ( .A(DP_OP_425J2_127_3477_n869), .B(
        DP_OP_425J2_127_3477_n1050), .CI(DP_OP_425J2_127_3477_n865), .CO(
        DP_OP_425J2_127_3477_n846), .S(DP_OP_425J2_127_3477_n847) );
  FADDX1_HVT DP_OP_425J2_127_3477_U603 ( .A(DP_OP_425J2_127_3477_n1046), .B(
        DP_OP_425J2_127_3477_n861), .CI(DP_OP_425J2_127_3477_n857), .CO(
        DP_OP_425J2_127_3477_n842), .S(DP_OP_425J2_127_3477_n843) );
  FADDX1_HVT DP_OP_425J2_127_3477_U602 ( .A(DP_OP_425J2_127_3477_n859), .B(
        DP_OP_425J2_127_3477_n1044), .CI(DP_OP_425J2_127_3477_n855), .CO(
        DP_OP_425J2_127_3477_n840), .S(DP_OP_425J2_127_3477_n841) );
  FADDX1_HVT DP_OP_425J2_127_3477_U601 ( .A(DP_OP_425J2_127_3477_n1042), .B(
        DP_OP_425J2_127_3477_n853), .CI(DP_OP_425J2_127_3477_n1040), .CO(
        DP_OP_425J2_127_3477_n838), .S(DP_OP_425J2_127_3477_n839) );
  FADDX1_HVT DP_OP_425J2_127_3477_U600 ( .A(DP_OP_425J2_127_3477_n851), .B(
        DP_OP_425J2_127_3477_n849), .CI(DP_OP_425J2_127_3477_n1038), .CO(
        DP_OP_425J2_127_3477_n836), .S(DP_OP_425J2_127_3477_n837) );
  FADDX1_HVT DP_OP_425J2_127_3477_U599 ( .A(DP_OP_425J2_127_3477_n1036), .B(
        DP_OP_425J2_127_3477_n847), .CI(DP_OP_425J2_127_3477_n1034), .CO(
        DP_OP_425J2_127_3477_n834), .S(DP_OP_425J2_127_3477_n835) );
  FADDX1_HVT DP_OP_425J2_127_3477_U598 ( .A(DP_OP_425J2_127_3477_n845), .B(
        DP_OP_425J2_127_3477_n843), .CI(DP_OP_425J2_127_3477_n1032), .CO(
        DP_OP_425J2_127_3477_n832), .S(DP_OP_425J2_127_3477_n833) );
  FADDX1_HVT DP_OP_425J2_127_3477_U597 ( .A(DP_OP_425J2_127_3477_n841), .B(
        DP_OP_425J2_127_3477_n1030), .CI(DP_OP_425J2_127_3477_n839), .CO(
        DP_OP_425J2_127_3477_n830), .S(DP_OP_425J2_127_3477_n831) );
  FADDX1_HVT DP_OP_425J2_127_3477_U595 ( .A(DP_OP_425J2_127_3477_n835), .B(
        DP_OP_425J2_127_3477_n833), .CI(DP_OP_425J2_127_3477_n1024), .CO(
        DP_OP_425J2_127_3477_n826), .S(DP_OP_425J2_127_3477_n827) );
  FADDX1_HVT DP_OP_425J2_127_3477_U591 ( .A(DP_OP_425J2_127_3477_n2236), .B(
        DP_OP_425J2_127_3477_n1972), .CI(DP_OP_425J2_127_3477_n1928), .CO(
        DP_OP_425J2_127_3477_n818), .S(DP_OP_425J2_127_3477_n819) );
  FADDX1_HVT DP_OP_425J2_127_3477_U590 ( .A(DP_OP_425J2_127_3477_n2808), .B(
        DP_OP_425J2_127_3477_n2030), .CI(DP_OP_425J2_127_3477_n2294), .CO(
        DP_OP_425J2_127_3477_n816), .S(DP_OP_425J2_127_3477_n817) );
  FADDX1_HVT DP_OP_425J2_127_3477_U589 ( .A(DP_OP_425J2_127_3477_n2280), .B(
        DP_OP_425J2_127_3477_n3040), .CI(DP_OP_425J2_127_3477_n2690), .CO(
        DP_OP_425J2_127_3477_n814), .S(DP_OP_425J2_127_3477_n815) );
  FADDX1_HVT DP_OP_425J2_127_3477_U588 ( .A(DP_OP_425J2_127_3477_n2500), .B(
        DP_OP_425J2_127_3477_n2074), .CI(DP_OP_425J2_127_3477_n2118), .CO(
        DP_OP_425J2_127_3477_n812), .S(DP_OP_425J2_127_3477_n813) );
  FADDX1_HVT DP_OP_425J2_127_3477_U587 ( .A(DP_OP_425J2_127_3477_n2060), .B(
        DP_OP_425J2_127_3477_n2162), .CI(DP_OP_425J2_127_3477_n2206), .CO(
        DP_OP_425J2_127_3477_n810), .S(DP_OP_425J2_127_3477_n811) );
  FADDX1_HVT DP_OP_425J2_127_3477_U586 ( .A(DP_OP_425J2_127_3477_n2764), .B(
        DP_OP_425J2_127_3477_n2866), .CI(DP_OP_425J2_127_3477_n2910), .CO(
        DP_OP_425J2_127_3477_n808), .S(DP_OP_425J2_127_3477_n809) );
  FADDX1_HVT DP_OP_425J2_127_3477_U585 ( .A(DP_OP_425J2_127_3477_n2104), .B(
        DP_OP_425J2_127_3477_n2822), .CI(DP_OP_425J2_127_3477_n2646), .CO(
        DP_OP_425J2_127_3477_n806), .S(DP_OP_425J2_127_3477_n807) );
  FADDX1_HVT DP_OP_425J2_127_3477_U584 ( .A(DP_OP_425J2_127_3477_n2192), .B(
        DP_OP_425J2_127_3477_n2470), .CI(DP_OP_425J2_127_3477_n2998), .CO(
        DP_OP_425J2_127_3477_n804), .S(DP_OP_425J2_127_3477_n805) );
  FADDX1_HVT DP_OP_425J2_127_3477_U583 ( .A(DP_OP_425J2_127_3477_n2720), .B(
        DP_OP_425J2_127_3477_n2954), .CI(DP_OP_425J2_127_3477_n2514), .CO(
        DP_OP_425J2_127_3477_n802), .S(DP_OP_425J2_127_3477_n803) );
  FADDX1_HVT DP_OP_425J2_127_3477_U582 ( .A(DP_OP_425J2_127_3477_n2676), .B(
        DP_OP_425J2_127_3477_n2426), .CI(DP_OP_425J2_127_3477_n2778), .CO(
        DP_OP_425J2_127_3477_n800), .S(DP_OP_425J2_127_3477_n801) );
  FADDX1_HVT DP_OP_425J2_127_3477_U581 ( .A(DP_OP_425J2_127_3477_n2896), .B(
        DP_OP_425J2_127_3477_n2558), .CI(DP_OP_425J2_127_3477_n2382), .CO(
        DP_OP_425J2_127_3477_n798), .S(DP_OP_425J2_127_3477_n799) );
  FADDX1_HVT DP_OP_425J2_127_3477_U580 ( .A(DP_OP_425J2_127_3477_n2368), .B(
        DP_OP_425J2_127_3477_n2338), .CI(DP_OP_425J2_127_3477_n1986), .CO(
        DP_OP_425J2_127_3477_n796), .S(DP_OP_425J2_127_3477_n797) );
  FADDX1_HVT DP_OP_425J2_127_3477_U579 ( .A(DP_OP_425J2_127_3477_n2588), .B(
        DP_OP_425J2_127_3477_n2250), .CI(DP_OP_425J2_127_3477_n2602), .CO(
        DP_OP_425J2_127_3477_n794), .S(DP_OP_425J2_127_3477_n795) );
  FADDX1_HVT DP_OP_425J2_127_3477_U578 ( .A(DP_OP_425J2_127_3477_n2544), .B(
        DP_OP_425J2_127_3477_n2412), .CI(DP_OP_425J2_127_3477_n2734), .CO(
        DP_OP_425J2_127_3477_n792), .S(DP_OP_425J2_127_3477_n793) );
  FADDX1_HVT DP_OP_425J2_127_3477_U577 ( .A(DP_OP_425J2_127_3477_n2852), .B(
        DP_OP_425J2_127_3477_n2148), .CI(DP_OP_425J2_127_3477_n2324), .CO(
        DP_OP_425J2_127_3477_n790), .S(DP_OP_425J2_127_3477_n791) );
  FADDX1_HVT DP_OP_425J2_127_3477_U576 ( .A(DP_OP_425J2_127_3477_n2016), .B(
        DP_OP_425J2_127_3477_n2632), .CI(DP_OP_425J2_127_3477_n2984), .CO(
        DP_OP_425J2_127_3477_n788), .S(DP_OP_425J2_127_3477_n789) );
  FADDX1_HVT DP_OP_425J2_127_3477_U575 ( .A(DP_OP_425J2_127_3477_n2940), .B(
        DP_OP_425J2_127_3477_n2456), .CI(DP_OP_425J2_127_3477_n821), .CO(
        DP_OP_425J2_127_3477_n786), .S(DP_OP_425J2_127_3477_n787) );
  FADDX1_HVT DP_OP_425J2_127_3477_U574 ( .A(DP_OP_425J2_127_3477_n2287), .B(
        DP_OP_425J2_127_3477_n2023), .CI(DP_OP_425J2_127_3477_n1979), .CO(
        DP_OP_425J2_127_3477_n784), .S(DP_OP_425J2_127_3477_n785) );
  FADDX1_HVT DP_OP_425J2_127_3477_U573 ( .A(DP_OP_425J2_127_3477_n3033), .B(
        DP_OP_425J2_127_3477_n2067), .CI(DP_OP_425J2_127_3477_n2111), .CO(
        DP_OP_425J2_127_3477_n782), .S(DP_OP_425J2_127_3477_n783) );
  FADDX1_HVT DP_OP_425J2_127_3477_U572 ( .A(DP_OP_425J2_127_3477_n2991), .B(
        DP_OP_425J2_127_3477_n2155), .CI(DP_OP_425J2_127_3477_n2199), .CO(
        DP_OP_425J2_127_3477_n780), .S(DP_OP_425J2_127_3477_n781) );
  FADDX1_HVT DP_OP_425J2_127_3477_U571 ( .A(DP_OP_425J2_127_3477_n2947), .B(
        DP_OP_425J2_127_3477_n2243), .CI(DP_OP_425J2_127_3477_n2331), .CO(
        DP_OP_425J2_127_3477_n778), .S(DP_OP_425J2_127_3477_n779) );
  FADDX1_HVT DP_OP_425J2_127_3477_U570 ( .A(DP_OP_425J2_127_3477_n2903), .B(
        DP_OP_425J2_127_3477_n2375), .CI(DP_OP_425J2_127_3477_n2419), .CO(
        DP_OP_425J2_127_3477_n776), .S(DP_OP_425J2_127_3477_n777) );
  FADDX1_HVT DP_OP_425J2_127_3477_U569 ( .A(DP_OP_425J2_127_3477_n2859), .B(
        DP_OP_425J2_127_3477_n2463), .CI(DP_OP_425J2_127_3477_n2507), .CO(
        DP_OP_425J2_127_3477_n774), .S(DP_OP_425J2_127_3477_n775) );
  FADDX1_HVT DP_OP_425J2_127_3477_U568 ( .A(DP_OP_425J2_127_3477_n2815), .B(
        DP_OP_425J2_127_3477_n2551), .CI(DP_OP_425J2_127_3477_n2595), .CO(
        DP_OP_425J2_127_3477_n772), .S(DP_OP_425J2_127_3477_n773) );
  FADDX1_HVT DP_OP_425J2_127_3477_U567 ( .A(DP_OP_425J2_127_3477_n2771), .B(
        DP_OP_425J2_127_3477_n2639), .CI(DP_OP_425J2_127_3477_n2683), .CO(
        DP_OP_425J2_127_3477_n770), .S(DP_OP_425J2_127_3477_n771) );
  FADDX1_HVT DP_OP_425J2_127_3477_U566 ( .A(DP_OP_425J2_127_3477_n2727), .B(
        DP_OP_425J2_127_3477_n1016), .CI(DP_OP_425J2_127_3477_n1014), .CO(
        DP_OP_425J2_127_3477_n768), .S(DP_OP_425J2_127_3477_n769) );
  FADDX1_HVT DP_OP_425J2_127_3477_U565 ( .A(DP_OP_425J2_127_3477_n1012), .B(
        DP_OP_425J2_127_3477_n984), .CI(DP_OP_425J2_127_3477_n986), .CO(
        DP_OP_425J2_127_3477_n766), .S(DP_OP_425J2_127_3477_n767) );
  FADDX1_HVT DP_OP_425J2_127_3477_U564 ( .A(DP_OP_425J2_127_3477_n1010), .B(
        DP_OP_425J2_127_3477_n988), .CI(DP_OP_425J2_127_3477_n990), .CO(
        DP_OP_425J2_127_3477_n764), .S(DP_OP_425J2_127_3477_n765) );
  FADDX1_HVT DP_OP_425J2_127_3477_U563 ( .A(DP_OP_425J2_127_3477_n1008), .B(
        DP_OP_425J2_127_3477_n992), .CI(DP_OP_425J2_127_3477_n994), .CO(
        DP_OP_425J2_127_3477_n762), .S(DP_OP_425J2_127_3477_n763) );
  FADDX1_HVT DP_OP_425J2_127_3477_U562 ( .A(DP_OP_425J2_127_3477_n1000), .B(
        DP_OP_425J2_127_3477_n1006), .CI(DP_OP_425J2_127_3477_n996), .CO(
        DP_OP_425J2_127_3477_n760), .S(DP_OP_425J2_127_3477_n761) );
  FADDX1_HVT DP_OP_425J2_127_3477_U561 ( .A(DP_OP_425J2_127_3477_n998), .B(
        DP_OP_425J2_127_3477_n1002), .CI(DP_OP_425J2_127_3477_n1004), .CO(
        DP_OP_425J2_127_3477_n758), .S(DP_OP_425J2_127_3477_n759) );
  FADDX1_HVT DP_OP_425J2_127_3477_U560 ( .A(DP_OP_425J2_127_3477_n982), .B(
        DP_OP_425J2_127_3477_n980), .CI(DP_OP_425J2_127_3477_n950), .CO(
        DP_OP_425J2_127_3477_n756), .S(DP_OP_425J2_127_3477_n757) );
  FADDX1_HVT DP_OP_425J2_127_3477_U559 ( .A(DP_OP_425J2_127_3477_n964), .B(
        DP_OP_425J2_127_3477_n952), .CI(DP_OP_425J2_127_3477_n954), .CO(
        DP_OP_425J2_127_3477_n754), .S(DP_OP_425J2_127_3477_n755) );
  FADDX1_HVT DP_OP_425J2_127_3477_U558 ( .A(DP_OP_425J2_127_3477_n962), .B(
        DP_OP_425J2_127_3477_n956), .CI(DP_OP_425J2_127_3477_n958), .CO(
        DP_OP_425J2_127_3477_n752), .S(DP_OP_425J2_127_3477_n753) );
  FADDX1_HVT DP_OP_425J2_127_3477_U557 ( .A(DP_OP_425J2_127_3477_n960), .B(
        DP_OP_425J2_127_3477_n978), .CI(DP_OP_425J2_127_3477_n976), .CO(
        DP_OP_425J2_127_3477_n750), .S(DP_OP_425J2_127_3477_n751) );
  FADDX1_HVT DP_OP_425J2_127_3477_U556 ( .A(DP_OP_425J2_127_3477_n970), .B(
        DP_OP_425J2_127_3477_n966), .CI(DP_OP_425J2_127_3477_n968), .CO(
        DP_OP_425J2_127_3477_n748), .S(DP_OP_425J2_127_3477_n749) );
  FADDX1_HVT DP_OP_425J2_127_3477_U555 ( .A(DP_OP_425J2_127_3477_n974), .B(
        DP_OP_425J2_127_3477_n972), .CI(DP_OP_425J2_127_3477_n813), .CO(
        DP_OP_425J2_127_3477_n746), .S(DP_OP_425J2_127_3477_n747) );
  FADDX1_HVT DP_OP_425J2_127_3477_U554 ( .A(DP_OP_425J2_127_3477_n809), .B(
        DP_OP_425J2_127_3477_n805), .CI(DP_OP_425J2_127_3477_n787), .CO(
        DP_OP_425J2_127_3477_n744), .S(DP_OP_425J2_127_3477_n745) );
  FADDX1_HVT DP_OP_425J2_127_3477_U553 ( .A(DP_OP_425J2_127_3477_n811), .B(
        DP_OP_425J2_127_3477_n793), .CI(DP_OP_425J2_127_3477_n791), .CO(
        DP_OP_425J2_127_3477_n742), .S(DP_OP_425J2_127_3477_n743) );
  FADDX1_HVT DP_OP_425J2_127_3477_U552 ( .A(DP_OP_425J2_127_3477_n803), .B(
        DP_OP_425J2_127_3477_n807), .CI(DP_OP_425J2_127_3477_n799), .CO(
        DP_OP_425J2_127_3477_n740), .S(DP_OP_425J2_127_3477_n741) );
  FADDX1_HVT DP_OP_425J2_127_3477_U551 ( .A(DP_OP_425J2_127_3477_n815), .B(
        DP_OP_425J2_127_3477_n795), .CI(DP_OP_425J2_127_3477_n789), .CO(
        DP_OP_425J2_127_3477_n738), .S(DP_OP_425J2_127_3477_n739) );
  FADDX1_HVT DP_OP_425J2_127_3477_U550 ( .A(DP_OP_425J2_127_3477_n797), .B(
        DP_OP_425J2_127_3477_n819), .CI(DP_OP_425J2_127_3477_n817), .CO(
        DP_OP_425J2_127_3477_n736), .S(DP_OP_425J2_127_3477_n737) );
  FADDX1_HVT DP_OP_425J2_127_3477_U549 ( .A(DP_OP_425J2_127_3477_n801), .B(
        DP_OP_425J2_127_3477_n781), .CI(DP_OP_425J2_127_3477_n777), .CO(
        DP_OP_425J2_127_3477_n734), .S(DP_OP_425J2_127_3477_n735) );
  FADDX1_HVT DP_OP_425J2_127_3477_U548 ( .A(DP_OP_425J2_127_3477_n773), .B(
        DP_OP_425J2_127_3477_n771), .CI(DP_OP_425J2_127_3477_n783), .CO(
        DP_OP_425J2_127_3477_n732), .S(DP_OP_425J2_127_3477_n733) );
  FADDX1_HVT DP_OP_425J2_127_3477_U547 ( .A(DP_OP_425J2_127_3477_n779), .B(
        DP_OP_425J2_127_3477_n775), .CI(DP_OP_425J2_127_3477_n785), .CO(
        DP_OP_425J2_127_3477_n730), .S(DP_OP_425J2_127_3477_n731) );
  FADDX1_HVT DP_OP_425J2_127_3477_U546 ( .A(DP_OP_425J2_127_3477_n948), .B(
        DP_OP_425J2_127_3477_n944), .CI(DP_OP_425J2_127_3477_n946), .CO(
        DP_OP_425J2_127_3477_n728), .S(DP_OP_425J2_127_3477_n729) );
  FADDX1_HVT DP_OP_425J2_127_3477_U545 ( .A(DP_OP_425J2_127_3477_n942), .B(
        DP_OP_425J2_127_3477_n928), .CI(DP_OP_425J2_127_3477_n930), .CO(
        DP_OP_425J2_127_3477_n726), .S(DP_OP_425J2_127_3477_n727) );
  FADDX1_HVT DP_OP_425J2_127_3477_U544 ( .A(DP_OP_425J2_127_3477_n940), .B(
        DP_OP_425J2_127_3477_n932), .CI(DP_OP_425J2_127_3477_n938), .CO(
        DP_OP_425J2_127_3477_n724), .S(DP_OP_425J2_127_3477_n725) );
  FADDX1_HVT DP_OP_425J2_127_3477_U543 ( .A(DP_OP_425J2_127_3477_n936), .B(
        DP_OP_425J2_127_3477_n934), .CI(DP_OP_425J2_127_3477_n769), .CO(
        DP_OP_425J2_127_3477_n722), .S(DP_OP_425J2_127_3477_n723) );
  FADDX1_HVT DP_OP_425J2_127_3477_U542 ( .A(DP_OP_425J2_127_3477_n926), .B(
        DP_OP_425J2_127_3477_n767), .CI(DP_OP_425J2_127_3477_n765), .CO(
        DP_OP_425J2_127_3477_n720), .S(DP_OP_425J2_127_3477_n721) );
  FADDX1_HVT DP_OP_425J2_127_3477_U541 ( .A(DP_OP_425J2_127_3477_n924), .B(
        DP_OP_425J2_127_3477_n761), .CI(DP_OP_425J2_127_3477_n763), .CO(
        DP_OP_425J2_127_3477_n718), .S(DP_OP_425J2_127_3477_n719) );
  FADDX1_HVT DP_OP_425J2_127_3477_U540 ( .A(DP_OP_425J2_127_3477_n922), .B(
        DP_OP_425J2_127_3477_n759), .CI(DP_OP_425J2_127_3477_n916), .CO(
        DP_OP_425J2_127_3477_n716), .S(DP_OP_425J2_127_3477_n717) );
  FADDX1_HVT DP_OP_425J2_127_3477_U539 ( .A(DP_OP_425J2_127_3477_n920), .B(
        DP_OP_425J2_127_3477_n918), .CI(DP_OP_425J2_127_3477_n906), .CO(
        DP_OP_425J2_127_3477_n714), .S(DP_OP_425J2_127_3477_n715) );
  FADDX1_HVT DP_OP_425J2_127_3477_U538 ( .A(DP_OP_425J2_127_3477_n914), .B(
        DP_OP_425J2_127_3477_n757), .CI(DP_OP_425J2_127_3477_n747), .CO(
        DP_OP_425J2_127_3477_n712), .S(DP_OP_425J2_127_3477_n713) );
  FADDX1_HVT DP_OP_425J2_127_3477_U537 ( .A(DP_OP_425J2_127_3477_n912), .B(
        DP_OP_425J2_127_3477_n753), .CI(DP_OP_425J2_127_3477_n749), .CO(
        DP_OP_425J2_127_3477_n710), .S(DP_OP_425J2_127_3477_n711) );
  FADDX1_HVT DP_OP_425J2_127_3477_U536 ( .A(DP_OP_425J2_127_3477_n910), .B(
        DP_OP_425J2_127_3477_n755), .CI(DP_OP_425J2_127_3477_n751), .CO(
        DP_OP_425J2_127_3477_n708), .S(DP_OP_425J2_127_3477_n709) );
  FADDX1_HVT DP_OP_425J2_127_3477_U535 ( .A(DP_OP_425J2_127_3477_n908), .B(
        DP_OP_425J2_127_3477_n743), .CI(DP_OP_425J2_127_3477_n739), .CO(
        DP_OP_425J2_127_3477_n706), .S(DP_OP_425J2_127_3477_n707) );
  FADDX1_HVT DP_OP_425J2_127_3477_U534 ( .A(DP_OP_425J2_127_3477_n741), .B(
        DP_OP_425J2_127_3477_n904), .CI(DP_OP_425J2_127_3477_n735), .CO(
        DP_OP_425J2_127_3477_n704), .S(DP_OP_425J2_127_3477_n705) );
  FADDX1_HVT DP_OP_425J2_127_3477_U533 ( .A(DP_OP_425J2_127_3477_n737), .B(
        DP_OP_425J2_127_3477_n745), .CI(DP_OP_425J2_127_3477_n731), .CO(
        DP_OP_425J2_127_3477_n702), .S(DP_OP_425J2_127_3477_n703) );
  FADDX1_HVT DP_OP_425J2_127_3477_U532 ( .A(DP_OP_425J2_127_3477_n733), .B(
        DP_OP_425J2_127_3477_n902), .CI(DP_OP_425J2_127_3477_n900), .CO(
        DP_OP_425J2_127_3477_n700), .S(DP_OP_425J2_127_3477_n701) );
  FADDX1_HVT DP_OP_425J2_127_3477_U531 ( .A(DP_OP_425J2_127_3477_n898), .B(
        DP_OP_425J2_127_3477_n896), .CI(DP_OP_425J2_127_3477_n729), .CO(
        DP_OP_425J2_127_3477_n698), .S(DP_OP_425J2_127_3477_n699) );
  FADDX1_HVT DP_OP_425J2_127_3477_U530 ( .A(DP_OP_425J2_127_3477_n894), .B(
        DP_OP_425J2_127_3477_n892), .CI(DP_OP_425J2_127_3477_n890), .CO(
        DP_OP_425J2_127_3477_n696), .S(DP_OP_425J2_127_3477_n697) );
  FADDX1_HVT DP_OP_425J2_127_3477_U529 ( .A(DP_OP_425J2_127_3477_n888), .B(
        DP_OP_425J2_127_3477_n723), .CI(DP_OP_425J2_127_3477_n882), .CO(
        DP_OP_425J2_127_3477_n694), .S(DP_OP_425J2_127_3477_n695) );
  FADDX1_HVT DP_OP_425J2_127_3477_U528 ( .A(DP_OP_425J2_127_3477_n886), .B(
        DP_OP_425J2_127_3477_n725), .CI(DP_OP_425J2_127_3477_n727), .CO(
        DP_OP_425J2_127_3477_n692), .S(DP_OP_425J2_127_3477_n693) );
  FADDX1_HVT DP_OP_425J2_127_3477_U527 ( .A(DP_OP_425J2_127_3477_n884), .B(
        DP_OP_425J2_127_3477_n721), .CI(DP_OP_425J2_127_3477_n717), .CO(
        DP_OP_425J2_127_3477_n690), .S(DP_OP_425J2_127_3477_n691) );
  FADDX1_HVT DP_OP_425J2_127_3477_U526 ( .A(DP_OP_425J2_127_3477_n880), .B(
        DP_OP_425J2_127_3477_n719), .CI(DP_OP_425J2_127_3477_n715), .CO(
        DP_OP_425J2_127_3477_n688), .S(DP_OP_425J2_127_3477_n689) );
  FADDX1_HVT DP_OP_425J2_127_3477_U525 ( .A(DP_OP_425J2_127_3477_n878), .B(
        DP_OP_425J2_127_3477_n876), .CI(DP_OP_425J2_127_3477_n711), .CO(
        DP_OP_425J2_127_3477_n686), .S(DP_OP_425J2_127_3477_n687) );
  FADDX1_HVT DP_OP_425J2_127_3477_U524 ( .A(DP_OP_425J2_127_3477_n709), .B(
        DP_OP_425J2_127_3477_n713), .CI(DP_OP_425J2_127_3477_n874), .CO(
        DP_OP_425J2_127_3477_n684), .S(DP_OP_425J2_127_3477_n685) );
  FADDX1_HVT DP_OP_425J2_127_3477_U523 ( .A(DP_OP_425J2_127_3477_n707), .B(
        DP_OP_425J2_127_3477_n872), .CI(DP_OP_425J2_127_3477_n703), .CO(
        DP_OP_425J2_127_3477_n682), .S(DP_OP_425J2_127_3477_n683) );
  FADDX1_HVT DP_OP_425J2_127_3477_U522 ( .A(DP_OP_425J2_127_3477_n705), .B(
        DP_OP_425J2_127_3477_n701), .CI(DP_OP_425J2_127_3477_n870), .CO(
        DP_OP_425J2_127_3477_n680), .S(DP_OP_425J2_127_3477_n681) );
  FADDX1_HVT DP_OP_425J2_127_3477_U521 ( .A(DP_OP_425J2_127_3477_n868), .B(
        DP_OP_425J2_127_3477_n866), .CI(DP_OP_425J2_127_3477_n699), .CO(
        DP_OP_425J2_127_3477_n678), .S(DP_OP_425J2_127_3477_n679) );
  FADDX1_HVT DP_OP_425J2_127_3477_U520 ( .A(DP_OP_425J2_127_3477_n864), .B(
        DP_OP_425J2_127_3477_n862), .CI(DP_OP_425J2_127_3477_n697), .CO(
        DP_OP_425J2_127_3477_n676), .S(DP_OP_425J2_127_3477_n677) );
  FADDX1_HVT DP_OP_425J2_127_3477_U519 ( .A(DP_OP_425J2_127_3477_n860), .B(
        DP_OP_425J2_127_3477_n693), .CI(DP_OP_425J2_127_3477_n856), .CO(
        DP_OP_425J2_127_3477_n674), .S(DP_OP_425J2_127_3477_n675) );
  FADDX1_HVT DP_OP_425J2_127_3477_U518 ( .A(DP_OP_425J2_127_3477_n858), .B(
        DP_OP_425J2_127_3477_n695), .CI(DP_OP_425J2_127_3477_n691), .CO(
        DP_OP_425J2_127_3477_n672), .S(DP_OP_425J2_127_3477_n673) );
  FADDX1_HVT DP_OP_425J2_127_3477_U517 ( .A(DP_OP_425J2_127_3477_n689), .B(
        DP_OP_425J2_127_3477_n687), .CI(DP_OP_425J2_127_3477_n854), .CO(
        DP_OP_425J2_127_3477_n670), .S(DP_OP_425J2_127_3477_n671) );
  FADDX1_HVT DP_OP_425J2_127_3477_U516 ( .A(DP_OP_425J2_127_3477_n685), .B(
        DP_OP_425J2_127_3477_n852), .CI(DP_OP_425J2_127_3477_n683), .CO(
        DP_OP_425J2_127_3477_n668), .S(DP_OP_425J2_127_3477_n669) );
  FADDX1_HVT DP_OP_425J2_127_3477_U515 ( .A(DP_OP_425J2_127_3477_n850), .B(
        DP_OP_425J2_127_3477_n681), .CI(DP_OP_425J2_127_3477_n848), .CO(
        DP_OP_425J2_127_3477_n666), .S(DP_OP_425J2_127_3477_n667) );
  FADDX1_HVT DP_OP_425J2_127_3477_U514 ( .A(DP_OP_425J2_127_3477_n846), .B(
        DP_OP_425J2_127_3477_n679), .CI(DP_OP_425J2_127_3477_n844), .CO(
        DP_OP_425J2_127_3477_n664), .S(DP_OP_425J2_127_3477_n665) );
  FADDX1_HVT DP_OP_425J2_127_3477_U513 ( .A(DP_OP_425J2_127_3477_n677), .B(
        DP_OP_425J2_127_3477_n842), .CI(DP_OP_425J2_127_3477_n675), .CO(
        DP_OP_425J2_127_3477_n662), .S(DP_OP_425J2_127_3477_n663) );
  FADDX1_HVT DP_OP_425J2_127_3477_U512 ( .A(DP_OP_425J2_127_3477_n673), .B(
        DP_OP_425J2_127_3477_n840), .CI(DP_OP_425J2_127_3477_n671), .CO(
        DP_OP_425J2_127_3477_n660), .S(DP_OP_425J2_127_3477_n661) );
  FADDX1_HVT DP_OP_425J2_127_3477_U511 ( .A(DP_OP_425J2_127_3477_n838), .B(
        DP_OP_425J2_127_3477_n669), .CI(DP_OP_425J2_127_3477_n836), .CO(
        DP_OP_425J2_127_3477_n658), .S(DP_OP_425J2_127_3477_n659) );
  FADDX1_HVT DP_OP_425J2_127_3477_U510 ( .A(DP_OP_425J2_127_3477_n667), .B(
        DP_OP_425J2_127_3477_n834), .CI(DP_OP_425J2_127_3477_n665), .CO(
        DP_OP_425J2_127_3477_n656), .S(DP_OP_425J2_127_3477_n657) );
  FADDX1_HVT DP_OP_425J2_127_3477_U509 ( .A(DP_OP_425J2_127_3477_n663), .B(
        DP_OP_425J2_127_3477_n832), .CI(DP_OP_425J2_127_3477_n661), .CO(
        DP_OP_425J2_127_3477_n654), .S(DP_OP_425J2_127_3477_n655) );
  FADDX1_HVT DP_OP_425J2_127_3477_U508 ( .A(DP_OP_425J2_127_3477_n830), .B(
        DP_OP_425J2_127_3477_n659), .CI(DP_OP_425J2_127_3477_n828), .CO(
        DP_OP_425J2_127_3477_n652), .S(DP_OP_425J2_127_3477_n653) );
  FADDX1_HVT DP_OP_425J2_127_3477_U507 ( .A(DP_OP_425J2_127_3477_n657), .B(
        DP_OP_425J2_127_3477_n826), .CI(DP_OP_425J2_127_3477_n655), .CO(
        DP_OP_425J2_127_3477_n650), .S(DP_OP_425J2_127_3477_n651) );
  FADDX1_HVT DP_OP_425J2_127_3477_U505 ( .A(DP_OP_425J2_127_3477_n3027), .B(
        DP_OP_425J2_127_3477_n1971), .CI(DP_OP_425J2_127_3477_n1927), .CO(
        DP_OP_425J2_127_3477_n646), .S(DP_OP_425J2_127_3477_n647) );
  FADDX1_HVT DP_OP_425J2_127_3477_U504 ( .A(DP_OP_425J2_127_3477_n820), .B(
        DP_OP_425J2_127_3477_n2286), .CI(DP_OP_425J2_127_3477_n1978), .CO(
        DP_OP_425J2_127_3477_n644), .S(DP_OP_425J2_127_3477_n645) );
  FADDX1_HVT DP_OP_425J2_127_3477_U503 ( .A(DP_OP_425J2_127_3477_n2367), .B(
        DP_OP_425J2_127_3477_n3032), .CI(DP_OP_425J2_127_3477_n2682), .CO(
        DP_OP_425J2_127_3477_n642), .S(DP_OP_425J2_127_3477_n643) );
  FADDX1_HVT DP_OP_425J2_127_3477_U502 ( .A(DP_OP_425J2_127_3477_n2059), .B(
        DP_OP_425J2_127_3477_n2594), .CI(DP_OP_425J2_127_3477_n2814), .CO(
        DP_OP_425J2_127_3477_n640), .S(DP_OP_425J2_127_3477_n641) );
  FADDX1_HVT DP_OP_425J2_127_3477_U501 ( .A(DP_OP_425J2_127_3477_n2279), .B(
        DP_OP_425J2_127_3477_n2374), .CI(DP_OP_425J2_127_3477_n2990), .CO(
        DP_OP_425J2_127_3477_n638), .S(DP_OP_425J2_127_3477_n639) );
  FADDX1_HVT DP_OP_425J2_127_3477_U500 ( .A(DP_OP_425J2_127_3477_n2015), .B(
        DP_OP_425J2_127_3477_n2902), .CI(DP_OP_425J2_127_3477_n2066), .CO(
        DP_OP_425J2_127_3477_n636), .S(DP_OP_425J2_127_3477_n637) );
  FADDX1_HVT DP_OP_425J2_127_3477_U499 ( .A(DP_OP_425J2_127_3477_n2147), .B(
        DP_OP_425J2_127_3477_n2022), .CI(DP_OP_425J2_127_3477_n2858), .CO(
        DP_OP_425J2_127_3477_n634), .S(DP_OP_425J2_127_3477_n635) );
  FADDX1_HVT DP_OP_425J2_127_3477_U498 ( .A(DP_OP_425J2_127_3477_n2983), .B(
        DP_OP_425J2_127_3477_n2418), .CI(DP_OP_425J2_127_3477_n2506), .CO(
        DP_OP_425J2_127_3477_n632), .S(DP_OP_425J2_127_3477_n633) );
  FADDX1_HVT DP_OP_425J2_127_3477_U497 ( .A(DP_OP_425J2_127_3477_n2499), .B(
        DP_OP_425J2_127_3477_n2550), .CI(DP_OP_425J2_127_3477_n2946), .CO(
        DP_OP_425J2_127_3477_n630), .S(DP_OP_425J2_127_3477_n631) );
  FADDX1_HVT DP_OP_425J2_127_3477_U496 ( .A(DP_OP_425J2_127_3477_n2763), .B(
        DP_OP_425J2_127_3477_n2242), .CI(DP_OP_425J2_127_3477_n2770), .CO(
        DP_OP_425J2_127_3477_n628), .S(DP_OP_425J2_127_3477_n629) );
  FADDX1_HVT DP_OP_425J2_127_3477_U495 ( .A(DP_OP_425J2_127_3477_n2939), .B(
        DP_OP_425J2_127_3477_n2462), .CI(DP_OP_425J2_127_3477_n2638), .CO(
        DP_OP_425J2_127_3477_n626), .S(DP_OP_425J2_127_3477_n627) );
  FADDX1_HVT DP_OP_425J2_127_3477_U494 ( .A(DP_OP_425J2_127_3477_n2235), .B(
        DP_OP_425J2_127_3477_n2110), .CI(DP_OP_425J2_127_3477_n2726), .CO(
        DP_OP_425J2_127_3477_n624), .S(DP_OP_425J2_127_3477_n625) );
  FADDX1_HVT DP_OP_425J2_127_3477_U493 ( .A(DP_OP_425J2_127_3477_n2191), .B(
        DP_OP_425J2_127_3477_n2330), .CI(DP_OP_425J2_127_3477_n2198), .CO(
        DP_OP_425J2_127_3477_n622), .S(DP_OP_425J2_127_3477_n623) );
  FADDX1_HVT DP_OP_425J2_127_3477_U492 ( .A(DP_OP_425J2_127_3477_n2587), .B(
        DP_OP_425J2_127_3477_n2411), .CI(DP_OP_425J2_127_3477_n2154), .CO(
        DP_OP_425J2_127_3477_n620), .S(DP_OP_425J2_127_3477_n621) );
  FADDX1_HVT DP_OP_425J2_127_3477_U491 ( .A(DP_OP_425J2_127_3477_n2895), .B(
        DP_OP_425J2_127_3477_n2103), .CI(DP_OP_425J2_127_3477_n2323), .CO(
        DP_OP_425J2_127_3477_n618), .S(DP_OP_425J2_127_3477_n619) );
  FADDX1_HVT DP_OP_425J2_127_3477_U490 ( .A(DP_OP_425J2_127_3477_n2851), .B(
        DP_OP_425J2_127_3477_n2455), .CI(DP_OP_425J2_127_3477_n2543), .CO(
        DP_OP_425J2_127_3477_n616), .S(DP_OP_425J2_127_3477_n617) );
  FADDX1_HVT DP_OP_425J2_127_3477_U489 ( .A(DP_OP_425J2_127_3477_n2807), .B(
        DP_OP_425J2_127_3477_n2631), .CI(DP_OP_425J2_127_3477_n2675), .CO(
        DP_OP_425J2_127_3477_n614), .S(DP_OP_425J2_127_3477_n615) );
  FADDX1_HVT DP_OP_425J2_127_3477_U488 ( .A(DP_OP_425J2_127_3477_n2719), .B(
        DP_OP_425J2_127_3477_n818), .CI(DP_OP_425J2_127_3477_n816), .CO(
        DP_OP_425J2_127_3477_n612), .S(DP_OP_425J2_127_3477_n613) );
  FADDX1_HVT DP_OP_425J2_127_3477_U487 ( .A(DP_OP_425J2_127_3477_n814), .B(
        DP_OP_425J2_127_3477_n786), .CI(DP_OP_425J2_127_3477_n788), .CO(
        DP_OP_425J2_127_3477_n610), .S(DP_OP_425J2_127_3477_n611) );
  FADDX1_HVT DP_OP_425J2_127_3477_U486 ( .A(DP_OP_425J2_127_3477_n812), .B(
        DP_OP_425J2_127_3477_n790), .CI(DP_OP_425J2_127_3477_n792), .CO(
        DP_OP_425J2_127_3477_n608), .S(DP_OP_425J2_127_3477_n609) );
  FADDX1_HVT DP_OP_425J2_127_3477_U485 ( .A(DP_OP_425J2_127_3477_n810), .B(
        DP_OP_425J2_127_3477_n794), .CI(DP_OP_425J2_127_3477_n796), .CO(
        DP_OP_425J2_127_3477_n606), .S(DP_OP_425J2_127_3477_n607) );
  FADDX1_HVT DP_OP_425J2_127_3477_U484 ( .A(DP_OP_425J2_127_3477_n808), .B(
        DP_OP_425J2_127_3477_n798), .CI(DP_OP_425J2_127_3477_n800), .CO(
        DP_OP_425J2_127_3477_n604), .S(DP_OP_425J2_127_3477_n605) );
  FADDX1_HVT DP_OP_425J2_127_3477_U483 ( .A(DP_OP_425J2_127_3477_n806), .B(
        DP_OP_425J2_127_3477_n802), .CI(DP_OP_425J2_127_3477_n804), .CO(
        DP_OP_425J2_127_3477_n602), .S(DP_OP_425J2_127_3477_n603) );
  FADDX1_HVT DP_OP_425J2_127_3477_U482 ( .A(DP_OP_425J2_127_3477_n784), .B(
        DP_OP_425J2_127_3477_n770), .CI(DP_OP_425J2_127_3477_n782), .CO(
        DP_OP_425J2_127_3477_n600), .S(DP_OP_425J2_127_3477_n601) );
  FADDX1_HVT DP_OP_425J2_127_3477_U481 ( .A(DP_OP_425J2_127_3477_n776), .B(
        DP_OP_425J2_127_3477_n772), .CI(DP_OP_425J2_127_3477_n774), .CO(
        DP_OP_425J2_127_3477_n598), .S(DP_OP_425J2_127_3477_n599) );
  FADDX1_HVT DP_OP_425J2_127_3477_U480 ( .A(DP_OP_425J2_127_3477_n780), .B(
        DP_OP_425J2_127_3477_n778), .CI(DP_OP_425J2_127_3477_n645), .CO(
        DP_OP_425J2_127_3477_n596), .S(DP_OP_425J2_127_3477_n597) );
  FADDX1_HVT DP_OP_425J2_127_3477_U479 ( .A(DP_OP_425J2_127_3477_n647), .B(
        DP_OP_425J2_127_3477_n633), .CI(DP_OP_425J2_127_3477_n639), .CO(
        DP_OP_425J2_127_3477_n594), .S(DP_OP_425J2_127_3477_n595) );
  FADDX1_HVT DP_OP_425J2_127_3477_U478 ( .A(DP_OP_425J2_127_3477_n615), .B(
        DP_OP_425J2_127_3477_n637), .CI(DP_OP_425J2_127_3477_n635), .CO(
        DP_OP_425J2_127_3477_n592), .S(DP_OP_425J2_127_3477_n593) );
  FADDX1_HVT DP_OP_425J2_127_3477_U477 ( .A(DP_OP_425J2_127_3477_n641), .B(
        DP_OP_425J2_127_3477_n623), .CI(DP_OP_425J2_127_3477_n625), .CO(
        DP_OP_425J2_127_3477_n590), .S(DP_OP_425J2_127_3477_n591) );
  FADDX1_HVT DP_OP_425J2_127_3477_U476 ( .A(DP_OP_425J2_127_3477_n627), .B(
        DP_OP_425J2_127_3477_n617), .CI(DP_OP_425J2_127_3477_n619), .CO(
        DP_OP_425J2_127_3477_n588), .S(DP_OP_425J2_127_3477_n589) );
  FADDX1_HVT DP_OP_425J2_127_3477_U475 ( .A(DP_OP_425J2_127_3477_n621), .B(
        DP_OP_425J2_127_3477_n643), .CI(DP_OP_425J2_127_3477_n631), .CO(
        DP_OP_425J2_127_3477_n586), .S(DP_OP_425J2_127_3477_n587) );
  FADDX1_HVT DP_OP_425J2_127_3477_U474 ( .A(DP_OP_425J2_127_3477_n629), .B(
        DP_OP_425J2_127_3477_n768), .CI(DP_OP_425J2_127_3477_n766), .CO(
        DP_OP_425J2_127_3477_n584), .S(DP_OP_425J2_127_3477_n585) );
  FADDX1_HVT DP_OP_425J2_127_3477_U473 ( .A(DP_OP_425J2_127_3477_n764), .B(
        DP_OP_425J2_127_3477_n758), .CI(DP_OP_425J2_127_3477_n760), .CO(
        DP_OP_425J2_127_3477_n582), .S(DP_OP_425J2_127_3477_n583) );
  FADDX1_HVT DP_OP_425J2_127_3477_U472 ( .A(DP_OP_425J2_127_3477_n762), .B(
        DP_OP_425J2_127_3477_n756), .CI(DP_OP_425J2_127_3477_n754), .CO(
        DP_OP_425J2_127_3477_n580), .S(DP_OP_425J2_127_3477_n581) );
  FADDX1_HVT DP_OP_425J2_127_3477_U471 ( .A(DP_OP_425J2_127_3477_n752), .B(
        DP_OP_425J2_127_3477_n748), .CI(DP_OP_425J2_127_3477_n746), .CO(
        DP_OP_425J2_127_3477_n578), .S(DP_OP_425J2_127_3477_n579) );
  FADDX1_HVT DP_OP_425J2_127_3477_U470 ( .A(DP_OP_425J2_127_3477_n750), .B(
        DP_OP_425J2_127_3477_n613), .CI(DP_OP_425J2_127_3477_n607), .CO(
        DP_OP_425J2_127_3477_n576), .S(DP_OP_425J2_127_3477_n577) );
  FADDX1_HVT DP_OP_425J2_127_3477_U469 ( .A(DP_OP_425J2_127_3477_n609), .B(
        DP_OP_425J2_127_3477_n603), .CI(DP_OP_425J2_127_3477_n734), .CO(
        DP_OP_425J2_127_3477_n574), .S(DP_OP_425J2_127_3477_n575) );
  FADDX1_HVT DP_OP_425J2_127_3477_U468 ( .A(DP_OP_425J2_127_3477_n744), .B(
        DP_OP_425J2_127_3477_n611), .CI(DP_OP_425J2_127_3477_n605), .CO(
        DP_OP_425J2_127_3477_n572), .S(DP_OP_425J2_127_3477_n573) );
  FADDX1_HVT DP_OP_425J2_127_3477_U467 ( .A(DP_OP_425J2_127_3477_n738), .B(
        DP_OP_425J2_127_3477_n742), .CI(DP_OP_425J2_127_3477_n736), .CO(
        DP_OP_425J2_127_3477_n570), .S(DP_OP_425J2_127_3477_n571) );
  FADDX1_HVT DP_OP_425J2_127_3477_U466 ( .A(DP_OP_425J2_127_3477_n740), .B(
        DP_OP_425J2_127_3477_n732), .CI(DP_OP_425J2_127_3477_n730), .CO(
        DP_OP_425J2_127_3477_n568), .S(DP_OP_425J2_127_3477_n569) );
  FADDX1_HVT DP_OP_425J2_127_3477_U465 ( .A(DP_OP_425J2_127_3477_n599), .B(
        DP_OP_425J2_127_3477_n601), .CI(DP_OP_425J2_127_3477_n597), .CO(
        DP_OP_425J2_127_3477_n566), .S(DP_OP_425J2_127_3477_n567) );
  FADDX1_HVT DP_OP_425J2_127_3477_U464 ( .A(DP_OP_425J2_127_3477_n595), .B(
        DP_OP_425J2_127_3477_n589), .CI(DP_OP_425J2_127_3477_n593), .CO(
        DP_OP_425J2_127_3477_n564), .S(DP_OP_425J2_127_3477_n565) );
  FADDX1_HVT DP_OP_425J2_127_3477_U463 ( .A(DP_OP_425J2_127_3477_n587), .B(
        DP_OP_425J2_127_3477_n591), .CI(DP_OP_425J2_127_3477_n728), .CO(
        DP_OP_425J2_127_3477_n562), .S(DP_OP_425J2_127_3477_n563) );
  FADDX1_HVT DP_OP_425J2_127_3477_U462 ( .A(DP_OP_425J2_127_3477_n726), .B(
        DP_OP_425J2_127_3477_n585), .CI(DP_OP_425J2_127_3477_n722), .CO(
        DP_OP_425J2_127_3477_n560), .S(DP_OP_425J2_127_3477_n561) );
  FADDX1_HVT DP_OP_425J2_127_3477_U461 ( .A(DP_OP_425J2_127_3477_n724), .B(
        DP_OP_425J2_127_3477_n720), .CI(DP_OP_425J2_127_3477_n718), .CO(
        DP_OP_425J2_127_3477_n558), .S(DP_OP_425J2_127_3477_n559) );
  FADDX1_HVT DP_OP_425J2_127_3477_U460 ( .A(DP_OP_425J2_127_3477_n716), .B(
        DP_OP_425J2_127_3477_n583), .CI(DP_OP_425J2_127_3477_n581), .CO(
        DP_OP_425J2_127_3477_n556), .S(DP_OP_425J2_127_3477_n557) );
  FADDX1_HVT DP_OP_425J2_127_3477_U459 ( .A(DP_OP_425J2_127_3477_n714), .B(
        DP_OP_425J2_127_3477_n712), .CI(DP_OP_425J2_127_3477_n710), .CO(
        DP_OP_425J2_127_3477_n554), .S(DP_OP_425J2_127_3477_n555) );
  FADDX1_HVT DP_OP_425J2_127_3477_U458 ( .A(DP_OP_425J2_127_3477_n708), .B(
        DP_OP_425J2_127_3477_n579), .CI(DP_OP_425J2_127_3477_n706), .CO(
        DP_OP_425J2_127_3477_n552), .S(DP_OP_425J2_127_3477_n553) );
  FADDX1_HVT DP_OP_425J2_127_3477_U457 ( .A(DP_OP_425J2_127_3477_n577), .B(
        DP_OP_425J2_127_3477_n704), .CI(DP_OP_425J2_127_3477_n575), .CO(
        DP_OP_425J2_127_3477_n550), .S(DP_OP_425J2_127_3477_n551) );
  FADDX1_HVT DP_OP_425J2_127_3477_U456 ( .A(DP_OP_425J2_127_3477_n702), .B(
        DP_OP_425J2_127_3477_n571), .CI(DP_OP_425J2_127_3477_n569), .CO(
        DP_OP_425J2_127_3477_n548), .S(DP_OP_425J2_127_3477_n549) );
  FADDX1_HVT DP_OP_425J2_127_3477_U455 ( .A(DP_OP_425J2_127_3477_n573), .B(
        DP_OP_425J2_127_3477_n567), .CI(DP_OP_425J2_127_3477_n700), .CO(
        DP_OP_425J2_127_3477_n546), .S(DP_OP_425J2_127_3477_n547) );
  FADDX1_HVT DP_OP_425J2_127_3477_U454 ( .A(DP_OP_425J2_127_3477_n565), .B(
        DP_OP_425J2_127_3477_n698), .CI(DP_OP_425J2_127_3477_n563), .CO(
        DP_OP_425J2_127_3477_n544), .S(DP_OP_425J2_127_3477_n545) );
  FADDX1_HVT DP_OP_425J2_127_3477_U453 ( .A(DP_OP_425J2_127_3477_n696), .B(
        DP_OP_425J2_127_3477_n694), .CI(DP_OP_425J2_127_3477_n692), .CO(
        DP_OP_425J2_127_3477_n542), .S(DP_OP_425J2_127_3477_n543) );
  FADDX1_HVT DP_OP_425J2_127_3477_U452 ( .A(DP_OP_425J2_127_3477_n561), .B(
        DP_OP_425J2_127_3477_n690), .CI(DP_OP_425J2_127_3477_n559), .CO(
        DP_OP_425J2_127_3477_n540), .S(DP_OP_425J2_127_3477_n541) );
  FADDX1_HVT DP_OP_425J2_127_3477_U451 ( .A(DP_OP_425J2_127_3477_n688), .B(
        DP_OP_425J2_127_3477_n557), .CI(DP_OP_425J2_127_3477_n555), .CO(
        DP_OP_425J2_127_3477_n538), .S(DP_OP_425J2_127_3477_n539) );
  FADDX1_HVT DP_OP_425J2_127_3477_U450 ( .A(DP_OP_425J2_127_3477_n686), .B(
        DP_OP_425J2_127_3477_n684), .CI(DP_OP_425J2_127_3477_n553), .CO(
        DP_OP_425J2_127_3477_n536), .S(DP_OP_425J2_127_3477_n537) );
  FADDX1_HVT DP_OP_425J2_127_3477_U449 ( .A(DP_OP_425J2_127_3477_n682), .B(
        DP_OP_425J2_127_3477_n551), .CI(DP_OP_425J2_127_3477_n549), .CO(
        DP_OP_425J2_127_3477_n534), .S(DP_OP_425J2_127_3477_n535) );
  FADDX1_HVT DP_OP_425J2_127_3477_U448 ( .A(DP_OP_425J2_127_3477_n680), .B(
        DP_OP_425J2_127_3477_n547), .CI(DP_OP_425J2_127_3477_n678), .CO(
        DP_OP_425J2_127_3477_n532), .S(DP_OP_425J2_127_3477_n533) );
  FADDX1_HVT DP_OP_425J2_127_3477_U447 ( .A(DP_OP_425J2_127_3477_n545), .B(
        DP_OP_425J2_127_3477_n676), .CI(DP_OP_425J2_127_3477_n543), .CO(
        DP_OP_425J2_127_3477_n530), .S(DP_OP_425J2_127_3477_n531) );
  FADDX1_HVT DP_OP_425J2_127_3477_U446 ( .A(DP_OP_425J2_127_3477_n674), .B(
        DP_OP_425J2_127_3477_n672), .CI(DP_OP_425J2_127_3477_n541), .CO(
        DP_OP_425J2_127_3477_n528), .S(DP_OP_425J2_127_3477_n529) );
  FADDX1_HVT DP_OP_425J2_127_3477_U445 ( .A(DP_OP_425J2_127_3477_n670), .B(
        DP_OP_425J2_127_3477_n539), .CI(DP_OP_425J2_127_3477_n537), .CO(
        DP_OP_425J2_127_3477_n526), .S(DP_OP_425J2_127_3477_n527) );
  FADDX1_HVT DP_OP_425J2_127_3477_U444 ( .A(DP_OP_425J2_127_3477_n535), .B(
        DP_OP_425J2_127_3477_n668), .CI(DP_OP_425J2_127_3477_n666), .CO(
        DP_OP_425J2_127_3477_n524), .S(DP_OP_425J2_127_3477_n525) );
  FADDX1_HVT DP_OP_425J2_127_3477_U443 ( .A(DP_OP_425J2_127_3477_n533), .B(
        DP_OP_425J2_127_3477_n664), .CI(DP_OP_425J2_127_3477_n531), .CO(
        DP_OP_425J2_127_3477_n522), .S(DP_OP_425J2_127_3477_n523) );
  FADDX1_HVT DP_OP_425J2_127_3477_U442 ( .A(DP_OP_425J2_127_3477_n662), .B(
        DP_OP_425J2_127_3477_n529), .CI(DP_OP_425J2_127_3477_n660), .CO(
        DP_OP_425J2_127_3477_n520), .S(DP_OP_425J2_127_3477_n521) );
  FADDX1_HVT DP_OP_425J2_127_3477_U441 ( .A(DP_OP_425J2_127_3477_n527), .B(
        DP_OP_425J2_127_3477_n658), .CI(DP_OP_425J2_127_3477_n525), .CO(
        DP_OP_425J2_127_3477_n518), .S(DP_OP_425J2_127_3477_n519) );
  FADDX1_HVT DP_OP_425J2_127_3477_U439 ( .A(DP_OP_425J2_127_3477_n521), .B(
        DP_OP_425J2_127_3477_n519), .CI(DP_OP_425J2_127_3477_n652), .CO(
        DP_OP_425J2_127_3477_n514), .S(DP_OP_425J2_127_3477_n515) );
  FADDX1_HVT DP_OP_425J2_127_3477_U436 ( .A(DP_OP_425J2_127_3477_n3026), .B(
        DP_OP_425J2_127_3477_n1970), .CI(DP_OP_425J2_127_3477_n511), .CO(
        DP_OP_425J2_127_3477_n508), .S(DP_OP_425J2_127_3477_n509) );
  FADDX1_HVT DP_OP_425J2_127_3477_U435 ( .A(DP_OP_425J2_127_3477_n2058), .B(
        DP_OP_425J2_127_3477_n2982), .CI(DP_OP_425J2_127_3477_n2410), .CO(
        DP_OP_425J2_127_3477_n506), .S(DP_OP_425J2_127_3477_n507) );
  FADDX1_HVT DP_OP_425J2_127_3477_U434 ( .A(DP_OP_425J2_127_3477_n2542), .B(
        DP_OP_425J2_127_3477_n2938), .CI(DP_OP_425J2_127_3477_n2894), .CO(
        DP_OP_425J2_127_3477_n504), .S(DP_OP_425J2_127_3477_n505) );
  FADDX1_HVT DP_OP_425J2_127_3477_U433 ( .A(DP_OP_425J2_127_3477_n2366), .B(
        DP_OP_425J2_127_3477_n2850), .CI(DP_OP_425J2_127_3477_n2806), .CO(
        DP_OP_425J2_127_3477_n502), .S(DP_OP_425J2_127_3477_n503) );
  FADDX1_HVT DP_OP_425J2_127_3477_U432 ( .A(DP_OP_425J2_127_3477_n2234), .B(
        DP_OP_425J2_127_3477_n2014), .CI(DP_OP_425J2_127_3477_n2762), .CO(
        DP_OP_425J2_127_3477_n500), .S(DP_OP_425J2_127_3477_n501) );
  FADDX1_HVT DP_OP_425J2_127_3477_U431 ( .A(DP_OP_425J2_127_3477_n2718), .B(
        DP_OP_425J2_127_3477_n2674), .CI(DP_OP_425J2_127_3477_n2630), .CO(
        DP_OP_425J2_127_3477_n498), .S(DP_OP_425J2_127_3477_n499) );
  FADDX1_HVT DP_OP_425J2_127_3477_U430 ( .A(DP_OP_425J2_127_3477_n2278), .B(
        DP_OP_425J2_127_3477_n2102), .CI(DP_OP_425J2_127_3477_n2146), .CO(
        DP_OP_425J2_127_3477_n496), .S(DP_OP_425J2_127_3477_n497) );
  FADDX1_HVT DP_OP_425J2_127_3477_U429 ( .A(DP_OP_425J2_127_3477_n2190), .B(
        DP_OP_425J2_127_3477_n2586), .CI(DP_OP_425J2_127_3477_n2498), .CO(
        DP_OP_425J2_127_3477_n494), .S(DP_OP_425J2_127_3477_n495) );
  FADDX1_HVT DP_OP_425J2_127_3477_U428 ( .A(DP_OP_425J2_127_3477_n2322), .B(
        DP_OP_425J2_127_3477_n2454), .CI(DP_OP_425J2_127_3477_n646), .CO(
        DP_OP_425J2_127_3477_n492), .S(DP_OP_425J2_127_3477_n493) );
  FADDX1_HVT DP_OP_425J2_127_3477_U427 ( .A(DP_OP_425J2_127_3477_n644), .B(
        DP_OP_425J2_127_3477_n614), .CI(DP_OP_425J2_127_3477_n642), .CO(
        DP_OP_425J2_127_3477_n490), .S(DP_OP_425J2_127_3477_n491) );
  FADDX1_HVT DP_OP_425J2_127_3477_U426 ( .A(DP_OP_425J2_127_3477_n640), .B(
        DP_OP_425J2_127_3477_n616), .CI(DP_OP_425J2_127_3477_n618), .CO(
        DP_OP_425J2_127_3477_n488), .S(DP_OP_425J2_127_3477_n489) );
  FADDX1_HVT DP_OP_425J2_127_3477_U425 ( .A(DP_OP_425J2_127_3477_n638), .B(
        DP_OP_425J2_127_3477_n620), .CI(DP_OP_425J2_127_3477_n622), .CO(
        DP_OP_425J2_127_3477_n486), .S(DP_OP_425J2_127_3477_n487) );
  FADDX1_HVT DP_OP_425J2_127_3477_U424 ( .A(DP_OP_425J2_127_3477_n636), .B(
        DP_OP_425J2_127_3477_n624), .CI(DP_OP_425J2_127_3477_n626), .CO(
        DP_OP_425J2_127_3477_n484), .S(DP_OP_425J2_127_3477_n485) );
  FADDX1_HVT DP_OP_425J2_127_3477_U423 ( .A(DP_OP_425J2_127_3477_n634), .B(
        DP_OP_425J2_127_3477_n628), .CI(DP_OP_425J2_127_3477_n630), .CO(
        DP_OP_425J2_127_3477_n482), .S(DP_OP_425J2_127_3477_n483) );
  FADDX1_HVT DP_OP_425J2_127_3477_U422 ( .A(DP_OP_425J2_127_3477_n632), .B(
        DP_OP_425J2_127_3477_n509), .CI(DP_OP_425J2_127_3477_n505), .CO(
        DP_OP_425J2_127_3477_n480), .S(DP_OP_425J2_127_3477_n481) );
  FADDX1_HVT DP_OP_425J2_127_3477_U421 ( .A(DP_OP_425J2_127_3477_n501), .B(
        DP_OP_425J2_127_3477_n495), .CI(DP_OP_425J2_127_3477_n497), .CO(
        DP_OP_425J2_127_3477_n478), .S(DP_OP_425J2_127_3477_n479) );
  FADDX1_HVT DP_OP_425J2_127_3477_U420 ( .A(DP_OP_425J2_127_3477_n499), .B(
        DP_OP_425J2_127_3477_n507), .CI(DP_OP_425J2_127_3477_n503), .CO(
        DP_OP_425J2_127_3477_n476), .S(DP_OP_425J2_127_3477_n477) );
  FADDX1_HVT DP_OP_425J2_127_3477_U419 ( .A(DP_OP_425J2_127_3477_n612), .B(
        DP_OP_425J2_127_3477_n610), .CI(DP_OP_425J2_127_3477_n602), .CO(
        DP_OP_425J2_127_3477_n474), .S(DP_OP_425J2_127_3477_n475) );
  FADDX1_HVT DP_OP_425J2_127_3477_U418 ( .A(DP_OP_425J2_127_3477_n608), .B(
        DP_OP_425J2_127_3477_n604), .CI(DP_OP_425J2_127_3477_n606), .CO(
        DP_OP_425J2_127_3477_n472), .S(DP_OP_425J2_127_3477_n473) );
  FADDX1_HVT DP_OP_425J2_127_3477_U417 ( .A(DP_OP_425J2_127_3477_n600), .B(
        DP_OP_425J2_127_3477_n596), .CI(DP_OP_425J2_127_3477_n493), .CO(
        DP_OP_425J2_127_3477_n470), .S(DP_OP_425J2_127_3477_n471) );
  FADDX1_HVT DP_OP_425J2_127_3477_U416 ( .A(DP_OP_425J2_127_3477_n598), .B(
        DP_OP_425J2_127_3477_n594), .CI(DP_OP_425J2_127_3477_n491), .CO(
        DP_OP_425J2_127_3477_n468), .S(DP_OP_425J2_127_3477_n469) );
  FADDX1_HVT DP_OP_425J2_127_3477_U415 ( .A(DP_OP_425J2_127_3477_n592), .B(
        DP_OP_425J2_127_3477_n485), .CI(DP_OP_425J2_127_3477_n487), .CO(
        DP_OP_425J2_127_3477_n466), .S(DP_OP_425J2_127_3477_n467) );
  FADDX1_HVT DP_OP_425J2_127_3477_U414 ( .A(DP_OP_425J2_127_3477_n590), .B(
        DP_OP_425J2_127_3477_n489), .CI(DP_OP_425J2_127_3477_n483), .CO(
        DP_OP_425J2_127_3477_n464), .S(DP_OP_425J2_127_3477_n465) );
  FADDX1_HVT DP_OP_425J2_127_3477_U413 ( .A(DP_OP_425J2_127_3477_n588), .B(
        DP_OP_425J2_127_3477_n586), .CI(DP_OP_425J2_127_3477_n584), .CO(
        DP_OP_425J2_127_3477_n462), .S(DP_OP_425J2_127_3477_n463) );
  FADDX1_HVT DP_OP_425J2_127_3477_U412 ( .A(DP_OP_425J2_127_3477_n481), .B(
        DP_OP_425J2_127_3477_n477), .CI(DP_OP_425J2_127_3477_n582), .CO(
        DP_OP_425J2_127_3477_n460), .S(DP_OP_425J2_127_3477_n461) );
  FADDX1_HVT DP_OP_425J2_127_3477_U411 ( .A(DP_OP_425J2_127_3477_n479), .B(
        DP_OP_425J2_127_3477_n580), .CI(DP_OP_425J2_127_3477_n578), .CO(
        DP_OP_425J2_127_3477_n458), .S(DP_OP_425J2_127_3477_n459) );
  FADDX1_HVT DP_OP_425J2_127_3477_U410 ( .A(DP_OP_425J2_127_3477_n576), .B(
        DP_OP_425J2_127_3477_n475), .CI(DP_OP_425J2_127_3477_n473), .CO(
        DP_OP_425J2_127_3477_n456), .S(DP_OP_425J2_127_3477_n457) );
  FADDX1_HVT DP_OP_425J2_127_3477_U409 ( .A(DP_OP_425J2_127_3477_n574), .B(
        DP_OP_425J2_127_3477_n570), .CI(DP_OP_425J2_127_3477_n568), .CO(
        DP_OP_425J2_127_3477_n454), .S(DP_OP_425J2_127_3477_n455) );
  FADDX1_HVT DP_OP_425J2_127_3477_U408 ( .A(DP_OP_425J2_127_3477_n572), .B(
        DP_OP_425J2_127_3477_n566), .CI(DP_OP_425J2_127_3477_n471), .CO(
        DP_OP_425J2_127_3477_n452), .S(DP_OP_425J2_127_3477_n453) );
  FADDX1_HVT DP_OP_425J2_127_3477_U407 ( .A(DP_OP_425J2_127_3477_n469), .B(
        DP_OP_425J2_127_3477_n564), .CI(DP_OP_425J2_127_3477_n562), .CO(
        DP_OP_425J2_127_3477_n450), .S(DP_OP_425J2_127_3477_n451) );
  FADDX1_HVT DP_OP_425J2_127_3477_U406 ( .A(DP_OP_425J2_127_3477_n467), .B(
        DP_OP_425J2_127_3477_n465), .CI(DP_OP_425J2_127_3477_n463), .CO(
        DP_OP_425J2_127_3477_n448), .S(DP_OP_425J2_127_3477_n449) );
  FADDX1_HVT DP_OP_425J2_127_3477_U405 ( .A(DP_OP_425J2_127_3477_n560), .B(
        DP_OP_425J2_127_3477_n558), .CI(DP_OP_425J2_127_3477_n461), .CO(
        DP_OP_425J2_127_3477_n446), .S(DP_OP_425J2_127_3477_n447) );
  FADDX1_HVT DP_OP_425J2_127_3477_U404 ( .A(DP_OP_425J2_127_3477_n556), .B(
        DP_OP_425J2_127_3477_n459), .CI(DP_OP_425J2_127_3477_n554), .CO(
        DP_OP_425J2_127_3477_n444), .S(DP_OP_425J2_127_3477_n445) );
  FADDX1_HVT DP_OP_425J2_127_3477_U403 ( .A(DP_OP_425J2_127_3477_n552), .B(
        DP_OP_425J2_127_3477_n457), .CI(DP_OP_425J2_127_3477_n550), .CO(
        DP_OP_425J2_127_3477_n442), .S(DP_OP_425J2_127_3477_n443) );
  FADDX1_HVT DP_OP_425J2_127_3477_U402 ( .A(DP_OP_425J2_127_3477_n548), .B(
        DP_OP_425J2_127_3477_n455), .CI(DP_OP_425J2_127_3477_n453), .CO(
        DP_OP_425J2_127_3477_n440), .S(DP_OP_425J2_127_3477_n441) );
  FADDX1_HVT DP_OP_425J2_127_3477_U401 ( .A(DP_OP_425J2_127_3477_n546), .B(
        DP_OP_425J2_127_3477_n451), .CI(DP_OP_425J2_127_3477_n544), .CO(
        DP_OP_425J2_127_3477_n438), .S(DP_OP_425J2_127_3477_n439) );
  FADDX1_HVT DP_OP_425J2_127_3477_U400 ( .A(DP_OP_425J2_127_3477_n449), .B(
        DP_OP_425J2_127_3477_n542), .CI(DP_OP_425J2_127_3477_n540), .CO(
        DP_OP_425J2_127_3477_n436), .S(DP_OP_425J2_127_3477_n437) );
  FADDX1_HVT DP_OP_425J2_127_3477_U399 ( .A(DP_OP_425J2_127_3477_n447), .B(
        DP_OP_425J2_127_3477_n538), .CI(DP_OP_425J2_127_3477_n445), .CO(
        DP_OP_425J2_127_3477_n434), .S(DP_OP_425J2_127_3477_n435) );
  FADDX1_HVT DP_OP_425J2_127_3477_U398 ( .A(DP_OP_425J2_127_3477_n536), .B(
        DP_OP_425J2_127_3477_n443), .CI(DP_OP_425J2_127_3477_n534), .CO(
        DP_OP_425J2_127_3477_n432), .S(DP_OP_425J2_127_3477_n433) );
  FADDX1_HVT DP_OP_425J2_127_3477_U397 ( .A(DP_OP_425J2_127_3477_n441), .B(
        DP_OP_425J2_127_3477_n532), .CI(DP_OP_425J2_127_3477_n439), .CO(
        DP_OP_425J2_127_3477_n430), .S(DP_OP_425J2_127_3477_n431) );
  FADDX1_HVT DP_OP_425J2_127_3477_U396 ( .A(DP_OP_425J2_127_3477_n530), .B(
        DP_OP_425J2_127_3477_n437), .CI(DP_OP_425J2_127_3477_n528), .CO(
        DP_OP_425J2_127_3477_n428), .S(DP_OP_425J2_127_3477_n429) );
  FADDX1_HVT DP_OP_425J2_127_3477_U395 ( .A(DP_OP_425J2_127_3477_n435), .B(
        DP_OP_425J2_127_3477_n526), .CI(DP_OP_425J2_127_3477_n433), .CO(
        DP_OP_425J2_127_3477_n426), .S(DP_OP_425J2_127_3477_n427) );
  FADDX1_HVT DP_OP_425J2_127_3477_U394 ( .A(DP_OP_425J2_127_3477_n524), .B(
        DP_OP_425J2_127_3477_n431), .CI(DP_OP_425J2_127_3477_n522), .CO(
        DP_OP_425J2_127_3477_n424), .S(DP_OP_425J2_127_3477_n425) );
  FADDX1_HVT DP_OP_425J2_127_3477_U393 ( .A(DP_OP_425J2_127_3477_n429), .B(
        DP_OP_425J2_127_3477_n520), .CI(DP_OP_425J2_127_3477_n427), .CO(
        DP_OP_425J2_127_3477_n422), .S(DP_OP_425J2_127_3477_n423) );
  FADDX1_HVT DP_OP_425J2_127_3477_U392 ( .A(DP_OP_425J2_127_3477_n518), .B(
        DP_OP_425J2_127_3477_n425), .CI(DP_OP_425J2_127_3477_n516), .CO(
        DP_OP_425J2_127_3477_n420), .S(DP_OP_425J2_127_3477_n421) );
  FADDX1_HVT DP_OP_425J2_127_3477_U390 ( .A(DP_OP_425J2_127_3477_n1926), .B(
        DP_OP_425J2_127_3477_n510), .CI(DP_OP_425J2_127_3477_n508), .CO(
        DP_OP_425J2_127_3477_n416), .S(DP_OP_425J2_127_3477_n417) );
  FADDX1_HVT DP_OP_425J2_127_3477_U389 ( .A(DP_OP_425J2_127_3477_n498), .B(
        DP_OP_425J2_127_3477_n494), .CI(DP_OP_425J2_127_3477_n506), .CO(
        DP_OP_425J2_127_3477_n414), .S(DP_OP_425J2_127_3477_n415) );
  FADDX1_HVT DP_OP_425J2_127_3477_U388 ( .A(DP_OP_425J2_127_3477_n504), .B(
        DP_OP_425J2_127_3477_n502), .CI(DP_OP_425J2_127_3477_n500), .CO(
        DP_OP_425J2_127_3477_n412), .S(DP_OP_425J2_127_3477_n413) );
  FADDX1_HVT DP_OP_425J2_127_3477_U387 ( .A(DP_OP_425J2_127_3477_n496), .B(
        DP_OP_425J2_127_3477_n492), .CI(DP_OP_425J2_127_3477_n490), .CO(
        DP_OP_425J2_127_3477_n410), .S(DP_OP_425J2_127_3477_n411) );
  FADDX1_HVT DP_OP_425J2_127_3477_U386 ( .A(DP_OP_425J2_127_3477_n488), .B(
        DP_OP_425J2_127_3477_n486), .CI(DP_OP_425J2_127_3477_n484), .CO(
        DP_OP_425J2_127_3477_n408), .S(DP_OP_425J2_127_3477_n409) );
  FADDX1_HVT DP_OP_425J2_127_3477_U385 ( .A(DP_OP_425J2_127_3477_n482), .B(
        DP_OP_425J2_127_3477_n417), .CI(DP_OP_425J2_127_3477_n480), .CO(
        DP_OP_425J2_127_3477_n406), .S(DP_OP_425J2_127_3477_n407) );
  FADDX1_HVT DP_OP_425J2_127_3477_U384 ( .A(DP_OP_425J2_127_3477_n478), .B(
        DP_OP_425J2_127_3477_n413), .CI(DP_OP_425J2_127_3477_n415), .CO(
        DP_OP_425J2_127_3477_n404), .S(DP_OP_425J2_127_3477_n405) );
  FADDX1_HVT DP_OP_425J2_127_3477_U383 ( .A(DP_OP_425J2_127_3477_n476), .B(
        DP_OP_425J2_127_3477_n474), .CI(DP_OP_425J2_127_3477_n472), .CO(
        DP_OP_425J2_127_3477_n402), .S(DP_OP_425J2_127_3477_n403) );
  FADDX1_HVT DP_OP_425J2_127_3477_U382 ( .A(DP_OP_425J2_127_3477_n470), .B(
        DP_OP_425J2_127_3477_n411), .CI(DP_OP_425J2_127_3477_n468), .CO(
        DP_OP_425J2_127_3477_n400), .S(DP_OP_425J2_127_3477_n401) );
  FADDX1_HVT DP_OP_425J2_127_3477_U381 ( .A(DP_OP_425J2_127_3477_n466), .B(
        DP_OP_425J2_127_3477_n409), .CI(DP_OP_425J2_127_3477_n464), .CO(
        DP_OP_425J2_127_3477_n398), .S(DP_OP_425J2_127_3477_n399) );
  FADDX1_HVT DP_OP_425J2_127_3477_U380 ( .A(DP_OP_425J2_127_3477_n462), .B(
        DP_OP_425J2_127_3477_n407), .CI(DP_OP_425J2_127_3477_n460), .CO(
        DP_OP_425J2_127_3477_n396), .S(DP_OP_425J2_127_3477_n397) );
  FADDX1_HVT DP_OP_425J2_127_3477_U379 ( .A(DP_OP_425J2_127_3477_n405), .B(
        DP_OP_425J2_127_3477_n458), .CI(DP_OP_425J2_127_3477_n456), .CO(
        DP_OP_425J2_127_3477_n394), .S(DP_OP_425J2_127_3477_n395) );
  FADDX1_HVT DP_OP_425J2_127_3477_U378 ( .A(DP_OP_425J2_127_3477_n403), .B(
        DP_OP_425J2_127_3477_n454), .CI(DP_OP_425J2_127_3477_n452), .CO(
        DP_OP_425J2_127_3477_n392), .S(DP_OP_425J2_127_3477_n393) );
  FADDX1_HVT DP_OP_425J2_127_3477_U377 ( .A(DP_OP_425J2_127_3477_n401), .B(
        DP_OP_425J2_127_3477_n450), .CI(DP_OP_425J2_127_3477_n399), .CO(
        DP_OP_425J2_127_3477_n390), .S(DP_OP_425J2_127_3477_n391) );
  FADDX1_HVT DP_OP_425J2_127_3477_U376 ( .A(DP_OP_425J2_127_3477_n448), .B(
        DP_OP_425J2_127_3477_n397), .CI(DP_OP_425J2_127_3477_n446), .CO(
        DP_OP_425J2_127_3477_n388), .S(DP_OP_425J2_127_3477_n389) );
  FADDX1_HVT DP_OP_425J2_127_3477_U375 ( .A(DP_OP_425J2_127_3477_n444), .B(
        DP_OP_425J2_127_3477_n395), .CI(DP_OP_425J2_127_3477_n442), .CO(
        DP_OP_425J2_127_3477_n386), .S(DP_OP_425J2_127_3477_n387) );
  FADDX1_HVT DP_OP_425J2_127_3477_U374 ( .A(DP_OP_425J2_127_3477_n393), .B(
        DP_OP_425J2_127_3477_n440), .CI(DP_OP_425J2_127_3477_n438), .CO(
        DP_OP_425J2_127_3477_n384), .S(DP_OP_425J2_127_3477_n385) );
  FADDX1_HVT DP_OP_425J2_127_3477_U373 ( .A(DP_OP_425J2_127_3477_n391), .B(
        DP_OP_425J2_127_3477_n436), .CI(DP_OP_425J2_127_3477_n389), .CO(
        DP_OP_425J2_127_3477_n382), .S(DP_OP_425J2_127_3477_n383) );
  FADDX1_HVT DP_OP_425J2_127_3477_U372 ( .A(DP_OP_425J2_127_3477_n434), .B(
        DP_OP_425J2_127_3477_n387), .CI(DP_OP_425J2_127_3477_n432), .CO(
        DP_OP_425J2_127_3477_n380), .S(DP_OP_425J2_127_3477_n381) );
  FADDX1_HVT DP_OP_425J2_127_3477_U368 ( .A(DP_OP_425J2_127_3477_n377), .B(
        DP_OP_425J2_127_3477_n420), .CI(DP_OP_425J2_127_3477_n375), .CO(
        DP_OP_425J2_127_3477_n372), .S(DP_OP_425J2_127_3477_n373) );
  FADDX1_HVT DP_OP_425J2_127_3477_U367 ( .A(DP_OP_425J2_127_3477_n1925), .B(
        DP_OP_425J2_127_3477_n416), .CI(DP_OP_425J2_127_3477_n414), .CO(
        DP_OP_425J2_127_3477_n370), .S(DP_OP_425J2_127_3477_n371) );
  FADDX1_HVT DP_OP_425J2_127_3477_U366 ( .A(DP_OP_425J2_127_3477_n412), .B(
        DP_OP_425J2_127_3477_n410), .CI(DP_OP_425J2_127_3477_n408), .CO(
        DP_OP_425J2_127_3477_n368), .S(DP_OP_425J2_127_3477_n369) );
  FADDX1_HVT DP_OP_425J2_127_3477_U365 ( .A(DP_OP_425J2_127_3477_n406), .B(
        DP_OP_425J2_127_3477_n371), .CI(DP_OP_425J2_127_3477_n404), .CO(
        DP_OP_425J2_127_3477_n366), .S(DP_OP_425J2_127_3477_n367) );
  FADDX1_HVT DP_OP_425J2_127_3477_U364 ( .A(DP_OP_425J2_127_3477_n402), .B(
        DP_OP_425J2_127_3477_n400), .CI(DP_OP_425J2_127_3477_n369), .CO(
        DP_OP_425J2_127_3477_n364), .S(DP_OP_425J2_127_3477_n365) );
  FADDX1_HVT DP_OP_425J2_127_3477_U363 ( .A(DP_OP_425J2_127_3477_n398), .B(
        DP_OP_425J2_127_3477_n396), .CI(DP_OP_425J2_127_3477_n367), .CO(
        DP_OP_425J2_127_3477_n362), .S(DP_OP_425J2_127_3477_n363) );
  FADDX1_HVT DP_OP_425J2_127_3477_U362 ( .A(DP_OP_425J2_127_3477_n394), .B(
        DP_OP_425J2_127_3477_n392), .CI(DP_OP_425J2_127_3477_n365), .CO(
        DP_OP_425J2_127_3477_n360), .S(DP_OP_425J2_127_3477_n361) );
  FADDX1_HVT DP_OP_425J2_127_3477_U361 ( .A(DP_OP_425J2_127_3477_n390), .B(
        DP_OP_425J2_127_3477_n363), .CI(DP_OP_425J2_127_3477_n388), .CO(
        DP_OP_425J2_127_3477_n358), .S(DP_OP_425J2_127_3477_n359) );
  FADDX1_HVT DP_OP_425J2_127_3477_U360 ( .A(DP_OP_425J2_127_3477_n386), .B(
        DP_OP_425J2_127_3477_n361), .CI(DP_OP_425J2_127_3477_n384), .CO(
        DP_OP_425J2_127_3477_n356), .S(DP_OP_425J2_127_3477_n357) );
  FADDX1_HVT DP_OP_425J2_127_3477_U359 ( .A(DP_OP_425J2_127_3477_n382), .B(
        DP_OP_425J2_127_3477_n359), .CI(DP_OP_425J2_127_3477_n380), .CO(
        DP_OP_425J2_127_3477_n354), .S(DP_OP_425J2_127_3477_n355) );
  FADDX1_HVT DP_OP_425J2_127_3477_U358 ( .A(DP_OP_425J2_127_3477_n357), .B(
        DP_OP_425J2_127_3477_n378), .CI(DP_OP_425J2_127_3477_n355), .CO(
        DP_OP_425J2_127_3477_n352), .S(DP_OP_425J2_127_3477_n353) );
  FADDX1_HVT DP_OP_425J2_127_3477_U356 ( .A(DP_OP_425J2_127_3477_n1924), .B(
        DP_OP_425J2_127_3477_n370), .CI(DP_OP_425J2_127_3477_n368), .CO(
        DP_OP_425J2_127_3477_n348), .S(DP_OP_425J2_127_3477_n349) );
  FADDX1_HVT DP_OP_425J2_127_3477_U355 ( .A(DP_OP_425J2_127_3477_n366), .B(
        DP_OP_425J2_127_3477_n349), .CI(DP_OP_425J2_127_3477_n364), .CO(
        DP_OP_425J2_127_3477_n346), .S(DP_OP_425J2_127_3477_n347) );
  FADDX1_HVT DP_OP_425J2_127_3477_U354 ( .A(DP_OP_425J2_127_3477_n362), .B(
        DP_OP_425J2_127_3477_n360), .CI(DP_OP_425J2_127_3477_n347), .CO(
        DP_OP_425J2_127_3477_n344), .S(DP_OP_425J2_127_3477_n345) );
  FADDX1_HVT DP_OP_425J2_127_3477_U353 ( .A(DP_OP_425J2_127_3477_n358), .B(
        DP_OP_425J2_127_3477_n345), .CI(DP_OP_425J2_127_3477_n356), .CO(
        DP_OP_425J2_127_3477_n342), .S(DP_OP_425J2_127_3477_n343) );
  FADDX1_HVT DP_OP_425J2_127_3477_U352 ( .A(DP_OP_425J2_127_3477_n354), .B(
        DP_OP_425J2_127_3477_n343), .CI(DP_OP_425J2_127_3477_n352), .CO(
        DP_OP_425J2_127_3477_n340), .S(DP_OP_425J2_127_3477_n341) );
  FADDX1_HVT DP_OP_425J2_127_3477_U350 ( .A(DP_OP_425J2_127_3477_n339), .B(
        DP_OP_425J2_127_3477_n348), .CI(DP_OP_425J2_127_3477_n346), .CO(
        DP_OP_425J2_127_3477_n336), .S(DP_OP_425J2_127_3477_n337) );
  FADDX1_HVT DP_OP_425J2_127_3477_U349 ( .A(DP_OP_425J2_127_3477_n337), .B(
        DP_OP_425J2_127_3477_n344), .CI(DP_OP_425J2_127_3477_n342), .CO(
        DP_OP_425J2_127_3477_n334), .S(DP_OP_425J2_127_3477_n335) );
  FADDX1_HVT DP_OP_425J2_127_3477_U348 ( .A(DP_OP_425J2_127_3477_n1923), .B(
        DP_OP_425J2_127_3477_n338), .CI(DP_OP_425J2_127_3477_n336), .CO(
        DP_OP_425J2_127_3477_n332), .S(DP_OP_425J2_127_3477_n333) );
  FADDX1_HVT DP_OP_425J2_127_3477_U331 ( .A(DP_OP_425J2_127_3477_n1903), .B(
        DP_OP_425J2_127_3477_n1901), .CI(DP_OP_425J2_127_3477_n1899), .CO(
        DP_OP_425J2_127_3477_n269), .S(n_conv2_sum_d[0]) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U330 ( .A1(DP_OP_425J2_127_3477_n1837), 
        .A2(DP_OP_425J2_127_3477_n1839), .Y(DP_OP_425J2_127_3477_n268) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U329 ( .A1(DP_OP_425J2_127_3477_n1839), .A2(
        DP_OP_425J2_127_3477_n1837), .Y(DP_OP_425J2_127_3477_n267) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U323 ( .A1(DP_OP_425J2_127_3477_n1731), 
        .A2(DP_OP_425J2_127_3477_n1733), .Y(DP_OP_425J2_127_3477_n265) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U315 ( .A1(DP_OP_425J2_127_3477_n1577), 
        .A2(DP_OP_425J2_127_3477_n1579), .Y(DP_OP_425J2_127_3477_n260) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U309 ( .A1(DP_OP_425J2_127_3477_n1401), 
        .A2(DP_OP_425J2_127_3477_n1403), .Y(DP_OP_425J2_127_3477_n257) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U301 ( .A1(DP_OP_425J2_127_3477_n1213), 
        .A2(DP_OP_425J2_127_3477_n1215), .Y(DP_OP_425J2_127_3477_n252) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U295 ( .A1(DP_OP_425J2_127_3477_n1019), 
        .A2(DP_OP_425J2_127_3477_n1021), .Y(DP_OP_425J2_127_3477_n249) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U287 ( .A1(DP_OP_425J2_127_3477_n823), .A2(
        DP_OP_425J2_127_3477_n1018), .Y(DP_OP_425J2_127_3477_n244) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U274 ( .A1(DP_OP_425J2_127_3477_n513), .A2(
        DP_OP_425J2_127_3477_n648), .Y(DP_OP_425J2_127_3477_n237) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U257 ( .A1(DP_OP_425J2_127_3477_n373), .A2(
        DP_OP_425J2_127_3477_n418), .Y(DP_OP_425J2_127_3477_n226) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U245 ( .A1(DP_OP_425J2_127_3477_n351), .A2(
        DP_OP_425J2_127_3477_n372), .Y(DP_OP_425J2_127_3477_n217) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U235 ( .A1(DP_OP_425J2_127_3477_n350), .A2(
        DP_OP_425J2_127_3477_n341), .Y(DP_OP_425J2_127_3477_n210) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U234 ( .A1(DP_OP_425J2_127_3477_n341), .A2(
        DP_OP_425J2_127_3477_n350), .Y(DP_OP_425J2_127_3477_n209) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U225 ( .A1(DP_OP_425J2_127_3477_n340), .A2(
        DP_OP_425J2_127_3477_n335), .Y(DP_OP_425J2_127_3477_n203) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U217 ( .A1(DP_OP_425J2_127_3477_n334), .A2(
        DP_OP_425J2_127_3477_n333), .Y(DP_OP_425J2_127_3477_n198) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U216 ( .A1(DP_OP_425J2_127_3477_n333), .A2(
        DP_OP_425J2_127_3477_n334), .Y(DP_OP_425J2_127_3477_n197) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U214 ( .A1(DP_OP_425J2_127_3477_n286), .A2(
        DP_OP_425J2_127_3477_n198), .Y(DP_OP_425J2_127_3477_n22) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U210 ( .A1(DP_OP_425J2_127_3477_n287), .A2(
        DP_OP_425J2_127_3477_n286), .Y(DP_OP_425J2_127_3477_n189) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U201 ( .A1(DP_OP_425J2_127_3477_n332), .A2(
        n1381), .Y(DP_OP_425J2_127_3477_n185) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U194 ( .A1(DP_OP_425J2_127_3477_n182), .A2(
        DP_OP_425J2_127_3477_n189), .Y(DP_OP_425J2_127_3477_n176) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U187 ( .A1(DP_OP_425J2_127_3477_n329), .A2(
        DP_OP_425J2_127_3477_n330), .Y(DP_OP_425J2_127_3477_n174) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U186 ( .A1(DP_OP_425J2_127_3477_n330), .A2(
        DP_OP_425J2_127_3477_n329), .Y(DP_OP_425J2_127_3477_n171) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U177 ( .A1(DP_OP_425J2_127_3477_n327), .A2(
        DP_OP_425J2_127_3477_n328), .Y(DP_OP_425J2_127_3477_n167) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U176 ( .A1(DP_OP_425J2_127_3477_n328), .A2(
        DP_OP_425J2_127_3477_n327), .Y(DP_OP_425J2_127_3477_n166) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U174 ( .A1(DP_OP_425J2_127_3477_n283), .A2(
        DP_OP_425J2_127_3477_n167), .Y(DP_OP_425J2_127_3477_n19) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U172 ( .A1(DP_OP_425J2_127_3477_n166), .A2(
        DP_OP_425J2_127_3477_n171), .Y(DP_OP_425J2_127_3477_n162) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U168 ( .A1(DP_OP_425J2_127_3477_n176), .A2(
        DP_OP_425J2_127_3477_n162), .Y(DP_OP_425J2_127_3477_n160) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U163 ( .A1(DP_OP_425J2_127_3477_n325), .A2(
        DP_OP_425J2_127_3477_n326), .Y(DP_OP_425J2_127_3477_n156) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U162 ( .A1(DP_OP_425J2_127_3477_n326), .A2(
        DP_OP_425J2_127_3477_n325), .Y(DP_OP_425J2_127_3477_n153) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U153 ( .A1(DP_OP_425J2_127_3477_n323), .A2(
        DP_OP_425J2_127_3477_n324), .Y(DP_OP_425J2_127_3477_n149) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U152 ( .A1(DP_OP_425J2_127_3477_n324), .A2(
        DP_OP_425J2_127_3477_n323), .Y(DP_OP_425J2_127_3477_n148) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U150 ( .A1(DP_OP_425J2_127_3477_n281), .A2(
        DP_OP_425J2_127_3477_n149), .Y(DP_OP_425J2_127_3477_n17) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U148 ( .A1(DP_OP_425J2_127_3477_n148), .A2(
        DP_OP_425J2_127_3477_n153), .Y(DP_OP_425J2_127_3477_n146) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U146 ( .A1(DP_OP_425J2_127_3477_n162), .A2(
        DP_OP_425J2_127_3477_n146), .Y(DP_OP_425J2_127_3477_n144) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U142 ( .A1(DP_OP_425J2_127_3477_n176), .A2(
        DP_OP_425J2_127_3477_n142), .Y(DP_OP_425J2_127_3477_n140) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U137 ( .A1(DP_OP_425J2_127_3477_n321), .A2(
        DP_OP_425J2_127_3477_n322), .Y(DP_OP_425J2_127_3477_n136) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U136 ( .A1(DP_OP_425J2_127_3477_n322), .A2(
        DP_OP_425J2_127_3477_n321), .Y(DP_OP_425J2_127_3477_n133) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U127 ( .A1(DP_OP_425J2_127_3477_n319), .A2(
        DP_OP_425J2_127_3477_n320), .Y(DP_OP_425J2_127_3477_n129) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U126 ( .A1(DP_OP_425J2_127_3477_n320), .A2(
        DP_OP_425J2_127_3477_n319), .Y(DP_OP_425J2_127_3477_n128) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U124 ( .A1(DP_OP_425J2_127_3477_n279), .A2(
        DP_OP_425J2_127_3477_n129), .Y(DP_OP_425J2_127_3477_n15) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U122 ( .A1(DP_OP_425J2_127_3477_n128), .A2(
        DP_OP_425J2_127_3477_n133), .Y(DP_OP_425J2_127_3477_n126) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U115 ( .A1(DP_OP_425J2_127_3477_n317), .A2(
        DP_OP_425J2_127_3477_n318), .Y(DP_OP_425J2_127_3477_n120) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U108 ( .A1(DP_OP_425J2_127_3477_n126), .A2(
        n1842), .Y(DP_OP_425J2_127_3477_n115) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U102 ( .A1(DP_OP_425J2_127_3477_n176), .A2(
        DP_OP_425J2_127_3477_n111), .Y(DP_OP_425J2_127_3477_n109) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U97 ( .A1(DP_OP_425J2_127_3477_n315), .A2(
        DP_OP_425J2_127_3477_n316), .Y(DP_OP_425J2_127_3477_n105) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U96 ( .A1(DP_OP_425J2_127_3477_n316), .A2(
        DP_OP_425J2_127_3477_n315), .Y(DP_OP_425J2_127_3477_n102) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U94 ( .A1(DP_OP_425J2_127_3477_n277), .A2(
        DP_OP_425J2_127_3477_n105), .Y(DP_OP_425J2_127_3477_n13) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U87 ( .A1(DP_OP_425J2_127_3477_n313), .A2(
        DP_OP_425J2_127_3477_n314), .Y(DP_OP_425J2_127_3477_n98) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U86 ( .A1(DP_OP_425J2_127_3477_n314), .A2(
        DP_OP_425J2_127_3477_n313), .Y(DP_OP_425J2_127_3477_n97) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U84 ( .A1(DP_OP_425J2_127_3477_n276), .A2(
        DP_OP_425J2_127_3477_n98), .Y(DP_OP_425J2_127_3477_n12) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U82 ( .A1(DP_OP_425J2_127_3477_n97), .A2(
        DP_OP_425J2_127_3477_n102), .Y(DP_OP_425J2_127_3477_n95) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U75 ( .A1(DP_OP_425J2_127_3477_n311), .A2(
        DP_OP_425J2_127_3477_n312), .Y(DP_OP_425J2_127_3477_n89) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U68 ( .A1(DP_OP_425J2_127_3477_n95), .A2(
        n1841), .Y(DP_OP_425J2_127_3477_n82) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U61 ( .A1(DP_OP_425J2_127_3477_n309), .A2(
        DP_OP_425J2_127_3477_n310), .Y(DP_OP_425J2_127_3477_n78) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U60 ( .A1(DP_OP_425J2_127_3477_n310), .A2(
        DP_OP_425J2_127_3477_n309), .Y(DP_OP_425J2_127_3477_n77) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U54 ( .A1(DP_OP_425J2_127_3477_n111), .A2(
        DP_OP_425J2_127_3477_n75), .Y(DP_OP_425J2_127_3477_n73) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U45 ( .A1(DP_OP_425J2_127_3477_n307), .A2(
        DP_OP_425J2_127_3477_n308), .Y(DP_OP_425J2_127_3477_n65) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U38 ( .A1(DP_OP_425J2_127_3477_n71), .A2(
        n1836), .Y(DP_OP_425J2_127_3477_n60) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U34 ( .A1(DP_OP_425J2_127_3477_n287), .A2(
        DP_OP_425J2_127_3477_n58), .Y(DP_OP_425J2_127_3477_n56) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U29 ( .A1(DP_OP_425J2_127_3477_n305), .A2(
        DP_OP_425J2_127_3477_n306), .Y(DP_OP_425J2_127_3477_n52) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U28 ( .A1(DP_OP_425J2_127_3477_n306), .A2(
        DP_OP_425J2_127_3477_n305), .Y(DP_OP_425J2_127_3477_n51) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U21 ( .A1(DP_OP_425J2_127_3477_n303), .A2(
        DP_OP_425J2_127_3477_n304), .Y(DP_OP_425J2_127_3477_n47) );
  NAND2X0_HVT DP_OP_425J2_127_3477_U9 ( .A1(n1834), .A2(
        DP_OP_425J2_127_3477_n302), .Y(DP_OP_425J2_127_3477_n38) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U200 ( .A1(DP_OP_424J2_126_3477_n331), .A2(
        DP_OP_424J2_126_3477_n332), .Y(DP_OP_424J2_126_3477_n182) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U325 ( .A1(DP_OP_424J2_126_3477_n5), .A2(
        DP_OP_424J2_126_3477_n267), .A3(DP_OP_424J2_126_3477_n268), .Y(
        DP_OP_424J2_126_3477_n266) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U173 ( .A1(DP_OP_424J2_126_3477_n174), .A2(
        DP_OP_424J2_126_3477_n166), .A3(DP_OP_424J2_126_3477_n167), .Y(
        DP_OP_424J2_126_3477_n165) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U83 ( .A1(DP_OP_424J2_126_3477_n105), .A2(
        DP_OP_424J2_126_3477_n97), .A3(DP_OP_424J2_126_3477_n98), .Y(
        DP_OP_424J2_126_3477_n96) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U123 ( .A1(DP_OP_424J2_126_3477_n136), .A2(
        DP_OP_424J2_126_3477_n128), .A3(DP_OP_424J2_126_3477_n129), .Y(
        DP_OP_424J2_126_3477_n127) );
  XNOR2X1_HVT DP_OP_424J2_126_3477_U787 ( .A1(DP_OP_424J2_126_3477_n2502), 
        .A2(DP_OP_424J2_126_3477_n3029), .Y(DP_OP_424J2_126_3477_n1211) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2291 ( .A1(DP_OP_424J2_126_3477_n3058), 
        .A2(n34), .Y(DP_OP_424J2_126_3477_n3050) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2290 ( .A1(DP_OP_424J2_126_3477_n3057), 
        .A2(n34), .Y(DP_OP_424J2_126_3477_n3049) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2289 ( .A1(DP_OP_425J2_127_3477_n2002), .A2(
        n693), .Y(DP_OP_424J2_126_3477_n3048) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2273 ( .A1(DP_OP_425J2_127_3477_n2002), .A2(
        DP_OP_424J2_126_3477_n3065), .Y(DP_OP_424J2_126_3477_n3032) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2271 ( .A1(DP_OP_425J2_127_3477_n2008), .A2(
        n213), .Y(DP_OP_424J2_126_3477_n3031) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2270 ( .A1(DP_OP_425J2_127_3477_n2007), .A2(
        n213), .Y(DP_OP_424J2_126_3477_n3030) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2269 ( .A1(DP_OP_424J2_126_3477_n3060), .A2(
        n215), .Y(DP_OP_424J2_126_3477_n3029) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2268 ( .A1(DP_OP_424J2_126_3477_n3059), .A2(
        n215), .Y(DP_OP_424J2_126_3477_n3028) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2267 ( .A1(DP_OP_424J2_126_3477_n3058), .A2(
        n210), .Y(DP_OP_424J2_126_3477_n820) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2266 ( .A1(DP_OP_424J2_126_3477_n3057), .A2(
        n213), .Y(DP_OP_424J2_126_3477_n3027) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2265 ( .A1(DP_OP_425J2_127_3477_n2002), 
        .A2(n212), .Y(DP_OP_424J2_126_3477_n3026) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2246 ( .A1(DP_OP_424J2_126_3477_n3015), 
        .A2(n846), .Y(DP_OP_424J2_126_3477_n3007) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2245 ( .A1(DP_OP_425J2_127_3477_n2046), .A2(
        DP_OP_424J2_126_3477_n3025), .Y(DP_OP_424J2_126_3477_n3006) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2238 ( .A1(DP_OP_424J2_126_3477_n3015), 
        .A2(n704), .Y(DP_OP_424J2_126_3477_n2999) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2237 ( .A1(DP_OP_425J2_127_3477_n2046), .A2(
        n704), .Y(DP_OP_424J2_126_3477_n2998) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2227 ( .A1(DP_OP_424J2_126_3477_n3020), .A2(
        n1507), .Y(DP_OP_424J2_126_3477_n2988) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2201 ( .A1(DP_OP_424J2_126_3477_n2970), .A2(
        n677), .Y(DP_OP_424J2_126_3477_n2962) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2193 ( .A1(DP_OP_424J2_126_3477_n2970), .A2(
        DP_OP_422J2_124_3477_n2980), .Y(DP_OP_424J2_126_3477_n2954) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2186 ( .A1(DP_OP_424J2_126_3477_n2971), 
        .A2(DP_OP_424J2_126_3477_n2979), .Y(DP_OP_424J2_126_3477_n2947) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2185 ( .A1(DP_OP_424J2_126_3477_n2970), .A2(
        DP_OP_424J2_126_3477_n2979), .Y(DP_OP_424J2_126_3477_n2946) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2184 ( .A1(DP_OP_424J2_126_3477_n2977), .A2(
        n254), .Y(DP_OP_424J2_126_3477_n2945) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2182 ( .A1(DP_OP_424J2_126_3477_n2975), .A2(
        n254), .Y(DP_OP_424J2_126_3477_n2943) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2181 ( .A1(DP_OP_424J2_126_3477_n2974), .A2(
        n254), .Y(DP_OP_424J2_126_3477_n2942) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2157 ( .A1(DP_OP_423J2_125_3477_n3014), .A2(
        n446), .Y(DP_OP_424J2_126_3477_n2918) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2149 ( .A1(DP_OP_423J2_125_3477_n3014), .A2(
        DP_OP_424J2_126_3477_n2936), .Y(DP_OP_424J2_126_3477_n2910) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2140 ( .A1(DP_OP_424J2_126_3477_n2933), .A2(
        n35), .Y(DP_OP_424J2_126_3477_n2901) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2139 ( .A1(DP_OP_424J2_126_3477_n2932), .A2(
        n35), .Y(DP_OP_424J2_126_3477_n2900) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2138 ( .A1(DP_OP_422J2_124_3477_n2007), .A2(
        n604), .Y(DP_OP_424J2_126_3477_n2899) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2137 ( .A1(DP_OP_422J2_124_3477_n2006), .A2(
        n35), .Y(DP_OP_424J2_126_3477_n2898) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2136 ( .A1(DP_OP_424J2_126_3477_n2929), .A2(
        n35), .Y(DP_OP_424J2_126_3477_n2897) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2135 ( .A1(DP_OP_424J2_126_3477_n2928), .A2(
        n35), .Y(DP_OP_424J2_126_3477_n2896) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2134 ( .A1(DP_OP_424J2_126_3477_n2927), .A2(
        n600), .Y(DP_OP_424J2_126_3477_n2895) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2133 ( .A1(DP_OP_423J2_125_3477_n3014), 
        .A2(n602), .Y(DP_OP_424J2_126_3477_n2894) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2114 ( .A1(DP_OP_424J2_126_3477_n2883), 
        .A2(DP_OP_424J2_126_3477_n2893), .Y(DP_OP_424J2_126_3477_n2875) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2113 ( .A1(DP_OP_424J2_126_3477_n2882), .A2(
        DP_OP_424J2_126_3477_n2893), .Y(DP_OP_424J2_126_3477_n2874) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2105 ( .A1(DP_OP_424J2_126_3477_n2882), .A2(
        DP_OP_423J2_125_3477_n2892), .Y(DP_OP_424J2_126_3477_n2866) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2098 ( .A1(DP_OP_424J2_126_3477_n2883), 
        .A2(DP_OP_423J2_125_3477_n2891), .Y(DP_OP_424J2_126_3477_n2859) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2097 ( .A1(DP_OP_424J2_126_3477_n2882), .A2(
        DP_OP_423J2_125_3477_n2891), .Y(DP_OP_424J2_126_3477_n2858) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2096 ( .A1(DP_OP_424J2_126_3477_n2889), .A2(
        DP_OP_422J2_124_3477_n2890), .Y(DP_OP_424J2_126_3477_n2857) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2095 ( .A1(DP_OP_423J2_125_3477_n2976), .A2(
        DP_OP_422J2_124_3477_n2890), .Y(DP_OP_424J2_126_3477_n2856) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2093 ( .A1(DP_OP_424J2_126_3477_n2886), .A2(
        DP_OP_424J2_126_3477_n2890), .Y(DP_OP_424J2_126_3477_n2854) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2092 ( .A1(DP_OP_423J2_125_3477_n2973), .A2(
        DP_OP_424J2_126_3477_n2890), .Y(DP_OP_424J2_126_3477_n2853) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2091 ( .A1(DP_OP_425J2_127_3477_n2180), .A2(
        DP_OP_422J2_124_3477_n2890), .Y(DP_OP_424J2_126_3477_n2852) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2090 ( .A1(DP_OP_424J2_126_3477_n2883), .A2(
        DP_OP_424J2_126_3477_n2890), .Y(DP_OP_424J2_126_3477_n2851) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2089 ( .A1(DP_OP_424J2_126_3477_n2882), 
        .A2(DP_OP_424J2_126_3477_n2890), .Y(DP_OP_424J2_126_3477_n2850) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2069 ( .A1(DP_OP_422J2_124_3477_n2090), .A2(
        DP_OP_424J2_126_3477_n2849), .Y(DP_OP_424J2_126_3477_n2830) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2055 ( .A1(DP_OP_422J2_124_3477_n2092), 
        .A2(n1438), .Y(DP_OP_424J2_126_3477_n2816) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2054 ( .A1(DP_OP_422J2_124_3477_n2091), 
        .A2(DP_OP_422J2_124_3477_n2847), .Y(DP_OP_424J2_126_3477_n2815) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2052 ( .A1(DP_OP_424J2_126_3477_n2845), .A2(
        DP_OP_424J2_126_3477_n2846), .Y(DP_OP_424J2_126_3477_n2813) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2051 ( .A1(DP_OP_423J2_125_3477_n2932), .A2(
        DP_OP_424J2_126_3477_n2846), .Y(DP_OP_424J2_126_3477_n2812) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2050 ( .A1(DP_OP_423J2_125_3477_n2931), .A2(
        DP_OP_424J2_126_3477_n2846), .Y(DP_OP_424J2_126_3477_n2811) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2049 ( .A1(DP_OP_425J2_127_3477_n2226), .A2(
        DP_OP_424J2_126_3477_n2846), .Y(DP_OP_424J2_126_3477_n2810) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2048 ( .A1(DP_OP_422J2_124_3477_n2093), .A2(
        DP_OP_424J2_126_3477_n2846), .Y(DP_OP_424J2_126_3477_n2809) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2047 ( .A1(DP_OP_422J2_124_3477_n2092), .A2(
        DP_OP_424J2_126_3477_n2846), .Y(DP_OP_424J2_126_3477_n2808) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2046 ( .A1(DP_OP_422J2_124_3477_n2091), .A2(
        DP_OP_424J2_126_3477_n2846), .Y(DP_OP_424J2_126_3477_n2807) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2045 ( .A1(DP_OP_422J2_124_3477_n2090), 
        .A2(DP_OP_424J2_126_3477_n2846), .Y(DP_OP_424J2_126_3477_n2806) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2026 ( .A1(DP_OP_424J2_126_3477_n2795), 
        .A2(DP_OP_424J2_126_3477_n2805), .Y(DP_OP_424J2_126_3477_n2787) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2025 ( .A1(DP_OP_424J2_126_3477_n2794), .A2(
        DP_OP_424J2_126_3477_n2805), .Y(DP_OP_424J2_126_3477_n2786) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2022 ( .A1(DP_OP_424J2_126_3477_n2799), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_424J2_126_3477_n2783) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2013 ( .A1(DP_OP_423J2_125_3477_n2886), 
        .A2(n1444), .Y(DP_OP_424J2_126_3477_n2774) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2011 ( .A1(DP_OP_424J2_126_3477_n2796), 
        .A2(n1444), .Y(DP_OP_424J2_126_3477_n2772) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2010 ( .A1(DP_OP_424J2_126_3477_n2795), 
        .A2(DP_OP_423J2_125_3477_n2803), .Y(DP_OP_424J2_126_3477_n2771) );
  OR2X1_HVT DP_OP_424J2_126_3477_U2008 ( .A1(DP_OP_424J2_126_3477_n2801), .A2(
        DP_OP_424J2_126_3477_n2802), .Y(DP_OP_424J2_126_3477_n2769) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1982 ( .A1(DP_OP_422J2_124_3477_n2179), 
        .A2(n66), .Y(DP_OP_424J2_126_3477_n2743) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1981 ( .A1(DP_OP_422J2_124_3477_n2178), .A2(
        n66), .Y(DP_OP_424J2_126_3477_n2742) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1964 ( .A1(DP_OP_422J2_124_3477_n2185), .A2(
        DP_OP_424J2_126_3477_n2758), .Y(DP_OP_424J2_126_3477_n2725) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1963 ( .A1(DP_OP_424J2_126_3477_n2756), .A2(
        DP_OP_424J2_126_3477_n2758), .Y(DP_OP_424J2_126_3477_n2724) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1961 ( .A1(DP_OP_424J2_126_3477_n2754), .A2(
        DP_OP_424J2_126_3477_n2758), .Y(DP_OP_424J2_126_3477_n2722) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1930 ( .A1(DP_OP_423J2_125_3477_n2795), 
        .A2(n1342), .Y(DP_OP_424J2_126_3477_n2691) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1929 ( .A1(DP_OP_422J2_124_3477_n2222), .A2(
        n1342), .Y(DP_OP_424J2_126_3477_n2690) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1923 ( .A1(DP_OP_425J2_127_3477_n2356), 
        .A2(DP_OP_422J2_124_3477_n2715), .Y(DP_OP_424J2_126_3477_n2684) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1885 ( .A1(DP_OP_423J2_125_3477_n2750), .A2(
        n279), .Y(DP_OP_424J2_126_3477_n2646) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1884 ( .A1(DP_OP_424J2_126_3477_n2669), 
        .A2(DP_OP_425J2_127_3477_n2671), .Y(DP_OP_424J2_126_3477_n2645) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1881 ( .A1(DP_OP_422J2_124_3477_n2270), 
        .A2(DP_OP_425J2_127_3477_n2671), .Y(DP_OP_424J2_126_3477_n2642) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1879 ( .A1(DP_OP_422J2_124_3477_n2268), 
        .A2(DP_OP_425J2_127_3477_n2671), .Y(DP_OP_424J2_126_3477_n2640) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1850 ( .A1(DP_OP_424J2_126_3477_n2619), 
        .A2(DP_OP_424J2_126_3477_n2629), .Y(DP_OP_424J2_126_3477_n2611) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1849 ( .A1(DP_OP_423J2_125_3477_n2706), .A2(
        DP_OP_424J2_126_3477_n2629), .Y(DP_OP_424J2_126_3477_n2610) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1834 ( .A1(DP_OP_424J2_126_3477_n2619), 
        .A2(DP_OP_424J2_126_3477_n2627), .Y(DP_OP_424J2_126_3477_n2595) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1833 ( .A1(DP_OP_422J2_124_3477_n2310), .A2(
        DP_OP_424J2_126_3477_n2627), .Y(DP_OP_424J2_126_3477_n2594) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1832 ( .A1(DP_OP_425J2_127_3477_n2449), .A2(
        n1331), .Y(DP_OP_424J2_126_3477_n2593) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1806 ( .A1(DP_OP_424J2_126_3477_n2575), 
        .A2(DP_OP_422J2_124_3477_n2585), .Y(DP_OP_424J2_126_3477_n2567) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1797 ( .A1(DP_OP_424J2_126_3477_n2574), .A2(
        n186), .Y(DP_OP_424J2_126_3477_n2558) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1788 ( .A1(DP_OP_423J2_125_3477_n2669), .A2(
        n424), .Y(DP_OP_424J2_126_3477_n2549) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1787 ( .A1(DP_OP_424J2_126_3477_n2580), .A2(
        n424), .Y(DP_OP_424J2_126_3477_n2548) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1786 ( .A1(DP_OP_424J2_126_3477_n2579), .A2(
        DP_OP_424J2_126_3477_n2582), .Y(DP_OP_424J2_126_3477_n2547) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1785 ( .A1(DP_OP_423J2_125_3477_n2666), .A2(
        n424), .Y(DP_OP_424J2_126_3477_n2546) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1784 ( .A1(DP_OP_423J2_125_3477_n2665), .A2(
        n424), .Y(DP_OP_424J2_126_3477_n2545) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1783 ( .A1(DP_OP_424J2_126_3477_n2576), .A2(
        n424), .Y(DP_OP_424J2_126_3477_n2544) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1782 ( .A1(DP_OP_424J2_126_3477_n2575), .A2(
        DP_OP_424J2_126_3477_n2582), .Y(DP_OP_424J2_126_3477_n2543) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1781 ( .A1(DP_OP_424J2_126_3477_n2574), 
        .A2(n424), .Y(DP_OP_424J2_126_3477_n2542) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1761 ( .A1(DP_OP_422J2_124_3477_n2398), .A2(
        DP_OP_424J2_126_3477_n2541), .Y(DP_OP_424J2_126_3477_n2522) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1754 ( .A1(DP_OP_422J2_124_3477_n2399), 
        .A2(DP_OP_424J2_126_3477_n2540), .Y(DP_OP_424J2_126_3477_n2515) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1745 ( .A1(DP_OP_422J2_124_3477_n2398), .A2(
        n772), .Y(DP_OP_424J2_126_3477_n2506) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1744 ( .A1(DP_OP_422J2_124_3477_n2405), .A2(
        n1337), .Y(DP_OP_424J2_126_3477_n2505) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1743 ( .A1(DP_OP_422J2_124_3477_n2404), .A2(
        n1335), .Y(DP_OP_424J2_126_3477_n2504) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1742 ( .A1(DP_OP_424J2_126_3477_n2535), .A2(
        n1334), .Y(DP_OP_424J2_126_3477_n2503) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1741 ( .A1(DP_OP_424J2_126_3477_n2534), .A2(
        n1362), .Y(DP_OP_424J2_126_3477_n2502) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1740 ( .A1(DP_OP_422J2_124_3477_n2401), .A2(
        n1335), .Y(DP_OP_424J2_126_3477_n2501) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1739 ( .A1(DP_OP_424J2_126_3477_n2532), .A2(
        n1334), .Y(DP_OP_424J2_126_3477_n2500) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1738 ( .A1(DP_OP_422J2_124_3477_n2399), .A2(
        n1336), .Y(DP_OP_424J2_126_3477_n2499) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1737 ( .A1(DP_OP_422J2_124_3477_n2398), 
        .A2(n1337), .Y(DP_OP_424J2_126_3477_n2498) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1717 ( .A1(DP_OP_424J2_126_3477_n2486), .A2(
        DP_OP_424J2_126_3477_n2497), .Y(DP_OP_424J2_126_3477_n2478) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1709 ( .A1(DP_OP_424J2_126_3477_n2486), .A2(
        n1491), .Y(DP_OP_424J2_126_3477_n2470) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1665 ( .A1(DP_OP_425J2_127_3477_n2574), .A2(
        DP_OP_423J2_125_3477_n2452), .Y(DP_OP_424J2_126_3477_n2426) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1631 ( .A1(DP_OP_424J2_126_3477_n2400), 
        .A2(DP_OP_423J2_125_3477_n2409), .Y(DP_OP_424J2_126_3477_n2392) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1614 ( .A1(DP_OP_422J2_124_3477_n2751), 
        .A2(n799), .Y(DP_OP_424J2_126_3477_n2375) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1613 ( .A1(DP_OP_422J2_124_3477_n2750), .A2(
        n799), .Y(DP_OP_424J2_126_3477_n2374) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1612 ( .A1(DP_OP_424J2_126_3477_n2405), .A2(
        n1433), .Y(DP_OP_424J2_126_3477_n2373) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1587 ( .A1(DP_OP_422J2_124_3477_n2796), 
        .A2(DP_OP_424J2_126_3477_n2365), .Y(DP_OP_424J2_126_3477_n2348) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1585 ( .A1(DP_OP_424J2_126_3477_n2354), .A2(
        DP_OP_425J2_127_3477_n2365), .Y(DP_OP_424J2_126_3477_n2346) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1577 ( .A1(DP_OP_424J2_126_3477_n2354), .A2(
        n1386), .Y(DP_OP_424J2_126_3477_n2338) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1542 ( .A1(DP_OP_424J2_126_3477_n2311), 
        .A2(DP_OP_425J2_127_3477_n2321), .Y(DP_OP_424J2_126_3477_n2303) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1541 ( .A1(DP_OP_423J2_125_3477_n2222), .A2(
        DP_OP_425J2_127_3477_n2321), .Y(DP_OP_424J2_126_3477_n2302) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1536 ( .A1(DP_OP_423J2_125_3477_n2225), 
        .A2(DP_OP_422J2_124_3477_n2320), .Y(DP_OP_424J2_126_3477_n2297) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1525 ( .A1(DP_OP_423J2_125_3477_n2222), .A2(
        n316), .Y(DP_OP_424J2_126_3477_n2286) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1524 ( .A1(DP_OP_424J2_126_3477_n2317), .A2(
        DP_OP_424J2_126_3477_n2318), .Y(DP_OP_424J2_126_3477_n2285) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1523 ( .A1(DP_OP_425J2_127_3477_n2712), .A2(
        DP_OP_424J2_126_3477_n2318), .Y(DP_OP_424J2_126_3477_n2284) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1522 ( .A1(DP_OP_424J2_126_3477_n2315), .A2(
        DP_OP_424J2_126_3477_n2318), .Y(DP_OP_424J2_126_3477_n2283) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1521 ( .A1(DP_OP_425J2_127_3477_n2710), .A2(
        DP_OP_424J2_126_3477_n2318), .Y(DP_OP_424J2_126_3477_n2282) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1520 ( .A1(DP_OP_423J2_125_3477_n2225), .A2(
        DP_OP_424J2_126_3477_n2318), .Y(DP_OP_424J2_126_3477_n2281) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1519 ( .A1(DP_OP_422J2_124_3477_n2840), .A2(
        DP_OP_424J2_126_3477_n2318), .Y(DP_OP_424J2_126_3477_n2280) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1518 ( .A1(DP_OP_424J2_126_3477_n2311), .A2(
        DP_OP_424J2_126_3477_n2318), .Y(DP_OP_424J2_126_3477_n2279) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1517 ( .A1(DP_OP_422J2_124_3477_n2838), 
        .A2(DP_OP_424J2_126_3477_n2318), .Y(DP_OP_424J2_126_3477_n2278) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1497 ( .A1(DP_OP_422J2_124_3477_n2882), .A2(
        DP_OP_424J2_126_3477_n2277), .Y(DP_OP_424J2_126_3477_n2258) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1489 ( .A1(DP_OP_422J2_124_3477_n2882), .A2(
        DP_OP_424J2_126_3477_n2276), .Y(DP_OP_424J2_126_3477_n2250) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1481 ( .A1(DP_OP_422J2_124_3477_n2882), .A2(
        DP_OP_424J2_126_3477_n2275), .Y(DP_OP_424J2_126_3477_n2242) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1480 ( .A1(DP_OP_423J2_125_3477_n2185), .A2(
        n1338), .Y(DP_OP_424J2_126_3477_n2241) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1479 ( .A1(DP_OP_422J2_124_3477_n2888), .A2(
        n1370), .Y(DP_OP_424J2_126_3477_n2240) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1478 ( .A1(DP_OP_425J2_127_3477_n2755), .A2(
        n1338), .Y(DP_OP_424J2_126_3477_n2239) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1477 ( .A1(DP_OP_423J2_125_3477_n2182), .A2(
        n1338), .Y(DP_OP_424J2_126_3477_n2238) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1476 ( .A1(DP_OP_424J2_126_3477_n2269), .A2(
        DP_OP_424J2_126_3477_n2274), .Y(DP_OP_424J2_126_3477_n2237) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1475 ( .A1(DP_OP_424J2_126_3477_n2268), .A2(
        n1370), .Y(DP_OP_424J2_126_3477_n2236) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1474 ( .A1(DP_OP_424J2_126_3477_n2267), .A2(
        n1370), .Y(DP_OP_424J2_126_3477_n2235) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1473 ( .A1(DP_OP_423J2_125_3477_n2178), 
        .A2(n1338), .Y(DP_OP_424J2_126_3477_n2234) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1454 ( .A1(DP_OP_422J2_124_3477_n2927), 
        .A2(DP_OP_423J2_125_3477_n2233), .Y(DP_OP_424J2_126_3477_n2215) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1453 ( .A1(DP_OP_424J2_126_3477_n2222), .A2(
        DP_OP_423J2_125_3477_n2233), .Y(DP_OP_424J2_126_3477_n2214) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1445 ( .A1(DP_OP_424J2_126_3477_n2222), .A2(
        n365), .Y(DP_OP_424J2_126_3477_n2206) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1435 ( .A1(DP_OP_423J2_125_3477_n2140), .A2(
        DP_OP_425J2_127_3477_n2230), .Y(DP_OP_424J2_126_3477_n2196) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1434 ( .A1(DP_OP_425J2_127_3477_n2799), .A2(
        DP_OP_422J2_124_3477_n2230), .Y(DP_OP_424J2_126_3477_n2195) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1433 ( .A1(DP_OP_422J2_124_3477_n2930), .A2(
        DP_OP_423J2_125_3477_n2230), .Y(DP_OP_424J2_126_3477_n2194) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1432 ( .A1(DP_OP_425J2_127_3477_n2797), .A2(
        DP_OP_423J2_125_3477_n2230), .Y(DP_OP_424J2_126_3477_n2193) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1431 ( .A1(DP_OP_425J2_127_3477_n2796), .A2(
        DP_OP_423J2_125_3477_n2230), .Y(DP_OP_424J2_126_3477_n2192) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1430 ( .A1(DP_OP_423J2_125_3477_n2135), .A2(
        DP_OP_425J2_127_3477_n2230), .Y(DP_OP_424J2_126_3477_n2191) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1429 ( .A1(DP_OP_424J2_126_3477_n2222), 
        .A2(DP_OP_422J2_124_3477_n2230), .Y(DP_OP_424J2_126_3477_n2190) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1409 ( .A1(DP_OP_422J2_124_3477_n2970), .A2(
        DP_OP_424J2_126_3477_n2189), .Y(DP_OP_424J2_126_3477_n2170) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1401 ( .A1(DP_OP_422J2_124_3477_n2970), .A2(
        n1344), .Y(DP_OP_424J2_126_3477_n2162) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1394 ( .A1(DP_OP_422J2_124_3477_n2971), 
        .A2(n1339), .Y(DP_OP_424J2_126_3477_n2155) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1393 ( .A1(DP_OP_422J2_124_3477_n2970), .A2(
        n1339), .Y(DP_OP_424J2_126_3477_n2154) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1392 ( .A1(DP_OP_424J2_126_3477_n2185), .A2(
        DP_OP_424J2_126_3477_n2186), .Y(DP_OP_424J2_126_3477_n2153) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1391 ( .A1(DP_OP_424J2_126_3477_n2184), .A2(
        DP_OP_422J2_124_3477_n2186), .Y(DP_OP_424J2_126_3477_n2152) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1389 ( .A1(DP_OP_422J2_124_3477_n2974), .A2(
        DP_OP_422J2_124_3477_n2186), .Y(DP_OP_424J2_126_3477_n2150) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1388 ( .A1(DP_OP_422J2_124_3477_n2973), .A2(
        DP_OP_422J2_124_3477_n2186), .Y(DP_OP_424J2_126_3477_n2149) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1387 ( .A1(DP_OP_422J2_124_3477_n2972), .A2(
        DP_OP_422J2_124_3477_n2186), .Y(DP_OP_424J2_126_3477_n2148) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1386 ( .A1(DP_OP_422J2_124_3477_n2971), .A2(
        DP_OP_422J2_124_3477_n2186), .Y(DP_OP_424J2_126_3477_n2147) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1385 ( .A1(DP_OP_422J2_124_3477_n2970), 
        .A2(DP_OP_425J2_127_3477_n2186), .Y(DP_OP_424J2_126_3477_n2146) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1358 ( .A1(DP_OP_422J2_124_3477_n3015), 
        .A2(DP_OP_425J2_127_3477_n2144), .Y(DP_OP_424J2_126_3477_n2119) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1357 ( .A1(DP_OP_422J2_124_3477_n3014), .A2(
        DP_OP_422J2_124_3477_n2144), .Y(DP_OP_424J2_126_3477_n2118) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1349 ( .A1(DP_OP_425J2_127_3477_n2882), .A2(
        DP_OP_424J2_126_3477_n2143), .Y(DP_OP_424J2_126_3477_n2110) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1313 ( .A1(DP_OP_424J2_126_3477_n2090), .A2(
        DP_OP_423J2_125_3477_n2100), .Y(DP_OP_424J2_126_3477_n2074) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1306 ( .A1(DP_OP_423J2_125_3477_n2003), 
        .A2(DP_OP_424J2_126_3477_n2099), .Y(DP_OP_424J2_126_3477_n2067) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1305 ( .A1(DP_OP_424J2_126_3477_n2090), .A2(
        DP_OP_424J2_126_3477_n2099), .Y(DP_OP_424J2_126_3477_n2066) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1278 ( .A1(DP_OP_425J2_127_3477_n2971), 
        .A2(DP_OP_425J2_127_3477_n2057), .Y(DP_OP_424J2_126_3477_n2039) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1269 ( .A1(DP_OP_425J2_127_3477_n2970), .A2(
        DP_OP_424J2_126_3477_n2056), .Y(DP_OP_424J2_126_3477_n2030) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1262 ( .A1(DP_OP_425J2_127_3477_n2971), 
        .A2(DP_OP_424J2_126_3477_n2055), .Y(DP_OP_424J2_126_3477_n2023) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1261 ( .A1(DP_OP_425J2_127_3477_n2970), .A2(
        DP_OP_424J2_126_3477_n2055), .Y(DP_OP_424J2_126_3477_n2022) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1259 ( .A1(DP_OP_425J2_127_3477_n2976), .A2(
        n30), .Y(DP_OP_424J2_126_3477_n2020) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1258 ( .A1(DP_OP_424J2_126_3477_n2051), .A2(
        n779), .Y(DP_OP_424J2_126_3477_n2019) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1257 ( .A1(DP_OP_425J2_127_3477_n2974), .A2(
        n30), .Y(DP_OP_424J2_126_3477_n2018) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1256 ( .A1(DP_OP_425J2_127_3477_n2973), .A2(
        n30), .Y(DP_OP_424J2_126_3477_n2017) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1255 ( .A1(DP_OP_425J2_127_3477_n2972), .A2(
        n30), .Y(DP_OP_424J2_126_3477_n2016) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1254 ( .A1(DP_OP_425J2_127_3477_n2971), .A2(
        n775), .Y(DP_OP_424J2_126_3477_n2015) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1253 ( .A1(DP_OP_425J2_127_3477_n2970), 
        .A2(n30), .Y(DP_OP_424J2_126_3477_n2014) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1225 ( .A1(DP_OP_424J2_126_3477_n2002), .A2(
        n557), .Y(DP_OP_424J2_126_3477_n1986) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1217 ( .A1(DP_OP_424J2_126_3477_n2002), .A2(
        DP_OP_424J2_126_3477_n2011), .Y(DP_OP_424J2_126_3477_n1978) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1216 ( .A1(DP_OP_425J2_127_3477_n3021), .A2(
        DP_OP_424J2_126_3477_n2010), .Y(DP_OP_424J2_126_3477_n1977) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1215 ( .A1(DP_OP_425J2_127_3477_n3020), .A2(
        DP_OP_424J2_126_3477_n2010), .Y(DP_OP_424J2_126_3477_n1976) );
  OR2X1_HVT DP_OP_424J2_126_3477_U1214 ( .A1(DP_OP_425J2_127_3477_n3019), .A2(
        DP_OP_424J2_126_3477_n2010), .Y(DP_OP_424J2_126_3477_n1975) );
  HADDX1_HVT DP_OP_424J2_126_3477_U1143 ( .A0(DP_OP_424J2_126_3477_n1936), 
        .B0(DP_OP_424J2_126_3477_n2045), .C1(DP_OP_424J2_126_3477_n1920), .SO(
        DP_OP_424J2_126_3477_n1921) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1142 ( .A(DP_OP_424J2_126_3477_n2089), .B(
        DP_OP_424J2_126_3477_n2001), .CI(DP_OP_424J2_126_3477_n2133), .CO(
        DP_OP_424J2_126_3477_n1918), .S(DP_OP_424J2_126_3477_n1919) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1141 ( .A(DP_OP_424J2_126_3477_n2221), .B(
        DP_OP_424J2_126_3477_n2177), .CI(DP_OP_424J2_126_3477_n2265), .CO(
        DP_OP_424J2_126_3477_n1916), .S(DP_OP_424J2_126_3477_n1917) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1140 ( .A(DP_OP_424J2_126_3477_n2353), .B(
        DP_OP_424J2_126_3477_n2309), .CI(DP_OP_424J2_126_3477_n2397), .CO(
        DP_OP_424J2_126_3477_n1914), .S(DP_OP_424J2_126_3477_n1915) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1139 ( .A(DP_OP_424J2_126_3477_n2485), .B(
        DP_OP_424J2_126_3477_n2441), .CI(DP_OP_424J2_126_3477_n2529), .CO(
        DP_OP_424J2_126_3477_n1912), .S(DP_OP_424J2_126_3477_n1913) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1138 ( .A(DP_OP_424J2_126_3477_n2617), .B(
        DP_OP_424J2_126_3477_n2573), .CI(DP_OP_424J2_126_3477_n2661), .CO(
        DP_OP_424J2_126_3477_n1910), .S(DP_OP_424J2_126_3477_n1911) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1137 ( .A(DP_OP_424J2_126_3477_n2749), .B(
        DP_OP_424J2_126_3477_n2705), .CI(DP_OP_424J2_126_3477_n2793), .CO(
        DP_OP_424J2_126_3477_n1908), .S(DP_OP_424J2_126_3477_n1909) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1136 ( .A(DP_OP_424J2_126_3477_n3055), .B(
        DP_OP_424J2_126_3477_n2837), .CI(DP_OP_424J2_126_3477_n2881), .CO(
        DP_OP_424J2_126_3477_n1906), .S(DP_OP_424J2_126_3477_n1907) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1135 ( .A(DP_OP_424J2_126_3477_n3013), .B(
        DP_OP_424J2_126_3477_n2925), .CI(DP_OP_424J2_126_3477_n2969), .CO(
        DP_OP_424J2_126_3477_n1904), .S(DP_OP_424J2_126_3477_n1905) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1134 ( .A(DP_OP_424J2_126_3477_n1921), .B(
        DP_OP_424J2_126_3477_n1907), .CI(DP_OP_424J2_126_3477_n1909), .CO(
        DP_OP_424J2_126_3477_n1902), .S(DP_OP_424J2_126_3477_n1903) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1133 ( .A(DP_OP_424J2_126_3477_n1911), .B(
        DP_OP_424J2_126_3477_n1905), .CI(DP_OP_424J2_126_3477_n1913), .CO(
        DP_OP_424J2_126_3477_n1900), .S(DP_OP_424J2_126_3477_n1901) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1132 ( .A(DP_OP_424J2_126_3477_n1919), .B(
        DP_OP_424J2_126_3477_n1915), .CI(DP_OP_424J2_126_3477_n1917), .CO(
        DP_OP_424J2_126_3477_n1898), .S(DP_OP_424J2_126_3477_n1899) );
  HADDX1_HVT DP_OP_424J2_126_3477_U1131 ( .A0(DP_OP_424J2_126_3477_n1935), 
        .B0(DP_OP_424J2_126_3477_n2000), .C1(DP_OP_424J2_126_3477_n1896), .SO(
        DP_OP_424J2_126_3477_n1897) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1130 ( .A(DP_OP_424J2_126_3477_n2037), .B(
        DP_OP_424J2_126_3477_n1993), .CI(DP_OP_424J2_126_3477_n2044), .CO(
        DP_OP_424J2_126_3477_n1894), .S(DP_OP_424J2_126_3477_n1895) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1129 ( .A(DP_OP_424J2_126_3477_n2088), .B(
        DP_OP_424J2_126_3477_n2081), .CI(DP_OP_424J2_126_3477_n2125), .CO(
        DP_OP_424J2_126_3477_n1892), .S(DP_OP_424J2_126_3477_n1893) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1128 ( .A(DP_OP_424J2_126_3477_n2169), .B(
        DP_OP_424J2_126_3477_n2132), .CI(DP_OP_424J2_126_3477_n2176), .CO(
        DP_OP_424J2_126_3477_n1890), .S(DP_OP_424J2_126_3477_n1891) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1127 ( .A(DP_OP_424J2_126_3477_n2220), .B(
        DP_OP_424J2_126_3477_n2213), .CI(DP_OP_424J2_126_3477_n2257), .CO(
        DP_OP_424J2_126_3477_n1888), .S(DP_OP_424J2_126_3477_n1889) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1126 ( .A(DP_OP_424J2_126_3477_n2301), .B(
        DP_OP_424J2_126_3477_n2264), .CI(DP_OP_424J2_126_3477_n2308), .CO(
        DP_OP_424J2_126_3477_n1886), .S(DP_OP_424J2_126_3477_n1887) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1125 ( .A(DP_OP_424J2_126_3477_n2352), .B(
        DP_OP_424J2_126_3477_n2345), .CI(DP_OP_424J2_126_3477_n2389), .CO(
        DP_OP_424J2_126_3477_n1884), .S(DP_OP_424J2_126_3477_n1885) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1124 ( .A(DP_OP_424J2_126_3477_n2433), .B(
        DP_OP_424J2_126_3477_n2396), .CI(DP_OP_424J2_126_3477_n2440), .CO(
        DP_OP_424J2_126_3477_n1882), .S(DP_OP_424J2_126_3477_n1883) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1123 ( .A(DP_OP_424J2_126_3477_n2484), .B(
        DP_OP_424J2_126_3477_n2477), .CI(DP_OP_424J2_126_3477_n2521), .CO(
        DP_OP_424J2_126_3477_n1880), .S(DP_OP_424J2_126_3477_n1881) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1122 ( .A(DP_OP_424J2_126_3477_n2565), .B(
        DP_OP_424J2_126_3477_n2528), .CI(DP_OP_424J2_126_3477_n2572), .CO(
        DP_OP_424J2_126_3477_n1878), .S(DP_OP_424J2_126_3477_n1879) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1121 ( .A(DP_OP_424J2_126_3477_n3054), .B(
        DP_OP_424J2_126_3477_n2609), .CI(DP_OP_424J2_126_3477_n3047), .CO(
        DP_OP_424J2_126_3477_n1876), .S(DP_OP_424J2_126_3477_n1877) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1120 ( .A(DP_OP_424J2_126_3477_n2792), .B(
        DP_OP_424J2_126_3477_n2616), .CI(DP_OP_424J2_126_3477_n2653), .CO(
        DP_OP_424J2_126_3477_n1874), .S(DP_OP_424J2_126_3477_n1875) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1119 ( .A(DP_OP_424J2_126_3477_n2829), .B(
        DP_OP_424J2_126_3477_n3012), .CI(DP_OP_424J2_126_3477_n3005), .CO(
        DP_OP_424J2_126_3477_n1872), .S(DP_OP_424J2_126_3477_n1873) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1118 ( .A(DP_OP_424J2_126_3477_n2748), .B(
        DP_OP_424J2_126_3477_n2968), .CI(DP_OP_424J2_126_3477_n2961), .CO(
        DP_OP_424J2_126_3477_n1870), .S(DP_OP_424J2_126_3477_n1871) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1117 ( .A(DP_OP_424J2_126_3477_n2741), .B(
        DP_OP_424J2_126_3477_n2924), .CI(DP_OP_424J2_126_3477_n2660), .CO(
        DP_OP_424J2_126_3477_n1868), .S(DP_OP_424J2_126_3477_n1869) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1116 ( .A(DP_OP_424J2_126_3477_n2917), .B(
        DP_OP_424J2_126_3477_n2697), .CI(DP_OP_424J2_126_3477_n2704), .CO(
        DP_OP_424J2_126_3477_n1866), .S(DP_OP_424J2_126_3477_n1867) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1115 ( .A(DP_OP_424J2_126_3477_n2873), .B(
        DP_OP_424J2_126_3477_n2785), .CI(DP_OP_424J2_126_3477_n2836), .CO(
        DP_OP_424J2_126_3477_n1864), .S(DP_OP_424J2_126_3477_n1865) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1114 ( .A(DP_OP_424J2_126_3477_n2880), .B(
        DP_OP_424J2_126_3477_n1920), .CI(DP_OP_424J2_126_3477_n1897), .CO(
        DP_OP_424J2_126_3477_n1862), .S(DP_OP_424J2_126_3477_n1863) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1113 ( .A(DP_OP_424J2_126_3477_n1904), .B(
        DP_OP_424J2_126_3477_n1918), .CI(DP_OP_424J2_126_3477_n1916), .CO(
        DP_OP_424J2_126_3477_n1860), .S(DP_OP_424J2_126_3477_n1861) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1112 ( .A(DP_OP_424J2_126_3477_n1910), .B(
        DP_OP_424J2_126_3477_n1906), .CI(DP_OP_424J2_126_3477_n1914), .CO(
        DP_OP_424J2_126_3477_n1858), .S(DP_OP_424J2_126_3477_n1859) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1111 ( .A(DP_OP_424J2_126_3477_n1912), .B(
        DP_OP_424J2_126_3477_n1908), .CI(DP_OP_424J2_126_3477_n1865), .CO(
        DP_OP_424J2_126_3477_n1856), .S(DP_OP_424J2_126_3477_n1857) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1110 ( .A(DP_OP_424J2_126_3477_n1887), .B(
        DP_OP_424J2_126_3477_n1873), .CI(DP_OP_424J2_126_3477_n1871), .CO(
        DP_OP_424J2_126_3477_n1854), .S(DP_OP_424J2_126_3477_n1855) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1109 ( .A(DP_OP_424J2_126_3477_n1891), .B(
        DP_OP_424J2_126_3477_n1875), .CI(DP_OP_424J2_126_3477_n1879), .CO(
        DP_OP_424J2_126_3477_n1852), .S(DP_OP_424J2_126_3477_n1853) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1108 ( .A(DP_OP_424J2_126_3477_n1893), .B(
        DP_OP_424J2_126_3477_n1881), .CI(DP_OP_424J2_126_3477_n1877), .CO(
        DP_OP_424J2_126_3477_n1850), .S(DP_OP_424J2_126_3477_n1851) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1107 ( .A(DP_OP_424J2_126_3477_n1895), .B(
        DP_OP_424J2_126_3477_n1885), .CI(DP_OP_424J2_126_3477_n1869), .CO(
        DP_OP_424J2_126_3477_n1848), .S(DP_OP_424J2_126_3477_n1849) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1106 ( .A(DP_OP_424J2_126_3477_n1889), .B(
        DP_OP_424J2_126_3477_n1883), .CI(DP_OP_424J2_126_3477_n1867), .CO(
        DP_OP_424J2_126_3477_n1846), .S(DP_OP_424J2_126_3477_n1847) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1105 ( .A(DP_OP_424J2_126_3477_n1863), .B(
        DP_OP_424J2_126_3477_n1902), .CI(DP_OP_424J2_126_3477_n1900), .CO(
        DP_OP_424J2_126_3477_n1844), .S(DP_OP_424J2_126_3477_n1845) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1104 ( .A(DP_OP_424J2_126_3477_n1898), .B(
        DP_OP_424J2_126_3477_n1859), .CI(DP_OP_424J2_126_3477_n1861), .CO(
        DP_OP_424J2_126_3477_n1842), .S(DP_OP_424J2_126_3477_n1843) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1103 ( .A(DP_OP_424J2_126_3477_n1857), .B(
        DP_OP_424J2_126_3477_n1849), .CI(DP_OP_424J2_126_3477_n1851), .CO(
        DP_OP_424J2_126_3477_n1840), .S(DP_OP_424J2_126_3477_n1841) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1102 ( .A(DP_OP_424J2_126_3477_n1855), .B(
        DP_OP_424J2_126_3477_n1847), .CI(DP_OP_424J2_126_3477_n1853), .CO(
        DP_OP_424J2_126_3477_n1838), .S(DP_OP_424J2_126_3477_n1839) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1101 ( .A(DP_OP_424J2_126_3477_n1845), .B(
        DP_OP_424J2_126_3477_n1843), .CI(DP_OP_424J2_126_3477_n1841), .CO(
        DP_OP_424J2_126_3477_n1836), .S(DP_OP_424J2_126_3477_n1837) );
  HADDX1_HVT DP_OP_424J2_126_3477_U1100 ( .A0(DP_OP_424J2_126_3477_n1934), 
        .B0(DP_OP_424J2_126_3477_n1999), .C1(DP_OP_424J2_126_3477_n1834), .SO(
        DP_OP_424J2_126_3477_n1835) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1099 ( .A(DP_OP_424J2_126_3477_n2029), .B(
        DP_OP_424J2_126_3477_n1992), .CI(DP_OP_424J2_126_3477_n1985), .CO(
        DP_OP_424J2_126_3477_n1832), .S(DP_OP_424J2_126_3477_n1833) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1098 ( .A(DP_OP_424J2_126_3477_n2043), .B(
        DP_OP_424J2_126_3477_n2036), .CI(DP_OP_424J2_126_3477_n2073), .CO(
        DP_OP_424J2_126_3477_n1830), .S(DP_OP_424J2_126_3477_n1831) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1097 ( .A(DP_OP_424J2_126_3477_n2087), .B(
        DP_OP_424J2_126_3477_n2080), .CI(DP_OP_424J2_126_3477_n2117), .CO(
        DP_OP_424J2_126_3477_n1828), .S(DP_OP_424J2_126_3477_n1829) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1096 ( .A(DP_OP_424J2_126_3477_n2131), .B(
        DP_OP_424J2_126_3477_n2124), .CI(DP_OP_424J2_126_3477_n2161), .CO(
        DP_OP_424J2_126_3477_n1826), .S(DP_OP_424J2_126_3477_n1827) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1095 ( .A(DP_OP_424J2_126_3477_n2175), .B(
        DP_OP_424J2_126_3477_n2168), .CI(DP_OP_424J2_126_3477_n2205), .CO(
        DP_OP_424J2_126_3477_n1824), .S(DP_OP_424J2_126_3477_n1825) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1094 ( .A(DP_OP_424J2_126_3477_n2219), .B(
        DP_OP_424J2_126_3477_n2212), .CI(DP_OP_424J2_126_3477_n2249), .CO(
        DP_OP_424J2_126_3477_n1822), .S(DP_OP_424J2_126_3477_n1823) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1093 ( .A(DP_OP_424J2_126_3477_n2263), .B(
        DP_OP_424J2_126_3477_n2256), .CI(DP_OP_424J2_126_3477_n2293), .CO(
        DP_OP_424J2_126_3477_n1820), .S(DP_OP_424J2_126_3477_n1821) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1092 ( .A(DP_OP_424J2_126_3477_n2307), .B(
        DP_OP_424J2_126_3477_n2300), .CI(DP_OP_424J2_126_3477_n2337), .CO(
        DP_OP_424J2_126_3477_n1818), .S(DP_OP_424J2_126_3477_n1819) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1091 ( .A(DP_OP_424J2_126_3477_n2351), .B(
        DP_OP_424J2_126_3477_n2344), .CI(DP_OP_424J2_126_3477_n2381), .CO(
        DP_OP_424J2_126_3477_n1816), .S(DP_OP_424J2_126_3477_n1817) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1090 ( .A(DP_OP_424J2_126_3477_n2395), .B(
        DP_OP_424J2_126_3477_n2388), .CI(DP_OP_424J2_126_3477_n2425), .CO(
        DP_OP_424J2_126_3477_n1814), .S(DP_OP_424J2_126_3477_n1815) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1089 ( .A(DP_OP_424J2_126_3477_n2439), .B(
        DP_OP_424J2_126_3477_n2432), .CI(DP_OP_424J2_126_3477_n2469), .CO(
        DP_OP_424J2_126_3477_n1812), .S(DP_OP_424J2_126_3477_n1813) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1088 ( .A(DP_OP_424J2_126_3477_n2740), .B(
        DP_OP_424J2_126_3477_n3053), .CI(DP_OP_424J2_126_3477_n3046), .CO(
        DP_OP_424J2_126_3477_n1810), .S(DP_OP_424J2_126_3477_n1811) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1087 ( .A(DP_OP_424J2_126_3477_n2703), .B(
        DP_OP_424J2_126_3477_n2476), .CI(DP_OP_424J2_126_3477_n3039), .CO(
        DP_OP_424J2_126_3477_n1808), .S(DP_OP_424J2_126_3477_n1809) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1086 ( .A(DP_OP_424J2_126_3477_n2696), .B(
        DP_OP_424J2_126_3477_n3011), .CI(DP_OP_424J2_126_3477_n2483), .CO(
        DP_OP_424J2_126_3477_n1806), .S(DP_OP_424J2_126_3477_n1807) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1085 ( .A(DP_OP_424J2_126_3477_n2733), .B(
        DP_OP_424J2_126_3477_n2513), .CI(DP_OP_424J2_126_3477_n2520), .CO(
        DP_OP_424J2_126_3477_n1804), .S(DP_OP_424J2_126_3477_n1805) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1084 ( .A(DP_OP_424J2_126_3477_n2747), .B(
        DP_OP_424J2_126_3477_n2527), .CI(DP_OP_424J2_126_3477_n3004), .CO(
        DP_OP_424J2_126_3477_n1802), .S(DP_OP_424J2_126_3477_n1803) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1083 ( .A(DP_OP_424J2_126_3477_n2777), .B(
        DP_OP_424J2_126_3477_n2557), .CI(DP_OP_424J2_126_3477_n2997), .CO(
        DP_OP_424J2_126_3477_n1800), .S(DP_OP_424J2_126_3477_n1801) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1082 ( .A(DP_OP_424J2_126_3477_n2689), .B(
        DP_OP_424J2_126_3477_n2564), .CI(DP_OP_424J2_126_3477_n2967), .CO(
        DP_OP_424J2_126_3477_n1798), .S(DP_OP_424J2_126_3477_n1799) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1081 ( .A(DP_OP_424J2_126_3477_n2659), .B(
        DP_OP_424J2_126_3477_n2571), .CI(DP_OP_424J2_126_3477_n2960), .CO(
        DP_OP_424J2_126_3477_n1796), .S(DP_OP_424J2_126_3477_n1797) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1080 ( .A(DP_OP_424J2_126_3477_n2953), .B(
        DP_OP_424J2_126_3477_n2601), .CI(DP_OP_424J2_126_3477_n2608), .CO(
        DP_OP_424J2_126_3477_n1794), .S(DP_OP_424J2_126_3477_n1795) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1079 ( .A(DP_OP_424J2_126_3477_n2923), .B(
        DP_OP_424J2_126_3477_n2615), .CI(DP_OP_424J2_126_3477_n2645), .CO(
        DP_OP_424J2_126_3477_n1792), .S(DP_OP_424J2_126_3477_n1793) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1078 ( .A(DP_OP_424J2_126_3477_n2916), .B(
        DP_OP_424J2_126_3477_n2652), .CI(DP_OP_424J2_126_3477_n2784), .CO(
        DP_OP_424J2_126_3477_n1790), .S(DP_OP_424J2_126_3477_n1791) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1076 ( .A(DP_OP_424J2_126_3477_n2879), .B(
        DP_OP_424J2_126_3477_n2828), .CI(DP_OP_424J2_126_3477_n2835), .CO(
        DP_OP_424J2_126_3477_n1786), .S(DP_OP_424J2_126_3477_n1787) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1075 ( .A(DP_OP_424J2_126_3477_n2872), .B(
        DP_OP_424J2_126_3477_n2865), .CI(DP_OP_424J2_126_3477_n1896), .CO(
        DP_OP_424J2_126_3477_n1784), .S(DP_OP_424J2_126_3477_n1785) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1074 ( .A(DP_OP_424J2_126_3477_n1835), .B(
        DP_OP_424J2_126_3477_n1864), .CI(DP_OP_424J2_126_3477_n1866), .CO(
        DP_OP_424J2_126_3477_n1782), .S(DP_OP_424J2_126_3477_n1783) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1073 ( .A(DP_OP_424J2_126_3477_n1882), .B(
        DP_OP_424J2_126_3477_n1894), .CI(DP_OP_424J2_126_3477_n1868), .CO(
        DP_OP_424J2_126_3477_n1780), .S(DP_OP_424J2_126_3477_n1781) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1072 ( .A(DP_OP_424J2_126_3477_n1880), .B(
        DP_OP_424J2_126_3477_n1892), .CI(DP_OP_424J2_126_3477_n1870), .CO(
        DP_OP_424J2_126_3477_n1778), .S(DP_OP_424J2_126_3477_n1779) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1071 ( .A(DP_OP_424J2_126_3477_n1876), .B(
        DP_OP_424J2_126_3477_n1890), .CI(DP_OP_424J2_126_3477_n1872), .CO(
        DP_OP_424J2_126_3477_n1776), .S(DP_OP_424J2_126_3477_n1777) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1070 ( .A(DP_OP_424J2_126_3477_n1888), .B(
        DP_OP_424J2_126_3477_n1886), .CI(DP_OP_424J2_126_3477_n1884), .CO(
        DP_OP_424J2_126_3477_n1774), .S(DP_OP_424J2_126_3477_n1775) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1069 ( .A(DP_OP_424J2_126_3477_n1878), .B(
        DP_OP_424J2_126_3477_n1874), .CI(DP_OP_424J2_126_3477_n1807), .CO(
        DP_OP_424J2_126_3477_n1772), .S(DP_OP_424J2_126_3477_n1773) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1068 ( .A(DP_OP_424J2_126_3477_n1801), .B(
        DP_OP_424J2_126_3477_n1815), .CI(DP_OP_424J2_126_3477_n1819), .CO(
        DP_OP_424J2_126_3477_n1770), .S(DP_OP_424J2_126_3477_n1771) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1067 ( .A(DP_OP_424J2_126_3477_n1797), .B(
        DP_OP_424J2_126_3477_n1825), .CI(DP_OP_424J2_126_3477_n1827), .CO(
        DP_OP_424J2_126_3477_n1768), .S(DP_OP_424J2_126_3477_n1769) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1066 ( .A(DP_OP_424J2_126_3477_n1795), .B(
        DP_OP_424J2_126_3477_n1817), .CI(DP_OP_424J2_126_3477_n1831), .CO(
        DP_OP_424J2_126_3477_n1766), .S(DP_OP_424J2_126_3477_n1767) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1065 ( .A(DP_OP_424J2_126_3477_n1793), .B(
        DP_OP_424J2_126_3477_n1811), .CI(DP_OP_424J2_126_3477_n1829), .CO(
        DP_OP_424J2_126_3477_n1764), .S(DP_OP_424J2_126_3477_n1765) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1064 ( .A(DP_OP_424J2_126_3477_n1791), .B(
        DP_OP_424J2_126_3477_n1821), .CI(DP_OP_424J2_126_3477_n1809), .CO(
        DP_OP_424J2_126_3477_n1762), .S(DP_OP_424J2_126_3477_n1763) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1063 ( .A(DP_OP_424J2_126_3477_n1789), .B(
        DP_OP_424J2_126_3477_n1823), .CI(DP_OP_424J2_126_3477_n1833), .CO(
        DP_OP_424J2_126_3477_n1760), .S(DP_OP_424J2_126_3477_n1761) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1062 ( .A(DP_OP_424J2_126_3477_n1787), .B(
        DP_OP_424J2_126_3477_n1813), .CI(DP_OP_424J2_126_3477_n1799), .CO(
        DP_OP_424J2_126_3477_n1758), .S(DP_OP_424J2_126_3477_n1759) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1061 ( .A(DP_OP_424J2_126_3477_n1805), .B(
        DP_OP_424J2_126_3477_n1803), .CI(DP_OP_424J2_126_3477_n1862), .CO(
        DP_OP_424J2_126_3477_n1756), .S(DP_OP_424J2_126_3477_n1757) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1060 ( .A(DP_OP_424J2_126_3477_n1785), .B(
        DP_OP_424J2_126_3477_n1860), .CI(DP_OP_424J2_126_3477_n1858), .CO(
        DP_OP_424J2_126_3477_n1754), .S(DP_OP_424J2_126_3477_n1755) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1059 ( .A(DP_OP_424J2_126_3477_n1856), .B(
        DP_OP_424J2_126_3477_n1783), .CI(DP_OP_424J2_126_3477_n1850), .CO(
        DP_OP_424J2_126_3477_n1752), .S(DP_OP_424J2_126_3477_n1753) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1058 ( .A(DP_OP_424J2_126_3477_n1854), .B(
        DP_OP_424J2_126_3477_n1775), .CI(DP_OP_424J2_126_3477_n1781), .CO(
        DP_OP_424J2_126_3477_n1750), .S(DP_OP_424J2_126_3477_n1751) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1057 ( .A(DP_OP_424J2_126_3477_n1852), .B(
        DP_OP_424J2_126_3477_n1779), .CI(DP_OP_424J2_126_3477_n1777), .CO(
        DP_OP_424J2_126_3477_n1748), .S(DP_OP_424J2_126_3477_n1749) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1056 ( .A(DP_OP_424J2_126_3477_n1848), .B(
        DP_OP_424J2_126_3477_n1846), .CI(DP_OP_424J2_126_3477_n1773), .CO(
        DP_OP_424J2_126_3477_n1746), .S(DP_OP_424J2_126_3477_n1747) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1055 ( .A(DP_OP_424J2_126_3477_n1771), .B(
        DP_OP_424J2_126_3477_n1759), .CI(DP_OP_424J2_126_3477_n1757), .CO(
        DP_OP_424J2_126_3477_n1744), .S(DP_OP_424J2_126_3477_n1745) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1054 ( .A(DP_OP_424J2_126_3477_n1761), .B(
        DP_OP_424J2_126_3477_n1769), .CI(DP_OP_424J2_126_3477_n1767), .CO(
        DP_OP_424J2_126_3477_n1742), .S(DP_OP_424J2_126_3477_n1743) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1053 ( .A(DP_OP_424J2_126_3477_n1763), .B(
        DP_OP_424J2_126_3477_n1765), .CI(DP_OP_424J2_126_3477_n1844), .CO(
        DP_OP_424J2_126_3477_n1740), .S(DP_OP_424J2_126_3477_n1741) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1052 ( .A(DP_OP_424J2_126_3477_n1755), .B(
        DP_OP_424J2_126_3477_n1842), .CI(DP_OP_424J2_126_3477_n1753), .CO(
        DP_OP_424J2_126_3477_n1738), .S(DP_OP_424J2_126_3477_n1739) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1051 ( .A(DP_OP_424J2_126_3477_n1840), .B(
        DP_OP_424J2_126_3477_n1838), .CI(DP_OP_424J2_126_3477_n1749), .CO(
        DP_OP_424J2_126_3477_n1736), .S(DP_OP_424J2_126_3477_n1737) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1050 ( .A(DP_OP_424J2_126_3477_n1751), .B(
        DP_OP_424J2_126_3477_n1747), .CI(DP_OP_424J2_126_3477_n1745), .CO(
        DP_OP_424J2_126_3477_n1734), .S(DP_OP_424J2_126_3477_n1735) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1049 ( .A(DP_OP_424J2_126_3477_n1743), .B(
        DP_OP_424J2_126_3477_n1741), .CI(DP_OP_424J2_126_3477_n1739), .CO(
        DP_OP_424J2_126_3477_n1732), .S(DP_OP_424J2_126_3477_n1733) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1048 ( .A(DP_OP_424J2_126_3477_n1836), .B(
        DP_OP_424J2_126_3477_n1737), .CI(DP_OP_424J2_126_3477_n1735), .CO(
        DP_OP_424J2_126_3477_n1730), .S(DP_OP_424J2_126_3477_n1731) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1046 ( .A(DP_OP_424J2_126_3477_n2505), .B(
        DP_OP_424J2_126_3477_n1977), .CI(DP_OP_424J2_126_3477_n1933), .CO(
        DP_OP_424J2_126_3477_n1726), .S(DP_OP_424J2_126_3477_n1727) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1045 ( .A(DP_OP_424J2_126_3477_n2197), .B(
        DP_OP_424J2_126_3477_n2637), .CI(DP_OP_424J2_126_3477_n2417), .CO(
        DP_OP_424J2_126_3477_n1724), .S(DP_OP_424J2_126_3477_n1725) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1044 ( .A(DP_OP_424J2_126_3477_n2945), .B(
        DP_OP_424J2_126_3477_n2153), .CI(DP_OP_424J2_126_3477_n2373), .CO(
        DP_OP_424J2_126_3477_n1722), .S(DP_OP_424J2_126_3477_n1723) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1043 ( .A(DP_OP_424J2_126_3477_n2549), .B(
        DP_OP_424J2_126_3477_n2857), .CI(DP_OP_424J2_126_3477_n2461), .CO(
        DP_OP_424J2_126_3477_n1720), .S(DP_OP_424J2_126_3477_n1721) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1042 ( .A(DP_OP_424J2_126_3477_n2285), .B(
        DP_OP_424J2_126_3477_n2329), .CI(DP_OP_424J2_126_3477_n2109), .CO(
        DP_OP_424J2_126_3477_n1718), .S(DP_OP_424J2_126_3477_n1719) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1041 ( .A(DP_OP_424J2_126_3477_n2813), .B(
        DP_OP_424J2_126_3477_n2681), .CI(DP_OP_424J2_126_3477_n2725), .CO(
        DP_OP_424J2_126_3477_n1716), .S(DP_OP_424J2_126_3477_n1717) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1040 ( .A(DP_OP_424J2_126_3477_n2065), .B(
        DP_OP_424J2_126_3477_n2901), .CI(DP_OP_424J2_126_3477_n2769), .CO(
        DP_OP_424J2_126_3477_n1714), .S(DP_OP_424J2_126_3477_n1715) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1039 ( .A(DP_OP_424J2_126_3477_n2593), .B(
        DP_OP_424J2_126_3477_n2989), .CI(DP_OP_424J2_126_3477_n2241), .CO(
        DP_OP_424J2_126_3477_n1712), .S(DP_OP_424J2_126_3477_n1713) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1038 ( .A(DP_OP_424J2_126_3477_n2021), .B(
        DP_OP_424J2_126_3477_n1729), .CI(DP_OP_424J2_126_3477_n1998), .CO(
        DP_OP_424J2_126_3477_n1710), .S(DP_OP_424J2_126_3477_n1711) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1037 ( .A(DP_OP_424J2_126_3477_n2028), .B(
        DP_OP_424J2_126_3477_n1991), .CI(DP_OP_424J2_126_3477_n1984), .CO(
        DP_OP_424J2_126_3477_n1708), .S(DP_OP_424J2_126_3477_n1709) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1036 ( .A(DP_OP_424J2_126_3477_n2042), .B(
        DP_OP_424J2_126_3477_n2035), .CI(DP_OP_424J2_126_3477_n2072), .CO(
        DP_OP_424J2_126_3477_n1706), .S(DP_OP_424J2_126_3477_n1707) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1035 ( .A(DP_OP_424J2_126_3477_n2086), .B(
        DP_OP_424J2_126_3477_n2079), .CI(DP_OP_424J2_126_3477_n2116), .CO(
        DP_OP_424J2_126_3477_n1704), .S(DP_OP_424J2_126_3477_n1705) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1034 ( .A(DP_OP_424J2_126_3477_n3052), .B(
        DP_OP_424J2_126_3477_n2123), .CI(DP_OP_424J2_126_3477_n2130), .CO(
        DP_OP_424J2_126_3477_n1702), .S(DP_OP_424J2_126_3477_n1703) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1033 ( .A(DP_OP_424J2_126_3477_n2563), .B(
        DP_OP_424J2_126_3477_n3045), .CI(DP_OP_424J2_126_3477_n3038), .CO(
        DP_OP_424J2_126_3477_n1700), .S(DP_OP_424J2_126_3477_n1701) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1032 ( .A(DP_OP_424J2_126_3477_n2526), .B(
        DP_OP_424J2_126_3477_n2160), .CI(DP_OP_424J2_126_3477_n3010), .CO(
        DP_OP_424J2_126_3477_n1698), .S(DP_OP_424J2_126_3477_n1699) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1031 ( .A(DP_OP_424J2_126_3477_n2556), .B(
        DP_OP_424J2_126_3477_n2167), .CI(DP_OP_424J2_126_3477_n3003), .CO(
        DP_OP_424J2_126_3477_n1696), .S(DP_OP_424J2_126_3477_n1697) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1030 ( .A(DP_OP_424J2_126_3477_n2996), .B(
        DP_OP_424J2_126_3477_n2174), .CI(DP_OP_424J2_126_3477_n2204), .CO(
        DP_OP_424J2_126_3477_n1694), .S(DP_OP_424J2_126_3477_n1695) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1029 ( .A(DP_OP_424J2_126_3477_n2519), .B(
        DP_OP_424J2_126_3477_n2211), .CI(DP_OP_424J2_126_3477_n2218), .CO(
        DP_OP_424J2_126_3477_n1692), .S(DP_OP_424J2_126_3477_n1693) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1028 ( .A(DP_OP_424J2_126_3477_n2600), .B(
        DP_OP_424J2_126_3477_n2248), .CI(DP_OP_424J2_126_3477_n2255), .CO(
        DP_OP_424J2_126_3477_n1690), .S(DP_OP_424J2_126_3477_n1691) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1027 ( .A(DP_OP_424J2_126_3477_n2607), .B(
        DP_OP_424J2_126_3477_n2262), .CI(DP_OP_424J2_126_3477_n2292), .CO(
        DP_OP_424J2_126_3477_n1688), .S(DP_OP_424J2_126_3477_n1689) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1026 ( .A(DP_OP_424J2_126_3477_n2614), .B(
        DP_OP_424J2_126_3477_n2966), .CI(DP_OP_424J2_126_3477_n2299), .CO(
        DP_OP_424J2_126_3477_n1686), .S(DP_OP_424J2_126_3477_n1687) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1025 ( .A(DP_OP_424J2_126_3477_n2644), .B(
        DP_OP_424J2_126_3477_n2306), .CI(DP_OP_424J2_126_3477_n2959), .CO(
        DP_OP_424J2_126_3477_n1684), .S(DP_OP_424J2_126_3477_n1685) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1023 ( .A(DP_OP_424J2_126_3477_n2482), .B(
        DP_OP_424J2_126_3477_n2915), .CI(DP_OP_424J2_126_3477_n2336), .CO(
        DP_OP_424J2_126_3477_n1680), .S(DP_OP_424J2_126_3477_n1681) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1022 ( .A(DP_OP_424J2_126_3477_n2908), .B(
        DP_OP_424J2_126_3477_n2343), .CI(DP_OP_424J2_126_3477_n2878), .CO(
        DP_OP_424J2_126_3477_n1678), .S(DP_OP_424J2_126_3477_n1679) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1021 ( .A(DP_OP_424J2_126_3477_n2871), .B(
        DP_OP_424J2_126_3477_n2864), .CI(DP_OP_424J2_126_3477_n2350), .CO(
        DP_OP_424J2_126_3477_n1676), .S(DP_OP_424J2_126_3477_n1677) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1020 ( .A(DP_OP_424J2_126_3477_n2475), .B(
        DP_OP_424J2_126_3477_n2380), .CI(DP_OP_424J2_126_3477_n2834), .CO(
        DP_OP_424J2_126_3477_n1674), .S(DP_OP_424J2_126_3477_n1675) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1019 ( .A(DP_OP_424J2_126_3477_n2468), .B(
        DP_OP_424J2_126_3477_n2827), .CI(DP_OP_424J2_126_3477_n2820), .CO(
        DP_OP_424J2_126_3477_n1672), .S(DP_OP_424J2_126_3477_n1673) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1018 ( .A(DP_OP_424J2_126_3477_n2424), .B(
        DP_OP_424J2_126_3477_n2790), .CI(DP_OP_424J2_126_3477_n2783), .CO(
        DP_OP_424J2_126_3477_n1670), .S(DP_OP_424J2_126_3477_n1671) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1017 ( .A(DP_OP_424J2_126_3477_n2387), .B(
        DP_OP_424J2_126_3477_n2776), .CI(DP_OP_424J2_126_3477_n2746), .CO(
        DP_OP_424J2_126_3477_n1668), .S(DP_OP_424J2_126_3477_n1669) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1016 ( .A(DP_OP_424J2_126_3477_n2658), .B(
        DP_OP_424J2_126_3477_n2739), .CI(DP_OP_424J2_126_3477_n2394), .CO(
        DP_OP_424J2_126_3477_n1666), .S(DP_OP_424J2_126_3477_n1667) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1015 ( .A(DP_OP_424J2_126_3477_n2512), .B(
        DP_OP_424J2_126_3477_n2431), .CI(DP_OP_424J2_126_3477_n2732), .CO(
        DP_OP_424J2_126_3477_n1664), .S(DP_OP_424J2_126_3477_n1665) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1014 ( .A(DP_OP_424J2_126_3477_n2702), .B(
        DP_OP_424J2_126_3477_n2438), .CI(DP_OP_424J2_126_3477_n2651), .CO(
        DP_OP_424J2_126_3477_n1662), .S(DP_OP_424J2_126_3477_n1663) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1013 ( .A(DP_OP_424J2_126_3477_n2695), .B(
        DP_OP_424J2_126_3477_n2688), .CI(DP_OP_424J2_126_3477_n1834), .CO(
        DP_OP_424J2_126_3477_n1660), .S(DP_OP_424J2_126_3477_n1661) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1012 ( .A(DP_OP_424J2_126_3477_n1810), .B(
        DP_OP_424J2_126_3477_n1832), .CI(DP_OP_424J2_126_3477_n1786), .CO(
        DP_OP_424J2_126_3477_n1658), .S(DP_OP_424J2_126_3477_n1659) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1011 ( .A(DP_OP_424J2_126_3477_n1808), .B(
        DP_OP_424J2_126_3477_n1830), .CI(DP_OP_424J2_126_3477_n1828), .CO(
        DP_OP_424J2_126_3477_n1656), .S(DP_OP_424J2_126_3477_n1657) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1010 ( .A(DP_OP_424J2_126_3477_n1802), .B(
        DP_OP_424J2_126_3477_n1826), .CI(DP_OP_424J2_126_3477_n1824), .CO(
        DP_OP_424J2_126_3477_n1654), .S(DP_OP_424J2_126_3477_n1655) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1009 ( .A(DP_OP_424J2_126_3477_n1798), .B(
        DP_OP_424J2_126_3477_n1788), .CI(DP_OP_424J2_126_3477_n1790), .CO(
        DP_OP_424J2_126_3477_n1652), .S(DP_OP_424J2_126_3477_n1653) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1008 ( .A(DP_OP_424J2_126_3477_n1796), .B(
        DP_OP_424J2_126_3477_n1822), .CI(DP_OP_424J2_126_3477_n1792), .CO(
        DP_OP_424J2_126_3477_n1650), .S(DP_OP_424J2_126_3477_n1651) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1007 ( .A(DP_OP_424J2_126_3477_n1794), .B(
        DP_OP_424J2_126_3477_n1820), .CI(DP_OP_424J2_126_3477_n1818), .CO(
        DP_OP_424J2_126_3477_n1648), .S(DP_OP_424J2_126_3477_n1649) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1006 ( .A(DP_OP_424J2_126_3477_n1806), .B(
        DP_OP_424J2_126_3477_n1816), .CI(DP_OP_424J2_126_3477_n1800), .CO(
        DP_OP_424J2_126_3477_n1646), .S(DP_OP_424J2_126_3477_n1647) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1005 ( .A(DP_OP_424J2_126_3477_n1814), .B(
        DP_OP_424J2_126_3477_n1804), .CI(DP_OP_424J2_126_3477_n1812), .CO(
        DP_OP_424J2_126_3477_n1644), .S(DP_OP_424J2_126_3477_n1645) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1004 ( .A(DP_OP_424J2_126_3477_n1723), .B(
        DP_OP_424J2_126_3477_n1725), .CI(DP_OP_424J2_126_3477_n1711), .CO(
        DP_OP_424J2_126_3477_n1642), .S(DP_OP_424J2_126_3477_n1643) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1003 ( .A(DP_OP_424J2_126_3477_n1717), .B(
        DP_OP_424J2_126_3477_n1719), .CI(DP_OP_424J2_126_3477_n1784), .CO(
        DP_OP_424J2_126_3477_n1640), .S(DP_OP_424J2_126_3477_n1641) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1002 ( .A(DP_OP_424J2_126_3477_n1713), .B(
        DP_OP_424J2_126_3477_n1715), .CI(DP_OP_424J2_126_3477_n1721), .CO(
        DP_OP_424J2_126_3477_n1638), .S(DP_OP_424J2_126_3477_n1639) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1001 ( .A(DP_OP_424J2_126_3477_n1727), .B(
        DP_OP_424J2_126_3477_n1677), .CI(DP_OP_424J2_126_3477_n1675), .CO(
        DP_OP_424J2_126_3477_n1636), .S(DP_OP_424J2_126_3477_n1637) );
  FADDX1_HVT DP_OP_424J2_126_3477_U1000 ( .A(DP_OP_424J2_126_3477_n1679), .B(
        DP_OP_424J2_126_3477_n1695), .CI(DP_OP_424J2_126_3477_n1703), .CO(
        DP_OP_424J2_126_3477_n1634), .S(DP_OP_424J2_126_3477_n1635) );
  FADDX1_HVT DP_OP_424J2_126_3477_U999 ( .A(DP_OP_424J2_126_3477_n1671), .B(
        DP_OP_424J2_126_3477_n1691), .CI(DP_OP_424J2_126_3477_n1689), .CO(
        DP_OP_424J2_126_3477_n1632), .S(DP_OP_424J2_126_3477_n1633) );
  FADDX1_HVT DP_OP_424J2_126_3477_U998 ( .A(DP_OP_424J2_126_3477_n1669), .B(
        DP_OP_424J2_126_3477_n1705), .CI(DP_OP_424J2_126_3477_n1693), .CO(
        DP_OP_424J2_126_3477_n1630), .S(DP_OP_424J2_126_3477_n1631) );
  FADDX1_HVT DP_OP_424J2_126_3477_U997 ( .A(DP_OP_424J2_126_3477_n1667), .B(
        DP_OP_424J2_126_3477_n1699), .CI(DP_OP_424J2_126_3477_n1701), .CO(
        DP_OP_424J2_126_3477_n1628), .S(DP_OP_424J2_126_3477_n1629) );
  FADDX1_HVT DP_OP_424J2_126_3477_U996 ( .A(DP_OP_424J2_126_3477_n1665), .B(
        DP_OP_424J2_126_3477_n1697), .CI(DP_OP_424J2_126_3477_n1709), .CO(
        DP_OP_424J2_126_3477_n1626), .S(DP_OP_424J2_126_3477_n1627) );
  FADDX1_HVT DP_OP_424J2_126_3477_U995 ( .A(DP_OP_424J2_126_3477_n1687), .B(
        DP_OP_424J2_126_3477_n1707), .CI(DP_OP_424J2_126_3477_n1663), .CO(
        DP_OP_424J2_126_3477_n1624), .S(DP_OP_424J2_126_3477_n1625) );
  FADDX1_HVT DP_OP_424J2_126_3477_U994 ( .A(DP_OP_424J2_126_3477_n1673), .B(
        DP_OP_424J2_126_3477_n1683), .CI(DP_OP_424J2_126_3477_n1685), .CO(
        DP_OP_424J2_126_3477_n1622), .S(DP_OP_424J2_126_3477_n1623) );
  FADDX1_HVT DP_OP_424J2_126_3477_U993 ( .A(DP_OP_424J2_126_3477_n1681), .B(
        DP_OP_424J2_126_3477_n1661), .CI(DP_OP_424J2_126_3477_n1782), .CO(
        DP_OP_424J2_126_3477_n1620), .S(DP_OP_424J2_126_3477_n1621) );
  FADDX1_HVT DP_OP_424J2_126_3477_U992 ( .A(DP_OP_424J2_126_3477_n1780), .B(
        DP_OP_424J2_126_3477_n1778), .CI(DP_OP_424J2_126_3477_n1776), .CO(
        DP_OP_424J2_126_3477_n1618), .S(DP_OP_424J2_126_3477_n1619) );
  FADDX1_HVT DP_OP_424J2_126_3477_U991 ( .A(DP_OP_424J2_126_3477_n1774), .B(
        DP_OP_424J2_126_3477_n1772), .CI(DP_OP_424J2_126_3477_n1760), .CO(
        DP_OP_424J2_126_3477_n1616), .S(DP_OP_424J2_126_3477_n1617) );
  FADDX1_HVT DP_OP_424J2_126_3477_U990 ( .A(DP_OP_424J2_126_3477_n1758), .B(
        DP_OP_424J2_126_3477_n1659), .CI(DP_OP_424J2_126_3477_n1756), .CO(
        DP_OP_424J2_126_3477_n1614), .S(DP_OP_424J2_126_3477_n1615) );
  FADDX1_HVT DP_OP_424J2_126_3477_U989 ( .A(DP_OP_424J2_126_3477_n1770), .B(
        DP_OP_424J2_126_3477_n1649), .CI(DP_OP_424J2_126_3477_n1657), .CO(
        DP_OP_424J2_126_3477_n1612), .S(DP_OP_424J2_126_3477_n1613) );
  FADDX1_HVT DP_OP_424J2_126_3477_U988 ( .A(DP_OP_424J2_126_3477_n1768), .B(
        DP_OP_424J2_126_3477_n1647), .CI(DP_OP_424J2_126_3477_n1651), .CO(
        DP_OP_424J2_126_3477_n1610), .S(DP_OP_424J2_126_3477_n1611) );
  FADDX1_HVT DP_OP_424J2_126_3477_U987 ( .A(DP_OP_424J2_126_3477_n1764), .B(
        DP_OP_424J2_126_3477_n1655), .CI(DP_OP_424J2_126_3477_n1653), .CO(
        DP_OP_424J2_126_3477_n1608), .S(DP_OP_424J2_126_3477_n1609) );
  FADDX1_HVT DP_OP_424J2_126_3477_U986 ( .A(DP_OP_424J2_126_3477_n1762), .B(
        DP_OP_424J2_126_3477_n1645), .CI(DP_OP_424J2_126_3477_n1766), .CO(
        DP_OP_424J2_126_3477_n1606), .S(DP_OP_424J2_126_3477_n1607) );
  FADDX1_HVT DP_OP_424J2_126_3477_U985 ( .A(DP_OP_424J2_126_3477_n1641), .B(
        DP_OP_424J2_126_3477_n1643), .CI(DP_OP_424J2_126_3477_n1637), .CO(
        DP_OP_424J2_126_3477_n1604), .S(DP_OP_424J2_126_3477_n1605) );
  FADDX1_HVT DP_OP_424J2_126_3477_U984 ( .A(DP_OP_424J2_126_3477_n1639), .B(
        DP_OP_424J2_126_3477_n1625), .CI(DP_OP_424J2_126_3477_n1627), .CO(
        DP_OP_424J2_126_3477_n1602), .S(DP_OP_424J2_126_3477_n1603) );
  FADDX1_HVT DP_OP_424J2_126_3477_U983 ( .A(DP_OP_424J2_126_3477_n1633), .B(
        DP_OP_424J2_126_3477_n1631), .CI(DP_OP_424J2_126_3477_n1754), .CO(
        DP_OP_424J2_126_3477_n1600), .S(DP_OP_424J2_126_3477_n1601) );
  FADDX1_HVT DP_OP_424J2_126_3477_U982 ( .A(DP_OP_424J2_126_3477_n1629), .B(
        DP_OP_424J2_126_3477_n1623), .CI(DP_OP_424J2_126_3477_n1635), .CO(
        DP_OP_424J2_126_3477_n1598), .S(DP_OP_424J2_126_3477_n1599) );
  FADDX1_HVT DP_OP_424J2_126_3477_U981 ( .A(DP_OP_424J2_126_3477_n1621), .B(
        DP_OP_424J2_126_3477_n1752), .CI(DP_OP_424J2_126_3477_n1748), .CO(
        DP_OP_424J2_126_3477_n1596), .S(DP_OP_424J2_126_3477_n1597) );
  FADDX1_HVT DP_OP_424J2_126_3477_U980 ( .A(DP_OP_424J2_126_3477_n1750), .B(
        DP_OP_424J2_126_3477_n1619), .CI(DP_OP_424J2_126_3477_n1746), .CO(
        DP_OP_424J2_126_3477_n1594), .S(DP_OP_424J2_126_3477_n1595) );
  FADDX1_HVT DP_OP_424J2_126_3477_U979 ( .A(DP_OP_424J2_126_3477_n1617), .B(
        DP_OP_424J2_126_3477_n1607), .CI(DP_OP_424J2_126_3477_n1609), .CO(
        DP_OP_424J2_126_3477_n1592), .S(DP_OP_424J2_126_3477_n1593) );
  FADDX1_HVT DP_OP_424J2_126_3477_U978 ( .A(DP_OP_424J2_126_3477_n1611), .B(
        DP_OP_424J2_126_3477_n1744), .CI(DP_OP_424J2_126_3477_n1742), .CO(
        DP_OP_424J2_126_3477_n1590), .S(DP_OP_424J2_126_3477_n1591) );
  FADDX1_HVT DP_OP_424J2_126_3477_U977 ( .A(DP_OP_424J2_126_3477_n1615), .B(
        DP_OP_424J2_126_3477_n1613), .CI(DP_OP_424J2_126_3477_n1605), .CO(
        DP_OP_424J2_126_3477_n1588), .S(DP_OP_424J2_126_3477_n1589) );
  FADDX1_HVT DP_OP_424J2_126_3477_U976 ( .A(DP_OP_424J2_126_3477_n1740), .B(
        DP_OP_424J2_126_3477_n1603), .CI(DP_OP_424J2_126_3477_n1599), .CO(
        DP_OP_424J2_126_3477_n1586), .S(DP_OP_424J2_126_3477_n1587) );
  FADDX1_HVT DP_OP_424J2_126_3477_U975 ( .A(DP_OP_424J2_126_3477_n1601), .B(
        DP_OP_424J2_126_3477_n1738), .CI(DP_OP_424J2_126_3477_n1597), .CO(
        DP_OP_424J2_126_3477_n1584), .S(DP_OP_424J2_126_3477_n1585) );
  FADDX1_HVT DP_OP_424J2_126_3477_U974 ( .A(DP_OP_424J2_126_3477_n1736), .B(
        DP_OP_424J2_126_3477_n1595), .CI(DP_OP_424J2_126_3477_n1734), .CO(
        DP_OP_424J2_126_3477_n1582), .S(DP_OP_424J2_126_3477_n1583) );
  FADDX1_HVT DP_OP_424J2_126_3477_U973 ( .A(DP_OP_424J2_126_3477_n1593), .B(
        DP_OP_424J2_126_3477_n1591), .CI(DP_OP_424J2_126_3477_n1589), .CO(
        DP_OP_424J2_126_3477_n1580), .S(DP_OP_424J2_126_3477_n1581) );
  FADDX1_HVT DP_OP_424J2_126_3477_U972 ( .A(DP_OP_424J2_126_3477_n1587), .B(
        DP_OP_424J2_126_3477_n1732), .CI(DP_OP_424J2_126_3477_n1585), .CO(
        DP_OP_424J2_126_3477_n1578), .S(DP_OP_424J2_126_3477_n1579) );
  FADDX1_HVT DP_OP_424J2_126_3477_U971 ( .A(DP_OP_424J2_126_3477_n1730), .B(
        DP_OP_424J2_126_3477_n1583), .CI(DP_OP_424J2_126_3477_n1581), .CO(
        DP_OP_424J2_126_3477_n1576), .S(DP_OP_424J2_126_3477_n1577) );
  FADDX1_HVT DP_OP_424J2_126_3477_U970 ( .A(DP_OP_424J2_126_3477_n1728), .B(
        DP_OP_424J2_126_3477_n1976), .CI(DP_OP_424J2_126_3477_n1932), .CO(
        DP_OP_424J2_126_3477_n1574), .S(DP_OP_424J2_126_3477_n1575) );
  FADDX1_HVT DP_OP_424J2_126_3477_U969 ( .A(DP_OP_424J2_126_3477_n3031), .B(
        DP_OP_424J2_126_3477_n2548), .CI(DP_OP_424J2_126_3477_n2416), .CO(
        DP_OP_424J2_126_3477_n1572), .S(DP_OP_424J2_126_3477_n1573) );
  FADDX1_HVT DP_OP_424J2_126_3477_U968 ( .A(DP_OP_424J2_126_3477_n2944), .B(
        DP_OP_424J2_126_3477_n2680), .CI(DP_OP_424J2_126_3477_n2328), .CO(
        DP_OP_424J2_126_3477_n1570), .S(DP_OP_424J2_126_3477_n1571) );
  FADDX1_HVT DP_OP_424J2_126_3477_U967 ( .A(DP_OP_424J2_126_3477_n2108), .B(
        DP_OP_424J2_126_3477_n2636), .CI(DP_OP_424J2_126_3477_n2856), .CO(
        DP_OP_424J2_126_3477_n1568), .S(DP_OP_424J2_126_3477_n1569) );
  FADDX1_HVT DP_OP_424J2_126_3477_U966 ( .A(DP_OP_424J2_126_3477_n2196), .B(
        DP_OP_424J2_126_3477_n2372), .CI(DP_OP_424J2_126_3477_n2460), .CO(
        DP_OP_424J2_126_3477_n1566), .S(DP_OP_424J2_126_3477_n1567) );
  FADDX1_HVT DP_OP_424J2_126_3477_U965 ( .A(DP_OP_424J2_126_3477_n2812), .B(
        DP_OP_424J2_126_3477_n2284), .CI(DP_OP_424J2_126_3477_n2900), .CO(
        DP_OP_424J2_126_3477_n1564), .S(DP_OP_424J2_126_3477_n1565) );
  FADDX1_HVT DP_OP_424J2_126_3477_U964 ( .A(DP_OP_424J2_126_3477_n2152), .B(
        DP_OP_424J2_126_3477_n2504), .CI(DP_OP_424J2_126_3477_n2592), .CO(
        DP_OP_424J2_126_3477_n1562), .S(DP_OP_424J2_126_3477_n1563) );
  FADDX1_HVT DP_OP_424J2_126_3477_U963 ( .A(DP_OP_424J2_126_3477_n2988), .B(
        DP_OP_424J2_126_3477_n2724), .CI(DP_OP_424J2_126_3477_n2768), .CO(
        DP_OP_424J2_126_3477_n1560), .S(DP_OP_424J2_126_3477_n1561) );
  FADDX1_HVT DP_OP_424J2_126_3477_U962 ( .A(DP_OP_424J2_126_3477_n2064), .B(
        DP_OP_424J2_126_3477_n2240), .CI(DP_OP_424J2_126_3477_n2020), .CO(
        DP_OP_424J2_126_3477_n1558), .S(DP_OP_424J2_126_3477_n1559) );
  FADDX1_HVT DP_OP_424J2_126_3477_U961 ( .A(DP_OP_424J2_126_3477_n2555), .B(
        DP_OP_424J2_126_3477_n1990), .CI(DP_OP_424J2_126_3477_n1983), .CO(
        DP_OP_424J2_126_3477_n1556), .S(DP_OP_424J2_126_3477_n1557) );
  FADDX1_HVT DP_OP_424J2_126_3477_U960 ( .A(DP_OP_424J2_126_3477_n3051), .B(
        DP_OP_424J2_126_3477_n1997), .CI(DP_OP_424J2_126_3477_n2027), .CO(
        DP_OP_424J2_126_3477_n1554), .S(DP_OP_424J2_126_3477_n1555) );
  FADDX1_HVT DP_OP_424J2_126_3477_U959 ( .A(DP_OP_424J2_126_3477_n2437), .B(
        DP_OP_424J2_126_3477_n3044), .CI(DP_OP_424J2_126_3477_n2034), .CO(
        DP_OP_424J2_126_3477_n1552), .S(DP_OP_424J2_126_3477_n1553) );
  FADDX1_HVT DP_OP_424J2_126_3477_U958 ( .A(DP_OP_424J2_126_3477_n2430), .B(
        DP_OP_424J2_126_3477_n3037), .CI(DP_OP_424J2_126_3477_n2041), .CO(
        DP_OP_424J2_126_3477_n1550), .S(DP_OP_424J2_126_3477_n1551) );
  FADDX1_HVT DP_OP_424J2_126_3477_U957 ( .A(DP_OP_424J2_126_3477_n3009), .B(
        DP_OP_424J2_126_3477_n2071), .CI(DP_OP_424J2_126_3477_n2078), .CO(
        DP_OP_424J2_126_3477_n1548), .S(DP_OP_424J2_126_3477_n1549) );
  FADDX1_HVT DP_OP_424J2_126_3477_U956 ( .A(DP_OP_424J2_126_3477_n2467), .B(
        DP_OP_424J2_126_3477_n3002), .CI(DP_OP_424J2_126_3477_n2995), .CO(
        DP_OP_424J2_126_3477_n1546), .S(DP_OP_424J2_126_3477_n1547) );
  FADDX1_HVT DP_OP_424J2_126_3477_U955 ( .A(DP_OP_424J2_126_3477_n2393), .B(
        DP_OP_424J2_126_3477_n2965), .CI(DP_OP_424J2_126_3477_n2958), .CO(
        DP_OP_424J2_126_3477_n1544), .S(DP_OP_424J2_126_3477_n1545) );
  FADDX1_HVT DP_OP_424J2_126_3477_U954 ( .A(DP_OP_424J2_126_3477_n2386), .B(
        DP_OP_424J2_126_3477_n2951), .CI(DP_OP_424J2_126_3477_n2085), .CO(
        DP_OP_424J2_126_3477_n1542), .S(DP_OP_424J2_126_3477_n1543) );
  FADDX1_HVT DP_OP_424J2_126_3477_U953 ( .A(DP_OP_424J2_126_3477_n2379), .B(
        DP_OP_424J2_126_3477_n2921), .CI(DP_OP_424J2_126_3477_n2914), .CO(
        DP_OP_424J2_126_3477_n1540), .S(DP_OP_424J2_126_3477_n1541) );
  FADDX1_HVT DP_OP_424J2_126_3477_U952 ( .A(DP_OP_424J2_126_3477_n2349), .B(
        DP_OP_424J2_126_3477_n2907), .CI(DP_OP_424J2_126_3477_n2115), .CO(
        DP_OP_424J2_126_3477_n1538), .S(DP_OP_424J2_126_3477_n1539) );
  FADDX1_HVT DP_OP_424J2_126_3477_U951 ( .A(DP_OP_424J2_126_3477_n2342), .B(
        DP_OP_424J2_126_3477_n2122), .CI(DP_OP_424J2_126_3477_n2129), .CO(
        DP_OP_424J2_126_3477_n1536), .S(DP_OP_424J2_126_3477_n1537) );
  FADDX1_HVT DP_OP_424J2_126_3477_U950 ( .A(DP_OP_424J2_126_3477_n2423), .B(
        DP_OP_424J2_126_3477_n2159), .CI(DP_OP_424J2_126_3477_n2877), .CO(
        DP_OP_424J2_126_3477_n1534), .S(DP_OP_424J2_126_3477_n1535) );
  FADDX1_HVT DP_OP_424J2_126_3477_U949 ( .A(DP_OP_424J2_126_3477_n2474), .B(
        DP_OP_424J2_126_3477_n2870), .CI(DP_OP_424J2_126_3477_n2863), .CO(
        DP_OP_424J2_126_3477_n1532), .S(DP_OP_424J2_126_3477_n1533) );
  FADDX1_HVT DP_OP_424J2_126_3477_U948 ( .A(DP_OP_424J2_126_3477_n2833), .B(
        DP_OP_424J2_126_3477_n2166), .CI(DP_OP_424J2_126_3477_n2173), .CO(
        DP_OP_424J2_126_3477_n1530), .S(DP_OP_424J2_126_3477_n1531) );
  FADDX1_HVT DP_OP_424J2_126_3477_U947 ( .A(DP_OP_424J2_126_3477_n2606), .B(
        DP_OP_424J2_126_3477_n2203), .CI(DP_OP_424J2_126_3477_n2210), .CO(
        DP_OP_424J2_126_3477_n1528), .S(DP_OP_424J2_126_3477_n1529) );
  FADDX1_HVT DP_OP_424J2_126_3477_U946 ( .A(DP_OP_424J2_126_3477_n2826), .B(
        DP_OP_424J2_126_3477_n2217), .CI(DP_OP_424J2_126_3477_n2247), .CO(
        DP_OP_424J2_126_3477_n1526), .S(DP_OP_424J2_126_3477_n1527) );
  FADDX1_HVT DP_OP_424J2_126_3477_U945 ( .A(DP_OP_424J2_126_3477_n2819), .B(
        DP_OP_424J2_126_3477_n2254), .CI(DP_OP_424J2_126_3477_n2261), .CO(
        DP_OP_424J2_126_3477_n1524), .S(DP_OP_424J2_126_3477_n1525) );
  FADDX1_HVT DP_OP_424J2_126_3477_U944 ( .A(DP_OP_424J2_126_3477_n2789), .B(
        DP_OP_424J2_126_3477_n2291), .CI(DP_OP_424J2_126_3477_n2298), .CO(
        DP_OP_424J2_126_3477_n1522), .S(DP_OP_424J2_126_3477_n1523) );
  FADDX1_HVT DP_OP_424J2_126_3477_U943 ( .A(DP_OP_424J2_126_3477_n2782), .B(
        DP_OP_424J2_126_3477_n2305), .CI(DP_OP_424J2_126_3477_n2335), .CO(
        DP_OP_424J2_126_3477_n1520), .S(DP_OP_424J2_126_3477_n1521) );
  FADDX1_HVT DP_OP_424J2_126_3477_U942 ( .A(DP_OP_424J2_126_3477_n2775), .B(
        DP_OP_424J2_126_3477_n2481), .CI(DP_OP_424J2_126_3477_n2511), .CO(
        DP_OP_424J2_126_3477_n1518), .S(DP_OP_424J2_126_3477_n1519) );
  FADDX1_HVT DP_OP_424J2_126_3477_U941 ( .A(DP_OP_424J2_126_3477_n2745), .B(
        DP_OP_424J2_126_3477_n2518), .CI(DP_OP_424J2_126_3477_n2738), .CO(
        DP_OP_424J2_126_3477_n1516), .S(DP_OP_424J2_126_3477_n1517) );
  FADDX1_HVT DP_OP_424J2_126_3477_U940 ( .A(DP_OP_424J2_126_3477_n2643), .B(
        DP_OP_424J2_126_3477_n2525), .CI(DP_OP_424J2_126_3477_n2562), .CO(
        DP_OP_424J2_126_3477_n1514), .S(DP_OP_424J2_126_3477_n1515) );
  FADDX1_HVT DP_OP_424J2_126_3477_U939 ( .A(DP_OP_424J2_126_3477_n2613), .B(
        DP_OP_424J2_126_3477_n2569), .CI(DP_OP_424J2_126_3477_n2731), .CO(
        DP_OP_424J2_126_3477_n1512), .S(DP_OP_424J2_126_3477_n1513) );
  FADDX1_HVT DP_OP_424J2_126_3477_U938 ( .A(DP_OP_424J2_126_3477_n2687), .B(
        DP_OP_424J2_126_3477_n2599), .CI(DP_OP_424J2_126_3477_n2701), .CO(
        DP_OP_424J2_126_3477_n1510), .S(DP_OP_424J2_126_3477_n1511) );
  FADDX1_HVT DP_OP_424J2_126_3477_U937 ( .A(DP_OP_424J2_126_3477_n2650), .B(
        DP_OP_424J2_126_3477_n2657), .CI(DP_OP_424J2_126_3477_n2694), .CO(
        DP_OP_424J2_126_3477_n1508), .S(DP_OP_424J2_126_3477_n1509) );
  FADDX1_HVT DP_OP_424J2_126_3477_U936 ( .A(DP_OP_424J2_126_3477_n1716), .B(
        DP_OP_424J2_126_3477_n1712), .CI(DP_OP_424J2_126_3477_n1710), .CO(
        DP_OP_424J2_126_3477_n1506), .S(DP_OP_424J2_126_3477_n1507) );
  FADDX1_HVT DP_OP_424J2_126_3477_U935 ( .A(DP_OP_424J2_126_3477_n1714), .B(
        DP_OP_424J2_126_3477_n1718), .CI(DP_OP_424J2_126_3477_n1720), .CO(
        DP_OP_424J2_126_3477_n1504), .S(DP_OP_424J2_126_3477_n1505) );
  FADDX1_HVT DP_OP_424J2_126_3477_U934 ( .A(DP_OP_424J2_126_3477_n1722), .B(
        DP_OP_424J2_126_3477_n1724), .CI(DP_OP_424J2_126_3477_n1726), .CO(
        DP_OP_424J2_126_3477_n1502), .S(DP_OP_424J2_126_3477_n1503) );
  FADDX1_HVT DP_OP_424J2_126_3477_U933 ( .A(DP_OP_424J2_126_3477_n1686), .B(
        DP_OP_424J2_126_3477_n1708), .CI(DP_OP_424J2_126_3477_n1706), .CO(
        DP_OP_424J2_126_3477_n1500), .S(DP_OP_424J2_126_3477_n1501) );
  FADDX1_HVT DP_OP_424J2_126_3477_U932 ( .A(DP_OP_424J2_126_3477_n1682), .B(
        DP_OP_424J2_126_3477_n1704), .CI(DP_OP_424J2_126_3477_n1702), .CO(
        DP_OP_424J2_126_3477_n1498), .S(DP_OP_424J2_126_3477_n1499) );
  FADDX1_HVT DP_OP_424J2_126_3477_U931 ( .A(DP_OP_424J2_126_3477_n1676), .B(
        DP_OP_424J2_126_3477_n1700), .CI(DP_OP_424J2_126_3477_n1698), .CO(
        DP_OP_424J2_126_3477_n1496), .S(DP_OP_424J2_126_3477_n1497) );
  FADDX1_HVT DP_OP_424J2_126_3477_U930 ( .A(DP_OP_424J2_126_3477_n1672), .B(
        DP_OP_424J2_126_3477_n1696), .CI(DP_OP_424J2_126_3477_n1662), .CO(
        DP_OP_424J2_126_3477_n1494), .S(DP_OP_424J2_126_3477_n1495) );
  FADDX1_HVT DP_OP_424J2_126_3477_U929 ( .A(DP_OP_424J2_126_3477_n1668), .B(
        DP_OP_424J2_126_3477_n1694), .CI(DP_OP_424J2_126_3477_n1692), .CO(
        DP_OP_424J2_126_3477_n1492), .S(DP_OP_424J2_126_3477_n1493) );
  FADDX1_HVT DP_OP_424J2_126_3477_U928 ( .A(DP_OP_424J2_126_3477_n1678), .B(
        DP_OP_424J2_126_3477_n1690), .CI(DP_OP_424J2_126_3477_n1688), .CO(
        DP_OP_424J2_126_3477_n1490), .S(DP_OP_424J2_126_3477_n1491) );
  FADDX1_HVT DP_OP_424J2_126_3477_U927 ( .A(DP_OP_424J2_126_3477_n1670), .B(
        DP_OP_424J2_126_3477_n1684), .CI(DP_OP_424J2_126_3477_n1680), .CO(
        DP_OP_424J2_126_3477_n1488), .S(DP_OP_424J2_126_3477_n1489) );
  FADDX1_HVT DP_OP_424J2_126_3477_U926 ( .A(DP_OP_424J2_126_3477_n1666), .B(
        DP_OP_424J2_126_3477_n1674), .CI(DP_OP_424J2_126_3477_n1664), .CO(
        DP_OP_424J2_126_3477_n1486), .S(DP_OP_424J2_126_3477_n1487) );
  FADDX1_HVT DP_OP_424J2_126_3477_U925 ( .A(DP_OP_424J2_126_3477_n1575), .B(
        DP_OP_424J2_126_3477_n1559), .CI(DP_OP_424J2_126_3477_n1660), .CO(
        DP_OP_424J2_126_3477_n1484), .S(DP_OP_424J2_126_3477_n1485) );
  FADDX1_HVT DP_OP_424J2_126_3477_U924 ( .A(DP_OP_424J2_126_3477_n1573), .B(
        DP_OP_424J2_126_3477_n1561), .CI(DP_OP_424J2_126_3477_n1563), .CO(
        DP_OP_424J2_126_3477_n1482), .S(DP_OP_424J2_126_3477_n1483) );
  FADDX1_HVT DP_OP_424J2_126_3477_U923 ( .A(DP_OP_424J2_126_3477_n1569), .B(
        DP_OP_424J2_126_3477_n1567), .CI(DP_OP_424J2_126_3477_n1571), .CO(
        DP_OP_424J2_126_3477_n1480), .S(DP_OP_424J2_126_3477_n1481) );
  FADDX1_HVT DP_OP_424J2_126_3477_U922 ( .A(DP_OP_424J2_126_3477_n1565), .B(
        DP_OP_424J2_126_3477_n1545), .CI(DP_OP_424J2_126_3477_n1549), .CO(
        DP_OP_424J2_126_3477_n1478), .S(DP_OP_424J2_126_3477_n1479) );
  FADDX1_HVT DP_OP_424J2_126_3477_U921 ( .A(DP_OP_424J2_126_3477_n1547), .B(
        DP_OP_424J2_126_3477_n1555), .CI(DP_OP_424J2_126_3477_n1553), .CO(
        DP_OP_424J2_126_3477_n1476), .S(DP_OP_424J2_126_3477_n1477) );
  FADDX1_HVT DP_OP_424J2_126_3477_U920 ( .A(DP_OP_424J2_126_3477_n1557), .B(
        DP_OP_424J2_126_3477_n1535), .CI(DP_OP_424J2_126_3477_n1529), .CO(
        DP_OP_424J2_126_3477_n1474), .S(DP_OP_424J2_126_3477_n1475) );
  FADDX1_HVT DP_OP_424J2_126_3477_U919 ( .A(DP_OP_424J2_126_3477_n1537), .B(
        DP_OP_424J2_126_3477_n1533), .CI(DP_OP_424J2_126_3477_n1527), .CO(
        DP_OP_424J2_126_3477_n1472), .S(DP_OP_424J2_126_3477_n1473) );
  FADDX1_HVT DP_OP_424J2_126_3477_U918 ( .A(DP_OP_424J2_126_3477_n1539), .B(
        DP_OP_424J2_126_3477_n1513), .CI(DP_OP_424J2_126_3477_n1511), .CO(
        DP_OP_424J2_126_3477_n1470), .S(DP_OP_424J2_126_3477_n1471) );
  FADDX1_HVT DP_OP_424J2_126_3477_U917 ( .A(DP_OP_424J2_126_3477_n1525), .B(
        DP_OP_424J2_126_3477_n1521), .CI(DP_OP_424J2_126_3477_n1523), .CO(
        DP_OP_424J2_126_3477_n1468), .S(DP_OP_424J2_126_3477_n1469) );
  FADDX1_HVT DP_OP_424J2_126_3477_U915 ( .A(DP_OP_424J2_126_3477_n1519), .B(
        DP_OP_424J2_126_3477_n1543), .CI(DP_OP_424J2_126_3477_n1551), .CO(
        DP_OP_424J2_126_3477_n1464), .S(DP_OP_424J2_126_3477_n1465) );
  FADDX1_HVT DP_OP_424J2_126_3477_U914 ( .A(DP_OP_424J2_126_3477_n1515), .B(
        DP_OP_424J2_126_3477_n1541), .CI(DP_OP_424J2_126_3477_n1658), .CO(
        DP_OP_424J2_126_3477_n1462), .S(DP_OP_424J2_126_3477_n1463) );
  FADDX1_HVT DP_OP_424J2_126_3477_U913 ( .A(DP_OP_424J2_126_3477_n1652), .B(
        DP_OP_424J2_126_3477_n1654), .CI(DP_OP_424J2_126_3477_n1656), .CO(
        DP_OP_424J2_126_3477_n1460), .S(DP_OP_424J2_126_3477_n1461) );
  FADDX1_HVT DP_OP_424J2_126_3477_U912 ( .A(DP_OP_424J2_126_3477_n1644), .B(
        DP_OP_424J2_126_3477_n1650), .CI(DP_OP_424J2_126_3477_n1646), .CO(
        DP_OP_424J2_126_3477_n1458), .S(DP_OP_424J2_126_3477_n1459) );
  FADDX1_HVT DP_OP_424J2_126_3477_U911 ( .A(DP_OP_424J2_126_3477_n1648), .B(
        DP_OP_424J2_126_3477_n1642), .CI(DP_OP_424J2_126_3477_n1503), .CO(
        DP_OP_424J2_126_3477_n1456), .S(DP_OP_424J2_126_3477_n1457) );
  FADDX1_HVT DP_OP_424J2_126_3477_U910 ( .A(DP_OP_424J2_126_3477_n1505), .B(
        DP_OP_424J2_126_3477_n1640), .CI(DP_OP_424J2_126_3477_n1636), .CO(
        DP_OP_424J2_126_3477_n1454), .S(DP_OP_424J2_126_3477_n1455) );
  FADDX1_HVT DP_OP_424J2_126_3477_U909 ( .A(DP_OP_424J2_126_3477_n1507), .B(
        DP_OP_424J2_126_3477_n1638), .CI(DP_OP_424J2_126_3477_n1634), .CO(
        DP_OP_424J2_126_3477_n1452), .S(DP_OP_424J2_126_3477_n1453) );
  FADDX1_HVT DP_OP_424J2_126_3477_U908 ( .A(DP_OP_424J2_126_3477_n1624), .B(
        DP_OP_424J2_126_3477_n1487), .CI(DP_OP_424J2_126_3477_n1499), .CO(
        DP_OP_424J2_126_3477_n1450), .S(DP_OP_424J2_126_3477_n1451) );
  FADDX1_HVT DP_OP_424J2_126_3477_U907 ( .A(DP_OP_424J2_126_3477_n1632), .B(
        DP_OP_424J2_126_3477_n1501), .CI(DP_OP_424J2_126_3477_n1497), .CO(
        DP_OP_424J2_126_3477_n1448), .S(DP_OP_424J2_126_3477_n1449) );
  FADDX1_HVT DP_OP_424J2_126_3477_U906 ( .A(DP_OP_424J2_126_3477_n1630), .B(
        DP_OP_424J2_126_3477_n1489), .CI(DP_OP_424J2_126_3477_n1491), .CO(
        DP_OP_424J2_126_3477_n1446), .S(DP_OP_424J2_126_3477_n1447) );
  FADDX1_HVT DP_OP_424J2_126_3477_U905 ( .A(DP_OP_424J2_126_3477_n1628), .B(
        DP_OP_424J2_126_3477_n1495), .CI(DP_OP_424J2_126_3477_n1493), .CO(
        DP_OP_424J2_126_3477_n1444), .S(DP_OP_424J2_126_3477_n1445) );
  FADDX1_HVT DP_OP_424J2_126_3477_U904 ( .A(DP_OP_424J2_126_3477_n1626), .B(
        DP_OP_424J2_126_3477_n1622), .CI(DP_OP_424J2_126_3477_n1483), .CO(
        DP_OP_424J2_126_3477_n1442), .S(DP_OP_424J2_126_3477_n1443) );
  FADDX1_HVT DP_OP_424J2_126_3477_U903 ( .A(DP_OP_424J2_126_3477_n1485), .B(
        DP_OP_424J2_126_3477_n1481), .CI(DP_OP_424J2_126_3477_n1479), .CO(
        DP_OP_424J2_126_3477_n1440), .S(DP_OP_424J2_126_3477_n1441) );
  FADDX1_HVT DP_OP_424J2_126_3477_U902 ( .A(DP_OP_424J2_126_3477_n1620), .B(
        DP_OP_424J2_126_3477_n1471), .CI(DP_OP_424J2_126_3477_n1469), .CO(
        DP_OP_424J2_126_3477_n1438), .S(DP_OP_424J2_126_3477_n1439) );
  FADDX1_HVT DP_OP_424J2_126_3477_U901 ( .A(DP_OP_424J2_126_3477_n1475), .B(
        DP_OP_424J2_126_3477_n1465), .CI(DP_OP_424J2_126_3477_n1467), .CO(
        DP_OP_424J2_126_3477_n1436), .S(DP_OP_424J2_126_3477_n1437) );
  FADDX1_HVT DP_OP_424J2_126_3477_U900 ( .A(DP_OP_424J2_126_3477_n1473), .B(
        DP_OP_424J2_126_3477_n1477), .CI(DP_OP_424J2_126_3477_n1618), .CO(
        DP_OP_424J2_126_3477_n1434), .S(DP_OP_424J2_126_3477_n1435) );
  FADDX1_HVT DP_OP_424J2_126_3477_U899 ( .A(DP_OP_424J2_126_3477_n1616), .B(
        DP_OP_424J2_126_3477_n1463), .CI(DP_OP_424J2_126_3477_n1614), .CO(
        DP_OP_424J2_126_3477_n1432), .S(DP_OP_424J2_126_3477_n1433) );
  FADDX1_HVT DP_OP_424J2_126_3477_U898 ( .A(DP_OP_424J2_126_3477_n1612), .B(
        DP_OP_424J2_126_3477_n1459), .CI(DP_OP_424J2_126_3477_n1461), .CO(
        DP_OP_424J2_126_3477_n1430), .S(DP_OP_424J2_126_3477_n1431) );
  FADDX1_HVT DP_OP_424J2_126_3477_U897 ( .A(DP_OP_424J2_126_3477_n1610), .B(
        DP_OP_424J2_126_3477_n1606), .CI(DP_OP_424J2_126_3477_n1608), .CO(
        DP_OP_424J2_126_3477_n1428), .S(DP_OP_424J2_126_3477_n1429) );
  FADDX1_HVT DP_OP_424J2_126_3477_U896 ( .A(DP_OP_424J2_126_3477_n1457), .B(
        DP_OP_424J2_126_3477_n1604), .CI(DP_OP_424J2_126_3477_n1602), .CO(
        DP_OP_424J2_126_3477_n1426), .S(DP_OP_424J2_126_3477_n1427) );
  FADDX1_HVT DP_OP_424J2_126_3477_U894 ( .A(DP_OP_424J2_126_3477_n1451), .B(
        DP_OP_424J2_126_3477_n1447), .CI(DP_OP_424J2_126_3477_n1443), .CO(
        DP_OP_424J2_126_3477_n1422), .S(DP_OP_424J2_126_3477_n1423) );
  FADDX1_HVT DP_OP_424J2_126_3477_U893 ( .A(DP_OP_424J2_126_3477_n1600), .B(
        DP_OP_424J2_126_3477_n1445), .CI(DP_OP_424J2_126_3477_n1598), .CO(
        DP_OP_424J2_126_3477_n1420), .S(DP_OP_424J2_126_3477_n1421) );
  FADDX1_HVT DP_OP_424J2_126_3477_U892 ( .A(DP_OP_424J2_126_3477_n1441), .B(
        DP_OP_424J2_126_3477_n1439), .CI(DP_OP_424J2_126_3477_n1437), .CO(
        DP_OP_424J2_126_3477_n1418), .S(DP_OP_424J2_126_3477_n1419) );
  FADDX1_HVT DP_OP_424J2_126_3477_U891 ( .A(DP_OP_424J2_126_3477_n1596), .B(
        DP_OP_424J2_126_3477_n1435), .CI(DP_OP_424J2_126_3477_n1594), .CO(
        DP_OP_424J2_126_3477_n1416), .S(DP_OP_424J2_126_3477_n1417) );
  FADDX1_HVT DP_OP_424J2_126_3477_U890 ( .A(DP_OP_424J2_126_3477_n1433), .B(
        DP_OP_424J2_126_3477_n1592), .CI(DP_OP_424J2_126_3477_n1590), .CO(
        DP_OP_424J2_126_3477_n1414), .S(DP_OP_424J2_126_3477_n1415) );
  FADDX1_HVT DP_OP_424J2_126_3477_U889 ( .A(DP_OP_424J2_126_3477_n1429), .B(
        DP_OP_424J2_126_3477_n1431), .CI(DP_OP_424J2_126_3477_n1588), .CO(
        DP_OP_424J2_126_3477_n1412), .S(DP_OP_424J2_126_3477_n1413) );
  FADDX1_HVT DP_OP_424J2_126_3477_U888 ( .A(DP_OP_424J2_126_3477_n1427), .B(
        DP_OP_424J2_126_3477_n1425), .CI(DP_OP_424J2_126_3477_n1586), .CO(
        DP_OP_424J2_126_3477_n1410), .S(DP_OP_424J2_126_3477_n1411) );
  FADDX1_HVT DP_OP_424J2_126_3477_U887 ( .A(DP_OP_424J2_126_3477_n1421), .B(
        DP_OP_424J2_126_3477_n1423), .CI(DP_OP_424J2_126_3477_n1584), .CO(
        DP_OP_424J2_126_3477_n1408), .S(DP_OP_424J2_126_3477_n1409) );
  FADDX1_HVT DP_OP_424J2_126_3477_U886 ( .A(DP_OP_424J2_126_3477_n1419), .B(
        DP_OP_424J2_126_3477_n1417), .CI(DP_OP_424J2_126_3477_n1582), .CO(
        DP_OP_424J2_126_3477_n1406), .S(DP_OP_424J2_126_3477_n1407) );
  FADDX1_HVT DP_OP_424J2_126_3477_U885 ( .A(DP_OP_424J2_126_3477_n1415), .B(
        DP_OP_424J2_126_3477_n1580), .CI(DP_OP_424J2_126_3477_n1413), .CO(
        DP_OP_424J2_126_3477_n1404), .S(DP_OP_424J2_126_3477_n1405) );
  FADDX1_HVT DP_OP_424J2_126_3477_U884 ( .A(DP_OP_424J2_126_3477_n1411), .B(
        DP_OP_424J2_126_3477_n1578), .CI(DP_OP_424J2_126_3477_n1409), .CO(
        DP_OP_424J2_126_3477_n1402), .S(DP_OP_424J2_126_3477_n1403) );
  FADDX1_HVT DP_OP_424J2_126_3477_U883 ( .A(DP_OP_424J2_126_3477_n1407), .B(
        DP_OP_424J2_126_3477_n1576), .CI(DP_OP_424J2_126_3477_n1405), .CO(
        DP_OP_424J2_126_3477_n1400), .S(DP_OP_424J2_126_3477_n1401) );
  HADDX1_HVT DP_OP_424J2_126_3477_U882 ( .A0(DP_OP_424J2_126_3477_n3030), .B0(
        DP_OP_424J2_126_3477_n1975), .C1(DP_OP_424J2_126_3477_n1398), .SO(
        DP_OP_424J2_126_3477_n1399) );
  FADDX1_HVT DP_OP_424J2_126_3477_U881 ( .A(DP_OP_424J2_126_3477_n2503), .B(
        DP_OP_424J2_126_3477_n2415), .CI(DP_OP_424J2_126_3477_n1931), .CO(
        DP_OP_424J2_126_3477_n1396), .S(DP_OP_424J2_126_3477_n1397) );
  FADDX1_HVT DP_OP_424J2_126_3477_U880 ( .A(DP_OP_424J2_126_3477_n2547), .B(
        DP_OP_424J2_126_3477_n2327), .CI(DP_OP_424J2_126_3477_n2371), .CO(
        DP_OP_424J2_126_3477_n1394), .S(DP_OP_424J2_126_3477_n1395) );
  FADDX1_HVT DP_OP_424J2_126_3477_U878 ( .A(DP_OP_424J2_126_3477_n2591), .B(
        DP_OP_424J2_126_3477_n2151), .CI(DP_OP_424J2_126_3477_n2679), .CO(
        DP_OP_424J2_126_3477_n1390), .S(DP_OP_424J2_126_3477_n1391) );
  FADDX1_HVT DP_OP_424J2_126_3477_U877 ( .A(DP_OP_424J2_126_3477_n2063), .B(
        DP_OP_424J2_126_3477_n2899), .CI(DP_OP_424J2_126_3477_n2195), .CO(
        DP_OP_424J2_126_3477_n1388), .S(DP_OP_424J2_126_3477_n1389) );
  FADDX1_HVT DP_OP_424J2_126_3477_U876 ( .A(DP_OP_424J2_126_3477_n2459), .B(
        DP_OP_424J2_126_3477_n2943), .CI(DP_OP_424J2_126_3477_n2767), .CO(
        DP_OP_424J2_126_3477_n1386), .S(DP_OP_424J2_126_3477_n1387) );
  FADDX1_HVT DP_OP_424J2_126_3477_U875 ( .A(DP_OP_424J2_126_3477_n2283), .B(
        DP_OP_424J2_126_3477_n2239), .CI(DP_OP_424J2_126_3477_n2723), .CO(
        DP_OP_424J2_126_3477_n1384), .S(DP_OP_424J2_126_3477_n1385) );
  FADDX1_HVT DP_OP_424J2_126_3477_U874 ( .A(DP_OP_424J2_126_3477_n2987), .B(
        DP_OP_424J2_126_3477_n2635), .CI(DP_OP_424J2_126_3477_n2811), .CO(
        DP_OP_424J2_126_3477_n1382), .S(DP_OP_424J2_126_3477_n1383) );
  FADDX1_HVT DP_OP_424J2_126_3477_U873 ( .A(DP_OP_424J2_126_3477_n2429), .B(
        DP_OP_424J2_126_3477_n3050), .CI(DP_OP_424J2_126_3477_n1982), .CO(
        DP_OP_424J2_126_3477_n1380), .S(DP_OP_424J2_126_3477_n1381) );
  FADDX1_HVT DP_OP_424J2_126_3477_U872 ( .A(DP_OP_424J2_126_3477_n2422), .B(
        DP_OP_424J2_126_3477_n1989), .CI(DP_OP_424J2_126_3477_n1996), .CO(
        DP_OP_424J2_126_3477_n1378), .S(DP_OP_424J2_126_3477_n1379) );
  FADDX1_HVT DP_OP_424J2_126_3477_U871 ( .A(DP_OP_424J2_126_3477_n2436), .B(
        DP_OP_424J2_126_3477_n2026), .CI(DP_OP_424J2_126_3477_n3043), .CO(
        DP_OP_424J2_126_3477_n1376), .S(DP_OP_424J2_126_3477_n1377) );
  FADDX1_HVT DP_OP_424J2_126_3477_U870 ( .A(DP_OP_424J2_126_3477_n2392), .B(
        DP_OP_424J2_126_3477_n3036), .CI(DP_OP_424J2_126_3477_n3008), .CO(
        DP_OP_424J2_126_3477_n1374), .S(DP_OP_424J2_126_3477_n1375) );
  FADDX1_HVT DP_OP_424J2_126_3477_U869 ( .A(DP_OP_424J2_126_3477_n2385), .B(
        DP_OP_424J2_126_3477_n3001), .CI(DP_OP_424J2_126_3477_n2994), .CO(
        DP_OP_424J2_126_3477_n1372), .S(DP_OP_424J2_126_3477_n1373) );
  FADDX1_HVT DP_OP_424J2_126_3477_U868 ( .A(DP_OP_424J2_126_3477_n2348), .B(
        DP_OP_424J2_126_3477_n2964), .CI(DP_OP_424J2_126_3477_n2957), .CO(
        DP_OP_424J2_126_3477_n1370), .S(DP_OP_424J2_126_3477_n1371) );
  FADDX1_HVT DP_OP_424J2_126_3477_U866 ( .A(DP_OP_424J2_126_3477_n2334), .B(
        DP_OP_424J2_126_3477_n2920), .CI(DP_OP_424J2_126_3477_n2913), .CO(
        DP_OP_424J2_126_3477_n1366), .S(DP_OP_424J2_126_3477_n1367) );
  FADDX1_HVT DP_OP_424J2_126_3477_U865 ( .A(DP_OP_424J2_126_3477_n2304), .B(
        DP_OP_424J2_126_3477_n2906), .CI(DP_OP_424J2_126_3477_n2040), .CO(
        DP_OP_424J2_126_3477_n1364), .S(DP_OP_424J2_126_3477_n1365) );
  FADDX1_HVT DP_OP_424J2_126_3477_U864 ( .A(DP_OP_424J2_126_3477_n2297), .B(
        DP_OP_424J2_126_3477_n2070), .CI(DP_OP_424J2_126_3477_n2077), .CO(
        DP_OP_424J2_126_3477_n1362), .S(DP_OP_424J2_126_3477_n1363) );
  FADDX1_HVT DP_OP_424J2_126_3477_U863 ( .A(DP_OP_424J2_126_3477_n2378), .B(
        DP_OP_424J2_126_3477_n2084), .CI(DP_OP_424J2_126_3477_n2876), .CO(
        DP_OP_424J2_126_3477_n1360), .S(DP_OP_424J2_126_3477_n1361) );
  FADDX1_HVT DP_OP_424J2_126_3477_U862 ( .A(DP_OP_424J2_126_3477_n2466), .B(
        DP_OP_424J2_126_3477_n2869), .CI(DP_OP_424J2_126_3477_n2114), .CO(
        DP_OP_424J2_126_3477_n1358), .S(DP_OP_424J2_126_3477_n1359) );
  FADDX1_HVT DP_OP_424J2_126_3477_U861 ( .A(DP_OP_424J2_126_3477_n2862), .B(
        DP_OP_424J2_126_3477_n2121), .CI(DP_OP_424J2_126_3477_n2128), .CO(
        DP_OP_424J2_126_3477_n1356), .S(DP_OP_424J2_126_3477_n1357) );
  FADDX1_HVT DP_OP_424J2_126_3477_U860 ( .A(DP_OP_424J2_126_3477_n2832), .B(
        DP_OP_424J2_126_3477_n2158), .CI(DP_OP_424J2_126_3477_n2165), .CO(
        DP_OP_424J2_126_3477_n1354), .S(DP_OP_424J2_126_3477_n1355) );
  FADDX1_HVT DP_OP_424J2_126_3477_U859 ( .A(DP_OP_424J2_126_3477_n2825), .B(
        DP_OP_424J2_126_3477_n2172), .CI(DP_OP_424J2_126_3477_n2202), .CO(
        DP_OP_424J2_126_3477_n1352), .S(DP_OP_424J2_126_3477_n1353) );
  FADDX1_HVT DP_OP_424J2_126_3477_U858 ( .A(DP_OP_424J2_126_3477_n2818), .B(
        DP_OP_424J2_126_3477_n2209), .CI(DP_OP_424J2_126_3477_n2216), .CO(
        DP_OP_424J2_126_3477_n1350), .S(DP_OP_424J2_126_3477_n1351) );
  FADDX1_HVT DP_OP_424J2_126_3477_U857 ( .A(DP_OP_424J2_126_3477_n2788), .B(
        DP_OP_424J2_126_3477_n2246), .CI(DP_OP_424J2_126_3477_n2253), .CO(
        DP_OP_424J2_126_3477_n1348), .S(DP_OP_424J2_126_3477_n1349) );
  FADDX1_HVT DP_OP_424J2_126_3477_U855 ( .A(DP_OP_424J2_126_3477_n2774), .B(
        DP_OP_424J2_126_3477_n2473), .CI(DP_OP_424J2_126_3477_n2480), .CO(
        DP_OP_424J2_126_3477_n1344), .S(DP_OP_424J2_126_3477_n1345) );
  FADDX1_HVT DP_OP_424J2_126_3477_U854 ( .A(DP_OP_424J2_126_3477_n2744), .B(
        DP_OP_424J2_126_3477_n2510), .CI(DP_OP_424J2_126_3477_n2517), .CO(
        DP_OP_424J2_126_3477_n1342), .S(DP_OP_424J2_126_3477_n1343) );
  FADDX1_HVT DP_OP_424J2_126_3477_U853 ( .A(DP_OP_424J2_126_3477_n2737), .B(
        DP_OP_424J2_126_3477_n2524), .CI(DP_OP_424J2_126_3477_n2554), .CO(
        DP_OP_424J2_126_3477_n1340), .S(DP_OP_424J2_126_3477_n1341) );
  FADDX1_HVT DP_OP_424J2_126_3477_U852 ( .A(DP_OP_424J2_126_3477_n2730), .B(
        DP_OP_424J2_126_3477_n2561), .CI(DP_OP_424J2_126_3477_n2568), .CO(
        DP_OP_424J2_126_3477_n1338), .S(DP_OP_424J2_126_3477_n1339) );
  FADDX1_HVT DP_OP_424J2_126_3477_U851 ( .A(DP_OP_424J2_126_3477_n2700), .B(
        DP_OP_424J2_126_3477_n2693), .CI(DP_OP_424J2_126_3477_n2686), .CO(
        DP_OP_424J2_126_3477_n1336), .S(DP_OP_424J2_126_3477_n1337) );
  FADDX1_HVT DP_OP_424J2_126_3477_U850 ( .A(DP_OP_424J2_126_3477_n2642), .B(
        DP_OP_424J2_126_3477_n2656), .CI(DP_OP_424J2_126_3477_n2598), .CO(
        DP_OP_424J2_126_3477_n1334), .S(DP_OP_424J2_126_3477_n1335) );
  FADDX1_HVT DP_OP_424J2_126_3477_U849 ( .A(DP_OP_424J2_126_3477_n2605), .B(
        DP_OP_424J2_126_3477_n2612), .CI(DP_OP_424J2_126_3477_n2649), .CO(
        DP_OP_424J2_126_3477_n1332), .S(DP_OP_424J2_126_3477_n1333) );
  FADDX1_HVT DP_OP_424J2_126_3477_U848 ( .A(DP_OP_424J2_126_3477_n1399), .B(
        DP_OP_424J2_126_3477_n1574), .CI(DP_OP_424J2_126_3477_n1564), .CO(
        DP_OP_424J2_126_3477_n1330), .S(DP_OP_424J2_126_3477_n1331) );
  FADDX1_HVT DP_OP_424J2_126_3477_U847 ( .A(DP_OP_424J2_126_3477_n1572), .B(
        DP_OP_424J2_126_3477_n1570), .CI(DP_OP_424J2_126_3477_n1568), .CO(
        DP_OP_424J2_126_3477_n1328), .S(DP_OP_424J2_126_3477_n1329) );
  FADDX1_HVT DP_OP_424J2_126_3477_U846 ( .A(DP_OP_424J2_126_3477_n1566), .B(
        DP_OP_424J2_126_3477_n1562), .CI(DP_OP_424J2_126_3477_n1558), .CO(
        DP_OP_424J2_126_3477_n1326), .S(DP_OP_424J2_126_3477_n1327) );
  FADDX1_HVT DP_OP_424J2_126_3477_U845 ( .A(DP_OP_424J2_126_3477_n1560), .B(
        DP_OP_424J2_126_3477_n1534), .CI(DP_OP_424J2_126_3477_n1532), .CO(
        DP_OP_424J2_126_3477_n1324), .S(DP_OP_424J2_126_3477_n1325) );
  FADDX1_HVT DP_OP_424J2_126_3477_U844 ( .A(DP_OP_424J2_126_3477_n1536), .B(
        DP_OP_424J2_126_3477_n1508), .CI(DP_OP_424J2_126_3477_n1556), .CO(
        DP_OP_424J2_126_3477_n1322), .S(DP_OP_424J2_126_3477_n1323) );
  FADDX1_HVT DP_OP_424J2_126_3477_U843 ( .A(DP_OP_424J2_126_3477_n1528), .B(
        DP_OP_424J2_126_3477_n1554), .CI(DP_OP_424J2_126_3477_n1552), .CO(
        DP_OP_424J2_126_3477_n1320), .S(DP_OP_424J2_126_3477_n1321) );
  FADDX1_HVT DP_OP_424J2_126_3477_U842 ( .A(DP_OP_424J2_126_3477_n1524), .B(
        DP_OP_424J2_126_3477_n1550), .CI(DP_OP_424J2_126_3477_n1548), .CO(
        DP_OP_424J2_126_3477_n1318), .S(DP_OP_424J2_126_3477_n1319) );
  FADDX1_HVT DP_OP_424J2_126_3477_U841 ( .A(DP_OP_424J2_126_3477_n1518), .B(
        DP_OP_424J2_126_3477_n1510), .CI(DP_OP_424J2_126_3477_n1512), .CO(
        DP_OP_424J2_126_3477_n1316), .S(DP_OP_424J2_126_3477_n1317) );
  FADDX1_HVT DP_OP_424J2_126_3477_U840 ( .A(DP_OP_424J2_126_3477_n1516), .B(
        DP_OP_424J2_126_3477_n1546), .CI(DP_OP_424J2_126_3477_n1544), .CO(
        DP_OP_424J2_126_3477_n1314), .S(DP_OP_424J2_126_3477_n1315) );
  FADDX1_HVT DP_OP_424J2_126_3477_U839 ( .A(DP_OP_424J2_126_3477_n1526), .B(
        DP_OP_424J2_126_3477_n1542), .CI(DP_OP_424J2_126_3477_n1514), .CO(
        DP_OP_424J2_126_3477_n1312), .S(DP_OP_424J2_126_3477_n1313) );
  FADDX1_HVT DP_OP_424J2_126_3477_U838 ( .A(DP_OP_424J2_126_3477_n1522), .B(
        DP_OP_424J2_126_3477_n1540), .CI(DP_OP_424J2_126_3477_n1538), .CO(
        DP_OP_424J2_126_3477_n1310), .S(DP_OP_424J2_126_3477_n1311) );
  FADDX1_HVT DP_OP_424J2_126_3477_U837 ( .A(DP_OP_424J2_126_3477_n1389), .B(
        DP_OP_424J2_126_3477_n1530), .CI(DP_OP_424J2_126_3477_n1520), .CO(
        DP_OP_424J2_126_3477_n1308), .S(DP_OP_424J2_126_3477_n1309) );
  FADDX1_HVT DP_OP_424J2_126_3477_U836 ( .A(DP_OP_424J2_126_3477_n1391), .B(
        DP_OP_424J2_126_3477_n1383), .CI(DP_OP_424J2_126_3477_n1385), .CO(
        DP_OP_424J2_126_3477_n1306), .S(DP_OP_424J2_126_3477_n1307) );
  FADDX1_HVT DP_OP_424J2_126_3477_U835 ( .A(DP_OP_424J2_126_3477_n1395), .B(
        DP_OP_424J2_126_3477_n1393), .CI(DP_OP_424J2_126_3477_n1397), .CO(
        DP_OP_424J2_126_3477_n1304), .S(DP_OP_424J2_126_3477_n1305) );
  FADDX1_HVT DP_OP_424J2_126_3477_U834 ( .A(DP_OP_424J2_126_3477_n1387), .B(
        DP_OP_424J2_126_3477_n1339), .CI(DP_OP_424J2_126_3477_n1337), .CO(
        DP_OP_424J2_126_3477_n1302), .S(DP_OP_424J2_126_3477_n1303) );
  FADDX1_HVT DP_OP_424J2_126_3477_U833 ( .A(DP_OP_424J2_126_3477_n1333), .B(
        DP_OP_424J2_126_3477_n1381), .CI(DP_OP_424J2_126_3477_n1379), .CO(
        DP_OP_424J2_126_3477_n1300), .S(DP_OP_424J2_126_3477_n1301) );
  FADDX1_HVT DP_OP_424J2_126_3477_U832 ( .A(DP_OP_424J2_126_3477_n1369), .B(
        DP_OP_424J2_126_3477_n1359), .CI(DP_OP_424J2_126_3477_n1365), .CO(
        DP_OP_424J2_126_3477_n1298), .S(DP_OP_424J2_126_3477_n1299) );
  FADDX1_HVT DP_OP_424J2_126_3477_U831 ( .A(DP_OP_424J2_126_3477_n1363), .B(
        DP_OP_424J2_126_3477_n1361), .CI(DP_OP_424J2_126_3477_n1345), .CO(
        DP_OP_424J2_126_3477_n1296), .S(DP_OP_424J2_126_3477_n1297) );
  FADDX1_HVT DP_OP_424J2_126_3477_U830 ( .A(DP_OP_424J2_126_3477_n1367), .B(
        DP_OP_424J2_126_3477_n1341), .CI(DP_OP_424J2_126_3477_n1335), .CO(
        DP_OP_424J2_126_3477_n1294), .S(DP_OP_424J2_126_3477_n1295) );
  FADDX1_HVT DP_OP_424J2_126_3477_U829 ( .A(DP_OP_424J2_126_3477_n1371), .B(
        DP_OP_424J2_126_3477_n1353), .CI(DP_OP_424J2_126_3477_n1355), .CO(
        DP_OP_424J2_126_3477_n1292), .S(DP_OP_424J2_126_3477_n1293) );
  FADDX1_HVT DP_OP_424J2_126_3477_U828 ( .A(DP_OP_424J2_126_3477_n1351), .B(
        DP_OP_424J2_126_3477_n1349), .CI(DP_OP_424J2_126_3477_n1343), .CO(
        DP_OP_424J2_126_3477_n1290), .S(DP_OP_424J2_126_3477_n1291) );
  FADDX1_HVT DP_OP_424J2_126_3477_U827 ( .A(DP_OP_424J2_126_3477_n1347), .B(
        DP_OP_424J2_126_3477_n1377), .CI(DP_OP_424J2_126_3477_n1373), .CO(
        DP_OP_424J2_126_3477_n1288), .S(DP_OP_424J2_126_3477_n1289) );
  FADDX1_HVT DP_OP_424J2_126_3477_U826 ( .A(DP_OP_424J2_126_3477_n1375), .B(
        DP_OP_424J2_126_3477_n1357), .CI(DP_OP_424J2_126_3477_n1506), .CO(
        DP_OP_424J2_126_3477_n1286), .S(DP_OP_424J2_126_3477_n1287) );
  FADDX1_HVT DP_OP_424J2_126_3477_U825 ( .A(DP_OP_424J2_126_3477_n1504), .B(
        DP_OP_424J2_126_3477_n1502), .CI(DP_OP_424J2_126_3477_n1500), .CO(
        DP_OP_424J2_126_3477_n1284), .S(DP_OP_424J2_126_3477_n1285) );
  FADDX1_HVT DP_OP_424J2_126_3477_U824 ( .A(DP_OP_424J2_126_3477_n1498), .B(
        DP_OP_424J2_126_3477_n1486), .CI(DP_OP_424J2_126_3477_n1488), .CO(
        DP_OP_424J2_126_3477_n1282), .S(DP_OP_424J2_126_3477_n1283) );
  FADDX1_HVT DP_OP_424J2_126_3477_U823 ( .A(DP_OP_424J2_126_3477_n1492), .B(
        DP_OP_424J2_126_3477_n1496), .CI(DP_OP_424J2_126_3477_n1490), .CO(
        DP_OP_424J2_126_3477_n1280), .S(DP_OP_424J2_126_3477_n1281) );
  FADDX1_HVT DP_OP_424J2_126_3477_U822 ( .A(DP_OP_424J2_126_3477_n1494), .B(
        DP_OP_424J2_126_3477_n1331), .CI(DP_OP_424J2_126_3477_n1484), .CO(
        DP_OP_424J2_126_3477_n1278), .S(DP_OP_424J2_126_3477_n1279) );
  FADDX1_HVT DP_OP_424J2_126_3477_U821 ( .A(DP_OP_424J2_126_3477_n1329), .B(
        DP_OP_424J2_126_3477_n1327), .CI(DP_OP_424J2_126_3477_n1325), .CO(
        DP_OP_424J2_126_3477_n1276), .S(DP_OP_424J2_126_3477_n1277) );
  FADDX1_HVT DP_OP_424J2_126_3477_U820 ( .A(DP_OP_424J2_126_3477_n1482), .B(
        DP_OP_424J2_126_3477_n1480), .CI(DP_OP_424J2_126_3477_n1478), .CO(
        DP_OP_424J2_126_3477_n1274), .S(DP_OP_424J2_126_3477_n1275) );
  FADDX1_HVT DP_OP_424J2_126_3477_U819 ( .A(DP_OP_424J2_126_3477_n1466), .B(
        DP_OP_424J2_126_3477_n1311), .CI(DP_OP_424J2_126_3477_n1309), .CO(
        DP_OP_424J2_126_3477_n1272), .S(DP_OP_424J2_126_3477_n1273) );
  FADDX1_HVT DP_OP_424J2_126_3477_U818 ( .A(DP_OP_424J2_126_3477_n1476), .B(
        DP_OP_424J2_126_3477_n1321), .CI(DP_OP_424J2_126_3477_n1323), .CO(
        DP_OP_424J2_126_3477_n1270), .S(DP_OP_424J2_126_3477_n1271) );
  FADDX1_HVT DP_OP_424J2_126_3477_U816 ( .A(DP_OP_424J2_126_3477_n1472), .B(
        DP_OP_424J2_126_3477_n1319), .CI(DP_OP_424J2_126_3477_n1315), .CO(
        DP_OP_424J2_126_3477_n1266), .S(DP_OP_424J2_126_3477_n1267) );
  FADDX1_HVT DP_OP_424J2_126_3477_U815 ( .A(DP_OP_424J2_126_3477_n1470), .B(
        DP_OP_424J2_126_3477_n1464), .CI(DP_OP_424J2_126_3477_n1468), .CO(
        DP_OP_424J2_126_3477_n1264), .S(DP_OP_424J2_126_3477_n1265) );
  FADDX1_HVT DP_OP_424J2_126_3477_U814 ( .A(DP_OP_424J2_126_3477_n1305), .B(
        DP_OP_424J2_126_3477_n1307), .CI(DP_OP_424J2_126_3477_n1303), .CO(
        DP_OP_424J2_126_3477_n1262), .S(DP_OP_424J2_126_3477_n1263) );
  FADDX1_HVT DP_OP_424J2_126_3477_U813 ( .A(DP_OP_424J2_126_3477_n1295), .B(
        DP_OP_424J2_126_3477_n1297), .CI(DP_OP_424J2_126_3477_n1462), .CO(
        DP_OP_424J2_126_3477_n1260), .S(DP_OP_424J2_126_3477_n1261) );
  FADDX1_HVT DP_OP_424J2_126_3477_U812 ( .A(DP_OP_424J2_126_3477_n1293), .B(
        DP_OP_424J2_126_3477_n1301), .CI(DP_OP_424J2_126_3477_n1299), .CO(
        DP_OP_424J2_126_3477_n1258), .S(DP_OP_424J2_126_3477_n1259) );
  FADDX1_HVT DP_OP_424J2_126_3477_U811 ( .A(DP_OP_424J2_126_3477_n1289), .B(
        DP_OP_424J2_126_3477_n1291), .CI(DP_OP_424J2_126_3477_n1458), .CO(
        DP_OP_424J2_126_3477_n1256), .S(DP_OP_424J2_126_3477_n1257) );
  FADDX1_HVT DP_OP_424J2_126_3477_U810 ( .A(DP_OP_424J2_126_3477_n1287), .B(
        DP_OP_424J2_126_3477_n1460), .CI(DP_OP_424J2_126_3477_n1456), .CO(
        DP_OP_424J2_126_3477_n1254), .S(DP_OP_424J2_126_3477_n1255) );
  FADDX1_HVT DP_OP_424J2_126_3477_U809 ( .A(DP_OP_424J2_126_3477_n1454), .B(
        DP_OP_424J2_126_3477_n1452), .CI(DP_OP_424J2_126_3477_n1285), .CO(
        DP_OP_424J2_126_3477_n1252), .S(DP_OP_424J2_126_3477_n1253) );
  FADDX1_HVT DP_OP_424J2_126_3477_U808 ( .A(DP_OP_424J2_126_3477_n1450), .B(
        DP_OP_424J2_126_3477_n1442), .CI(DP_OP_424J2_126_3477_n1279), .CO(
        DP_OP_424J2_126_3477_n1250), .S(DP_OP_424J2_126_3477_n1251) );
  FADDX1_HVT DP_OP_424J2_126_3477_U807 ( .A(DP_OP_424J2_126_3477_n1448), .B(
        DP_OP_424J2_126_3477_n1281), .CI(DP_OP_424J2_126_3477_n1283), .CO(
        DP_OP_424J2_126_3477_n1248), .S(DP_OP_424J2_126_3477_n1249) );
  FADDX1_HVT DP_OP_424J2_126_3477_U806 ( .A(DP_OP_424J2_126_3477_n1446), .B(
        DP_OP_424J2_126_3477_n1444), .CI(DP_OP_424J2_126_3477_n1440), .CO(
        DP_OP_424J2_126_3477_n1246), .S(DP_OP_424J2_126_3477_n1247) );
  FADDX1_HVT DP_OP_424J2_126_3477_U805 ( .A(DP_OP_424J2_126_3477_n1275), .B(
        DP_OP_424J2_126_3477_n1277), .CI(DP_OP_424J2_126_3477_n1438), .CO(
        DP_OP_424J2_126_3477_n1244), .S(DP_OP_424J2_126_3477_n1245) );
  FADDX1_HVT DP_OP_424J2_126_3477_U804 ( .A(DP_OP_424J2_126_3477_n1436), .B(
        DP_OP_424J2_126_3477_n1269), .CI(DP_OP_424J2_126_3477_n1434), .CO(
        DP_OP_424J2_126_3477_n1242), .S(DP_OP_424J2_126_3477_n1243) );
  FADDX1_HVT DP_OP_424J2_126_3477_U802 ( .A(DP_OP_424J2_126_3477_n1265), .B(
        DP_OP_424J2_126_3477_n1263), .CI(DP_OP_424J2_126_3477_n1259), .CO(
        DP_OP_424J2_126_3477_n1238), .S(DP_OP_424J2_126_3477_n1239) );
  FADDX1_HVT DP_OP_424J2_126_3477_U801 ( .A(DP_OP_424J2_126_3477_n1261), .B(
        DP_OP_424J2_126_3477_n1432), .CI(DP_OP_424J2_126_3477_n1257), .CO(
        DP_OP_424J2_126_3477_n1236), .S(DP_OP_424J2_126_3477_n1237) );
  FADDX1_HVT DP_OP_424J2_126_3477_U800 ( .A(DP_OP_424J2_126_3477_n1430), .B(
        DP_OP_424J2_126_3477_n1428), .CI(DP_OP_424J2_126_3477_n1255), .CO(
        DP_OP_424J2_126_3477_n1234), .S(DP_OP_424J2_126_3477_n1235) );
  FADDX1_HVT DP_OP_424J2_126_3477_U799 ( .A(DP_OP_424J2_126_3477_n1426), .B(
        DP_OP_424J2_126_3477_n1424), .CI(DP_OP_424J2_126_3477_n1253), .CO(
        DP_OP_424J2_126_3477_n1232), .S(DP_OP_424J2_126_3477_n1233) );
  FADDX1_HVT DP_OP_424J2_126_3477_U798 ( .A(DP_OP_424J2_126_3477_n1422), .B(
        DP_OP_424J2_126_3477_n1249), .CI(DP_OP_424J2_126_3477_n1247), .CO(
        DP_OP_424J2_126_3477_n1230), .S(DP_OP_424J2_126_3477_n1231) );
  FADDX1_HVT DP_OP_424J2_126_3477_U797 ( .A(DP_OP_424J2_126_3477_n1420), .B(
        DP_OP_424J2_126_3477_n1251), .CI(DP_OP_424J2_126_3477_n1245), .CO(
        DP_OP_424J2_126_3477_n1228), .S(DP_OP_424J2_126_3477_n1229) );
  FADDX1_HVT DP_OP_424J2_126_3477_U796 ( .A(DP_OP_424J2_126_3477_n1418), .B(
        DP_OP_424J2_126_3477_n1241), .CI(DP_OP_424J2_126_3477_n1416), .CO(
        DP_OP_424J2_126_3477_n1226), .S(DP_OP_424J2_126_3477_n1227) );
  FADDX1_HVT DP_OP_424J2_126_3477_U795 ( .A(DP_OP_424J2_126_3477_n1243), .B(
        DP_OP_424J2_126_3477_n1239), .CI(DP_OP_424J2_126_3477_n1237), .CO(
        DP_OP_424J2_126_3477_n1224), .S(DP_OP_424J2_126_3477_n1225) );
  FADDX1_HVT DP_OP_424J2_126_3477_U794 ( .A(DP_OP_424J2_126_3477_n1414), .B(
        DP_OP_424J2_126_3477_n1235), .CI(DP_OP_424J2_126_3477_n1412), .CO(
        DP_OP_424J2_126_3477_n1222), .S(DP_OP_424J2_126_3477_n1223) );
  FADDX1_HVT DP_OP_424J2_126_3477_U793 ( .A(DP_OP_424J2_126_3477_n1233), .B(
        DP_OP_424J2_126_3477_n1410), .CI(DP_OP_424J2_126_3477_n1231), .CO(
        DP_OP_424J2_126_3477_n1220), .S(DP_OP_424J2_126_3477_n1221) );
  FADDX1_HVT DP_OP_424J2_126_3477_U792 ( .A(DP_OP_424J2_126_3477_n1229), .B(
        DP_OP_424J2_126_3477_n1408), .CI(DP_OP_424J2_126_3477_n1227), .CO(
        DP_OP_424J2_126_3477_n1218), .S(DP_OP_424J2_126_3477_n1219) );
  FADDX1_HVT DP_OP_424J2_126_3477_U791 ( .A(DP_OP_424J2_126_3477_n1406), .B(
        DP_OP_424J2_126_3477_n1225), .CI(DP_OP_424J2_126_3477_n1404), .CO(
        DP_OP_424J2_126_3477_n1216), .S(DP_OP_424J2_126_3477_n1217) );
  FADDX1_HVT DP_OP_424J2_126_3477_U790 ( .A(DP_OP_424J2_126_3477_n1223), .B(
        DP_OP_424J2_126_3477_n1221), .CI(DP_OP_424J2_126_3477_n1402), .CO(
        DP_OP_424J2_126_3477_n1214), .S(DP_OP_424J2_126_3477_n1215) );
  FADDX1_HVT DP_OP_424J2_126_3477_U789 ( .A(DP_OP_424J2_126_3477_n1219), .B(
        DP_OP_424J2_126_3477_n1217), .CI(DP_OP_424J2_126_3477_n1400), .CO(
        DP_OP_424J2_126_3477_n1212), .S(DP_OP_424J2_126_3477_n1213) );
  OR2X1_HVT DP_OP_424J2_126_3477_U788 ( .A1(DP_OP_424J2_126_3477_n3029), .A2(
        DP_OP_424J2_126_3477_n2502), .Y(DP_OP_424J2_126_3477_n1210) );
  FADDX1_HVT DP_OP_424J2_126_3477_U786 ( .A(DP_OP_424J2_126_3477_n2194), .B(
        DP_OP_424J2_126_3477_n1974), .CI(DP_OP_424J2_126_3477_n1930), .CO(
        DP_OP_424J2_126_3477_n1208), .S(DP_OP_424J2_126_3477_n1209) );
  FADDX1_HVT DP_OP_424J2_126_3477_U785 ( .A(DP_OP_424J2_126_3477_n2634), .B(
        DP_OP_424J2_126_3477_n2062), .CI(DP_OP_424J2_126_3477_n2414), .CO(
        DP_OP_424J2_126_3477_n1206), .S(DP_OP_424J2_126_3477_n1207) );
  FADDX1_HVT DP_OP_424J2_126_3477_U784 ( .A(DP_OP_424J2_126_3477_n2854), .B(
        DP_OP_424J2_126_3477_n2678), .CI(DP_OP_424J2_126_3477_n2238), .CO(
        DP_OP_424J2_126_3477_n1204), .S(DP_OP_424J2_126_3477_n1205) );
  FADDX1_HVT DP_OP_424J2_126_3477_U783 ( .A(DP_OP_424J2_126_3477_n2326), .B(
        DP_OP_424J2_126_3477_n2150), .CI(DP_OP_424J2_126_3477_n2898), .CO(
        DP_OP_424J2_126_3477_n1202), .S(DP_OP_424J2_126_3477_n1203) );
  FADDX1_HVT DP_OP_424J2_126_3477_U782 ( .A(DP_OP_424J2_126_3477_n2458), .B(
        DP_OP_424J2_126_3477_n2942), .CI(DP_OP_424J2_126_3477_n2722), .CO(
        DP_OP_424J2_126_3477_n1200), .S(DP_OP_424J2_126_3477_n1201) );
  FADDX1_HVT DP_OP_424J2_126_3477_U781 ( .A(DP_OP_424J2_126_3477_n2546), .B(
        DP_OP_424J2_126_3477_n2766), .CI(DP_OP_424J2_126_3477_n2590), .CO(
        DP_OP_424J2_126_3477_n1198), .S(DP_OP_424J2_126_3477_n1199) );
  FADDX1_HVT DP_OP_424J2_126_3477_U780 ( .A(DP_OP_424J2_126_3477_n2282), .B(
        DP_OP_424J2_126_3477_n2106), .CI(DP_OP_424J2_126_3477_n2986), .CO(
        DP_OP_424J2_126_3477_n1196), .S(DP_OP_424J2_126_3477_n1197) );
  FADDX1_HVT DP_OP_424J2_126_3477_U779 ( .A(DP_OP_424J2_126_3477_n2810), .B(
        DP_OP_424J2_126_3477_n2018), .CI(DP_OP_424J2_126_3477_n2370), .CO(
        DP_OP_424J2_126_3477_n1194), .S(DP_OP_424J2_126_3477_n1195) );
  FADDX1_HVT DP_OP_424J2_126_3477_U778 ( .A(DP_OP_424J2_126_3477_n2421), .B(
        DP_OP_424J2_126_3477_n3049), .CI(DP_OP_424J2_126_3477_n1981), .CO(
        DP_OP_424J2_126_3477_n1192), .S(DP_OP_424J2_126_3477_n1193) );
  FADDX1_HVT DP_OP_424J2_126_3477_U777 ( .A(DP_OP_424J2_126_3477_n2428), .B(
        DP_OP_424J2_126_3477_n3042), .CI(DP_OP_424J2_126_3477_n3035), .CO(
        DP_OP_424J2_126_3477_n1190), .S(DP_OP_424J2_126_3477_n1191) );
  FADDX1_HVT DP_OP_424J2_126_3477_U776 ( .A(DP_OP_424J2_126_3477_n2384), .B(
        DP_OP_424J2_126_3477_n3007), .CI(DP_OP_424J2_126_3477_n3000), .CO(
        DP_OP_424J2_126_3477_n1188), .S(DP_OP_424J2_126_3477_n1189) );
  FADDX1_HVT DP_OP_424J2_126_3477_U775 ( .A(DP_OP_424J2_126_3477_n2347), .B(
        DP_OP_424J2_126_3477_n2993), .CI(DP_OP_424J2_126_3477_n2963), .CO(
        DP_OP_424J2_126_3477_n1186), .S(DP_OP_424J2_126_3477_n1187) );
  FADDX1_HVT DP_OP_424J2_126_3477_U774 ( .A(DP_OP_424J2_126_3477_n2340), .B(
        DP_OP_424J2_126_3477_n1988), .CI(DP_OP_424J2_126_3477_n2956), .CO(
        DP_OP_424J2_126_3477_n1184), .S(DP_OP_424J2_126_3477_n1185) );
  FADDX1_HVT DP_OP_424J2_126_3477_U773 ( .A(DP_OP_424J2_126_3477_n2377), .B(
        DP_OP_424J2_126_3477_n2949), .CI(DP_OP_424J2_126_3477_n1995), .CO(
        DP_OP_424J2_126_3477_n1182), .S(DP_OP_424J2_126_3477_n1183) );
  FADDX1_HVT DP_OP_424J2_126_3477_U771 ( .A(DP_OP_424J2_126_3477_n2303), .B(
        DP_OP_424J2_126_3477_n2912), .CI(DP_OP_424J2_126_3477_n2905), .CO(
        DP_OP_424J2_126_3477_n1178), .S(DP_OP_424J2_126_3477_n1179) );
  FADDX1_HVT DP_OP_424J2_126_3477_U770 ( .A(DP_OP_424J2_126_3477_n2296), .B(
        DP_OP_424J2_126_3477_n2032), .CI(DP_OP_424J2_126_3477_n2875), .CO(
        DP_OP_424J2_126_3477_n1176), .S(DP_OP_424J2_126_3477_n1177) );
  FADDX1_HVT DP_OP_424J2_126_3477_U769 ( .A(DP_OP_424J2_126_3477_n2289), .B(
        DP_OP_424J2_126_3477_n2039), .CI(DP_OP_424J2_126_3477_n2868), .CO(
        DP_OP_424J2_126_3477_n1174), .S(DP_OP_424J2_126_3477_n1175) );
  FADDX1_HVT DP_OP_424J2_126_3477_U768 ( .A(DP_OP_424J2_126_3477_n2069), .B(
        DP_OP_424J2_126_3477_n2076), .CI(DP_OP_424J2_126_3477_n2083), .CO(
        DP_OP_424J2_126_3477_n1172), .S(DP_OP_424J2_126_3477_n1173) );
  FADDX1_HVT DP_OP_424J2_126_3477_U767 ( .A(DP_OP_424J2_126_3477_n2861), .B(
        DP_OP_424J2_126_3477_n2113), .CI(DP_OP_424J2_126_3477_n2120), .CO(
        DP_OP_424J2_126_3477_n1170), .S(DP_OP_424J2_126_3477_n1171) );
  FADDX1_HVT DP_OP_424J2_126_3477_U766 ( .A(DP_OP_424J2_126_3477_n2831), .B(
        DP_OP_424J2_126_3477_n2127), .CI(DP_OP_424J2_126_3477_n2157), .CO(
        DP_OP_424J2_126_3477_n1168), .S(DP_OP_424J2_126_3477_n1169) );
  FADDX1_HVT DP_OP_424J2_126_3477_U765 ( .A(DP_OP_424J2_126_3477_n2824), .B(
        DP_OP_424J2_126_3477_n2164), .CI(DP_OP_424J2_126_3477_n2171), .CO(
        DP_OP_424J2_126_3477_n1166), .S(DP_OP_424J2_126_3477_n1167) );
  FADDX1_HVT DP_OP_424J2_126_3477_U764 ( .A(DP_OP_424J2_126_3477_n2817), .B(
        DP_OP_424J2_126_3477_n2201), .CI(DP_OP_424J2_126_3477_n2208), .CO(
        DP_OP_424J2_126_3477_n1164), .S(DP_OP_424J2_126_3477_n1165) );
  FADDX1_HVT DP_OP_424J2_126_3477_U763 ( .A(DP_OP_424J2_126_3477_n2787), .B(
        DP_OP_424J2_126_3477_n2215), .CI(DP_OP_424J2_126_3477_n2245), .CO(
        DP_OP_424J2_126_3477_n1162), .S(DP_OP_424J2_126_3477_n1163) );
  FADDX1_HVT DP_OP_424J2_126_3477_U762 ( .A(DP_OP_424J2_126_3477_n2780), .B(
        DP_OP_424J2_126_3477_n2252), .CI(DP_OP_424J2_126_3477_n2259), .CO(
        DP_OP_424J2_126_3477_n1160), .S(DP_OP_424J2_126_3477_n1161) );
  FADDX1_HVT DP_OP_424J2_126_3477_U761 ( .A(DP_OP_424J2_126_3477_n2773), .B(
        DP_OP_424J2_126_3477_n2391), .CI(DP_OP_424J2_126_3477_n2435), .CO(
        DP_OP_424J2_126_3477_n1158), .S(DP_OP_424J2_126_3477_n1159) );
  FADDX1_HVT DP_OP_424J2_126_3477_U760 ( .A(DP_OP_424J2_126_3477_n2743), .B(
        DP_OP_424J2_126_3477_n2465), .CI(DP_OP_424J2_126_3477_n2472), .CO(
        DP_OP_424J2_126_3477_n1156), .S(DP_OP_424J2_126_3477_n1157) );
  FADDX1_HVT DP_OP_424J2_126_3477_U759 ( .A(DP_OP_424J2_126_3477_n2736), .B(
        DP_OP_424J2_126_3477_n2479), .CI(DP_OP_424J2_126_3477_n2509), .CO(
        DP_OP_424J2_126_3477_n1154), .S(DP_OP_424J2_126_3477_n1155) );
  FADDX1_HVT DP_OP_424J2_126_3477_U758 ( .A(DP_OP_424J2_126_3477_n2729), .B(
        DP_OP_424J2_126_3477_n2516), .CI(DP_OP_424J2_126_3477_n2523), .CO(
        DP_OP_424J2_126_3477_n1152), .S(DP_OP_424J2_126_3477_n1153) );
  FADDX1_HVT DP_OP_424J2_126_3477_U757 ( .A(DP_OP_424J2_126_3477_n2699), .B(
        DP_OP_424J2_126_3477_n2553), .CI(DP_OP_424J2_126_3477_n2560), .CO(
        DP_OP_424J2_126_3477_n1150), .S(DP_OP_424J2_126_3477_n1151) );
  FADDX1_HVT DP_OP_424J2_126_3477_U756 ( .A(DP_OP_424J2_126_3477_n2692), .B(
        DP_OP_424J2_126_3477_n2567), .CI(DP_OP_424J2_126_3477_n2597), .CO(
        DP_OP_424J2_126_3477_n1148), .S(DP_OP_424J2_126_3477_n1149) );
  FADDX1_HVT DP_OP_424J2_126_3477_U755 ( .A(DP_OP_424J2_126_3477_n2685), .B(
        DP_OP_424J2_126_3477_n2604), .CI(DP_OP_424J2_126_3477_n2611), .CO(
        DP_OP_424J2_126_3477_n1146), .S(DP_OP_424J2_126_3477_n1147) );
  FADDX1_HVT DP_OP_424J2_126_3477_U754 ( .A(DP_OP_424J2_126_3477_n2641), .B(
        DP_OP_424J2_126_3477_n2648), .CI(DP_OP_424J2_126_3477_n2655), .CO(
        DP_OP_424J2_126_3477_n1144), .S(DP_OP_424J2_126_3477_n1145) );
  FADDX1_HVT DP_OP_424J2_126_3477_U753 ( .A(DP_OP_424J2_126_3477_n1398), .B(
        DP_OP_424J2_126_3477_n1386), .CI(DP_OP_424J2_126_3477_n1384), .CO(
        DP_OP_424J2_126_3477_n1142), .S(DP_OP_424J2_126_3477_n1143) );
  FADDX1_HVT DP_OP_424J2_126_3477_U752 ( .A(DP_OP_424J2_126_3477_n1382), .B(
        DP_OP_424J2_126_3477_n1211), .CI(DP_OP_424J2_126_3477_n1388), .CO(
        DP_OP_424J2_126_3477_n1140), .S(DP_OP_424J2_126_3477_n1141) );
  FADDX1_HVT DP_OP_424J2_126_3477_U751 ( .A(DP_OP_424J2_126_3477_n1392), .B(
        DP_OP_424J2_126_3477_n1396), .CI(DP_OP_424J2_126_3477_n1390), .CO(
        DP_OP_424J2_126_3477_n1138), .S(DP_OP_424J2_126_3477_n1139) );
  FADDX1_HVT DP_OP_424J2_126_3477_U750 ( .A(DP_OP_424J2_126_3477_n1394), .B(
        DP_OP_424J2_126_3477_n1358), .CI(DP_OP_424J2_126_3477_n1356), .CO(
        DP_OP_424J2_126_3477_n1136), .S(DP_OP_424J2_126_3477_n1137) );
  FADDX1_HVT DP_OP_424J2_126_3477_U749 ( .A(DP_OP_424J2_126_3477_n1360), .B(
        DP_OP_424J2_126_3477_n1332), .CI(DP_OP_424J2_126_3477_n1380), .CO(
        DP_OP_424J2_126_3477_n1134), .S(DP_OP_424J2_126_3477_n1135) );
  FADDX1_HVT DP_OP_424J2_126_3477_U748 ( .A(DP_OP_424J2_126_3477_n1352), .B(
        DP_OP_424J2_126_3477_n1334), .CI(DP_OP_424J2_126_3477_n1378), .CO(
        DP_OP_424J2_126_3477_n1132), .S(DP_OP_424J2_126_3477_n1133) );
  FADDX1_HVT DP_OP_424J2_126_3477_U747 ( .A(DP_OP_424J2_126_3477_n1350), .B(
        DP_OP_424J2_126_3477_n1336), .CI(DP_OP_424J2_126_3477_n1376), .CO(
        DP_OP_424J2_126_3477_n1130), .S(DP_OP_424J2_126_3477_n1131) );
  FADDX1_HVT DP_OP_424J2_126_3477_U746 ( .A(DP_OP_424J2_126_3477_n1346), .B(
        DP_OP_424J2_126_3477_n1374), .CI(DP_OP_424J2_126_3477_n1372), .CO(
        DP_OP_424J2_126_3477_n1128), .S(DP_OP_424J2_126_3477_n1129) );
  FADDX1_HVT DP_OP_424J2_126_3477_U745 ( .A(DP_OP_424J2_126_3477_n1340), .B(
        DP_OP_424J2_126_3477_n1370), .CI(DP_OP_424J2_126_3477_n1368), .CO(
        DP_OP_424J2_126_3477_n1126), .S(DP_OP_424J2_126_3477_n1127) );
  FADDX1_HVT DP_OP_424J2_126_3477_U744 ( .A(DP_OP_424J2_126_3477_n1348), .B(
        DP_OP_424J2_126_3477_n1366), .CI(DP_OP_424J2_126_3477_n1364), .CO(
        DP_OP_424J2_126_3477_n1124), .S(DP_OP_424J2_126_3477_n1125) );
  FADDX1_HVT DP_OP_424J2_126_3477_U743 ( .A(DP_OP_424J2_126_3477_n1342), .B(
        DP_OP_424J2_126_3477_n1362), .CI(DP_OP_424J2_126_3477_n1354), .CO(
        DP_OP_424J2_126_3477_n1122), .S(DP_OP_424J2_126_3477_n1123) );
  FADDX1_HVT DP_OP_424J2_126_3477_U742 ( .A(DP_OP_424J2_126_3477_n1344), .B(
        DP_OP_424J2_126_3477_n1338), .CI(DP_OP_424J2_126_3477_n1201), .CO(
        DP_OP_424J2_126_3477_n1120), .S(DP_OP_424J2_126_3477_n1121) );
  FADDX1_HVT DP_OP_424J2_126_3477_U741 ( .A(DP_OP_424J2_126_3477_n1197), .B(
        DP_OP_424J2_126_3477_n1195), .CI(DP_OP_424J2_126_3477_n1199), .CO(
        DP_OP_424J2_126_3477_n1118), .S(DP_OP_424J2_126_3477_n1119) );
  FADDX1_HVT DP_OP_424J2_126_3477_U740 ( .A(DP_OP_424J2_126_3477_n1207), .B(
        DP_OP_424J2_126_3477_n1205), .CI(DP_OP_424J2_126_3477_n1209), .CO(
        DP_OP_424J2_126_3477_n1116), .S(DP_OP_424J2_126_3477_n1117) );
  FADDX1_HVT DP_OP_424J2_126_3477_U739 ( .A(DP_OP_424J2_126_3477_n1203), .B(
        DP_OP_424J2_126_3477_n1151), .CI(DP_OP_424J2_126_3477_n1153), .CO(
        DP_OP_424J2_126_3477_n1114), .S(DP_OP_424J2_126_3477_n1115) );
  FADDX1_HVT DP_OP_424J2_126_3477_U738 ( .A(DP_OP_424J2_126_3477_n1149), .B(
        DP_OP_424J2_126_3477_n1185), .CI(DP_OP_424J2_126_3477_n1181), .CO(
        DP_OP_424J2_126_3477_n1112), .S(DP_OP_424J2_126_3477_n1113) );
  FADDX1_HVT DP_OP_424J2_126_3477_U737 ( .A(DP_OP_424J2_126_3477_n1187), .B(
        DP_OP_424J2_126_3477_n1171), .CI(DP_OP_424J2_126_3477_n1177), .CO(
        DP_OP_424J2_126_3477_n1110), .S(DP_OP_424J2_126_3477_n1111) );
  FADDX1_HVT DP_OP_424J2_126_3477_U736 ( .A(DP_OP_424J2_126_3477_n1175), .B(
        DP_OP_424J2_126_3477_n1173), .CI(DP_OP_424J2_126_3477_n1157), .CO(
        DP_OP_424J2_126_3477_n1108), .S(DP_OP_424J2_126_3477_n1109) );
  FADDX1_HVT DP_OP_424J2_126_3477_U735 ( .A(DP_OP_424J2_126_3477_n1179), .B(
        DP_OP_424J2_126_3477_n1147), .CI(DP_OP_424J2_126_3477_n1145), .CO(
        DP_OP_424J2_126_3477_n1106), .S(DP_OP_424J2_126_3477_n1107) );
  FADDX1_HVT DP_OP_424J2_126_3477_U734 ( .A(DP_OP_424J2_126_3477_n1183), .B(
        DP_OP_424J2_126_3477_n1165), .CI(DP_OP_424J2_126_3477_n1167), .CO(
        DP_OP_424J2_126_3477_n1104), .S(DP_OP_424J2_126_3477_n1105) );
  FADDX1_HVT DP_OP_424J2_126_3477_U733 ( .A(DP_OP_424J2_126_3477_n1163), .B(
        DP_OP_424J2_126_3477_n1161), .CI(DP_OP_424J2_126_3477_n1155), .CO(
        DP_OP_424J2_126_3477_n1102), .S(DP_OP_424J2_126_3477_n1103) );
  FADDX1_HVT DP_OP_424J2_126_3477_U732 ( .A(DP_OP_424J2_126_3477_n1193), .B(
        DP_OP_424J2_126_3477_n1159), .CI(DP_OP_424J2_126_3477_n1191), .CO(
        DP_OP_424J2_126_3477_n1100), .S(DP_OP_424J2_126_3477_n1101) );
  FADDX1_HVT DP_OP_424J2_126_3477_U731 ( .A(DP_OP_424J2_126_3477_n1189), .B(
        DP_OP_424J2_126_3477_n1169), .CI(DP_OP_424J2_126_3477_n1330), .CO(
        DP_OP_424J2_126_3477_n1098), .S(DP_OP_424J2_126_3477_n1099) );
  FADDX1_HVT DP_OP_424J2_126_3477_U730 ( .A(DP_OP_424J2_126_3477_n1328), .B(
        DP_OP_424J2_126_3477_n1326), .CI(DP_OP_424J2_126_3477_n1324), .CO(
        DP_OP_424J2_126_3477_n1096), .S(DP_OP_424J2_126_3477_n1097) );
  FADDX1_HVT DP_OP_424J2_126_3477_U729 ( .A(DP_OP_424J2_126_3477_n1322), .B(
        DP_OP_424J2_126_3477_n1310), .CI(DP_OP_424J2_126_3477_n1308), .CO(
        DP_OP_424J2_126_3477_n1094), .S(DP_OP_424J2_126_3477_n1095) );
  FADDX1_HVT DP_OP_424J2_126_3477_U728 ( .A(DP_OP_424J2_126_3477_n1314), .B(
        DP_OP_424J2_126_3477_n1312), .CI(DP_OP_424J2_126_3477_n1320), .CO(
        DP_OP_424J2_126_3477_n1092), .S(DP_OP_424J2_126_3477_n1093) );
  FADDX1_HVT DP_OP_424J2_126_3477_U727 ( .A(DP_OP_424J2_126_3477_n1143), .B(
        DP_OP_424J2_126_3477_n1318), .CI(DP_OP_424J2_126_3477_n1316), .CO(
        DP_OP_424J2_126_3477_n1090), .S(DP_OP_424J2_126_3477_n1091) );
  FADDX1_HVT DP_OP_424J2_126_3477_U726 ( .A(DP_OP_424J2_126_3477_n1306), .B(
        DP_OP_424J2_126_3477_n1304), .CI(DP_OP_424J2_126_3477_n1137), .CO(
        DP_OP_424J2_126_3477_n1088), .S(DP_OP_424J2_126_3477_n1089) );
  FADDX1_HVT DP_OP_424J2_126_3477_U725 ( .A(DP_OP_424J2_126_3477_n1141), .B(
        DP_OP_424J2_126_3477_n1139), .CI(DP_OP_424J2_126_3477_n1302), .CO(
        DP_OP_424J2_126_3477_n1086), .S(DP_OP_424J2_126_3477_n1087) );
  FADDX1_HVT DP_OP_424J2_126_3477_U724 ( .A(DP_OP_424J2_126_3477_n1290), .B(
        DP_OP_424J2_126_3477_n1135), .CI(DP_OP_424J2_126_3477_n1121), .CO(
        DP_OP_424J2_126_3477_n1084), .S(DP_OP_424J2_126_3477_n1085) );
  FADDX1_HVT DP_OP_424J2_126_3477_U723 ( .A(DP_OP_424J2_126_3477_n1288), .B(
        DP_OP_424J2_126_3477_n1131), .CI(DP_OP_424J2_126_3477_n1133), .CO(
        DP_OP_424J2_126_3477_n1082), .S(DP_OP_424J2_126_3477_n1083) );
  FADDX1_HVT DP_OP_424J2_126_3477_U722 ( .A(DP_OP_424J2_126_3477_n1292), .B(
        DP_OP_424J2_126_3477_n1129), .CI(DP_OP_424J2_126_3477_n1127), .CO(
        DP_OP_424J2_126_3477_n1080), .S(DP_OP_424J2_126_3477_n1081) );
  FADDX1_HVT DP_OP_424J2_126_3477_U721 ( .A(DP_OP_424J2_126_3477_n1300), .B(
        DP_OP_424J2_126_3477_n1123), .CI(DP_OP_424J2_126_3477_n1125), .CO(
        DP_OP_424J2_126_3477_n1078), .S(DP_OP_424J2_126_3477_n1079) );
  FADDX1_HVT DP_OP_424J2_126_3477_U720 ( .A(DP_OP_424J2_126_3477_n1298), .B(
        DP_OP_424J2_126_3477_n1294), .CI(DP_OP_424J2_126_3477_n1296), .CO(
        DP_OP_424J2_126_3477_n1076), .S(DP_OP_424J2_126_3477_n1077) );
  FADDX1_HVT DP_OP_424J2_126_3477_U719 ( .A(DP_OP_424J2_126_3477_n1117), .B(
        DP_OP_424J2_126_3477_n1286), .CI(DP_OP_424J2_126_3477_n1115), .CO(
        DP_OP_424J2_126_3477_n1074), .S(DP_OP_424J2_126_3477_n1075) );
  FADDX1_HVT DP_OP_424J2_126_3477_U718 ( .A(DP_OP_424J2_126_3477_n1119), .B(
        DP_OP_424J2_126_3477_n1109), .CI(DP_OP_424J2_126_3477_n1111), .CO(
        DP_OP_424J2_126_3477_n1072), .S(DP_OP_424J2_126_3477_n1073) );
  FADDX1_HVT DP_OP_424J2_126_3477_U717 ( .A(DP_OP_424J2_126_3477_n1107), .B(
        DP_OP_424J2_126_3477_n1101), .CI(DP_OP_424J2_126_3477_n1284), .CO(
        DP_OP_424J2_126_3477_n1070), .S(DP_OP_424J2_126_3477_n1071) );
  FADDX1_HVT DP_OP_424J2_126_3477_U716 ( .A(DP_OP_424J2_126_3477_n1103), .B(
        DP_OP_424J2_126_3477_n1113), .CI(DP_OP_424J2_126_3477_n1105), .CO(
        DP_OP_424J2_126_3477_n1068), .S(DP_OP_424J2_126_3477_n1069) );
  FADDX1_HVT DP_OP_424J2_126_3477_U715 ( .A(DP_OP_424J2_126_3477_n1099), .B(
        DP_OP_424J2_126_3477_n1282), .CI(DP_OP_424J2_126_3477_n1278), .CO(
        DP_OP_424J2_126_3477_n1066), .S(DP_OP_424J2_126_3477_n1067) );
  FADDX1_HVT DP_OP_424J2_126_3477_U714 ( .A(DP_OP_424J2_126_3477_n1280), .B(
        DP_OP_424J2_126_3477_n1276), .CI(DP_OP_424J2_126_3477_n1274), .CO(
        DP_OP_424J2_126_3477_n1064), .S(DP_OP_424J2_126_3477_n1065) );
  FADDX1_HVT DP_OP_424J2_126_3477_U713 ( .A(DP_OP_424J2_126_3477_n1097), .B(
        DP_OP_424J2_126_3477_n1272), .CI(DP_OP_424J2_126_3477_n1270), .CO(
        DP_OP_424J2_126_3477_n1062), .S(DP_OP_424J2_126_3477_n1063) );
  FADDX1_HVT DP_OP_424J2_126_3477_U712 ( .A(DP_OP_424J2_126_3477_n1268), .B(
        DP_OP_424J2_126_3477_n1093), .CI(DP_OP_424J2_126_3477_n1091), .CO(
        DP_OP_424J2_126_3477_n1060), .S(DP_OP_424J2_126_3477_n1061) );
  FADDX1_HVT DP_OP_424J2_126_3477_U711 ( .A(DP_OP_424J2_126_3477_n1266), .B(
        DP_OP_424J2_126_3477_n1264), .CI(DP_OP_424J2_126_3477_n1095), .CO(
        DP_OP_424J2_126_3477_n1058), .S(DP_OP_424J2_126_3477_n1059) );
  FADDX1_HVT DP_OP_424J2_126_3477_U710 ( .A(DP_OP_424J2_126_3477_n1087), .B(
        DP_OP_424J2_126_3477_n1262), .CI(DP_OP_424J2_126_3477_n1089), .CO(
        DP_OP_424J2_126_3477_n1056), .S(DP_OP_424J2_126_3477_n1057) );
  FADDX1_HVT DP_OP_424J2_126_3477_U709 ( .A(DP_OP_424J2_126_3477_n1081), .B(
        DP_OP_424J2_126_3477_n1085), .CI(DP_OP_424J2_126_3477_n1256), .CO(
        DP_OP_424J2_126_3477_n1054), .S(DP_OP_424J2_126_3477_n1055) );
  FADDX1_HVT DP_OP_424J2_126_3477_U708 ( .A(DP_OP_424J2_126_3477_n1083), .B(
        DP_OP_424J2_126_3477_n1079), .CI(DP_OP_424J2_126_3477_n1260), .CO(
        DP_OP_424J2_126_3477_n1052), .S(DP_OP_424J2_126_3477_n1053) );
  FADDX1_HVT DP_OP_424J2_126_3477_U707 ( .A(DP_OP_424J2_126_3477_n1258), .B(
        DP_OP_424J2_126_3477_n1077), .CI(DP_OP_424J2_126_3477_n1254), .CO(
        DP_OP_424J2_126_3477_n1050), .S(DP_OP_424J2_126_3477_n1051) );
  FADDX1_HVT DP_OP_424J2_126_3477_U706 ( .A(DP_OP_424J2_126_3477_n1075), .B(
        DP_OP_424J2_126_3477_n1073), .CI(DP_OP_424J2_126_3477_n1071), .CO(
        DP_OP_424J2_126_3477_n1048), .S(DP_OP_424J2_126_3477_n1049) );
  FADDX1_HVT DP_OP_424J2_126_3477_U705 ( .A(DP_OP_424J2_126_3477_n1069), .B(
        DP_OP_424J2_126_3477_n1252), .CI(DP_OP_424J2_126_3477_n1067), .CO(
        DP_OP_424J2_126_3477_n1046), .S(DP_OP_424J2_126_3477_n1047) );
  FADDX1_HVT DP_OP_424J2_126_3477_U704 ( .A(DP_OP_424J2_126_3477_n1250), .B(
        DP_OP_424J2_126_3477_n1248), .CI(DP_OP_424J2_126_3477_n1246), .CO(
        DP_OP_424J2_126_3477_n1044), .S(DP_OP_424J2_126_3477_n1045) );
  FADDX1_HVT DP_OP_424J2_126_3477_U703 ( .A(DP_OP_424J2_126_3477_n1065), .B(
        DP_OP_424J2_126_3477_n1244), .CI(DP_OP_424J2_126_3477_n1063), .CO(
        DP_OP_424J2_126_3477_n1042), .S(DP_OP_424J2_126_3477_n1043) );
  FADDX1_HVT DP_OP_424J2_126_3477_U702 ( .A(DP_OP_424J2_126_3477_n1059), .B(
        DP_OP_424J2_126_3477_n1242), .CI(DP_OP_424J2_126_3477_n1061), .CO(
        DP_OP_424J2_126_3477_n1040), .S(DP_OP_424J2_126_3477_n1041) );
  FADDX1_HVT DP_OP_424J2_126_3477_U701 ( .A(DP_OP_424J2_126_3477_n1240), .B(
        DP_OP_424J2_126_3477_n1238), .CI(DP_OP_424J2_126_3477_n1057), .CO(
        DP_OP_424J2_126_3477_n1038), .S(DP_OP_424J2_126_3477_n1039) );
  FADDX1_HVT DP_OP_424J2_126_3477_U700 ( .A(DP_OP_424J2_126_3477_n1236), .B(
        DP_OP_424J2_126_3477_n1053), .CI(DP_OP_424J2_126_3477_n1051), .CO(
        DP_OP_424J2_126_3477_n1036), .S(DP_OP_424J2_126_3477_n1037) );
  FADDX1_HVT DP_OP_424J2_126_3477_U699 ( .A(DP_OP_424J2_126_3477_n1055), .B(
        DP_OP_424J2_126_3477_n1234), .CI(DP_OP_424J2_126_3477_n1049), .CO(
        DP_OP_424J2_126_3477_n1034), .S(DP_OP_424J2_126_3477_n1035) );
  FADDX1_HVT DP_OP_424J2_126_3477_U698 ( .A(DP_OP_424J2_126_3477_n1047), .B(
        DP_OP_424J2_126_3477_n1232), .CI(DP_OP_424J2_126_3477_n1230), .CO(
        DP_OP_424J2_126_3477_n1032), .S(DP_OP_424J2_126_3477_n1033) );
  FADDX1_HVT DP_OP_424J2_126_3477_U697 ( .A(DP_OP_424J2_126_3477_n1045), .B(
        DP_OP_424J2_126_3477_n1228), .CI(DP_OP_424J2_126_3477_n1043), .CO(
        DP_OP_424J2_126_3477_n1030), .S(DP_OP_424J2_126_3477_n1031) );
  FADDX1_HVT DP_OP_424J2_126_3477_U696 ( .A(DP_OP_424J2_126_3477_n1226), .B(
        DP_OP_424J2_126_3477_n1041), .CI(DP_OP_424J2_126_3477_n1039), .CO(
        DP_OP_424J2_126_3477_n1028), .S(DP_OP_424J2_126_3477_n1029) );
  FADDX1_HVT DP_OP_424J2_126_3477_U695 ( .A(DP_OP_424J2_126_3477_n1224), .B(
        DP_OP_424J2_126_3477_n1037), .CI(DP_OP_424J2_126_3477_n1222), .CO(
        DP_OP_424J2_126_3477_n1026), .S(DP_OP_424J2_126_3477_n1027) );
  FADDX1_HVT DP_OP_424J2_126_3477_U694 ( .A(DP_OP_424J2_126_3477_n1035), .B(
        DP_OP_424J2_126_3477_n1220), .CI(DP_OP_424J2_126_3477_n1033), .CO(
        DP_OP_424J2_126_3477_n1024), .S(DP_OP_424J2_126_3477_n1025) );
  FADDX1_HVT DP_OP_424J2_126_3477_U692 ( .A(DP_OP_424J2_126_3477_n1216), .B(
        DP_OP_424J2_126_3477_n1027), .CI(DP_OP_424J2_126_3477_n1025), .CO(
        DP_OP_424J2_126_3477_n1020), .S(DP_OP_424J2_126_3477_n1021) );
  FADDX1_HVT DP_OP_424J2_126_3477_U691 ( .A(DP_OP_424J2_126_3477_n1214), .B(
        DP_OP_424J2_126_3477_n1023), .CI(DP_OP_424J2_126_3477_n1212), .CO(
        DP_OP_424J2_126_3477_n1018), .S(DP_OP_424J2_126_3477_n1019) );
  FADDX1_HVT DP_OP_424J2_126_3477_U690 ( .A(DP_OP_424J2_126_3477_n3028), .B(
        DP_OP_424J2_126_3477_n1973), .CI(DP_OP_424J2_126_3477_n1929), .CO(
        DP_OP_424J2_126_3477_n1016), .S(DP_OP_424J2_126_3477_n1017) );
  FADDX1_HVT DP_OP_424J2_126_3477_U689 ( .A(DP_OP_424J2_126_3477_n2853), .B(
        DP_OP_424J2_126_3477_n2170), .CI(DP_OP_424J2_126_3477_n2434), .CO(
        DP_OP_424J2_126_3477_n1014), .S(DP_OP_424J2_126_3477_n1015) );
  FADDX1_HVT DP_OP_424J2_126_3477_U688 ( .A(DP_OP_424J2_126_3477_n2061), .B(
        DP_OP_424J2_126_3477_n2478), .CI(DP_OP_424J2_126_3477_n2038), .CO(
        DP_OP_424J2_126_3477_n1012), .S(DP_OP_424J2_126_3477_n1013) );
  FADDX1_HVT DP_OP_424J2_126_3477_U687 ( .A(DP_OP_424J2_126_3477_n2369), .B(
        DP_OP_424J2_126_3477_n1994), .CI(DP_OP_424J2_126_3477_n2962), .CO(
        DP_OP_424J2_126_3477_n1010), .S(DP_OP_424J2_126_3477_n1011) );
  FADDX1_HVT DP_OP_424J2_126_3477_U686 ( .A(DP_OP_424J2_126_3477_n2325), .B(
        DP_OP_424J2_126_3477_n2302), .CI(DP_OP_424J2_126_3477_n2654), .CO(
        DP_OP_424J2_126_3477_n1008), .S(DP_OP_424J2_126_3477_n1009) );
  FADDX1_HVT DP_OP_424J2_126_3477_U685 ( .A(DP_OP_424J2_126_3477_n2237), .B(
        DP_OP_424J2_126_3477_n2346), .CI(DP_OP_424J2_126_3477_n3006), .CO(
        DP_OP_424J2_126_3477_n1006), .S(DP_OP_424J2_126_3477_n1007) );
  FADDX1_HVT DP_OP_424J2_126_3477_U684 ( .A(DP_OP_424J2_126_3477_n2017), .B(
        DP_OP_424J2_126_3477_n2082), .CI(DP_OP_424J2_126_3477_n2522), .CO(
        DP_OP_424J2_126_3477_n1004), .S(DP_OP_424J2_126_3477_n1005) );
  FADDX1_HVT DP_OP_424J2_126_3477_U683 ( .A(DP_OP_424J2_126_3477_n2105), .B(
        DP_OP_424J2_126_3477_n2786), .CI(DP_OP_424J2_126_3477_n2830), .CO(
        DP_OP_424J2_126_3477_n1002), .S(DP_OP_424J2_126_3477_n1003) );
  FADDX1_HVT DP_OP_424J2_126_3477_U682 ( .A(DP_OP_424J2_126_3477_n2193), .B(
        DP_OP_424J2_126_3477_n2742), .CI(DP_OP_424J2_126_3477_n2610), .CO(
        DP_OP_424J2_126_3477_n1000), .S(DP_OP_424J2_126_3477_n1001) );
  FADDX1_HVT DP_OP_424J2_126_3477_U681 ( .A(DP_OP_424J2_126_3477_n2545), .B(
        DP_OP_424J2_126_3477_n2390), .CI(DP_OP_424J2_126_3477_n2874), .CO(
        DP_OP_424J2_126_3477_n998), .S(DP_OP_424J2_126_3477_n999) );
  FADDX1_HVT DP_OP_424J2_126_3477_U680 ( .A(DP_OP_424J2_126_3477_n2941), .B(
        DP_OP_424J2_126_3477_n2214), .CI(DP_OP_424J2_126_3477_n2126), .CO(
        DP_OP_424J2_126_3477_n996), .S(DP_OP_424J2_126_3477_n997) );
  FADDX1_HVT DP_OP_424J2_126_3477_U679 ( .A(DP_OP_424J2_126_3477_n2677), .B(
        DP_OP_424J2_126_3477_n2918), .CI(DP_OP_424J2_126_3477_n2566), .CO(
        DP_OP_424J2_126_3477_n994), .S(DP_OP_424J2_126_3477_n995) );
  FADDX1_HVT DP_OP_424J2_126_3477_U678 ( .A(DP_OP_424J2_126_3477_n2457), .B(
        DP_OP_424J2_126_3477_n3048), .CI(DP_OP_424J2_126_3477_n2258), .CO(
        DP_OP_424J2_126_3477_n992), .S(DP_OP_424J2_126_3477_n993) );
  FADDX1_HVT DP_OP_424J2_126_3477_U677 ( .A(DP_OP_424J2_126_3477_n2149), .B(
        DP_OP_424J2_126_3477_n2413), .CI(DP_OP_424J2_126_3477_n2698), .CO(
        DP_OP_424J2_126_3477_n990), .S(DP_OP_424J2_126_3477_n991) );
  FADDX1_HVT DP_OP_424J2_126_3477_U676 ( .A(DP_OP_424J2_126_3477_n2765), .B(
        DP_OP_424J2_126_3477_n2809), .CI(DP_OP_424J2_126_3477_n2897), .CO(
        DP_OP_424J2_126_3477_n988), .S(DP_OP_424J2_126_3477_n989) );
  FADDX1_HVT DP_OP_424J2_126_3477_U675 ( .A(DP_OP_424J2_126_3477_n2501), .B(
        DP_OP_424J2_126_3477_n2589), .CI(DP_OP_424J2_126_3477_n2985), .CO(
        DP_OP_424J2_126_3477_n986), .S(DP_OP_424J2_126_3477_n987) );
  FADDX1_HVT DP_OP_424J2_126_3477_U674 ( .A(DP_OP_424J2_126_3477_n2633), .B(
        DP_OP_424J2_126_3477_n2281), .CI(DP_OP_424J2_126_3477_n2721), .CO(
        DP_OP_424J2_126_3477_n984), .S(DP_OP_424J2_126_3477_n985) );
  FADDX1_HVT DP_OP_424J2_126_3477_U673 ( .A(DP_OP_424J2_126_3477_n3041), .B(
        DP_OP_424J2_126_3477_n1987), .CI(DP_OP_424J2_126_3477_n1980), .CO(
        DP_OP_424J2_126_3477_n982), .S(DP_OP_424J2_126_3477_n983) );
  FADDX1_HVT DP_OP_424J2_126_3477_U672 ( .A(DP_OP_424J2_126_3477_n3034), .B(
        DP_OP_424J2_126_3477_n2999), .CI(DP_OP_424J2_126_3477_n2992), .CO(
        DP_OP_424J2_126_3477_n980), .S(DP_OP_424J2_126_3477_n981) );
  FADDX1_HVT DP_OP_424J2_126_3477_U671 ( .A(DP_OP_424J2_126_3477_n2515), .B(
        DP_OP_424J2_126_3477_n2955), .CI(DP_OP_424J2_126_3477_n2948), .CO(
        DP_OP_424J2_126_3477_n978), .S(DP_OP_424J2_126_3477_n979) );
  FADDX1_HVT DP_OP_424J2_126_3477_U670 ( .A(DP_OP_424J2_126_3477_n2911), .B(
        DP_OP_424J2_126_3477_n2024), .CI(DP_OP_424J2_126_3477_n2031), .CO(
        DP_OP_424J2_126_3477_n976), .S(DP_OP_424J2_126_3477_n977) );
  FADDX1_HVT DP_OP_424J2_126_3477_U669 ( .A(DP_OP_424J2_126_3477_n2904), .B(
        DP_OP_424J2_126_3477_n2068), .CI(DP_OP_424J2_126_3477_n2075), .CO(
        DP_OP_424J2_126_3477_n974), .S(DP_OP_424J2_126_3477_n975) );
  FADDX1_HVT DP_OP_424J2_126_3477_U668 ( .A(DP_OP_424J2_126_3477_n2867), .B(
        DP_OP_424J2_126_3477_n2112), .CI(DP_OP_424J2_126_3477_n2119), .CO(
        DP_OP_424J2_126_3477_n972), .S(DP_OP_424J2_126_3477_n973) );
  FADDX1_HVT DP_OP_424J2_126_3477_U667 ( .A(DP_OP_424J2_126_3477_n2860), .B(
        DP_OP_424J2_126_3477_n2156), .CI(DP_OP_424J2_126_3477_n2163), .CO(
        DP_OP_424J2_126_3477_n970), .S(DP_OP_424J2_126_3477_n971) );
  FADDX1_HVT DP_OP_424J2_126_3477_U666 ( .A(DP_OP_424J2_126_3477_n2823), .B(
        DP_OP_424J2_126_3477_n2200), .CI(DP_OP_424J2_126_3477_n2207), .CO(
        DP_OP_424J2_126_3477_n968), .S(DP_OP_424J2_126_3477_n969) );
  FADDX1_HVT DP_OP_424J2_126_3477_U665 ( .A(DP_OP_424J2_126_3477_n2816), .B(
        DP_OP_424J2_126_3477_n2244), .CI(DP_OP_424J2_126_3477_n2251), .CO(
        DP_OP_424J2_126_3477_n966), .S(DP_OP_424J2_126_3477_n967) );
  FADDX1_HVT DP_OP_424J2_126_3477_U664 ( .A(DP_OP_424J2_126_3477_n2779), .B(
        DP_OP_424J2_126_3477_n2288), .CI(DP_OP_424J2_126_3477_n2295), .CO(
        DP_OP_424J2_126_3477_n964), .S(DP_OP_424J2_126_3477_n965) );
  FADDX1_HVT DP_OP_424J2_126_3477_U663 ( .A(DP_OP_424J2_126_3477_n2772), .B(
        DP_OP_424J2_126_3477_n2332), .CI(DP_OP_424J2_126_3477_n2339), .CO(
        DP_OP_424J2_126_3477_n962), .S(DP_OP_424J2_126_3477_n963) );
  FADDX1_HVT DP_OP_424J2_126_3477_U662 ( .A(DP_OP_424J2_126_3477_n2735), .B(
        DP_OP_424J2_126_3477_n2376), .CI(DP_OP_424J2_126_3477_n2383), .CO(
        DP_OP_424J2_126_3477_n960), .S(DP_OP_424J2_126_3477_n961) );
  FADDX1_HVT DP_OP_424J2_126_3477_U661 ( .A(DP_OP_424J2_126_3477_n2728), .B(
        DP_OP_424J2_126_3477_n2420), .CI(DP_OP_424J2_126_3477_n2427), .CO(
        DP_OP_424J2_126_3477_n958), .S(DP_OP_424J2_126_3477_n959) );
  FADDX1_HVT DP_OP_424J2_126_3477_U660 ( .A(DP_OP_424J2_126_3477_n2691), .B(
        DP_OP_424J2_126_3477_n2464), .CI(DP_OP_424J2_126_3477_n2471), .CO(
        DP_OP_424J2_126_3477_n956), .S(DP_OP_424J2_126_3477_n957) );
  FADDX1_HVT DP_OP_424J2_126_3477_U659 ( .A(DP_OP_424J2_126_3477_n2684), .B(
        DP_OP_424J2_126_3477_n2508), .CI(DP_OP_424J2_126_3477_n2552), .CO(
        DP_OP_424J2_126_3477_n954), .S(DP_OP_424J2_126_3477_n955) );
  FADDX1_HVT DP_OP_424J2_126_3477_U658 ( .A(DP_OP_424J2_126_3477_n2647), .B(
        DP_OP_424J2_126_3477_n2559), .CI(DP_OP_424J2_126_3477_n2596), .CO(
        DP_OP_424J2_126_3477_n952), .S(DP_OP_424J2_126_3477_n953) );
  FADDX1_HVT DP_OP_424J2_126_3477_U657 ( .A(DP_OP_424J2_126_3477_n2640), .B(
        DP_OP_424J2_126_3477_n2603), .CI(DP_OP_424J2_126_3477_n1210), .CO(
        DP_OP_424J2_126_3477_n950), .S(DP_OP_424J2_126_3477_n951) );
  FADDX1_HVT DP_OP_424J2_126_3477_U656 ( .A(DP_OP_424J2_126_3477_n1198), .B(
        DP_OP_424J2_126_3477_n1194), .CI(DP_OP_424J2_126_3477_n1208), .CO(
        DP_OP_424J2_126_3477_n948), .S(DP_OP_424J2_126_3477_n949) );
  FADDX1_HVT DP_OP_424J2_126_3477_U655 ( .A(DP_OP_424J2_126_3477_n1206), .B(
        DP_OP_424J2_126_3477_n1196), .CI(DP_OP_424J2_126_3477_n1204), .CO(
        DP_OP_424J2_126_3477_n946), .S(DP_OP_424J2_126_3477_n947) );
  FADDX1_HVT DP_OP_424J2_126_3477_U654 ( .A(DP_OP_424J2_126_3477_n1202), .B(
        DP_OP_424J2_126_3477_n1200), .CI(DP_OP_424J2_126_3477_n1170), .CO(
        DP_OP_424J2_126_3477_n944), .S(DP_OP_424J2_126_3477_n945) );
  FADDX1_HVT DP_OP_424J2_126_3477_U653 ( .A(DP_OP_424J2_126_3477_n1168), .B(
        DP_OP_424J2_126_3477_n1144), .CI(DP_OP_424J2_126_3477_n1192), .CO(
        DP_OP_424J2_126_3477_n942), .S(DP_OP_424J2_126_3477_n943) );
  FADDX1_HVT DP_OP_424J2_126_3477_U652 ( .A(DP_OP_424J2_126_3477_n1166), .B(
        DP_OP_424J2_126_3477_n1190), .CI(DP_OP_424J2_126_3477_n1188), .CO(
        DP_OP_424J2_126_3477_n940), .S(DP_OP_424J2_126_3477_n941) );
  FADDX1_HVT DP_OP_424J2_126_3477_U651 ( .A(DP_OP_424J2_126_3477_n1160), .B(
        DP_OP_424J2_126_3477_n1186), .CI(DP_OP_424J2_126_3477_n1184), .CO(
        DP_OP_424J2_126_3477_n938), .S(DP_OP_424J2_126_3477_n939) );
  FADDX1_HVT DP_OP_424J2_126_3477_U650 ( .A(DP_OP_424J2_126_3477_n1182), .B(
        DP_OP_424J2_126_3477_n1180), .CI(DP_OP_424J2_126_3477_n1178), .CO(
        DP_OP_424J2_126_3477_n936), .S(DP_OP_424J2_126_3477_n937) );
  FADDX1_HVT DP_OP_424J2_126_3477_U649 ( .A(DP_OP_424J2_126_3477_n1150), .B(
        DP_OP_424J2_126_3477_n1176), .CI(DP_OP_424J2_126_3477_n1174), .CO(
        DP_OP_424J2_126_3477_n934), .S(DP_OP_424J2_126_3477_n935) );
  FADDX1_HVT DP_OP_424J2_126_3477_U648 ( .A(DP_OP_424J2_126_3477_n1156), .B(
        DP_OP_424J2_126_3477_n1172), .CI(DP_OP_424J2_126_3477_n1164), .CO(
        DP_OP_424J2_126_3477_n932), .S(DP_OP_424J2_126_3477_n933) );
  FADDX1_HVT DP_OP_424J2_126_3477_U647 ( .A(DP_OP_424J2_126_3477_n1148), .B(
        DP_OP_424J2_126_3477_n1162), .CI(DP_OP_424J2_126_3477_n1158), .CO(
        DP_OP_424J2_126_3477_n930), .S(DP_OP_424J2_126_3477_n931) );
  FADDX1_HVT DP_OP_424J2_126_3477_U646 ( .A(DP_OP_424J2_126_3477_n1152), .B(
        DP_OP_424J2_126_3477_n1146), .CI(DP_OP_424J2_126_3477_n1154), .CO(
        DP_OP_424J2_126_3477_n928), .S(DP_OP_424J2_126_3477_n929) );
  FADDX1_HVT DP_OP_424J2_126_3477_U645 ( .A(DP_OP_424J2_126_3477_n1017), .B(
        DP_OP_424J2_126_3477_n1003), .CI(DP_OP_424J2_126_3477_n1005), .CO(
        DP_OP_424J2_126_3477_n926), .S(DP_OP_424J2_126_3477_n927) );
  FADDX1_HVT DP_OP_424J2_126_3477_U644 ( .A(DP_OP_424J2_126_3477_n1009), .B(
        DP_OP_424J2_126_3477_n987), .CI(DP_OP_424J2_126_3477_n985), .CO(
        DP_OP_424J2_126_3477_n924), .S(DP_OP_424J2_126_3477_n925) );
  FADDX1_HVT DP_OP_424J2_126_3477_U643 ( .A(DP_OP_424J2_126_3477_n1001), .B(
        DP_OP_424J2_126_3477_n999), .CI(DP_OP_424J2_126_3477_n995), .CO(
        DP_OP_424J2_126_3477_n922), .S(DP_OP_424J2_126_3477_n923) );
  FADDX1_HVT DP_OP_424J2_126_3477_U642 ( .A(DP_OP_424J2_126_3477_n1007), .B(
        DP_OP_424J2_126_3477_n989), .CI(DP_OP_424J2_126_3477_n993), .CO(
        DP_OP_424J2_126_3477_n920), .S(DP_OP_424J2_126_3477_n921) );
  FADDX1_HVT DP_OP_424J2_126_3477_U641 ( .A(DP_OP_424J2_126_3477_n997), .B(
        DP_OP_424J2_126_3477_n1015), .CI(DP_OP_424J2_126_3477_n1011), .CO(
        DP_OP_424J2_126_3477_n918), .S(DP_OP_424J2_126_3477_n919) );
  FADDX1_HVT DP_OP_424J2_126_3477_U640 ( .A(DP_OP_424J2_126_3477_n991), .B(
        DP_OP_424J2_126_3477_n1013), .CI(DP_OP_424J2_126_3477_n973), .CO(
        DP_OP_424J2_126_3477_n916), .S(DP_OP_424J2_126_3477_n917) );
  FADDX1_HVT DP_OP_424J2_126_3477_U639 ( .A(DP_OP_424J2_126_3477_n975), .B(
        DP_OP_424J2_126_3477_n957), .CI(DP_OP_424J2_126_3477_n951), .CO(
        DP_OP_424J2_126_3477_n914), .S(DP_OP_424J2_126_3477_n915) );
  FADDX1_HVT DP_OP_424J2_126_3477_U638 ( .A(DP_OP_424J2_126_3477_n977), .B(
        DP_OP_424J2_126_3477_n953), .CI(DP_OP_424J2_126_3477_n969), .CO(
        DP_OP_424J2_126_3477_n912), .S(DP_OP_424J2_126_3477_n913) );
  FADDX1_HVT DP_OP_424J2_126_3477_U637 ( .A(DP_OP_424J2_126_3477_n967), .B(
        DP_OP_424J2_126_3477_n965), .CI(DP_OP_424J2_126_3477_n955), .CO(
        DP_OP_424J2_126_3477_n910), .S(DP_OP_424J2_126_3477_n911) );
  FADDX1_HVT DP_OP_424J2_126_3477_U636 ( .A(DP_OP_424J2_126_3477_n971), .B(
        DP_OP_424J2_126_3477_n959), .CI(DP_OP_424J2_126_3477_n961), .CO(
        DP_OP_424J2_126_3477_n908), .S(DP_OP_424J2_126_3477_n909) );
  FADDX1_HVT DP_OP_424J2_126_3477_U635 ( .A(DP_OP_424J2_126_3477_n979), .B(
        DP_OP_424J2_126_3477_n981), .CI(DP_OP_424J2_126_3477_n983), .CO(
        DP_OP_424J2_126_3477_n906), .S(DP_OP_424J2_126_3477_n907) );
  FADDX1_HVT DP_OP_424J2_126_3477_U634 ( .A(DP_OP_424J2_126_3477_n963), .B(
        DP_OP_424J2_126_3477_n1142), .CI(DP_OP_424J2_126_3477_n1140), .CO(
        DP_OP_424J2_126_3477_n904), .S(DP_OP_424J2_126_3477_n905) );
  FADDX1_HVT DP_OP_424J2_126_3477_U633 ( .A(DP_OP_424J2_126_3477_n1138), .B(
        DP_OP_424J2_126_3477_n1136), .CI(DP_OP_424J2_126_3477_n1122), .CO(
        DP_OP_424J2_126_3477_n902), .S(DP_OP_424J2_126_3477_n903) );
  FADDX1_HVT DP_OP_424J2_126_3477_U632 ( .A(DP_OP_424J2_126_3477_n1134), .B(
        DP_OP_424J2_126_3477_n1132), .CI(DP_OP_424J2_126_3477_n1120), .CO(
        DP_OP_424J2_126_3477_n900), .S(DP_OP_424J2_126_3477_n901) );
  FADDX1_HVT DP_OP_424J2_126_3477_U631 ( .A(DP_OP_424J2_126_3477_n1130), .B(
        DP_OP_424J2_126_3477_n1124), .CI(DP_OP_424J2_126_3477_n1126), .CO(
        DP_OP_424J2_126_3477_n898), .S(DP_OP_424J2_126_3477_n899) );
  FADDX1_HVT DP_OP_424J2_126_3477_U630 ( .A(DP_OP_424J2_126_3477_n1128), .B(
        DP_OP_424J2_126_3477_n1118), .CI(DP_OP_424J2_126_3477_n1116), .CO(
        DP_OP_424J2_126_3477_n896), .S(DP_OP_424J2_126_3477_n897) );
  FADDX1_HVT DP_OP_424J2_126_3477_U629 ( .A(DP_OP_424J2_126_3477_n949), .B(
        DP_OP_424J2_126_3477_n945), .CI(DP_OP_424J2_126_3477_n1114), .CO(
        DP_OP_424J2_126_3477_n894), .S(DP_OP_424J2_126_3477_n895) );
  FADDX1_HVT DP_OP_424J2_126_3477_U628 ( .A(DP_OP_424J2_126_3477_n947), .B(
        DP_OP_424J2_126_3477_n1102), .CI(DP_OP_424J2_126_3477_n1100), .CO(
        DP_OP_424J2_126_3477_n892), .S(DP_OP_424J2_126_3477_n893) );
  FADDX1_HVT DP_OP_424J2_126_3477_U627 ( .A(DP_OP_424J2_126_3477_n1108), .B(
        DP_OP_424J2_126_3477_n943), .CI(DP_OP_424J2_126_3477_n1098), .CO(
        DP_OP_424J2_126_3477_n890), .S(DP_OP_424J2_126_3477_n891) );
  FADDX1_HVT DP_OP_424J2_126_3477_U626 ( .A(DP_OP_424J2_126_3477_n1106), .B(
        DP_OP_424J2_126_3477_n939), .CI(DP_OP_424J2_126_3477_n929), .CO(
        DP_OP_424J2_126_3477_n888), .S(DP_OP_424J2_126_3477_n889) );
  FADDX1_HVT DP_OP_424J2_126_3477_U625 ( .A(DP_OP_424J2_126_3477_n1112), .B(
        DP_OP_424J2_126_3477_n935), .CI(DP_OP_424J2_126_3477_n937), .CO(
        DP_OP_424J2_126_3477_n886), .S(DP_OP_424J2_126_3477_n887) );
  FADDX1_HVT DP_OP_424J2_126_3477_U624 ( .A(DP_OP_424J2_126_3477_n1110), .B(
        DP_OP_424J2_126_3477_n931), .CI(DP_OP_424J2_126_3477_n933), .CO(
        DP_OP_424J2_126_3477_n884), .S(DP_OP_424J2_126_3477_n885) );
  FADDX1_HVT DP_OP_424J2_126_3477_U623 ( .A(DP_OP_424J2_126_3477_n1104), .B(
        DP_OP_424J2_126_3477_n941), .CI(DP_OP_424J2_126_3477_n927), .CO(
        DP_OP_424J2_126_3477_n882), .S(DP_OP_424J2_126_3477_n883) );
  FADDX1_HVT DP_OP_424J2_126_3477_U622 ( .A(DP_OP_424J2_126_3477_n921), .B(
        DP_OP_424J2_126_3477_n925), .CI(DP_OP_424J2_126_3477_n917), .CO(
        DP_OP_424J2_126_3477_n880), .S(DP_OP_424J2_126_3477_n881) );
  FADDX1_HVT DP_OP_424J2_126_3477_U621 ( .A(DP_OP_424J2_126_3477_n919), .B(
        DP_OP_424J2_126_3477_n923), .CI(DP_OP_424J2_126_3477_n911), .CO(
        DP_OP_424J2_126_3477_n878), .S(DP_OP_424J2_126_3477_n879) );
  FADDX1_HVT DP_OP_424J2_126_3477_U620 ( .A(DP_OP_424J2_126_3477_n909), .B(
        DP_OP_424J2_126_3477_n915), .CI(DP_OP_424J2_126_3477_n1096), .CO(
        DP_OP_424J2_126_3477_n876), .S(DP_OP_424J2_126_3477_n877) );
  FADDX1_HVT DP_OP_424J2_126_3477_U619 ( .A(DP_OP_424J2_126_3477_n907), .B(
        DP_OP_424J2_126_3477_n913), .CI(DP_OP_424J2_126_3477_n1092), .CO(
        DP_OP_424J2_126_3477_n874), .S(DP_OP_424J2_126_3477_n875) );
  FADDX1_HVT DP_OP_424J2_126_3477_U618 ( .A(DP_OP_424J2_126_3477_n1090), .B(
        DP_OP_424J2_126_3477_n905), .CI(DP_OP_424J2_126_3477_n1094), .CO(
        DP_OP_424J2_126_3477_n872), .S(DP_OP_424J2_126_3477_n873) );
  FADDX1_HVT DP_OP_424J2_126_3477_U617 ( .A(DP_OP_424J2_126_3477_n1088), .B(
        DP_OP_424J2_126_3477_n1086), .CI(DP_OP_424J2_126_3477_n903), .CO(
        DP_OP_424J2_126_3477_n870), .S(DP_OP_424J2_126_3477_n871) );
  FADDX1_HVT DP_OP_424J2_126_3477_U616 ( .A(DP_OP_424J2_126_3477_n1084), .B(
        DP_OP_424J2_126_3477_n901), .CI(DP_OP_424J2_126_3477_n899), .CO(
        DP_OP_424J2_126_3477_n868), .S(DP_OP_424J2_126_3477_n869) );
  FADDX1_HVT DP_OP_424J2_126_3477_U615 ( .A(DP_OP_424J2_126_3477_n1082), .B(
        DP_OP_424J2_126_3477_n1076), .CI(DP_OP_424J2_126_3477_n1078), .CO(
        DP_OP_424J2_126_3477_n866), .S(DP_OP_424J2_126_3477_n867) );
  FADDX1_HVT DP_OP_424J2_126_3477_U614 ( .A(DP_OP_424J2_126_3477_n1080), .B(
        DP_OP_424J2_126_3477_n897), .CI(DP_OP_424J2_126_3477_n1074), .CO(
        DP_OP_424J2_126_3477_n864), .S(DP_OP_424J2_126_3477_n865) );
  FADDX1_HVT DP_OP_424J2_126_3477_U613 ( .A(DP_OP_424J2_126_3477_n895), .B(
        DP_OP_424J2_126_3477_n1072), .CI(DP_OP_424J2_126_3477_n893), .CO(
        DP_OP_424J2_126_3477_n862), .S(DP_OP_424J2_126_3477_n863) );
  FADDX1_HVT DP_OP_424J2_126_3477_U612 ( .A(DP_OP_424J2_126_3477_n1070), .B(
        DP_OP_424J2_126_3477_n887), .CI(DP_OP_424J2_126_3477_n883), .CO(
        DP_OP_424J2_126_3477_n860), .S(DP_OP_424J2_126_3477_n861) );
  FADDX1_HVT DP_OP_424J2_126_3477_U611 ( .A(DP_OP_424J2_126_3477_n1068), .B(
        DP_OP_424J2_126_3477_n891), .CI(DP_OP_424J2_126_3477_n889), .CO(
        DP_OP_424J2_126_3477_n858), .S(DP_OP_424J2_126_3477_n859) );
  FADDX1_HVT DP_OP_424J2_126_3477_U610 ( .A(DP_OP_424J2_126_3477_n885), .B(
        DP_OP_424J2_126_3477_n1066), .CI(DP_OP_424J2_126_3477_n881), .CO(
        DP_OP_424J2_126_3477_n856), .S(DP_OP_424J2_126_3477_n857) );
  FADDX1_HVT DP_OP_424J2_126_3477_U609 ( .A(DP_OP_424J2_126_3477_n879), .B(
        DP_OP_424J2_126_3477_n1064), .CI(DP_OP_424J2_126_3477_n877), .CO(
        DP_OP_424J2_126_3477_n854), .S(DP_OP_424J2_126_3477_n855) );
  FADDX1_HVT DP_OP_424J2_126_3477_U608 ( .A(DP_OP_424J2_126_3477_n875), .B(
        DP_OP_424J2_126_3477_n1062), .CI(DP_OP_424J2_126_3477_n1058), .CO(
        DP_OP_424J2_126_3477_n852), .S(DP_OP_424J2_126_3477_n853) );
  FADDX1_HVT DP_OP_424J2_126_3477_U607 ( .A(DP_OP_424J2_126_3477_n1060), .B(
        DP_OP_424J2_126_3477_n873), .CI(DP_OP_424J2_126_3477_n1056), .CO(
        DP_OP_424J2_126_3477_n850), .S(DP_OP_424J2_126_3477_n851) );
  FADDX1_HVT DP_OP_424J2_126_3477_U606 ( .A(DP_OP_424J2_126_3477_n871), .B(
        DP_OP_424J2_126_3477_n1054), .CI(DP_OP_424J2_126_3477_n1052), .CO(
        DP_OP_424J2_126_3477_n848), .S(DP_OP_424J2_126_3477_n849) );
  FADDX1_HVT DP_OP_424J2_126_3477_U605 ( .A(DP_OP_424J2_126_3477_n869), .B(
        DP_OP_424J2_126_3477_n1050), .CI(DP_OP_424J2_126_3477_n865), .CO(
        DP_OP_424J2_126_3477_n846), .S(DP_OP_424J2_126_3477_n847) );
  FADDX1_HVT DP_OP_424J2_126_3477_U604 ( .A(DP_OP_424J2_126_3477_n867), .B(
        DP_OP_424J2_126_3477_n1048), .CI(DP_OP_424J2_126_3477_n863), .CO(
        DP_OP_424J2_126_3477_n844), .S(DP_OP_424J2_126_3477_n845) );
  FADDX1_HVT DP_OP_424J2_126_3477_U603 ( .A(DP_OP_424J2_126_3477_n1046), .B(
        DP_OP_424J2_126_3477_n857), .CI(DP_OP_424J2_126_3477_n861), .CO(
        DP_OP_424J2_126_3477_n842), .S(DP_OP_424J2_126_3477_n843) );
  FADDX1_HVT DP_OP_424J2_126_3477_U602 ( .A(DP_OP_424J2_126_3477_n859), .B(
        DP_OP_424J2_126_3477_n1044), .CI(DP_OP_424J2_126_3477_n855), .CO(
        DP_OP_424J2_126_3477_n840), .S(DP_OP_424J2_126_3477_n841) );
  FADDX1_HVT DP_OP_424J2_126_3477_U601 ( .A(DP_OP_424J2_126_3477_n1042), .B(
        DP_OP_424J2_126_3477_n853), .CI(DP_OP_424J2_126_3477_n1040), .CO(
        DP_OP_424J2_126_3477_n838), .S(DP_OP_424J2_126_3477_n839) );
  FADDX1_HVT DP_OP_424J2_126_3477_U600 ( .A(DP_OP_424J2_126_3477_n851), .B(
        DP_OP_424J2_126_3477_n849), .CI(DP_OP_424J2_126_3477_n1038), .CO(
        DP_OP_424J2_126_3477_n836), .S(DP_OP_424J2_126_3477_n837) );
  FADDX1_HVT DP_OP_424J2_126_3477_U599 ( .A(DP_OP_424J2_126_3477_n1036), .B(
        DP_OP_424J2_126_3477_n847), .CI(DP_OP_424J2_126_3477_n1034), .CO(
        DP_OP_424J2_126_3477_n834), .S(DP_OP_424J2_126_3477_n835) );
  FADDX1_HVT DP_OP_424J2_126_3477_U598 ( .A(DP_OP_424J2_126_3477_n845), .B(
        DP_OP_424J2_126_3477_n843), .CI(DP_OP_424J2_126_3477_n1032), .CO(
        DP_OP_424J2_126_3477_n832), .S(DP_OP_424J2_126_3477_n833) );
  FADDX1_HVT DP_OP_424J2_126_3477_U597 ( .A(DP_OP_424J2_126_3477_n841), .B(
        DP_OP_424J2_126_3477_n1030), .CI(DP_OP_424J2_126_3477_n839), .CO(
        DP_OP_424J2_126_3477_n830), .S(DP_OP_424J2_126_3477_n831) );
  FADDX1_HVT DP_OP_424J2_126_3477_U596 ( .A(DP_OP_424J2_126_3477_n1028), .B(
        DP_OP_424J2_126_3477_n837), .CI(DP_OP_424J2_126_3477_n1026), .CO(
        DP_OP_424J2_126_3477_n828), .S(DP_OP_424J2_126_3477_n829) );
  FADDX1_HVT DP_OP_424J2_126_3477_U595 ( .A(DP_OP_424J2_126_3477_n835), .B(
        DP_OP_424J2_126_3477_n833), .CI(DP_OP_424J2_126_3477_n1024), .CO(
        DP_OP_424J2_126_3477_n826), .S(DP_OP_424J2_126_3477_n827) );
  FADDX1_HVT DP_OP_424J2_126_3477_U594 ( .A(DP_OP_424J2_126_3477_n831), .B(
        DP_OP_424J2_126_3477_n829), .CI(DP_OP_424J2_126_3477_n1022), .CO(
        DP_OP_424J2_126_3477_n824), .S(DP_OP_424J2_126_3477_n825) );
  FADDX1_HVT DP_OP_424J2_126_3477_U591 ( .A(DP_OP_424J2_126_3477_n2236), .B(
        DP_OP_424J2_126_3477_n1972), .CI(DP_OP_424J2_126_3477_n1928), .CO(
        DP_OP_424J2_126_3477_n818), .S(DP_OP_424J2_126_3477_n819) );
  FADDX1_HVT DP_OP_424J2_126_3477_U590 ( .A(DP_OP_424J2_126_3477_n2808), .B(
        DP_OP_424J2_126_3477_n2030), .CI(DP_OP_424J2_126_3477_n2294), .CO(
        DP_OP_424J2_126_3477_n816), .S(DP_OP_424J2_126_3477_n817) );
  FADDX1_HVT DP_OP_424J2_126_3477_U589 ( .A(DP_OP_424J2_126_3477_n2280), .B(
        DP_OP_424J2_126_3477_n3040), .CI(DP_OP_424J2_126_3477_n2690), .CO(
        DP_OP_424J2_126_3477_n814), .S(DP_OP_424J2_126_3477_n815) );
  FADDX1_HVT DP_OP_424J2_126_3477_U588 ( .A(DP_OP_424J2_126_3477_n2500), .B(
        DP_OP_424J2_126_3477_n2074), .CI(DP_OP_424J2_126_3477_n2118), .CO(
        DP_OP_424J2_126_3477_n812), .S(DP_OP_424J2_126_3477_n813) );
  FADDX1_HVT DP_OP_424J2_126_3477_U587 ( .A(DP_OP_424J2_126_3477_n2060), .B(
        DP_OP_424J2_126_3477_n2162), .CI(DP_OP_424J2_126_3477_n2206), .CO(
        DP_OP_424J2_126_3477_n810), .S(DP_OP_424J2_126_3477_n811) );
  FADDX1_HVT DP_OP_424J2_126_3477_U586 ( .A(DP_OP_424J2_126_3477_n2764), .B(
        DP_OP_424J2_126_3477_n2866), .CI(DP_OP_424J2_126_3477_n2910), .CO(
        DP_OP_424J2_126_3477_n808), .S(DP_OP_424J2_126_3477_n809) );
  FADDX1_HVT DP_OP_424J2_126_3477_U585 ( .A(DP_OP_424J2_126_3477_n2104), .B(
        DP_OP_424J2_126_3477_n2822), .CI(DP_OP_424J2_126_3477_n2646), .CO(
        DP_OP_424J2_126_3477_n806), .S(DP_OP_424J2_126_3477_n807) );
  FADDX1_HVT DP_OP_424J2_126_3477_U584 ( .A(DP_OP_424J2_126_3477_n2192), .B(
        DP_OP_424J2_126_3477_n2470), .CI(DP_OP_424J2_126_3477_n2998), .CO(
        DP_OP_424J2_126_3477_n804), .S(DP_OP_424J2_126_3477_n805) );
  FADDX1_HVT DP_OP_424J2_126_3477_U583 ( .A(DP_OP_424J2_126_3477_n2720), .B(
        DP_OP_424J2_126_3477_n2954), .CI(DP_OP_424J2_126_3477_n2514), .CO(
        DP_OP_424J2_126_3477_n802), .S(DP_OP_424J2_126_3477_n803) );
  FADDX1_HVT DP_OP_424J2_126_3477_U582 ( .A(DP_OP_424J2_126_3477_n2676), .B(
        DP_OP_424J2_126_3477_n2426), .CI(DP_OP_424J2_126_3477_n2778), .CO(
        DP_OP_424J2_126_3477_n800), .S(DP_OP_424J2_126_3477_n801) );
  FADDX1_HVT DP_OP_424J2_126_3477_U581 ( .A(DP_OP_424J2_126_3477_n2896), .B(
        DP_OP_424J2_126_3477_n2558), .CI(DP_OP_424J2_126_3477_n2382), .CO(
        DP_OP_424J2_126_3477_n798), .S(DP_OP_424J2_126_3477_n799) );
  FADDX1_HVT DP_OP_424J2_126_3477_U580 ( .A(DP_OP_424J2_126_3477_n2368), .B(
        DP_OP_424J2_126_3477_n2338), .CI(DP_OP_424J2_126_3477_n1986), .CO(
        DP_OP_424J2_126_3477_n796), .S(DP_OP_424J2_126_3477_n797) );
  FADDX1_HVT DP_OP_424J2_126_3477_U579 ( .A(DP_OP_424J2_126_3477_n2588), .B(
        DP_OP_424J2_126_3477_n2250), .CI(DP_OP_424J2_126_3477_n2602), .CO(
        DP_OP_424J2_126_3477_n794), .S(DP_OP_424J2_126_3477_n795) );
  FADDX1_HVT DP_OP_424J2_126_3477_U578 ( .A(DP_OP_424J2_126_3477_n2544), .B(
        DP_OP_424J2_126_3477_n2412), .CI(DP_OP_424J2_126_3477_n2734), .CO(
        DP_OP_424J2_126_3477_n792), .S(DP_OP_424J2_126_3477_n793) );
  FADDX1_HVT DP_OP_424J2_126_3477_U577 ( .A(DP_OP_424J2_126_3477_n2852), .B(
        DP_OP_424J2_126_3477_n2148), .CI(DP_OP_424J2_126_3477_n2324), .CO(
        DP_OP_424J2_126_3477_n790), .S(DP_OP_424J2_126_3477_n791) );
  FADDX1_HVT DP_OP_424J2_126_3477_U576 ( .A(DP_OP_424J2_126_3477_n2016), .B(
        DP_OP_424J2_126_3477_n2632), .CI(DP_OP_424J2_126_3477_n2984), .CO(
        DP_OP_424J2_126_3477_n788), .S(DP_OP_424J2_126_3477_n789) );
  FADDX1_HVT DP_OP_424J2_126_3477_U575 ( .A(DP_OP_424J2_126_3477_n2940), .B(
        DP_OP_424J2_126_3477_n2456), .CI(DP_OP_424J2_126_3477_n821), .CO(
        DP_OP_424J2_126_3477_n786), .S(DP_OP_424J2_126_3477_n787) );
  FADDX1_HVT DP_OP_424J2_126_3477_U574 ( .A(DP_OP_424J2_126_3477_n2287), .B(
        DP_OP_424J2_126_3477_n2023), .CI(DP_OP_424J2_126_3477_n1979), .CO(
        DP_OP_424J2_126_3477_n784), .S(DP_OP_424J2_126_3477_n785) );
  FADDX1_HVT DP_OP_424J2_126_3477_U573 ( .A(DP_OP_424J2_126_3477_n3033), .B(
        DP_OP_424J2_126_3477_n2067), .CI(DP_OP_424J2_126_3477_n2111), .CO(
        DP_OP_424J2_126_3477_n782), .S(DP_OP_424J2_126_3477_n783) );
  FADDX1_HVT DP_OP_424J2_126_3477_U572 ( .A(DP_OP_424J2_126_3477_n2991), .B(
        DP_OP_424J2_126_3477_n2155), .CI(DP_OP_424J2_126_3477_n2199), .CO(
        DP_OP_424J2_126_3477_n780), .S(DP_OP_424J2_126_3477_n781) );
  FADDX1_HVT DP_OP_424J2_126_3477_U571 ( .A(DP_OP_424J2_126_3477_n2947), .B(
        DP_OP_424J2_126_3477_n2243), .CI(DP_OP_424J2_126_3477_n2331), .CO(
        DP_OP_424J2_126_3477_n778), .S(DP_OP_424J2_126_3477_n779) );
  FADDX1_HVT DP_OP_424J2_126_3477_U570 ( .A(DP_OP_424J2_126_3477_n2903), .B(
        DP_OP_424J2_126_3477_n2375), .CI(DP_OP_424J2_126_3477_n2419), .CO(
        DP_OP_424J2_126_3477_n776), .S(DP_OP_424J2_126_3477_n777) );
  FADDX1_HVT DP_OP_424J2_126_3477_U569 ( .A(DP_OP_424J2_126_3477_n2859), .B(
        DP_OP_424J2_126_3477_n2463), .CI(DP_OP_424J2_126_3477_n2507), .CO(
        DP_OP_424J2_126_3477_n774), .S(DP_OP_424J2_126_3477_n775) );
  FADDX1_HVT DP_OP_424J2_126_3477_U568 ( .A(DP_OP_424J2_126_3477_n2815), .B(
        DP_OP_424J2_126_3477_n2551), .CI(DP_OP_424J2_126_3477_n2595), .CO(
        DP_OP_424J2_126_3477_n772), .S(DP_OP_424J2_126_3477_n773) );
  FADDX1_HVT DP_OP_424J2_126_3477_U567 ( .A(DP_OP_424J2_126_3477_n2771), .B(
        DP_OP_424J2_126_3477_n2639), .CI(DP_OP_424J2_126_3477_n2683), .CO(
        DP_OP_424J2_126_3477_n770), .S(DP_OP_424J2_126_3477_n771) );
  FADDX1_HVT DP_OP_424J2_126_3477_U566 ( .A(DP_OP_424J2_126_3477_n2727), .B(
        DP_OP_424J2_126_3477_n1016), .CI(DP_OP_424J2_126_3477_n1014), .CO(
        DP_OP_424J2_126_3477_n768), .S(DP_OP_424J2_126_3477_n769) );
  FADDX1_HVT DP_OP_424J2_126_3477_U565 ( .A(DP_OP_424J2_126_3477_n1012), .B(
        DP_OP_424J2_126_3477_n984), .CI(DP_OP_424J2_126_3477_n986), .CO(
        DP_OP_424J2_126_3477_n766), .S(DP_OP_424J2_126_3477_n767) );
  FADDX1_HVT DP_OP_424J2_126_3477_U564 ( .A(DP_OP_424J2_126_3477_n1010), .B(
        DP_OP_424J2_126_3477_n988), .CI(DP_OP_424J2_126_3477_n990), .CO(
        DP_OP_424J2_126_3477_n764), .S(DP_OP_424J2_126_3477_n765) );
  FADDX1_HVT DP_OP_424J2_126_3477_U563 ( .A(DP_OP_424J2_126_3477_n1008), .B(
        DP_OP_424J2_126_3477_n992), .CI(DP_OP_424J2_126_3477_n994), .CO(
        DP_OP_424J2_126_3477_n762), .S(DP_OP_424J2_126_3477_n763) );
  FADDX1_HVT DP_OP_424J2_126_3477_U562 ( .A(DP_OP_424J2_126_3477_n1000), .B(
        DP_OP_424J2_126_3477_n1006), .CI(DP_OP_424J2_126_3477_n996), .CO(
        DP_OP_424J2_126_3477_n760), .S(DP_OP_424J2_126_3477_n761) );
  FADDX1_HVT DP_OP_424J2_126_3477_U561 ( .A(DP_OP_424J2_126_3477_n998), .B(
        DP_OP_424J2_126_3477_n1002), .CI(DP_OP_424J2_126_3477_n1004), .CO(
        DP_OP_424J2_126_3477_n758), .S(DP_OP_424J2_126_3477_n759) );
  FADDX1_HVT DP_OP_424J2_126_3477_U560 ( .A(DP_OP_424J2_126_3477_n982), .B(
        DP_OP_424J2_126_3477_n980), .CI(DP_OP_424J2_126_3477_n950), .CO(
        DP_OP_424J2_126_3477_n756), .S(DP_OP_424J2_126_3477_n757) );
  FADDX1_HVT DP_OP_424J2_126_3477_U559 ( .A(DP_OP_424J2_126_3477_n964), .B(
        DP_OP_424J2_126_3477_n952), .CI(DP_OP_424J2_126_3477_n954), .CO(
        DP_OP_424J2_126_3477_n754), .S(DP_OP_424J2_126_3477_n755) );
  FADDX1_HVT DP_OP_424J2_126_3477_U557 ( .A(DP_OP_424J2_126_3477_n960), .B(
        DP_OP_424J2_126_3477_n978), .CI(DP_OP_424J2_126_3477_n976), .CO(
        DP_OP_424J2_126_3477_n750), .S(DP_OP_424J2_126_3477_n751) );
  FADDX1_HVT DP_OP_424J2_126_3477_U556 ( .A(DP_OP_424J2_126_3477_n970), .B(
        DP_OP_424J2_126_3477_n966), .CI(DP_OP_424J2_126_3477_n968), .CO(
        DP_OP_424J2_126_3477_n748), .S(DP_OP_424J2_126_3477_n749) );
  FADDX1_HVT DP_OP_424J2_126_3477_U555 ( .A(DP_OP_424J2_126_3477_n974), .B(
        DP_OP_424J2_126_3477_n972), .CI(DP_OP_424J2_126_3477_n813), .CO(
        DP_OP_424J2_126_3477_n746), .S(DP_OP_424J2_126_3477_n747) );
  FADDX1_HVT DP_OP_424J2_126_3477_U554 ( .A(DP_OP_424J2_126_3477_n809), .B(
        DP_OP_424J2_126_3477_n805), .CI(DP_OP_424J2_126_3477_n787), .CO(
        DP_OP_424J2_126_3477_n744), .S(DP_OP_424J2_126_3477_n745) );
  FADDX1_HVT DP_OP_424J2_126_3477_U553 ( .A(DP_OP_424J2_126_3477_n811), .B(
        DP_OP_424J2_126_3477_n793), .CI(DP_OP_424J2_126_3477_n791), .CO(
        DP_OP_424J2_126_3477_n742), .S(DP_OP_424J2_126_3477_n743) );
  FADDX1_HVT DP_OP_424J2_126_3477_U552 ( .A(DP_OP_424J2_126_3477_n803), .B(
        DP_OP_424J2_126_3477_n807), .CI(DP_OP_424J2_126_3477_n799), .CO(
        DP_OP_424J2_126_3477_n740), .S(DP_OP_424J2_126_3477_n741) );
  FADDX1_HVT DP_OP_424J2_126_3477_U551 ( .A(DP_OP_424J2_126_3477_n815), .B(
        DP_OP_424J2_126_3477_n795), .CI(DP_OP_424J2_126_3477_n789), .CO(
        DP_OP_424J2_126_3477_n738), .S(DP_OP_424J2_126_3477_n739) );
  FADDX1_HVT DP_OP_424J2_126_3477_U550 ( .A(DP_OP_424J2_126_3477_n797), .B(
        DP_OP_424J2_126_3477_n819), .CI(DP_OP_424J2_126_3477_n817), .CO(
        DP_OP_424J2_126_3477_n736), .S(DP_OP_424J2_126_3477_n737) );
  FADDX1_HVT DP_OP_424J2_126_3477_U549 ( .A(DP_OP_424J2_126_3477_n801), .B(
        DP_OP_424J2_126_3477_n781), .CI(DP_OP_424J2_126_3477_n777), .CO(
        DP_OP_424J2_126_3477_n734), .S(DP_OP_424J2_126_3477_n735) );
  FADDX1_HVT DP_OP_424J2_126_3477_U548 ( .A(DP_OP_424J2_126_3477_n773), .B(
        DP_OP_424J2_126_3477_n771), .CI(DP_OP_424J2_126_3477_n783), .CO(
        DP_OP_424J2_126_3477_n732), .S(DP_OP_424J2_126_3477_n733) );
  FADDX1_HVT DP_OP_424J2_126_3477_U547 ( .A(DP_OP_424J2_126_3477_n779), .B(
        DP_OP_424J2_126_3477_n775), .CI(DP_OP_424J2_126_3477_n785), .CO(
        DP_OP_424J2_126_3477_n730), .S(DP_OP_424J2_126_3477_n731) );
  FADDX1_HVT DP_OP_424J2_126_3477_U546 ( .A(DP_OP_424J2_126_3477_n948), .B(
        DP_OP_424J2_126_3477_n944), .CI(DP_OP_424J2_126_3477_n946), .CO(
        DP_OP_424J2_126_3477_n728), .S(DP_OP_424J2_126_3477_n729) );
  FADDX1_HVT DP_OP_424J2_126_3477_U545 ( .A(DP_OP_424J2_126_3477_n942), .B(
        DP_OP_424J2_126_3477_n928), .CI(DP_OP_424J2_126_3477_n930), .CO(
        DP_OP_424J2_126_3477_n726), .S(DP_OP_424J2_126_3477_n727) );
  FADDX1_HVT DP_OP_424J2_126_3477_U544 ( .A(DP_OP_424J2_126_3477_n940), .B(
        DP_OP_424J2_126_3477_n932), .CI(DP_OP_424J2_126_3477_n938), .CO(
        DP_OP_424J2_126_3477_n724), .S(DP_OP_424J2_126_3477_n725) );
  FADDX1_HVT DP_OP_424J2_126_3477_U543 ( .A(DP_OP_424J2_126_3477_n936), .B(
        DP_OP_424J2_126_3477_n934), .CI(DP_OP_424J2_126_3477_n769), .CO(
        DP_OP_424J2_126_3477_n722), .S(DP_OP_424J2_126_3477_n723) );
  FADDX1_HVT DP_OP_424J2_126_3477_U542 ( .A(DP_OP_424J2_126_3477_n926), .B(
        DP_OP_424J2_126_3477_n767), .CI(DP_OP_424J2_126_3477_n765), .CO(
        DP_OP_424J2_126_3477_n720), .S(DP_OP_424J2_126_3477_n721) );
  FADDX1_HVT DP_OP_424J2_126_3477_U541 ( .A(DP_OP_424J2_126_3477_n924), .B(
        DP_OP_424J2_126_3477_n761), .CI(DP_OP_424J2_126_3477_n763), .CO(
        DP_OP_424J2_126_3477_n718), .S(DP_OP_424J2_126_3477_n719) );
  FADDX1_HVT DP_OP_424J2_126_3477_U540 ( .A(DP_OP_424J2_126_3477_n922), .B(
        DP_OP_424J2_126_3477_n759), .CI(DP_OP_424J2_126_3477_n916), .CO(
        DP_OP_424J2_126_3477_n716), .S(DP_OP_424J2_126_3477_n717) );
  FADDX1_HVT DP_OP_424J2_126_3477_U539 ( .A(DP_OP_424J2_126_3477_n920), .B(
        DP_OP_424J2_126_3477_n918), .CI(DP_OP_424J2_126_3477_n906), .CO(
        DP_OP_424J2_126_3477_n714), .S(DP_OP_424J2_126_3477_n715) );
  FADDX1_HVT DP_OP_424J2_126_3477_U538 ( .A(DP_OP_424J2_126_3477_n914), .B(
        DP_OP_424J2_126_3477_n757), .CI(DP_OP_424J2_126_3477_n747), .CO(
        DP_OP_424J2_126_3477_n712), .S(DP_OP_424J2_126_3477_n713) );
  FADDX1_HVT DP_OP_424J2_126_3477_U537 ( .A(DP_OP_424J2_126_3477_n912), .B(
        DP_OP_424J2_126_3477_n753), .CI(DP_OP_424J2_126_3477_n749), .CO(
        DP_OP_424J2_126_3477_n710), .S(DP_OP_424J2_126_3477_n711) );
  FADDX1_HVT DP_OP_424J2_126_3477_U536 ( .A(DP_OP_424J2_126_3477_n910), .B(
        DP_OP_424J2_126_3477_n755), .CI(DP_OP_424J2_126_3477_n751), .CO(
        DP_OP_424J2_126_3477_n708), .S(DP_OP_424J2_126_3477_n709) );
  FADDX1_HVT DP_OP_424J2_126_3477_U535 ( .A(DP_OP_424J2_126_3477_n908), .B(
        DP_OP_424J2_126_3477_n743), .CI(DP_OP_424J2_126_3477_n739), .CO(
        DP_OP_424J2_126_3477_n706), .S(DP_OP_424J2_126_3477_n707) );
  FADDX1_HVT DP_OP_424J2_126_3477_U534 ( .A(DP_OP_424J2_126_3477_n741), .B(
        DP_OP_424J2_126_3477_n904), .CI(DP_OP_424J2_126_3477_n735), .CO(
        DP_OP_424J2_126_3477_n704), .S(DP_OP_424J2_126_3477_n705) );
  FADDX1_HVT DP_OP_424J2_126_3477_U533 ( .A(DP_OP_424J2_126_3477_n737), .B(
        DP_OP_424J2_126_3477_n745), .CI(DP_OP_424J2_126_3477_n731), .CO(
        DP_OP_424J2_126_3477_n702), .S(DP_OP_424J2_126_3477_n703) );
  FADDX1_HVT DP_OP_424J2_126_3477_U532 ( .A(DP_OP_424J2_126_3477_n733), .B(
        DP_OP_424J2_126_3477_n902), .CI(DP_OP_424J2_126_3477_n900), .CO(
        DP_OP_424J2_126_3477_n700), .S(DP_OP_424J2_126_3477_n701) );
  FADDX1_HVT DP_OP_424J2_126_3477_U531 ( .A(DP_OP_424J2_126_3477_n898), .B(
        DP_OP_424J2_126_3477_n896), .CI(DP_OP_424J2_126_3477_n729), .CO(
        DP_OP_424J2_126_3477_n698), .S(DP_OP_424J2_126_3477_n699) );
  FADDX1_HVT DP_OP_424J2_126_3477_U530 ( .A(DP_OP_424J2_126_3477_n894), .B(
        DP_OP_424J2_126_3477_n892), .CI(DP_OP_424J2_126_3477_n890), .CO(
        DP_OP_424J2_126_3477_n696), .S(DP_OP_424J2_126_3477_n697) );
  FADDX1_HVT DP_OP_424J2_126_3477_U529 ( .A(DP_OP_424J2_126_3477_n888), .B(
        DP_OP_424J2_126_3477_n723), .CI(DP_OP_424J2_126_3477_n882), .CO(
        DP_OP_424J2_126_3477_n694), .S(DP_OP_424J2_126_3477_n695) );
  FADDX1_HVT DP_OP_424J2_126_3477_U528 ( .A(DP_OP_424J2_126_3477_n886), .B(
        DP_OP_424J2_126_3477_n725), .CI(DP_OP_424J2_126_3477_n727), .CO(
        DP_OP_424J2_126_3477_n692), .S(DP_OP_424J2_126_3477_n693) );
  FADDX1_HVT DP_OP_424J2_126_3477_U527 ( .A(DP_OP_424J2_126_3477_n884), .B(
        DP_OP_424J2_126_3477_n721), .CI(DP_OP_424J2_126_3477_n717), .CO(
        DP_OP_424J2_126_3477_n690), .S(DP_OP_424J2_126_3477_n691) );
  FADDX1_HVT DP_OP_424J2_126_3477_U526 ( .A(DP_OP_424J2_126_3477_n880), .B(
        DP_OP_424J2_126_3477_n719), .CI(DP_OP_424J2_126_3477_n715), .CO(
        DP_OP_424J2_126_3477_n688), .S(DP_OP_424J2_126_3477_n689) );
  FADDX1_HVT DP_OP_424J2_126_3477_U525 ( .A(DP_OP_424J2_126_3477_n878), .B(
        DP_OP_424J2_126_3477_n876), .CI(DP_OP_424J2_126_3477_n711), .CO(
        DP_OP_424J2_126_3477_n686), .S(DP_OP_424J2_126_3477_n687) );
  FADDX1_HVT DP_OP_424J2_126_3477_U524 ( .A(DP_OP_424J2_126_3477_n709), .B(
        DP_OP_424J2_126_3477_n713), .CI(DP_OP_424J2_126_3477_n874), .CO(
        DP_OP_424J2_126_3477_n684), .S(DP_OP_424J2_126_3477_n685) );
  FADDX1_HVT DP_OP_424J2_126_3477_U523 ( .A(DP_OP_424J2_126_3477_n707), .B(
        DP_OP_424J2_126_3477_n872), .CI(DP_OP_424J2_126_3477_n703), .CO(
        DP_OP_424J2_126_3477_n682), .S(DP_OP_424J2_126_3477_n683) );
  FADDX1_HVT DP_OP_424J2_126_3477_U522 ( .A(DP_OP_424J2_126_3477_n705), .B(
        DP_OP_424J2_126_3477_n870), .CI(DP_OP_424J2_126_3477_n701), .CO(
        DP_OP_424J2_126_3477_n680), .S(DP_OP_424J2_126_3477_n681) );
  FADDX1_HVT DP_OP_424J2_126_3477_U521 ( .A(DP_OP_424J2_126_3477_n868), .B(
        DP_OP_424J2_126_3477_n866), .CI(DP_OP_424J2_126_3477_n699), .CO(
        DP_OP_424J2_126_3477_n678), .S(DP_OP_424J2_126_3477_n679) );
  FADDX1_HVT DP_OP_424J2_126_3477_U520 ( .A(DP_OP_424J2_126_3477_n864), .B(
        DP_OP_424J2_126_3477_n862), .CI(DP_OP_424J2_126_3477_n697), .CO(
        DP_OP_424J2_126_3477_n676), .S(DP_OP_424J2_126_3477_n677) );
  FADDX1_HVT DP_OP_424J2_126_3477_U519 ( .A(DP_OP_424J2_126_3477_n860), .B(
        DP_OP_424J2_126_3477_n693), .CI(DP_OP_424J2_126_3477_n856), .CO(
        DP_OP_424J2_126_3477_n674), .S(DP_OP_424J2_126_3477_n675) );
  FADDX1_HVT DP_OP_424J2_126_3477_U518 ( .A(DP_OP_424J2_126_3477_n858), .B(
        DP_OP_424J2_126_3477_n695), .CI(DP_OP_424J2_126_3477_n691), .CO(
        DP_OP_424J2_126_3477_n672), .S(DP_OP_424J2_126_3477_n673) );
  FADDX1_HVT DP_OP_424J2_126_3477_U517 ( .A(DP_OP_424J2_126_3477_n689), .B(
        DP_OP_424J2_126_3477_n854), .CI(DP_OP_424J2_126_3477_n687), .CO(
        DP_OP_424J2_126_3477_n670), .S(DP_OP_424J2_126_3477_n671) );
  FADDX1_HVT DP_OP_424J2_126_3477_U516 ( .A(DP_OP_424J2_126_3477_n685), .B(
        DP_OP_424J2_126_3477_n852), .CI(DP_OP_424J2_126_3477_n683), .CO(
        DP_OP_424J2_126_3477_n668), .S(DP_OP_424J2_126_3477_n669) );
  FADDX1_HVT DP_OP_424J2_126_3477_U515 ( .A(DP_OP_424J2_126_3477_n850), .B(
        DP_OP_424J2_126_3477_n681), .CI(DP_OP_424J2_126_3477_n848), .CO(
        DP_OP_424J2_126_3477_n666), .S(DP_OP_424J2_126_3477_n667) );
  FADDX1_HVT DP_OP_424J2_126_3477_U514 ( .A(DP_OP_424J2_126_3477_n846), .B(
        DP_OP_424J2_126_3477_n679), .CI(DP_OP_424J2_126_3477_n844), .CO(
        DP_OP_424J2_126_3477_n664), .S(DP_OP_424J2_126_3477_n665) );
  FADDX1_HVT DP_OP_424J2_126_3477_U513 ( .A(DP_OP_424J2_126_3477_n677), .B(
        DP_OP_424J2_126_3477_n675), .CI(DP_OP_424J2_126_3477_n842), .CO(
        DP_OP_424J2_126_3477_n662), .S(DP_OP_424J2_126_3477_n663) );
  FADDX1_HVT DP_OP_424J2_126_3477_U512 ( .A(DP_OP_424J2_126_3477_n673), .B(
        DP_OP_424J2_126_3477_n671), .CI(DP_OP_424J2_126_3477_n840), .CO(
        DP_OP_424J2_126_3477_n660), .S(DP_OP_424J2_126_3477_n661) );
  FADDX1_HVT DP_OP_424J2_126_3477_U511 ( .A(DP_OP_424J2_126_3477_n669), .B(
        DP_OP_424J2_126_3477_n838), .CI(DP_OP_424J2_126_3477_n836), .CO(
        DP_OP_424J2_126_3477_n658), .S(DP_OP_424J2_126_3477_n659) );
  FADDX1_HVT DP_OP_424J2_126_3477_U510 ( .A(DP_OP_424J2_126_3477_n667), .B(
        DP_OP_424J2_126_3477_n834), .CI(DP_OP_424J2_126_3477_n665), .CO(
        DP_OP_424J2_126_3477_n656), .S(DP_OP_424J2_126_3477_n657) );
  FADDX1_HVT DP_OP_424J2_126_3477_U509 ( .A(DP_OP_424J2_126_3477_n663), .B(
        DP_OP_424J2_126_3477_n832), .CI(DP_OP_424J2_126_3477_n661), .CO(
        DP_OP_424J2_126_3477_n654), .S(DP_OP_424J2_126_3477_n655) );
  FADDX1_HVT DP_OP_424J2_126_3477_U508 ( .A(DP_OP_424J2_126_3477_n830), .B(
        DP_OP_424J2_126_3477_n659), .CI(DP_OP_424J2_126_3477_n828), .CO(
        DP_OP_424J2_126_3477_n652), .S(DP_OP_424J2_126_3477_n653) );
  FADDX1_HVT DP_OP_424J2_126_3477_U507 ( .A(DP_OP_424J2_126_3477_n657), .B(
        DP_OP_424J2_126_3477_n826), .CI(DP_OP_424J2_126_3477_n655), .CO(
        DP_OP_424J2_126_3477_n650), .S(DP_OP_424J2_126_3477_n651) );
  FADDX1_HVT DP_OP_424J2_126_3477_U506 ( .A(DP_OP_424J2_126_3477_n824), .B(
        DP_OP_424J2_126_3477_n651), .CI(DP_OP_424J2_126_3477_n653), .CO(
        DP_OP_424J2_126_3477_n648), .S(DP_OP_424J2_126_3477_n649) );
  FADDX1_HVT DP_OP_424J2_126_3477_U505 ( .A(DP_OP_424J2_126_3477_n3027), .B(
        DP_OP_424J2_126_3477_n1971), .CI(DP_OP_424J2_126_3477_n1927), .CO(
        DP_OP_424J2_126_3477_n646), .S(DP_OP_424J2_126_3477_n647) );
  FADDX1_HVT DP_OP_424J2_126_3477_U504 ( .A(DP_OP_424J2_126_3477_n820), .B(
        DP_OP_424J2_126_3477_n2286), .CI(DP_OP_424J2_126_3477_n1978), .CO(
        DP_OP_424J2_126_3477_n644), .S(DP_OP_424J2_126_3477_n645) );
  FADDX1_HVT DP_OP_424J2_126_3477_U503 ( .A(DP_OP_424J2_126_3477_n2367), .B(
        DP_OP_424J2_126_3477_n3032), .CI(DP_OP_424J2_126_3477_n2682), .CO(
        DP_OP_424J2_126_3477_n642), .S(DP_OP_424J2_126_3477_n643) );
  FADDX1_HVT DP_OP_424J2_126_3477_U502 ( .A(DP_OP_424J2_126_3477_n2059), .B(
        DP_OP_424J2_126_3477_n2594), .CI(DP_OP_424J2_126_3477_n2814), .CO(
        DP_OP_424J2_126_3477_n640), .S(DP_OP_424J2_126_3477_n641) );
  FADDX1_HVT DP_OP_424J2_126_3477_U501 ( .A(DP_OP_424J2_126_3477_n2279), .B(
        DP_OP_424J2_126_3477_n2374), .CI(DP_OP_424J2_126_3477_n2990), .CO(
        DP_OP_424J2_126_3477_n638), .S(DP_OP_424J2_126_3477_n639) );
  FADDX1_HVT DP_OP_424J2_126_3477_U500 ( .A(DP_OP_424J2_126_3477_n2015), .B(
        DP_OP_424J2_126_3477_n2902), .CI(DP_OP_424J2_126_3477_n2066), .CO(
        DP_OP_424J2_126_3477_n636), .S(DP_OP_424J2_126_3477_n637) );
  FADDX1_HVT DP_OP_424J2_126_3477_U499 ( .A(DP_OP_424J2_126_3477_n2147), .B(
        DP_OP_424J2_126_3477_n2022), .CI(DP_OP_424J2_126_3477_n2858), .CO(
        DP_OP_424J2_126_3477_n634), .S(DP_OP_424J2_126_3477_n635) );
  FADDX1_HVT DP_OP_424J2_126_3477_U498 ( .A(DP_OP_424J2_126_3477_n2983), .B(
        DP_OP_424J2_126_3477_n2418), .CI(DP_OP_424J2_126_3477_n2506), .CO(
        DP_OP_424J2_126_3477_n632), .S(DP_OP_424J2_126_3477_n633) );
  FADDX1_HVT DP_OP_424J2_126_3477_U497 ( .A(DP_OP_424J2_126_3477_n2499), .B(
        DP_OP_424J2_126_3477_n2550), .CI(DP_OP_424J2_126_3477_n2946), .CO(
        DP_OP_424J2_126_3477_n630), .S(DP_OP_424J2_126_3477_n631) );
  FADDX1_HVT DP_OP_424J2_126_3477_U496 ( .A(DP_OP_424J2_126_3477_n2763), .B(
        DP_OP_424J2_126_3477_n2242), .CI(DP_OP_424J2_126_3477_n2770), .CO(
        DP_OP_424J2_126_3477_n628), .S(DP_OP_424J2_126_3477_n629) );
  FADDX1_HVT DP_OP_424J2_126_3477_U495 ( .A(DP_OP_424J2_126_3477_n2939), .B(
        DP_OP_424J2_126_3477_n2462), .CI(DP_OP_424J2_126_3477_n2638), .CO(
        DP_OP_424J2_126_3477_n626), .S(DP_OP_424J2_126_3477_n627) );
  FADDX1_HVT DP_OP_424J2_126_3477_U494 ( .A(DP_OP_424J2_126_3477_n2235), .B(
        DP_OP_424J2_126_3477_n2110), .CI(DP_OP_424J2_126_3477_n2726), .CO(
        DP_OP_424J2_126_3477_n624), .S(DP_OP_424J2_126_3477_n625) );
  FADDX1_HVT DP_OP_424J2_126_3477_U493 ( .A(DP_OP_424J2_126_3477_n2191), .B(
        DP_OP_424J2_126_3477_n2330), .CI(DP_OP_424J2_126_3477_n2198), .CO(
        DP_OP_424J2_126_3477_n622), .S(DP_OP_424J2_126_3477_n623) );
  FADDX1_HVT DP_OP_424J2_126_3477_U492 ( .A(DP_OP_424J2_126_3477_n2587), .B(
        DP_OP_424J2_126_3477_n2411), .CI(DP_OP_424J2_126_3477_n2154), .CO(
        DP_OP_424J2_126_3477_n620), .S(DP_OP_424J2_126_3477_n621) );
  FADDX1_HVT DP_OP_424J2_126_3477_U491 ( .A(DP_OP_424J2_126_3477_n2895), .B(
        DP_OP_424J2_126_3477_n2103), .CI(DP_OP_424J2_126_3477_n2323), .CO(
        DP_OP_424J2_126_3477_n618), .S(DP_OP_424J2_126_3477_n619) );
  FADDX1_HVT DP_OP_424J2_126_3477_U490 ( .A(DP_OP_424J2_126_3477_n2851), .B(
        DP_OP_424J2_126_3477_n2455), .CI(DP_OP_424J2_126_3477_n2543), .CO(
        DP_OP_424J2_126_3477_n616), .S(DP_OP_424J2_126_3477_n617) );
  FADDX1_HVT DP_OP_424J2_126_3477_U489 ( .A(DP_OP_424J2_126_3477_n2807), .B(
        DP_OP_424J2_126_3477_n2631), .CI(DP_OP_424J2_126_3477_n2675), .CO(
        DP_OP_424J2_126_3477_n614), .S(DP_OP_424J2_126_3477_n615) );
  FADDX1_HVT DP_OP_424J2_126_3477_U488 ( .A(DP_OP_424J2_126_3477_n2719), .B(
        DP_OP_424J2_126_3477_n818), .CI(DP_OP_424J2_126_3477_n816), .CO(
        DP_OP_424J2_126_3477_n612), .S(DP_OP_424J2_126_3477_n613) );
  FADDX1_HVT DP_OP_424J2_126_3477_U487 ( .A(DP_OP_424J2_126_3477_n814), .B(
        DP_OP_424J2_126_3477_n786), .CI(DP_OP_424J2_126_3477_n788), .CO(
        DP_OP_424J2_126_3477_n610), .S(DP_OP_424J2_126_3477_n611) );
  FADDX1_HVT DP_OP_424J2_126_3477_U486 ( .A(DP_OP_424J2_126_3477_n812), .B(
        DP_OP_424J2_126_3477_n790), .CI(DP_OP_424J2_126_3477_n792), .CO(
        DP_OP_424J2_126_3477_n608), .S(DP_OP_424J2_126_3477_n609) );
  FADDX1_HVT DP_OP_424J2_126_3477_U485 ( .A(DP_OP_424J2_126_3477_n810), .B(
        DP_OP_424J2_126_3477_n794), .CI(DP_OP_424J2_126_3477_n796), .CO(
        DP_OP_424J2_126_3477_n606), .S(DP_OP_424J2_126_3477_n607) );
  FADDX1_HVT DP_OP_424J2_126_3477_U484 ( .A(DP_OP_424J2_126_3477_n808), .B(
        DP_OP_424J2_126_3477_n798), .CI(DP_OP_424J2_126_3477_n800), .CO(
        DP_OP_424J2_126_3477_n604), .S(DP_OP_424J2_126_3477_n605) );
  FADDX1_HVT DP_OP_424J2_126_3477_U483 ( .A(DP_OP_424J2_126_3477_n806), .B(
        DP_OP_424J2_126_3477_n802), .CI(DP_OP_424J2_126_3477_n804), .CO(
        DP_OP_424J2_126_3477_n602), .S(DP_OP_424J2_126_3477_n603) );
  FADDX1_HVT DP_OP_424J2_126_3477_U482 ( .A(DP_OP_424J2_126_3477_n784), .B(
        DP_OP_424J2_126_3477_n770), .CI(DP_OP_424J2_126_3477_n782), .CO(
        DP_OP_424J2_126_3477_n600), .S(DP_OP_424J2_126_3477_n601) );
  FADDX1_HVT DP_OP_424J2_126_3477_U481 ( .A(DP_OP_424J2_126_3477_n776), .B(
        DP_OP_424J2_126_3477_n772), .CI(DP_OP_424J2_126_3477_n774), .CO(
        DP_OP_424J2_126_3477_n598), .S(DP_OP_424J2_126_3477_n599) );
  FADDX1_HVT DP_OP_424J2_126_3477_U480 ( .A(DP_OP_424J2_126_3477_n780), .B(
        DP_OP_424J2_126_3477_n778), .CI(DP_OP_424J2_126_3477_n645), .CO(
        DP_OP_424J2_126_3477_n596), .S(DP_OP_424J2_126_3477_n597) );
  FADDX1_HVT DP_OP_424J2_126_3477_U479 ( .A(DP_OP_424J2_126_3477_n647), .B(
        DP_OP_424J2_126_3477_n633), .CI(DP_OP_424J2_126_3477_n639), .CO(
        DP_OP_424J2_126_3477_n594), .S(DP_OP_424J2_126_3477_n595) );
  FADDX1_HVT DP_OP_424J2_126_3477_U478 ( .A(DP_OP_424J2_126_3477_n615), .B(
        DP_OP_424J2_126_3477_n637), .CI(DP_OP_424J2_126_3477_n635), .CO(
        DP_OP_424J2_126_3477_n592), .S(DP_OP_424J2_126_3477_n593) );
  FADDX1_HVT DP_OP_424J2_126_3477_U477 ( .A(DP_OP_424J2_126_3477_n641), .B(
        DP_OP_424J2_126_3477_n623), .CI(DP_OP_424J2_126_3477_n625), .CO(
        DP_OP_424J2_126_3477_n590), .S(DP_OP_424J2_126_3477_n591) );
  FADDX1_HVT DP_OP_424J2_126_3477_U476 ( .A(DP_OP_424J2_126_3477_n627), .B(
        DP_OP_424J2_126_3477_n617), .CI(DP_OP_424J2_126_3477_n619), .CO(
        DP_OP_424J2_126_3477_n588), .S(DP_OP_424J2_126_3477_n589) );
  FADDX1_HVT DP_OP_424J2_126_3477_U475 ( .A(DP_OP_424J2_126_3477_n621), .B(
        DP_OP_424J2_126_3477_n643), .CI(DP_OP_424J2_126_3477_n631), .CO(
        DP_OP_424J2_126_3477_n586), .S(DP_OP_424J2_126_3477_n587) );
  FADDX1_HVT DP_OP_424J2_126_3477_U474 ( .A(DP_OP_424J2_126_3477_n629), .B(
        DP_OP_424J2_126_3477_n768), .CI(DP_OP_424J2_126_3477_n766), .CO(
        DP_OP_424J2_126_3477_n584), .S(DP_OP_424J2_126_3477_n585) );
  FADDX1_HVT DP_OP_424J2_126_3477_U473 ( .A(DP_OP_424J2_126_3477_n764), .B(
        DP_OP_424J2_126_3477_n758), .CI(DP_OP_424J2_126_3477_n760), .CO(
        DP_OP_424J2_126_3477_n582), .S(DP_OP_424J2_126_3477_n583) );
  FADDX1_HVT DP_OP_424J2_126_3477_U472 ( .A(DP_OP_424J2_126_3477_n762), .B(
        DP_OP_424J2_126_3477_n756), .CI(DP_OP_424J2_126_3477_n754), .CO(
        DP_OP_424J2_126_3477_n580), .S(DP_OP_424J2_126_3477_n581) );
  FADDX1_HVT DP_OP_424J2_126_3477_U470 ( .A(DP_OP_424J2_126_3477_n750), .B(
        DP_OP_424J2_126_3477_n613), .CI(DP_OP_424J2_126_3477_n607), .CO(
        DP_OP_424J2_126_3477_n576), .S(DP_OP_424J2_126_3477_n577) );
  FADDX1_HVT DP_OP_424J2_126_3477_U469 ( .A(DP_OP_424J2_126_3477_n609), .B(
        DP_OP_424J2_126_3477_n603), .CI(DP_OP_424J2_126_3477_n734), .CO(
        DP_OP_424J2_126_3477_n574), .S(DP_OP_424J2_126_3477_n575) );
  FADDX1_HVT DP_OP_424J2_126_3477_U468 ( .A(DP_OP_424J2_126_3477_n744), .B(
        DP_OP_424J2_126_3477_n611), .CI(DP_OP_424J2_126_3477_n605), .CO(
        DP_OP_424J2_126_3477_n572), .S(DP_OP_424J2_126_3477_n573) );
  FADDX1_HVT DP_OP_424J2_126_3477_U467 ( .A(DP_OP_424J2_126_3477_n738), .B(
        DP_OP_424J2_126_3477_n742), .CI(DP_OP_424J2_126_3477_n736), .CO(
        DP_OP_424J2_126_3477_n570), .S(DP_OP_424J2_126_3477_n571) );
  FADDX1_HVT DP_OP_424J2_126_3477_U466 ( .A(DP_OP_424J2_126_3477_n740), .B(
        DP_OP_424J2_126_3477_n732), .CI(DP_OP_424J2_126_3477_n730), .CO(
        DP_OP_424J2_126_3477_n568), .S(DP_OP_424J2_126_3477_n569) );
  FADDX1_HVT DP_OP_424J2_126_3477_U465 ( .A(DP_OP_424J2_126_3477_n599), .B(
        DP_OP_424J2_126_3477_n601), .CI(DP_OP_424J2_126_3477_n597), .CO(
        DP_OP_424J2_126_3477_n566), .S(DP_OP_424J2_126_3477_n567) );
  FADDX1_HVT DP_OP_424J2_126_3477_U464 ( .A(DP_OP_424J2_126_3477_n595), .B(
        DP_OP_424J2_126_3477_n589), .CI(DP_OP_424J2_126_3477_n593), .CO(
        DP_OP_424J2_126_3477_n564), .S(DP_OP_424J2_126_3477_n565) );
  FADDX1_HVT DP_OP_424J2_126_3477_U463 ( .A(DP_OP_424J2_126_3477_n587), .B(
        DP_OP_424J2_126_3477_n591), .CI(DP_OP_424J2_126_3477_n728), .CO(
        DP_OP_424J2_126_3477_n562), .S(DP_OP_424J2_126_3477_n563) );
  FADDX1_HVT DP_OP_424J2_126_3477_U462 ( .A(DP_OP_424J2_126_3477_n726), .B(
        DP_OP_424J2_126_3477_n585), .CI(DP_OP_424J2_126_3477_n722), .CO(
        DP_OP_424J2_126_3477_n560), .S(DP_OP_424J2_126_3477_n561) );
  FADDX1_HVT DP_OP_424J2_126_3477_U461 ( .A(DP_OP_424J2_126_3477_n724), .B(
        DP_OP_424J2_126_3477_n720), .CI(DP_OP_424J2_126_3477_n718), .CO(
        DP_OP_424J2_126_3477_n558), .S(DP_OP_424J2_126_3477_n559) );
  FADDX1_HVT DP_OP_424J2_126_3477_U460 ( .A(DP_OP_424J2_126_3477_n716), .B(
        DP_OP_424J2_126_3477_n583), .CI(DP_OP_424J2_126_3477_n581), .CO(
        DP_OP_424J2_126_3477_n556), .S(DP_OP_424J2_126_3477_n557) );
  FADDX1_HVT DP_OP_424J2_126_3477_U459 ( .A(DP_OP_424J2_126_3477_n714), .B(
        DP_OP_424J2_126_3477_n712), .CI(DP_OP_424J2_126_3477_n710), .CO(
        DP_OP_424J2_126_3477_n554), .S(DP_OP_424J2_126_3477_n555) );
  FADDX1_HVT DP_OP_424J2_126_3477_U458 ( .A(DP_OP_424J2_126_3477_n708), .B(
        DP_OP_424J2_126_3477_n579), .CI(DP_OP_424J2_126_3477_n706), .CO(
        DP_OP_424J2_126_3477_n552), .S(DP_OP_424J2_126_3477_n553) );
  FADDX1_HVT DP_OP_424J2_126_3477_U457 ( .A(DP_OP_424J2_126_3477_n577), .B(
        DP_OP_424J2_126_3477_n704), .CI(DP_OP_424J2_126_3477_n575), .CO(
        DP_OP_424J2_126_3477_n550), .S(DP_OP_424J2_126_3477_n551) );
  FADDX1_HVT DP_OP_424J2_126_3477_U456 ( .A(DP_OP_424J2_126_3477_n702), .B(
        DP_OP_424J2_126_3477_n571), .CI(DP_OP_424J2_126_3477_n569), .CO(
        DP_OP_424J2_126_3477_n548), .S(DP_OP_424J2_126_3477_n549) );
  FADDX1_HVT DP_OP_424J2_126_3477_U455 ( .A(DP_OP_424J2_126_3477_n573), .B(
        DP_OP_424J2_126_3477_n567), .CI(DP_OP_424J2_126_3477_n700), .CO(
        DP_OP_424J2_126_3477_n546), .S(DP_OP_424J2_126_3477_n547) );
  FADDX1_HVT DP_OP_424J2_126_3477_U454 ( .A(DP_OP_424J2_126_3477_n565), .B(
        DP_OP_424J2_126_3477_n698), .CI(DP_OP_424J2_126_3477_n563), .CO(
        DP_OP_424J2_126_3477_n544), .S(DP_OP_424J2_126_3477_n545) );
  FADDX1_HVT DP_OP_424J2_126_3477_U453 ( .A(DP_OP_424J2_126_3477_n696), .B(
        DP_OP_424J2_126_3477_n694), .CI(DP_OP_424J2_126_3477_n692), .CO(
        DP_OP_424J2_126_3477_n542), .S(DP_OP_424J2_126_3477_n543) );
  FADDX1_HVT DP_OP_424J2_126_3477_U452 ( .A(DP_OP_424J2_126_3477_n561), .B(
        DP_OP_424J2_126_3477_n690), .CI(DP_OP_424J2_126_3477_n559), .CO(
        DP_OP_424J2_126_3477_n540), .S(DP_OP_424J2_126_3477_n541) );
  FADDX1_HVT DP_OP_424J2_126_3477_U451 ( .A(DP_OP_424J2_126_3477_n688), .B(
        DP_OP_424J2_126_3477_n557), .CI(DP_OP_424J2_126_3477_n555), .CO(
        DP_OP_424J2_126_3477_n538), .S(DP_OP_424J2_126_3477_n539) );
  FADDX1_HVT DP_OP_424J2_126_3477_U449 ( .A(DP_OP_424J2_126_3477_n682), .B(
        DP_OP_424J2_126_3477_n551), .CI(DP_OP_424J2_126_3477_n549), .CO(
        DP_OP_424J2_126_3477_n534), .S(DP_OP_424J2_126_3477_n535) );
  FADDX1_HVT DP_OP_424J2_126_3477_U448 ( .A(DP_OP_424J2_126_3477_n680), .B(
        DP_OP_424J2_126_3477_n547), .CI(DP_OP_424J2_126_3477_n678), .CO(
        DP_OP_424J2_126_3477_n532), .S(DP_OP_424J2_126_3477_n533) );
  FADDX1_HVT DP_OP_424J2_126_3477_U447 ( .A(DP_OP_424J2_126_3477_n545), .B(
        DP_OP_424J2_126_3477_n676), .CI(DP_OP_424J2_126_3477_n543), .CO(
        DP_OP_424J2_126_3477_n530), .S(DP_OP_424J2_126_3477_n531) );
  FADDX1_HVT DP_OP_424J2_126_3477_U446 ( .A(DP_OP_424J2_126_3477_n674), .B(
        DP_OP_424J2_126_3477_n672), .CI(DP_OP_424J2_126_3477_n541), .CO(
        DP_OP_424J2_126_3477_n528), .S(DP_OP_424J2_126_3477_n529) );
  FADDX1_HVT DP_OP_424J2_126_3477_U445 ( .A(DP_OP_424J2_126_3477_n670), .B(
        DP_OP_424J2_126_3477_n539), .CI(DP_OP_424J2_126_3477_n537), .CO(
        DP_OP_424J2_126_3477_n526), .S(DP_OP_424J2_126_3477_n527) );
  FADDX1_HVT DP_OP_424J2_126_3477_U443 ( .A(DP_OP_424J2_126_3477_n533), .B(
        DP_OP_424J2_126_3477_n664), .CI(DP_OP_424J2_126_3477_n531), .CO(
        DP_OP_424J2_126_3477_n522), .S(DP_OP_424J2_126_3477_n523) );
  FADDX1_HVT DP_OP_424J2_126_3477_U442 ( .A(DP_OP_424J2_126_3477_n662), .B(
        DP_OP_424J2_126_3477_n529), .CI(DP_OP_424J2_126_3477_n660), .CO(
        DP_OP_424J2_126_3477_n520), .S(DP_OP_424J2_126_3477_n521) );
  FADDX1_HVT DP_OP_424J2_126_3477_U441 ( .A(DP_OP_424J2_126_3477_n527), .B(
        DP_OP_424J2_126_3477_n525), .CI(DP_OP_424J2_126_3477_n658), .CO(
        DP_OP_424J2_126_3477_n518), .S(DP_OP_424J2_126_3477_n519) );
  FADDX1_HVT DP_OP_424J2_126_3477_U440 ( .A(DP_OP_424J2_126_3477_n523), .B(
        DP_OP_424J2_126_3477_n656), .CI(DP_OP_424J2_126_3477_n654), .CO(
        DP_OP_424J2_126_3477_n516), .S(DP_OP_424J2_126_3477_n517) );
  FADDX1_HVT DP_OP_424J2_126_3477_U439 ( .A(DP_OP_424J2_126_3477_n521), .B(
        DP_OP_424J2_126_3477_n519), .CI(DP_OP_424J2_126_3477_n652), .CO(
        DP_OP_424J2_126_3477_n514), .S(DP_OP_424J2_126_3477_n515) );
  FADDX1_HVT DP_OP_424J2_126_3477_U438 ( .A(DP_OP_424J2_126_3477_n650), .B(
        DP_OP_424J2_126_3477_n517), .CI(DP_OP_424J2_126_3477_n515), .CO(
        DP_OP_424J2_126_3477_n512), .S(DP_OP_424J2_126_3477_n513) );
  FADDX1_HVT DP_OP_424J2_126_3477_U435 ( .A(DP_OP_424J2_126_3477_n2058), .B(
        DP_OP_424J2_126_3477_n2982), .CI(DP_OP_424J2_126_3477_n2410), .CO(
        DP_OP_424J2_126_3477_n506), .S(DP_OP_424J2_126_3477_n507) );
  FADDX1_HVT DP_OP_424J2_126_3477_U434 ( .A(DP_OP_424J2_126_3477_n2542), .B(
        DP_OP_424J2_126_3477_n2938), .CI(DP_OP_424J2_126_3477_n2894), .CO(
        DP_OP_424J2_126_3477_n504), .S(DP_OP_424J2_126_3477_n505) );
  FADDX1_HVT DP_OP_424J2_126_3477_U433 ( .A(DP_OP_424J2_126_3477_n2366), .B(
        DP_OP_424J2_126_3477_n2850), .CI(DP_OP_424J2_126_3477_n2806), .CO(
        DP_OP_424J2_126_3477_n502), .S(DP_OP_424J2_126_3477_n503) );
  FADDX1_HVT DP_OP_424J2_126_3477_U432 ( .A(DP_OP_424J2_126_3477_n2234), .B(
        DP_OP_424J2_126_3477_n2014), .CI(DP_OP_424J2_126_3477_n2762), .CO(
        DP_OP_424J2_126_3477_n500), .S(DP_OP_424J2_126_3477_n501) );
  FADDX1_HVT DP_OP_424J2_126_3477_U431 ( .A(DP_OP_424J2_126_3477_n2718), .B(
        DP_OP_424J2_126_3477_n2674), .CI(DP_OP_424J2_126_3477_n2630), .CO(
        DP_OP_424J2_126_3477_n498), .S(DP_OP_424J2_126_3477_n499) );
  FADDX1_HVT DP_OP_424J2_126_3477_U430 ( .A(DP_OP_424J2_126_3477_n2278), .B(
        DP_OP_424J2_126_3477_n2102), .CI(DP_OP_424J2_126_3477_n2146), .CO(
        DP_OP_424J2_126_3477_n496), .S(DP_OP_424J2_126_3477_n497) );
  FADDX1_HVT DP_OP_424J2_126_3477_U429 ( .A(DP_OP_424J2_126_3477_n2190), .B(
        DP_OP_424J2_126_3477_n2586), .CI(DP_OP_424J2_126_3477_n2498), .CO(
        DP_OP_424J2_126_3477_n494), .S(DP_OP_424J2_126_3477_n495) );
  FADDX1_HVT DP_OP_424J2_126_3477_U428 ( .A(DP_OP_424J2_126_3477_n2322), .B(
        DP_OP_424J2_126_3477_n2454), .CI(DP_OP_424J2_126_3477_n646), .CO(
        DP_OP_424J2_126_3477_n492), .S(DP_OP_424J2_126_3477_n493) );
  FADDX1_HVT DP_OP_424J2_126_3477_U427 ( .A(DP_OP_424J2_126_3477_n644), .B(
        DP_OP_424J2_126_3477_n614), .CI(DP_OP_424J2_126_3477_n642), .CO(
        DP_OP_424J2_126_3477_n490), .S(DP_OP_424J2_126_3477_n491) );
  FADDX1_HVT DP_OP_424J2_126_3477_U426 ( .A(DP_OP_424J2_126_3477_n640), .B(
        DP_OP_424J2_126_3477_n616), .CI(DP_OP_424J2_126_3477_n618), .CO(
        DP_OP_424J2_126_3477_n488), .S(DP_OP_424J2_126_3477_n489) );
  FADDX1_HVT DP_OP_424J2_126_3477_U425 ( .A(DP_OP_424J2_126_3477_n638), .B(
        DP_OP_424J2_126_3477_n620), .CI(DP_OP_424J2_126_3477_n622), .CO(
        DP_OP_424J2_126_3477_n486), .S(DP_OP_424J2_126_3477_n487) );
  FADDX1_HVT DP_OP_424J2_126_3477_U424 ( .A(DP_OP_424J2_126_3477_n636), .B(
        DP_OP_424J2_126_3477_n624), .CI(DP_OP_424J2_126_3477_n626), .CO(
        DP_OP_424J2_126_3477_n484), .S(DP_OP_424J2_126_3477_n485) );
  FADDX1_HVT DP_OP_424J2_126_3477_U423 ( .A(DP_OP_424J2_126_3477_n634), .B(
        DP_OP_424J2_126_3477_n628), .CI(DP_OP_424J2_126_3477_n630), .CO(
        DP_OP_424J2_126_3477_n482), .S(DP_OP_424J2_126_3477_n483) );
  FADDX1_HVT DP_OP_424J2_126_3477_U422 ( .A(DP_OP_424J2_126_3477_n632), .B(
        DP_OP_424J2_126_3477_n509), .CI(DP_OP_424J2_126_3477_n505), .CO(
        DP_OP_424J2_126_3477_n480), .S(DP_OP_424J2_126_3477_n481) );
  FADDX1_HVT DP_OP_424J2_126_3477_U421 ( .A(DP_OP_424J2_126_3477_n501), .B(
        DP_OP_424J2_126_3477_n495), .CI(DP_OP_424J2_126_3477_n497), .CO(
        DP_OP_424J2_126_3477_n478), .S(DP_OP_424J2_126_3477_n479) );
  FADDX1_HVT DP_OP_424J2_126_3477_U420 ( .A(DP_OP_424J2_126_3477_n499), .B(
        DP_OP_424J2_126_3477_n507), .CI(DP_OP_424J2_126_3477_n503), .CO(
        DP_OP_424J2_126_3477_n476), .S(DP_OP_424J2_126_3477_n477) );
  FADDX1_HVT DP_OP_424J2_126_3477_U419 ( .A(DP_OP_424J2_126_3477_n612), .B(
        DP_OP_424J2_126_3477_n610), .CI(DP_OP_424J2_126_3477_n602), .CO(
        DP_OP_424J2_126_3477_n474), .S(DP_OP_424J2_126_3477_n475) );
  FADDX1_HVT DP_OP_424J2_126_3477_U418 ( .A(DP_OP_424J2_126_3477_n608), .B(
        DP_OP_424J2_126_3477_n604), .CI(DP_OP_424J2_126_3477_n606), .CO(
        DP_OP_424J2_126_3477_n472), .S(DP_OP_424J2_126_3477_n473) );
  FADDX1_HVT DP_OP_424J2_126_3477_U417 ( .A(DP_OP_424J2_126_3477_n600), .B(
        DP_OP_424J2_126_3477_n596), .CI(DP_OP_424J2_126_3477_n493), .CO(
        DP_OP_424J2_126_3477_n470), .S(DP_OP_424J2_126_3477_n471) );
  FADDX1_HVT DP_OP_424J2_126_3477_U416 ( .A(DP_OP_424J2_126_3477_n598), .B(
        DP_OP_424J2_126_3477_n594), .CI(DP_OP_424J2_126_3477_n491), .CO(
        DP_OP_424J2_126_3477_n468), .S(DP_OP_424J2_126_3477_n469) );
  FADDX1_HVT DP_OP_424J2_126_3477_U415 ( .A(DP_OP_424J2_126_3477_n592), .B(
        DP_OP_424J2_126_3477_n485), .CI(DP_OP_424J2_126_3477_n487), .CO(
        DP_OP_424J2_126_3477_n466), .S(DP_OP_424J2_126_3477_n467) );
  FADDX1_HVT DP_OP_424J2_126_3477_U414 ( .A(DP_OP_424J2_126_3477_n590), .B(
        DP_OP_424J2_126_3477_n489), .CI(DP_OP_424J2_126_3477_n483), .CO(
        DP_OP_424J2_126_3477_n464), .S(DP_OP_424J2_126_3477_n465) );
  FADDX1_HVT DP_OP_424J2_126_3477_U413 ( .A(DP_OP_424J2_126_3477_n588), .B(
        DP_OP_424J2_126_3477_n586), .CI(DP_OP_424J2_126_3477_n584), .CO(
        DP_OP_424J2_126_3477_n462), .S(DP_OP_424J2_126_3477_n463) );
  FADDX1_HVT DP_OP_424J2_126_3477_U412 ( .A(DP_OP_424J2_126_3477_n481), .B(
        DP_OP_424J2_126_3477_n477), .CI(DP_OP_424J2_126_3477_n582), .CO(
        DP_OP_424J2_126_3477_n460), .S(DP_OP_424J2_126_3477_n461) );
  FADDX1_HVT DP_OP_424J2_126_3477_U411 ( .A(DP_OP_424J2_126_3477_n479), .B(
        DP_OP_424J2_126_3477_n580), .CI(DP_OP_424J2_126_3477_n578), .CO(
        DP_OP_424J2_126_3477_n458), .S(DP_OP_424J2_126_3477_n459) );
  FADDX1_HVT DP_OP_424J2_126_3477_U410 ( .A(DP_OP_424J2_126_3477_n576), .B(
        DP_OP_424J2_126_3477_n475), .CI(DP_OP_424J2_126_3477_n473), .CO(
        DP_OP_424J2_126_3477_n456), .S(DP_OP_424J2_126_3477_n457) );
  FADDX1_HVT DP_OP_424J2_126_3477_U409 ( .A(DP_OP_424J2_126_3477_n574), .B(
        DP_OP_424J2_126_3477_n570), .CI(DP_OP_424J2_126_3477_n568), .CO(
        DP_OP_424J2_126_3477_n454), .S(DP_OP_424J2_126_3477_n455) );
  FADDX1_HVT DP_OP_424J2_126_3477_U408 ( .A(DP_OP_424J2_126_3477_n572), .B(
        DP_OP_424J2_126_3477_n566), .CI(DP_OP_424J2_126_3477_n471), .CO(
        DP_OP_424J2_126_3477_n452), .S(DP_OP_424J2_126_3477_n453) );
  FADDX1_HVT DP_OP_424J2_126_3477_U407 ( .A(DP_OP_424J2_126_3477_n469), .B(
        DP_OP_424J2_126_3477_n564), .CI(DP_OP_424J2_126_3477_n562), .CO(
        DP_OP_424J2_126_3477_n450), .S(DP_OP_424J2_126_3477_n451) );
  FADDX1_HVT DP_OP_424J2_126_3477_U406 ( .A(DP_OP_424J2_126_3477_n467), .B(
        DP_OP_424J2_126_3477_n465), .CI(DP_OP_424J2_126_3477_n463), .CO(
        DP_OP_424J2_126_3477_n448), .S(DP_OP_424J2_126_3477_n449) );
  FADDX1_HVT DP_OP_424J2_126_3477_U405 ( .A(DP_OP_424J2_126_3477_n560), .B(
        DP_OP_424J2_126_3477_n558), .CI(DP_OP_424J2_126_3477_n461), .CO(
        DP_OP_424J2_126_3477_n446), .S(DP_OP_424J2_126_3477_n447) );
  FADDX1_HVT DP_OP_424J2_126_3477_U404 ( .A(DP_OP_424J2_126_3477_n556), .B(
        DP_OP_424J2_126_3477_n459), .CI(DP_OP_424J2_126_3477_n554), .CO(
        DP_OP_424J2_126_3477_n444), .S(DP_OP_424J2_126_3477_n445) );
  FADDX1_HVT DP_OP_424J2_126_3477_U403 ( .A(DP_OP_424J2_126_3477_n552), .B(
        DP_OP_424J2_126_3477_n457), .CI(DP_OP_424J2_126_3477_n550), .CO(
        DP_OP_424J2_126_3477_n442), .S(DP_OP_424J2_126_3477_n443) );
  FADDX1_HVT DP_OP_424J2_126_3477_U402 ( .A(DP_OP_424J2_126_3477_n548), .B(
        DP_OP_424J2_126_3477_n455), .CI(DP_OP_424J2_126_3477_n453), .CO(
        DP_OP_424J2_126_3477_n440), .S(DP_OP_424J2_126_3477_n441) );
  FADDX1_HVT DP_OP_424J2_126_3477_U401 ( .A(DP_OP_424J2_126_3477_n546), .B(
        DP_OP_424J2_126_3477_n451), .CI(DP_OP_424J2_126_3477_n544), .CO(
        DP_OP_424J2_126_3477_n438), .S(DP_OP_424J2_126_3477_n439) );
  FADDX1_HVT DP_OP_424J2_126_3477_U400 ( .A(DP_OP_424J2_126_3477_n449), .B(
        DP_OP_424J2_126_3477_n542), .CI(DP_OP_424J2_126_3477_n540), .CO(
        DP_OP_424J2_126_3477_n436), .S(DP_OP_424J2_126_3477_n437) );
  FADDX1_HVT DP_OP_424J2_126_3477_U399 ( .A(DP_OP_424J2_126_3477_n447), .B(
        DP_OP_424J2_126_3477_n538), .CI(DP_OP_424J2_126_3477_n445), .CO(
        DP_OP_424J2_126_3477_n434), .S(DP_OP_424J2_126_3477_n435) );
  FADDX1_HVT DP_OP_424J2_126_3477_U398 ( .A(DP_OP_424J2_126_3477_n536), .B(
        DP_OP_424J2_126_3477_n443), .CI(DP_OP_424J2_126_3477_n534), .CO(
        DP_OP_424J2_126_3477_n432), .S(DP_OP_424J2_126_3477_n433) );
  FADDX1_HVT DP_OP_424J2_126_3477_U397 ( .A(DP_OP_424J2_126_3477_n441), .B(
        DP_OP_424J2_126_3477_n532), .CI(DP_OP_424J2_126_3477_n439), .CO(
        DP_OP_424J2_126_3477_n430), .S(DP_OP_424J2_126_3477_n431) );
  FADDX1_HVT DP_OP_424J2_126_3477_U396 ( .A(DP_OP_424J2_126_3477_n530), .B(
        DP_OP_424J2_126_3477_n437), .CI(DP_OP_424J2_126_3477_n528), .CO(
        DP_OP_424J2_126_3477_n428), .S(DP_OP_424J2_126_3477_n429) );
  FADDX1_HVT DP_OP_424J2_126_3477_U395 ( .A(DP_OP_424J2_126_3477_n435), .B(
        DP_OP_424J2_126_3477_n526), .CI(DP_OP_424J2_126_3477_n433), .CO(
        DP_OP_424J2_126_3477_n426), .S(DP_OP_424J2_126_3477_n427) );
  FADDX1_HVT DP_OP_424J2_126_3477_U394 ( .A(DP_OP_424J2_126_3477_n524), .B(
        DP_OP_424J2_126_3477_n431), .CI(DP_OP_424J2_126_3477_n522), .CO(
        DP_OP_424J2_126_3477_n424), .S(DP_OP_424J2_126_3477_n425) );
  FADDX1_HVT DP_OP_424J2_126_3477_U393 ( .A(DP_OP_424J2_126_3477_n429), .B(
        DP_OP_424J2_126_3477_n520), .CI(DP_OP_424J2_126_3477_n427), .CO(
        DP_OP_424J2_126_3477_n422), .S(DP_OP_424J2_126_3477_n423) );
  FADDX1_HVT DP_OP_424J2_126_3477_U392 ( .A(DP_OP_424J2_126_3477_n518), .B(
        DP_OP_424J2_126_3477_n425), .CI(DP_OP_424J2_126_3477_n516), .CO(
        DP_OP_424J2_126_3477_n420), .S(DP_OP_424J2_126_3477_n421) );
  FADDX1_HVT DP_OP_424J2_126_3477_U390 ( .A(DP_OP_424J2_126_3477_n1926), .B(
        DP_OP_424J2_126_3477_n510), .CI(DP_OP_424J2_126_3477_n508), .CO(
        DP_OP_424J2_126_3477_n416), .S(DP_OP_424J2_126_3477_n417) );
  FADDX1_HVT DP_OP_424J2_126_3477_U389 ( .A(DP_OP_424J2_126_3477_n498), .B(
        DP_OP_424J2_126_3477_n494), .CI(DP_OP_424J2_126_3477_n506), .CO(
        DP_OP_424J2_126_3477_n414), .S(DP_OP_424J2_126_3477_n415) );
  FADDX1_HVT DP_OP_424J2_126_3477_U388 ( .A(DP_OP_424J2_126_3477_n504), .B(
        DP_OP_424J2_126_3477_n502), .CI(DP_OP_424J2_126_3477_n500), .CO(
        DP_OP_424J2_126_3477_n412), .S(DP_OP_424J2_126_3477_n413) );
  FADDX1_HVT DP_OP_424J2_126_3477_U387 ( .A(DP_OP_424J2_126_3477_n496), .B(
        DP_OP_424J2_126_3477_n492), .CI(DP_OP_424J2_126_3477_n490), .CO(
        DP_OP_424J2_126_3477_n410), .S(DP_OP_424J2_126_3477_n411) );
  FADDX1_HVT DP_OP_424J2_126_3477_U386 ( .A(DP_OP_424J2_126_3477_n488), .B(
        DP_OP_424J2_126_3477_n486), .CI(DP_OP_424J2_126_3477_n484), .CO(
        DP_OP_424J2_126_3477_n408), .S(DP_OP_424J2_126_3477_n409) );
  FADDX1_HVT DP_OP_424J2_126_3477_U385 ( .A(DP_OP_424J2_126_3477_n482), .B(
        DP_OP_424J2_126_3477_n417), .CI(DP_OP_424J2_126_3477_n480), .CO(
        DP_OP_424J2_126_3477_n406), .S(DP_OP_424J2_126_3477_n407) );
  FADDX1_HVT DP_OP_424J2_126_3477_U384 ( .A(DP_OP_424J2_126_3477_n478), .B(
        DP_OP_424J2_126_3477_n413), .CI(DP_OP_424J2_126_3477_n415), .CO(
        DP_OP_424J2_126_3477_n404), .S(DP_OP_424J2_126_3477_n405) );
  FADDX1_HVT DP_OP_424J2_126_3477_U383 ( .A(DP_OP_424J2_126_3477_n476), .B(
        DP_OP_424J2_126_3477_n474), .CI(DP_OP_424J2_126_3477_n472), .CO(
        DP_OP_424J2_126_3477_n402), .S(DP_OP_424J2_126_3477_n403) );
  FADDX1_HVT DP_OP_424J2_126_3477_U382 ( .A(DP_OP_424J2_126_3477_n470), .B(
        DP_OP_424J2_126_3477_n411), .CI(DP_OP_424J2_126_3477_n468), .CO(
        DP_OP_424J2_126_3477_n400), .S(DP_OP_424J2_126_3477_n401) );
  FADDX1_HVT DP_OP_424J2_126_3477_U381 ( .A(DP_OP_424J2_126_3477_n466), .B(
        DP_OP_424J2_126_3477_n409), .CI(DP_OP_424J2_126_3477_n464), .CO(
        DP_OP_424J2_126_3477_n398), .S(DP_OP_424J2_126_3477_n399) );
  FADDX1_HVT DP_OP_424J2_126_3477_U380 ( .A(DP_OP_424J2_126_3477_n462), .B(
        DP_OP_424J2_126_3477_n407), .CI(DP_OP_424J2_126_3477_n460), .CO(
        DP_OP_424J2_126_3477_n396), .S(DP_OP_424J2_126_3477_n397) );
  FADDX1_HVT DP_OP_424J2_126_3477_U379 ( .A(DP_OP_424J2_126_3477_n405), .B(
        DP_OP_424J2_126_3477_n458), .CI(DP_OP_424J2_126_3477_n456), .CO(
        DP_OP_424J2_126_3477_n394), .S(DP_OP_424J2_126_3477_n395) );
  FADDX1_HVT DP_OP_424J2_126_3477_U378 ( .A(DP_OP_424J2_126_3477_n403), .B(
        DP_OP_424J2_126_3477_n454), .CI(DP_OP_424J2_126_3477_n452), .CO(
        DP_OP_424J2_126_3477_n392), .S(DP_OP_424J2_126_3477_n393) );
  FADDX1_HVT DP_OP_424J2_126_3477_U377 ( .A(DP_OP_424J2_126_3477_n401), .B(
        DP_OP_424J2_126_3477_n450), .CI(DP_OP_424J2_126_3477_n399), .CO(
        DP_OP_424J2_126_3477_n390), .S(DP_OP_424J2_126_3477_n391) );
  FADDX1_HVT DP_OP_424J2_126_3477_U376 ( .A(DP_OP_424J2_126_3477_n448), .B(
        DP_OP_424J2_126_3477_n397), .CI(DP_OP_424J2_126_3477_n446), .CO(
        DP_OP_424J2_126_3477_n388), .S(DP_OP_424J2_126_3477_n389) );
  FADDX1_HVT DP_OP_424J2_126_3477_U375 ( .A(DP_OP_424J2_126_3477_n444), .B(
        DP_OP_424J2_126_3477_n395), .CI(DP_OP_424J2_126_3477_n442), .CO(
        DP_OP_424J2_126_3477_n386), .S(DP_OP_424J2_126_3477_n387) );
  FADDX1_HVT DP_OP_424J2_126_3477_U374 ( .A(DP_OP_424J2_126_3477_n393), .B(
        DP_OP_424J2_126_3477_n440), .CI(DP_OP_424J2_126_3477_n438), .CO(
        DP_OP_424J2_126_3477_n384), .S(DP_OP_424J2_126_3477_n385) );
  FADDX1_HVT DP_OP_424J2_126_3477_U373 ( .A(DP_OP_424J2_126_3477_n391), .B(
        DP_OP_424J2_126_3477_n436), .CI(DP_OP_424J2_126_3477_n389), .CO(
        DP_OP_424J2_126_3477_n382), .S(DP_OP_424J2_126_3477_n383) );
  FADDX1_HVT DP_OP_424J2_126_3477_U372 ( .A(DP_OP_424J2_126_3477_n434), .B(
        DP_OP_424J2_126_3477_n387), .CI(DP_OP_424J2_126_3477_n432), .CO(
        DP_OP_424J2_126_3477_n380), .S(DP_OP_424J2_126_3477_n381) );
  FADDX1_HVT DP_OP_424J2_126_3477_U370 ( .A(DP_OP_424J2_126_3477_n428), .B(
        DP_OP_424J2_126_3477_n381), .CI(DP_OP_424J2_126_3477_n426), .CO(
        DP_OP_424J2_126_3477_n376), .S(DP_OP_424J2_126_3477_n377) );
  FADDX1_HVT DP_OP_424J2_126_3477_U368 ( .A(DP_OP_424J2_126_3477_n377), .B(
        DP_OP_424J2_126_3477_n420), .CI(DP_OP_424J2_126_3477_n375), .CO(
        DP_OP_424J2_126_3477_n372), .S(DP_OP_424J2_126_3477_n373) );
  FADDX1_HVT DP_OP_424J2_126_3477_U367 ( .A(DP_OP_424J2_126_3477_n1925), .B(
        DP_OP_424J2_126_3477_n416), .CI(DP_OP_424J2_126_3477_n414), .CO(
        DP_OP_424J2_126_3477_n370), .S(DP_OP_424J2_126_3477_n371) );
  FADDX1_HVT DP_OP_424J2_126_3477_U366 ( .A(DP_OP_424J2_126_3477_n412), .B(
        DP_OP_424J2_126_3477_n410), .CI(DP_OP_424J2_126_3477_n408), .CO(
        DP_OP_424J2_126_3477_n368), .S(DP_OP_424J2_126_3477_n369) );
  FADDX1_HVT DP_OP_424J2_126_3477_U365 ( .A(DP_OP_424J2_126_3477_n406), .B(
        DP_OP_424J2_126_3477_n371), .CI(DP_OP_424J2_126_3477_n404), .CO(
        DP_OP_424J2_126_3477_n366), .S(DP_OP_424J2_126_3477_n367) );
  FADDX1_HVT DP_OP_424J2_126_3477_U364 ( .A(DP_OP_424J2_126_3477_n402), .B(
        DP_OP_424J2_126_3477_n400), .CI(DP_OP_424J2_126_3477_n369), .CO(
        DP_OP_424J2_126_3477_n364), .S(DP_OP_424J2_126_3477_n365) );
  FADDX1_HVT DP_OP_424J2_126_3477_U363 ( .A(DP_OP_424J2_126_3477_n398), .B(
        DP_OP_424J2_126_3477_n396), .CI(DP_OP_424J2_126_3477_n367), .CO(
        DP_OP_424J2_126_3477_n362), .S(DP_OP_424J2_126_3477_n363) );
  FADDX1_HVT DP_OP_424J2_126_3477_U362 ( .A(DP_OP_424J2_126_3477_n394), .B(
        DP_OP_424J2_126_3477_n392), .CI(DP_OP_424J2_126_3477_n365), .CO(
        DP_OP_424J2_126_3477_n360), .S(DP_OP_424J2_126_3477_n361) );
  FADDX1_HVT DP_OP_424J2_126_3477_U361 ( .A(DP_OP_424J2_126_3477_n390), .B(
        DP_OP_424J2_126_3477_n363), .CI(DP_OP_424J2_126_3477_n388), .CO(
        DP_OP_424J2_126_3477_n358), .S(DP_OP_424J2_126_3477_n359) );
  FADDX1_HVT DP_OP_424J2_126_3477_U360 ( .A(DP_OP_424J2_126_3477_n386), .B(
        DP_OP_424J2_126_3477_n361), .CI(DP_OP_424J2_126_3477_n384), .CO(
        DP_OP_424J2_126_3477_n356), .S(DP_OP_424J2_126_3477_n357) );
  FADDX1_HVT DP_OP_424J2_126_3477_U359 ( .A(DP_OP_424J2_126_3477_n382), .B(
        DP_OP_424J2_126_3477_n359), .CI(DP_OP_424J2_126_3477_n380), .CO(
        DP_OP_424J2_126_3477_n354), .S(DP_OP_424J2_126_3477_n355) );
  FADDX1_HVT DP_OP_424J2_126_3477_U358 ( .A(DP_OP_424J2_126_3477_n357), .B(
        DP_OP_424J2_126_3477_n378), .CI(DP_OP_424J2_126_3477_n355), .CO(
        DP_OP_424J2_126_3477_n352), .S(DP_OP_424J2_126_3477_n353) );
  FADDX1_HVT DP_OP_424J2_126_3477_U357 ( .A(DP_OP_424J2_126_3477_n376), .B(
        DP_OP_424J2_126_3477_n374), .CI(DP_OP_424J2_126_3477_n353), .CO(
        DP_OP_424J2_126_3477_n350), .S(DP_OP_424J2_126_3477_n351) );
  FADDX1_HVT DP_OP_424J2_126_3477_U356 ( .A(DP_OP_424J2_126_3477_n1924), .B(
        DP_OP_424J2_126_3477_n370), .CI(DP_OP_424J2_126_3477_n368), .CO(
        DP_OP_424J2_126_3477_n348), .S(DP_OP_424J2_126_3477_n349) );
  FADDX1_HVT DP_OP_424J2_126_3477_U355 ( .A(DP_OP_424J2_126_3477_n366), .B(
        DP_OP_424J2_126_3477_n349), .CI(DP_OP_424J2_126_3477_n364), .CO(
        DP_OP_424J2_126_3477_n346), .S(DP_OP_424J2_126_3477_n347) );
  FADDX1_HVT DP_OP_424J2_126_3477_U354 ( .A(DP_OP_424J2_126_3477_n362), .B(
        DP_OP_424J2_126_3477_n360), .CI(DP_OP_424J2_126_3477_n347), .CO(
        DP_OP_424J2_126_3477_n344), .S(DP_OP_424J2_126_3477_n345) );
  FADDX1_HVT DP_OP_424J2_126_3477_U353 ( .A(DP_OP_424J2_126_3477_n358), .B(
        DP_OP_424J2_126_3477_n345), .CI(DP_OP_424J2_126_3477_n356), .CO(
        DP_OP_424J2_126_3477_n342), .S(DP_OP_424J2_126_3477_n343) );
  FADDX1_HVT DP_OP_424J2_126_3477_U352 ( .A(DP_OP_424J2_126_3477_n354), .B(
        DP_OP_424J2_126_3477_n343), .CI(DP_OP_424J2_126_3477_n352), .CO(
        DP_OP_424J2_126_3477_n340), .S(DP_OP_424J2_126_3477_n341) );
  FADDX1_HVT DP_OP_424J2_126_3477_U350 ( .A(DP_OP_424J2_126_3477_n339), .B(
        DP_OP_424J2_126_3477_n348), .CI(DP_OP_424J2_126_3477_n346), .CO(
        DP_OP_424J2_126_3477_n336), .S(DP_OP_424J2_126_3477_n337) );
  FADDX1_HVT DP_OP_424J2_126_3477_U349 ( .A(DP_OP_424J2_126_3477_n337), .B(
        DP_OP_424J2_126_3477_n344), .CI(DP_OP_424J2_126_3477_n342), .CO(
        DP_OP_424J2_126_3477_n334), .S(DP_OP_424J2_126_3477_n335) );
  FADDX1_HVT DP_OP_424J2_126_3477_U348 ( .A(DP_OP_424J2_126_3477_n1923), .B(
        DP_OP_424J2_126_3477_n338), .CI(DP_OP_424J2_126_3477_n336), .CO(
        DP_OP_424J2_126_3477_n332), .S(DP_OP_424J2_126_3477_n333) );
  FADDX1_HVT DP_OP_424J2_126_3477_U331 ( .A(DP_OP_424J2_126_3477_n1903), .B(
        DP_OP_424J2_126_3477_n1901), .CI(DP_OP_424J2_126_3477_n1899), .CO(
        DP_OP_424J2_126_3477_n269), .S(n_conv2_sum_c[0]) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U330 ( .A1(DP_OP_424J2_126_3477_n1837), 
        .A2(DP_OP_424J2_126_3477_n1839), .Y(DP_OP_424J2_126_3477_n268) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U329 ( .A1(DP_OP_424J2_126_3477_n1839), .A2(
        DP_OP_424J2_126_3477_n1837), .Y(DP_OP_424J2_126_3477_n267) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U323 ( .A1(DP_OP_424J2_126_3477_n1731), 
        .A2(DP_OP_424J2_126_3477_n1733), .Y(DP_OP_424J2_126_3477_n265) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U315 ( .A1(DP_OP_424J2_126_3477_n1577), 
        .A2(DP_OP_424J2_126_3477_n1579), .Y(DP_OP_424J2_126_3477_n260) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U309 ( .A1(DP_OP_424J2_126_3477_n1401), 
        .A2(DP_OP_424J2_126_3477_n1403), .Y(DP_OP_424J2_126_3477_n257) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U301 ( .A1(DP_OP_424J2_126_3477_n1213), 
        .A2(DP_OP_424J2_126_3477_n1215), .Y(DP_OP_424J2_126_3477_n252) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U274 ( .A1(DP_OP_424J2_126_3477_n513), .A2(
        DP_OP_424J2_126_3477_n648), .Y(DP_OP_424J2_126_3477_n237) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U235 ( .A1(DP_OP_424J2_126_3477_n350), .A2(
        DP_OP_424J2_126_3477_n341), .Y(DP_OP_424J2_126_3477_n210) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U234 ( .A1(DP_OP_424J2_126_3477_n341), .A2(
        DP_OP_424J2_126_3477_n350), .Y(DP_OP_424J2_126_3477_n209) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U225 ( .A1(DP_OP_424J2_126_3477_n340), .A2(
        DP_OP_424J2_126_3477_n335), .Y(DP_OP_424J2_126_3477_n203) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U217 ( .A1(DP_OP_424J2_126_3477_n334), .A2(
        DP_OP_424J2_126_3477_n333), .Y(DP_OP_424J2_126_3477_n198) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U216 ( .A1(DP_OP_424J2_126_3477_n333), .A2(
        DP_OP_424J2_126_3477_n334), .Y(DP_OP_424J2_126_3477_n197) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U214 ( .A1(DP_OP_424J2_126_3477_n286), .A2(
        DP_OP_424J2_126_3477_n198), .Y(DP_OP_424J2_126_3477_n22) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U210 ( .A1(DP_OP_424J2_126_3477_n287), .A2(
        DP_OP_424J2_126_3477_n286), .Y(DP_OP_424J2_126_3477_n189) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U201 ( .A1(DP_OP_424J2_126_3477_n332), .A2(
        DP_OP_424J2_126_3477_n331), .Y(DP_OP_424J2_126_3477_n185) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U194 ( .A1(DP_OP_424J2_126_3477_n182), .A2(
        DP_OP_424J2_126_3477_n189), .Y(DP_OP_424J2_126_3477_n176) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U187 ( .A1(DP_OP_424J2_126_3477_n329), .A2(
        DP_OP_424J2_126_3477_n330), .Y(DP_OP_424J2_126_3477_n174) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U186 ( .A1(DP_OP_424J2_126_3477_n330), .A2(
        DP_OP_424J2_126_3477_n329), .Y(DP_OP_424J2_126_3477_n171) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U177 ( .A1(DP_OP_424J2_126_3477_n327), .A2(
        DP_OP_424J2_126_3477_n328), .Y(DP_OP_424J2_126_3477_n167) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U176 ( .A1(DP_OP_424J2_126_3477_n328), .A2(
        DP_OP_424J2_126_3477_n327), .Y(DP_OP_424J2_126_3477_n166) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U172 ( .A1(DP_OP_424J2_126_3477_n166), .A2(
        DP_OP_424J2_126_3477_n171), .Y(DP_OP_424J2_126_3477_n162) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U168 ( .A1(DP_OP_424J2_126_3477_n176), .A2(
        DP_OP_424J2_126_3477_n162), .Y(DP_OP_424J2_126_3477_n160) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U163 ( .A1(DP_OP_424J2_126_3477_n325), .A2(
        DP_OP_424J2_126_3477_n326), .Y(DP_OP_424J2_126_3477_n156) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U162 ( .A1(DP_OP_424J2_126_3477_n326), .A2(
        DP_OP_424J2_126_3477_n325), .Y(DP_OP_424J2_126_3477_n153) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U153 ( .A1(DP_OP_424J2_126_3477_n323), .A2(
        DP_OP_424J2_126_3477_n324), .Y(DP_OP_424J2_126_3477_n149) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U152 ( .A1(DP_OP_424J2_126_3477_n324), .A2(
        DP_OP_424J2_126_3477_n323), .Y(DP_OP_424J2_126_3477_n148) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U150 ( .A1(DP_OP_424J2_126_3477_n281), .A2(
        DP_OP_424J2_126_3477_n149), .Y(DP_OP_424J2_126_3477_n17) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U148 ( .A1(DP_OP_424J2_126_3477_n148), .A2(
        DP_OP_424J2_126_3477_n153), .Y(DP_OP_424J2_126_3477_n146) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U146 ( .A1(DP_OP_424J2_126_3477_n162), .A2(
        DP_OP_424J2_126_3477_n146), .Y(DP_OP_424J2_126_3477_n144) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U142 ( .A1(DP_OP_424J2_126_3477_n176), .A2(
        DP_OP_424J2_126_3477_n142), .Y(DP_OP_424J2_126_3477_n140) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U137 ( .A1(n1380), .A2(
        DP_OP_424J2_126_3477_n322), .Y(DP_OP_424J2_126_3477_n136) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U136 ( .A1(DP_OP_424J2_126_3477_n322), .A2(
        n1380), .Y(DP_OP_424J2_126_3477_n133) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U127 ( .A1(DP_OP_424J2_126_3477_n319), .A2(
        DP_OP_424J2_126_3477_n320), .Y(DP_OP_424J2_126_3477_n129) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U126 ( .A1(DP_OP_424J2_126_3477_n320), .A2(
        DP_OP_424J2_126_3477_n319), .Y(DP_OP_424J2_126_3477_n128) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U124 ( .A1(DP_OP_424J2_126_3477_n279), .A2(
        DP_OP_424J2_126_3477_n129), .Y(DP_OP_424J2_126_3477_n15) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U122 ( .A1(DP_OP_424J2_126_3477_n128), .A2(
        DP_OP_424J2_126_3477_n133), .Y(DP_OP_424J2_126_3477_n126) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U115 ( .A1(DP_OP_424J2_126_3477_n317), .A2(
        DP_OP_424J2_126_3477_n318), .Y(DP_OP_424J2_126_3477_n120) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U108 ( .A1(DP_OP_424J2_126_3477_n126), .A2(
        n1764), .Y(DP_OP_424J2_126_3477_n115) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U102 ( .A1(DP_OP_424J2_126_3477_n176), .A2(
        DP_OP_424J2_126_3477_n111), .Y(DP_OP_424J2_126_3477_n109) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U97 ( .A1(DP_OP_424J2_126_3477_n315), .A2(
        DP_OP_424J2_126_3477_n316), .Y(DP_OP_424J2_126_3477_n105) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U96 ( .A1(DP_OP_424J2_126_3477_n316), .A2(
        DP_OP_424J2_126_3477_n315), .Y(DP_OP_424J2_126_3477_n102) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U94 ( .A1(DP_OP_424J2_126_3477_n277), .A2(
        DP_OP_424J2_126_3477_n105), .Y(DP_OP_424J2_126_3477_n13) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U87 ( .A1(DP_OP_424J2_126_3477_n313), .A2(
        DP_OP_424J2_126_3477_n314), .Y(DP_OP_424J2_126_3477_n98) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U86 ( .A1(DP_OP_424J2_126_3477_n314), .A2(
        DP_OP_424J2_126_3477_n313), .Y(DP_OP_424J2_126_3477_n97) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U82 ( .A1(DP_OP_424J2_126_3477_n97), .A2(
        DP_OP_424J2_126_3477_n102), .Y(DP_OP_424J2_126_3477_n95) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U75 ( .A1(DP_OP_424J2_126_3477_n311), .A2(
        DP_OP_424J2_126_3477_n312), .Y(DP_OP_424J2_126_3477_n89) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U68 ( .A1(DP_OP_424J2_126_3477_n95), .A2(
        n1763), .Y(DP_OP_424J2_126_3477_n82) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U61 ( .A1(DP_OP_424J2_126_3477_n309), .A2(
        DP_OP_424J2_126_3477_n310), .Y(DP_OP_424J2_126_3477_n78) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U60 ( .A1(DP_OP_424J2_126_3477_n310), .A2(
        DP_OP_424J2_126_3477_n309), .Y(DP_OP_424J2_126_3477_n77) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U54 ( .A1(DP_OP_424J2_126_3477_n111), .A2(
        DP_OP_424J2_126_3477_n75), .Y(DP_OP_424J2_126_3477_n73) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U45 ( .A1(DP_OP_424J2_126_3477_n307), .A2(
        DP_OP_424J2_126_3477_n308), .Y(DP_OP_424J2_126_3477_n65) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U38 ( .A1(DP_OP_424J2_126_3477_n71), .A2(
        n1759), .Y(DP_OP_424J2_126_3477_n60) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U34 ( .A1(DP_OP_424J2_126_3477_n287), .A2(
        DP_OP_424J2_126_3477_n58), .Y(DP_OP_424J2_126_3477_n56) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U29 ( .A1(DP_OP_424J2_126_3477_n305), .A2(
        DP_OP_424J2_126_3477_n306), .Y(DP_OP_424J2_126_3477_n52) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U28 ( .A1(DP_OP_424J2_126_3477_n306), .A2(
        DP_OP_424J2_126_3477_n305), .Y(DP_OP_424J2_126_3477_n51) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U21 ( .A1(DP_OP_424J2_126_3477_n303), .A2(
        DP_OP_424J2_126_3477_n304), .Y(DP_OP_424J2_126_3477_n47) );
  NAND2X0_HVT DP_OP_424J2_126_3477_U9 ( .A1(n1757), .A2(
        DP_OP_424J2_126_3477_n302), .Y(DP_OP_424J2_126_3477_n38) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U325 ( .A1(DP_OP_423J2_125_3477_n5), .A2(
        DP_OP_423J2_125_3477_n267), .A3(DP_OP_423J2_125_3477_n268), .Y(
        DP_OP_423J2_125_3477_n266) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U173 ( .A1(DP_OP_423J2_125_3477_n174), .A2(
        DP_OP_423J2_125_3477_n166), .A3(DP_OP_423J2_125_3477_n167), .Y(
        DP_OP_423J2_125_3477_n165) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1161 ( .A1(n1977), .A2(n1508), .Y(
        DP_OP_423J2_125_3477_n338) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U83 ( .A1(DP_OP_423J2_125_3477_n105), .A2(
        DP_OP_423J2_125_3477_n97), .A3(DP_OP_423J2_125_3477_n98), .Y(
        DP_OP_423J2_125_3477_n96) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U123 ( .A1(DP_OP_423J2_125_3477_n136), .A2(
        DP_OP_423J2_125_3477_n128), .A3(DP_OP_423J2_125_3477_n129), .Y(
        DP_OP_423J2_125_3477_n127) );
  XNOR2X1_HVT DP_OP_423J2_125_3477_U787 ( .A1(DP_OP_423J2_125_3477_n2502), 
        .A2(DP_OP_423J2_125_3477_n3029), .Y(DP_OP_423J2_125_3477_n1211) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2291 ( .A1(DP_OP_425J2_127_3477_n2092), 
        .A2(n34), .Y(DP_OP_423J2_125_3477_n3050) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2290 ( .A1(DP_OP_423J2_125_3477_n3057), 
        .A2(n34), .Y(DP_OP_423J2_125_3477_n3049) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2289 ( .A1(DP_OP_423J2_125_3477_n3056), .A2(
        n34), .Y(DP_OP_423J2_125_3477_n3048) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2283 ( .A1(DP_OP_425J2_127_3477_n2092), 
        .A2(DP_OP_424J2_126_3477_n3066), .Y(DP_OP_423J2_125_3477_n3042) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2282 ( .A1(DP_OP_423J2_125_3477_n3057), 
        .A2(DP_OP_424J2_126_3477_n3066), .Y(DP_OP_423J2_125_3477_n3041) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2274 ( .A1(DP_OP_423J2_125_3477_n3057), 
        .A2(DP_OP_423J2_125_3477_n3065), .Y(DP_OP_423J2_125_3477_n3033) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2273 ( .A1(DP_OP_423J2_125_3477_n3056), .A2(
        DP_OP_423J2_125_3477_n3065), .Y(DP_OP_423J2_125_3477_n3032) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2272 ( .A1(DP_OP_423J2_125_3477_n3063), .A2(
        n215), .Y(DP_OP_423J2_125_3477_n1728) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2271 ( .A1(DP_OP_423J2_125_3477_n3062), .A2(
        n215), .Y(DP_OP_423J2_125_3477_n3031) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2270 ( .A1(DP_OP_423J2_125_3477_n3061), .A2(
        n215), .Y(DP_OP_423J2_125_3477_n3030) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2268 ( .A1(DP_OP_423J2_125_3477_n3059), .A2(
        n215), .Y(DP_OP_423J2_125_3477_n3028) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2267 ( .A1(DP_OP_425J2_127_3477_n2092), .A2(
        n213), .Y(DP_OP_423J2_125_3477_n820) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2266 ( .A1(DP_OP_423J2_125_3477_n3057), .A2(
        n215), .Y(DP_OP_423J2_125_3477_n3027) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2265 ( .A1(DP_OP_423J2_125_3477_n3056), 
        .A2(n215), .Y(DP_OP_423J2_125_3477_n3026) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2245 ( .A1(DP_OP_423J2_125_3477_n3014), .A2(
        DP_OP_423J2_125_3477_n3025), .Y(DP_OP_423J2_125_3477_n3006) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2238 ( .A1(DP_OP_424J2_126_3477_n2927), 
        .A2(n704), .Y(DP_OP_423J2_125_3477_n2999) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2237 ( .A1(DP_OP_423J2_125_3477_n3014), .A2(
        n699), .Y(DP_OP_423J2_125_3477_n2998) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2231 ( .A1(DP_OP_424J2_126_3477_n2928), 
        .A2(DP_OP_425J2_127_3477_n3023), .Y(DP_OP_423J2_125_3477_n2992) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2229 ( .A1(DP_OP_423J2_125_3477_n3014), .A2(
        DP_OP_424J2_126_3477_n3023), .Y(DP_OP_423J2_125_3477_n2990) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2208 ( .A1(DP_OP_424J2_126_3477_n2889), 
        .A2(n677), .Y(DP_OP_423J2_125_3477_n2969) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2207 ( .A1(DP_OP_423J2_125_3477_n2976), 
        .A2(n674), .Y(DP_OP_423J2_125_3477_n2968) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2206 ( .A1(DP_OP_422J2_124_3477_n2051), 
        .A2(n677), .Y(DP_OP_423J2_125_3477_n2967) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2205 ( .A1(DP_OP_425J2_127_3477_n2182), 
        .A2(n677), .Y(DP_OP_423J2_125_3477_n2966) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2204 ( .A1(DP_OP_423J2_125_3477_n2973), 
        .A2(n677), .Y(DP_OP_423J2_125_3477_n2965) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2203 ( .A1(DP_OP_422J2_124_3477_n2048), 
        .A2(n677), .Y(DP_OP_423J2_125_3477_n2964) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2202 ( .A1(DP_OP_424J2_126_3477_n2883), 
        .A2(n677), .Y(DP_OP_423J2_125_3477_n2963) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2201 ( .A1(DP_OP_424J2_126_3477_n2882), .A2(
        n677), .Y(DP_OP_423J2_125_3477_n2962) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2200 ( .A1(DP_OP_425J2_127_3477_n2185), 
        .A2(DP_OP_422J2_124_3477_n2980), .Y(DP_OP_423J2_125_3477_n2961) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2199 ( .A1(DP_OP_423J2_125_3477_n2976), 
        .A2(DP_OP_424J2_126_3477_n2980), .Y(DP_OP_423J2_125_3477_n2960) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2198 ( .A1(DP_OP_422J2_124_3477_n2051), 
        .A2(DP_OP_422J2_124_3477_n2980), .Y(DP_OP_423J2_125_3477_n2959) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2197 ( .A1(DP_OP_425J2_127_3477_n2182), 
        .A2(DP_OP_424J2_126_3477_n2980), .Y(DP_OP_423J2_125_3477_n2958) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2196 ( .A1(DP_OP_423J2_125_3477_n2973), 
        .A2(DP_OP_424J2_126_3477_n2980), .Y(DP_OP_423J2_125_3477_n2957) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2195 ( .A1(DP_OP_422J2_124_3477_n2048), 
        .A2(DP_OP_425J2_127_3477_n2980), .Y(DP_OP_423J2_125_3477_n2956) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2194 ( .A1(DP_OP_424J2_126_3477_n2883), 
        .A2(DP_OP_425J2_127_3477_n2980), .Y(DP_OP_423J2_125_3477_n2955) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2193 ( .A1(DP_OP_424J2_126_3477_n2882), .A2(
        DP_OP_425J2_127_3477_n2980), .Y(DP_OP_423J2_125_3477_n2954) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2186 ( .A1(DP_OP_424J2_126_3477_n2883), 
        .A2(DP_OP_424J2_126_3477_n2979), .Y(DP_OP_423J2_125_3477_n2947) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2185 ( .A1(DP_OP_424J2_126_3477_n2882), .A2(
        DP_OP_424J2_126_3477_n2979), .Y(DP_OP_423J2_125_3477_n2946) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2183 ( .A1(DP_OP_423J2_125_3477_n2976), .A2(
        n663), .Y(DP_OP_423J2_125_3477_n2944) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2177 ( .A1(DP_OP_424J2_126_3477_n2882), 
        .A2(n663), .Y(DP_OP_423J2_125_3477_n2938) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2158 ( .A1(DP_OP_422J2_124_3477_n2091), 
        .A2(n445), .Y(DP_OP_423J2_125_3477_n2919) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2157 ( .A1(DP_OP_422J2_124_3477_n2090), .A2(
        n446), .Y(DP_OP_423J2_125_3477_n2918) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2150 ( .A1(DP_OP_422J2_124_3477_n2091), 
        .A2(DP_OP_423J2_125_3477_n2936), .Y(DP_OP_423J2_125_3477_n2911) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2149 ( .A1(DP_OP_422J2_124_3477_n2090), .A2(
        DP_OP_423J2_125_3477_n2936), .Y(DP_OP_423J2_125_3477_n2910) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2139 ( .A1(DP_OP_423J2_125_3477_n2932), .A2(
        n35), .Y(DP_OP_423J2_125_3477_n2900) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2138 ( .A1(DP_OP_423J2_125_3477_n2931), .A2(
        n35), .Y(DP_OP_423J2_125_3477_n2899) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2137 ( .A1(DP_OP_425J2_127_3477_n2226), .A2(
        n35), .Y(DP_OP_423J2_125_3477_n2898) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2136 ( .A1(DP_OP_422J2_124_3477_n2093), .A2(
        n35), .Y(DP_OP_423J2_125_3477_n2897) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2135 ( .A1(DP_OP_422J2_124_3477_n2092), .A2(
        n35), .Y(DP_OP_423J2_125_3477_n2896) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2134 ( .A1(DP_OP_422J2_124_3477_n2091), .A2(
        n35), .Y(DP_OP_423J2_125_3477_n2895) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2133 ( .A1(DP_OP_422J2_124_3477_n2090), 
        .A2(n35), .Y(DP_OP_423J2_125_3477_n2894) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2114 ( .A1(DP_OP_424J2_126_3477_n2795), 
        .A2(DP_OP_424J2_126_3477_n2893), .Y(DP_OP_423J2_125_3477_n2875) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2113 ( .A1(DP_OP_424J2_126_3477_n2794), .A2(
        DP_OP_425J2_127_3477_n2893), .Y(DP_OP_423J2_125_3477_n2874) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2109 ( .A1(DP_OP_423J2_125_3477_n2886), 
        .A2(DP_OP_423J2_125_3477_n2892), .Y(DP_OP_423J2_125_3477_n2870) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2108 ( .A1(DP_OP_422J2_124_3477_n2137), 
        .A2(DP_OP_423J2_125_3477_n2892), .Y(DP_OP_423J2_125_3477_n2869) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2107 ( .A1(DP_OP_425J2_127_3477_n2268), 
        .A2(DP_OP_423J2_125_3477_n2892), .Y(DP_OP_423J2_125_3477_n2868) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2106 ( .A1(DP_OP_422J2_124_3477_n2135), 
        .A2(DP_OP_423J2_125_3477_n2892), .Y(DP_OP_423J2_125_3477_n2867) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2105 ( .A1(DP_OP_422J2_124_3477_n2134), .A2(
        DP_OP_423J2_125_3477_n2892), .Y(DP_OP_423J2_125_3477_n2866) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2096 ( .A1(DP_OP_423J2_125_3477_n2889), .A2(
        DP_OP_424J2_126_3477_n2890), .Y(DP_OP_423J2_125_3477_n2857) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2095 ( .A1(DP_OP_422J2_124_3477_n2140), .A2(
        DP_OP_424J2_126_3477_n2890), .Y(DP_OP_423J2_125_3477_n2856) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2094 ( .A1(DP_OP_423J2_125_3477_n2887), .A2(
        DP_OP_423J2_125_3477_n2890), .Y(DP_OP_423J2_125_3477_n2855) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2093 ( .A1(DP_OP_423J2_125_3477_n2886), .A2(
        DP_OP_423J2_125_3477_n2890), .Y(DP_OP_423J2_125_3477_n2854) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2092 ( .A1(DP_OP_422J2_124_3477_n2137), .A2(
        DP_OP_424J2_126_3477_n2890), .Y(DP_OP_423J2_125_3477_n2853) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2091 ( .A1(DP_OP_424J2_126_3477_n2796), .A2(
        DP_OP_422J2_124_3477_n2890), .Y(DP_OP_423J2_125_3477_n2852) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2090 ( .A1(DP_OP_422J2_124_3477_n2135), .A2(
        DP_OP_422J2_124_3477_n2890), .Y(DP_OP_423J2_125_3477_n2851) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2089 ( .A1(DP_OP_422J2_124_3477_n2134), 
        .A2(DP_OP_422J2_124_3477_n2890), .Y(DP_OP_423J2_125_3477_n2850) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2075 ( .A1(DP_OP_423J2_125_3477_n2844), 
        .A2(DP_OP_423J2_125_3477_n2849), .Y(DP_OP_423J2_125_3477_n2836) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2074 ( .A1(DP_OP_423J2_125_3477_n2843), 
        .A2(DP_OP_423J2_125_3477_n2849), .Y(DP_OP_423J2_125_3477_n2835) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2073 ( .A1(DP_OP_423J2_125_3477_n2842), 
        .A2(n1428), .Y(DP_OP_423J2_125_3477_n2834) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2072 ( .A1(DP_OP_423J2_125_3477_n2841), 
        .A2(DP_OP_424J2_126_3477_n2849), .Y(DP_OP_423J2_125_3477_n2833) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2070 ( .A1(DP_OP_425J2_127_3477_n2311), 
        .A2(n1428), .Y(DP_OP_423J2_125_3477_n2831) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2052 ( .A1(DP_OP_423J2_125_3477_n2845), .A2(
        DP_OP_422J2_124_3477_n2846), .Y(DP_OP_423J2_125_3477_n2813) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2051 ( .A1(DP_OP_423J2_125_3477_n2844), .A2(
        DP_OP_425J2_127_3477_n2846), .Y(DP_OP_423J2_125_3477_n2812) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2050 ( .A1(DP_OP_423J2_125_3477_n2843), .A2(
        DP_OP_425J2_127_3477_n2846), .Y(DP_OP_423J2_125_3477_n2811) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2049 ( .A1(DP_OP_423J2_125_3477_n2842), .A2(
        DP_OP_425J2_127_3477_n2846), .Y(DP_OP_423J2_125_3477_n2810) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2048 ( .A1(DP_OP_423J2_125_3477_n2841), .A2(
        DP_OP_422J2_124_3477_n2846), .Y(DP_OP_423J2_125_3477_n2809) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2047 ( .A1(DP_OP_425J2_127_3477_n2312), .A2(
        DP_OP_424J2_126_3477_n2846), .Y(DP_OP_423J2_125_3477_n2808) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2046 ( .A1(DP_OP_425J2_127_3477_n2311), .A2(
        DP_OP_422J2_124_3477_n2846), .Y(DP_OP_423J2_125_3477_n2807) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2045 ( .A1(DP_OP_425J2_127_3477_n2310), 
        .A2(DP_OP_424J2_126_3477_n2846), .Y(DP_OP_423J2_125_3477_n2806) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2026 ( .A1(DP_OP_423J2_125_3477_n2795), 
        .A2(DP_OP_423J2_125_3477_n2805), .Y(DP_OP_423J2_125_3477_n2787) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2025 ( .A1(DP_OP_423J2_125_3477_n2794), .A2(
        DP_OP_423J2_125_3477_n2805), .Y(DP_OP_423J2_125_3477_n2786) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2020 ( .A1(DP_OP_422J2_124_3477_n2225), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_423J2_125_3477_n2781) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2017 ( .A1(DP_OP_423J2_125_3477_n2794), .A2(
        DP_OP_423J2_125_3477_n2804), .Y(DP_OP_423J2_125_3477_n2778) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2013 ( .A1(DP_OP_423J2_125_3477_n2798), 
        .A2(n1444), .Y(DP_OP_423J2_125_3477_n2774) );
  OR2X1_HVT DP_OP_423J2_125_3477_U2009 ( .A1(DP_OP_423J2_125_3477_n2794), .A2(
        DP_OP_422J2_124_3477_n2803), .Y(DP_OP_423J2_125_3477_n2770) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1983 ( .A1(DP_OP_422J2_124_3477_n2268), 
        .A2(n66), .Y(DP_OP_423J2_125_3477_n2744) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1982 ( .A1(DP_OP_423J2_125_3477_n2751), 
        .A2(DP_OP_425J2_127_3477_n2761), .Y(DP_OP_423J2_125_3477_n2743) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1981 ( .A1(DP_OP_423J2_125_3477_n2750), .A2(
        n66), .Y(DP_OP_423J2_125_3477_n2742) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1964 ( .A1(DP_OP_423J2_125_3477_n2757), .A2(
        DP_OP_423J2_125_3477_n2758), .Y(DP_OP_423J2_125_3477_n2725) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1963 ( .A1(DP_OP_423J2_125_3477_n2756), .A2(
        DP_OP_423J2_125_3477_n2758), .Y(DP_OP_423J2_125_3477_n2724) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1962 ( .A1(DP_OP_425J2_127_3477_n2403), .A2(
        DP_OP_423J2_125_3477_n2758), .Y(DP_OP_423J2_125_3477_n2723) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1961 ( .A1(DP_OP_423J2_125_3477_n2754), .A2(
        DP_OP_423J2_125_3477_n2758), .Y(DP_OP_423J2_125_3477_n2722) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1960 ( .A1(DP_OP_425J2_127_3477_n2401), .A2(
        DP_OP_423J2_125_3477_n2758), .Y(DP_OP_423J2_125_3477_n2721) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1959 ( .A1(DP_OP_425J2_127_3477_n2400), .A2(
        DP_OP_423J2_125_3477_n2758), .Y(DP_OP_423J2_125_3477_n2720) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1958 ( .A1(DP_OP_423J2_125_3477_n2751), .A2(
        DP_OP_423J2_125_3477_n2758), .Y(DP_OP_423J2_125_3477_n2719) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1957 ( .A1(DP_OP_423J2_125_3477_n2750), 
        .A2(DP_OP_423J2_125_3477_n2758), .Y(DP_OP_423J2_125_3477_n2718) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1938 ( .A1(DP_OP_424J2_126_3477_n2619), 
        .A2(n596), .Y(DP_OP_423J2_125_3477_n2699) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1937 ( .A1(DP_OP_423J2_125_3477_n2706), .A2(
        n597), .Y(DP_OP_423J2_125_3477_n2698) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1930 ( .A1(DP_OP_424J2_126_3477_n2619), 
        .A2(n1340), .Y(DP_OP_423J2_125_3477_n2691) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1929 ( .A1(DP_OP_423J2_125_3477_n2706), .A2(
        n1342), .Y(DP_OP_423J2_125_3477_n2690) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1920 ( .A1(DP_OP_423J2_125_3477_n2713), .A2(
        DP_OP_425J2_127_3477_n2714), .Y(DP_OP_423J2_125_3477_n2681) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1894 ( .A1(DP_OP_424J2_126_3477_n2575), 
        .A2(n1), .Y(DP_OP_423J2_125_3477_n2655) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1893 ( .A1(DP_OP_424J2_126_3477_n2574), .A2(
        DP_OP_422J2_124_3477_n2673), .Y(DP_OP_423J2_125_3477_n2654) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1886 ( .A1(DP_OP_424J2_126_3477_n2575), 
        .A2(n278), .Y(DP_OP_423J2_125_3477_n2647) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1885 ( .A1(DP_OP_424J2_126_3477_n2574), .A2(
        n279), .Y(DP_OP_423J2_125_3477_n2646) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1880 ( .A1(DP_OP_423J2_125_3477_n2665), 
        .A2(n1400), .Y(DP_OP_423J2_125_3477_n2641) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1876 ( .A1(DP_OP_423J2_125_3477_n2669), .A2(
        DP_OP_422J2_124_3477_n2670), .Y(DP_OP_423J2_125_3477_n2637) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1875 ( .A1(DP_OP_423J2_125_3477_n2668), .A2(
        DP_OP_422J2_124_3477_n2670), .Y(DP_OP_423J2_125_3477_n2636) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1874 ( .A1(DP_OP_423J2_125_3477_n2667), .A2(
        DP_OP_422J2_124_3477_n2670), .Y(DP_OP_423J2_125_3477_n2635) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1873 ( .A1(DP_OP_423J2_125_3477_n2666), .A2(
        DP_OP_422J2_124_3477_n2670), .Y(DP_OP_423J2_125_3477_n2634) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1872 ( .A1(DP_OP_423J2_125_3477_n2665), .A2(
        DP_OP_422J2_124_3477_n2670), .Y(DP_OP_423J2_125_3477_n2633) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1871 ( .A1(DP_OP_424J2_126_3477_n2576), .A2(
        n86), .Y(DP_OP_423J2_125_3477_n2632) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1870 ( .A1(DP_OP_424J2_126_3477_n2575), .A2(
        DP_OP_422J2_124_3477_n2670), .Y(DP_OP_423J2_125_3477_n2631) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1869 ( .A1(DP_OP_422J2_124_3477_n2354), 
        .A2(n86), .Y(DP_OP_423J2_125_3477_n2630) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1846 ( .A1(n1441), .A2(
        DP_OP_423J2_125_3477_n2623), .Y(DP_OP_423J2_125_3477_n2607) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1845 ( .A1(n1441), .A2(
        DP_OP_423J2_125_3477_n2622), .Y(DP_OP_423J2_125_3477_n2606) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1833 ( .A1(DP_OP_423J2_125_3477_n2618), .A2(
        DP_OP_423J2_125_3477_n2627), .Y(DP_OP_423J2_125_3477_n2594) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1832 ( .A1(DP_OP_423J2_125_3477_n2625), .A2(
        n1331), .Y(DP_OP_423J2_125_3477_n2593) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1831 ( .A1(DP_OP_423J2_125_3477_n2624), .A2(
        n1331), .Y(DP_OP_423J2_125_3477_n2592) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1829 ( .A1(DP_OP_423J2_125_3477_n2622), .A2(
        n1331), .Y(DP_OP_423J2_125_3477_n2590) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1828 ( .A1(DP_OP_423J2_125_3477_n2621), .A2(
        DP_OP_422J2_124_3477_n2626), .Y(DP_OP_423J2_125_3477_n2589) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1827 ( .A1(DP_OP_423J2_125_3477_n2620), .A2(
        DP_OP_422J2_124_3477_n2626), .Y(DP_OP_423J2_125_3477_n2588) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1826 ( .A1(DP_OP_423J2_125_3477_n2619), .A2(
        DP_OP_422J2_124_3477_n2626), .Y(DP_OP_423J2_125_3477_n2587) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1825 ( .A1(DP_OP_423J2_125_3477_n2618), 
        .A2(DP_OP_422J2_124_3477_n2626), .Y(DP_OP_423J2_125_3477_n2586) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1806 ( .A1(DP_OP_422J2_124_3477_n2443), 
        .A2(DP_OP_423J2_125_3477_n2585), .Y(DP_OP_423J2_125_3477_n2567) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1805 ( .A1(DP_OP_422J2_124_3477_n2442), .A2(
        DP_OP_422J2_124_3477_n2585), .Y(DP_OP_423J2_125_3477_n2566) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1798 ( .A1(DP_OP_422J2_124_3477_n2443), 
        .A2(n185), .Y(DP_OP_423J2_125_3477_n2559) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1797 ( .A1(DP_OP_422J2_124_3477_n2442), .A2(
        n186), .Y(DP_OP_423J2_125_3477_n2558) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1790 ( .A1(DP_OP_422J2_124_3477_n2443), 
        .A2(n671), .Y(DP_OP_423J2_125_3477_n2551) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1788 ( .A1(DP_OP_423J2_125_3477_n2581), .A2(
        DP_OP_422J2_124_3477_n2582), .Y(DP_OP_423J2_125_3477_n2549) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1787 ( .A1(DP_OP_422J2_124_3477_n2448), .A2(
        DP_OP_425J2_127_3477_n2582), .Y(DP_OP_423J2_125_3477_n2548) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1786 ( .A1(DP_OP_423J2_125_3477_n2579), .A2(
        n424), .Y(DP_OP_423J2_125_3477_n2547) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1785 ( .A1(DP_OP_422J2_124_3477_n2446), .A2(
        DP_OP_422J2_124_3477_n2582), .Y(DP_OP_423J2_125_3477_n2546) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1784 ( .A1(DP_OP_422J2_124_3477_n2445), .A2(
        n424), .Y(DP_OP_423J2_125_3477_n2545) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1783 ( .A1(DP_OP_422J2_124_3477_n2444), .A2(
        DP_OP_425J2_127_3477_n2582), .Y(DP_OP_423J2_125_3477_n2544) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1782 ( .A1(DP_OP_422J2_124_3477_n2443), .A2(
        DP_OP_422J2_124_3477_n2582), .Y(DP_OP_423J2_125_3477_n2543) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1781 ( .A1(DP_OP_422J2_124_3477_n2442), 
        .A2(n424), .Y(DP_OP_423J2_125_3477_n2542) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1763 ( .A1(DP_OP_422J2_124_3477_n2488), 
        .A2(DP_OP_425J2_127_3477_n2541), .Y(DP_OP_423J2_125_3477_n2524) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1762 ( .A1(DP_OP_423J2_125_3477_n2531), 
        .A2(DP_OP_425J2_127_3477_n2541), .Y(DP_OP_423J2_125_3477_n2523) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1761 ( .A1(DP_OP_422J2_124_3477_n2486), .A2(
        DP_OP_424J2_126_3477_n2541), .Y(DP_OP_423J2_125_3477_n2522) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1754 ( .A1(DP_OP_423J2_125_3477_n2531), 
        .A2(DP_OP_424J2_126_3477_n2540), .Y(DP_OP_423J2_125_3477_n2515) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1746 ( .A1(DP_OP_423J2_125_3477_n2531), 
        .A2(n770), .Y(DP_OP_423J2_125_3477_n2507) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1745 ( .A1(DP_OP_422J2_124_3477_n2486), .A2(
        n772), .Y(DP_OP_423J2_125_3477_n2506) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1744 ( .A1(DP_OP_423J2_125_3477_n2537), .A2(
        n1334), .Y(DP_OP_423J2_125_3477_n2505) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1743 ( .A1(DP_OP_423J2_125_3477_n2536), .A2(
        n1337), .Y(DP_OP_423J2_125_3477_n2504) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1742 ( .A1(DP_OP_422J2_124_3477_n2491), .A2(
        n1336), .Y(DP_OP_423J2_125_3477_n2503) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1740 ( .A1(DP_OP_422J2_124_3477_n2489), .A2(
        n1337), .Y(DP_OP_423J2_125_3477_n2501) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1739 ( .A1(DP_OP_422J2_124_3477_n2488), .A2(
        n1334), .Y(DP_OP_423J2_125_3477_n2500) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1738 ( .A1(DP_OP_423J2_125_3477_n2531), .A2(
        n1336), .Y(DP_OP_423J2_125_3477_n2499) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1737 ( .A1(DP_OP_422J2_124_3477_n2486), 
        .A2(n1336), .Y(DP_OP_423J2_125_3477_n2498) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1724 ( .A1(DP_OP_423J2_125_3477_n2493), 
        .A2(DP_OP_425J2_127_3477_n2497), .Y(DP_OP_423J2_125_3477_n2485) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1723 ( .A1(DP_OP_422J2_124_3477_n2580), 
        .A2(DP_OP_424J2_126_3477_n2497), .Y(DP_OP_423J2_125_3477_n2484) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1722 ( .A1(DP_OP_422J2_124_3477_n2579), 
        .A2(DP_OP_422J2_124_3477_n2497), .Y(DP_OP_423J2_125_3477_n2483) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1721 ( .A1(DP_OP_422J2_124_3477_n2578), 
        .A2(DP_OP_424J2_126_3477_n2497), .Y(DP_OP_423J2_125_3477_n2482) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1720 ( .A1(DP_OP_422J2_124_3477_n2577), 
        .A2(DP_OP_422J2_124_3477_n2497), .Y(DP_OP_423J2_125_3477_n2481) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1719 ( .A1(DP_OP_422J2_124_3477_n2576), 
        .A2(DP_OP_424J2_126_3477_n2497), .Y(DP_OP_423J2_125_3477_n2480) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1718 ( .A1(DP_OP_422J2_124_3477_n2575), 
        .A2(DP_OP_422J2_124_3477_n2497), .Y(DP_OP_423J2_125_3477_n2479) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1717 ( .A1(DP_OP_422J2_124_3477_n2574), .A2(
        DP_OP_422J2_124_3477_n2497), .Y(DP_OP_423J2_125_3477_n2478) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1710 ( .A1(DP_OP_422J2_124_3477_n2575), 
        .A2(DP_OP_423J2_125_3477_n2496), .Y(DP_OP_423J2_125_3477_n2471) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1673 ( .A1(DP_OP_422J2_124_3477_n2618), .A2(
        DP_OP_425J2_127_3477_n2453), .Y(DP_OP_423J2_125_3477_n2434) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1657 ( .A1(DP_OP_422J2_124_3477_n2618), .A2(
        n789), .Y(DP_OP_423J2_125_3477_n2418) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1634 ( .A1(DP_OP_424J2_126_3477_n2491), 
        .A2(DP_OP_423J2_125_3477_n2409), .Y(DP_OP_423J2_125_3477_n2395) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1633 ( .A1(DP_OP_425J2_127_3477_n2534), 
        .A2(DP_OP_423J2_125_3477_n2409), .Y(DP_OP_423J2_125_3477_n2394) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1631 ( .A1(DP_OP_423J2_125_3477_n2400), 
        .A2(DP_OP_423J2_125_3477_n2409), .Y(DP_OP_423J2_125_3477_n2392) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1630 ( .A1(DP_OP_423J2_125_3477_n2399), 
        .A2(DP_OP_423J2_125_3477_n2409), .Y(DP_OP_423J2_125_3477_n2391) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1629 ( .A1(DP_OP_424J2_126_3477_n2486), .A2(
        DP_OP_424J2_126_3477_n2409), .Y(DP_OP_423J2_125_3477_n2390) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1624 ( .A1(DP_OP_423J2_125_3477_n2401), 
        .A2(n1346), .Y(DP_OP_423J2_125_3477_n2385) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1623 ( .A1(DP_OP_423J2_125_3477_n2400), 
        .A2(DP_OP_424J2_126_3477_n2408), .Y(DP_OP_423J2_125_3477_n2384) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1621 ( .A1(DP_OP_424J2_126_3477_n2486), .A2(
        n1333), .Y(DP_OP_423J2_125_3477_n2382) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1614 ( .A1(DP_OP_423J2_125_3477_n2399), 
        .A2(n795), .Y(DP_OP_423J2_125_3477_n2375) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1613 ( .A1(DP_OP_424J2_126_3477_n2486), .A2(
        n799), .Y(DP_OP_423J2_125_3477_n2374) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1612 ( .A1(DP_OP_423J2_125_3477_n2405), .A2(
        n1433), .Y(DP_OP_423J2_125_3477_n2373) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1610 ( .A1(DP_OP_424J2_126_3477_n2491), .A2(
        DP_OP_422J2_124_3477_n2406), .Y(DP_OP_423J2_125_3477_n2371) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1605 ( .A1(DP_OP_424J2_126_3477_n2486), 
        .A2(n1433), .Y(DP_OP_423J2_125_3477_n2366) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1568 ( .A1(DP_OP_423J2_125_3477_n2361), .A2(
        DP_OP_423J2_125_3477_n2362), .Y(DP_OP_423J2_125_3477_n2329) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1567 ( .A1(DP_OP_422J2_124_3477_n2712), .A2(
        DP_OP_423J2_125_3477_n2362), .Y(DP_OP_423J2_125_3477_n2328) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1566 ( .A1(DP_OP_425J2_127_3477_n2579), .A2(
        DP_OP_423J2_125_3477_n2362), .Y(DP_OP_423J2_125_3477_n2327) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1565 ( .A1(DP_OP_422J2_124_3477_n2710), .A2(
        DP_OP_423J2_125_3477_n2362), .Y(DP_OP_423J2_125_3477_n2326) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1564 ( .A1(DP_OP_425J2_127_3477_n2577), .A2(
        DP_OP_423J2_125_3477_n2362), .Y(DP_OP_423J2_125_3477_n2325) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1563 ( .A1(DP_OP_425J2_127_3477_n2576), .A2(
        DP_OP_423J2_125_3477_n2362), .Y(DP_OP_423J2_125_3477_n2324) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1562 ( .A1(DP_OP_424J2_126_3477_n2443), .A2(
        DP_OP_423J2_125_3477_n2362), .Y(DP_OP_423J2_125_3477_n2323) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1561 ( .A1(DP_OP_423J2_125_3477_n2354), 
        .A2(DP_OP_423J2_125_3477_n2362), .Y(DP_OP_423J2_125_3477_n2322) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1542 ( .A1(DP_OP_423J2_125_3477_n2311), 
        .A2(DP_OP_423J2_125_3477_n2321), .Y(DP_OP_423J2_125_3477_n2303) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1536 ( .A1(DP_OP_425J2_127_3477_n2621), 
        .A2(DP_OP_425J2_127_3477_n2320), .Y(DP_OP_423J2_125_3477_n2297) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1534 ( .A1(DP_OP_423J2_125_3477_n2311), 
        .A2(DP_OP_422J2_124_3477_n2320), .Y(DP_OP_423J2_125_3477_n2295) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1533 ( .A1(DP_OP_423J2_125_3477_n2310), .A2(
        DP_OP_423J2_125_3477_n2320), .Y(DP_OP_423J2_125_3477_n2294) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1524 ( .A1(DP_OP_423J2_125_3477_n2317), .A2(
        DP_OP_423J2_125_3477_n2318), .Y(DP_OP_423J2_125_3477_n2285) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1523 ( .A1(DP_OP_423J2_125_3477_n2316), .A2(
        DP_OP_423J2_125_3477_n2318), .Y(DP_OP_423J2_125_3477_n2284) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1522 ( .A1(DP_OP_423J2_125_3477_n2315), .A2(
        DP_OP_423J2_125_3477_n2318), .Y(DP_OP_423J2_125_3477_n2283) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1521 ( .A1(DP_OP_425J2_127_3477_n2622), .A2(
        DP_OP_423J2_125_3477_n2318), .Y(DP_OP_423J2_125_3477_n2282) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1520 ( .A1(DP_OP_425J2_127_3477_n2621), .A2(
        DP_OP_423J2_125_3477_n2318), .Y(DP_OP_423J2_125_3477_n2281) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1519 ( .A1(DP_OP_425J2_127_3477_n2620), .A2(
        DP_OP_423J2_125_3477_n2318), .Y(DP_OP_423J2_125_3477_n2280) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1518 ( .A1(DP_OP_423J2_125_3477_n2311), .A2(
        DP_OP_423J2_125_3477_n2318), .Y(DP_OP_423J2_125_3477_n2279) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1517 ( .A1(DP_OP_423J2_125_3477_n2310), 
        .A2(DP_OP_423J2_125_3477_n2318), .Y(DP_OP_423J2_125_3477_n2278) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1498 ( .A1(DP_OP_423J2_125_3477_n2267), 
        .A2(DP_OP_423J2_125_3477_n2277), .Y(DP_OP_423J2_125_3477_n2259) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1497 ( .A1(DP_OP_424J2_126_3477_n2354), .A2(
        DP_OP_423J2_125_3477_n2277), .Y(DP_OP_423J2_125_3477_n2258) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1489 ( .A1(DP_OP_424J2_126_3477_n2354), .A2(
        DP_OP_423J2_125_3477_n2276), .Y(DP_OP_423J2_125_3477_n2250) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1488 ( .A1(DP_OP_423J2_125_3477_n2273), 
        .A2(DP_OP_422J2_124_3477_n2275), .Y(DP_OP_423J2_125_3477_n2249) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1487 ( .A1(DP_OP_423J2_125_3477_n2272), 
        .A2(n1427), .Y(DP_OP_423J2_125_3477_n2248) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1486 ( .A1(DP_OP_423J2_125_3477_n2271), 
        .A2(DP_OP_422J2_124_3477_n2275), .Y(DP_OP_423J2_125_3477_n2247) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1485 ( .A1(DP_OP_422J2_124_3477_n2798), 
        .A2(DP_OP_422J2_124_3477_n2275), .Y(DP_OP_423J2_125_3477_n2246) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1484 ( .A1(DP_OP_423J2_125_3477_n2269), 
        .A2(n1427), .Y(DP_OP_423J2_125_3477_n2245) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1483 ( .A1(DP_OP_423J2_125_3477_n2268), 
        .A2(DP_OP_424J2_126_3477_n2275), .Y(DP_OP_423J2_125_3477_n2244) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1482 ( .A1(DP_OP_423J2_125_3477_n2267), 
        .A2(DP_OP_424J2_126_3477_n2275), .Y(DP_OP_423J2_125_3477_n2243) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1481 ( .A1(DP_OP_424J2_126_3477_n2354), .A2(
        DP_OP_422J2_124_3477_n2275), .Y(DP_OP_423J2_125_3477_n2242) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1480 ( .A1(DP_OP_423J2_125_3477_n2273), .A2(
        n1370), .Y(DP_OP_423J2_125_3477_n2241) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1479 ( .A1(DP_OP_423J2_125_3477_n2272), .A2(
        n1338), .Y(DP_OP_423J2_125_3477_n2240) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1478 ( .A1(DP_OP_423J2_125_3477_n2271), .A2(
        n1338), .Y(DP_OP_423J2_125_3477_n2239) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1477 ( .A1(DP_OP_424J2_126_3477_n2358), .A2(
        n1338), .Y(DP_OP_423J2_125_3477_n2238) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1476 ( .A1(DP_OP_423J2_125_3477_n2269), .A2(
        DP_OP_424J2_126_3477_n2274), .Y(DP_OP_423J2_125_3477_n2237) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1475 ( .A1(DP_OP_423J2_125_3477_n2268), .A2(
        n1370), .Y(DP_OP_423J2_125_3477_n2236) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1474 ( .A1(DP_OP_423J2_125_3477_n2267), .A2(
        n1370), .Y(DP_OP_423J2_125_3477_n2235) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1473 ( .A1(DP_OP_424J2_126_3477_n2354), 
        .A2(n1370), .Y(DP_OP_423J2_125_3477_n2234) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1454 ( .A1(DP_OP_422J2_124_3477_n2839), 
        .A2(DP_OP_423J2_125_3477_n2233), .Y(DP_OP_423J2_125_3477_n2215) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1453 ( .A1(DP_OP_423J2_125_3477_n2222), .A2(
        DP_OP_423J2_125_3477_n2233), .Y(DP_OP_423J2_125_3477_n2214) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1445 ( .A1(DP_OP_423J2_125_3477_n2222), .A2(
        n365), .Y(DP_OP_423J2_125_3477_n2206) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1439 ( .A1(DP_OP_425J2_127_3477_n2708), 
        .A2(DP_OP_424J2_126_3477_n2231), .Y(DP_OP_423J2_125_3477_n2200) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1437 ( .A1(DP_OP_423J2_125_3477_n2222), .A2(
        DP_OP_424J2_126_3477_n2231), .Y(DP_OP_423J2_125_3477_n2198) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1436 ( .A1(DP_OP_423J2_125_3477_n2229), .A2(
        DP_OP_422J2_124_3477_n2230), .Y(DP_OP_423J2_125_3477_n2197) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1432 ( .A1(DP_OP_423J2_125_3477_n2225), .A2(
        DP_OP_423J2_125_3477_n2230), .Y(DP_OP_423J2_125_3477_n2193) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1416 ( .A1(DP_OP_423J2_125_3477_n2185), 
        .A2(DP_OP_424J2_126_3477_n2189), .Y(DP_OP_423J2_125_3477_n2177) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1415 ( .A1(DP_OP_425J2_127_3477_n2756), 
        .A2(DP_OP_424J2_126_3477_n2189), .Y(DP_OP_423J2_125_3477_n2176) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1414 ( .A1(DP_OP_425J2_127_3477_n2755), 
        .A2(DP_OP_425J2_127_3477_n2189), .Y(DP_OP_423J2_125_3477_n2175) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1413 ( .A1(DP_OP_423J2_125_3477_n2182), 
        .A2(DP_OP_425J2_127_3477_n2189), .Y(DP_OP_423J2_125_3477_n2174) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1412 ( .A1(DP_OP_424J2_126_3477_n2269), 
        .A2(DP_OP_424J2_126_3477_n2189), .Y(DP_OP_423J2_125_3477_n2173) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1411 ( .A1(DP_OP_424J2_126_3477_n2268), 
        .A2(DP_OP_424J2_126_3477_n2189), .Y(DP_OP_423J2_125_3477_n2172) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1410 ( .A1(DP_OP_424J2_126_3477_n2267), 
        .A2(DP_OP_425J2_127_3477_n2189), .Y(DP_OP_423J2_125_3477_n2171) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1409 ( .A1(DP_OP_423J2_125_3477_n2178), .A2(
        DP_OP_425J2_127_3477_n2189), .Y(DP_OP_423J2_125_3477_n2170) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1401 ( .A1(DP_OP_423J2_125_3477_n2178), .A2(
        n1344), .Y(DP_OP_423J2_125_3477_n2162) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1394 ( .A1(DP_OP_422J2_124_3477_n2883), 
        .A2(n1339), .Y(DP_OP_423J2_125_3477_n2155) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1393 ( .A1(DP_OP_423J2_125_3477_n2178), .A2(
        n1339), .Y(DP_OP_423J2_125_3477_n2154) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1392 ( .A1(DP_OP_423J2_125_3477_n2185), .A2(
        DP_OP_424J2_126_3477_n2186), .Y(DP_OP_423J2_125_3477_n2153) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1391 ( .A1(DP_OP_425J2_127_3477_n2756), .A2(
        DP_OP_422J2_124_3477_n2186), .Y(DP_OP_423J2_125_3477_n2152) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1390 ( .A1(DP_OP_422J2_124_3477_n2887), .A2(
        DP_OP_425J2_127_3477_n2186), .Y(DP_OP_423J2_125_3477_n2151) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1389 ( .A1(DP_OP_423J2_125_3477_n2182), .A2(
        DP_OP_424J2_126_3477_n2186), .Y(DP_OP_423J2_125_3477_n2150) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1388 ( .A1(DP_OP_424J2_126_3477_n2269), .A2(
        DP_OP_425J2_127_3477_n2186), .Y(DP_OP_423J2_125_3477_n2149) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1386 ( .A1(DP_OP_424J2_126_3477_n2267), .A2(
        DP_OP_422J2_124_3477_n2186), .Y(DP_OP_423J2_125_3477_n2147) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1385 ( .A1(DP_OP_423J2_125_3477_n2178), 
        .A2(DP_OP_425J2_127_3477_n2186), .Y(DP_OP_423J2_125_3477_n2146) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1366 ( .A1(DP_OP_423J2_125_3477_n2135), 
        .A2(n1442), .Y(DP_OP_423J2_125_3477_n2127) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1358 ( .A1(DP_OP_423J2_125_3477_n2135), 
        .A2(DP_OP_424J2_126_3477_n2144), .Y(DP_OP_423J2_125_3477_n2119) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1357 ( .A1(DP_OP_422J2_124_3477_n2926), .A2(
        DP_OP_425J2_127_3477_n2144), .Y(DP_OP_423J2_125_3477_n2118) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1350 ( .A1(DP_OP_423J2_125_3477_n2135), 
        .A2(DP_OP_425J2_127_3477_n2143), .Y(DP_OP_423J2_125_3477_n2111) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1349 ( .A1(DP_OP_424J2_126_3477_n2222), .A2(
        DP_OP_424J2_126_3477_n2143), .Y(DP_OP_423J2_125_3477_n2110) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1322 ( .A1(DP_OP_425J2_127_3477_n2839), 
        .A2(n621), .Y(DP_OP_423J2_125_3477_n2083) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1315 ( .A1(DP_OP_425J2_127_3477_n2840), 
        .A2(DP_OP_422J2_124_3477_n2100), .Y(DP_OP_423J2_125_3477_n2076) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1314 ( .A1(DP_OP_425J2_127_3477_n2839), 
        .A2(DP_OP_423J2_125_3477_n2100), .Y(DP_OP_423J2_125_3477_n2075) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1313 ( .A1(DP_OP_423J2_125_3477_n2090), .A2(
        DP_OP_424J2_126_3477_n2100), .Y(DP_OP_423J2_125_3477_n2074) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1306 ( .A1(DP_OP_425J2_127_3477_n2839), 
        .A2(DP_OP_423J2_125_3477_n2099), .Y(DP_OP_423J2_125_3477_n2067) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1303 ( .A1(DP_OP_423J2_125_3477_n2096), .A2(
        DP_OP_425J2_127_3477_n2098), .Y(DP_OP_423J2_125_3477_n2064) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1300 ( .A1(DP_OP_425J2_127_3477_n2841), .A2(
        n1439), .Y(DP_OP_423J2_125_3477_n2061) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1279 ( .A1(DP_OP_423J2_125_3477_n2048), 
        .A2(DP_OP_425J2_127_3477_n2057), .Y(DP_OP_423J2_125_3477_n2040) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1278 ( .A1(DP_OP_425J2_127_3477_n2883), 
        .A2(DP_OP_425J2_127_3477_n2057), .Y(DP_OP_423J2_125_3477_n2039) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1277 ( .A1(DP_OP_425J2_127_3477_n2882), .A2(
        n1475), .Y(DP_OP_423J2_125_3477_n2038) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1270 ( .A1(DP_OP_422J2_124_3477_n3015), 
        .A2(DP_OP_425J2_127_3477_n2056), .Y(DP_OP_423J2_125_3477_n2031) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1269 ( .A1(DP_OP_422J2_124_3477_n3014), .A2(
        DP_OP_424J2_126_3477_n2056), .Y(DP_OP_423J2_125_3477_n2030) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1262 ( .A1(DP_OP_425J2_127_3477_n2883), 
        .A2(DP_OP_425J2_127_3477_n2055), .Y(DP_OP_423J2_125_3477_n2023) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1261 ( .A1(DP_OP_422J2_124_3477_n3014), .A2(
        DP_OP_424J2_126_3477_n2055), .Y(DP_OP_423J2_125_3477_n2022) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1259 ( .A1(DP_OP_423J2_125_3477_n2052), .A2(
        n30), .Y(DP_OP_423J2_125_3477_n2020) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1258 ( .A1(DP_OP_423J2_125_3477_n2051), .A2(
        n30), .Y(DP_OP_423J2_125_3477_n2019) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1257 ( .A1(DP_OP_425J2_127_3477_n2886), .A2(
        n779), .Y(DP_OP_423J2_125_3477_n2018) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1256 ( .A1(DP_OP_425J2_127_3477_n2885), .A2(
        n30), .Y(DP_OP_423J2_125_3477_n2017) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1255 ( .A1(DP_OP_423J2_125_3477_n2048), .A2(
        n776), .Y(DP_OP_423J2_125_3477_n2016) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1254 ( .A1(DP_OP_422J2_124_3477_n3015), .A2(
        n30), .Y(DP_OP_423J2_125_3477_n2015) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1253 ( .A1(DP_OP_422J2_124_3477_n3014), 
        .A2(n30), .Y(DP_OP_423J2_125_3477_n2014) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1240 ( .A1(DP_OP_425J2_127_3477_n2933), 
        .A2(n1431), .Y(DP_OP_423J2_125_3477_n2001) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1238 ( .A1(DP_OP_423J2_125_3477_n2007), 
        .A2(DP_OP_423J2_125_3477_n2013), .Y(DP_OP_423J2_125_3477_n1999) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1237 ( .A1(DP_OP_423J2_125_3477_n2006), 
        .A2(DP_OP_423J2_125_3477_n2013), .Y(DP_OP_423J2_125_3477_n1998) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1235 ( .A1(DP_OP_422J2_124_3477_n3058), 
        .A2(DP_OP_423J2_125_3477_n2013), .Y(DP_OP_423J2_125_3477_n1996) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1234 ( .A1(DP_OP_423J2_125_3477_n2003), 
        .A2(DP_OP_423J2_125_3477_n2013), .Y(DP_OP_423J2_125_3477_n1995) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1233 ( .A1(DP_OP_424J2_126_3477_n2090), .A2(
        DP_OP_423J2_125_3477_n2013), .Y(DP_OP_423J2_125_3477_n1994) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1226 ( .A1(DP_OP_423J2_125_3477_n2003), 
        .A2(n558), .Y(DP_OP_423J2_125_3477_n1987) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1225 ( .A1(DP_OP_424J2_126_3477_n2090), .A2(
        n558), .Y(DP_OP_423J2_125_3477_n1986) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1217 ( .A1(DP_OP_424J2_126_3477_n2090), .A2(
        DP_OP_422J2_124_3477_n2011), .Y(DP_OP_423J2_125_3477_n1978) );
  OR2X1_HVT DP_OP_423J2_125_3477_U1214 ( .A1(DP_OP_423J2_125_3477_n2007), .A2(
        DP_OP_423J2_125_3477_n2010), .Y(DP_OP_423J2_125_3477_n1975) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1165 ( .A1(n1850), .A2(n1508), .Y(
        DP_OP_423J2_125_3477_n510) );
  HADDX1_HVT DP_OP_423J2_125_3477_U1143 ( .A0(DP_OP_423J2_125_3477_n1936), 
        .B0(DP_OP_423J2_125_3477_n2045), .C1(DP_OP_423J2_125_3477_n1920), .SO(
        DP_OP_423J2_125_3477_n1921) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1142 ( .A(DP_OP_423J2_125_3477_n2089), .B(
        DP_OP_423J2_125_3477_n2001), .CI(DP_OP_423J2_125_3477_n2133), .CO(
        DP_OP_423J2_125_3477_n1918), .S(DP_OP_423J2_125_3477_n1919) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1141 ( .A(DP_OP_423J2_125_3477_n2221), .B(
        DP_OP_423J2_125_3477_n2177), .CI(DP_OP_423J2_125_3477_n2265), .CO(
        DP_OP_423J2_125_3477_n1916), .S(DP_OP_423J2_125_3477_n1917) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1140 ( .A(DP_OP_423J2_125_3477_n2353), .B(
        DP_OP_423J2_125_3477_n2309), .CI(DP_OP_423J2_125_3477_n2397), .CO(
        DP_OP_423J2_125_3477_n1914), .S(DP_OP_423J2_125_3477_n1915) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1139 ( .A(DP_OP_423J2_125_3477_n2485), .B(
        DP_OP_423J2_125_3477_n2441), .CI(DP_OP_423J2_125_3477_n2529), .CO(
        DP_OP_423J2_125_3477_n1912), .S(DP_OP_423J2_125_3477_n1913) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1138 ( .A(DP_OP_423J2_125_3477_n2617), .B(
        DP_OP_423J2_125_3477_n2573), .CI(DP_OP_423J2_125_3477_n2661), .CO(
        DP_OP_423J2_125_3477_n1910), .S(DP_OP_423J2_125_3477_n1911) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1137 ( .A(DP_OP_423J2_125_3477_n2749), .B(
        DP_OP_423J2_125_3477_n2705), .CI(DP_OP_423J2_125_3477_n2793), .CO(
        DP_OP_423J2_125_3477_n1908), .S(DP_OP_423J2_125_3477_n1909) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1136 ( .A(DP_OP_423J2_125_3477_n3055), .B(
        DP_OP_423J2_125_3477_n2837), .CI(DP_OP_423J2_125_3477_n2881), .CO(
        DP_OP_423J2_125_3477_n1906), .S(DP_OP_423J2_125_3477_n1907) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1135 ( .A(DP_OP_423J2_125_3477_n3013), .B(
        DP_OP_423J2_125_3477_n2925), .CI(DP_OP_423J2_125_3477_n2969), .CO(
        DP_OP_423J2_125_3477_n1904), .S(DP_OP_423J2_125_3477_n1905) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1134 ( .A(DP_OP_423J2_125_3477_n1921), .B(
        DP_OP_423J2_125_3477_n1907), .CI(DP_OP_423J2_125_3477_n1909), .CO(
        DP_OP_423J2_125_3477_n1902), .S(DP_OP_423J2_125_3477_n1903) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1133 ( .A(DP_OP_423J2_125_3477_n1911), .B(
        DP_OP_423J2_125_3477_n1905), .CI(DP_OP_423J2_125_3477_n1913), .CO(
        DP_OP_423J2_125_3477_n1900), .S(DP_OP_423J2_125_3477_n1901) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1132 ( .A(DP_OP_423J2_125_3477_n1919), .B(
        DP_OP_423J2_125_3477_n1915), .CI(DP_OP_423J2_125_3477_n1917), .CO(
        DP_OP_423J2_125_3477_n1898), .S(DP_OP_423J2_125_3477_n1899) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1130 ( .A(DP_OP_423J2_125_3477_n2037), .B(
        DP_OP_423J2_125_3477_n1993), .CI(DP_OP_423J2_125_3477_n2044), .CO(
        DP_OP_423J2_125_3477_n1894), .S(DP_OP_423J2_125_3477_n1895) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1129 ( .A(DP_OP_423J2_125_3477_n2088), .B(
        DP_OP_423J2_125_3477_n2081), .CI(DP_OP_423J2_125_3477_n2125), .CO(
        DP_OP_423J2_125_3477_n1892), .S(DP_OP_423J2_125_3477_n1893) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1128 ( .A(DP_OP_423J2_125_3477_n2169), .B(
        DP_OP_423J2_125_3477_n2132), .CI(DP_OP_423J2_125_3477_n2176), .CO(
        DP_OP_423J2_125_3477_n1890), .S(DP_OP_423J2_125_3477_n1891) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1127 ( .A(DP_OP_423J2_125_3477_n2220), .B(
        DP_OP_423J2_125_3477_n2213), .CI(DP_OP_423J2_125_3477_n2257), .CO(
        DP_OP_423J2_125_3477_n1888), .S(DP_OP_423J2_125_3477_n1889) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1126 ( .A(DP_OP_423J2_125_3477_n2301), .B(
        DP_OP_423J2_125_3477_n2264), .CI(DP_OP_423J2_125_3477_n2308), .CO(
        DP_OP_423J2_125_3477_n1886), .S(DP_OP_423J2_125_3477_n1887) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1125 ( .A(DP_OP_423J2_125_3477_n2352), .B(
        DP_OP_423J2_125_3477_n2345), .CI(DP_OP_423J2_125_3477_n2389), .CO(
        DP_OP_423J2_125_3477_n1884), .S(DP_OP_423J2_125_3477_n1885) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1124 ( .A(DP_OP_423J2_125_3477_n2433), .B(
        DP_OP_423J2_125_3477_n2396), .CI(DP_OP_423J2_125_3477_n2440), .CO(
        DP_OP_423J2_125_3477_n1882), .S(DP_OP_423J2_125_3477_n1883) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1123 ( .A(DP_OP_423J2_125_3477_n2484), .B(
        DP_OP_423J2_125_3477_n2477), .CI(DP_OP_423J2_125_3477_n2521), .CO(
        DP_OP_423J2_125_3477_n1880), .S(DP_OP_423J2_125_3477_n1881) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1122 ( .A(DP_OP_423J2_125_3477_n2565), .B(
        DP_OP_423J2_125_3477_n2528), .CI(DP_OP_423J2_125_3477_n2572), .CO(
        DP_OP_423J2_125_3477_n1878), .S(DP_OP_423J2_125_3477_n1879) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1121 ( .A(DP_OP_423J2_125_3477_n3054), .B(
        DP_OP_423J2_125_3477_n2609), .CI(DP_OP_423J2_125_3477_n3047), .CO(
        DP_OP_423J2_125_3477_n1876), .S(DP_OP_423J2_125_3477_n1877) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1120 ( .A(DP_OP_423J2_125_3477_n2792), .B(
        DP_OP_423J2_125_3477_n2616), .CI(DP_OP_423J2_125_3477_n2653), .CO(
        DP_OP_423J2_125_3477_n1874), .S(DP_OP_423J2_125_3477_n1875) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1119 ( .A(DP_OP_423J2_125_3477_n2829), .B(
        DP_OP_423J2_125_3477_n3012), .CI(DP_OP_423J2_125_3477_n3005), .CO(
        DP_OP_423J2_125_3477_n1872), .S(DP_OP_423J2_125_3477_n1873) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1118 ( .A(DP_OP_423J2_125_3477_n2748), .B(
        DP_OP_423J2_125_3477_n2968), .CI(DP_OP_423J2_125_3477_n2961), .CO(
        DP_OP_423J2_125_3477_n1870), .S(DP_OP_423J2_125_3477_n1871) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1117 ( .A(DP_OP_423J2_125_3477_n2741), .B(
        DP_OP_423J2_125_3477_n2924), .CI(DP_OP_423J2_125_3477_n2660), .CO(
        DP_OP_423J2_125_3477_n1868), .S(DP_OP_423J2_125_3477_n1869) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1116 ( .A(DP_OP_423J2_125_3477_n2917), .B(
        DP_OP_423J2_125_3477_n2697), .CI(DP_OP_423J2_125_3477_n2704), .CO(
        DP_OP_423J2_125_3477_n1866), .S(DP_OP_423J2_125_3477_n1867) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1115 ( .A(DP_OP_423J2_125_3477_n2873), .B(
        DP_OP_423J2_125_3477_n2785), .CI(DP_OP_423J2_125_3477_n2836), .CO(
        DP_OP_423J2_125_3477_n1864), .S(DP_OP_423J2_125_3477_n1865) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1114 ( .A(DP_OP_423J2_125_3477_n2880), .B(
        DP_OP_423J2_125_3477_n1920), .CI(DP_OP_423J2_125_3477_n1897), .CO(
        DP_OP_423J2_125_3477_n1862), .S(DP_OP_423J2_125_3477_n1863) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1113 ( .A(DP_OP_423J2_125_3477_n1904), .B(
        DP_OP_423J2_125_3477_n1918), .CI(DP_OP_423J2_125_3477_n1916), .CO(
        DP_OP_423J2_125_3477_n1860), .S(DP_OP_423J2_125_3477_n1861) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1112 ( .A(DP_OP_423J2_125_3477_n1910), .B(
        DP_OP_423J2_125_3477_n1906), .CI(DP_OP_423J2_125_3477_n1914), .CO(
        DP_OP_423J2_125_3477_n1858), .S(DP_OP_423J2_125_3477_n1859) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1111 ( .A(DP_OP_423J2_125_3477_n1912), .B(
        DP_OP_423J2_125_3477_n1908), .CI(DP_OP_423J2_125_3477_n1865), .CO(
        DP_OP_423J2_125_3477_n1856), .S(DP_OP_423J2_125_3477_n1857) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1110 ( .A(DP_OP_423J2_125_3477_n1887), .B(
        DP_OP_423J2_125_3477_n1873), .CI(DP_OP_423J2_125_3477_n1871), .CO(
        DP_OP_423J2_125_3477_n1854), .S(DP_OP_423J2_125_3477_n1855) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1109 ( .A(DP_OP_423J2_125_3477_n1891), .B(
        DP_OP_423J2_125_3477_n1875), .CI(DP_OP_423J2_125_3477_n1879), .CO(
        DP_OP_423J2_125_3477_n1852), .S(DP_OP_423J2_125_3477_n1853) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1108 ( .A(DP_OP_423J2_125_3477_n1893), .B(
        DP_OP_423J2_125_3477_n1881), .CI(DP_OP_423J2_125_3477_n1877), .CO(
        DP_OP_423J2_125_3477_n1850), .S(DP_OP_423J2_125_3477_n1851) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1107 ( .A(DP_OP_423J2_125_3477_n1895), .B(
        DP_OP_423J2_125_3477_n1885), .CI(DP_OP_423J2_125_3477_n1869), .CO(
        DP_OP_423J2_125_3477_n1848), .S(DP_OP_423J2_125_3477_n1849) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1106 ( .A(DP_OP_423J2_125_3477_n1889), .B(
        DP_OP_423J2_125_3477_n1883), .CI(DP_OP_423J2_125_3477_n1867), .CO(
        DP_OP_423J2_125_3477_n1846), .S(DP_OP_423J2_125_3477_n1847) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1105 ( .A(DP_OP_423J2_125_3477_n1863), .B(
        DP_OP_423J2_125_3477_n1902), .CI(DP_OP_423J2_125_3477_n1900), .CO(
        DP_OP_423J2_125_3477_n1844), .S(DP_OP_423J2_125_3477_n1845) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1104 ( .A(DP_OP_423J2_125_3477_n1898), .B(
        DP_OP_423J2_125_3477_n1859), .CI(DP_OP_423J2_125_3477_n1861), .CO(
        DP_OP_423J2_125_3477_n1842), .S(DP_OP_423J2_125_3477_n1843) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1103 ( .A(DP_OP_423J2_125_3477_n1857), .B(
        DP_OP_423J2_125_3477_n1849), .CI(DP_OP_423J2_125_3477_n1851), .CO(
        DP_OP_423J2_125_3477_n1840), .S(DP_OP_423J2_125_3477_n1841) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1102 ( .A(DP_OP_423J2_125_3477_n1855), .B(
        DP_OP_423J2_125_3477_n1847), .CI(DP_OP_423J2_125_3477_n1853), .CO(
        DP_OP_423J2_125_3477_n1838), .S(DP_OP_423J2_125_3477_n1839) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1101 ( .A(DP_OP_423J2_125_3477_n1845), .B(
        DP_OP_423J2_125_3477_n1843), .CI(DP_OP_423J2_125_3477_n1841), .CO(
        DP_OP_423J2_125_3477_n1836), .S(DP_OP_423J2_125_3477_n1837) );
  HADDX1_HVT DP_OP_423J2_125_3477_U1100 ( .A0(DP_OP_423J2_125_3477_n1934), 
        .B0(DP_OP_423J2_125_3477_n1999), .C1(DP_OP_423J2_125_3477_n1834), .SO(
        DP_OP_423J2_125_3477_n1835) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1099 ( .A(DP_OP_423J2_125_3477_n2029), .B(
        DP_OP_423J2_125_3477_n1992), .CI(DP_OP_423J2_125_3477_n1985), .CO(
        DP_OP_423J2_125_3477_n1832), .S(DP_OP_423J2_125_3477_n1833) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1098 ( .A(DP_OP_423J2_125_3477_n2043), .B(
        DP_OP_423J2_125_3477_n2036), .CI(DP_OP_423J2_125_3477_n2073), .CO(
        DP_OP_423J2_125_3477_n1830), .S(DP_OP_423J2_125_3477_n1831) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1096 ( .A(DP_OP_423J2_125_3477_n2131), .B(
        DP_OP_423J2_125_3477_n2124), .CI(DP_OP_423J2_125_3477_n2161), .CO(
        DP_OP_423J2_125_3477_n1826), .S(DP_OP_423J2_125_3477_n1827) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1095 ( .A(DP_OP_423J2_125_3477_n2175), .B(
        DP_OP_423J2_125_3477_n2168), .CI(DP_OP_423J2_125_3477_n2205), .CO(
        DP_OP_423J2_125_3477_n1824), .S(DP_OP_423J2_125_3477_n1825) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1094 ( .A(DP_OP_423J2_125_3477_n2219), .B(
        DP_OP_423J2_125_3477_n2212), .CI(DP_OP_423J2_125_3477_n2249), .CO(
        DP_OP_423J2_125_3477_n1822), .S(DP_OP_423J2_125_3477_n1823) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1093 ( .A(DP_OP_423J2_125_3477_n2263), .B(
        DP_OP_423J2_125_3477_n2256), .CI(DP_OP_423J2_125_3477_n2293), .CO(
        DP_OP_423J2_125_3477_n1820), .S(DP_OP_423J2_125_3477_n1821) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1092 ( .A(DP_OP_423J2_125_3477_n2307), .B(
        DP_OP_423J2_125_3477_n2300), .CI(DP_OP_423J2_125_3477_n2337), .CO(
        DP_OP_423J2_125_3477_n1818), .S(DP_OP_423J2_125_3477_n1819) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1091 ( .A(DP_OP_423J2_125_3477_n2351), .B(
        DP_OP_423J2_125_3477_n2344), .CI(DP_OP_423J2_125_3477_n2381), .CO(
        DP_OP_423J2_125_3477_n1816), .S(DP_OP_423J2_125_3477_n1817) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1090 ( .A(DP_OP_423J2_125_3477_n2395), .B(
        DP_OP_423J2_125_3477_n2388), .CI(DP_OP_423J2_125_3477_n2425), .CO(
        DP_OP_423J2_125_3477_n1814), .S(DP_OP_423J2_125_3477_n1815) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1089 ( .A(DP_OP_423J2_125_3477_n2439), .B(
        DP_OP_423J2_125_3477_n2432), .CI(DP_OP_423J2_125_3477_n2469), .CO(
        DP_OP_423J2_125_3477_n1812), .S(DP_OP_423J2_125_3477_n1813) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1088 ( .A(DP_OP_423J2_125_3477_n2740), .B(
        DP_OP_423J2_125_3477_n3053), .CI(DP_OP_423J2_125_3477_n3046), .CO(
        DP_OP_423J2_125_3477_n1810), .S(DP_OP_423J2_125_3477_n1811) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1087 ( .A(DP_OP_423J2_125_3477_n2703), .B(
        DP_OP_423J2_125_3477_n2476), .CI(DP_OP_423J2_125_3477_n3039), .CO(
        DP_OP_423J2_125_3477_n1808), .S(DP_OP_423J2_125_3477_n1809) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1086 ( .A(DP_OP_423J2_125_3477_n2696), .B(
        DP_OP_423J2_125_3477_n3011), .CI(DP_OP_423J2_125_3477_n2483), .CO(
        DP_OP_423J2_125_3477_n1806), .S(DP_OP_423J2_125_3477_n1807) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1083 ( .A(DP_OP_423J2_125_3477_n2777), .B(
        DP_OP_423J2_125_3477_n2557), .CI(DP_OP_423J2_125_3477_n2997), .CO(
        DP_OP_423J2_125_3477_n1800), .S(DP_OP_423J2_125_3477_n1801) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1082 ( .A(DP_OP_423J2_125_3477_n2689), .B(
        DP_OP_423J2_125_3477_n2564), .CI(DP_OP_423J2_125_3477_n2967), .CO(
        DP_OP_423J2_125_3477_n1798), .S(DP_OP_423J2_125_3477_n1799) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1081 ( .A(DP_OP_423J2_125_3477_n2659), .B(
        DP_OP_423J2_125_3477_n2571), .CI(DP_OP_423J2_125_3477_n2960), .CO(
        DP_OP_423J2_125_3477_n1796), .S(DP_OP_423J2_125_3477_n1797) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1080 ( .A(DP_OP_423J2_125_3477_n2953), .B(
        DP_OP_423J2_125_3477_n2601), .CI(DP_OP_423J2_125_3477_n2608), .CO(
        DP_OP_423J2_125_3477_n1794), .S(DP_OP_423J2_125_3477_n1795) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1079 ( .A(DP_OP_423J2_125_3477_n2923), .B(
        DP_OP_423J2_125_3477_n2615), .CI(DP_OP_423J2_125_3477_n2645), .CO(
        DP_OP_423J2_125_3477_n1792), .S(DP_OP_423J2_125_3477_n1793) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1078 ( .A(DP_OP_423J2_125_3477_n2916), .B(
        DP_OP_423J2_125_3477_n2652), .CI(DP_OP_423J2_125_3477_n2784), .CO(
        DP_OP_423J2_125_3477_n1790), .S(DP_OP_423J2_125_3477_n1791) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1077 ( .A(DP_OP_423J2_125_3477_n2909), .B(
        DP_OP_423J2_125_3477_n2791), .CI(DP_OP_423J2_125_3477_n2821), .CO(
        DP_OP_423J2_125_3477_n1788), .S(DP_OP_423J2_125_3477_n1789) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1076 ( .A(DP_OP_423J2_125_3477_n2879), .B(
        DP_OP_423J2_125_3477_n2828), .CI(DP_OP_423J2_125_3477_n2835), .CO(
        DP_OP_423J2_125_3477_n1786), .S(DP_OP_423J2_125_3477_n1787) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1074 ( .A(DP_OP_423J2_125_3477_n1835), .B(
        DP_OP_423J2_125_3477_n1864), .CI(DP_OP_423J2_125_3477_n1866), .CO(
        DP_OP_423J2_125_3477_n1782), .S(DP_OP_423J2_125_3477_n1783) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1073 ( .A(DP_OP_423J2_125_3477_n1882), .B(
        DP_OP_423J2_125_3477_n1894), .CI(DP_OP_423J2_125_3477_n1868), .CO(
        DP_OP_423J2_125_3477_n1780), .S(DP_OP_423J2_125_3477_n1781) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1072 ( .A(DP_OP_423J2_125_3477_n1880), .B(
        DP_OP_423J2_125_3477_n1892), .CI(DP_OP_423J2_125_3477_n1870), .CO(
        DP_OP_423J2_125_3477_n1778), .S(DP_OP_423J2_125_3477_n1779) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1071 ( .A(DP_OP_423J2_125_3477_n1876), .B(
        DP_OP_423J2_125_3477_n1890), .CI(DP_OP_423J2_125_3477_n1872), .CO(
        DP_OP_423J2_125_3477_n1776), .S(DP_OP_423J2_125_3477_n1777) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1070 ( .A(DP_OP_423J2_125_3477_n1886), .B(
        DP_OP_423J2_125_3477_n1888), .CI(DP_OP_423J2_125_3477_n1884), .CO(
        DP_OP_423J2_125_3477_n1774), .S(DP_OP_423J2_125_3477_n1775) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1069 ( .A(DP_OP_423J2_125_3477_n1878), .B(
        DP_OP_423J2_125_3477_n1874), .CI(DP_OP_423J2_125_3477_n1807), .CO(
        DP_OP_423J2_125_3477_n1772), .S(DP_OP_423J2_125_3477_n1773) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1068 ( .A(DP_OP_423J2_125_3477_n1801), .B(
        DP_OP_423J2_125_3477_n1819), .CI(DP_OP_423J2_125_3477_n1815), .CO(
        DP_OP_423J2_125_3477_n1770), .S(DP_OP_423J2_125_3477_n1771) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1067 ( .A(DP_OP_423J2_125_3477_n1797), .B(
        DP_OP_423J2_125_3477_n1825), .CI(DP_OP_423J2_125_3477_n1827), .CO(
        DP_OP_423J2_125_3477_n1768), .S(DP_OP_423J2_125_3477_n1769) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1066 ( .A(DP_OP_423J2_125_3477_n1831), .B(
        DP_OP_423J2_125_3477_n1817), .CI(DP_OP_423J2_125_3477_n1795), .CO(
        DP_OP_423J2_125_3477_n1766), .S(DP_OP_423J2_125_3477_n1767) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1065 ( .A(DP_OP_423J2_125_3477_n1793), .B(
        DP_OP_423J2_125_3477_n1811), .CI(DP_OP_423J2_125_3477_n1829), .CO(
        DP_OP_423J2_125_3477_n1764), .S(DP_OP_423J2_125_3477_n1765) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1064 ( .A(DP_OP_423J2_125_3477_n1791), .B(
        DP_OP_423J2_125_3477_n1821), .CI(DP_OP_423J2_125_3477_n1809), .CO(
        DP_OP_423J2_125_3477_n1762), .S(DP_OP_423J2_125_3477_n1763) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1063 ( .A(DP_OP_423J2_125_3477_n1789), .B(
        DP_OP_423J2_125_3477_n1823), .CI(DP_OP_423J2_125_3477_n1833), .CO(
        DP_OP_423J2_125_3477_n1760), .S(DP_OP_423J2_125_3477_n1761) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1062 ( .A(DP_OP_423J2_125_3477_n1787), .B(
        DP_OP_423J2_125_3477_n1813), .CI(DP_OP_423J2_125_3477_n1799), .CO(
        DP_OP_423J2_125_3477_n1758), .S(DP_OP_423J2_125_3477_n1759) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1061 ( .A(DP_OP_423J2_125_3477_n1803), .B(
        DP_OP_423J2_125_3477_n1805), .CI(DP_OP_423J2_125_3477_n1862), .CO(
        DP_OP_423J2_125_3477_n1756), .S(DP_OP_423J2_125_3477_n1757) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1060 ( .A(DP_OP_423J2_125_3477_n1785), .B(
        DP_OP_423J2_125_3477_n1860), .CI(DP_OP_423J2_125_3477_n1858), .CO(
        DP_OP_423J2_125_3477_n1754), .S(DP_OP_423J2_125_3477_n1755) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1059 ( .A(DP_OP_423J2_125_3477_n1856), .B(
        DP_OP_423J2_125_3477_n1783), .CI(DP_OP_423J2_125_3477_n1850), .CO(
        DP_OP_423J2_125_3477_n1752), .S(DP_OP_423J2_125_3477_n1753) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1058 ( .A(DP_OP_423J2_125_3477_n1854), .B(
        DP_OP_423J2_125_3477_n1775), .CI(DP_OP_423J2_125_3477_n1781), .CO(
        DP_OP_423J2_125_3477_n1750), .S(DP_OP_423J2_125_3477_n1751) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1057 ( .A(DP_OP_423J2_125_3477_n1852), .B(
        DP_OP_423J2_125_3477_n1779), .CI(DP_OP_423J2_125_3477_n1777), .CO(
        DP_OP_423J2_125_3477_n1748), .S(DP_OP_423J2_125_3477_n1749) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1056 ( .A(DP_OP_423J2_125_3477_n1848), .B(
        DP_OP_423J2_125_3477_n1846), .CI(DP_OP_423J2_125_3477_n1773), .CO(
        DP_OP_423J2_125_3477_n1746), .S(DP_OP_423J2_125_3477_n1747) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1055 ( .A(DP_OP_423J2_125_3477_n1771), .B(
        DP_OP_423J2_125_3477_n1759), .CI(DP_OP_423J2_125_3477_n1757), .CO(
        DP_OP_423J2_125_3477_n1744), .S(DP_OP_423J2_125_3477_n1745) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1054 ( .A(DP_OP_423J2_125_3477_n1767), .B(
        DP_OP_423J2_125_3477_n1769), .CI(DP_OP_423J2_125_3477_n1761), .CO(
        DP_OP_423J2_125_3477_n1742), .S(DP_OP_423J2_125_3477_n1743) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1053 ( .A(DP_OP_423J2_125_3477_n1763), .B(
        DP_OP_423J2_125_3477_n1765), .CI(DP_OP_423J2_125_3477_n1844), .CO(
        DP_OP_423J2_125_3477_n1740), .S(DP_OP_423J2_125_3477_n1741) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1052 ( .A(DP_OP_423J2_125_3477_n1755), .B(
        DP_OP_423J2_125_3477_n1842), .CI(DP_OP_423J2_125_3477_n1753), .CO(
        DP_OP_423J2_125_3477_n1738), .S(DP_OP_423J2_125_3477_n1739) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1051 ( .A(DP_OP_423J2_125_3477_n1840), .B(
        DP_OP_423J2_125_3477_n1838), .CI(DP_OP_423J2_125_3477_n1749), .CO(
        DP_OP_423J2_125_3477_n1736), .S(DP_OP_423J2_125_3477_n1737) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1050 ( .A(DP_OP_423J2_125_3477_n1751), .B(
        DP_OP_423J2_125_3477_n1747), .CI(DP_OP_423J2_125_3477_n1745), .CO(
        DP_OP_423J2_125_3477_n1734), .S(DP_OP_423J2_125_3477_n1735) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1049 ( .A(DP_OP_423J2_125_3477_n1743), .B(
        DP_OP_423J2_125_3477_n1741), .CI(DP_OP_423J2_125_3477_n1739), .CO(
        DP_OP_423J2_125_3477_n1732), .S(DP_OP_423J2_125_3477_n1733) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1048 ( .A(DP_OP_423J2_125_3477_n1836), .B(
        DP_OP_423J2_125_3477_n1737), .CI(DP_OP_423J2_125_3477_n1735), .CO(
        DP_OP_423J2_125_3477_n1730), .S(DP_OP_423J2_125_3477_n1731) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1046 ( .A(DP_OP_423J2_125_3477_n2505), .B(
        DP_OP_423J2_125_3477_n1977), .CI(DP_OP_423J2_125_3477_n1933), .CO(
        DP_OP_423J2_125_3477_n1726), .S(DP_OP_423J2_125_3477_n1727) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1045 ( .A(DP_OP_423J2_125_3477_n2197), .B(
        DP_OP_423J2_125_3477_n2637), .CI(DP_OP_423J2_125_3477_n2417), .CO(
        DP_OP_423J2_125_3477_n1724), .S(DP_OP_423J2_125_3477_n1725) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1044 ( .A(DP_OP_423J2_125_3477_n2945), .B(
        DP_OP_423J2_125_3477_n2153), .CI(DP_OP_423J2_125_3477_n2373), .CO(
        DP_OP_423J2_125_3477_n1722), .S(DP_OP_423J2_125_3477_n1723) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1043 ( .A(DP_OP_423J2_125_3477_n2549), .B(
        DP_OP_423J2_125_3477_n2857), .CI(DP_OP_423J2_125_3477_n2461), .CO(
        DP_OP_423J2_125_3477_n1720), .S(DP_OP_423J2_125_3477_n1721) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1042 ( .A(DP_OP_423J2_125_3477_n2285), .B(
        DP_OP_423J2_125_3477_n2329), .CI(DP_OP_423J2_125_3477_n2109), .CO(
        DP_OP_423J2_125_3477_n1718), .S(DP_OP_423J2_125_3477_n1719) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1041 ( .A(DP_OP_423J2_125_3477_n2813), .B(
        DP_OP_423J2_125_3477_n2681), .CI(DP_OP_423J2_125_3477_n2725), .CO(
        DP_OP_423J2_125_3477_n1716), .S(DP_OP_423J2_125_3477_n1717) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1039 ( .A(DP_OP_423J2_125_3477_n2593), .B(
        DP_OP_423J2_125_3477_n2989), .CI(DP_OP_423J2_125_3477_n2241), .CO(
        DP_OP_423J2_125_3477_n1712), .S(DP_OP_423J2_125_3477_n1713) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1038 ( .A(DP_OP_423J2_125_3477_n1729), .B(
        DP_OP_423J2_125_3477_n2021), .CI(DP_OP_423J2_125_3477_n1998), .CO(
        DP_OP_423J2_125_3477_n1710), .S(DP_OP_423J2_125_3477_n1711) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1037 ( .A(DP_OP_423J2_125_3477_n2028), .B(
        DP_OP_423J2_125_3477_n1991), .CI(DP_OP_423J2_125_3477_n1984), .CO(
        DP_OP_423J2_125_3477_n1708), .S(DP_OP_423J2_125_3477_n1709) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1036 ( .A(DP_OP_423J2_125_3477_n2042), .B(
        DP_OP_423J2_125_3477_n2035), .CI(DP_OP_423J2_125_3477_n2072), .CO(
        DP_OP_423J2_125_3477_n1706), .S(DP_OP_423J2_125_3477_n1707) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1035 ( .A(DP_OP_423J2_125_3477_n2086), .B(
        DP_OP_423J2_125_3477_n2079), .CI(DP_OP_423J2_125_3477_n2116), .CO(
        DP_OP_423J2_125_3477_n1704), .S(DP_OP_423J2_125_3477_n1705) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1034 ( .A(DP_OP_423J2_125_3477_n3052), .B(
        DP_OP_423J2_125_3477_n2123), .CI(DP_OP_423J2_125_3477_n2130), .CO(
        DP_OP_423J2_125_3477_n1702), .S(DP_OP_423J2_125_3477_n1703) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1033 ( .A(DP_OP_423J2_125_3477_n2563), .B(
        DP_OP_423J2_125_3477_n3045), .CI(DP_OP_423J2_125_3477_n3038), .CO(
        DP_OP_423J2_125_3477_n1700), .S(DP_OP_423J2_125_3477_n1701) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1032 ( .A(DP_OP_423J2_125_3477_n2526), .B(
        DP_OP_423J2_125_3477_n2160), .CI(DP_OP_423J2_125_3477_n3010), .CO(
        DP_OP_423J2_125_3477_n1698), .S(DP_OP_423J2_125_3477_n1699) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1031 ( .A(DP_OP_423J2_125_3477_n2556), .B(
        DP_OP_423J2_125_3477_n2167), .CI(DP_OP_423J2_125_3477_n3003), .CO(
        DP_OP_423J2_125_3477_n1696), .S(DP_OP_423J2_125_3477_n1697) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1030 ( .A(DP_OP_423J2_125_3477_n2996), .B(
        DP_OP_423J2_125_3477_n2174), .CI(DP_OP_423J2_125_3477_n2204), .CO(
        DP_OP_423J2_125_3477_n1694), .S(DP_OP_423J2_125_3477_n1695) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1029 ( .A(DP_OP_423J2_125_3477_n2519), .B(
        DP_OP_423J2_125_3477_n2211), .CI(DP_OP_423J2_125_3477_n2218), .CO(
        DP_OP_423J2_125_3477_n1692), .S(DP_OP_423J2_125_3477_n1693) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1028 ( .A(DP_OP_423J2_125_3477_n2600), .B(
        DP_OP_423J2_125_3477_n2248), .CI(DP_OP_423J2_125_3477_n2255), .CO(
        DP_OP_423J2_125_3477_n1690), .S(DP_OP_423J2_125_3477_n1691) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1027 ( .A(DP_OP_423J2_125_3477_n2607), .B(
        DP_OP_423J2_125_3477_n2262), .CI(DP_OP_423J2_125_3477_n2292), .CO(
        DP_OP_423J2_125_3477_n1688), .S(DP_OP_423J2_125_3477_n1689) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1026 ( .A(DP_OP_423J2_125_3477_n2614), .B(
        DP_OP_423J2_125_3477_n2966), .CI(DP_OP_423J2_125_3477_n2299), .CO(
        DP_OP_423J2_125_3477_n1686), .S(DP_OP_423J2_125_3477_n1687) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1025 ( .A(DP_OP_423J2_125_3477_n2644), .B(
        DP_OP_423J2_125_3477_n2306), .CI(DP_OP_423J2_125_3477_n2959), .CO(
        DP_OP_423J2_125_3477_n1684), .S(DP_OP_423J2_125_3477_n1685) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1024 ( .A(DP_OP_423J2_125_3477_n2570), .B(
        DP_OP_423J2_125_3477_n2952), .CI(DP_OP_423J2_125_3477_n2922), .CO(
        DP_OP_423J2_125_3477_n1682), .S(DP_OP_423J2_125_3477_n1683) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1023 ( .A(DP_OP_423J2_125_3477_n2482), .B(
        DP_OP_423J2_125_3477_n2915), .CI(DP_OP_423J2_125_3477_n2336), .CO(
        DP_OP_423J2_125_3477_n1680), .S(DP_OP_423J2_125_3477_n1681) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1022 ( .A(DP_OP_423J2_125_3477_n2908), .B(
        DP_OP_423J2_125_3477_n2343), .CI(DP_OP_423J2_125_3477_n2878), .CO(
        DP_OP_423J2_125_3477_n1678), .S(DP_OP_423J2_125_3477_n1679) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1021 ( .A(DP_OP_423J2_125_3477_n2871), .B(
        DP_OP_423J2_125_3477_n2864), .CI(DP_OP_423J2_125_3477_n2350), .CO(
        DP_OP_423J2_125_3477_n1676), .S(DP_OP_423J2_125_3477_n1677) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1020 ( .A(DP_OP_423J2_125_3477_n2475), .B(
        DP_OP_423J2_125_3477_n2380), .CI(DP_OP_423J2_125_3477_n2834), .CO(
        DP_OP_423J2_125_3477_n1674), .S(DP_OP_423J2_125_3477_n1675) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1019 ( .A(DP_OP_423J2_125_3477_n2468), .B(
        DP_OP_423J2_125_3477_n2827), .CI(DP_OP_423J2_125_3477_n2820), .CO(
        DP_OP_423J2_125_3477_n1672), .S(DP_OP_423J2_125_3477_n1673) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1018 ( .A(DP_OP_423J2_125_3477_n2424), .B(
        DP_OP_423J2_125_3477_n2790), .CI(DP_OP_423J2_125_3477_n2783), .CO(
        DP_OP_423J2_125_3477_n1670), .S(DP_OP_423J2_125_3477_n1671) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1017 ( .A(DP_OP_423J2_125_3477_n2387), .B(
        DP_OP_423J2_125_3477_n2776), .CI(DP_OP_423J2_125_3477_n2746), .CO(
        DP_OP_423J2_125_3477_n1668), .S(DP_OP_423J2_125_3477_n1669) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1016 ( .A(DP_OP_423J2_125_3477_n2658), .B(
        DP_OP_423J2_125_3477_n2739), .CI(DP_OP_423J2_125_3477_n2394), .CO(
        DP_OP_423J2_125_3477_n1666), .S(DP_OP_423J2_125_3477_n1667) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1015 ( .A(DP_OP_423J2_125_3477_n2512), .B(
        DP_OP_423J2_125_3477_n2431), .CI(DP_OP_423J2_125_3477_n2732), .CO(
        DP_OP_423J2_125_3477_n1664), .S(DP_OP_423J2_125_3477_n1665) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1014 ( .A(DP_OP_423J2_125_3477_n2702), .B(
        DP_OP_423J2_125_3477_n2438), .CI(DP_OP_423J2_125_3477_n2651), .CO(
        DP_OP_423J2_125_3477_n1662), .S(DP_OP_423J2_125_3477_n1663) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1013 ( .A(DP_OP_423J2_125_3477_n2695), .B(
        DP_OP_423J2_125_3477_n2688), .CI(DP_OP_423J2_125_3477_n1834), .CO(
        DP_OP_423J2_125_3477_n1660), .S(DP_OP_423J2_125_3477_n1661) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1012 ( .A(DP_OP_423J2_125_3477_n1810), .B(
        DP_OP_423J2_125_3477_n1832), .CI(DP_OP_423J2_125_3477_n1786), .CO(
        DP_OP_423J2_125_3477_n1658), .S(DP_OP_423J2_125_3477_n1659) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1010 ( .A(DP_OP_423J2_125_3477_n1802), .B(
        DP_OP_423J2_125_3477_n1826), .CI(DP_OP_423J2_125_3477_n1824), .CO(
        DP_OP_423J2_125_3477_n1654), .S(DP_OP_423J2_125_3477_n1655) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1009 ( .A(DP_OP_423J2_125_3477_n1790), .B(
        DP_OP_423J2_125_3477_n1798), .CI(DP_OP_423J2_125_3477_n1788), .CO(
        DP_OP_423J2_125_3477_n1652), .S(DP_OP_423J2_125_3477_n1653) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1008 ( .A(DP_OP_423J2_125_3477_n1792), .B(
        DP_OP_423J2_125_3477_n1822), .CI(DP_OP_423J2_125_3477_n1796), .CO(
        DP_OP_423J2_125_3477_n1650), .S(DP_OP_423J2_125_3477_n1651) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1007 ( .A(DP_OP_423J2_125_3477_n1794), .B(
        DP_OP_423J2_125_3477_n1820), .CI(DP_OP_423J2_125_3477_n1818), .CO(
        DP_OP_423J2_125_3477_n1648), .S(DP_OP_423J2_125_3477_n1649) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1006 ( .A(DP_OP_423J2_125_3477_n1806), .B(
        DP_OP_423J2_125_3477_n1816), .CI(DP_OP_423J2_125_3477_n1800), .CO(
        DP_OP_423J2_125_3477_n1646), .S(DP_OP_423J2_125_3477_n1647) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1005 ( .A(DP_OP_423J2_125_3477_n1814), .B(
        DP_OP_423J2_125_3477_n1804), .CI(DP_OP_423J2_125_3477_n1812), .CO(
        DP_OP_423J2_125_3477_n1644), .S(DP_OP_423J2_125_3477_n1645) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1004 ( .A(DP_OP_423J2_125_3477_n1723), .B(
        DP_OP_423J2_125_3477_n1711), .CI(DP_OP_423J2_125_3477_n1725), .CO(
        DP_OP_423J2_125_3477_n1642), .S(DP_OP_423J2_125_3477_n1643) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1003 ( .A(DP_OP_423J2_125_3477_n1717), .B(
        DP_OP_423J2_125_3477_n1719), .CI(DP_OP_423J2_125_3477_n1784), .CO(
        DP_OP_423J2_125_3477_n1640), .S(DP_OP_423J2_125_3477_n1641) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1002 ( .A(DP_OP_423J2_125_3477_n1713), .B(
        DP_OP_423J2_125_3477_n1715), .CI(DP_OP_423J2_125_3477_n1721), .CO(
        DP_OP_423J2_125_3477_n1638), .S(DP_OP_423J2_125_3477_n1639) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1001 ( .A(DP_OP_423J2_125_3477_n1727), .B(
        DP_OP_423J2_125_3477_n1677), .CI(DP_OP_423J2_125_3477_n1675), .CO(
        DP_OP_423J2_125_3477_n1636), .S(DP_OP_423J2_125_3477_n1637) );
  FADDX1_HVT DP_OP_423J2_125_3477_U1000 ( .A(DP_OP_423J2_125_3477_n1679), .B(
        DP_OP_423J2_125_3477_n1695), .CI(DP_OP_423J2_125_3477_n1703), .CO(
        DP_OP_423J2_125_3477_n1634), .S(DP_OP_423J2_125_3477_n1635) );
  FADDX1_HVT DP_OP_423J2_125_3477_U999 ( .A(DP_OP_423J2_125_3477_n1671), .B(
        DP_OP_423J2_125_3477_n1691), .CI(DP_OP_423J2_125_3477_n1689), .CO(
        DP_OP_423J2_125_3477_n1632), .S(DP_OP_423J2_125_3477_n1633) );
  FADDX1_HVT DP_OP_423J2_125_3477_U998 ( .A(DP_OP_423J2_125_3477_n1669), .B(
        DP_OP_423J2_125_3477_n1705), .CI(DP_OP_423J2_125_3477_n1693), .CO(
        DP_OP_423J2_125_3477_n1630), .S(DP_OP_423J2_125_3477_n1631) );
  FADDX1_HVT DP_OP_423J2_125_3477_U997 ( .A(DP_OP_423J2_125_3477_n1667), .B(
        DP_OP_423J2_125_3477_n1699), .CI(DP_OP_423J2_125_3477_n1701), .CO(
        DP_OP_423J2_125_3477_n1628), .S(DP_OP_423J2_125_3477_n1629) );
  FADDX1_HVT DP_OP_423J2_125_3477_U996 ( .A(DP_OP_423J2_125_3477_n1665), .B(
        DP_OP_423J2_125_3477_n1697), .CI(DP_OP_423J2_125_3477_n1709), .CO(
        DP_OP_423J2_125_3477_n1626), .S(DP_OP_423J2_125_3477_n1627) );
  FADDX1_HVT DP_OP_423J2_125_3477_U995 ( .A(DP_OP_423J2_125_3477_n1687), .B(
        DP_OP_423J2_125_3477_n1707), .CI(DP_OP_423J2_125_3477_n1663), .CO(
        DP_OP_423J2_125_3477_n1624), .S(DP_OP_423J2_125_3477_n1625) );
  FADDX1_HVT DP_OP_423J2_125_3477_U994 ( .A(DP_OP_423J2_125_3477_n1673), .B(
        DP_OP_423J2_125_3477_n1683), .CI(DP_OP_423J2_125_3477_n1685), .CO(
        DP_OP_423J2_125_3477_n1622), .S(DP_OP_423J2_125_3477_n1623) );
  FADDX1_HVT DP_OP_423J2_125_3477_U993 ( .A(DP_OP_423J2_125_3477_n1681), .B(
        DP_OP_423J2_125_3477_n1661), .CI(DP_OP_423J2_125_3477_n1782), .CO(
        DP_OP_423J2_125_3477_n1620), .S(DP_OP_423J2_125_3477_n1621) );
  FADDX1_HVT DP_OP_423J2_125_3477_U992 ( .A(DP_OP_423J2_125_3477_n1780), .B(
        DP_OP_423J2_125_3477_n1778), .CI(DP_OP_423J2_125_3477_n1776), .CO(
        DP_OP_423J2_125_3477_n1618), .S(DP_OP_423J2_125_3477_n1619) );
  FADDX1_HVT DP_OP_423J2_125_3477_U991 ( .A(DP_OP_423J2_125_3477_n1774), .B(
        DP_OP_423J2_125_3477_n1772), .CI(DP_OP_423J2_125_3477_n1760), .CO(
        DP_OP_423J2_125_3477_n1616), .S(DP_OP_423J2_125_3477_n1617) );
  FADDX1_HVT DP_OP_423J2_125_3477_U990 ( .A(DP_OP_423J2_125_3477_n1758), .B(
        DP_OP_423J2_125_3477_n1659), .CI(DP_OP_423J2_125_3477_n1756), .CO(
        DP_OP_423J2_125_3477_n1614), .S(DP_OP_423J2_125_3477_n1615) );
  FADDX1_HVT DP_OP_423J2_125_3477_U989 ( .A(DP_OP_423J2_125_3477_n1770), .B(
        DP_OP_423J2_125_3477_n1649), .CI(DP_OP_423J2_125_3477_n1657), .CO(
        DP_OP_423J2_125_3477_n1612), .S(DP_OP_423J2_125_3477_n1613) );
  FADDX1_HVT DP_OP_423J2_125_3477_U988 ( .A(DP_OP_423J2_125_3477_n1768), .B(
        DP_OP_423J2_125_3477_n1647), .CI(DP_OP_423J2_125_3477_n1651), .CO(
        DP_OP_423J2_125_3477_n1610), .S(DP_OP_423J2_125_3477_n1611) );
  FADDX1_HVT DP_OP_423J2_125_3477_U987 ( .A(DP_OP_423J2_125_3477_n1764), .B(
        DP_OP_423J2_125_3477_n1655), .CI(DP_OP_423J2_125_3477_n1653), .CO(
        DP_OP_423J2_125_3477_n1608), .S(DP_OP_423J2_125_3477_n1609) );
  FADDX1_HVT DP_OP_423J2_125_3477_U986 ( .A(DP_OP_423J2_125_3477_n1762), .B(
        DP_OP_423J2_125_3477_n1766), .CI(DP_OP_423J2_125_3477_n1645), .CO(
        DP_OP_423J2_125_3477_n1606), .S(DP_OP_423J2_125_3477_n1607) );
  FADDX1_HVT DP_OP_423J2_125_3477_U985 ( .A(DP_OP_423J2_125_3477_n1641), .B(
        DP_OP_423J2_125_3477_n1643), .CI(DP_OP_423J2_125_3477_n1637), .CO(
        DP_OP_423J2_125_3477_n1604), .S(DP_OP_423J2_125_3477_n1605) );
  FADDX1_HVT DP_OP_423J2_125_3477_U984 ( .A(DP_OP_423J2_125_3477_n1639), .B(
        DP_OP_423J2_125_3477_n1625), .CI(DP_OP_423J2_125_3477_n1627), .CO(
        DP_OP_423J2_125_3477_n1602), .S(DP_OP_423J2_125_3477_n1603) );
  FADDX1_HVT DP_OP_423J2_125_3477_U983 ( .A(DP_OP_423J2_125_3477_n1633), .B(
        DP_OP_423J2_125_3477_n1631), .CI(DP_OP_423J2_125_3477_n1754), .CO(
        DP_OP_423J2_125_3477_n1600), .S(DP_OP_423J2_125_3477_n1601) );
  FADDX1_HVT DP_OP_423J2_125_3477_U982 ( .A(DP_OP_423J2_125_3477_n1629), .B(
        DP_OP_423J2_125_3477_n1623), .CI(DP_OP_423J2_125_3477_n1635), .CO(
        DP_OP_423J2_125_3477_n1598), .S(DP_OP_423J2_125_3477_n1599) );
  FADDX1_HVT DP_OP_423J2_125_3477_U981 ( .A(DP_OP_423J2_125_3477_n1621), .B(
        DP_OP_423J2_125_3477_n1752), .CI(DP_OP_423J2_125_3477_n1748), .CO(
        DP_OP_423J2_125_3477_n1596), .S(DP_OP_423J2_125_3477_n1597) );
  FADDX1_HVT DP_OP_423J2_125_3477_U980 ( .A(DP_OP_423J2_125_3477_n1750), .B(
        DP_OP_423J2_125_3477_n1619), .CI(DP_OP_423J2_125_3477_n1746), .CO(
        DP_OP_423J2_125_3477_n1594), .S(DP_OP_423J2_125_3477_n1595) );
  FADDX1_HVT DP_OP_423J2_125_3477_U979 ( .A(DP_OP_423J2_125_3477_n1617), .B(
        DP_OP_423J2_125_3477_n1607), .CI(DP_OP_423J2_125_3477_n1609), .CO(
        DP_OP_423J2_125_3477_n1592), .S(DP_OP_423J2_125_3477_n1593) );
  FADDX1_HVT DP_OP_423J2_125_3477_U978 ( .A(DP_OP_423J2_125_3477_n1744), .B(
        DP_OP_423J2_125_3477_n1742), .CI(DP_OP_423J2_125_3477_n1611), .CO(
        DP_OP_423J2_125_3477_n1590), .S(DP_OP_423J2_125_3477_n1591) );
  FADDX1_HVT DP_OP_423J2_125_3477_U977 ( .A(DP_OP_423J2_125_3477_n1615), .B(
        DP_OP_423J2_125_3477_n1613), .CI(DP_OP_423J2_125_3477_n1605), .CO(
        DP_OP_423J2_125_3477_n1588), .S(DP_OP_423J2_125_3477_n1589) );
  FADDX1_HVT DP_OP_423J2_125_3477_U976 ( .A(DP_OP_423J2_125_3477_n1740), .B(
        DP_OP_423J2_125_3477_n1603), .CI(DP_OP_423J2_125_3477_n1599), .CO(
        DP_OP_423J2_125_3477_n1586), .S(DP_OP_423J2_125_3477_n1587) );
  FADDX1_HVT DP_OP_423J2_125_3477_U975 ( .A(DP_OP_423J2_125_3477_n1601), .B(
        DP_OP_423J2_125_3477_n1738), .CI(DP_OP_423J2_125_3477_n1597), .CO(
        DP_OP_423J2_125_3477_n1584), .S(DP_OP_423J2_125_3477_n1585) );
  FADDX1_HVT DP_OP_423J2_125_3477_U974 ( .A(DP_OP_423J2_125_3477_n1736), .B(
        DP_OP_423J2_125_3477_n1595), .CI(DP_OP_423J2_125_3477_n1734), .CO(
        DP_OP_423J2_125_3477_n1582), .S(DP_OP_423J2_125_3477_n1583) );
  FADDX1_HVT DP_OP_423J2_125_3477_U973 ( .A(DP_OP_423J2_125_3477_n1593), .B(
        DP_OP_423J2_125_3477_n1591), .CI(DP_OP_423J2_125_3477_n1589), .CO(
        DP_OP_423J2_125_3477_n1580), .S(DP_OP_423J2_125_3477_n1581) );
  FADDX1_HVT DP_OP_423J2_125_3477_U972 ( .A(DP_OP_423J2_125_3477_n1587), .B(
        DP_OP_423J2_125_3477_n1732), .CI(DP_OP_423J2_125_3477_n1585), .CO(
        DP_OP_423J2_125_3477_n1578), .S(DP_OP_423J2_125_3477_n1579) );
  FADDX1_HVT DP_OP_423J2_125_3477_U971 ( .A(DP_OP_423J2_125_3477_n1730), .B(
        DP_OP_423J2_125_3477_n1583), .CI(DP_OP_423J2_125_3477_n1581), .CO(
        DP_OP_423J2_125_3477_n1576), .S(DP_OP_423J2_125_3477_n1577) );
  FADDX1_HVT DP_OP_423J2_125_3477_U970 ( .A(DP_OP_423J2_125_3477_n1728), .B(
        DP_OP_423J2_125_3477_n1976), .CI(DP_OP_423J2_125_3477_n1932), .CO(
        DP_OP_423J2_125_3477_n1574), .S(DP_OP_423J2_125_3477_n1575) );
  FADDX1_HVT DP_OP_423J2_125_3477_U969 ( .A(DP_OP_423J2_125_3477_n3031), .B(
        DP_OP_423J2_125_3477_n2548), .CI(DP_OP_423J2_125_3477_n2416), .CO(
        DP_OP_423J2_125_3477_n1572), .S(DP_OP_423J2_125_3477_n1573) );
  FADDX1_HVT DP_OP_423J2_125_3477_U968 ( .A(DP_OP_423J2_125_3477_n2944), .B(
        DP_OP_423J2_125_3477_n2680), .CI(DP_OP_423J2_125_3477_n2328), .CO(
        DP_OP_423J2_125_3477_n1570), .S(DP_OP_423J2_125_3477_n1571) );
  FADDX1_HVT DP_OP_423J2_125_3477_U967 ( .A(DP_OP_423J2_125_3477_n2108), .B(
        DP_OP_423J2_125_3477_n2636), .CI(DP_OP_423J2_125_3477_n2856), .CO(
        DP_OP_423J2_125_3477_n1568), .S(DP_OP_423J2_125_3477_n1569) );
  FADDX1_HVT DP_OP_423J2_125_3477_U966 ( .A(DP_OP_423J2_125_3477_n2196), .B(
        DP_OP_423J2_125_3477_n2372), .CI(DP_OP_423J2_125_3477_n2460), .CO(
        DP_OP_423J2_125_3477_n1566), .S(DP_OP_423J2_125_3477_n1567) );
  FADDX1_HVT DP_OP_423J2_125_3477_U965 ( .A(DP_OP_423J2_125_3477_n2812), .B(
        DP_OP_423J2_125_3477_n2284), .CI(DP_OP_423J2_125_3477_n2900), .CO(
        DP_OP_423J2_125_3477_n1564), .S(DP_OP_423J2_125_3477_n1565) );
  FADDX1_HVT DP_OP_423J2_125_3477_U964 ( .A(DP_OP_423J2_125_3477_n2152), .B(
        DP_OP_423J2_125_3477_n2504), .CI(DP_OP_423J2_125_3477_n2592), .CO(
        DP_OP_423J2_125_3477_n1562), .S(DP_OP_423J2_125_3477_n1563) );
  FADDX1_HVT DP_OP_423J2_125_3477_U963 ( .A(DP_OP_423J2_125_3477_n2988), .B(
        DP_OP_423J2_125_3477_n2724), .CI(DP_OP_423J2_125_3477_n2768), .CO(
        DP_OP_423J2_125_3477_n1560), .S(DP_OP_423J2_125_3477_n1561) );
  FADDX1_HVT DP_OP_423J2_125_3477_U962 ( .A(DP_OP_423J2_125_3477_n2064), .B(
        DP_OP_423J2_125_3477_n2240), .CI(DP_OP_423J2_125_3477_n2020), .CO(
        DP_OP_423J2_125_3477_n1558), .S(DP_OP_423J2_125_3477_n1559) );
  FADDX1_HVT DP_OP_423J2_125_3477_U961 ( .A(DP_OP_423J2_125_3477_n2555), .B(
        DP_OP_423J2_125_3477_n1990), .CI(DP_OP_423J2_125_3477_n1983), .CO(
        DP_OP_423J2_125_3477_n1556), .S(DP_OP_423J2_125_3477_n1557) );
  FADDX1_HVT DP_OP_423J2_125_3477_U960 ( .A(DP_OP_423J2_125_3477_n3051), .B(
        DP_OP_423J2_125_3477_n1997), .CI(DP_OP_423J2_125_3477_n2027), .CO(
        DP_OP_423J2_125_3477_n1554), .S(DP_OP_423J2_125_3477_n1555) );
  FADDX1_HVT DP_OP_423J2_125_3477_U959 ( .A(DP_OP_423J2_125_3477_n2437), .B(
        DP_OP_423J2_125_3477_n3044), .CI(DP_OP_423J2_125_3477_n2034), .CO(
        DP_OP_423J2_125_3477_n1552), .S(DP_OP_423J2_125_3477_n1553) );
  FADDX1_HVT DP_OP_423J2_125_3477_U958 ( .A(DP_OP_423J2_125_3477_n2430), .B(
        DP_OP_423J2_125_3477_n3037), .CI(DP_OP_423J2_125_3477_n2041), .CO(
        DP_OP_423J2_125_3477_n1550), .S(DP_OP_423J2_125_3477_n1551) );
  FADDX1_HVT DP_OP_423J2_125_3477_U957 ( .A(DP_OP_423J2_125_3477_n3009), .B(
        DP_OP_423J2_125_3477_n2071), .CI(DP_OP_423J2_125_3477_n2078), .CO(
        DP_OP_423J2_125_3477_n1548), .S(DP_OP_423J2_125_3477_n1549) );
  FADDX1_HVT DP_OP_423J2_125_3477_U956 ( .A(DP_OP_423J2_125_3477_n2467), .B(
        DP_OP_423J2_125_3477_n3002), .CI(DP_OP_423J2_125_3477_n2995), .CO(
        DP_OP_423J2_125_3477_n1546), .S(DP_OP_423J2_125_3477_n1547) );
  FADDX1_HVT DP_OP_423J2_125_3477_U955 ( .A(DP_OP_423J2_125_3477_n2393), .B(
        DP_OP_423J2_125_3477_n2965), .CI(DP_OP_423J2_125_3477_n2958), .CO(
        DP_OP_423J2_125_3477_n1544), .S(DP_OP_423J2_125_3477_n1545) );
  FADDX1_HVT DP_OP_423J2_125_3477_U954 ( .A(DP_OP_423J2_125_3477_n2386), .B(
        DP_OP_423J2_125_3477_n2951), .CI(DP_OP_423J2_125_3477_n2085), .CO(
        DP_OP_423J2_125_3477_n1542), .S(DP_OP_423J2_125_3477_n1543) );
  FADDX1_HVT DP_OP_423J2_125_3477_U953 ( .A(DP_OP_423J2_125_3477_n2379), .B(
        DP_OP_423J2_125_3477_n2921), .CI(DP_OP_423J2_125_3477_n2914), .CO(
        DP_OP_423J2_125_3477_n1540), .S(DP_OP_423J2_125_3477_n1541) );
  FADDX1_HVT DP_OP_423J2_125_3477_U952 ( .A(DP_OP_423J2_125_3477_n2349), .B(
        DP_OP_423J2_125_3477_n2907), .CI(DP_OP_423J2_125_3477_n2115), .CO(
        DP_OP_423J2_125_3477_n1538), .S(DP_OP_423J2_125_3477_n1539) );
  FADDX1_HVT DP_OP_423J2_125_3477_U951 ( .A(DP_OP_423J2_125_3477_n2342), .B(
        DP_OP_423J2_125_3477_n2122), .CI(DP_OP_423J2_125_3477_n2129), .CO(
        DP_OP_423J2_125_3477_n1536), .S(DP_OP_423J2_125_3477_n1537) );
  FADDX1_HVT DP_OP_423J2_125_3477_U950 ( .A(DP_OP_423J2_125_3477_n2423), .B(
        DP_OP_423J2_125_3477_n2159), .CI(DP_OP_423J2_125_3477_n2877), .CO(
        DP_OP_423J2_125_3477_n1534), .S(DP_OP_423J2_125_3477_n1535) );
  FADDX1_HVT DP_OP_423J2_125_3477_U949 ( .A(DP_OP_423J2_125_3477_n2474), .B(
        DP_OP_423J2_125_3477_n2870), .CI(DP_OP_423J2_125_3477_n2863), .CO(
        DP_OP_423J2_125_3477_n1532), .S(DP_OP_423J2_125_3477_n1533) );
  FADDX1_HVT DP_OP_423J2_125_3477_U948 ( .A(DP_OP_423J2_125_3477_n2833), .B(
        DP_OP_423J2_125_3477_n2166), .CI(DP_OP_423J2_125_3477_n2173), .CO(
        DP_OP_423J2_125_3477_n1530), .S(DP_OP_423J2_125_3477_n1531) );
  FADDX1_HVT DP_OP_423J2_125_3477_U947 ( .A(DP_OP_423J2_125_3477_n2606), .B(
        DP_OP_423J2_125_3477_n2203), .CI(DP_OP_423J2_125_3477_n2210), .CO(
        DP_OP_423J2_125_3477_n1528), .S(DP_OP_423J2_125_3477_n1529) );
  FADDX1_HVT DP_OP_423J2_125_3477_U946 ( .A(DP_OP_423J2_125_3477_n2826), .B(
        DP_OP_423J2_125_3477_n2217), .CI(DP_OP_423J2_125_3477_n2247), .CO(
        DP_OP_423J2_125_3477_n1526), .S(DP_OP_423J2_125_3477_n1527) );
  FADDX1_HVT DP_OP_423J2_125_3477_U945 ( .A(DP_OP_423J2_125_3477_n2819), .B(
        DP_OP_423J2_125_3477_n2254), .CI(DP_OP_423J2_125_3477_n2261), .CO(
        DP_OP_423J2_125_3477_n1524), .S(DP_OP_423J2_125_3477_n1525) );
  FADDX1_HVT DP_OP_423J2_125_3477_U944 ( .A(DP_OP_423J2_125_3477_n2789), .B(
        DP_OP_423J2_125_3477_n2291), .CI(DP_OP_423J2_125_3477_n2298), .CO(
        DP_OP_423J2_125_3477_n1522), .S(DP_OP_423J2_125_3477_n1523) );
  FADDX1_HVT DP_OP_423J2_125_3477_U943 ( .A(DP_OP_423J2_125_3477_n2782), .B(
        DP_OP_423J2_125_3477_n2305), .CI(DP_OP_423J2_125_3477_n2335), .CO(
        DP_OP_423J2_125_3477_n1520), .S(DP_OP_423J2_125_3477_n1521) );
  FADDX1_HVT DP_OP_423J2_125_3477_U942 ( .A(DP_OP_423J2_125_3477_n2775), .B(
        DP_OP_423J2_125_3477_n2481), .CI(DP_OP_423J2_125_3477_n2511), .CO(
        DP_OP_423J2_125_3477_n1518), .S(DP_OP_423J2_125_3477_n1519) );
  FADDX1_HVT DP_OP_423J2_125_3477_U941 ( .A(DP_OP_423J2_125_3477_n2745), .B(
        DP_OP_423J2_125_3477_n2518), .CI(DP_OP_423J2_125_3477_n2738), .CO(
        DP_OP_423J2_125_3477_n1516), .S(DP_OP_423J2_125_3477_n1517) );
  FADDX1_HVT DP_OP_423J2_125_3477_U940 ( .A(DP_OP_423J2_125_3477_n2643), .B(
        DP_OP_423J2_125_3477_n2525), .CI(DP_OP_423J2_125_3477_n2562), .CO(
        DP_OP_423J2_125_3477_n1514), .S(DP_OP_423J2_125_3477_n1515) );
  FADDX1_HVT DP_OP_423J2_125_3477_U939 ( .A(DP_OP_423J2_125_3477_n2613), .B(
        DP_OP_423J2_125_3477_n2569), .CI(DP_OP_423J2_125_3477_n2731), .CO(
        DP_OP_423J2_125_3477_n1512), .S(DP_OP_423J2_125_3477_n1513) );
  FADDX1_HVT DP_OP_423J2_125_3477_U938 ( .A(DP_OP_423J2_125_3477_n2687), .B(
        DP_OP_423J2_125_3477_n2599), .CI(DP_OP_423J2_125_3477_n2701), .CO(
        DP_OP_423J2_125_3477_n1510), .S(DP_OP_423J2_125_3477_n1511) );
  FADDX1_HVT DP_OP_423J2_125_3477_U937 ( .A(DP_OP_423J2_125_3477_n2650), .B(
        DP_OP_423J2_125_3477_n2657), .CI(DP_OP_423J2_125_3477_n2694), .CO(
        DP_OP_423J2_125_3477_n1508), .S(DP_OP_423J2_125_3477_n1509) );
  FADDX1_HVT DP_OP_423J2_125_3477_U936 ( .A(DP_OP_423J2_125_3477_n1716), .B(
        DP_OP_423J2_125_3477_n1712), .CI(DP_OP_423J2_125_3477_n1710), .CO(
        DP_OP_423J2_125_3477_n1506), .S(DP_OP_423J2_125_3477_n1507) );
  FADDX1_HVT DP_OP_423J2_125_3477_U935 ( .A(DP_OP_423J2_125_3477_n1714), .B(
        DP_OP_423J2_125_3477_n1718), .CI(DP_OP_423J2_125_3477_n1720), .CO(
        DP_OP_423J2_125_3477_n1504), .S(DP_OP_423J2_125_3477_n1505) );
  FADDX1_HVT DP_OP_423J2_125_3477_U934 ( .A(DP_OP_423J2_125_3477_n1722), .B(
        DP_OP_423J2_125_3477_n1724), .CI(DP_OP_423J2_125_3477_n1726), .CO(
        DP_OP_423J2_125_3477_n1502), .S(DP_OP_423J2_125_3477_n1503) );
  FADDX1_HVT DP_OP_423J2_125_3477_U933 ( .A(DP_OP_423J2_125_3477_n1686), .B(
        DP_OP_423J2_125_3477_n1708), .CI(DP_OP_423J2_125_3477_n1706), .CO(
        DP_OP_423J2_125_3477_n1500), .S(DP_OP_423J2_125_3477_n1501) );
  FADDX1_HVT DP_OP_423J2_125_3477_U932 ( .A(DP_OP_423J2_125_3477_n1682), .B(
        DP_OP_423J2_125_3477_n1704), .CI(DP_OP_423J2_125_3477_n1702), .CO(
        DP_OP_423J2_125_3477_n1498), .S(DP_OP_423J2_125_3477_n1499) );
  FADDX1_HVT DP_OP_423J2_125_3477_U931 ( .A(DP_OP_423J2_125_3477_n1676), .B(
        DP_OP_423J2_125_3477_n1700), .CI(DP_OP_423J2_125_3477_n1698), .CO(
        DP_OP_423J2_125_3477_n1496), .S(DP_OP_423J2_125_3477_n1497) );
  FADDX1_HVT DP_OP_423J2_125_3477_U930 ( .A(DP_OP_423J2_125_3477_n1672), .B(
        DP_OP_423J2_125_3477_n1696), .CI(DP_OP_423J2_125_3477_n1662), .CO(
        DP_OP_423J2_125_3477_n1494), .S(DP_OP_423J2_125_3477_n1495) );
  FADDX1_HVT DP_OP_423J2_125_3477_U928 ( .A(DP_OP_423J2_125_3477_n1678), .B(
        DP_OP_423J2_125_3477_n1690), .CI(DP_OP_423J2_125_3477_n1688), .CO(
        DP_OP_423J2_125_3477_n1490), .S(DP_OP_423J2_125_3477_n1491) );
  FADDX1_HVT DP_OP_423J2_125_3477_U927 ( .A(DP_OP_423J2_125_3477_n1670), .B(
        DP_OP_423J2_125_3477_n1684), .CI(DP_OP_423J2_125_3477_n1680), .CO(
        DP_OP_423J2_125_3477_n1488), .S(DP_OP_423J2_125_3477_n1489) );
  FADDX1_HVT DP_OP_423J2_125_3477_U926 ( .A(DP_OP_423J2_125_3477_n1666), .B(
        DP_OP_423J2_125_3477_n1674), .CI(DP_OP_423J2_125_3477_n1664), .CO(
        DP_OP_423J2_125_3477_n1486), .S(DP_OP_423J2_125_3477_n1487) );
  FADDX1_HVT DP_OP_423J2_125_3477_U925 ( .A(DP_OP_423J2_125_3477_n1575), .B(
        DP_OP_423J2_125_3477_n1559), .CI(DP_OP_423J2_125_3477_n1660), .CO(
        DP_OP_423J2_125_3477_n1484), .S(DP_OP_423J2_125_3477_n1485) );
  FADDX1_HVT DP_OP_423J2_125_3477_U924 ( .A(DP_OP_423J2_125_3477_n1573), .B(
        DP_OP_423J2_125_3477_n1561), .CI(DP_OP_423J2_125_3477_n1563), .CO(
        DP_OP_423J2_125_3477_n1482), .S(DP_OP_423J2_125_3477_n1483) );
  FADDX1_HVT DP_OP_423J2_125_3477_U923 ( .A(DP_OP_423J2_125_3477_n1569), .B(
        DP_OP_423J2_125_3477_n1567), .CI(DP_OP_423J2_125_3477_n1571), .CO(
        DP_OP_423J2_125_3477_n1480), .S(DP_OP_423J2_125_3477_n1481) );
  FADDX1_HVT DP_OP_423J2_125_3477_U922 ( .A(DP_OP_423J2_125_3477_n1565), .B(
        DP_OP_423J2_125_3477_n1545), .CI(DP_OP_423J2_125_3477_n1549), .CO(
        DP_OP_423J2_125_3477_n1478), .S(DP_OP_423J2_125_3477_n1479) );
  FADDX1_HVT DP_OP_423J2_125_3477_U921 ( .A(DP_OP_423J2_125_3477_n1547), .B(
        DP_OP_423J2_125_3477_n1555), .CI(DP_OP_423J2_125_3477_n1553), .CO(
        DP_OP_423J2_125_3477_n1476), .S(DP_OP_423J2_125_3477_n1477) );
  FADDX1_HVT DP_OP_423J2_125_3477_U920 ( .A(DP_OP_423J2_125_3477_n1557), .B(
        DP_OP_423J2_125_3477_n1535), .CI(DP_OP_423J2_125_3477_n1529), .CO(
        DP_OP_423J2_125_3477_n1474), .S(DP_OP_423J2_125_3477_n1475) );
  FADDX1_HVT DP_OP_423J2_125_3477_U919 ( .A(DP_OP_423J2_125_3477_n1537), .B(
        DP_OP_423J2_125_3477_n1533), .CI(DP_OP_423J2_125_3477_n1527), .CO(
        DP_OP_423J2_125_3477_n1472), .S(DP_OP_423J2_125_3477_n1473) );
  FADDX1_HVT DP_OP_423J2_125_3477_U918 ( .A(DP_OP_423J2_125_3477_n1539), .B(
        DP_OP_423J2_125_3477_n1513), .CI(DP_OP_423J2_125_3477_n1511), .CO(
        DP_OP_423J2_125_3477_n1470), .S(DP_OP_423J2_125_3477_n1471) );
  FADDX1_HVT DP_OP_423J2_125_3477_U917 ( .A(DP_OP_423J2_125_3477_n1525), .B(
        DP_OP_423J2_125_3477_n1521), .CI(DP_OP_423J2_125_3477_n1523), .CO(
        DP_OP_423J2_125_3477_n1468), .S(DP_OP_423J2_125_3477_n1469) );
  FADDX1_HVT DP_OP_423J2_125_3477_U916 ( .A(DP_OP_423J2_125_3477_n1531), .B(
        DP_OP_423J2_125_3477_n1509), .CI(DP_OP_423J2_125_3477_n1517), .CO(
        DP_OP_423J2_125_3477_n1466), .S(DP_OP_423J2_125_3477_n1467) );
  FADDX1_HVT DP_OP_423J2_125_3477_U915 ( .A(DP_OP_423J2_125_3477_n1519), .B(
        DP_OP_423J2_125_3477_n1543), .CI(DP_OP_423J2_125_3477_n1551), .CO(
        DP_OP_423J2_125_3477_n1464), .S(DP_OP_423J2_125_3477_n1465) );
  FADDX1_HVT DP_OP_423J2_125_3477_U914 ( .A(DP_OP_423J2_125_3477_n1515), .B(
        DP_OP_423J2_125_3477_n1541), .CI(DP_OP_423J2_125_3477_n1658), .CO(
        DP_OP_423J2_125_3477_n1462), .S(DP_OP_423J2_125_3477_n1463) );
  FADDX1_HVT DP_OP_423J2_125_3477_U913 ( .A(DP_OP_423J2_125_3477_n1652), .B(
        DP_OP_423J2_125_3477_n1656), .CI(DP_OP_423J2_125_3477_n1654), .CO(
        DP_OP_423J2_125_3477_n1460), .S(DP_OP_423J2_125_3477_n1461) );
  FADDX1_HVT DP_OP_423J2_125_3477_U912 ( .A(DP_OP_423J2_125_3477_n1644), .B(
        DP_OP_423J2_125_3477_n1650), .CI(DP_OP_423J2_125_3477_n1646), .CO(
        DP_OP_423J2_125_3477_n1458), .S(DP_OP_423J2_125_3477_n1459) );
  FADDX1_HVT DP_OP_423J2_125_3477_U911 ( .A(DP_OP_423J2_125_3477_n1648), .B(
        DP_OP_423J2_125_3477_n1642), .CI(DP_OP_423J2_125_3477_n1503), .CO(
        DP_OP_423J2_125_3477_n1456), .S(DP_OP_423J2_125_3477_n1457) );
  FADDX1_HVT DP_OP_423J2_125_3477_U910 ( .A(DP_OP_423J2_125_3477_n1505), .B(
        DP_OP_423J2_125_3477_n1640), .CI(DP_OP_423J2_125_3477_n1636), .CO(
        DP_OP_423J2_125_3477_n1454), .S(DP_OP_423J2_125_3477_n1455) );
  FADDX1_HVT DP_OP_423J2_125_3477_U909 ( .A(DP_OP_423J2_125_3477_n1507), .B(
        DP_OP_423J2_125_3477_n1638), .CI(DP_OP_423J2_125_3477_n1634), .CO(
        DP_OP_423J2_125_3477_n1452), .S(DP_OP_423J2_125_3477_n1453) );
  FADDX1_HVT DP_OP_423J2_125_3477_U908 ( .A(DP_OP_423J2_125_3477_n1624), .B(
        DP_OP_423J2_125_3477_n1487), .CI(DP_OP_423J2_125_3477_n1499), .CO(
        DP_OP_423J2_125_3477_n1450), .S(DP_OP_423J2_125_3477_n1451) );
  FADDX1_HVT DP_OP_423J2_125_3477_U907 ( .A(DP_OP_423J2_125_3477_n1632), .B(
        DP_OP_423J2_125_3477_n1501), .CI(DP_OP_423J2_125_3477_n1497), .CO(
        DP_OP_423J2_125_3477_n1448), .S(DP_OP_423J2_125_3477_n1449) );
  FADDX1_HVT DP_OP_423J2_125_3477_U906 ( .A(DP_OP_423J2_125_3477_n1630), .B(
        DP_OP_423J2_125_3477_n1489), .CI(DP_OP_423J2_125_3477_n1491), .CO(
        DP_OP_423J2_125_3477_n1446), .S(DP_OP_423J2_125_3477_n1447) );
  FADDX1_HVT DP_OP_423J2_125_3477_U905 ( .A(DP_OP_423J2_125_3477_n1628), .B(
        DP_OP_423J2_125_3477_n1495), .CI(DP_OP_423J2_125_3477_n1493), .CO(
        DP_OP_423J2_125_3477_n1444), .S(DP_OP_423J2_125_3477_n1445) );
  FADDX1_HVT DP_OP_423J2_125_3477_U904 ( .A(DP_OP_423J2_125_3477_n1626), .B(
        DP_OP_423J2_125_3477_n1622), .CI(DP_OP_423J2_125_3477_n1483), .CO(
        DP_OP_423J2_125_3477_n1442), .S(DP_OP_423J2_125_3477_n1443) );
  FADDX1_HVT DP_OP_423J2_125_3477_U903 ( .A(DP_OP_423J2_125_3477_n1485), .B(
        DP_OP_423J2_125_3477_n1481), .CI(DP_OP_423J2_125_3477_n1479), .CO(
        DP_OP_423J2_125_3477_n1440), .S(DP_OP_423J2_125_3477_n1441) );
  FADDX1_HVT DP_OP_423J2_125_3477_U902 ( .A(DP_OP_423J2_125_3477_n1620), .B(
        DP_OP_423J2_125_3477_n1471), .CI(DP_OP_423J2_125_3477_n1469), .CO(
        DP_OP_423J2_125_3477_n1438), .S(DP_OP_423J2_125_3477_n1439) );
  FADDX1_HVT DP_OP_423J2_125_3477_U901 ( .A(DP_OP_423J2_125_3477_n1475), .B(
        DP_OP_423J2_125_3477_n1465), .CI(DP_OP_423J2_125_3477_n1467), .CO(
        DP_OP_423J2_125_3477_n1436), .S(DP_OP_423J2_125_3477_n1437) );
  FADDX1_HVT DP_OP_423J2_125_3477_U900 ( .A(DP_OP_423J2_125_3477_n1473), .B(
        DP_OP_423J2_125_3477_n1477), .CI(DP_OP_423J2_125_3477_n1618), .CO(
        DP_OP_423J2_125_3477_n1434), .S(DP_OP_423J2_125_3477_n1435) );
  FADDX1_HVT DP_OP_423J2_125_3477_U899 ( .A(DP_OP_423J2_125_3477_n1616), .B(
        DP_OP_423J2_125_3477_n1463), .CI(DP_OP_423J2_125_3477_n1614), .CO(
        DP_OP_423J2_125_3477_n1432), .S(DP_OP_423J2_125_3477_n1433) );
  FADDX1_HVT DP_OP_423J2_125_3477_U898 ( .A(DP_OP_423J2_125_3477_n1612), .B(
        DP_OP_423J2_125_3477_n1459), .CI(DP_OP_423J2_125_3477_n1461), .CO(
        DP_OP_423J2_125_3477_n1430), .S(DP_OP_423J2_125_3477_n1431) );
  FADDX1_HVT DP_OP_423J2_125_3477_U897 ( .A(DP_OP_423J2_125_3477_n1610), .B(
        DP_OP_423J2_125_3477_n1606), .CI(DP_OP_423J2_125_3477_n1608), .CO(
        DP_OP_423J2_125_3477_n1428), .S(DP_OP_423J2_125_3477_n1429) );
  FADDX1_HVT DP_OP_423J2_125_3477_U896 ( .A(DP_OP_423J2_125_3477_n1457), .B(
        DP_OP_423J2_125_3477_n1604), .CI(DP_OP_423J2_125_3477_n1602), .CO(
        DP_OP_423J2_125_3477_n1426), .S(DP_OP_423J2_125_3477_n1427) );
  FADDX1_HVT DP_OP_423J2_125_3477_U895 ( .A(DP_OP_423J2_125_3477_n1455), .B(
        DP_OP_423J2_125_3477_n1453), .CI(DP_OP_423J2_125_3477_n1449), .CO(
        DP_OP_423J2_125_3477_n1424), .S(DP_OP_423J2_125_3477_n1425) );
  FADDX1_HVT DP_OP_423J2_125_3477_U894 ( .A(DP_OP_423J2_125_3477_n1451), .B(
        DP_OP_423J2_125_3477_n1447), .CI(DP_OP_423J2_125_3477_n1443), .CO(
        DP_OP_423J2_125_3477_n1422), .S(DP_OP_423J2_125_3477_n1423) );
  FADDX1_HVT DP_OP_423J2_125_3477_U893 ( .A(DP_OP_423J2_125_3477_n1600), .B(
        DP_OP_423J2_125_3477_n1445), .CI(DP_OP_423J2_125_3477_n1598), .CO(
        DP_OP_423J2_125_3477_n1420), .S(DP_OP_423J2_125_3477_n1421) );
  FADDX1_HVT DP_OP_423J2_125_3477_U892 ( .A(DP_OP_423J2_125_3477_n1441), .B(
        DP_OP_423J2_125_3477_n1439), .CI(DP_OP_423J2_125_3477_n1437), .CO(
        DP_OP_423J2_125_3477_n1418), .S(DP_OP_423J2_125_3477_n1419) );
  FADDX1_HVT DP_OP_423J2_125_3477_U891 ( .A(DP_OP_423J2_125_3477_n1596), .B(
        DP_OP_423J2_125_3477_n1435), .CI(DP_OP_423J2_125_3477_n1594), .CO(
        DP_OP_423J2_125_3477_n1416), .S(DP_OP_423J2_125_3477_n1417) );
  FADDX1_HVT DP_OP_423J2_125_3477_U889 ( .A(DP_OP_423J2_125_3477_n1429), .B(
        DP_OP_423J2_125_3477_n1431), .CI(DP_OP_423J2_125_3477_n1588), .CO(
        DP_OP_423J2_125_3477_n1412), .S(DP_OP_423J2_125_3477_n1413) );
  FADDX1_HVT DP_OP_423J2_125_3477_U888 ( .A(DP_OP_423J2_125_3477_n1427), .B(
        DP_OP_423J2_125_3477_n1425), .CI(DP_OP_423J2_125_3477_n1586), .CO(
        DP_OP_423J2_125_3477_n1410), .S(DP_OP_423J2_125_3477_n1411) );
  FADDX1_HVT DP_OP_423J2_125_3477_U887 ( .A(DP_OP_423J2_125_3477_n1421), .B(
        DP_OP_423J2_125_3477_n1423), .CI(DP_OP_423J2_125_3477_n1584), .CO(
        DP_OP_423J2_125_3477_n1408), .S(DP_OP_423J2_125_3477_n1409) );
  FADDX1_HVT DP_OP_423J2_125_3477_U886 ( .A(DP_OP_423J2_125_3477_n1419), .B(
        DP_OP_423J2_125_3477_n1417), .CI(DP_OP_423J2_125_3477_n1582), .CO(
        DP_OP_423J2_125_3477_n1406), .S(DP_OP_423J2_125_3477_n1407) );
  FADDX1_HVT DP_OP_423J2_125_3477_U885 ( .A(DP_OP_423J2_125_3477_n1415), .B(
        DP_OP_423J2_125_3477_n1580), .CI(DP_OP_423J2_125_3477_n1413), .CO(
        DP_OP_423J2_125_3477_n1404), .S(DP_OP_423J2_125_3477_n1405) );
  FADDX1_HVT DP_OP_423J2_125_3477_U884 ( .A(DP_OP_423J2_125_3477_n1411), .B(
        DP_OP_423J2_125_3477_n1578), .CI(DP_OP_423J2_125_3477_n1409), .CO(
        DP_OP_423J2_125_3477_n1402), .S(DP_OP_423J2_125_3477_n1403) );
  FADDX1_HVT DP_OP_423J2_125_3477_U883 ( .A(DP_OP_423J2_125_3477_n1407), .B(
        DP_OP_423J2_125_3477_n1576), .CI(DP_OP_423J2_125_3477_n1405), .CO(
        DP_OP_423J2_125_3477_n1400), .S(DP_OP_423J2_125_3477_n1401) );
  HADDX1_HVT DP_OP_423J2_125_3477_U882 ( .A0(DP_OP_423J2_125_3477_n3030), .B0(
        DP_OP_423J2_125_3477_n1975), .C1(DP_OP_423J2_125_3477_n1398), .SO(
        DP_OP_423J2_125_3477_n1399) );
  FADDX1_HVT DP_OP_423J2_125_3477_U881 ( .A(DP_OP_423J2_125_3477_n2503), .B(
        DP_OP_423J2_125_3477_n2415), .CI(DP_OP_423J2_125_3477_n1931), .CO(
        DP_OP_423J2_125_3477_n1396), .S(DP_OP_423J2_125_3477_n1397) );
  FADDX1_HVT DP_OP_423J2_125_3477_U880 ( .A(DP_OP_423J2_125_3477_n2547), .B(
        DP_OP_423J2_125_3477_n2327), .CI(DP_OP_423J2_125_3477_n2371), .CO(
        DP_OP_423J2_125_3477_n1394), .S(DP_OP_423J2_125_3477_n1395) );
  FADDX1_HVT DP_OP_423J2_125_3477_U879 ( .A(DP_OP_423J2_125_3477_n2855), .B(
        DP_OP_423J2_125_3477_n2019), .CI(DP_OP_423J2_125_3477_n2107), .CO(
        DP_OP_423J2_125_3477_n1392), .S(DP_OP_423J2_125_3477_n1393) );
  FADDX1_HVT DP_OP_423J2_125_3477_U878 ( .A(DP_OP_423J2_125_3477_n2591), .B(
        DP_OP_423J2_125_3477_n2151), .CI(DP_OP_423J2_125_3477_n2679), .CO(
        DP_OP_423J2_125_3477_n1390), .S(DP_OP_423J2_125_3477_n1391) );
  FADDX1_HVT DP_OP_423J2_125_3477_U877 ( .A(DP_OP_423J2_125_3477_n2063), .B(
        DP_OP_423J2_125_3477_n2899), .CI(DP_OP_423J2_125_3477_n2195), .CO(
        DP_OP_423J2_125_3477_n1388), .S(DP_OP_423J2_125_3477_n1389) );
  FADDX1_HVT DP_OP_423J2_125_3477_U876 ( .A(DP_OP_423J2_125_3477_n2459), .B(
        DP_OP_423J2_125_3477_n2943), .CI(DP_OP_423J2_125_3477_n2767), .CO(
        DP_OP_423J2_125_3477_n1386), .S(DP_OP_423J2_125_3477_n1387) );
  FADDX1_HVT DP_OP_423J2_125_3477_U875 ( .A(DP_OP_423J2_125_3477_n2283), .B(
        DP_OP_423J2_125_3477_n2239), .CI(DP_OP_423J2_125_3477_n2723), .CO(
        DP_OP_423J2_125_3477_n1384), .S(DP_OP_423J2_125_3477_n1385) );
  FADDX1_HVT DP_OP_423J2_125_3477_U874 ( .A(DP_OP_423J2_125_3477_n2987), .B(
        DP_OP_423J2_125_3477_n2635), .CI(DP_OP_423J2_125_3477_n2811), .CO(
        DP_OP_423J2_125_3477_n1382), .S(DP_OP_423J2_125_3477_n1383) );
  FADDX1_HVT DP_OP_423J2_125_3477_U873 ( .A(DP_OP_423J2_125_3477_n2429), .B(
        DP_OP_423J2_125_3477_n3050), .CI(DP_OP_423J2_125_3477_n1982), .CO(
        DP_OP_423J2_125_3477_n1380), .S(DP_OP_423J2_125_3477_n1381) );
  FADDX1_HVT DP_OP_423J2_125_3477_U872 ( .A(DP_OP_423J2_125_3477_n2422), .B(
        DP_OP_423J2_125_3477_n1989), .CI(DP_OP_423J2_125_3477_n1996), .CO(
        DP_OP_423J2_125_3477_n1378), .S(DP_OP_423J2_125_3477_n1379) );
  FADDX1_HVT DP_OP_423J2_125_3477_U871 ( .A(DP_OP_423J2_125_3477_n2436), .B(
        DP_OP_423J2_125_3477_n2026), .CI(DP_OP_423J2_125_3477_n3043), .CO(
        DP_OP_423J2_125_3477_n1376), .S(DP_OP_423J2_125_3477_n1377) );
  FADDX1_HVT DP_OP_423J2_125_3477_U870 ( .A(DP_OP_423J2_125_3477_n2392), .B(
        DP_OP_423J2_125_3477_n3036), .CI(DP_OP_423J2_125_3477_n3008), .CO(
        DP_OP_423J2_125_3477_n1374), .S(DP_OP_423J2_125_3477_n1375) );
  FADDX1_HVT DP_OP_423J2_125_3477_U869 ( .A(DP_OP_423J2_125_3477_n2385), .B(
        DP_OP_423J2_125_3477_n3001), .CI(DP_OP_423J2_125_3477_n2994), .CO(
        DP_OP_423J2_125_3477_n1372), .S(DP_OP_423J2_125_3477_n1373) );
  FADDX1_HVT DP_OP_423J2_125_3477_U868 ( .A(DP_OP_423J2_125_3477_n2348), .B(
        DP_OP_423J2_125_3477_n2964), .CI(DP_OP_423J2_125_3477_n2957), .CO(
        DP_OP_423J2_125_3477_n1370), .S(DP_OP_423J2_125_3477_n1371) );
  FADDX1_HVT DP_OP_423J2_125_3477_U867 ( .A(DP_OP_423J2_125_3477_n2341), .B(
        DP_OP_423J2_125_3477_n2033), .CI(DP_OP_423J2_125_3477_n2950), .CO(
        DP_OP_423J2_125_3477_n1368), .S(DP_OP_423J2_125_3477_n1369) );
  FADDX1_HVT DP_OP_423J2_125_3477_U866 ( .A(DP_OP_423J2_125_3477_n2334), .B(
        DP_OP_423J2_125_3477_n2920), .CI(DP_OP_423J2_125_3477_n2913), .CO(
        DP_OP_423J2_125_3477_n1366), .S(DP_OP_423J2_125_3477_n1367) );
  FADDX1_HVT DP_OP_423J2_125_3477_U865 ( .A(DP_OP_423J2_125_3477_n2304), .B(
        DP_OP_423J2_125_3477_n2906), .CI(DP_OP_423J2_125_3477_n2040), .CO(
        DP_OP_423J2_125_3477_n1364), .S(DP_OP_423J2_125_3477_n1365) );
  FADDX1_HVT DP_OP_423J2_125_3477_U864 ( .A(DP_OP_423J2_125_3477_n2297), .B(
        DP_OP_423J2_125_3477_n2070), .CI(DP_OP_423J2_125_3477_n2077), .CO(
        DP_OP_423J2_125_3477_n1362), .S(DP_OP_423J2_125_3477_n1363) );
  FADDX1_HVT DP_OP_423J2_125_3477_U863 ( .A(DP_OP_423J2_125_3477_n2378), .B(
        DP_OP_423J2_125_3477_n2084), .CI(DP_OP_423J2_125_3477_n2876), .CO(
        DP_OP_423J2_125_3477_n1360), .S(DP_OP_423J2_125_3477_n1361) );
  FADDX1_HVT DP_OP_423J2_125_3477_U862 ( .A(DP_OP_423J2_125_3477_n2466), .B(
        DP_OP_423J2_125_3477_n2869), .CI(DP_OP_423J2_125_3477_n2114), .CO(
        DP_OP_423J2_125_3477_n1358), .S(DP_OP_423J2_125_3477_n1359) );
  FADDX1_HVT DP_OP_423J2_125_3477_U861 ( .A(DP_OP_423J2_125_3477_n2862), .B(
        DP_OP_423J2_125_3477_n2121), .CI(DP_OP_423J2_125_3477_n2128), .CO(
        DP_OP_423J2_125_3477_n1356), .S(DP_OP_423J2_125_3477_n1357) );
  FADDX1_HVT DP_OP_423J2_125_3477_U860 ( .A(DP_OP_423J2_125_3477_n2832), .B(
        DP_OP_423J2_125_3477_n2158), .CI(DP_OP_423J2_125_3477_n2165), .CO(
        DP_OP_423J2_125_3477_n1354), .S(DP_OP_423J2_125_3477_n1355) );
  FADDX1_HVT DP_OP_423J2_125_3477_U859 ( .A(DP_OP_423J2_125_3477_n2825), .B(
        DP_OP_423J2_125_3477_n2172), .CI(DP_OP_423J2_125_3477_n2202), .CO(
        DP_OP_423J2_125_3477_n1352), .S(DP_OP_423J2_125_3477_n1353) );
  FADDX1_HVT DP_OP_423J2_125_3477_U858 ( .A(DP_OP_423J2_125_3477_n2818), .B(
        DP_OP_423J2_125_3477_n2209), .CI(DP_OP_423J2_125_3477_n2216), .CO(
        DP_OP_423J2_125_3477_n1350), .S(DP_OP_423J2_125_3477_n1351) );
  FADDX1_HVT DP_OP_423J2_125_3477_U857 ( .A(DP_OP_423J2_125_3477_n2788), .B(
        DP_OP_423J2_125_3477_n2246), .CI(DP_OP_423J2_125_3477_n2253), .CO(
        DP_OP_423J2_125_3477_n1348), .S(DP_OP_423J2_125_3477_n1349) );
  FADDX1_HVT DP_OP_423J2_125_3477_U856 ( .A(DP_OP_423J2_125_3477_n2781), .B(
        DP_OP_423J2_125_3477_n2260), .CI(DP_OP_423J2_125_3477_n2290), .CO(
        DP_OP_423J2_125_3477_n1346), .S(DP_OP_423J2_125_3477_n1347) );
  FADDX1_HVT DP_OP_423J2_125_3477_U855 ( .A(DP_OP_423J2_125_3477_n2774), .B(
        DP_OP_423J2_125_3477_n2473), .CI(DP_OP_423J2_125_3477_n2480), .CO(
        DP_OP_423J2_125_3477_n1344), .S(DP_OP_423J2_125_3477_n1345) );
  FADDX1_HVT DP_OP_423J2_125_3477_U854 ( .A(DP_OP_423J2_125_3477_n2744), .B(
        DP_OP_423J2_125_3477_n2510), .CI(DP_OP_423J2_125_3477_n2517), .CO(
        DP_OP_423J2_125_3477_n1342), .S(DP_OP_423J2_125_3477_n1343) );
  FADDX1_HVT DP_OP_423J2_125_3477_U853 ( .A(DP_OP_423J2_125_3477_n2737), .B(
        DP_OP_423J2_125_3477_n2524), .CI(DP_OP_423J2_125_3477_n2554), .CO(
        DP_OP_423J2_125_3477_n1340), .S(DP_OP_423J2_125_3477_n1341) );
  FADDX1_HVT DP_OP_423J2_125_3477_U852 ( .A(DP_OP_423J2_125_3477_n2730), .B(
        DP_OP_423J2_125_3477_n2561), .CI(DP_OP_423J2_125_3477_n2568), .CO(
        DP_OP_423J2_125_3477_n1338), .S(DP_OP_423J2_125_3477_n1339) );
  FADDX1_HVT DP_OP_423J2_125_3477_U851 ( .A(DP_OP_423J2_125_3477_n2700), .B(
        DP_OP_423J2_125_3477_n2693), .CI(DP_OP_423J2_125_3477_n2686), .CO(
        DP_OP_423J2_125_3477_n1336), .S(DP_OP_423J2_125_3477_n1337) );
  FADDX1_HVT DP_OP_423J2_125_3477_U850 ( .A(DP_OP_423J2_125_3477_n2642), .B(
        DP_OP_423J2_125_3477_n2656), .CI(DP_OP_423J2_125_3477_n2598), .CO(
        DP_OP_423J2_125_3477_n1334), .S(DP_OP_423J2_125_3477_n1335) );
  FADDX1_HVT DP_OP_423J2_125_3477_U849 ( .A(DP_OP_423J2_125_3477_n2605), .B(
        DP_OP_423J2_125_3477_n2612), .CI(DP_OP_423J2_125_3477_n2649), .CO(
        DP_OP_423J2_125_3477_n1332), .S(DP_OP_423J2_125_3477_n1333) );
  FADDX1_HVT DP_OP_423J2_125_3477_U848 ( .A(DP_OP_423J2_125_3477_n1399), .B(
        DP_OP_423J2_125_3477_n1574), .CI(DP_OP_423J2_125_3477_n1564), .CO(
        DP_OP_423J2_125_3477_n1330), .S(DP_OP_423J2_125_3477_n1331) );
  FADDX1_HVT DP_OP_423J2_125_3477_U847 ( .A(DP_OP_423J2_125_3477_n1572), .B(
        DP_OP_423J2_125_3477_n1570), .CI(DP_OP_423J2_125_3477_n1568), .CO(
        DP_OP_423J2_125_3477_n1328), .S(DP_OP_423J2_125_3477_n1329) );
  FADDX1_HVT DP_OP_423J2_125_3477_U846 ( .A(DP_OP_423J2_125_3477_n1566), .B(
        DP_OP_423J2_125_3477_n1562), .CI(DP_OP_423J2_125_3477_n1558), .CO(
        DP_OP_423J2_125_3477_n1326), .S(DP_OP_423J2_125_3477_n1327) );
  FADDX1_HVT DP_OP_423J2_125_3477_U845 ( .A(DP_OP_423J2_125_3477_n1560), .B(
        DP_OP_423J2_125_3477_n1534), .CI(DP_OP_423J2_125_3477_n1532), .CO(
        DP_OP_423J2_125_3477_n1324), .S(DP_OP_423J2_125_3477_n1325) );
  FADDX1_HVT DP_OP_423J2_125_3477_U844 ( .A(DP_OP_423J2_125_3477_n1536), .B(
        DP_OP_423J2_125_3477_n1508), .CI(DP_OP_423J2_125_3477_n1556), .CO(
        DP_OP_423J2_125_3477_n1322), .S(DP_OP_423J2_125_3477_n1323) );
  FADDX1_HVT DP_OP_423J2_125_3477_U843 ( .A(DP_OP_423J2_125_3477_n1528), .B(
        DP_OP_423J2_125_3477_n1554), .CI(DP_OP_423J2_125_3477_n1552), .CO(
        DP_OP_423J2_125_3477_n1320), .S(DP_OP_423J2_125_3477_n1321) );
  FADDX1_HVT DP_OP_423J2_125_3477_U842 ( .A(DP_OP_423J2_125_3477_n1524), .B(
        DP_OP_423J2_125_3477_n1550), .CI(DP_OP_423J2_125_3477_n1548), .CO(
        DP_OP_423J2_125_3477_n1318), .S(DP_OP_423J2_125_3477_n1319) );
  FADDX1_HVT DP_OP_423J2_125_3477_U841 ( .A(DP_OP_423J2_125_3477_n1518), .B(
        DP_OP_423J2_125_3477_n1510), .CI(DP_OP_423J2_125_3477_n1512), .CO(
        DP_OP_423J2_125_3477_n1316), .S(DP_OP_423J2_125_3477_n1317) );
  FADDX1_HVT DP_OP_423J2_125_3477_U840 ( .A(DP_OP_423J2_125_3477_n1516), .B(
        DP_OP_423J2_125_3477_n1546), .CI(DP_OP_423J2_125_3477_n1544), .CO(
        DP_OP_423J2_125_3477_n1314), .S(DP_OP_423J2_125_3477_n1315) );
  FADDX1_HVT DP_OP_423J2_125_3477_U839 ( .A(DP_OP_423J2_125_3477_n1526), .B(
        DP_OP_423J2_125_3477_n1542), .CI(DP_OP_423J2_125_3477_n1514), .CO(
        DP_OP_423J2_125_3477_n1312), .S(DP_OP_423J2_125_3477_n1313) );
  FADDX1_HVT DP_OP_423J2_125_3477_U838 ( .A(DP_OP_423J2_125_3477_n1522), .B(
        DP_OP_423J2_125_3477_n1540), .CI(DP_OP_423J2_125_3477_n1538), .CO(
        DP_OP_423J2_125_3477_n1310), .S(DP_OP_423J2_125_3477_n1311) );
  FADDX1_HVT DP_OP_423J2_125_3477_U837 ( .A(DP_OP_423J2_125_3477_n1520), .B(
        DP_OP_423J2_125_3477_n1530), .CI(DP_OP_423J2_125_3477_n1389), .CO(
        DP_OP_423J2_125_3477_n1308), .S(DP_OP_423J2_125_3477_n1309) );
  FADDX1_HVT DP_OP_423J2_125_3477_U836 ( .A(DP_OP_423J2_125_3477_n1391), .B(
        DP_OP_423J2_125_3477_n1383), .CI(DP_OP_423J2_125_3477_n1385), .CO(
        DP_OP_423J2_125_3477_n1306), .S(DP_OP_423J2_125_3477_n1307) );
  FADDX1_HVT DP_OP_423J2_125_3477_U835 ( .A(DP_OP_423J2_125_3477_n1395), .B(
        DP_OP_423J2_125_3477_n1393), .CI(DP_OP_423J2_125_3477_n1397), .CO(
        DP_OP_423J2_125_3477_n1304), .S(DP_OP_423J2_125_3477_n1305) );
  FADDX1_HVT DP_OP_423J2_125_3477_U834 ( .A(DP_OP_423J2_125_3477_n1387), .B(
        DP_OP_423J2_125_3477_n1339), .CI(DP_OP_423J2_125_3477_n1337), .CO(
        DP_OP_423J2_125_3477_n1302), .S(DP_OP_423J2_125_3477_n1303) );
  FADDX1_HVT DP_OP_423J2_125_3477_U833 ( .A(DP_OP_423J2_125_3477_n1333), .B(
        DP_OP_423J2_125_3477_n1381), .CI(DP_OP_423J2_125_3477_n1379), .CO(
        DP_OP_423J2_125_3477_n1300), .S(DP_OP_423J2_125_3477_n1301) );
  FADDX1_HVT DP_OP_423J2_125_3477_U832 ( .A(DP_OP_423J2_125_3477_n1369), .B(
        DP_OP_423J2_125_3477_n1359), .CI(DP_OP_423J2_125_3477_n1365), .CO(
        DP_OP_423J2_125_3477_n1298), .S(DP_OP_423J2_125_3477_n1299) );
  FADDX1_HVT DP_OP_423J2_125_3477_U831 ( .A(DP_OP_423J2_125_3477_n1363), .B(
        DP_OP_423J2_125_3477_n1361), .CI(DP_OP_423J2_125_3477_n1345), .CO(
        DP_OP_423J2_125_3477_n1296), .S(DP_OP_423J2_125_3477_n1297) );
  FADDX1_HVT DP_OP_423J2_125_3477_U830 ( .A(DP_OP_423J2_125_3477_n1367), .B(
        DP_OP_423J2_125_3477_n1341), .CI(DP_OP_423J2_125_3477_n1335), .CO(
        DP_OP_423J2_125_3477_n1294), .S(DP_OP_423J2_125_3477_n1295) );
  FADDX1_HVT DP_OP_423J2_125_3477_U829 ( .A(DP_OP_423J2_125_3477_n1371), .B(
        DP_OP_423J2_125_3477_n1353), .CI(DP_OP_423J2_125_3477_n1355), .CO(
        DP_OP_423J2_125_3477_n1292), .S(DP_OP_423J2_125_3477_n1293) );
  FADDX1_HVT DP_OP_423J2_125_3477_U828 ( .A(DP_OP_423J2_125_3477_n1351), .B(
        DP_OP_423J2_125_3477_n1349), .CI(DP_OP_423J2_125_3477_n1343), .CO(
        DP_OP_423J2_125_3477_n1290), .S(DP_OP_423J2_125_3477_n1291) );
  FADDX1_HVT DP_OP_423J2_125_3477_U827 ( .A(DP_OP_423J2_125_3477_n1347), .B(
        DP_OP_423J2_125_3477_n1373), .CI(DP_OP_423J2_125_3477_n1377), .CO(
        DP_OP_423J2_125_3477_n1288), .S(DP_OP_423J2_125_3477_n1289) );
  FADDX1_HVT DP_OP_423J2_125_3477_U826 ( .A(DP_OP_423J2_125_3477_n1375), .B(
        DP_OP_423J2_125_3477_n1357), .CI(DP_OP_423J2_125_3477_n1506), .CO(
        DP_OP_423J2_125_3477_n1286), .S(DP_OP_423J2_125_3477_n1287) );
  FADDX1_HVT DP_OP_423J2_125_3477_U825 ( .A(DP_OP_423J2_125_3477_n1504), .B(
        DP_OP_423J2_125_3477_n1502), .CI(DP_OP_423J2_125_3477_n1500), .CO(
        DP_OP_423J2_125_3477_n1284), .S(DP_OP_423J2_125_3477_n1285) );
  FADDX1_HVT DP_OP_423J2_125_3477_U823 ( .A(DP_OP_423J2_125_3477_n1492), .B(
        DP_OP_423J2_125_3477_n1496), .CI(DP_OP_423J2_125_3477_n1490), .CO(
        DP_OP_423J2_125_3477_n1280), .S(DP_OP_423J2_125_3477_n1281) );
  FADDX1_HVT DP_OP_423J2_125_3477_U822 ( .A(DP_OP_423J2_125_3477_n1494), .B(
        DP_OP_423J2_125_3477_n1331), .CI(DP_OP_423J2_125_3477_n1484), .CO(
        DP_OP_423J2_125_3477_n1278), .S(DP_OP_423J2_125_3477_n1279) );
  FADDX1_HVT DP_OP_423J2_125_3477_U821 ( .A(DP_OP_423J2_125_3477_n1329), .B(
        DP_OP_423J2_125_3477_n1327), .CI(DP_OP_423J2_125_3477_n1325), .CO(
        DP_OP_423J2_125_3477_n1276), .S(DP_OP_423J2_125_3477_n1277) );
  FADDX1_HVT DP_OP_423J2_125_3477_U820 ( .A(DP_OP_423J2_125_3477_n1482), .B(
        DP_OP_423J2_125_3477_n1480), .CI(DP_OP_423J2_125_3477_n1478), .CO(
        DP_OP_423J2_125_3477_n1274), .S(DP_OP_423J2_125_3477_n1275) );
  FADDX1_HVT DP_OP_423J2_125_3477_U819 ( .A(DP_OP_423J2_125_3477_n1466), .B(
        DP_OP_423J2_125_3477_n1311), .CI(DP_OP_423J2_125_3477_n1309), .CO(
        DP_OP_423J2_125_3477_n1272), .S(DP_OP_423J2_125_3477_n1273) );
  FADDX1_HVT DP_OP_423J2_125_3477_U818 ( .A(DP_OP_423J2_125_3477_n1476), .B(
        DP_OP_423J2_125_3477_n1321), .CI(DP_OP_423J2_125_3477_n1323), .CO(
        DP_OP_423J2_125_3477_n1270), .S(DP_OP_423J2_125_3477_n1271) );
  FADDX1_HVT DP_OP_423J2_125_3477_U817 ( .A(DP_OP_423J2_125_3477_n1474), .B(
        DP_OP_423J2_125_3477_n1317), .CI(DP_OP_423J2_125_3477_n1313), .CO(
        DP_OP_423J2_125_3477_n1268), .S(DP_OP_423J2_125_3477_n1269) );
  FADDX1_HVT DP_OP_423J2_125_3477_U816 ( .A(DP_OP_423J2_125_3477_n1472), .B(
        DP_OP_423J2_125_3477_n1319), .CI(DP_OP_423J2_125_3477_n1315), .CO(
        DP_OP_423J2_125_3477_n1266), .S(DP_OP_423J2_125_3477_n1267) );
  FADDX1_HVT DP_OP_423J2_125_3477_U815 ( .A(DP_OP_423J2_125_3477_n1470), .B(
        DP_OP_423J2_125_3477_n1464), .CI(DP_OP_423J2_125_3477_n1468), .CO(
        DP_OP_423J2_125_3477_n1264), .S(DP_OP_423J2_125_3477_n1265) );
  FADDX1_HVT DP_OP_423J2_125_3477_U814 ( .A(DP_OP_423J2_125_3477_n1305), .B(
        DP_OP_423J2_125_3477_n1307), .CI(DP_OP_423J2_125_3477_n1303), .CO(
        DP_OP_423J2_125_3477_n1262), .S(DP_OP_423J2_125_3477_n1263) );
  FADDX1_HVT DP_OP_423J2_125_3477_U813 ( .A(DP_OP_423J2_125_3477_n1295), .B(
        DP_OP_423J2_125_3477_n1297), .CI(DP_OP_423J2_125_3477_n1462), .CO(
        DP_OP_423J2_125_3477_n1260), .S(DP_OP_423J2_125_3477_n1261) );
  FADDX1_HVT DP_OP_423J2_125_3477_U812 ( .A(DP_OP_423J2_125_3477_n1293), .B(
        DP_OP_423J2_125_3477_n1301), .CI(DP_OP_423J2_125_3477_n1299), .CO(
        DP_OP_423J2_125_3477_n1258), .S(DP_OP_423J2_125_3477_n1259) );
  FADDX1_HVT DP_OP_423J2_125_3477_U810 ( .A(DP_OP_423J2_125_3477_n1287), .B(
        DP_OP_423J2_125_3477_n1460), .CI(DP_OP_423J2_125_3477_n1456), .CO(
        DP_OP_423J2_125_3477_n1254), .S(DP_OP_423J2_125_3477_n1255) );
  FADDX1_HVT DP_OP_423J2_125_3477_U809 ( .A(DP_OP_423J2_125_3477_n1285), .B(
        DP_OP_423J2_125_3477_n1452), .CI(DP_OP_423J2_125_3477_n1454), .CO(
        DP_OP_423J2_125_3477_n1252), .S(DP_OP_423J2_125_3477_n1253) );
  FADDX1_HVT DP_OP_423J2_125_3477_U808 ( .A(DP_OP_423J2_125_3477_n1450), .B(
        DP_OP_423J2_125_3477_n1442), .CI(DP_OP_423J2_125_3477_n1279), .CO(
        DP_OP_423J2_125_3477_n1250), .S(DP_OP_423J2_125_3477_n1251) );
  FADDX1_HVT DP_OP_423J2_125_3477_U807 ( .A(DP_OP_423J2_125_3477_n1448), .B(
        DP_OP_423J2_125_3477_n1281), .CI(DP_OP_423J2_125_3477_n1283), .CO(
        DP_OP_423J2_125_3477_n1248), .S(DP_OP_423J2_125_3477_n1249) );
  FADDX1_HVT DP_OP_423J2_125_3477_U806 ( .A(DP_OP_423J2_125_3477_n1446), .B(
        DP_OP_423J2_125_3477_n1444), .CI(DP_OP_423J2_125_3477_n1440), .CO(
        DP_OP_423J2_125_3477_n1246), .S(DP_OP_423J2_125_3477_n1247) );
  FADDX1_HVT DP_OP_423J2_125_3477_U805 ( .A(DP_OP_423J2_125_3477_n1275), .B(
        DP_OP_423J2_125_3477_n1277), .CI(DP_OP_423J2_125_3477_n1438), .CO(
        DP_OP_423J2_125_3477_n1244), .S(DP_OP_423J2_125_3477_n1245) );
  FADDX1_HVT DP_OP_423J2_125_3477_U804 ( .A(DP_OP_423J2_125_3477_n1436), .B(
        DP_OP_423J2_125_3477_n1269), .CI(DP_OP_423J2_125_3477_n1434), .CO(
        DP_OP_423J2_125_3477_n1242), .S(DP_OP_423J2_125_3477_n1243) );
  FADDX1_HVT DP_OP_423J2_125_3477_U803 ( .A(DP_OP_423J2_125_3477_n1267), .B(
        DP_OP_423J2_125_3477_n1273), .CI(DP_OP_423J2_125_3477_n1271), .CO(
        DP_OP_423J2_125_3477_n1240), .S(DP_OP_423J2_125_3477_n1241) );
  FADDX1_HVT DP_OP_423J2_125_3477_U802 ( .A(DP_OP_423J2_125_3477_n1265), .B(
        DP_OP_423J2_125_3477_n1263), .CI(DP_OP_423J2_125_3477_n1259), .CO(
        DP_OP_423J2_125_3477_n1238), .S(DP_OP_423J2_125_3477_n1239) );
  FADDX1_HVT DP_OP_423J2_125_3477_U801 ( .A(DP_OP_423J2_125_3477_n1261), .B(
        DP_OP_423J2_125_3477_n1432), .CI(DP_OP_423J2_125_3477_n1257), .CO(
        DP_OP_423J2_125_3477_n1236), .S(DP_OP_423J2_125_3477_n1237) );
  FADDX1_HVT DP_OP_423J2_125_3477_U800 ( .A(DP_OP_423J2_125_3477_n1430), .B(
        DP_OP_423J2_125_3477_n1428), .CI(DP_OP_423J2_125_3477_n1255), .CO(
        DP_OP_423J2_125_3477_n1234), .S(DP_OP_423J2_125_3477_n1235) );
  FADDX1_HVT DP_OP_423J2_125_3477_U799 ( .A(DP_OP_423J2_125_3477_n1426), .B(
        DP_OP_423J2_125_3477_n1424), .CI(DP_OP_423J2_125_3477_n1253), .CO(
        DP_OP_423J2_125_3477_n1232), .S(DP_OP_423J2_125_3477_n1233) );
  FADDX1_HVT DP_OP_423J2_125_3477_U798 ( .A(DP_OP_423J2_125_3477_n1422), .B(
        DP_OP_423J2_125_3477_n1249), .CI(DP_OP_423J2_125_3477_n1247), .CO(
        DP_OP_423J2_125_3477_n1230), .S(DP_OP_423J2_125_3477_n1231) );
  FADDX1_HVT DP_OP_423J2_125_3477_U797 ( .A(DP_OP_423J2_125_3477_n1420), .B(
        DP_OP_423J2_125_3477_n1251), .CI(DP_OP_423J2_125_3477_n1245), .CO(
        DP_OP_423J2_125_3477_n1228), .S(DP_OP_423J2_125_3477_n1229) );
  FADDX1_HVT DP_OP_423J2_125_3477_U796 ( .A(DP_OP_423J2_125_3477_n1418), .B(
        DP_OP_423J2_125_3477_n1241), .CI(DP_OP_423J2_125_3477_n1416), .CO(
        DP_OP_423J2_125_3477_n1226), .S(DP_OP_423J2_125_3477_n1227) );
  FADDX1_HVT DP_OP_423J2_125_3477_U795 ( .A(DP_OP_423J2_125_3477_n1243), .B(
        DP_OP_423J2_125_3477_n1239), .CI(DP_OP_423J2_125_3477_n1237), .CO(
        DP_OP_423J2_125_3477_n1224), .S(DP_OP_423J2_125_3477_n1225) );
  FADDX1_HVT DP_OP_423J2_125_3477_U793 ( .A(DP_OP_423J2_125_3477_n1410), .B(
        DP_OP_423J2_125_3477_n1233), .CI(DP_OP_423J2_125_3477_n1231), .CO(
        DP_OP_423J2_125_3477_n1220), .S(DP_OP_423J2_125_3477_n1221) );
  FADDX1_HVT DP_OP_423J2_125_3477_U792 ( .A(DP_OP_423J2_125_3477_n1229), .B(
        DP_OP_423J2_125_3477_n1408), .CI(DP_OP_423J2_125_3477_n1227), .CO(
        DP_OP_423J2_125_3477_n1218), .S(DP_OP_423J2_125_3477_n1219) );
  FADDX1_HVT DP_OP_423J2_125_3477_U791 ( .A(DP_OP_423J2_125_3477_n1406), .B(
        DP_OP_423J2_125_3477_n1225), .CI(DP_OP_423J2_125_3477_n1404), .CO(
        DP_OP_423J2_125_3477_n1216), .S(DP_OP_423J2_125_3477_n1217) );
  FADDX1_HVT DP_OP_423J2_125_3477_U790 ( .A(DP_OP_423J2_125_3477_n1223), .B(
        DP_OP_423J2_125_3477_n1221), .CI(DP_OP_423J2_125_3477_n1402), .CO(
        DP_OP_423J2_125_3477_n1214), .S(DP_OP_423J2_125_3477_n1215) );
  FADDX1_HVT DP_OP_423J2_125_3477_U789 ( .A(DP_OP_423J2_125_3477_n1219), .B(
        DP_OP_423J2_125_3477_n1217), .CI(DP_OP_423J2_125_3477_n1400), .CO(
        DP_OP_423J2_125_3477_n1212), .S(DP_OP_423J2_125_3477_n1213) );
  FADDX1_HVT DP_OP_423J2_125_3477_U786 ( .A(DP_OP_423J2_125_3477_n2194), .B(
        DP_OP_423J2_125_3477_n1974), .CI(DP_OP_423J2_125_3477_n1930), .CO(
        DP_OP_423J2_125_3477_n1208), .S(DP_OP_423J2_125_3477_n1209) );
  FADDX1_HVT DP_OP_423J2_125_3477_U785 ( .A(DP_OP_423J2_125_3477_n2634), .B(
        DP_OP_423J2_125_3477_n2062), .CI(DP_OP_423J2_125_3477_n2414), .CO(
        DP_OP_423J2_125_3477_n1206), .S(DP_OP_423J2_125_3477_n1207) );
  FADDX1_HVT DP_OP_423J2_125_3477_U784 ( .A(DP_OP_423J2_125_3477_n2854), .B(
        DP_OP_423J2_125_3477_n2678), .CI(DP_OP_423J2_125_3477_n2238), .CO(
        DP_OP_423J2_125_3477_n1204), .S(DP_OP_423J2_125_3477_n1205) );
  FADDX1_HVT DP_OP_423J2_125_3477_U783 ( .A(DP_OP_423J2_125_3477_n2326), .B(
        DP_OP_423J2_125_3477_n2150), .CI(DP_OP_423J2_125_3477_n2898), .CO(
        DP_OP_423J2_125_3477_n1202), .S(DP_OP_423J2_125_3477_n1203) );
  FADDX1_HVT DP_OP_423J2_125_3477_U782 ( .A(DP_OP_423J2_125_3477_n2458), .B(
        DP_OP_423J2_125_3477_n2942), .CI(DP_OP_423J2_125_3477_n2722), .CO(
        DP_OP_423J2_125_3477_n1200), .S(DP_OP_423J2_125_3477_n1201) );
  FADDX1_HVT DP_OP_423J2_125_3477_U781 ( .A(DP_OP_423J2_125_3477_n2546), .B(
        DP_OP_423J2_125_3477_n2766), .CI(DP_OP_423J2_125_3477_n2590), .CO(
        DP_OP_423J2_125_3477_n1198), .S(DP_OP_423J2_125_3477_n1199) );
  FADDX1_HVT DP_OP_423J2_125_3477_U780 ( .A(DP_OP_423J2_125_3477_n2282), .B(
        DP_OP_423J2_125_3477_n2106), .CI(DP_OP_423J2_125_3477_n2986), .CO(
        DP_OP_423J2_125_3477_n1196), .S(DP_OP_423J2_125_3477_n1197) );
  FADDX1_HVT DP_OP_423J2_125_3477_U779 ( .A(DP_OP_423J2_125_3477_n2810), .B(
        DP_OP_423J2_125_3477_n2018), .CI(DP_OP_423J2_125_3477_n2370), .CO(
        DP_OP_423J2_125_3477_n1194), .S(DP_OP_423J2_125_3477_n1195) );
  FADDX1_HVT DP_OP_423J2_125_3477_U778 ( .A(DP_OP_423J2_125_3477_n2421), .B(
        DP_OP_423J2_125_3477_n3049), .CI(DP_OP_423J2_125_3477_n1981), .CO(
        DP_OP_423J2_125_3477_n1192), .S(DP_OP_423J2_125_3477_n1193) );
  FADDX1_HVT DP_OP_423J2_125_3477_U777 ( .A(DP_OP_423J2_125_3477_n2428), .B(
        DP_OP_423J2_125_3477_n3042), .CI(DP_OP_423J2_125_3477_n3035), .CO(
        DP_OP_423J2_125_3477_n1190), .S(DP_OP_423J2_125_3477_n1191) );
  FADDX1_HVT DP_OP_423J2_125_3477_U776 ( .A(DP_OP_423J2_125_3477_n2384), .B(
        DP_OP_423J2_125_3477_n3007), .CI(DP_OP_423J2_125_3477_n3000), .CO(
        DP_OP_423J2_125_3477_n1188), .S(DP_OP_423J2_125_3477_n1189) );
  FADDX1_HVT DP_OP_423J2_125_3477_U775 ( .A(DP_OP_423J2_125_3477_n2347), .B(
        DP_OP_423J2_125_3477_n2993), .CI(DP_OP_423J2_125_3477_n2963), .CO(
        DP_OP_423J2_125_3477_n1186), .S(DP_OP_423J2_125_3477_n1187) );
  FADDX1_HVT DP_OP_423J2_125_3477_U774 ( .A(DP_OP_423J2_125_3477_n2340), .B(
        DP_OP_423J2_125_3477_n1988), .CI(DP_OP_423J2_125_3477_n2956), .CO(
        DP_OP_423J2_125_3477_n1184), .S(DP_OP_423J2_125_3477_n1185) );
  FADDX1_HVT DP_OP_423J2_125_3477_U773 ( .A(DP_OP_423J2_125_3477_n2377), .B(
        DP_OP_423J2_125_3477_n2949), .CI(DP_OP_423J2_125_3477_n1995), .CO(
        DP_OP_423J2_125_3477_n1182), .S(DP_OP_423J2_125_3477_n1183) );
  FADDX1_HVT DP_OP_423J2_125_3477_U772 ( .A(DP_OP_423J2_125_3477_n2333), .B(
        DP_OP_423J2_125_3477_n2919), .CI(DP_OP_423J2_125_3477_n2025), .CO(
        DP_OP_423J2_125_3477_n1180), .S(DP_OP_423J2_125_3477_n1181) );
  FADDX1_HVT DP_OP_423J2_125_3477_U771 ( .A(DP_OP_423J2_125_3477_n2303), .B(
        DP_OP_423J2_125_3477_n2912), .CI(DP_OP_423J2_125_3477_n2905), .CO(
        DP_OP_423J2_125_3477_n1178), .S(DP_OP_423J2_125_3477_n1179) );
  FADDX1_HVT DP_OP_423J2_125_3477_U770 ( .A(DP_OP_423J2_125_3477_n2296), .B(
        DP_OP_423J2_125_3477_n2032), .CI(DP_OP_423J2_125_3477_n2875), .CO(
        DP_OP_423J2_125_3477_n1176), .S(DP_OP_423J2_125_3477_n1177) );
  FADDX1_HVT DP_OP_423J2_125_3477_U769 ( .A(DP_OP_423J2_125_3477_n2289), .B(
        DP_OP_423J2_125_3477_n2039), .CI(DP_OP_423J2_125_3477_n2868), .CO(
        DP_OP_423J2_125_3477_n1174), .S(DP_OP_423J2_125_3477_n1175) );
  FADDX1_HVT DP_OP_423J2_125_3477_U768 ( .A(DP_OP_423J2_125_3477_n2069), .B(
        DP_OP_423J2_125_3477_n2076), .CI(DP_OP_423J2_125_3477_n2083), .CO(
        DP_OP_423J2_125_3477_n1172), .S(DP_OP_423J2_125_3477_n1173) );
  FADDX1_HVT DP_OP_423J2_125_3477_U767 ( .A(DP_OP_423J2_125_3477_n2861), .B(
        DP_OP_423J2_125_3477_n2113), .CI(DP_OP_423J2_125_3477_n2120), .CO(
        DP_OP_423J2_125_3477_n1170), .S(DP_OP_423J2_125_3477_n1171) );
  FADDX1_HVT DP_OP_423J2_125_3477_U766 ( .A(DP_OP_423J2_125_3477_n2831), .B(
        DP_OP_423J2_125_3477_n2127), .CI(DP_OP_423J2_125_3477_n2157), .CO(
        DP_OP_423J2_125_3477_n1168), .S(DP_OP_423J2_125_3477_n1169) );
  FADDX1_HVT DP_OP_423J2_125_3477_U765 ( .A(DP_OP_423J2_125_3477_n2824), .B(
        DP_OP_423J2_125_3477_n2164), .CI(DP_OP_423J2_125_3477_n2171), .CO(
        DP_OP_423J2_125_3477_n1166), .S(DP_OP_423J2_125_3477_n1167) );
  FADDX1_HVT DP_OP_423J2_125_3477_U764 ( .A(DP_OP_423J2_125_3477_n2817), .B(
        DP_OP_423J2_125_3477_n2201), .CI(DP_OP_423J2_125_3477_n2208), .CO(
        DP_OP_423J2_125_3477_n1164), .S(DP_OP_423J2_125_3477_n1165) );
  FADDX1_HVT DP_OP_423J2_125_3477_U763 ( .A(DP_OP_423J2_125_3477_n2787), .B(
        DP_OP_423J2_125_3477_n2215), .CI(DP_OP_423J2_125_3477_n2245), .CO(
        DP_OP_423J2_125_3477_n1162), .S(DP_OP_423J2_125_3477_n1163) );
  FADDX1_HVT DP_OP_423J2_125_3477_U762 ( .A(DP_OP_423J2_125_3477_n2780), .B(
        DP_OP_423J2_125_3477_n2252), .CI(DP_OP_423J2_125_3477_n2259), .CO(
        DP_OP_423J2_125_3477_n1160), .S(DP_OP_423J2_125_3477_n1161) );
  FADDX1_HVT DP_OP_423J2_125_3477_U761 ( .A(DP_OP_423J2_125_3477_n2773), .B(
        DP_OP_423J2_125_3477_n2391), .CI(DP_OP_423J2_125_3477_n2435), .CO(
        DP_OP_423J2_125_3477_n1158), .S(DP_OP_423J2_125_3477_n1159) );
  FADDX1_HVT DP_OP_423J2_125_3477_U760 ( .A(DP_OP_423J2_125_3477_n2743), .B(
        DP_OP_423J2_125_3477_n2465), .CI(DP_OP_423J2_125_3477_n2472), .CO(
        DP_OP_423J2_125_3477_n1156), .S(DP_OP_423J2_125_3477_n1157) );
  FADDX1_HVT DP_OP_423J2_125_3477_U759 ( .A(DP_OP_423J2_125_3477_n2736), .B(
        DP_OP_423J2_125_3477_n2479), .CI(DP_OP_423J2_125_3477_n2509), .CO(
        DP_OP_423J2_125_3477_n1154), .S(DP_OP_423J2_125_3477_n1155) );
  FADDX1_HVT DP_OP_423J2_125_3477_U758 ( .A(DP_OP_423J2_125_3477_n2729), .B(
        DP_OP_423J2_125_3477_n2516), .CI(DP_OP_423J2_125_3477_n2523), .CO(
        DP_OP_423J2_125_3477_n1152), .S(DP_OP_423J2_125_3477_n1153) );
  FADDX1_HVT DP_OP_423J2_125_3477_U757 ( .A(DP_OP_423J2_125_3477_n2699), .B(
        DP_OP_423J2_125_3477_n2553), .CI(DP_OP_423J2_125_3477_n2560), .CO(
        DP_OP_423J2_125_3477_n1150), .S(DP_OP_423J2_125_3477_n1151) );
  FADDX1_HVT DP_OP_423J2_125_3477_U756 ( .A(DP_OP_423J2_125_3477_n2692), .B(
        DP_OP_423J2_125_3477_n2567), .CI(DP_OP_423J2_125_3477_n2597), .CO(
        DP_OP_423J2_125_3477_n1148), .S(DP_OP_423J2_125_3477_n1149) );
  FADDX1_HVT DP_OP_423J2_125_3477_U755 ( .A(DP_OP_423J2_125_3477_n2685), .B(
        DP_OP_423J2_125_3477_n2604), .CI(DP_OP_423J2_125_3477_n2611), .CO(
        DP_OP_423J2_125_3477_n1146), .S(DP_OP_423J2_125_3477_n1147) );
  FADDX1_HVT DP_OP_423J2_125_3477_U754 ( .A(DP_OP_423J2_125_3477_n2641), .B(
        DP_OP_423J2_125_3477_n2648), .CI(DP_OP_423J2_125_3477_n2655), .CO(
        DP_OP_423J2_125_3477_n1144), .S(DP_OP_423J2_125_3477_n1145) );
  FADDX1_HVT DP_OP_423J2_125_3477_U753 ( .A(DP_OP_423J2_125_3477_n1398), .B(
        DP_OP_423J2_125_3477_n1386), .CI(DP_OP_423J2_125_3477_n1384), .CO(
        DP_OP_423J2_125_3477_n1142), .S(DP_OP_423J2_125_3477_n1143) );
  FADDX1_HVT DP_OP_423J2_125_3477_U752 ( .A(DP_OP_423J2_125_3477_n1382), .B(
        DP_OP_423J2_125_3477_n1388), .CI(DP_OP_423J2_125_3477_n1211), .CO(
        DP_OP_423J2_125_3477_n1140), .S(DP_OP_423J2_125_3477_n1141) );
  FADDX1_HVT DP_OP_423J2_125_3477_U751 ( .A(DP_OP_423J2_125_3477_n1392), .B(
        DP_OP_423J2_125_3477_n1396), .CI(DP_OP_423J2_125_3477_n1390), .CO(
        DP_OP_423J2_125_3477_n1138), .S(DP_OP_423J2_125_3477_n1139) );
  FADDX1_HVT DP_OP_423J2_125_3477_U750 ( .A(DP_OP_423J2_125_3477_n1394), .B(
        DP_OP_423J2_125_3477_n1358), .CI(DP_OP_423J2_125_3477_n1356), .CO(
        DP_OP_423J2_125_3477_n1136), .S(DP_OP_423J2_125_3477_n1137) );
  FADDX1_HVT DP_OP_423J2_125_3477_U749 ( .A(DP_OP_423J2_125_3477_n1360), .B(
        DP_OP_423J2_125_3477_n1332), .CI(DP_OP_423J2_125_3477_n1380), .CO(
        DP_OP_423J2_125_3477_n1134), .S(DP_OP_423J2_125_3477_n1135) );
  FADDX1_HVT DP_OP_423J2_125_3477_U748 ( .A(DP_OP_423J2_125_3477_n1352), .B(
        DP_OP_423J2_125_3477_n1334), .CI(DP_OP_423J2_125_3477_n1378), .CO(
        DP_OP_423J2_125_3477_n1132), .S(DP_OP_423J2_125_3477_n1133) );
  FADDX1_HVT DP_OP_423J2_125_3477_U747 ( .A(DP_OP_423J2_125_3477_n1350), .B(
        DP_OP_423J2_125_3477_n1336), .CI(DP_OP_423J2_125_3477_n1376), .CO(
        DP_OP_423J2_125_3477_n1130), .S(DP_OP_423J2_125_3477_n1131) );
  FADDX1_HVT DP_OP_423J2_125_3477_U746 ( .A(DP_OP_423J2_125_3477_n1346), .B(
        DP_OP_423J2_125_3477_n1374), .CI(DP_OP_423J2_125_3477_n1372), .CO(
        DP_OP_423J2_125_3477_n1128), .S(DP_OP_423J2_125_3477_n1129) );
  FADDX1_HVT DP_OP_423J2_125_3477_U745 ( .A(DP_OP_423J2_125_3477_n1340), .B(
        DP_OP_423J2_125_3477_n1370), .CI(DP_OP_423J2_125_3477_n1368), .CO(
        DP_OP_423J2_125_3477_n1126), .S(DP_OP_423J2_125_3477_n1127) );
  FADDX1_HVT DP_OP_423J2_125_3477_U744 ( .A(DP_OP_423J2_125_3477_n1348), .B(
        DP_OP_423J2_125_3477_n1366), .CI(DP_OP_423J2_125_3477_n1364), .CO(
        DP_OP_423J2_125_3477_n1124), .S(DP_OP_423J2_125_3477_n1125) );
  FADDX1_HVT DP_OP_423J2_125_3477_U743 ( .A(DP_OP_423J2_125_3477_n1342), .B(
        DP_OP_423J2_125_3477_n1362), .CI(DP_OP_423J2_125_3477_n1354), .CO(
        DP_OP_423J2_125_3477_n1122), .S(DP_OP_423J2_125_3477_n1123) );
  FADDX1_HVT DP_OP_423J2_125_3477_U742 ( .A(DP_OP_423J2_125_3477_n1344), .B(
        DP_OP_423J2_125_3477_n1338), .CI(DP_OP_423J2_125_3477_n1201), .CO(
        DP_OP_423J2_125_3477_n1120), .S(DP_OP_423J2_125_3477_n1121) );
  FADDX1_HVT DP_OP_423J2_125_3477_U741 ( .A(DP_OP_423J2_125_3477_n1197), .B(
        DP_OP_423J2_125_3477_n1195), .CI(DP_OP_423J2_125_3477_n1199), .CO(
        DP_OP_423J2_125_3477_n1118), .S(DP_OP_423J2_125_3477_n1119) );
  FADDX1_HVT DP_OP_423J2_125_3477_U740 ( .A(DP_OP_423J2_125_3477_n1207), .B(
        DP_OP_423J2_125_3477_n1205), .CI(DP_OP_423J2_125_3477_n1209), .CO(
        DP_OP_423J2_125_3477_n1116), .S(DP_OP_423J2_125_3477_n1117) );
  FADDX1_HVT DP_OP_423J2_125_3477_U739 ( .A(DP_OP_423J2_125_3477_n1203), .B(
        DP_OP_423J2_125_3477_n1151), .CI(DP_OP_423J2_125_3477_n1153), .CO(
        DP_OP_423J2_125_3477_n1114), .S(DP_OP_423J2_125_3477_n1115) );
  FADDX1_HVT DP_OP_423J2_125_3477_U738 ( .A(DP_OP_423J2_125_3477_n1149), .B(
        DP_OP_423J2_125_3477_n1185), .CI(DP_OP_423J2_125_3477_n1181), .CO(
        DP_OP_423J2_125_3477_n1112), .S(DP_OP_423J2_125_3477_n1113) );
  FADDX1_HVT DP_OP_423J2_125_3477_U737 ( .A(DP_OP_423J2_125_3477_n1187), .B(
        DP_OP_423J2_125_3477_n1171), .CI(DP_OP_423J2_125_3477_n1177), .CO(
        DP_OP_423J2_125_3477_n1110), .S(DP_OP_423J2_125_3477_n1111) );
  FADDX1_HVT DP_OP_423J2_125_3477_U736 ( .A(DP_OP_423J2_125_3477_n1175), .B(
        DP_OP_423J2_125_3477_n1173), .CI(DP_OP_423J2_125_3477_n1157), .CO(
        DP_OP_423J2_125_3477_n1108), .S(DP_OP_423J2_125_3477_n1109) );
  FADDX1_HVT DP_OP_423J2_125_3477_U735 ( .A(DP_OP_423J2_125_3477_n1179), .B(
        DP_OP_423J2_125_3477_n1147), .CI(DP_OP_423J2_125_3477_n1145), .CO(
        DP_OP_423J2_125_3477_n1106), .S(DP_OP_423J2_125_3477_n1107) );
  FADDX1_HVT DP_OP_423J2_125_3477_U734 ( .A(DP_OP_423J2_125_3477_n1183), .B(
        DP_OP_423J2_125_3477_n1165), .CI(DP_OP_423J2_125_3477_n1167), .CO(
        DP_OP_423J2_125_3477_n1104), .S(DP_OP_423J2_125_3477_n1105) );
  FADDX1_HVT DP_OP_423J2_125_3477_U733 ( .A(DP_OP_423J2_125_3477_n1163), .B(
        DP_OP_423J2_125_3477_n1161), .CI(DP_OP_423J2_125_3477_n1155), .CO(
        DP_OP_423J2_125_3477_n1102), .S(DP_OP_423J2_125_3477_n1103) );
  FADDX1_HVT DP_OP_423J2_125_3477_U732 ( .A(DP_OP_423J2_125_3477_n1159), .B(
        DP_OP_423J2_125_3477_n1193), .CI(DP_OP_423J2_125_3477_n1191), .CO(
        DP_OP_423J2_125_3477_n1100), .S(DP_OP_423J2_125_3477_n1101) );
  FADDX1_HVT DP_OP_423J2_125_3477_U731 ( .A(DP_OP_423J2_125_3477_n1189), .B(
        DP_OP_423J2_125_3477_n1169), .CI(DP_OP_423J2_125_3477_n1330), .CO(
        DP_OP_423J2_125_3477_n1098), .S(DP_OP_423J2_125_3477_n1099) );
  FADDX1_HVT DP_OP_423J2_125_3477_U730 ( .A(DP_OP_423J2_125_3477_n1328), .B(
        DP_OP_423J2_125_3477_n1326), .CI(DP_OP_423J2_125_3477_n1324), .CO(
        DP_OP_423J2_125_3477_n1096), .S(DP_OP_423J2_125_3477_n1097) );
  FADDX1_HVT DP_OP_423J2_125_3477_U729 ( .A(DP_OP_423J2_125_3477_n1322), .B(
        DP_OP_423J2_125_3477_n1310), .CI(DP_OP_423J2_125_3477_n1308), .CO(
        DP_OP_423J2_125_3477_n1094), .S(DP_OP_423J2_125_3477_n1095) );
  FADDX1_HVT DP_OP_423J2_125_3477_U728 ( .A(DP_OP_423J2_125_3477_n1314), .B(
        DP_OP_423J2_125_3477_n1312), .CI(DP_OP_423J2_125_3477_n1320), .CO(
        DP_OP_423J2_125_3477_n1092), .S(DP_OP_423J2_125_3477_n1093) );
  FADDX1_HVT DP_OP_423J2_125_3477_U727 ( .A(DP_OP_423J2_125_3477_n1143), .B(
        DP_OP_423J2_125_3477_n1316), .CI(DP_OP_423J2_125_3477_n1318), .CO(
        DP_OP_423J2_125_3477_n1090), .S(DP_OP_423J2_125_3477_n1091) );
  FADDX1_HVT DP_OP_423J2_125_3477_U726 ( .A(DP_OP_423J2_125_3477_n1306), .B(
        DP_OP_423J2_125_3477_n1304), .CI(DP_OP_423J2_125_3477_n1137), .CO(
        DP_OP_423J2_125_3477_n1088), .S(DP_OP_423J2_125_3477_n1089) );
  FADDX1_HVT DP_OP_423J2_125_3477_U725 ( .A(DP_OP_423J2_125_3477_n1141), .B(
        DP_OP_423J2_125_3477_n1139), .CI(DP_OP_423J2_125_3477_n1302), .CO(
        DP_OP_423J2_125_3477_n1086), .S(DP_OP_423J2_125_3477_n1087) );
  FADDX1_HVT DP_OP_423J2_125_3477_U724 ( .A(DP_OP_423J2_125_3477_n1290), .B(
        DP_OP_423J2_125_3477_n1135), .CI(DP_OP_423J2_125_3477_n1121), .CO(
        DP_OP_423J2_125_3477_n1084), .S(DP_OP_423J2_125_3477_n1085) );
  FADDX1_HVT DP_OP_423J2_125_3477_U723 ( .A(DP_OP_423J2_125_3477_n1288), .B(
        DP_OP_423J2_125_3477_n1131), .CI(DP_OP_423J2_125_3477_n1133), .CO(
        DP_OP_423J2_125_3477_n1082), .S(DP_OP_423J2_125_3477_n1083) );
  FADDX1_HVT DP_OP_423J2_125_3477_U722 ( .A(DP_OP_423J2_125_3477_n1292), .B(
        DP_OP_423J2_125_3477_n1129), .CI(DP_OP_423J2_125_3477_n1127), .CO(
        DP_OP_423J2_125_3477_n1080), .S(DP_OP_423J2_125_3477_n1081) );
  FADDX1_HVT DP_OP_423J2_125_3477_U721 ( .A(DP_OP_423J2_125_3477_n1300), .B(
        DP_OP_423J2_125_3477_n1123), .CI(DP_OP_423J2_125_3477_n1125), .CO(
        DP_OP_423J2_125_3477_n1078), .S(DP_OP_423J2_125_3477_n1079) );
  FADDX1_HVT DP_OP_423J2_125_3477_U720 ( .A(DP_OP_423J2_125_3477_n1298), .B(
        DP_OP_423J2_125_3477_n1294), .CI(DP_OP_423J2_125_3477_n1296), .CO(
        DP_OP_423J2_125_3477_n1076), .S(DP_OP_423J2_125_3477_n1077) );
  FADDX1_HVT DP_OP_423J2_125_3477_U719 ( .A(DP_OP_423J2_125_3477_n1117), .B(
        DP_OP_423J2_125_3477_n1286), .CI(DP_OP_423J2_125_3477_n1115), .CO(
        DP_OP_423J2_125_3477_n1074), .S(DP_OP_423J2_125_3477_n1075) );
  FADDX1_HVT DP_OP_423J2_125_3477_U718 ( .A(DP_OP_423J2_125_3477_n1119), .B(
        DP_OP_423J2_125_3477_n1109), .CI(DP_OP_423J2_125_3477_n1111), .CO(
        DP_OP_423J2_125_3477_n1072), .S(DP_OP_423J2_125_3477_n1073) );
  FADDX1_HVT DP_OP_423J2_125_3477_U717 ( .A(DP_OP_423J2_125_3477_n1107), .B(
        DP_OP_423J2_125_3477_n1101), .CI(DP_OP_423J2_125_3477_n1284), .CO(
        DP_OP_423J2_125_3477_n1070), .S(DP_OP_423J2_125_3477_n1071) );
  FADDX1_HVT DP_OP_423J2_125_3477_U716 ( .A(DP_OP_423J2_125_3477_n1103), .B(
        DP_OP_423J2_125_3477_n1113), .CI(DP_OP_423J2_125_3477_n1105), .CO(
        DP_OP_423J2_125_3477_n1068), .S(DP_OP_423J2_125_3477_n1069) );
  FADDX1_HVT DP_OP_423J2_125_3477_U715 ( .A(DP_OP_423J2_125_3477_n1099), .B(
        DP_OP_423J2_125_3477_n1282), .CI(DP_OP_423J2_125_3477_n1278), .CO(
        DP_OP_423J2_125_3477_n1066), .S(DP_OP_423J2_125_3477_n1067) );
  FADDX1_HVT DP_OP_423J2_125_3477_U714 ( .A(DP_OP_423J2_125_3477_n1280), .B(
        DP_OP_423J2_125_3477_n1276), .CI(DP_OP_423J2_125_3477_n1274), .CO(
        DP_OP_423J2_125_3477_n1064), .S(DP_OP_423J2_125_3477_n1065) );
  FADDX1_HVT DP_OP_423J2_125_3477_U713 ( .A(DP_OP_423J2_125_3477_n1097), .B(
        DP_OP_423J2_125_3477_n1272), .CI(DP_OP_423J2_125_3477_n1270), .CO(
        DP_OP_423J2_125_3477_n1062), .S(DP_OP_423J2_125_3477_n1063) );
  FADDX1_HVT DP_OP_423J2_125_3477_U712 ( .A(DP_OP_423J2_125_3477_n1268), .B(
        DP_OP_423J2_125_3477_n1093), .CI(DP_OP_423J2_125_3477_n1091), .CO(
        DP_OP_423J2_125_3477_n1060), .S(DP_OP_423J2_125_3477_n1061) );
  FADDX1_HVT DP_OP_423J2_125_3477_U711 ( .A(DP_OP_423J2_125_3477_n1266), .B(
        DP_OP_423J2_125_3477_n1264), .CI(DP_OP_423J2_125_3477_n1095), .CO(
        DP_OP_423J2_125_3477_n1058), .S(DP_OP_423J2_125_3477_n1059) );
  FADDX1_HVT DP_OP_423J2_125_3477_U710 ( .A(DP_OP_423J2_125_3477_n1087), .B(
        DP_OP_423J2_125_3477_n1262), .CI(DP_OP_423J2_125_3477_n1089), .CO(
        DP_OP_423J2_125_3477_n1056), .S(DP_OP_423J2_125_3477_n1057) );
  FADDX1_HVT DP_OP_423J2_125_3477_U709 ( .A(DP_OP_423J2_125_3477_n1081), .B(
        DP_OP_423J2_125_3477_n1085), .CI(DP_OP_423J2_125_3477_n1256), .CO(
        DP_OP_423J2_125_3477_n1054), .S(DP_OP_423J2_125_3477_n1055) );
  FADDX1_HVT DP_OP_423J2_125_3477_U708 ( .A(DP_OP_423J2_125_3477_n1083), .B(
        DP_OP_423J2_125_3477_n1079), .CI(DP_OP_423J2_125_3477_n1260), .CO(
        DP_OP_423J2_125_3477_n1052), .S(DP_OP_423J2_125_3477_n1053) );
  FADDX1_HVT DP_OP_423J2_125_3477_U707 ( .A(DP_OP_423J2_125_3477_n1258), .B(
        DP_OP_423J2_125_3477_n1077), .CI(DP_OP_423J2_125_3477_n1254), .CO(
        DP_OP_423J2_125_3477_n1050), .S(DP_OP_423J2_125_3477_n1051) );
  FADDX1_HVT DP_OP_423J2_125_3477_U706 ( .A(DP_OP_423J2_125_3477_n1075), .B(
        DP_OP_423J2_125_3477_n1073), .CI(DP_OP_423J2_125_3477_n1071), .CO(
        DP_OP_423J2_125_3477_n1048), .S(DP_OP_423J2_125_3477_n1049) );
  FADDX1_HVT DP_OP_423J2_125_3477_U705 ( .A(DP_OP_423J2_125_3477_n1069), .B(
        DP_OP_423J2_125_3477_n1252), .CI(DP_OP_423J2_125_3477_n1067), .CO(
        DP_OP_423J2_125_3477_n1046), .S(DP_OP_423J2_125_3477_n1047) );
  FADDX1_HVT DP_OP_423J2_125_3477_U703 ( .A(DP_OP_423J2_125_3477_n1065), .B(
        DP_OP_423J2_125_3477_n1244), .CI(DP_OP_423J2_125_3477_n1063), .CO(
        DP_OP_423J2_125_3477_n1042), .S(DP_OP_423J2_125_3477_n1043) );
  FADDX1_HVT DP_OP_423J2_125_3477_U702 ( .A(DP_OP_423J2_125_3477_n1061), .B(
        DP_OP_423J2_125_3477_n1059), .CI(DP_OP_423J2_125_3477_n1242), .CO(
        DP_OP_423J2_125_3477_n1040), .S(DP_OP_423J2_125_3477_n1041) );
  FADDX1_HVT DP_OP_423J2_125_3477_U701 ( .A(DP_OP_423J2_125_3477_n1240), .B(
        DP_OP_423J2_125_3477_n1238), .CI(DP_OP_423J2_125_3477_n1057), .CO(
        DP_OP_423J2_125_3477_n1038), .S(DP_OP_423J2_125_3477_n1039) );
  FADDX1_HVT DP_OP_423J2_125_3477_U700 ( .A(DP_OP_423J2_125_3477_n1236), .B(
        DP_OP_423J2_125_3477_n1051), .CI(DP_OP_423J2_125_3477_n1053), .CO(
        DP_OP_423J2_125_3477_n1036), .S(DP_OP_423J2_125_3477_n1037) );
  FADDX1_HVT DP_OP_423J2_125_3477_U699 ( .A(DP_OP_423J2_125_3477_n1055), .B(
        DP_OP_423J2_125_3477_n1234), .CI(DP_OP_423J2_125_3477_n1049), .CO(
        DP_OP_423J2_125_3477_n1034), .S(DP_OP_423J2_125_3477_n1035) );
  FADDX1_HVT DP_OP_423J2_125_3477_U697 ( .A(DP_OP_423J2_125_3477_n1045), .B(
        DP_OP_423J2_125_3477_n1228), .CI(DP_OP_423J2_125_3477_n1043), .CO(
        DP_OP_423J2_125_3477_n1030), .S(DP_OP_423J2_125_3477_n1031) );
  FADDX1_HVT DP_OP_423J2_125_3477_U696 ( .A(DP_OP_423J2_125_3477_n1226), .B(
        DP_OP_423J2_125_3477_n1041), .CI(DP_OP_423J2_125_3477_n1039), .CO(
        DP_OP_423J2_125_3477_n1028), .S(DP_OP_423J2_125_3477_n1029) );
  FADDX1_HVT DP_OP_423J2_125_3477_U695 ( .A(DP_OP_423J2_125_3477_n1224), .B(
        DP_OP_423J2_125_3477_n1037), .CI(DP_OP_423J2_125_3477_n1222), .CO(
        DP_OP_423J2_125_3477_n1026), .S(DP_OP_423J2_125_3477_n1027) );
  FADDX1_HVT DP_OP_423J2_125_3477_U694 ( .A(DP_OP_423J2_125_3477_n1035), .B(
        DP_OP_423J2_125_3477_n1220), .CI(DP_OP_423J2_125_3477_n1033), .CO(
        DP_OP_423J2_125_3477_n1024), .S(DP_OP_423J2_125_3477_n1025) );
  FADDX1_HVT DP_OP_423J2_125_3477_U693 ( .A(DP_OP_423J2_125_3477_n1031), .B(
        DP_OP_423J2_125_3477_n1218), .CI(DP_OP_423J2_125_3477_n1029), .CO(
        DP_OP_423J2_125_3477_n1022), .S(DP_OP_423J2_125_3477_n1023) );
  FADDX1_HVT DP_OP_423J2_125_3477_U692 ( .A(DP_OP_423J2_125_3477_n1216), .B(
        DP_OP_423J2_125_3477_n1027), .CI(DP_OP_423J2_125_3477_n1025), .CO(
        DP_OP_423J2_125_3477_n1020), .S(DP_OP_423J2_125_3477_n1021) );
  FADDX1_HVT DP_OP_423J2_125_3477_U691 ( .A(DP_OP_423J2_125_3477_n1214), .B(
        DP_OP_423J2_125_3477_n1023), .CI(DP_OP_423J2_125_3477_n1212), .CO(
        DP_OP_423J2_125_3477_n1018), .S(DP_OP_423J2_125_3477_n1019) );
  FADDX1_HVT DP_OP_423J2_125_3477_U690 ( .A(DP_OP_423J2_125_3477_n3028), .B(
        DP_OP_423J2_125_3477_n1973), .CI(DP_OP_423J2_125_3477_n1929), .CO(
        DP_OP_423J2_125_3477_n1016), .S(DP_OP_423J2_125_3477_n1017) );
  FADDX1_HVT DP_OP_423J2_125_3477_U689 ( .A(DP_OP_423J2_125_3477_n2853), .B(
        DP_OP_423J2_125_3477_n2170), .CI(DP_OP_423J2_125_3477_n2434), .CO(
        DP_OP_423J2_125_3477_n1014), .S(DP_OP_423J2_125_3477_n1015) );
  FADDX1_HVT DP_OP_423J2_125_3477_U688 ( .A(DP_OP_423J2_125_3477_n2061), .B(
        DP_OP_423J2_125_3477_n2478), .CI(DP_OP_423J2_125_3477_n2038), .CO(
        DP_OP_423J2_125_3477_n1012), .S(DP_OP_423J2_125_3477_n1013) );
  FADDX1_HVT DP_OP_423J2_125_3477_U687 ( .A(DP_OP_423J2_125_3477_n2369), .B(
        DP_OP_423J2_125_3477_n1994), .CI(DP_OP_423J2_125_3477_n2962), .CO(
        DP_OP_423J2_125_3477_n1010), .S(DP_OP_423J2_125_3477_n1011) );
  FADDX1_HVT DP_OP_423J2_125_3477_U686 ( .A(DP_OP_423J2_125_3477_n2325), .B(
        DP_OP_423J2_125_3477_n2302), .CI(DP_OP_423J2_125_3477_n2654), .CO(
        DP_OP_423J2_125_3477_n1008), .S(DP_OP_423J2_125_3477_n1009) );
  FADDX1_HVT DP_OP_423J2_125_3477_U685 ( .A(DP_OP_423J2_125_3477_n2237), .B(
        DP_OP_423J2_125_3477_n2346), .CI(DP_OP_423J2_125_3477_n3006), .CO(
        DP_OP_423J2_125_3477_n1006), .S(DP_OP_423J2_125_3477_n1007) );
  FADDX1_HVT DP_OP_423J2_125_3477_U684 ( .A(DP_OP_423J2_125_3477_n2017), .B(
        DP_OP_423J2_125_3477_n2082), .CI(DP_OP_423J2_125_3477_n2522), .CO(
        DP_OP_423J2_125_3477_n1004), .S(DP_OP_423J2_125_3477_n1005) );
  FADDX1_HVT DP_OP_423J2_125_3477_U683 ( .A(DP_OP_423J2_125_3477_n2105), .B(
        DP_OP_423J2_125_3477_n2786), .CI(DP_OP_423J2_125_3477_n2830), .CO(
        DP_OP_423J2_125_3477_n1002), .S(DP_OP_423J2_125_3477_n1003) );
  FADDX1_HVT DP_OP_423J2_125_3477_U682 ( .A(DP_OP_423J2_125_3477_n2193), .B(
        DP_OP_423J2_125_3477_n2742), .CI(DP_OP_423J2_125_3477_n2610), .CO(
        DP_OP_423J2_125_3477_n1000), .S(DP_OP_423J2_125_3477_n1001) );
  FADDX1_HVT DP_OP_423J2_125_3477_U681 ( .A(DP_OP_423J2_125_3477_n2545), .B(
        DP_OP_423J2_125_3477_n2390), .CI(DP_OP_423J2_125_3477_n2874), .CO(
        DP_OP_423J2_125_3477_n998), .S(DP_OP_423J2_125_3477_n999) );
  FADDX1_HVT DP_OP_423J2_125_3477_U680 ( .A(DP_OP_423J2_125_3477_n2941), .B(
        DP_OP_423J2_125_3477_n2214), .CI(DP_OP_423J2_125_3477_n2126), .CO(
        DP_OP_423J2_125_3477_n996), .S(DP_OP_423J2_125_3477_n997) );
  FADDX1_HVT DP_OP_423J2_125_3477_U679 ( .A(DP_OP_423J2_125_3477_n2677), .B(
        DP_OP_423J2_125_3477_n2918), .CI(DP_OP_423J2_125_3477_n2566), .CO(
        DP_OP_423J2_125_3477_n994), .S(DP_OP_423J2_125_3477_n995) );
  FADDX1_HVT DP_OP_423J2_125_3477_U678 ( .A(DP_OP_423J2_125_3477_n2457), .B(
        DP_OP_423J2_125_3477_n3048), .CI(DP_OP_423J2_125_3477_n2258), .CO(
        DP_OP_423J2_125_3477_n992), .S(DP_OP_423J2_125_3477_n993) );
  FADDX1_HVT DP_OP_423J2_125_3477_U677 ( .A(DP_OP_423J2_125_3477_n2149), .B(
        DP_OP_423J2_125_3477_n2413), .CI(DP_OP_423J2_125_3477_n2698), .CO(
        DP_OP_423J2_125_3477_n990), .S(DP_OP_423J2_125_3477_n991) );
  FADDX1_HVT DP_OP_423J2_125_3477_U676 ( .A(DP_OP_423J2_125_3477_n2765), .B(
        DP_OP_423J2_125_3477_n2809), .CI(DP_OP_423J2_125_3477_n2897), .CO(
        DP_OP_423J2_125_3477_n988), .S(DP_OP_423J2_125_3477_n989) );
  FADDX1_HVT DP_OP_423J2_125_3477_U675 ( .A(DP_OP_423J2_125_3477_n2501), .B(
        DP_OP_423J2_125_3477_n2589), .CI(DP_OP_423J2_125_3477_n2985), .CO(
        DP_OP_423J2_125_3477_n986), .S(DP_OP_423J2_125_3477_n987) );
  FADDX1_HVT DP_OP_423J2_125_3477_U674 ( .A(DP_OP_423J2_125_3477_n2633), .B(
        DP_OP_423J2_125_3477_n2281), .CI(DP_OP_423J2_125_3477_n2721), .CO(
        DP_OP_423J2_125_3477_n984), .S(DP_OP_423J2_125_3477_n985) );
  FADDX1_HVT DP_OP_423J2_125_3477_U673 ( .A(DP_OP_423J2_125_3477_n3041), .B(
        DP_OP_423J2_125_3477_n1987), .CI(DP_OP_423J2_125_3477_n1980), .CO(
        DP_OP_423J2_125_3477_n982), .S(DP_OP_423J2_125_3477_n983) );
  FADDX1_HVT DP_OP_423J2_125_3477_U672 ( .A(DP_OP_423J2_125_3477_n3034), .B(
        DP_OP_423J2_125_3477_n2999), .CI(DP_OP_423J2_125_3477_n2992), .CO(
        DP_OP_423J2_125_3477_n980), .S(DP_OP_423J2_125_3477_n981) );
  FADDX1_HVT DP_OP_423J2_125_3477_U671 ( .A(DP_OP_423J2_125_3477_n2515), .B(
        DP_OP_423J2_125_3477_n2955), .CI(DP_OP_423J2_125_3477_n2948), .CO(
        DP_OP_423J2_125_3477_n978), .S(DP_OP_423J2_125_3477_n979) );
  FADDX1_HVT DP_OP_423J2_125_3477_U670 ( .A(DP_OP_423J2_125_3477_n2911), .B(
        DP_OP_423J2_125_3477_n2024), .CI(DP_OP_423J2_125_3477_n2031), .CO(
        DP_OP_423J2_125_3477_n976), .S(DP_OP_423J2_125_3477_n977) );
  FADDX1_HVT DP_OP_423J2_125_3477_U669 ( .A(DP_OP_423J2_125_3477_n2904), .B(
        DP_OP_423J2_125_3477_n2068), .CI(DP_OP_423J2_125_3477_n2075), .CO(
        DP_OP_423J2_125_3477_n974), .S(DP_OP_423J2_125_3477_n975) );
  FADDX1_HVT DP_OP_423J2_125_3477_U668 ( .A(DP_OP_423J2_125_3477_n2867), .B(
        DP_OP_423J2_125_3477_n2112), .CI(DP_OP_423J2_125_3477_n2119), .CO(
        DP_OP_423J2_125_3477_n972), .S(DP_OP_423J2_125_3477_n973) );
  FADDX1_HVT DP_OP_423J2_125_3477_U667 ( .A(DP_OP_423J2_125_3477_n2860), .B(
        DP_OP_423J2_125_3477_n2156), .CI(DP_OP_423J2_125_3477_n2163), .CO(
        DP_OP_423J2_125_3477_n970), .S(DP_OP_423J2_125_3477_n971) );
  FADDX1_HVT DP_OP_423J2_125_3477_U666 ( .A(DP_OP_423J2_125_3477_n2823), .B(
        DP_OP_423J2_125_3477_n2200), .CI(DP_OP_423J2_125_3477_n2207), .CO(
        DP_OP_423J2_125_3477_n968), .S(DP_OP_423J2_125_3477_n969) );
  FADDX1_HVT DP_OP_423J2_125_3477_U664 ( .A(DP_OP_423J2_125_3477_n2779), .B(
        DP_OP_423J2_125_3477_n2288), .CI(DP_OP_423J2_125_3477_n2295), .CO(
        DP_OP_423J2_125_3477_n964), .S(DP_OP_423J2_125_3477_n965) );
  FADDX1_HVT DP_OP_423J2_125_3477_U663 ( .A(DP_OP_423J2_125_3477_n2772), .B(
        DP_OP_423J2_125_3477_n2332), .CI(DP_OP_423J2_125_3477_n2339), .CO(
        DP_OP_423J2_125_3477_n962), .S(DP_OP_423J2_125_3477_n963) );
  FADDX1_HVT DP_OP_423J2_125_3477_U662 ( .A(DP_OP_423J2_125_3477_n2735), .B(
        DP_OP_423J2_125_3477_n2376), .CI(DP_OP_423J2_125_3477_n2383), .CO(
        DP_OP_423J2_125_3477_n960), .S(DP_OP_423J2_125_3477_n961) );
  FADDX1_HVT DP_OP_423J2_125_3477_U661 ( .A(DP_OP_423J2_125_3477_n2728), .B(
        DP_OP_423J2_125_3477_n2420), .CI(DP_OP_423J2_125_3477_n2427), .CO(
        DP_OP_423J2_125_3477_n958), .S(DP_OP_423J2_125_3477_n959) );
  FADDX1_HVT DP_OP_423J2_125_3477_U660 ( .A(DP_OP_423J2_125_3477_n2691), .B(
        DP_OP_423J2_125_3477_n2464), .CI(DP_OP_423J2_125_3477_n2471), .CO(
        DP_OP_423J2_125_3477_n956), .S(DP_OP_423J2_125_3477_n957) );
  FADDX1_HVT DP_OP_423J2_125_3477_U659 ( .A(DP_OP_423J2_125_3477_n2684), .B(
        DP_OP_423J2_125_3477_n2508), .CI(DP_OP_423J2_125_3477_n2552), .CO(
        DP_OP_423J2_125_3477_n954), .S(DP_OP_423J2_125_3477_n955) );
  FADDX1_HVT DP_OP_423J2_125_3477_U658 ( .A(DP_OP_423J2_125_3477_n2647), .B(
        DP_OP_423J2_125_3477_n2559), .CI(DP_OP_423J2_125_3477_n2596), .CO(
        DP_OP_423J2_125_3477_n952), .S(DP_OP_423J2_125_3477_n953) );
  FADDX1_HVT DP_OP_423J2_125_3477_U657 ( .A(DP_OP_423J2_125_3477_n2640), .B(
        DP_OP_423J2_125_3477_n2603), .CI(DP_OP_423J2_125_3477_n1210), .CO(
        DP_OP_423J2_125_3477_n950), .S(DP_OP_423J2_125_3477_n951) );
  FADDX1_HVT DP_OP_423J2_125_3477_U656 ( .A(DP_OP_423J2_125_3477_n1198), .B(
        DP_OP_423J2_125_3477_n1194), .CI(DP_OP_423J2_125_3477_n1208), .CO(
        DP_OP_423J2_125_3477_n948), .S(DP_OP_423J2_125_3477_n949) );
  FADDX1_HVT DP_OP_423J2_125_3477_U655 ( .A(DP_OP_423J2_125_3477_n1206), .B(
        DP_OP_423J2_125_3477_n1196), .CI(DP_OP_423J2_125_3477_n1204), .CO(
        DP_OP_423J2_125_3477_n946), .S(DP_OP_423J2_125_3477_n947) );
  FADDX1_HVT DP_OP_423J2_125_3477_U654 ( .A(DP_OP_423J2_125_3477_n1202), .B(
        DP_OP_423J2_125_3477_n1200), .CI(DP_OP_423J2_125_3477_n1170), .CO(
        DP_OP_423J2_125_3477_n944), .S(DP_OP_423J2_125_3477_n945) );
  FADDX1_HVT DP_OP_423J2_125_3477_U653 ( .A(DP_OP_423J2_125_3477_n1168), .B(
        DP_OP_423J2_125_3477_n1144), .CI(DP_OP_423J2_125_3477_n1192), .CO(
        DP_OP_423J2_125_3477_n942), .S(DP_OP_423J2_125_3477_n943) );
  FADDX1_HVT DP_OP_423J2_125_3477_U652 ( .A(DP_OP_423J2_125_3477_n1166), .B(
        DP_OP_423J2_125_3477_n1190), .CI(DP_OP_423J2_125_3477_n1188), .CO(
        DP_OP_423J2_125_3477_n940), .S(DP_OP_423J2_125_3477_n941) );
  FADDX1_HVT DP_OP_423J2_125_3477_U651 ( .A(DP_OP_423J2_125_3477_n1160), .B(
        DP_OP_423J2_125_3477_n1186), .CI(DP_OP_423J2_125_3477_n1184), .CO(
        DP_OP_423J2_125_3477_n938), .S(DP_OP_423J2_125_3477_n939) );
  FADDX1_HVT DP_OP_423J2_125_3477_U650 ( .A(DP_OP_423J2_125_3477_n1182), .B(
        DP_OP_423J2_125_3477_n1180), .CI(DP_OP_423J2_125_3477_n1178), .CO(
        DP_OP_423J2_125_3477_n936), .S(DP_OP_423J2_125_3477_n937) );
  FADDX1_HVT DP_OP_423J2_125_3477_U649 ( .A(DP_OP_423J2_125_3477_n1150), .B(
        DP_OP_423J2_125_3477_n1176), .CI(DP_OP_423J2_125_3477_n1174), .CO(
        DP_OP_423J2_125_3477_n934), .S(DP_OP_423J2_125_3477_n935) );
  FADDX1_HVT DP_OP_423J2_125_3477_U648 ( .A(DP_OP_423J2_125_3477_n1156), .B(
        DP_OP_423J2_125_3477_n1172), .CI(DP_OP_423J2_125_3477_n1164), .CO(
        DP_OP_423J2_125_3477_n932), .S(DP_OP_423J2_125_3477_n933) );
  FADDX1_HVT DP_OP_423J2_125_3477_U647 ( .A(DP_OP_423J2_125_3477_n1148), .B(
        DP_OP_423J2_125_3477_n1162), .CI(DP_OP_423J2_125_3477_n1158), .CO(
        DP_OP_423J2_125_3477_n930), .S(DP_OP_423J2_125_3477_n931) );
  FADDX1_HVT DP_OP_423J2_125_3477_U646 ( .A(DP_OP_423J2_125_3477_n1152), .B(
        DP_OP_423J2_125_3477_n1146), .CI(DP_OP_423J2_125_3477_n1154), .CO(
        DP_OP_423J2_125_3477_n928), .S(DP_OP_423J2_125_3477_n929) );
  FADDX1_HVT DP_OP_423J2_125_3477_U645 ( .A(DP_OP_423J2_125_3477_n1017), .B(
        DP_OP_423J2_125_3477_n1003), .CI(DP_OP_423J2_125_3477_n1005), .CO(
        DP_OP_423J2_125_3477_n926), .S(DP_OP_423J2_125_3477_n927) );
  FADDX1_HVT DP_OP_423J2_125_3477_U644 ( .A(DP_OP_423J2_125_3477_n1009), .B(
        DP_OP_423J2_125_3477_n987), .CI(DP_OP_423J2_125_3477_n985), .CO(
        DP_OP_423J2_125_3477_n924), .S(DP_OP_423J2_125_3477_n925) );
  FADDX1_HVT DP_OP_423J2_125_3477_U643 ( .A(DP_OP_423J2_125_3477_n1001), .B(
        DP_OP_423J2_125_3477_n999), .CI(DP_OP_423J2_125_3477_n995), .CO(
        DP_OP_423J2_125_3477_n922), .S(DP_OP_423J2_125_3477_n923) );
  FADDX1_HVT DP_OP_423J2_125_3477_U642 ( .A(DP_OP_423J2_125_3477_n1007), .B(
        DP_OP_423J2_125_3477_n989), .CI(DP_OP_423J2_125_3477_n993), .CO(
        DP_OP_423J2_125_3477_n920), .S(DP_OP_423J2_125_3477_n921) );
  FADDX1_HVT DP_OP_423J2_125_3477_U641 ( .A(DP_OP_423J2_125_3477_n997), .B(
        DP_OP_423J2_125_3477_n1015), .CI(DP_OP_423J2_125_3477_n1011), .CO(
        DP_OP_423J2_125_3477_n918), .S(DP_OP_423J2_125_3477_n919) );
  FADDX1_HVT DP_OP_423J2_125_3477_U640 ( .A(DP_OP_423J2_125_3477_n991), .B(
        DP_OP_423J2_125_3477_n1013), .CI(DP_OP_423J2_125_3477_n973), .CO(
        DP_OP_423J2_125_3477_n916), .S(DP_OP_423J2_125_3477_n917) );
  FADDX1_HVT DP_OP_423J2_125_3477_U639 ( .A(DP_OP_423J2_125_3477_n975), .B(
        DP_OP_423J2_125_3477_n957), .CI(DP_OP_423J2_125_3477_n951), .CO(
        DP_OP_423J2_125_3477_n914), .S(DP_OP_423J2_125_3477_n915) );
  FADDX1_HVT DP_OP_423J2_125_3477_U637 ( .A(DP_OP_423J2_125_3477_n967), .B(
        DP_OP_423J2_125_3477_n965), .CI(DP_OP_423J2_125_3477_n955), .CO(
        DP_OP_423J2_125_3477_n910), .S(DP_OP_423J2_125_3477_n911) );
  FADDX1_HVT DP_OP_423J2_125_3477_U636 ( .A(DP_OP_423J2_125_3477_n971), .B(
        DP_OP_423J2_125_3477_n959), .CI(DP_OP_423J2_125_3477_n961), .CO(
        DP_OP_423J2_125_3477_n908), .S(DP_OP_423J2_125_3477_n909) );
  FADDX1_HVT DP_OP_423J2_125_3477_U634 ( .A(DP_OP_423J2_125_3477_n963), .B(
        DP_OP_423J2_125_3477_n1142), .CI(DP_OP_423J2_125_3477_n1140), .CO(
        DP_OP_423J2_125_3477_n904), .S(DP_OP_423J2_125_3477_n905) );
  FADDX1_HVT DP_OP_423J2_125_3477_U633 ( .A(DP_OP_423J2_125_3477_n1138), .B(
        DP_OP_423J2_125_3477_n1136), .CI(DP_OP_423J2_125_3477_n1122), .CO(
        DP_OP_423J2_125_3477_n902), .S(DP_OP_423J2_125_3477_n903) );
  FADDX1_HVT DP_OP_423J2_125_3477_U632 ( .A(DP_OP_423J2_125_3477_n1134), .B(
        DP_OP_423J2_125_3477_n1132), .CI(DP_OP_423J2_125_3477_n1120), .CO(
        DP_OP_423J2_125_3477_n900), .S(DP_OP_423J2_125_3477_n901) );
  FADDX1_HVT DP_OP_423J2_125_3477_U631 ( .A(DP_OP_423J2_125_3477_n1130), .B(
        DP_OP_423J2_125_3477_n1124), .CI(DP_OP_423J2_125_3477_n1126), .CO(
        DP_OP_423J2_125_3477_n898), .S(DP_OP_423J2_125_3477_n899) );
  FADDX1_HVT DP_OP_423J2_125_3477_U630 ( .A(DP_OP_423J2_125_3477_n1128), .B(
        DP_OP_423J2_125_3477_n1118), .CI(DP_OP_423J2_125_3477_n1116), .CO(
        DP_OP_423J2_125_3477_n896), .S(DP_OP_423J2_125_3477_n897) );
  FADDX1_HVT DP_OP_423J2_125_3477_U629 ( .A(DP_OP_423J2_125_3477_n949), .B(
        DP_OP_423J2_125_3477_n945), .CI(DP_OP_423J2_125_3477_n1114), .CO(
        DP_OP_423J2_125_3477_n894), .S(DP_OP_423J2_125_3477_n895) );
  FADDX1_HVT DP_OP_423J2_125_3477_U628 ( .A(DP_OP_423J2_125_3477_n947), .B(
        DP_OP_423J2_125_3477_n1102), .CI(DP_OP_423J2_125_3477_n1100), .CO(
        DP_OP_423J2_125_3477_n892), .S(DP_OP_423J2_125_3477_n893) );
  FADDX1_HVT DP_OP_423J2_125_3477_U627 ( .A(DP_OP_423J2_125_3477_n1108), .B(
        DP_OP_423J2_125_3477_n943), .CI(DP_OP_423J2_125_3477_n1098), .CO(
        DP_OP_423J2_125_3477_n890), .S(DP_OP_423J2_125_3477_n891) );
  FADDX1_HVT DP_OP_423J2_125_3477_U626 ( .A(DP_OP_423J2_125_3477_n1106), .B(
        DP_OP_423J2_125_3477_n939), .CI(DP_OP_423J2_125_3477_n929), .CO(
        DP_OP_423J2_125_3477_n888), .S(DP_OP_423J2_125_3477_n889) );
  FADDX1_HVT DP_OP_423J2_125_3477_U625 ( .A(DP_OP_423J2_125_3477_n1112), .B(
        DP_OP_423J2_125_3477_n935), .CI(DP_OP_423J2_125_3477_n937), .CO(
        DP_OP_423J2_125_3477_n886), .S(DP_OP_423J2_125_3477_n887) );
  FADDX1_HVT DP_OP_423J2_125_3477_U624 ( .A(DP_OP_423J2_125_3477_n1110), .B(
        DP_OP_423J2_125_3477_n931), .CI(DP_OP_423J2_125_3477_n933), .CO(
        DP_OP_423J2_125_3477_n884), .S(DP_OP_423J2_125_3477_n885) );
  FADDX1_HVT DP_OP_423J2_125_3477_U623 ( .A(DP_OP_423J2_125_3477_n1104), .B(
        DP_OP_423J2_125_3477_n941), .CI(DP_OP_423J2_125_3477_n927), .CO(
        DP_OP_423J2_125_3477_n882), .S(DP_OP_423J2_125_3477_n883) );
  FADDX1_HVT DP_OP_423J2_125_3477_U622 ( .A(DP_OP_423J2_125_3477_n921), .B(
        DP_OP_423J2_125_3477_n925), .CI(DP_OP_423J2_125_3477_n917), .CO(
        DP_OP_423J2_125_3477_n880), .S(DP_OP_423J2_125_3477_n881) );
  FADDX1_HVT DP_OP_423J2_125_3477_U621 ( .A(DP_OP_423J2_125_3477_n919), .B(
        DP_OP_423J2_125_3477_n923), .CI(DP_OP_423J2_125_3477_n911), .CO(
        DP_OP_423J2_125_3477_n878), .S(DP_OP_423J2_125_3477_n879) );
  FADDX1_HVT DP_OP_423J2_125_3477_U620 ( .A(DP_OP_423J2_125_3477_n909), .B(
        DP_OP_423J2_125_3477_n915), .CI(DP_OP_423J2_125_3477_n1096), .CO(
        DP_OP_423J2_125_3477_n876), .S(DP_OP_423J2_125_3477_n877) );
  FADDX1_HVT DP_OP_423J2_125_3477_U619 ( .A(DP_OP_423J2_125_3477_n913), .B(
        DP_OP_423J2_125_3477_n907), .CI(DP_OP_423J2_125_3477_n1092), .CO(
        DP_OP_423J2_125_3477_n874), .S(DP_OP_423J2_125_3477_n875) );
  FADDX1_HVT DP_OP_423J2_125_3477_U618 ( .A(DP_OP_423J2_125_3477_n905), .B(
        DP_OP_423J2_125_3477_n1090), .CI(DP_OP_423J2_125_3477_n1094), .CO(
        DP_OP_423J2_125_3477_n872), .S(DP_OP_423J2_125_3477_n873) );
  FADDX1_HVT DP_OP_423J2_125_3477_U617 ( .A(DP_OP_423J2_125_3477_n1086), .B(
        DP_OP_423J2_125_3477_n1088), .CI(DP_OP_423J2_125_3477_n903), .CO(
        DP_OP_423J2_125_3477_n870), .S(DP_OP_423J2_125_3477_n871) );
  FADDX1_HVT DP_OP_423J2_125_3477_U616 ( .A(DP_OP_423J2_125_3477_n1084), .B(
        DP_OP_423J2_125_3477_n901), .CI(DP_OP_423J2_125_3477_n899), .CO(
        DP_OP_423J2_125_3477_n868), .S(DP_OP_423J2_125_3477_n869) );
  FADDX1_HVT DP_OP_423J2_125_3477_U615 ( .A(DP_OP_423J2_125_3477_n1082), .B(
        DP_OP_423J2_125_3477_n1076), .CI(DP_OP_423J2_125_3477_n1078), .CO(
        DP_OP_423J2_125_3477_n866), .S(DP_OP_423J2_125_3477_n867) );
  FADDX1_HVT DP_OP_423J2_125_3477_U614 ( .A(DP_OP_423J2_125_3477_n1080), .B(
        DP_OP_423J2_125_3477_n897), .CI(DP_OP_423J2_125_3477_n1074), .CO(
        DP_OP_423J2_125_3477_n864), .S(DP_OP_423J2_125_3477_n865) );
  FADDX1_HVT DP_OP_423J2_125_3477_U613 ( .A(DP_OP_423J2_125_3477_n893), .B(
        DP_OP_423J2_125_3477_n1072), .CI(DP_OP_423J2_125_3477_n895), .CO(
        DP_OP_423J2_125_3477_n862), .S(DP_OP_423J2_125_3477_n863) );
  FADDX1_HVT DP_OP_423J2_125_3477_U612 ( .A(DP_OP_423J2_125_3477_n1070), .B(
        DP_OP_423J2_125_3477_n887), .CI(DP_OP_423J2_125_3477_n883), .CO(
        DP_OP_423J2_125_3477_n860), .S(DP_OP_423J2_125_3477_n861) );
  FADDX1_HVT DP_OP_423J2_125_3477_U611 ( .A(DP_OP_423J2_125_3477_n1068), .B(
        DP_OP_423J2_125_3477_n891), .CI(DP_OP_423J2_125_3477_n889), .CO(
        DP_OP_423J2_125_3477_n858), .S(DP_OP_423J2_125_3477_n859) );
  FADDX1_HVT DP_OP_423J2_125_3477_U610 ( .A(DP_OP_423J2_125_3477_n885), .B(
        DP_OP_423J2_125_3477_n1066), .CI(DP_OP_423J2_125_3477_n881), .CO(
        DP_OP_423J2_125_3477_n856), .S(DP_OP_423J2_125_3477_n857) );
  FADDX1_HVT DP_OP_423J2_125_3477_U609 ( .A(DP_OP_423J2_125_3477_n879), .B(
        DP_OP_423J2_125_3477_n1064), .CI(DP_OP_423J2_125_3477_n877), .CO(
        DP_OP_423J2_125_3477_n854), .S(DP_OP_423J2_125_3477_n855) );
  FADDX1_HVT DP_OP_423J2_125_3477_U608 ( .A(DP_OP_423J2_125_3477_n1062), .B(
        DP_OP_423J2_125_3477_n875), .CI(DP_OP_423J2_125_3477_n1058), .CO(
        DP_OP_423J2_125_3477_n852), .S(DP_OP_423J2_125_3477_n853) );
  FADDX1_HVT DP_OP_423J2_125_3477_U607 ( .A(DP_OP_423J2_125_3477_n1060), .B(
        DP_OP_423J2_125_3477_n873), .CI(DP_OP_423J2_125_3477_n1056), .CO(
        DP_OP_423J2_125_3477_n850), .S(DP_OP_423J2_125_3477_n851) );
  FADDX1_HVT DP_OP_423J2_125_3477_U606 ( .A(DP_OP_423J2_125_3477_n871), .B(
        DP_OP_423J2_125_3477_n1054), .CI(DP_OP_423J2_125_3477_n1052), .CO(
        DP_OP_423J2_125_3477_n848), .S(DP_OP_423J2_125_3477_n849) );
  FADDX1_HVT DP_OP_423J2_125_3477_U605 ( .A(DP_OP_423J2_125_3477_n869), .B(
        DP_OP_423J2_125_3477_n1050), .CI(DP_OP_423J2_125_3477_n865), .CO(
        DP_OP_423J2_125_3477_n846), .S(DP_OP_423J2_125_3477_n847) );
  FADDX1_HVT DP_OP_423J2_125_3477_U604 ( .A(DP_OP_423J2_125_3477_n867), .B(
        DP_OP_423J2_125_3477_n1048), .CI(DP_OP_423J2_125_3477_n863), .CO(
        DP_OP_423J2_125_3477_n844), .S(DP_OP_423J2_125_3477_n845) );
  FADDX1_HVT DP_OP_423J2_125_3477_U603 ( .A(DP_OP_423J2_125_3477_n861), .B(
        DP_OP_423J2_125_3477_n1046), .CI(DP_OP_423J2_125_3477_n857), .CO(
        DP_OP_423J2_125_3477_n842), .S(DP_OP_423J2_125_3477_n843) );
  FADDX1_HVT DP_OP_423J2_125_3477_U602 ( .A(DP_OP_423J2_125_3477_n859), .B(
        DP_OP_423J2_125_3477_n1044), .CI(DP_OP_423J2_125_3477_n855), .CO(
        DP_OP_423J2_125_3477_n840), .S(DP_OP_423J2_125_3477_n841) );
  FADDX1_HVT DP_OP_423J2_125_3477_U601 ( .A(DP_OP_423J2_125_3477_n1042), .B(
        DP_OP_423J2_125_3477_n853), .CI(DP_OP_423J2_125_3477_n1040), .CO(
        DP_OP_423J2_125_3477_n838), .S(DP_OP_423J2_125_3477_n839) );
  FADDX1_HVT DP_OP_423J2_125_3477_U600 ( .A(DP_OP_423J2_125_3477_n851), .B(
        DP_OP_423J2_125_3477_n1038), .CI(DP_OP_423J2_125_3477_n849), .CO(
        DP_OP_423J2_125_3477_n836), .S(DP_OP_423J2_125_3477_n837) );
  FADDX1_HVT DP_OP_423J2_125_3477_U598 ( .A(DP_OP_423J2_125_3477_n845), .B(
        DP_OP_423J2_125_3477_n843), .CI(DP_OP_423J2_125_3477_n1032), .CO(
        DP_OP_423J2_125_3477_n832), .S(DP_OP_423J2_125_3477_n833) );
  FADDX1_HVT DP_OP_423J2_125_3477_U597 ( .A(DP_OP_423J2_125_3477_n841), .B(
        DP_OP_423J2_125_3477_n1030), .CI(DP_OP_423J2_125_3477_n839), .CO(
        DP_OP_423J2_125_3477_n830), .S(DP_OP_423J2_125_3477_n831) );
  FADDX1_HVT DP_OP_423J2_125_3477_U596 ( .A(DP_OP_423J2_125_3477_n1028), .B(
        DP_OP_423J2_125_3477_n837), .CI(DP_OP_423J2_125_3477_n1026), .CO(
        DP_OP_423J2_125_3477_n828), .S(DP_OP_423J2_125_3477_n829) );
  FADDX1_HVT DP_OP_423J2_125_3477_U595 ( .A(DP_OP_423J2_125_3477_n835), .B(
        DP_OP_423J2_125_3477_n833), .CI(DP_OP_423J2_125_3477_n1024), .CO(
        DP_OP_423J2_125_3477_n826), .S(DP_OP_423J2_125_3477_n827) );
  FADDX1_HVT DP_OP_423J2_125_3477_U594 ( .A(DP_OP_423J2_125_3477_n831), .B(
        DP_OP_423J2_125_3477_n1022), .CI(DP_OP_423J2_125_3477_n829), .CO(
        DP_OP_423J2_125_3477_n824), .S(DP_OP_423J2_125_3477_n825) );
  FADDX1_HVT DP_OP_423J2_125_3477_U591 ( .A(DP_OP_423J2_125_3477_n2236), .B(
        DP_OP_423J2_125_3477_n1972), .CI(DP_OP_423J2_125_3477_n1928), .CO(
        DP_OP_423J2_125_3477_n818), .S(DP_OP_423J2_125_3477_n819) );
  FADDX1_HVT DP_OP_423J2_125_3477_U590 ( .A(DP_OP_423J2_125_3477_n2808), .B(
        DP_OP_423J2_125_3477_n2030), .CI(DP_OP_423J2_125_3477_n2294), .CO(
        DP_OP_423J2_125_3477_n816), .S(DP_OP_423J2_125_3477_n817) );
  FADDX1_HVT DP_OP_423J2_125_3477_U589 ( .A(DP_OP_423J2_125_3477_n2280), .B(
        DP_OP_423J2_125_3477_n3040), .CI(DP_OP_423J2_125_3477_n2690), .CO(
        DP_OP_423J2_125_3477_n814), .S(DP_OP_423J2_125_3477_n815) );
  FADDX1_HVT DP_OP_423J2_125_3477_U588 ( .A(DP_OP_423J2_125_3477_n2500), .B(
        DP_OP_423J2_125_3477_n2074), .CI(DP_OP_423J2_125_3477_n2118), .CO(
        DP_OP_423J2_125_3477_n812), .S(DP_OP_423J2_125_3477_n813) );
  FADDX1_HVT DP_OP_423J2_125_3477_U587 ( .A(DP_OP_423J2_125_3477_n2060), .B(
        DP_OP_423J2_125_3477_n2162), .CI(DP_OP_423J2_125_3477_n2206), .CO(
        DP_OP_423J2_125_3477_n810), .S(DP_OP_423J2_125_3477_n811) );
  FADDX1_HVT DP_OP_423J2_125_3477_U586 ( .A(DP_OP_423J2_125_3477_n2764), .B(
        DP_OP_423J2_125_3477_n2866), .CI(DP_OP_423J2_125_3477_n2910), .CO(
        DP_OP_423J2_125_3477_n808), .S(DP_OP_423J2_125_3477_n809) );
  FADDX1_HVT DP_OP_423J2_125_3477_U585 ( .A(DP_OP_423J2_125_3477_n2104), .B(
        DP_OP_423J2_125_3477_n2822), .CI(DP_OP_423J2_125_3477_n2646), .CO(
        DP_OP_423J2_125_3477_n806), .S(DP_OP_423J2_125_3477_n807) );
  FADDX1_HVT DP_OP_423J2_125_3477_U584 ( .A(DP_OP_423J2_125_3477_n2192), .B(
        DP_OP_423J2_125_3477_n2470), .CI(DP_OP_423J2_125_3477_n2998), .CO(
        DP_OP_423J2_125_3477_n804), .S(DP_OP_423J2_125_3477_n805) );
  FADDX1_HVT DP_OP_423J2_125_3477_U583 ( .A(DP_OP_423J2_125_3477_n2720), .B(
        DP_OP_423J2_125_3477_n2954), .CI(DP_OP_423J2_125_3477_n2514), .CO(
        DP_OP_423J2_125_3477_n802), .S(DP_OP_423J2_125_3477_n803) );
  FADDX1_HVT DP_OP_423J2_125_3477_U582 ( .A(DP_OP_423J2_125_3477_n2676), .B(
        DP_OP_423J2_125_3477_n2426), .CI(DP_OP_423J2_125_3477_n2778), .CO(
        DP_OP_423J2_125_3477_n800), .S(DP_OP_423J2_125_3477_n801) );
  FADDX1_HVT DP_OP_423J2_125_3477_U581 ( .A(DP_OP_423J2_125_3477_n2896), .B(
        DP_OP_423J2_125_3477_n2558), .CI(DP_OP_423J2_125_3477_n2382), .CO(
        DP_OP_423J2_125_3477_n798), .S(DP_OP_423J2_125_3477_n799) );
  FADDX1_HVT DP_OP_423J2_125_3477_U580 ( .A(DP_OP_423J2_125_3477_n2368), .B(
        DP_OP_423J2_125_3477_n2338), .CI(DP_OP_423J2_125_3477_n1986), .CO(
        DP_OP_423J2_125_3477_n796), .S(DP_OP_423J2_125_3477_n797) );
  FADDX1_HVT DP_OP_423J2_125_3477_U579 ( .A(DP_OP_423J2_125_3477_n2588), .B(
        DP_OP_423J2_125_3477_n2250), .CI(DP_OP_423J2_125_3477_n2602), .CO(
        DP_OP_423J2_125_3477_n794), .S(DP_OP_423J2_125_3477_n795) );
  FADDX1_HVT DP_OP_423J2_125_3477_U578 ( .A(DP_OP_423J2_125_3477_n2544), .B(
        DP_OP_423J2_125_3477_n2412), .CI(DP_OP_423J2_125_3477_n2734), .CO(
        DP_OP_423J2_125_3477_n792), .S(DP_OP_423J2_125_3477_n793) );
  FADDX1_HVT DP_OP_423J2_125_3477_U577 ( .A(DP_OP_423J2_125_3477_n2852), .B(
        DP_OP_423J2_125_3477_n2148), .CI(DP_OP_423J2_125_3477_n2324), .CO(
        DP_OP_423J2_125_3477_n790), .S(DP_OP_423J2_125_3477_n791) );
  FADDX1_HVT DP_OP_423J2_125_3477_U576 ( .A(DP_OP_423J2_125_3477_n2016), .B(
        DP_OP_423J2_125_3477_n2632), .CI(DP_OP_423J2_125_3477_n2984), .CO(
        DP_OP_423J2_125_3477_n788), .S(DP_OP_423J2_125_3477_n789) );
  FADDX1_HVT DP_OP_423J2_125_3477_U575 ( .A(DP_OP_423J2_125_3477_n2940), .B(
        DP_OP_423J2_125_3477_n2456), .CI(DP_OP_423J2_125_3477_n821), .CO(
        DP_OP_423J2_125_3477_n786), .S(DP_OP_423J2_125_3477_n787) );
  FADDX1_HVT DP_OP_423J2_125_3477_U574 ( .A(DP_OP_423J2_125_3477_n2287), .B(
        DP_OP_423J2_125_3477_n2023), .CI(DP_OP_423J2_125_3477_n1979), .CO(
        DP_OP_423J2_125_3477_n784), .S(DP_OP_423J2_125_3477_n785) );
  FADDX1_HVT DP_OP_423J2_125_3477_U573 ( .A(DP_OP_423J2_125_3477_n3033), .B(
        DP_OP_423J2_125_3477_n2067), .CI(DP_OP_423J2_125_3477_n2111), .CO(
        DP_OP_423J2_125_3477_n782), .S(DP_OP_423J2_125_3477_n783) );
  FADDX1_HVT DP_OP_423J2_125_3477_U572 ( .A(DP_OP_423J2_125_3477_n2991), .B(
        DP_OP_423J2_125_3477_n2155), .CI(DP_OP_423J2_125_3477_n2199), .CO(
        DP_OP_423J2_125_3477_n780), .S(DP_OP_423J2_125_3477_n781) );
  FADDX1_HVT DP_OP_423J2_125_3477_U571 ( .A(DP_OP_423J2_125_3477_n2947), .B(
        DP_OP_423J2_125_3477_n2243), .CI(DP_OP_423J2_125_3477_n2331), .CO(
        DP_OP_423J2_125_3477_n778), .S(DP_OP_423J2_125_3477_n779) );
  FADDX1_HVT DP_OP_423J2_125_3477_U570 ( .A(DP_OP_423J2_125_3477_n2903), .B(
        DP_OP_423J2_125_3477_n2375), .CI(DP_OP_423J2_125_3477_n2419), .CO(
        DP_OP_423J2_125_3477_n776), .S(DP_OP_423J2_125_3477_n777) );
  FADDX1_HVT DP_OP_423J2_125_3477_U569 ( .A(DP_OP_423J2_125_3477_n2859), .B(
        DP_OP_423J2_125_3477_n2463), .CI(DP_OP_423J2_125_3477_n2507), .CO(
        DP_OP_423J2_125_3477_n774), .S(DP_OP_423J2_125_3477_n775) );
  FADDX1_HVT DP_OP_423J2_125_3477_U568 ( .A(DP_OP_423J2_125_3477_n2815), .B(
        DP_OP_423J2_125_3477_n2551), .CI(DP_OP_423J2_125_3477_n2595), .CO(
        DP_OP_423J2_125_3477_n772), .S(DP_OP_423J2_125_3477_n773) );
  FADDX1_HVT DP_OP_423J2_125_3477_U567 ( .A(DP_OP_423J2_125_3477_n2771), .B(
        DP_OP_423J2_125_3477_n2639), .CI(DP_OP_423J2_125_3477_n2683), .CO(
        DP_OP_423J2_125_3477_n770), .S(DP_OP_423J2_125_3477_n771) );
  FADDX1_HVT DP_OP_423J2_125_3477_U566 ( .A(DP_OP_423J2_125_3477_n2727), .B(
        DP_OP_423J2_125_3477_n1016), .CI(DP_OP_423J2_125_3477_n1014), .CO(
        DP_OP_423J2_125_3477_n768), .S(DP_OP_423J2_125_3477_n769) );
  FADDX1_HVT DP_OP_423J2_125_3477_U565 ( .A(DP_OP_423J2_125_3477_n1012), .B(
        DP_OP_423J2_125_3477_n984), .CI(DP_OP_423J2_125_3477_n986), .CO(
        DP_OP_423J2_125_3477_n766), .S(DP_OP_423J2_125_3477_n767) );
  FADDX1_HVT DP_OP_423J2_125_3477_U564 ( .A(DP_OP_423J2_125_3477_n1010), .B(
        DP_OP_423J2_125_3477_n988), .CI(DP_OP_423J2_125_3477_n990), .CO(
        DP_OP_423J2_125_3477_n764), .S(DP_OP_423J2_125_3477_n765) );
  FADDX1_HVT DP_OP_423J2_125_3477_U563 ( .A(DP_OP_423J2_125_3477_n1008), .B(
        DP_OP_423J2_125_3477_n992), .CI(DP_OP_423J2_125_3477_n994), .CO(
        DP_OP_423J2_125_3477_n762), .S(DP_OP_423J2_125_3477_n763) );
  FADDX1_HVT DP_OP_423J2_125_3477_U562 ( .A(DP_OP_423J2_125_3477_n1000), .B(
        DP_OP_423J2_125_3477_n1006), .CI(DP_OP_423J2_125_3477_n996), .CO(
        DP_OP_423J2_125_3477_n760), .S(DP_OP_423J2_125_3477_n761) );
  FADDX1_HVT DP_OP_423J2_125_3477_U561 ( .A(DP_OP_423J2_125_3477_n998), .B(
        DP_OP_423J2_125_3477_n1002), .CI(DP_OP_423J2_125_3477_n1004), .CO(
        DP_OP_423J2_125_3477_n758), .S(DP_OP_423J2_125_3477_n759) );
  FADDX1_HVT DP_OP_423J2_125_3477_U560 ( .A(DP_OP_423J2_125_3477_n982), .B(
        DP_OP_423J2_125_3477_n980), .CI(DP_OP_423J2_125_3477_n950), .CO(
        DP_OP_423J2_125_3477_n756), .S(DP_OP_423J2_125_3477_n757) );
  FADDX1_HVT DP_OP_423J2_125_3477_U559 ( .A(DP_OP_423J2_125_3477_n964), .B(
        DP_OP_423J2_125_3477_n952), .CI(DP_OP_423J2_125_3477_n954), .CO(
        DP_OP_423J2_125_3477_n754), .S(DP_OP_423J2_125_3477_n755) );
  FADDX1_HVT DP_OP_423J2_125_3477_U558 ( .A(DP_OP_423J2_125_3477_n962), .B(
        DP_OP_423J2_125_3477_n956), .CI(DP_OP_423J2_125_3477_n958), .CO(
        DP_OP_423J2_125_3477_n752), .S(DP_OP_423J2_125_3477_n753) );
  FADDX1_HVT DP_OP_423J2_125_3477_U557 ( .A(DP_OP_423J2_125_3477_n960), .B(
        DP_OP_423J2_125_3477_n978), .CI(DP_OP_423J2_125_3477_n976), .CO(
        DP_OP_423J2_125_3477_n750), .S(DP_OP_423J2_125_3477_n751) );
  FADDX1_HVT DP_OP_423J2_125_3477_U555 ( .A(DP_OP_423J2_125_3477_n974), .B(
        DP_OP_423J2_125_3477_n972), .CI(DP_OP_423J2_125_3477_n813), .CO(
        DP_OP_423J2_125_3477_n746), .S(DP_OP_423J2_125_3477_n747) );
  FADDX1_HVT DP_OP_423J2_125_3477_U554 ( .A(DP_OP_423J2_125_3477_n809), .B(
        DP_OP_423J2_125_3477_n805), .CI(DP_OP_423J2_125_3477_n787), .CO(
        DP_OP_423J2_125_3477_n744), .S(DP_OP_423J2_125_3477_n745) );
  FADDX1_HVT DP_OP_423J2_125_3477_U553 ( .A(DP_OP_423J2_125_3477_n811), .B(
        DP_OP_423J2_125_3477_n793), .CI(DP_OP_423J2_125_3477_n791), .CO(
        DP_OP_423J2_125_3477_n742), .S(DP_OP_423J2_125_3477_n743) );
  FADDX1_HVT DP_OP_423J2_125_3477_U552 ( .A(DP_OP_423J2_125_3477_n803), .B(
        DP_OP_423J2_125_3477_n807), .CI(DP_OP_423J2_125_3477_n799), .CO(
        DP_OP_423J2_125_3477_n740), .S(DP_OP_423J2_125_3477_n741) );
  FADDX1_HVT DP_OP_423J2_125_3477_U551 ( .A(DP_OP_423J2_125_3477_n815), .B(
        DP_OP_423J2_125_3477_n795), .CI(DP_OP_423J2_125_3477_n789), .CO(
        DP_OP_423J2_125_3477_n738), .S(DP_OP_423J2_125_3477_n739) );
  FADDX1_HVT DP_OP_423J2_125_3477_U550 ( .A(DP_OP_423J2_125_3477_n797), .B(
        DP_OP_423J2_125_3477_n819), .CI(DP_OP_423J2_125_3477_n817), .CO(
        DP_OP_423J2_125_3477_n736), .S(DP_OP_423J2_125_3477_n737) );
  FADDX1_HVT DP_OP_423J2_125_3477_U549 ( .A(DP_OP_423J2_125_3477_n801), .B(
        DP_OP_423J2_125_3477_n781), .CI(DP_OP_423J2_125_3477_n777), .CO(
        DP_OP_423J2_125_3477_n734), .S(DP_OP_423J2_125_3477_n735) );
  FADDX1_HVT DP_OP_423J2_125_3477_U548 ( .A(DP_OP_423J2_125_3477_n773), .B(
        DP_OP_423J2_125_3477_n771), .CI(DP_OP_423J2_125_3477_n783), .CO(
        DP_OP_423J2_125_3477_n732), .S(DP_OP_423J2_125_3477_n733) );
  FADDX1_HVT DP_OP_423J2_125_3477_U547 ( .A(DP_OP_423J2_125_3477_n779), .B(
        DP_OP_423J2_125_3477_n775), .CI(DP_OP_423J2_125_3477_n785), .CO(
        DP_OP_423J2_125_3477_n730), .S(DP_OP_423J2_125_3477_n731) );
  FADDX1_HVT DP_OP_423J2_125_3477_U546 ( .A(DP_OP_423J2_125_3477_n948), .B(
        DP_OP_423J2_125_3477_n944), .CI(DP_OP_423J2_125_3477_n946), .CO(
        DP_OP_423J2_125_3477_n728), .S(DP_OP_423J2_125_3477_n729) );
  FADDX1_HVT DP_OP_423J2_125_3477_U545 ( .A(DP_OP_423J2_125_3477_n942), .B(
        DP_OP_423J2_125_3477_n928), .CI(DP_OP_423J2_125_3477_n930), .CO(
        DP_OP_423J2_125_3477_n726), .S(DP_OP_423J2_125_3477_n727) );
  FADDX1_HVT DP_OP_423J2_125_3477_U544 ( .A(DP_OP_423J2_125_3477_n940), .B(
        DP_OP_423J2_125_3477_n932), .CI(DP_OP_423J2_125_3477_n938), .CO(
        DP_OP_423J2_125_3477_n724), .S(DP_OP_423J2_125_3477_n725) );
  FADDX1_HVT DP_OP_423J2_125_3477_U543 ( .A(DP_OP_423J2_125_3477_n936), .B(
        DP_OP_423J2_125_3477_n934), .CI(DP_OP_423J2_125_3477_n769), .CO(
        DP_OP_423J2_125_3477_n722), .S(DP_OP_423J2_125_3477_n723) );
  FADDX1_HVT DP_OP_423J2_125_3477_U542 ( .A(DP_OP_423J2_125_3477_n926), .B(
        DP_OP_423J2_125_3477_n767), .CI(DP_OP_423J2_125_3477_n765), .CO(
        DP_OP_423J2_125_3477_n720), .S(DP_OP_423J2_125_3477_n721) );
  FADDX1_HVT DP_OP_423J2_125_3477_U541 ( .A(DP_OP_423J2_125_3477_n924), .B(
        DP_OP_423J2_125_3477_n761), .CI(DP_OP_423J2_125_3477_n763), .CO(
        DP_OP_423J2_125_3477_n718), .S(DP_OP_423J2_125_3477_n719) );
  FADDX1_HVT DP_OP_423J2_125_3477_U540 ( .A(DP_OP_423J2_125_3477_n922), .B(
        DP_OP_423J2_125_3477_n759), .CI(DP_OP_423J2_125_3477_n916), .CO(
        DP_OP_423J2_125_3477_n716), .S(DP_OP_423J2_125_3477_n717) );
  FADDX1_HVT DP_OP_423J2_125_3477_U539 ( .A(DP_OP_423J2_125_3477_n920), .B(
        DP_OP_423J2_125_3477_n918), .CI(DP_OP_423J2_125_3477_n906), .CO(
        DP_OP_423J2_125_3477_n714), .S(DP_OP_423J2_125_3477_n715) );
  FADDX1_HVT DP_OP_423J2_125_3477_U538 ( .A(DP_OP_423J2_125_3477_n914), .B(
        DP_OP_423J2_125_3477_n757), .CI(DP_OP_423J2_125_3477_n747), .CO(
        DP_OP_423J2_125_3477_n712), .S(DP_OP_423J2_125_3477_n713) );
  FADDX1_HVT DP_OP_423J2_125_3477_U536 ( .A(DP_OP_423J2_125_3477_n910), .B(
        DP_OP_423J2_125_3477_n755), .CI(DP_OP_423J2_125_3477_n751), .CO(
        DP_OP_423J2_125_3477_n708), .S(DP_OP_423J2_125_3477_n709) );
  FADDX1_HVT DP_OP_423J2_125_3477_U535 ( .A(DP_OP_423J2_125_3477_n908), .B(
        DP_OP_423J2_125_3477_n743), .CI(DP_OP_423J2_125_3477_n739), .CO(
        DP_OP_423J2_125_3477_n706), .S(DP_OP_423J2_125_3477_n707) );
  FADDX1_HVT DP_OP_423J2_125_3477_U534 ( .A(DP_OP_423J2_125_3477_n741), .B(
        DP_OP_423J2_125_3477_n904), .CI(DP_OP_423J2_125_3477_n735), .CO(
        DP_OP_423J2_125_3477_n704), .S(DP_OP_423J2_125_3477_n705) );
  FADDX1_HVT DP_OP_423J2_125_3477_U533 ( .A(DP_OP_423J2_125_3477_n737), .B(
        DP_OP_423J2_125_3477_n745), .CI(DP_OP_423J2_125_3477_n731), .CO(
        DP_OP_423J2_125_3477_n702), .S(DP_OP_423J2_125_3477_n703) );
  FADDX1_HVT DP_OP_423J2_125_3477_U532 ( .A(DP_OP_423J2_125_3477_n733), .B(
        DP_OP_423J2_125_3477_n902), .CI(DP_OP_423J2_125_3477_n900), .CO(
        DP_OP_423J2_125_3477_n700), .S(DP_OP_423J2_125_3477_n701) );
  FADDX1_HVT DP_OP_423J2_125_3477_U531 ( .A(DP_OP_423J2_125_3477_n898), .B(
        DP_OP_423J2_125_3477_n896), .CI(DP_OP_423J2_125_3477_n729), .CO(
        DP_OP_423J2_125_3477_n698), .S(DP_OP_423J2_125_3477_n699) );
  FADDX1_HVT DP_OP_423J2_125_3477_U530 ( .A(DP_OP_423J2_125_3477_n894), .B(
        DP_OP_423J2_125_3477_n892), .CI(DP_OP_423J2_125_3477_n890), .CO(
        DP_OP_423J2_125_3477_n696), .S(DP_OP_423J2_125_3477_n697) );
  FADDX1_HVT DP_OP_423J2_125_3477_U529 ( .A(DP_OP_423J2_125_3477_n888), .B(
        DP_OP_423J2_125_3477_n723), .CI(DP_OP_423J2_125_3477_n882), .CO(
        DP_OP_423J2_125_3477_n694), .S(DP_OP_423J2_125_3477_n695) );
  FADDX1_HVT DP_OP_423J2_125_3477_U528 ( .A(DP_OP_423J2_125_3477_n886), .B(
        DP_OP_423J2_125_3477_n725), .CI(DP_OP_423J2_125_3477_n727), .CO(
        DP_OP_423J2_125_3477_n692), .S(DP_OP_423J2_125_3477_n693) );
  FADDX1_HVT DP_OP_423J2_125_3477_U527 ( .A(DP_OP_423J2_125_3477_n884), .B(
        DP_OP_423J2_125_3477_n721), .CI(DP_OP_423J2_125_3477_n717), .CO(
        DP_OP_423J2_125_3477_n690), .S(DP_OP_423J2_125_3477_n691) );
  FADDX1_HVT DP_OP_423J2_125_3477_U526 ( .A(DP_OP_423J2_125_3477_n880), .B(
        DP_OP_423J2_125_3477_n719), .CI(DP_OP_423J2_125_3477_n715), .CO(
        DP_OP_423J2_125_3477_n688), .S(DP_OP_423J2_125_3477_n689) );
  FADDX1_HVT DP_OP_423J2_125_3477_U524 ( .A(DP_OP_423J2_125_3477_n709), .B(
        DP_OP_423J2_125_3477_n713), .CI(DP_OP_423J2_125_3477_n874), .CO(
        DP_OP_423J2_125_3477_n684), .S(DP_OP_423J2_125_3477_n685) );
  FADDX1_HVT DP_OP_423J2_125_3477_U523 ( .A(DP_OP_423J2_125_3477_n707), .B(
        DP_OP_423J2_125_3477_n872), .CI(DP_OP_423J2_125_3477_n703), .CO(
        DP_OP_423J2_125_3477_n682), .S(DP_OP_423J2_125_3477_n683) );
  FADDX1_HVT DP_OP_423J2_125_3477_U522 ( .A(DP_OP_423J2_125_3477_n705), .B(
        DP_OP_423J2_125_3477_n870), .CI(DP_OP_423J2_125_3477_n701), .CO(
        DP_OP_423J2_125_3477_n680), .S(DP_OP_423J2_125_3477_n681) );
  FADDX1_HVT DP_OP_423J2_125_3477_U521 ( .A(DP_OP_423J2_125_3477_n868), .B(
        DP_OP_423J2_125_3477_n866), .CI(DP_OP_423J2_125_3477_n699), .CO(
        DP_OP_423J2_125_3477_n678), .S(DP_OP_423J2_125_3477_n679) );
  FADDX1_HVT DP_OP_423J2_125_3477_U520 ( .A(DP_OP_423J2_125_3477_n864), .B(
        DP_OP_423J2_125_3477_n862), .CI(DP_OP_423J2_125_3477_n697), .CO(
        DP_OP_423J2_125_3477_n676), .S(DP_OP_423J2_125_3477_n677) );
  FADDX1_HVT DP_OP_423J2_125_3477_U519 ( .A(DP_OP_423J2_125_3477_n693), .B(
        DP_OP_423J2_125_3477_n860), .CI(DP_OP_423J2_125_3477_n856), .CO(
        DP_OP_423J2_125_3477_n674), .S(DP_OP_423J2_125_3477_n675) );
  FADDX1_HVT DP_OP_423J2_125_3477_U518 ( .A(DP_OP_423J2_125_3477_n858), .B(
        DP_OP_423J2_125_3477_n695), .CI(DP_OP_423J2_125_3477_n691), .CO(
        DP_OP_423J2_125_3477_n672), .S(DP_OP_423J2_125_3477_n673) );
  FADDX1_HVT DP_OP_423J2_125_3477_U517 ( .A(DP_OP_423J2_125_3477_n689), .B(
        DP_OP_423J2_125_3477_n687), .CI(DP_OP_423J2_125_3477_n854), .CO(
        DP_OP_423J2_125_3477_n670), .S(DP_OP_423J2_125_3477_n671) );
  FADDX1_HVT DP_OP_423J2_125_3477_U516 ( .A(DP_OP_423J2_125_3477_n685), .B(
        DP_OP_423J2_125_3477_n852), .CI(DP_OP_423J2_125_3477_n683), .CO(
        DP_OP_423J2_125_3477_n668), .S(DP_OP_423J2_125_3477_n669) );
  FADDX1_HVT DP_OP_423J2_125_3477_U515 ( .A(DP_OP_423J2_125_3477_n850), .B(
        DP_OP_423J2_125_3477_n681), .CI(DP_OP_423J2_125_3477_n848), .CO(
        DP_OP_423J2_125_3477_n666), .S(DP_OP_423J2_125_3477_n667) );
  FADDX1_HVT DP_OP_423J2_125_3477_U514 ( .A(DP_OP_423J2_125_3477_n846), .B(
        DP_OP_423J2_125_3477_n679), .CI(DP_OP_423J2_125_3477_n844), .CO(
        DP_OP_423J2_125_3477_n664), .S(DP_OP_423J2_125_3477_n665) );
  FADDX1_HVT DP_OP_423J2_125_3477_U513 ( .A(DP_OP_423J2_125_3477_n677), .B(
        DP_OP_423J2_125_3477_n842), .CI(DP_OP_423J2_125_3477_n675), .CO(
        DP_OP_423J2_125_3477_n662), .S(DP_OP_423J2_125_3477_n663) );
  FADDX1_HVT DP_OP_423J2_125_3477_U512 ( .A(DP_OP_423J2_125_3477_n673), .B(
        DP_OP_423J2_125_3477_n840), .CI(DP_OP_423J2_125_3477_n671), .CO(
        DP_OP_423J2_125_3477_n660), .S(DP_OP_423J2_125_3477_n661) );
  FADDX1_HVT DP_OP_423J2_125_3477_U511 ( .A(DP_OP_423J2_125_3477_n838), .B(
        DP_OP_423J2_125_3477_n669), .CI(DP_OP_423J2_125_3477_n836), .CO(
        DP_OP_423J2_125_3477_n658), .S(DP_OP_423J2_125_3477_n659) );
  FADDX1_HVT DP_OP_423J2_125_3477_U510 ( .A(DP_OP_423J2_125_3477_n667), .B(
        DP_OP_423J2_125_3477_n834), .CI(DP_OP_423J2_125_3477_n665), .CO(
        DP_OP_423J2_125_3477_n656), .S(DP_OP_423J2_125_3477_n657) );
  FADDX1_HVT DP_OP_423J2_125_3477_U509 ( .A(DP_OP_423J2_125_3477_n663), .B(
        DP_OP_423J2_125_3477_n832), .CI(DP_OP_423J2_125_3477_n661), .CO(
        DP_OP_423J2_125_3477_n654), .S(DP_OP_423J2_125_3477_n655) );
  FADDX1_HVT DP_OP_423J2_125_3477_U508 ( .A(DP_OP_423J2_125_3477_n830), .B(
        DP_OP_423J2_125_3477_n659), .CI(DP_OP_423J2_125_3477_n828), .CO(
        DP_OP_423J2_125_3477_n652), .S(DP_OP_423J2_125_3477_n653) );
  FADDX1_HVT DP_OP_423J2_125_3477_U507 ( .A(DP_OP_423J2_125_3477_n657), .B(
        DP_OP_423J2_125_3477_n826), .CI(DP_OP_423J2_125_3477_n655), .CO(
        DP_OP_423J2_125_3477_n650), .S(DP_OP_423J2_125_3477_n651) );
  FADDX1_HVT DP_OP_423J2_125_3477_U505 ( .A(DP_OP_423J2_125_3477_n3027), .B(
        DP_OP_423J2_125_3477_n1971), .CI(DP_OP_423J2_125_3477_n1927), .CO(
        DP_OP_423J2_125_3477_n646), .S(DP_OP_423J2_125_3477_n647) );
  FADDX1_HVT DP_OP_423J2_125_3477_U504 ( .A(DP_OP_423J2_125_3477_n820), .B(
        DP_OP_423J2_125_3477_n2286), .CI(DP_OP_423J2_125_3477_n1978), .CO(
        DP_OP_423J2_125_3477_n644), .S(DP_OP_423J2_125_3477_n645) );
  FADDX1_HVT DP_OP_423J2_125_3477_U503 ( .A(DP_OP_423J2_125_3477_n2367), .B(
        DP_OP_423J2_125_3477_n3032), .CI(DP_OP_423J2_125_3477_n2682), .CO(
        DP_OP_423J2_125_3477_n642), .S(DP_OP_423J2_125_3477_n643) );
  FADDX1_HVT DP_OP_423J2_125_3477_U502 ( .A(DP_OP_423J2_125_3477_n2059), .B(
        DP_OP_423J2_125_3477_n2594), .CI(DP_OP_423J2_125_3477_n2814), .CO(
        DP_OP_423J2_125_3477_n640), .S(DP_OP_423J2_125_3477_n641) );
  FADDX1_HVT DP_OP_423J2_125_3477_U501 ( .A(DP_OP_423J2_125_3477_n2279), .B(
        DP_OP_423J2_125_3477_n2374), .CI(DP_OP_423J2_125_3477_n2990), .CO(
        DP_OP_423J2_125_3477_n638), .S(DP_OP_423J2_125_3477_n639) );
  FADDX1_HVT DP_OP_423J2_125_3477_U500 ( .A(DP_OP_423J2_125_3477_n2015), .B(
        DP_OP_423J2_125_3477_n2902), .CI(DP_OP_423J2_125_3477_n2066), .CO(
        DP_OP_423J2_125_3477_n636), .S(DP_OP_423J2_125_3477_n637) );
  FADDX1_HVT DP_OP_423J2_125_3477_U499 ( .A(DP_OP_423J2_125_3477_n2147), .B(
        DP_OP_423J2_125_3477_n2022), .CI(DP_OP_423J2_125_3477_n2858), .CO(
        DP_OP_423J2_125_3477_n634), .S(DP_OP_423J2_125_3477_n635) );
  FADDX1_HVT DP_OP_423J2_125_3477_U498 ( .A(DP_OP_423J2_125_3477_n2983), .B(
        DP_OP_423J2_125_3477_n2418), .CI(DP_OP_423J2_125_3477_n2506), .CO(
        DP_OP_423J2_125_3477_n632), .S(DP_OP_423J2_125_3477_n633) );
  FADDX1_HVT DP_OP_423J2_125_3477_U497 ( .A(DP_OP_423J2_125_3477_n2499), .B(
        DP_OP_423J2_125_3477_n2550), .CI(DP_OP_423J2_125_3477_n2946), .CO(
        DP_OP_423J2_125_3477_n630), .S(DP_OP_423J2_125_3477_n631) );
  FADDX1_HVT DP_OP_423J2_125_3477_U496 ( .A(DP_OP_423J2_125_3477_n2763), .B(
        DP_OP_423J2_125_3477_n2242), .CI(DP_OP_423J2_125_3477_n2770), .CO(
        DP_OP_423J2_125_3477_n628), .S(DP_OP_423J2_125_3477_n629) );
  FADDX1_HVT DP_OP_423J2_125_3477_U495 ( .A(DP_OP_423J2_125_3477_n2939), .B(
        DP_OP_423J2_125_3477_n2462), .CI(DP_OP_423J2_125_3477_n2638), .CO(
        DP_OP_423J2_125_3477_n626), .S(DP_OP_423J2_125_3477_n627) );
  FADDX1_HVT DP_OP_423J2_125_3477_U494 ( .A(DP_OP_423J2_125_3477_n2235), .B(
        DP_OP_423J2_125_3477_n2110), .CI(DP_OP_423J2_125_3477_n2726), .CO(
        DP_OP_423J2_125_3477_n624), .S(DP_OP_423J2_125_3477_n625) );
  FADDX1_HVT DP_OP_423J2_125_3477_U493 ( .A(DP_OP_423J2_125_3477_n2191), .B(
        DP_OP_423J2_125_3477_n2330), .CI(DP_OP_423J2_125_3477_n2198), .CO(
        DP_OP_423J2_125_3477_n622), .S(DP_OP_423J2_125_3477_n623) );
  FADDX1_HVT DP_OP_423J2_125_3477_U492 ( .A(DP_OP_423J2_125_3477_n2587), .B(
        DP_OP_423J2_125_3477_n2411), .CI(DP_OP_423J2_125_3477_n2154), .CO(
        DP_OP_423J2_125_3477_n620), .S(DP_OP_423J2_125_3477_n621) );
  FADDX1_HVT DP_OP_423J2_125_3477_U491 ( .A(DP_OP_423J2_125_3477_n2895), .B(
        DP_OP_423J2_125_3477_n2103), .CI(DP_OP_423J2_125_3477_n2323), .CO(
        DP_OP_423J2_125_3477_n618), .S(DP_OP_423J2_125_3477_n619) );
  FADDX1_HVT DP_OP_423J2_125_3477_U490 ( .A(DP_OP_423J2_125_3477_n2851), .B(
        DP_OP_423J2_125_3477_n2455), .CI(DP_OP_423J2_125_3477_n2543), .CO(
        DP_OP_423J2_125_3477_n616), .S(DP_OP_423J2_125_3477_n617) );
  FADDX1_HVT DP_OP_423J2_125_3477_U489 ( .A(DP_OP_423J2_125_3477_n2807), .B(
        DP_OP_423J2_125_3477_n2631), .CI(DP_OP_423J2_125_3477_n2675), .CO(
        DP_OP_423J2_125_3477_n614), .S(DP_OP_423J2_125_3477_n615) );
  FADDX1_HVT DP_OP_423J2_125_3477_U488 ( .A(DP_OP_423J2_125_3477_n2719), .B(
        DP_OP_423J2_125_3477_n818), .CI(DP_OP_423J2_125_3477_n816), .CO(
        DP_OP_423J2_125_3477_n612), .S(DP_OP_423J2_125_3477_n613) );
  FADDX1_HVT DP_OP_423J2_125_3477_U487 ( .A(DP_OP_423J2_125_3477_n814), .B(
        DP_OP_423J2_125_3477_n786), .CI(DP_OP_423J2_125_3477_n788), .CO(
        DP_OP_423J2_125_3477_n610), .S(DP_OP_423J2_125_3477_n611) );
  FADDX1_HVT DP_OP_423J2_125_3477_U486 ( .A(DP_OP_423J2_125_3477_n812), .B(
        DP_OP_423J2_125_3477_n790), .CI(DP_OP_423J2_125_3477_n792), .CO(
        DP_OP_423J2_125_3477_n608), .S(DP_OP_423J2_125_3477_n609) );
  FADDX1_HVT DP_OP_423J2_125_3477_U485 ( .A(DP_OP_423J2_125_3477_n810), .B(
        DP_OP_423J2_125_3477_n794), .CI(DP_OP_423J2_125_3477_n796), .CO(
        DP_OP_423J2_125_3477_n606), .S(DP_OP_423J2_125_3477_n607) );
  FADDX1_HVT DP_OP_423J2_125_3477_U484 ( .A(DP_OP_423J2_125_3477_n808), .B(
        DP_OP_423J2_125_3477_n798), .CI(DP_OP_423J2_125_3477_n800), .CO(
        DP_OP_423J2_125_3477_n604), .S(DP_OP_423J2_125_3477_n605) );
  FADDX1_HVT DP_OP_423J2_125_3477_U483 ( .A(DP_OP_423J2_125_3477_n806), .B(
        DP_OP_423J2_125_3477_n802), .CI(DP_OP_423J2_125_3477_n804), .CO(
        DP_OP_423J2_125_3477_n602), .S(DP_OP_423J2_125_3477_n603) );
  FADDX1_HVT DP_OP_423J2_125_3477_U482 ( .A(DP_OP_423J2_125_3477_n784), .B(
        DP_OP_423J2_125_3477_n770), .CI(DP_OP_423J2_125_3477_n782), .CO(
        DP_OP_423J2_125_3477_n600), .S(DP_OP_423J2_125_3477_n601) );
  FADDX1_HVT DP_OP_423J2_125_3477_U481 ( .A(DP_OP_423J2_125_3477_n776), .B(
        DP_OP_423J2_125_3477_n772), .CI(DP_OP_423J2_125_3477_n774), .CO(
        DP_OP_423J2_125_3477_n598), .S(DP_OP_423J2_125_3477_n599) );
  FADDX1_HVT DP_OP_423J2_125_3477_U480 ( .A(DP_OP_423J2_125_3477_n780), .B(
        DP_OP_423J2_125_3477_n778), .CI(DP_OP_423J2_125_3477_n645), .CO(
        DP_OP_423J2_125_3477_n596), .S(DP_OP_423J2_125_3477_n597) );
  FADDX1_HVT DP_OP_423J2_125_3477_U479 ( .A(DP_OP_423J2_125_3477_n647), .B(
        DP_OP_423J2_125_3477_n633), .CI(DP_OP_423J2_125_3477_n639), .CO(
        DP_OP_423J2_125_3477_n594), .S(DP_OP_423J2_125_3477_n595) );
  FADDX1_HVT DP_OP_423J2_125_3477_U478 ( .A(DP_OP_423J2_125_3477_n615), .B(
        DP_OP_423J2_125_3477_n637), .CI(DP_OP_423J2_125_3477_n635), .CO(
        DP_OP_423J2_125_3477_n592), .S(DP_OP_423J2_125_3477_n593) );
  FADDX1_HVT DP_OP_423J2_125_3477_U477 ( .A(DP_OP_423J2_125_3477_n641), .B(
        DP_OP_423J2_125_3477_n623), .CI(DP_OP_423J2_125_3477_n625), .CO(
        DP_OP_423J2_125_3477_n590), .S(DP_OP_423J2_125_3477_n591) );
  FADDX1_HVT DP_OP_423J2_125_3477_U476 ( .A(DP_OP_423J2_125_3477_n627), .B(
        DP_OP_423J2_125_3477_n617), .CI(DP_OP_423J2_125_3477_n619), .CO(
        DP_OP_423J2_125_3477_n588), .S(DP_OP_423J2_125_3477_n589) );
  FADDX1_HVT DP_OP_423J2_125_3477_U475 ( .A(DP_OP_423J2_125_3477_n621), .B(
        DP_OP_423J2_125_3477_n643), .CI(DP_OP_423J2_125_3477_n631), .CO(
        DP_OP_423J2_125_3477_n586), .S(DP_OP_423J2_125_3477_n587) );
  FADDX1_HVT DP_OP_423J2_125_3477_U474 ( .A(DP_OP_423J2_125_3477_n629), .B(
        DP_OP_423J2_125_3477_n768), .CI(DP_OP_423J2_125_3477_n766), .CO(
        DP_OP_423J2_125_3477_n584), .S(DP_OP_423J2_125_3477_n585) );
  FADDX1_HVT DP_OP_423J2_125_3477_U473 ( .A(DP_OP_423J2_125_3477_n764), .B(
        DP_OP_423J2_125_3477_n758), .CI(DP_OP_423J2_125_3477_n760), .CO(
        DP_OP_423J2_125_3477_n582), .S(DP_OP_423J2_125_3477_n583) );
  FADDX1_HVT DP_OP_423J2_125_3477_U472 ( .A(DP_OP_423J2_125_3477_n762), .B(
        DP_OP_423J2_125_3477_n756), .CI(DP_OP_423J2_125_3477_n754), .CO(
        DP_OP_423J2_125_3477_n580), .S(DP_OP_423J2_125_3477_n581) );
  FADDX1_HVT DP_OP_423J2_125_3477_U471 ( .A(DP_OP_423J2_125_3477_n752), .B(
        DP_OP_423J2_125_3477_n748), .CI(DP_OP_423J2_125_3477_n746), .CO(
        DP_OP_423J2_125_3477_n578), .S(DP_OP_423J2_125_3477_n579) );
  FADDX1_HVT DP_OP_423J2_125_3477_U470 ( .A(DP_OP_423J2_125_3477_n750), .B(
        DP_OP_423J2_125_3477_n613), .CI(DP_OP_423J2_125_3477_n607), .CO(
        DP_OP_423J2_125_3477_n576), .S(DP_OP_423J2_125_3477_n577) );
  FADDX1_HVT DP_OP_423J2_125_3477_U469 ( .A(DP_OP_423J2_125_3477_n609), .B(
        DP_OP_423J2_125_3477_n603), .CI(DP_OP_423J2_125_3477_n734), .CO(
        DP_OP_423J2_125_3477_n574), .S(DP_OP_423J2_125_3477_n575) );
  FADDX1_HVT DP_OP_423J2_125_3477_U468 ( .A(DP_OP_423J2_125_3477_n744), .B(
        DP_OP_423J2_125_3477_n611), .CI(DP_OP_423J2_125_3477_n605), .CO(
        DP_OP_423J2_125_3477_n572), .S(DP_OP_423J2_125_3477_n573) );
  FADDX1_HVT DP_OP_423J2_125_3477_U467 ( .A(DP_OP_423J2_125_3477_n738), .B(
        DP_OP_423J2_125_3477_n742), .CI(DP_OP_423J2_125_3477_n736), .CO(
        DP_OP_423J2_125_3477_n570), .S(DP_OP_423J2_125_3477_n571) );
  FADDX1_HVT DP_OP_423J2_125_3477_U466 ( .A(DP_OP_423J2_125_3477_n740), .B(
        DP_OP_423J2_125_3477_n732), .CI(DP_OP_423J2_125_3477_n730), .CO(
        DP_OP_423J2_125_3477_n568), .S(DP_OP_423J2_125_3477_n569) );
  FADDX1_HVT DP_OP_423J2_125_3477_U465 ( .A(DP_OP_423J2_125_3477_n599), .B(
        DP_OP_423J2_125_3477_n601), .CI(DP_OP_423J2_125_3477_n597), .CO(
        DP_OP_423J2_125_3477_n566), .S(DP_OP_423J2_125_3477_n567) );
  FADDX1_HVT DP_OP_423J2_125_3477_U464 ( .A(DP_OP_423J2_125_3477_n595), .B(
        DP_OP_423J2_125_3477_n589), .CI(DP_OP_423J2_125_3477_n593), .CO(
        DP_OP_423J2_125_3477_n564), .S(DP_OP_423J2_125_3477_n565) );
  FADDX1_HVT DP_OP_423J2_125_3477_U463 ( .A(DP_OP_423J2_125_3477_n587), .B(
        DP_OP_423J2_125_3477_n591), .CI(DP_OP_423J2_125_3477_n728), .CO(
        DP_OP_423J2_125_3477_n562), .S(DP_OP_423J2_125_3477_n563) );
  FADDX1_HVT DP_OP_423J2_125_3477_U462 ( .A(DP_OP_423J2_125_3477_n726), .B(
        DP_OP_423J2_125_3477_n722), .CI(DP_OP_423J2_125_3477_n585), .CO(
        DP_OP_423J2_125_3477_n560), .S(DP_OP_423J2_125_3477_n561) );
  FADDX1_HVT DP_OP_423J2_125_3477_U461 ( .A(DP_OP_423J2_125_3477_n724), .B(
        DP_OP_423J2_125_3477_n720), .CI(DP_OP_423J2_125_3477_n718), .CO(
        DP_OP_423J2_125_3477_n558), .S(DP_OP_423J2_125_3477_n559) );
  FADDX1_HVT DP_OP_423J2_125_3477_U460 ( .A(DP_OP_423J2_125_3477_n716), .B(
        DP_OP_423J2_125_3477_n583), .CI(DP_OP_423J2_125_3477_n581), .CO(
        DP_OP_423J2_125_3477_n556), .S(DP_OP_423J2_125_3477_n557) );
  FADDX1_HVT DP_OP_423J2_125_3477_U459 ( .A(DP_OP_423J2_125_3477_n714), .B(
        DP_OP_423J2_125_3477_n712), .CI(DP_OP_423J2_125_3477_n710), .CO(
        DP_OP_423J2_125_3477_n554), .S(DP_OP_423J2_125_3477_n555) );
  FADDX1_HVT DP_OP_423J2_125_3477_U458 ( .A(DP_OP_423J2_125_3477_n708), .B(
        DP_OP_423J2_125_3477_n579), .CI(DP_OP_423J2_125_3477_n706), .CO(
        DP_OP_423J2_125_3477_n552), .S(DP_OP_423J2_125_3477_n553) );
  FADDX1_HVT DP_OP_423J2_125_3477_U457 ( .A(DP_OP_423J2_125_3477_n577), .B(
        DP_OP_423J2_125_3477_n704), .CI(DP_OP_423J2_125_3477_n575), .CO(
        DP_OP_423J2_125_3477_n550), .S(DP_OP_423J2_125_3477_n551) );
  FADDX1_HVT DP_OP_423J2_125_3477_U456 ( .A(DP_OP_423J2_125_3477_n702), .B(
        DP_OP_423J2_125_3477_n571), .CI(DP_OP_423J2_125_3477_n569), .CO(
        DP_OP_423J2_125_3477_n548), .S(DP_OP_423J2_125_3477_n549) );
  FADDX1_HVT DP_OP_423J2_125_3477_U455 ( .A(DP_OP_423J2_125_3477_n573), .B(
        DP_OP_423J2_125_3477_n567), .CI(DP_OP_423J2_125_3477_n700), .CO(
        DP_OP_423J2_125_3477_n546), .S(DP_OP_423J2_125_3477_n547) );
  FADDX1_HVT DP_OP_423J2_125_3477_U454 ( .A(DP_OP_423J2_125_3477_n565), .B(
        DP_OP_423J2_125_3477_n698), .CI(DP_OP_423J2_125_3477_n563), .CO(
        DP_OP_423J2_125_3477_n544), .S(DP_OP_423J2_125_3477_n545) );
  FADDX1_HVT DP_OP_423J2_125_3477_U453 ( .A(DP_OP_423J2_125_3477_n696), .B(
        DP_OP_423J2_125_3477_n694), .CI(DP_OP_423J2_125_3477_n692), .CO(
        DP_OP_423J2_125_3477_n542), .S(DP_OP_423J2_125_3477_n543) );
  FADDX1_HVT DP_OP_423J2_125_3477_U452 ( .A(DP_OP_423J2_125_3477_n561), .B(
        DP_OP_423J2_125_3477_n690), .CI(DP_OP_423J2_125_3477_n559), .CO(
        DP_OP_423J2_125_3477_n540), .S(DP_OP_423J2_125_3477_n541) );
  FADDX1_HVT DP_OP_423J2_125_3477_U451 ( .A(DP_OP_423J2_125_3477_n688), .B(
        DP_OP_423J2_125_3477_n557), .CI(DP_OP_423J2_125_3477_n555), .CO(
        DP_OP_423J2_125_3477_n538), .S(DP_OP_423J2_125_3477_n539) );
  FADDX1_HVT DP_OP_423J2_125_3477_U450 ( .A(DP_OP_423J2_125_3477_n686), .B(
        DP_OP_423J2_125_3477_n684), .CI(DP_OP_423J2_125_3477_n553), .CO(
        DP_OP_423J2_125_3477_n536), .S(DP_OP_423J2_125_3477_n537) );
  FADDX1_HVT DP_OP_423J2_125_3477_U449 ( .A(DP_OP_423J2_125_3477_n682), .B(
        DP_OP_423J2_125_3477_n551), .CI(DP_OP_423J2_125_3477_n549), .CO(
        DP_OP_423J2_125_3477_n534), .S(DP_OP_423J2_125_3477_n535) );
  FADDX1_HVT DP_OP_423J2_125_3477_U448 ( .A(DP_OP_423J2_125_3477_n680), .B(
        DP_OP_423J2_125_3477_n547), .CI(DP_OP_423J2_125_3477_n678), .CO(
        DP_OP_423J2_125_3477_n532), .S(DP_OP_423J2_125_3477_n533) );
  FADDX1_HVT DP_OP_423J2_125_3477_U447 ( .A(DP_OP_423J2_125_3477_n545), .B(
        DP_OP_423J2_125_3477_n676), .CI(DP_OP_423J2_125_3477_n543), .CO(
        DP_OP_423J2_125_3477_n530), .S(DP_OP_423J2_125_3477_n531) );
  FADDX1_HVT DP_OP_423J2_125_3477_U446 ( .A(DP_OP_423J2_125_3477_n674), .B(
        DP_OP_423J2_125_3477_n672), .CI(DP_OP_423J2_125_3477_n541), .CO(
        DP_OP_423J2_125_3477_n528), .S(DP_OP_423J2_125_3477_n529) );
  FADDX1_HVT DP_OP_423J2_125_3477_U445 ( .A(DP_OP_423J2_125_3477_n670), .B(
        DP_OP_423J2_125_3477_n539), .CI(DP_OP_423J2_125_3477_n537), .CO(
        DP_OP_423J2_125_3477_n526), .S(DP_OP_423J2_125_3477_n527) );
  FADDX1_HVT DP_OP_423J2_125_3477_U444 ( .A(DP_OP_423J2_125_3477_n668), .B(
        DP_OP_423J2_125_3477_n535), .CI(DP_OP_423J2_125_3477_n666), .CO(
        DP_OP_423J2_125_3477_n524), .S(DP_OP_423J2_125_3477_n525) );
  FADDX1_HVT DP_OP_423J2_125_3477_U443 ( .A(DP_OP_423J2_125_3477_n533), .B(
        DP_OP_423J2_125_3477_n664), .CI(DP_OP_423J2_125_3477_n531), .CO(
        DP_OP_423J2_125_3477_n522), .S(DP_OP_423J2_125_3477_n523) );
  FADDX1_HVT DP_OP_423J2_125_3477_U442 ( .A(DP_OP_423J2_125_3477_n662), .B(
        DP_OP_423J2_125_3477_n529), .CI(DP_OP_423J2_125_3477_n660), .CO(
        DP_OP_423J2_125_3477_n520), .S(DP_OP_423J2_125_3477_n521) );
  FADDX1_HVT DP_OP_423J2_125_3477_U439 ( .A(DP_OP_423J2_125_3477_n521), .B(
        DP_OP_423J2_125_3477_n519), .CI(DP_OP_423J2_125_3477_n652), .CO(
        DP_OP_423J2_125_3477_n514), .S(DP_OP_423J2_125_3477_n515) );
  FADDX1_HVT DP_OP_423J2_125_3477_U436 ( .A(DP_OP_423J2_125_3477_n3026), .B(
        DP_OP_423J2_125_3477_n1970), .CI(DP_OP_423J2_125_3477_n511), .CO(
        DP_OP_423J2_125_3477_n508), .S(DP_OP_423J2_125_3477_n509) );
  FADDX1_HVT DP_OP_423J2_125_3477_U435 ( .A(DP_OP_423J2_125_3477_n2058), .B(
        DP_OP_423J2_125_3477_n2982), .CI(DP_OP_423J2_125_3477_n2410), .CO(
        DP_OP_423J2_125_3477_n506), .S(DP_OP_423J2_125_3477_n507) );
  FADDX1_HVT DP_OP_423J2_125_3477_U434 ( .A(DP_OP_423J2_125_3477_n2542), .B(
        DP_OP_423J2_125_3477_n2938), .CI(DP_OP_423J2_125_3477_n2894), .CO(
        DP_OP_423J2_125_3477_n504), .S(DP_OP_423J2_125_3477_n505) );
  FADDX1_HVT DP_OP_423J2_125_3477_U433 ( .A(DP_OP_423J2_125_3477_n2366), .B(
        DP_OP_423J2_125_3477_n2850), .CI(DP_OP_423J2_125_3477_n2806), .CO(
        DP_OP_423J2_125_3477_n502), .S(DP_OP_423J2_125_3477_n503) );
  FADDX1_HVT DP_OP_423J2_125_3477_U432 ( .A(DP_OP_423J2_125_3477_n2234), .B(
        DP_OP_423J2_125_3477_n2014), .CI(DP_OP_423J2_125_3477_n2762), .CO(
        DP_OP_423J2_125_3477_n500), .S(DP_OP_423J2_125_3477_n501) );
  FADDX1_HVT DP_OP_423J2_125_3477_U431 ( .A(DP_OP_423J2_125_3477_n2718), .B(
        DP_OP_423J2_125_3477_n2674), .CI(DP_OP_423J2_125_3477_n2630), .CO(
        DP_OP_423J2_125_3477_n498), .S(DP_OP_423J2_125_3477_n499) );
  FADDX1_HVT DP_OP_423J2_125_3477_U430 ( .A(DP_OP_423J2_125_3477_n2278), .B(
        DP_OP_423J2_125_3477_n2102), .CI(DP_OP_423J2_125_3477_n2146), .CO(
        DP_OP_423J2_125_3477_n496), .S(DP_OP_423J2_125_3477_n497) );
  FADDX1_HVT DP_OP_423J2_125_3477_U429 ( .A(DP_OP_423J2_125_3477_n2190), .B(
        DP_OP_423J2_125_3477_n2586), .CI(DP_OP_423J2_125_3477_n2498), .CO(
        DP_OP_423J2_125_3477_n494), .S(DP_OP_423J2_125_3477_n495) );
  FADDX1_HVT DP_OP_423J2_125_3477_U428 ( .A(DP_OP_423J2_125_3477_n2322), .B(
        DP_OP_423J2_125_3477_n2454), .CI(DP_OP_423J2_125_3477_n646), .CO(
        DP_OP_423J2_125_3477_n492), .S(DP_OP_423J2_125_3477_n493) );
  FADDX1_HVT DP_OP_423J2_125_3477_U427 ( .A(DP_OP_423J2_125_3477_n644), .B(
        DP_OP_423J2_125_3477_n614), .CI(DP_OP_423J2_125_3477_n642), .CO(
        DP_OP_423J2_125_3477_n490), .S(DP_OP_423J2_125_3477_n491) );
  FADDX1_HVT DP_OP_423J2_125_3477_U426 ( .A(DP_OP_423J2_125_3477_n640), .B(
        DP_OP_423J2_125_3477_n616), .CI(DP_OP_423J2_125_3477_n618), .CO(
        DP_OP_423J2_125_3477_n488), .S(DP_OP_423J2_125_3477_n489) );
  FADDX1_HVT DP_OP_423J2_125_3477_U425 ( .A(DP_OP_423J2_125_3477_n638), .B(
        DP_OP_423J2_125_3477_n620), .CI(DP_OP_423J2_125_3477_n622), .CO(
        DP_OP_423J2_125_3477_n486), .S(DP_OP_423J2_125_3477_n487) );
  FADDX1_HVT DP_OP_423J2_125_3477_U424 ( .A(DP_OP_423J2_125_3477_n636), .B(
        DP_OP_423J2_125_3477_n624), .CI(DP_OP_423J2_125_3477_n626), .CO(
        DP_OP_423J2_125_3477_n484), .S(DP_OP_423J2_125_3477_n485) );
  FADDX1_HVT DP_OP_423J2_125_3477_U423 ( .A(DP_OP_423J2_125_3477_n634), .B(
        DP_OP_423J2_125_3477_n628), .CI(DP_OP_423J2_125_3477_n630), .CO(
        DP_OP_423J2_125_3477_n482), .S(DP_OP_423J2_125_3477_n483) );
  FADDX1_HVT DP_OP_423J2_125_3477_U422 ( .A(DP_OP_423J2_125_3477_n632), .B(
        DP_OP_423J2_125_3477_n509), .CI(DP_OP_423J2_125_3477_n505), .CO(
        DP_OP_423J2_125_3477_n480), .S(DP_OP_423J2_125_3477_n481) );
  FADDX1_HVT DP_OP_423J2_125_3477_U421 ( .A(DP_OP_423J2_125_3477_n501), .B(
        DP_OP_423J2_125_3477_n495), .CI(DP_OP_423J2_125_3477_n497), .CO(
        DP_OP_423J2_125_3477_n478), .S(DP_OP_423J2_125_3477_n479) );
  FADDX1_HVT DP_OP_423J2_125_3477_U420 ( .A(DP_OP_423J2_125_3477_n499), .B(
        DP_OP_423J2_125_3477_n507), .CI(DP_OP_423J2_125_3477_n503), .CO(
        DP_OP_423J2_125_3477_n476), .S(DP_OP_423J2_125_3477_n477) );
  FADDX1_HVT DP_OP_423J2_125_3477_U419 ( .A(DP_OP_423J2_125_3477_n612), .B(
        DP_OP_423J2_125_3477_n610), .CI(DP_OP_423J2_125_3477_n602), .CO(
        DP_OP_423J2_125_3477_n474), .S(DP_OP_423J2_125_3477_n475) );
  FADDX1_HVT DP_OP_423J2_125_3477_U418 ( .A(DP_OP_423J2_125_3477_n608), .B(
        DP_OP_423J2_125_3477_n604), .CI(DP_OP_423J2_125_3477_n606), .CO(
        DP_OP_423J2_125_3477_n472), .S(DP_OP_423J2_125_3477_n473) );
  FADDX1_HVT DP_OP_423J2_125_3477_U417 ( .A(DP_OP_423J2_125_3477_n600), .B(
        DP_OP_423J2_125_3477_n596), .CI(DP_OP_423J2_125_3477_n493), .CO(
        DP_OP_423J2_125_3477_n470), .S(DP_OP_423J2_125_3477_n471) );
  FADDX1_HVT DP_OP_423J2_125_3477_U416 ( .A(DP_OP_423J2_125_3477_n598), .B(
        DP_OP_423J2_125_3477_n594), .CI(DP_OP_423J2_125_3477_n491), .CO(
        DP_OP_423J2_125_3477_n468), .S(DP_OP_423J2_125_3477_n469) );
  FADDX1_HVT DP_OP_423J2_125_3477_U415 ( .A(DP_OP_423J2_125_3477_n592), .B(
        DP_OP_423J2_125_3477_n485), .CI(DP_OP_423J2_125_3477_n487), .CO(
        DP_OP_423J2_125_3477_n466), .S(DP_OP_423J2_125_3477_n467) );
  FADDX1_HVT DP_OP_423J2_125_3477_U414 ( .A(DP_OP_423J2_125_3477_n590), .B(
        DP_OP_423J2_125_3477_n489), .CI(DP_OP_423J2_125_3477_n483), .CO(
        DP_OP_423J2_125_3477_n464), .S(DP_OP_423J2_125_3477_n465) );
  FADDX1_HVT DP_OP_423J2_125_3477_U413 ( .A(DP_OP_423J2_125_3477_n588), .B(
        DP_OP_423J2_125_3477_n586), .CI(DP_OP_423J2_125_3477_n584), .CO(
        DP_OP_423J2_125_3477_n462), .S(DP_OP_423J2_125_3477_n463) );
  FADDX1_HVT DP_OP_423J2_125_3477_U412 ( .A(DP_OP_423J2_125_3477_n481), .B(
        DP_OP_423J2_125_3477_n477), .CI(DP_OP_423J2_125_3477_n582), .CO(
        DP_OP_423J2_125_3477_n460), .S(DP_OP_423J2_125_3477_n461) );
  FADDX1_HVT DP_OP_423J2_125_3477_U411 ( .A(DP_OP_423J2_125_3477_n479), .B(
        DP_OP_423J2_125_3477_n580), .CI(DP_OP_423J2_125_3477_n578), .CO(
        DP_OP_423J2_125_3477_n458), .S(DP_OP_423J2_125_3477_n459) );
  FADDX1_HVT DP_OP_423J2_125_3477_U410 ( .A(DP_OP_423J2_125_3477_n576), .B(
        DP_OP_423J2_125_3477_n475), .CI(DP_OP_423J2_125_3477_n473), .CO(
        DP_OP_423J2_125_3477_n456), .S(DP_OP_423J2_125_3477_n457) );
  FADDX1_HVT DP_OP_423J2_125_3477_U409 ( .A(DP_OP_423J2_125_3477_n574), .B(
        DP_OP_423J2_125_3477_n570), .CI(DP_OP_423J2_125_3477_n568), .CO(
        DP_OP_423J2_125_3477_n454), .S(DP_OP_423J2_125_3477_n455) );
  FADDX1_HVT DP_OP_423J2_125_3477_U408 ( .A(DP_OP_423J2_125_3477_n572), .B(
        DP_OP_423J2_125_3477_n566), .CI(DP_OP_423J2_125_3477_n471), .CO(
        DP_OP_423J2_125_3477_n452), .S(DP_OP_423J2_125_3477_n453) );
  FADDX1_HVT DP_OP_423J2_125_3477_U407 ( .A(DP_OP_423J2_125_3477_n469), .B(
        DP_OP_423J2_125_3477_n564), .CI(DP_OP_423J2_125_3477_n562), .CO(
        DP_OP_423J2_125_3477_n450), .S(DP_OP_423J2_125_3477_n451) );
  FADDX1_HVT DP_OP_423J2_125_3477_U406 ( .A(DP_OP_423J2_125_3477_n467), .B(
        DP_OP_423J2_125_3477_n465), .CI(DP_OP_423J2_125_3477_n463), .CO(
        DP_OP_423J2_125_3477_n448), .S(DP_OP_423J2_125_3477_n449) );
  FADDX1_HVT DP_OP_423J2_125_3477_U405 ( .A(DP_OP_423J2_125_3477_n560), .B(
        DP_OP_423J2_125_3477_n558), .CI(DP_OP_423J2_125_3477_n461), .CO(
        DP_OP_423J2_125_3477_n446), .S(DP_OP_423J2_125_3477_n447) );
  FADDX1_HVT DP_OP_423J2_125_3477_U404 ( .A(DP_OP_423J2_125_3477_n556), .B(
        DP_OP_423J2_125_3477_n459), .CI(DP_OP_423J2_125_3477_n554), .CO(
        DP_OP_423J2_125_3477_n444), .S(DP_OP_423J2_125_3477_n445) );
  FADDX1_HVT DP_OP_423J2_125_3477_U402 ( .A(DP_OP_423J2_125_3477_n548), .B(
        DP_OP_423J2_125_3477_n455), .CI(DP_OP_423J2_125_3477_n453), .CO(
        DP_OP_423J2_125_3477_n440), .S(DP_OP_423J2_125_3477_n441) );
  FADDX1_HVT DP_OP_423J2_125_3477_U401 ( .A(DP_OP_423J2_125_3477_n546), .B(
        DP_OP_423J2_125_3477_n451), .CI(DP_OP_423J2_125_3477_n544), .CO(
        DP_OP_423J2_125_3477_n438), .S(DP_OP_423J2_125_3477_n439) );
  FADDX1_HVT DP_OP_423J2_125_3477_U400 ( .A(DP_OP_423J2_125_3477_n449), .B(
        DP_OP_423J2_125_3477_n542), .CI(DP_OP_423J2_125_3477_n540), .CO(
        DP_OP_423J2_125_3477_n436), .S(DP_OP_423J2_125_3477_n437) );
  FADDX1_HVT DP_OP_423J2_125_3477_U399 ( .A(DP_OP_423J2_125_3477_n447), .B(
        DP_OP_423J2_125_3477_n538), .CI(DP_OP_423J2_125_3477_n445), .CO(
        DP_OP_423J2_125_3477_n434), .S(DP_OP_423J2_125_3477_n435) );
  FADDX1_HVT DP_OP_423J2_125_3477_U397 ( .A(DP_OP_423J2_125_3477_n441), .B(
        DP_OP_423J2_125_3477_n532), .CI(DP_OP_423J2_125_3477_n439), .CO(
        DP_OP_423J2_125_3477_n430), .S(DP_OP_423J2_125_3477_n431) );
  FADDX1_HVT DP_OP_423J2_125_3477_U396 ( .A(DP_OP_423J2_125_3477_n530), .B(
        DP_OP_423J2_125_3477_n437), .CI(DP_OP_423J2_125_3477_n528), .CO(
        DP_OP_423J2_125_3477_n428), .S(DP_OP_423J2_125_3477_n429) );
  FADDX1_HVT DP_OP_423J2_125_3477_U395 ( .A(DP_OP_423J2_125_3477_n435), .B(
        DP_OP_423J2_125_3477_n526), .CI(DP_OP_423J2_125_3477_n433), .CO(
        DP_OP_423J2_125_3477_n426), .S(DP_OP_423J2_125_3477_n427) );
  FADDX1_HVT DP_OP_423J2_125_3477_U394 ( .A(DP_OP_423J2_125_3477_n524), .B(
        DP_OP_423J2_125_3477_n431), .CI(DP_OP_423J2_125_3477_n522), .CO(
        DP_OP_423J2_125_3477_n424), .S(DP_OP_423J2_125_3477_n425) );
  FADDX1_HVT DP_OP_423J2_125_3477_U393 ( .A(DP_OP_423J2_125_3477_n429), .B(
        DP_OP_423J2_125_3477_n520), .CI(DP_OP_423J2_125_3477_n427), .CO(
        DP_OP_423J2_125_3477_n422), .S(DP_OP_423J2_125_3477_n423) );
  FADDX1_HVT DP_OP_423J2_125_3477_U392 ( .A(DP_OP_423J2_125_3477_n518), .B(
        DP_OP_423J2_125_3477_n425), .CI(DP_OP_423J2_125_3477_n516), .CO(
        DP_OP_423J2_125_3477_n420), .S(DP_OP_423J2_125_3477_n421) );
  FADDX1_HVT DP_OP_423J2_125_3477_U391 ( .A(DP_OP_423J2_125_3477_n423), .B(
        DP_OP_423J2_125_3477_n514), .CI(DP_OP_423J2_125_3477_n421), .CO(
        DP_OP_423J2_125_3477_n418), .S(DP_OP_423J2_125_3477_n419) );
  FADDX1_HVT DP_OP_423J2_125_3477_U390 ( .A(DP_OP_423J2_125_3477_n1926), .B(
        DP_OP_423J2_125_3477_n510), .CI(DP_OP_423J2_125_3477_n508), .CO(
        DP_OP_423J2_125_3477_n416), .S(DP_OP_423J2_125_3477_n417) );
  FADDX1_HVT DP_OP_423J2_125_3477_U389 ( .A(DP_OP_423J2_125_3477_n498), .B(
        DP_OP_423J2_125_3477_n494), .CI(DP_OP_423J2_125_3477_n506), .CO(
        DP_OP_423J2_125_3477_n414), .S(DP_OP_423J2_125_3477_n415) );
  FADDX1_HVT DP_OP_423J2_125_3477_U388 ( .A(DP_OP_423J2_125_3477_n504), .B(
        DP_OP_423J2_125_3477_n502), .CI(DP_OP_423J2_125_3477_n500), .CO(
        DP_OP_423J2_125_3477_n412), .S(DP_OP_423J2_125_3477_n413) );
  FADDX1_HVT DP_OP_423J2_125_3477_U387 ( .A(DP_OP_423J2_125_3477_n496), .B(
        DP_OP_423J2_125_3477_n492), .CI(DP_OP_423J2_125_3477_n490), .CO(
        DP_OP_423J2_125_3477_n410), .S(DP_OP_423J2_125_3477_n411) );
  FADDX1_HVT DP_OP_423J2_125_3477_U386 ( .A(DP_OP_423J2_125_3477_n488), .B(
        DP_OP_423J2_125_3477_n486), .CI(DP_OP_423J2_125_3477_n484), .CO(
        DP_OP_423J2_125_3477_n408), .S(DP_OP_423J2_125_3477_n409) );
  FADDX1_HVT DP_OP_423J2_125_3477_U385 ( .A(DP_OP_423J2_125_3477_n482), .B(
        DP_OP_423J2_125_3477_n417), .CI(DP_OP_423J2_125_3477_n480), .CO(
        DP_OP_423J2_125_3477_n406), .S(DP_OP_423J2_125_3477_n407) );
  FADDX1_HVT DP_OP_423J2_125_3477_U384 ( .A(DP_OP_423J2_125_3477_n478), .B(
        DP_OP_423J2_125_3477_n413), .CI(DP_OP_423J2_125_3477_n415), .CO(
        DP_OP_423J2_125_3477_n404), .S(DP_OP_423J2_125_3477_n405) );
  FADDX1_HVT DP_OP_423J2_125_3477_U383 ( .A(DP_OP_423J2_125_3477_n476), .B(
        DP_OP_423J2_125_3477_n474), .CI(DP_OP_423J2_125_3477_n472), .CO(
        DP_OP_423J2_125_3477_n402), .S(DP_OP_423J2_125_3477_n403) );
  FADDX1_HVT DP_OP_423J2_125_3477_U382 ( .A(DP_OP_423J2_125_3477_n470), .B(
        DP_OP_423J2_125_3477_n411), .CI(DP_OP_423J2_125_3477_n468), .CO(
        DP_OP_423J2_125_3477_n400), .S(DP_OP_423J2_125_3477_n401) );
  FADDX1_HVT DP_OP_423J2_125_3477_U381 ( .A(DP_OP_423J2_125_3477_n466), .B(
        DP_OP_423J2_125_3477_n409), .CI(DP_OP_423J2_125_3477_n464), .CO(
        DP_OP_423J2_125_3477_n398), .S(DP_OP_423J2_125_3477_n399) );
  FADDX1_HVT DP_OP_423J2_125_3477_U380 ( .A(DP_OP_423J2_125_3477_n462), .B(
        DP_OP_423J2_125_3477_n407), .CI(DP_OP_423J2_125_3477_n460), .CO(
        DP_OP_423J2_125_3477_n396), .S(DP_OP_423J2_125_3477_n397) );
  FADDX1_HVT DP_OP_423J2_125_3477_U379 ( .A(DP_OP_423J2_125_3477_n405), .B(
        DP_OP_423J2_125_3477_n458), .CI(DP_OP_423J2_125_3477_n456), .CO(
        DP_OP_423J2_125_3477_n394), .S(DP_OP_423J2_125_3477_n395) );
  FADDX1_HVT DP_OP_423J2_125_3477_U378 ( .A(DP_OP_423J2_125_3477_n403), .B(
        DP_OP_423J2_125_3477_n454), .CI(DP_OP_423J2_125_3477_n452), .CO(
        DP_OP_423J2_125_3477_n392), .S(DP_OP_423J2_125_3477_n393) );
  FADDX1_HVT DP_OP_423J2_125_3477_U377 ( .A(DP_OP_423J2_125_3477_n401), .B(
        DP_OP_423J2_125_3477_n450), .CI(DP_OP_423J2_125_3477_n399), .CO(
        DP_OP_423J2_125_3477_n390), .S(DP_OP_423J2_125_3477_n391) );
  FADDX1_HVT DP_OP_423J2_125_3477_U376 ( .A(DP_OP_423J2_125_3477_n448), .B(
        DP_OP_423J2_125_3477_n397), .CI(DP_OP_423J2_125_3477_n446), .CO(
        DP_OP_423J2_125_3477_n388), .S(DP_OP_423J2_125_3477_n389) );
  FADDX1_HVT DP_OP_423J2_125_3477_U375 ( .A(DP_OP_423J2_125_3477_n395), .B(
        DP_OP_423J2_125_3477_n444), .CI(DP_OP_423J2_125_3477_n442), .CO(
        DP_OP_423J2_125_3477_n386), .S(DP_OP_423J2_125_3477_n387) );
  FADDX1_HVT DP_OP_423J2_125_3477_U374 ( .A(DP_OP_423J2_125_3477_n393), .B(
        DP_OP_423J2_125_3477_n440), .CI(DP_OP_423J2_125_3477_n438), .CO(
        DP_OP_423J2_125_3477_n384), .S(DP_OP_423J2_125_3477_n385) );
  FADDX1_HVT DP_OP_423J2_125_3477_U373 ( .A(DP_OP_423J2_125_3477_n391), .B(
        DP_OP_423J2_125_3477_n436), .CI(DP_OP_423J2_125_3477_n389), .CO(
        DP_OP_423J2_125_3477_n382), .S(DP_OP_423J2_125_3477_n383) );
  FADDX1_HVT DP_OP_423J2_125_3477_U372 ( .A(DP_OP_423J2_125_3477_n434), .B(
        DP_OP_423J2_125_3477_n387), .CI(DP_OP_423J2_125_3477_n432), .CO(
        DP_OP_423J2_125_3477_n380), .S(DP_OP_423J2_125_3477_n381) );
  FADDX1_HVT DP_OP_423J2_125_3477_U371 ( .A(DP_OP_423J2_125_3477_n430), .B(
        DP_OP_423J2_125_3477_n385), .CI(DP_OP_423J2_125_3477_n383), .CO(
        DP_OP_423J2_125_3477_n378), .S(DP_OP_423J2_125_3477_n379) );
  FADDX1_HVT DP_OP_423J2_125_3477_U370 ( .A(DP_OP_423J2_125_3477_n428), .B(
        DP_OP_423J2_125_3477_n381), .CI(DP_OP_423J2_125_3477_n426), .CO(
        DP_OP_423J2_125_3477_n376), .S(DP_OP_423J2_125_3477_n377) );
  FADDX1_HVT DP_OP_423J2_125_3477_U368 ( .A(DP_OP_423J2_125_3477_n377), .B(
        DP_OP_423J2_125_3477_n420), .CI(DP_OP_423J2_125_3477_n375), .CO(
        DP_OP_423J2_125_3477_n372), .S(DP_OP_423J2_125_3477_n373) );
  FADDX1_HVT DP_OP_423J2_125_3477_U367 ( .A(DP_OP_423J2_125_3477_n1925), .B(
        DP_OP_423J2_125_3477_n416), .CI(DP_OP_423J2_125_3477_n414), .CO(
        DP_OP_423J2_125_3477_n370), .S(DP_OP_423J2_125_3477_n371) );
  FADDX1_HVT DP_OP_423J2_125_3477_U366 ( .A(DP_OP_423J2_125_3477_n412), .B(
        DP_OP_423J2_125_3477_n410), .CI(DP_OP_423J2_125_3477_n408), .CO(
        DP_OP_423J2_125_3477_n368), .S(DP_OP_423J2_125_3477_n369) );
  FADDX1_HVT DP_OP_423J2_125_3477_U365 ( .A(DP_OP_423J2_125_3477_n406), .B(
        DP_OP_423J2_125_3477_n371), .CI(DP_OP_423J2_125_3477_n404), .CO(
        DP_OP_423J2_125_3477_n366), .S(DP_OP_423J2_125_3477_n367) );
  FADDX1_HVT DP_OP_423J2_125_3477_U364 ( .A(DP_OP_423J2_125_3477_n402), .B(
        DP_OP_423J2_125_3477_n400), .CI(DP_OP_423J2_125_3477_n369), .CO(
        DP_OP_423J2_125_3477_n364), .S(DP_OP_423J2_125_3477_n365) );
  FADDX1_HVT DP_OP_423J2_125_3477_U363 ( .A(DP_OP_423J2_125_3477_n398), .B(
        DP_OP_423J2_125_3477_n396), .CI(DP_OP_423J2_125_3477_n367), .CO(
        DP_OP_423J2_125_3477_n362), .S(DP_OP_423J2_125_3477_n363) );
  FADDX1_HVT DP_OP_423J2_125_3477_U362 ( .A(DP_OP_423J2_125_3477_n394), .B(
        DP_OP_423J2_125_3477_n392), .CI(DP_OP_423J2_125_3477_n365), .CO(
        DP_OP_423J2_125_3477_n360), .S(DP_OP_423J2_125_3477_n361) );
  FADDX1_HVT DP_OP_423J2_125_3477_U361 ( .A(DP_OP_423J2_125_3477_n390), .B(
        DP_OP_423J2_125_3477_n363), .CI(DP_OP_423J2_125_3477_n388), .CO(
        DP_OP_423J2_125_3477_n358), .S(DP_OP_423J2_125_3477_n359) );
  FADDX1_HVT DP_OP_423J2_125_3477_U360 ( .A(DP_OP_423J2_125_3477_n386), .B(
        DP_OP_423J2_125_3477_n361), .CI(DP_OP_423J2_125_3477_n384), .CO(
        DP_OP_423J2_125_3477_n356), .S(DP_OP_423J2_125_3477_n357) );
  FADDX1_HVT DP_OP_423J2_125_3477_U358 ( .A(DP_OP_423J2_125_3477_n357), .B(
        DP_OP_423J2_125_3477_n378), .CI(DP_OP_423J2_125_3477_n355), .CO(
        DP_OP_423J2_125_3477_n352), .S(DP_OP_423J2_125_3477_n353) );
  FADDX1_HVT DP_OP_423J2_125_3477_U357 ( .A(DP_OP_423J2_125_3477_n376), .B(
        DP_OP_423J2_125_3477_n374), .CI(DP_OP_423J2_125_3477_n353), .CO(
        DP_OP_423J2_125_3477_n350), .S(DP_OP_423J2_125_3477_n351) );
  FADDX1_HVT DP_OP_423J2_125_3477_U356 ( .A(DP_OP_423J2_125_3477_n1924), .B(
        DP_OP_423J2_125_3477_n370), .CI(DP_OP_423J2_125_3477_n368), .CO(
        DP_OP_423J2_125_3477_n348), .S(DP_OP_423J2_125_3477_n349) );
  FADDX1_HVT DP_OP_423J2_125_3477_U355 ( .A(DP_OP_423J2_125_3477_n366), .B(
        DP_OP_423J2_125_3477_n349), .CI(DP_OP_423J2_125_3477_n364), .CO(
        DP_OP_423J2_125_3477_n346), .S(DP_OP_423J2_125_3477_n347) );
  FADDX1_HVT DP_OP_423J2_125_3477_U354 ( .A(DP_OP_423J2_125_3477_n362), .B(
        DP_OP_423J2_125_3477_n360), .CI(DP_OP_423J2_125_3477_n347), .CO(
        DP_OP_423J2_125_3477_n344), .S(DP_OP_423J2_125_3477_n345) );
  FADDX1_HVT DP_OP_423J2_125_3477_U353 ( .A(DP_OP_423J2_125_3477_n358), .B(
        DP_OP_423J2_125_3477_n345), .CI(DP_OP_423J2_125_3477_n356), .CO(
        DP_OP_423J2_125_3477_n342), .S(DP_OP_423J2_125_3477_n343) );
  FADDX1_HVT DP_OP_423J2_125_3477_U350 ( .A(DP_OP_423J2_125_3477_n339), .B(
        DP_OP_423J2_125_3477_n348), .CI(DP_OP_423J2_125_3477_n346), .CO(
        DP_OP_423J2_125_3477_n336), .S(DP_OP_423J2_125_3477_n337) );
  FADDX1_HVT DP_OP_423J2_125_3477_U349 ( .A(DP_OP_423J2_125_3477_n337), .B(
        DP_OP_423J2_125_3477_n344), .CI(DP_OP_423J2_125_3477_n342), .CO(
        DP_OP_423J2_125_3477_n334), .S(DP_OP_423J2_125_3477_n335) );
  FADDX1_HVT DP_OP_423J2_125_3477_U348 ( .A(DP_OP_423J2_125_3477_n1923), .B(
        DP_OP_423J2_125_3477_n338), .CI(DP_OP_423J2_125_3477_n336), .CO(
        DP_OP_423J2_125_3477_n332), .S(DP_OP_423J2_125_3477_n333) );
  FADDX1_HVT DP_OP_423J2_125_3477_U331 ( .A(DP_OP_423J2_125_3477_n1903), .B(
        DP_OP_423J2_125_3477_n1901), .CI(DP_OP_423J2_125_3477_n1899), .CO(
        DP_OP_423J2_125_3477_n269), .S(n_conv2_sum_b[0]) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U330 ( .A1(DP_OP_423J2_125_3477_n1837), 
        .A2(DP_OP_423J2_125_3477_n1839), .Y(DP_OP_423J2_125_3477_n268) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U329 ( .A1(DP_OP_423J2_125_3477_n1839), .A2(
        DP_OP_423J2_125_3477_n1837), .Y(DP_OP_423J2_125_3477_n267) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U323 ( .A1(DP_OP_423J2_125_3477_n1731), 
        .A2(DP_OP_423J2_125_3477_n1733), .Y(DP_OP_423J2_125_3477_n265) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U315 ( .A1(DP_OP_423J2_125_3477_n1577), 
        .A2(DP_OP_423J2_125_3477_n1579), .Y(DP_OP_423J2_125_3477_n260) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U314 ( .A1(DP_OP_423J2_125_3477_n1579), .A2(
        DP_OP_423J2_125_3477_n1577), .Y(DP_OP_423J2_125_3477_n259) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U309 ( .A1(DP_OP_423J2_125_3477_n1401), 
        .A2(DP_OP_423J2_125_3477_n1403), .Y(DP_OP_423J2_125_3477_n257) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U308 ( .A1(DP_OP_423J2_125_3477_n1403), .A2(
        DP_OP_423J2_125_3477_n1401), .Y(DP_OP_423J2_125_3477_n256) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U301 ( .A1(DP_OP_423J2_125_3477_n1213), 
        .A2(DP_OP_423J2_125_3477_n1215), .Y(DP_OP_423J2_125_3477_n252) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U287 ( .A1(DP_OP_423J2_125_3477_n1018), 
        .A2(DP_OP_423J2_125_3477_n823), .Y(DP_OP_423J2_125_3477_n244) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U274 ( .A1(DP_OP_423J2_125_3477_n513), .A2(
        n891), .Y(DP_OP_423J2_125_3477_n237) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U257 ( .A1(DP_OP_423J2_125_3477_n373), .A2(
        DP_OP_423J2_125_3477_n418), .Y(DP_OP_423J2_125_3477_n226) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U245 ( .A1(DP_OP_423J2_125_3477_n351), .A2(
        DP_OP_423J2_125_3477_n372), .Y(DP_OP_423J2_125_3477_n217) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U235 ( .A1(DP_OP_423J2_125_3477_n350), .A2(
        DP_OP_423J2_125_3477_n341), .Y(DP_OP_423J2_125_3477_n210) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U234 ( .A1(DP_OP_423J2_125_3477_n341), .A2(
        DP_OP_423J2_125_3477_n350), .Y(DP_OP_423J2_125_3477_n209) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U217 ( .A1(DP_OP_423J2_125_3477_n334), .A2(
        DP_OP_423J2_125_3477_n333), .Y(DP_OP_423J2_125_3477_n198) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U216 ( .A1(DP_OP_423J2_125_3477_n333), .A2(
        DP_OP_423J2_125_3477_n334), .Y(DP_OP_423J2_125_3477_n197) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U210 ( .A1(n1677), .A2(
        DP_OP_423J2_125_3477_n286), .Y(DP_OP_423J2_125_3477_n189) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U201 ( .A1(DP_OP_423J2_125_3477_n332), .A2(
        DP_OP_423J2_125_3477_n331), .Y(DP_OP_423J2_125_3477_n185) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U200 ( .A1(DP_OP_423J2_125_3477_n331), .A2(
        DP_OP_423J2_125_3477_n332), .Y(DP_OP_423J2_125_3477_n182) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U194 ( .A1(DP_OP_423J2_125_3477_n182), .A2(
        DP_OP_423J2_125_3477_n189), .Y(DP_OP_423J2_125_3477_n176) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U187 ( .A1(DP_OP_423J2_125_3477_n329), .A2(
        DP_OP_423J2_125_3477_n330), .Y(DP_OP_423J2_125_3477_n174) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U186 ( .A1(DP_OP_423J2_125_3477_n330), .A2(
        DP_OP_423J2_125_3477_n329), .Y(DP_OP_423J2_125_3477_n171) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U177 ( .A1(DP_OP_423J2_125_3477_n327), .A2(
        DP_OP_423J2_125_3477_n328), .Y(DP_OP_423J2_125_3477_n167) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U176 ( .A1(DP_OP_423J2_125_3477_n328), .A2(
        DP_OP_423J2_125_3477_n327), .Y(DP_OP_423J2_125_3477_n166) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U172 ( .A1(DP_OP_423J2_125_3477_n166), .A2(
        DP_OP_423J2_125_3477_n171), .Y(DP_OP_423J2_125_3477_n162) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U168 ( .A1(DP_OP_423J2_125_3477_n176), .A2(
        DP_OP_423J2_125_3477_n162), .Y(DP_OP_423J2_125_3477_n160) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U163 ( .A1(DP_OP_423J2_125_3477_n325), .A2(
        DP_OP_423J2_125_3477_n326), .Y(DP_OP_423J2_125_3477_n156) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U162 ( .A1(DP_OP_423J2_125_3477_n326), .A2(
        DP_OP_423J2_125_3477_n325), .Y(DP_OP_423J2_125_3477_n153) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U153 ( .A1(DP_OP_423J2_125_3477_n323), .A2(
        DP_OP_423J2_125_3477_n324), .Y(DP_OP_423J2_125_3477_n149) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U152 ( .A1(DP_OP_423J2_125_3477_n324), .A2(
        DP_OP_423J2_125_3477_n323), .Y(DP_OP_423J2_125_3477_n148) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U150 ( .A1(DP_OP_423J2_125_3477_n281), .A2(
        DP_OP_423J2_125_3477_n149), .Y(DP_OP_423J2_125_3477_n17) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U148 ( .A1(DP_OP_423J2_125_3477_n148), .A2(
        DP_OP_423J2_125_3477_n153), .Y(DP_OP_423J2_125_3477_n146) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U146 ( .A1(DP_OP_423J2_125_3477_n162), .A2(
        DP_OP_423J2_125_3477_n146), .Y(DP_OP_423J2_125_3477_n144) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U142 ( .A1(DP_OP_423J2_125_3477_n176), .A2(
        DP_OP_423J2_125_3477_n142), .Y(DP_OP_423J2_125_3477_n140) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U137 ( .A1(DP_OP_423J2_125_3477_n321), .A2(
        DP_OP_423J2_125_3477_n322), .Y(DP_OP_423J2_125_3477_n136) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U136 ( .A1(DP_OP_423J2_125_3477_n322), .A2(
        DP_OP_423J2_125_3477_n321), .Y(DP_OP_423J2_125_3477_n133) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U127 ( .A1(DP_OP_423J2_125_3477_n319), .A2(
        DP_OP_423J2_125_3477_n320), .Y(DP_OP_423J2_125_3477_n129) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U126 ( .A1(DP_OP_423J2_125_3477_n320), .A2(
        DP_OP_423J2_125_3477_n319), .Y(DP_OP_423J2_125_3477_n128) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U122 ( .A1(DP_OP_423J2_125_3477_n128), .A2(
        DP_OP_423J2_125_3477_n133), .Y(DP_OP_423J2_125_3477_n126) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U115 ( .A1(DP_OP_423J2_125_3477_n317), .A2(
        DP_OP_423J2_125_3477_n318), .Y(DP_OP_423J2_125_3477_n120) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U112 ( .A1(n1673), .A2(
        DP_OP_423J2_125_3477_n120), .Y(DP_OP_423J2_125_3477_n14) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U108 ( .A1(DP_OP_423J2_125_3477_n126), .A2(
        n1673), .Y(DP_OP_423J2_125_3477_n115) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U106 ( .A1(DP_OP_423J2_125_3477_n115), .A2(
        DP_OP_423J2_125_3477_n144), .Y(DP_OP_423J2_125_3477_n111) );
  AOI21X1_HVT DP_OP_423J2_125_3477_U103 ( .A1(DP_OP_423J2_125_3477_n177), .A2(
        DP_OP_423J2_125_3477_n111), .A3(DP_OP_423J2_125_3477_n114), .Y(
        DP_OP_423J2_125_3477_n110) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U102 ( .A1(DP_OP_423J2_125_3477_n176), .A2(
        DP_OP_423J2_125_3477_n111), .Y(DP_OP_423J2_125_3477_n109) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U97 ( .A1(DP_OP_423J2_125_3477_n315), .A2(
        DP_OP_423J2_125_3477_n316), .Y(DP_OP_423J2_125_3477_n105) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U96 ( .A1(DP_OP_423J2_125_3477_n316), .A2(
        DP_OP_423J2_125_3477_n315), .Y(DP_OP_423J2_125_3477_n102) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U87 ( .A1(n1382), .A2(
        DP_OP_423J2_125_3477_n314), .Y(DP_OP_423J2_125_3477_n98) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U86 ( .A1(DP_OP_423J2_125_3477_n314), .A2(
        n1382), .Y(DP_OP_423J2_125_3477_n97) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U82 ( .A1(DP_OP_423J2_125_3477_n97), .A2(
        DP_OP_423J2_125_3477_n102), .Y(DP_OP_423J2_125_3477_n95) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U75 ( .A1(DP_OP_423J2_125_3477_n311), .A2(
        DP_OP_423J2_125_3477_n312), .Y(DP_OP_423J2_125_3477_n89) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U68 ( .A1(DP_OP_423J2_125_3477_n95), .A2(
        n1672), .Y(DP_OP_423J2_125_3477_n82) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U61 ( .A1(DP_OP_423J2_125_3477_n309), .A2(
        DP_OP_423J2_125_3477_n310), .Y(DP_OP_423J2_125_3477_n78) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U60 ( .A1(DP_OP_423J2_125_3477_n310), .A2(
        DP_OP_423J2_125_3477_n309), .Y(DP_OP_423J2_125_3477_n77) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U54 ( .A1(DP_OP_423J2_125_3477_n111), .A2(
        DP_OP_423J2_125_3477_n75), .Y(DP_OP_423J2_125_3477_n73) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U45 ( .A1(DP_OP_423J2_125_3477_n307), .A2(
        DP_OP_423J2_125_3477_n308), .Y(DP_OP_423J2_125_3477_n65) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U42 ( .A1(n1671), .A2(
        DP_OP_423J2_125_3477_n65), .Y(DP_OP_423J2_125_3477_n9) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U38 ( .A1(DP_OP_423J2_125_3477_n71), .A2(
        n1671), .Y(DP_OP_423J2_125_3477_n60) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U34 ( .A1(n1677), .A2(
        DP_OP_423J2_125_3477_n58), .Y(DP_OP_423J2_125_3477_n56) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U29 ( .A1(DP_OP_423J2_125_3477_n305), .A2(
        DP_OP_423J2_125_3477_n306), .Y(DP_OP_423J2_125_3477_n52) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U28 ( .A1(DP_OP_423J2_125_3477_n306), .A2(
        DP_OP_423J2_125_3477_n305), .Y(DP_OP_423J2_125_3477_n51) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U21 ( .A1(DP_OP_423J2_125_3477_n303), .A2(
        DP_OP_423J2_125_3477_n304), .Y(DP_OP_423J2_125_3477_n47) );
  NAND2X0_HVT DP_OP_423J2_125_3477_U9 ( .A1(n1669), .A2(
        DP_OP_423J2_125_3477_n302), .Y(DP_OP_423J2_125_3477_n38) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U311 ( .A1(DP_OP_422J2_124_3477_n261), .A2(
        DP_OP_422J2_124_3477_n259), .A3(DP_OP_422J2_124_3477_n260), .Y(
        DP_OP_422J2_124_3477_n258) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U325 ( .A1(DP_OP_422J2_124_3477_n5), .A2(
        DP_OP_422J2_124_3477_n267), .A3(DP_OP_422J2_124_3477_n268), .Y(
        DP_OP_422J2_124_3477_n266) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U173 ( .A1(DP_OP_422J2_124_3477_n174), .A2(
        DP_OP_422J2_124_3477_n166), .A3(DP_OP_422J2_124_3477_n167), .Y(
        DP_OP_422J2_124_3477_n165) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U83 ( .A1(DP_OP_422J2_124_3477_n105), .A2(
        DP_OP_422J2_124_3477_n97), .A3(DP_OP_422J2_124_3477_n98), .Y(
        DP_OP_422J2_124_3477_n96) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U123 ( .A1(DP_OP_422J2_124_3477_n136), .A2(
        DP_OP_422J2_124_3477_n128), .A3(DP_OP_422J2_124_3477_n129), .Y(
        DP_OP_422J2_124_3477_n127) );
  XNOR2X1_HVT DP_OP_422J2_124_3477_U787 ( .A1(DP_OP_422J2_124_3477_n2502), 
        .A2(DP_OP_422J2_124_3477_n3029), .Y(DP_OP_422J2_124_3477_n1211) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2291 ( .A1(DP_OP_422J2_124_3477_n3058), 
        .A2(n34), .Y(DP_OP_422J2_124_3477_n3050) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2290 ( .A1(DP_OP_422J2_124_3477_n3057), 
        .A2(n34), .Y(DP_OP_422J2_124_3477_n3049) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2289 ( .A1(DP_OP_422J2_124_3477_n3056), .A2(
        n32), .Y(DP_OP_422J2_124_3477_n3048) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2273 ( .A1(DP_OP_422J2_124_3477_n3056), .A2(
        DP_OP_424J2_126_3477_n3065), .Y(DP_OP_422J2_124_3477_n3032) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2272 ( .A1(DP_OP_422J2_124_3477_n3063), .A2(
        n215), .Y(DP_OP_422J2_124_3477_n1728) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2271 ( .A1(DP_OP_423J2_125_3477_n2008), .A2(
        n215), .Y(DP_OP_422J2_124_3477_n3031) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2270 ( .A1(DP_OP_424J2_126_3477_n2095), .A2(
        n215), .Y(DP_OP_422J2_124_3477_n3030) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2269 ( .A1(DP_OP_422J2_124_3477_n3060), .A2(
        n215), .Y(DP_OP_422J2_124_3477_n3029) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2268 ( .A1(DP_OP_422J2_124_3477_n3059), .A2(
        n214), .Y(DP_OP_422J2_124_3477_n3028) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2267 ( .A1(DP_OP_422J2_124_3477_n3058), .A2(
        n215), .Y(DP_OP_422J2_124_3477_n820) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2266 ( .A1(DP_OP_422J2_124_3477_n3057), .A2(
        n215), .Y(DP_OP_422J2_124_3477_n3027) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2265 ( .A1(DP_OP_422J2_124_3477_n3056), 
        .A2(n211), .Y(DP_OP_422J2_124_3477_n3026) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2246 ( .A1(DP_OP_422J2_124_3477_n3015), 
        .A2(n846), .Y(DP_OP_422J2_124_3477_n3007) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2245 ( .A1(DP_OP_422J2_124_3477_n3014), .A2(
        DP_OP_423J2_125_3477_n3025), .Y(DP_OP_422J2_124_3477_n3006) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2202 ( .A1(DP_OP_422J2_124_3477_n2971), 
        .A2(n675), .Y(DP_OP_422J2_124_3477_n2963) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2201 ( .A1(DP_OP_422J2_124_3477_n2970), .A2(
        n677), .Y(DP_OP_422J2_124_3477_n2962) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2158 ( .A1(DP_OP_422J2_124_3477_n2927), 
        .A2(n445), .Y(DP_OP_422J2_124_3477_n2919) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2157 ( .A1(DP_OP_422J2_124_3477_n2926), .A2(
        n445), .Y(DP_OP_422J2_124_3477_n2918) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2142 ( .A1(DP_OP_422J2_124_3477_n2927), 
        .A2(DP_OP_425J2_127_3477_n2935), .Y(DP_OP_422J2_124_3477_n2903) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2139 ( .A1(DP_OP_423J2_125_3477_n2140), .A2(
        n35), .Y(DP_OP_422J2_124_3477_n2900) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2138 ( .A1(DP_OP_425J2_127_3477_n2799), .A2(
        n35), .Y(DP_OP_422J2_124_3477_n2899) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2137 ( .A1(DP_OP_422J2_124_3477_n2930), .A2(
        n35), .Y(DP_OP_422J2_124_3477_n2898) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2136 ( .A1(DP_OP_422J2_124_3477_n2929), .A2(
        n35), .Y(DP_OP_422J2_124_3477_n2897) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2135 ( .A1(DP_OP_422J2_124_3477_n2928), .A2(
        n35), .Y(DP_OP_422J2_124_3477_n2896) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2134 ( .A1(DP_OP_422J2_124_3477_n2927), .A2(
        n35), .Y(DP_OP_422J2_124_3477_n2895) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2133 ( .A1(DP_OP_422J2_124_3477_n2926), 
        .A2(n35), .Y(DP_OP_422J2_124_3477_n2894) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2114 ( .A1(DP_OP_422J2_124_3477_n2883), 
        .A2(DP_OP_422J2_124_3477_n2893), .Y(DP_OP_422J2_124_3477_n2875) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2113 ( .A1(DP_OP_422J2_124_3477_n2882), .A2(
        DP_OP_422J2_124_3477_n2893), .Y(DP_OP_422J2_124_3477_n2874) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2098 ( .A1(DP_OP_422J2_124_3477_n2883), 
        .A2(DP_OP_423J2_125_3477_n2891), .Y(DP_OP_422J2_124_3477_n2859) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2097 ( .A1(DP_OP_422J2_124_3477_n2882), .A2(
        DP_OP_423J2_125_3477_n2891), .Y(DP_OP_422J2_124_3477_n2858) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2096 ( .A1(DP_OP_422J2_124_3477_n2889), .A2(
        DP_OP_423J2_125_3477_n2890), .Y(DP_OP_422J2_124_3477_n2857) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2095 ( .A1(DP_OP_422J2_124_3477_n2888), .A2(
        DP_OP_423J2_125_3477_n2890), .Y(DP_OP_422J2_124_3477_n2856) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2094 ( .A1(DP_OP_422J2_124_3477_n2887), .A2(
        DP_OP_424J2_126_3477_n2890), .Y(DP_OP_422J2_124_3477_n2855) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2093 ( .A1(DP_OP_423J2_125_3477_n2182), .A2(
        DP_OP_423J2_125_3477_n2890), .Y(DP_OP_422J2_124_3477_n2854) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2092 ( .A1(DP_OP_422J2_124_3477_n2885), .A2(
        DP_OP_422J2_124_3477_n2890), .Y(DP_OP_422J2_124_3477_n2853) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2091 ( .A1(DP_OP_422J2_124_3477_n2884), .A2(
        DP_OP_422J2_124_3477_n2890), .Y(DP_OP_422J2_124_3477_n2852) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2090 ( .A1(DP_OP_422J2_124_3477_n2883), .A2(
        DP_OP_422J2_124_3477_n2890), .Y(DP_OP_422J2_124_3477_n2851) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2089 ( .A1(DP_OP_422J2_124_3477_n2882), 
        .A2(DP_OP_422J2_124_3477_n2890), .Y(DP_OP_422J2_124_3477_n2850) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2070 ( .A1(DP_OP_422J2_124_3477_n2839), 
        .A2(DP_OP_423J2_125_3477_n2849), .Y(DP_OP_422J2_124_3477_n2831) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2069 ( .A1(DP_OP_422J2_124_3477_n2838), .A2(
        DP_OP_424J2_126_3477_n2849), .Y(DP_OP_422J2_124_3477_n2830) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2054 ( .A1(DP_OP_422J2_124_3477_n2839), 
        .A2(DP_OP_422J2_124_3477_n2847), .Y(DP_OP_422J2_124_3477_n2815) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2051 ( .A1(DP_OP_423J2_125_3477_n2228), .A2(
        DP_OP_422J2_124_3477_n2846), .Y(DP_OP_422J2_124_3477_n2812) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2050 ( .A1(DP_OP_424J2_126_3477_n2315), .A2(
        DP_OP_422J2_124_3477_n2846), .Y(DP_OP_422J2_124_3477_n2811) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2049 ( .A1(DP_OP_422J2_124_3477_n2842), .A2(
        DP_OP_422J2_124_3477_n2846), .Y(DP_OP_422J2_124_3477_n2810) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2048 ( .A1(DP_OP_422J2_124_3477_n2841), .A2(
        DP_OP_422J2_124_3477_n2846), .Y(DP_OP_422J2_124_3477_n2809) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2047 ( .A1(DP_OP_422J2_124_3477_n2840), .A2(
        DP_OP_422J2_124_3477_n2846), .Y(DP_OP_422J2_124_3477_n2808) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2046 ( .A1(DP_OP_422J2_124_3477_n2839), .A2(
        DP_OP_422J2_124_3477_n2846), .Y(DP_OP_422J2_124_3477_n2807) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2045 ( .A1(DP_OP_422J2_124_3477_n2838), 
        .A2(DP_OP_422J2_124_3477_n2846), .Y(DP_OP_422J2_124_3477_n2806) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2025 ( .A1(DP_OP_422J2_124_3477_n2794), .A2(
        DP_OP_422J2_124_3477_n2805), .Y(DP_OP_422J2_124_3477_n2786) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2019 ( .A1(DP_OP_422J2_124_3477_n2796), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_422J2_124_3477_n2780) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2017 ( .A1(DP_OP_422J2_124_3477_n2794), .A2(
        DP_OP_423J2_125_3477_n2804), .Y(DP_OP_422J2_124_3477_n2778) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2013 ( .A1(DP_OP_422J2_124_3477_n2798), 
        .A2(DP_OP_423J2_125_3477_n2803), .Y(DP_OP_422J2_124_3477_n2774) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2011 ( .A1(DP_OP_422J2_124_3477_n2796), 
        .A2(DP_OP_423J2_125_3477_n2803), .Y(DP_OP_422J2_124_3477_n2772) );
  OR2X1_HVT DP_OP_422J2_124_3477_U2007 ( .A1(DP_OP_422J2_124_3477_n2800), .A2(
        DP_OP_423J2_125_3477_n2802), .Y(DP_OP_422J2_124_3477_n2768) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1982 ( .A1(DP_OP_422J2_124_3477_n2751), 
        .A2(DP_OP_425J2_127_3477_n2761), .Y(DP_OP_422J2_124_3477_n2743) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1981 ( .A1(DP_OP_422J2_124_3477_n2750), .A2(
        n66), .Y(DP_OP_422J2_124_3477_n2742) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1964 ( .A1(DP_OP_424J2_126_3477_n2405), .A2(
        DP_OP_422J2_124_3477_n2758), .Y(DP_OP_422J2_124_3477_n2725) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1961 ( .A1(DP_OP_422J2_124_3477_n2754), .A2(
        DP_OP_422J2_124_3477_n2758), .Y(DP_OP_422J2_124_3477_n2722) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1960 ( .A1(DP_OP_422J2_124_3477_n2753), .A2(
        DP_OP_422J2_124_3477_n2758), .Y(DP_OP_422J2_124_3477_n2721) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1957 ( .A1(DP_OP_422J2_124_3477_n2750), 
        .A2(DP_OP_422J2_124_3477_n2758), .Y(DP_OP_422J2_124_3477_n2718) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1940 ( .A1(DP_OP_422J2_124_3477_n2709), 
        .A2(n597), .Y(DP_OP_422J2_124_3477_n2701) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1938 ( .A1(DP_OP_422J2_124_3477_n2707), 
        .A2(DP_OP_422J2_124_3477_n2717), .Y(DP_OP_422J2_124_3477_n2699) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1937 ( .A1(DP_OP_423J2_125_3477_n2354), .A2(
        n597), .Y(DP_OP_422J2_124_3477_n2698) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1930 ( .A1(DP_OP_422J2_124_3477_n2707), 
        .A2(DP_OP_424J2_126_3477_n2716), .Y(DP_OP_422J2_124_3477_n2691) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1929 ( .A1(DP_OP_423J2_125_3477_n2354), .A2(
        n1341), .Y(DP_OP_422J2_124_3477_n2690) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1924 ( .A1(DP_OP_422J2_124_3477_n2709), 
        .A2(n1440), .Y(DP_OP_422J2_124_3477_n2685) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1923 ( .A1(DP_OP_422J2_124_3477_n2708), 
        .A2(n1440), .Y(DP_OP_422J2_124_3477_n2684) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1920 ( .A1(DP_OP_425J2_127_3477_n2581), .A2(
        DP_OP_422J2_124_3477_n2714), .Y(DP_OP_422J2_124_3477_n2681) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1919 ( .A1(DP_OP_422J2_124_3477_n2712), .A2(
        DP_OP_422J2_124_3477_n2714), .Y(DP_OP_422J2_124_3477_n2680) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1918 ( .A1(DP_OP_424J2_126_3477_n2447), .A2(
        DP_OP_422J2_124_3477_n2714), .Y(DP_OP_422J2_124_3477_n2679) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1917 ( .A1(DP_OP_422J2_124_3477_n2710), .A2(
        DP_OP_422J2_124_3477_n2714), .Y(DP_OP_422J2_124_3477_n2678) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1916 ( .A1(DP_OP_422J2_124_3477_n2709), .A2(
        DP_OP_422J2_124_3477_n2714), .Y(DP_OP_422J2_124_3477_n2677) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1915 ( .A1(DP_OP_422J2_124_3477_n2708), .A2(
        DP_OP_422J2_124_3477_n2714), .Y(DP_OP_422J2_124_3477_n2676) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1914 ( .A1(DP_OP_422J2_124_3477_n2707), .A2(
        DP_OP_422J2_124_3477_n2714), .Y(DP_OP_422J2_124_3477_n2675) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1913 ( .A1(DP_OP_425J2_127_3477_n2574), 
        .A2(DP_OP_422J2_124_3477_n2714), .Y(DP_OP_422J2_124_3477_n2674) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1894 ( .A1(DP_OP_422J2_124_3477_n2663), 
        .A2(DP_OP_422J2_124_3477_n2673), .Y(DP_OP_422J2_124_3477_n2655) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1893 ( .A1(DP_OP_422J2_124_3477_n2662), .A2(
        DP_OP_424J2_126_3477_n2673), .Y(DP_OP_422J2_124_3477_n2654) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1885 ( .A1(DP_OP_422J2_124_3477_n2662), .A2(
        n279), .Y(DP_OP_422J2_124_3477_n2646) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1879 ( .A1(DP_OP_422J2_124_3477_n2664), 
        .A2(DP_OP_425J2_127_3477_n2671), .Y(DP_OP_422J2_124_3477_n2640) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1876 ( .A1(DP_OP_422J2_124_3477_n2669), .A2(
        DP_OP_422J2_124_3477_n2670), .Y(DP_OP_422J2_124_3477_n2637) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1875 ( .A1(DP_OP_425J2_127_3477_n2536), .A2(
        DP_OP_422J2_124_3477_n2670), .Y(DP_OP_422J2_124_3477_n2636) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1874 ( .A1(DP_OP_422J2_124_3477_n2667), .A2(
        DP_OP_422J2_124_3477_n2670), .Y(DP_OP_422J2_124_3477_n2635) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1873 ( .A1(DP_OP_425J2_127_3477_n2534), .A2(
        DP_OP_422J2_124_3477_n2670), .Y(DP_OP_422J2_124_3477_n2634) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1872 ( .A1(DP_OP_422J2_124_3477_n2665), .A2(
        DP_OP_422J2_124_3477_n2670), .Y(DP_OP_422J2_124_3477_n2633) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1871 ( .A1(DP_OP_422J2_124_3477_n2664), .A2(
        n86), .Y(DP_OP_422J2_124_3477_n2632) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1870 ( .A1(DP_OP_422J2_124_3477_n2663), .A2(
        DP_OP_422J2_124_3477_n2670), .Y(DP_OP_422J2_124_3477_n2631) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1869 ( .A1(DP_OP_422J2_124_3477_n2662), 
        .A2(n86), .Y(DP_OP_422J2_124_3477_n2630) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1834 ( .A1(DP_OP_422J2_124_3477_n2619), 
        .A2(DP_OP_422J2_124_3477_n2627), .Y(DP_OP_422J2_124_3477_n2595) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1833 ( .A1(DP_OP_422J2_124_3477_n2618), .A2(
        DP_OP_422J2_124_3477_n2627), .Y(DP_OP_422J2_124_3477_n2594) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1832 ( .A1(DP_OP_422J2_124_3477_n2625), .A2(
        n1331), .Y(DP_OP_422J2_124_3477_n2593) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1831 ( .A1(DP_OP_423J2_125_3477_n2448), .A2(
        DP_OP_422J2_124_3477_n2626), .Y(DP_OP_422J2_124_3477_n2592) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1829 ( .A1(DP_OP_422J2_124_3477_n2622), .A2(
        DP_OP_422J2_124_3477_n2626), .Y(DP_OP_422J2_124_3477_n2590) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1828 ( .A1(DP_OP_422J2_124_3477_n2621), .A2(
        n1331), .Y(DP_OP_422J2_124_3477_n2589) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1827 ( .A1(DP_OP_422J2_124_3477_n2620), .A2(
        DP_OP_422J2_124_3477_n2626), .Y(DP_OP_422J2_124_3477_n2588) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1826 ( .A1(DP_OP_422J2_124_3477_n2619), .A2(
        n1331), .Y(DP_OP_422J2_124_3477_n2587) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1825 ( .A1(DP_OP_422J2_124_3477_n2618), 
        .A2(n1331), .Y(DP_OP_422J2_124_3477_n2586) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1806 ( .A1(DP_OP_422J2_124_3477_n2575), 
        .A2(DP_OP_423J2_125_3477_n2585), .Y(DP_OP_422J2_124_3477_n2567) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1805 ( .A1(DP_OP_422J2_124_3477_n2574), .A2(
        DP_OP_422J2_124_3477_n2585), .Y(DP_OP_422J2_124_3477_n2566) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1797 ( .A1(DP_OP_422J2_124_3477_n2574), .A2(
        n186), .Y(DP_OP_422J2_124_3477_n2558) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1788 ( .A1(DP_OP_423J2_125_3477_n2493), .A2(
        DP_OP_422J2_124_3477_n2582), .Y(DP_OP_422J2_124_3477_n2549) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1787 ( .A1(DP_OP_422J2_124_3477_n2580), .A2(
        DP_OP_422J2_124_3477_n2582), .Y(DP_OP_422J2_124_3477_n2548) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1786 ( .A1(DP_OP_422J2_124_3477_n2579), .A2(
        DP_OP_422J2_124_3477_n2582), .Y(DP_OP_422J2_124_3477_n2547) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1785 ( .A1(DP_OP_422J2_124_3477_n2578), .A2(
        DP_OP_422J2_124_3477_n2582), .Y(DP_OP_422J2_124_3477_n2546) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1784 ( .A1(DP_OP_422J2_124_3477_n2577), .A2(
        DP_OP_422J2_124_3477_n2582), .Y(DP_OP_422J2_124_3477_n2545) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1783 ( .A1(DP_OP_422J2_124_3477_n2576), .A2(
        DP_OP_422J2_124_3477_n2582), .Y(DP_OP_422J2_124_3477_n2544) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1782 ( .A1(DP_OP_422J2_124_3477_n2575), .A2(
        DP_OP_422J2_124_3477_n2582), .Y(DP_OP_422J2_124_3477_n2543) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1781 ( .A1(DP_OP_422J2_124_3477_n2574), 
        .A2(DP_OP_422J2_124_3477_n2582), .Y(DP_OP_422J2_124_3477_n2542) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1761 ( .A1(DP_OP_422J2_124_3477_n2530), .A2(
        DP_OP_422J2_124_3477_n2541), .Y(DP_OP_422J2_124_3477_n2522) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1754 ( .A1(DP_OP_422J2_124_3477_n2531), 
        .A2(DP_OP_424J2_126_3477_n2540), .Y(DP_OP_422J2_124_3477_n2515) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1746 ( .A1(DP_OP_422J2_124_3477_n2531), 
        .A2(n772), .Y(DP_OP_422J2_124_3477_n2507) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1745 ( .A1(DP_OP_422J2_124_3477_n2530), .A2(
        n772), .Y(DP_OP_422J2_124_3477_n2506) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1741 ( .A1(DP_OP_422J2_124_3477_n2534), .A2(
        DP_OP_423J2_125_3477_n2538), .Y(DP_OP_422J2_124_3477_n2502) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1739 ( .A1(DP_OP_422J2_124_3477_n2532), .A2(
        n1335), .Y(DP_OP_422J2_124_3477_n2500) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1738 ( .A1(DP_OP_422J2_124_3477_n2531), .A2(
        n1335), .Y(DP_OP_422J2_124_3477_n2499) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1718 ( .A1(DP_OP_423J2_125_3477_n2531), 
        .A2(DP_OP_425J2_127_3477_n2497), .Y(DP_OP_422J2_124_3477_n2479) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1717 ( .A1(DP_OP_422J2_124_3477_n2486), .A2(
        DP_OP_422J2_124_3477_n2497), .Y(DP_OP_422J2_124_3477_n2478) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1709 ( .A1(DP_OP_422J2_124_3477_n2486), .A2(
        n1491), .Y(DP_OP_422J2_124_3477_n2470) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1702 ( .A1(DP_OP_423J2_125_3477_n2531), 
        .A2(DP_OP_422J2_124_3477_n2495), .Y(DP_OP_422J2_124_3477_n2463) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1701 ( .A1(DP_OP_422J2_124_3477_n2486), .A2(
        DP_OP_422J2_124_3477_n2495), .Y(DP_OP_422J2_124_3477_n2462) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1665 ( .A1(DP_OP_422J2_124_3477_n2442), .A2(
        n1488), .Y(DP_OP_422J2_124_3477_n2426) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1657 ( .A1(DP_OP_422J2_124_3477_n2442), .A2(
        n789), .Y(DP_OP_422J2_124_3477_n2418) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1656 ( .A1(DP_OP_423J2_125_3477_n2581), .A2(
        DP_OP_422J2_124_3477_n2450), .Y(DP_OP_422J2_124_3477_n2417) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1654 ( .A1(DP_OP_423J2_125_3477_n2579), .A2(
        DP_OP_422J2_124_3477_n2450), .Y(DP_OP_422J2_124_3477_n2415) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1653 ( .A1(DP_OP_422J2_124_3477_n2446), .A2(
        DP_OP_422J2_124_3477_n2450), .Y(DP_OP_422J2_124_3477_n2414) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1652 ( .A1(DP_OP_422J2_124_3477_n2445), .A2(
        DP_OP_422J2_124_3477_n2450), .Y(DP_OP_422J2_124_3477_n2413) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1651 ( .A1(DP_OP_422J2_124_3477_n2444), .A2(
        DP_OP_422J2_124_3477_n2450), .Y(DP_OP_422J2_124_3477_n2412) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1650 ( .A1(DP_OP_422J2_124_3477_n2443), .A2(
        DP_OP_422J2_124_3477_n2450), .Y(DP_OP_422J2_124_3477_n2411) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1649 ( .A1(DP_OP_422J2_124_3477_n2442), 
        .A2(DP_OP_422J2_124_3477_n2450), .Y(DP_OP_422J2_124_3477_n2410) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1631 ( .A1(DP_OP_424J2_126_3477_n2532), 
        .A2(DP_OP_422J2_124_3477_n2409), .Y(DP_OP_422J2_124_3477_n2392) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1630 ( .A1(DP_OP_422J2_124_3477_n2399), 
        .A2(DP_OP_422J2_124_3477_n2409), .Y(DP_OP_422J2_124_3477_n2391) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1629 ( .A1(DP_OP_422J2_124_3477_n2398), .A2(
        DP_OP_424J2_126_3477_n2409), .Y(DP_OP_422J2_124_3477_n2390) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1622 ( .A1(DP_OP_422J2_124_3477_n2399), 
        .A2(DP_OP_424J2_126_3477_n2408), .Y(DP_OP_422J2_124_3477_n2383) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1621 ( .A1(DP_OP_422J2_124_3477_n2398), .A2(
        n1333), .Y(DP_OP_422J2_124_3477_n2382) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1614 ( .A1(DP_OP_422J2_124_3477_n2399), 
        .A2(n799), .Y(DP_OP_422J2_124_3477_n2375) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1613 ( .A1(DP_OP_422J2_124_3477_n2398), .A2(
        n799), .Y(DP_OP_422J2_124_3477_n2374) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1612 ( .A1(DP_OP_422J2_124_3477_n2405), .A2(
        n1433), .Y(DP_OP_422J2_124_3477_n2373) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1611 ( .A1(DP_OP_422J2_124_3477_n2404), .A2(
        DP_OP_422J2_124_3477_n2406), .Y(DP_OP_422J2_124_3477_n2372) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1610 ( .A1(DP_OP_424J2_126_3477_n2535), .A2(
        DP_OP_422J2_124_3477_n2406), .Y(DP_OP_422J2_124_3477_n2371) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1609 ( .A1(DP_OP_424J2_126_3477_n2534), .A2(
        n1426), .Y(DP_OP_422J2_124_3477_n2370) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1607 ( .A1(DP_OP_424J2_126_3477_n2532), .A2(
        DP_OP_422J2_124_3477_n2406), .Y(DP_OP_422J2_124_3477_n2368) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1606 ( .A1(DP_OP_422J2_124_3477_n2399), .A2(
        n1426), .Y(DP_OP_422J2_124_3477_n2367) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1605 ( .A1(DP_OP_422J2_124_3477_n2398), 
        .A2(DP_OP_422J2_124_3477_n2406), .Y(DP_OP_422J2_124_3477_n2366) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1587 ( .A1(DP_OP_422J2_124_3477_n2356), 
        .A2(DP_OP_424J2_126_3477_n2365), .Y(DP_OP_422J2_124_3477_n2348) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1586 ( .A1(DP_OP_422J2_124_3477_n2355), 
        .A2(DP_OP_424J2_126_3477_n2365), .Y(DP_OP_422J2_124_3477_n2347) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1568 ( .A1(DP_OP_425J2_127_3477_n2493), .A2(
        DP_OP_422J2_124_3477_n2362), .Y(DP_OP_422J2_124_3477_n2329) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1567 ( .A1(DP_OP_423J2_125_3477_n2668), .A2(
        DP_OP_422J2_124_3477_n2362), .Y(DP_OP_422J2_124_3477_n2328) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1566 ( .A1(DP_OP_424J2_126_3477_n2579), .A2(
        DP_OP_422J2_124_3477_n2362), .Y(DP_OP_422J2_124_3477_n2327) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1565 ( .A1(DP_OP_422J2_124_3477_n2358), .A2(
        DP_OP_422J2_124_3477_n2362), .Y(DP_OP_422J2_124_3477_n2326) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1564 ( .A1(DP_OP_422J2_124_3477_n2357), .A2(
        DP_OP_422J2_124_3477_n2362), .Y(DP_OP_422J2_124_3477_n2325) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1563 ( .A1(DP_OP_422J2_124_3477_n2356), .A2(
        DP_OP_422J2_124_3477_n2362), .Y(DP_OP_422J2_124_3477_n2324) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1562 ( .A1(DP_OP_422J2_124_3477_n2355), .A2(
        DP_OP_422J2_124_3477_n2362), .Y(DP_OP_422J2_124_3477_n2323) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1561 ( .A1(DP_OP_422J2_124_3477_n2354), 
        .A2(DP_OP_422J2_124_3477_n2362), .Y(DP_OP_422J2_124_3477_n2322) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1541 ( .A1(DP_OP_422J2_124_3477_n2310), .A2(
        DP_OP_422J2_124_3477_n2321), .Y(DP_OP_422J2_124_3477_n2302) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1524 ( .A1(DP_OP_425J2_127_3477_n2449), .A2(
        DP_OP_422J2_124_3477_n2318), .Y(DP_OP_422J2_124_3477_n2285) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1523 ( .A1(DP_OP_425J2_127_3477_n2448), .A2(
        DP_OP_422J2_124_3477_n2318), .Y(DP_OP_422J2_124_3477_n2284) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1522 ( .A1(DP_OP_424J2_126_3477_n2623), .A2(
        DP_OP_422J2_124_3477_n2318), .Y(DP_OP_422J2_124_3477_n2283) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1521 ( .A1(DP_OP_422J2_124_3477_n2314), .A2(
        DP_OP_422J2_124_3477_n2318), .Y(DP_OP_422J2_124_3477_n2282) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1520 ( .A1(DP_OP_422J2_124_3477_n2313), .A2(
        DP_OP_422J2_124_3477_n2318), .Y(DP_OP_422J2_124_3477_n2281) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1519 ( .A1(DP_OP_422J2_124_3477_n2312), .A2(
        DP_OP_422J2_124_3477_n2318), .Y(DP_OP_422J2_124_3477_n2280) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1518 ( .A1(DP_OP_422J2_124_3477_n2311), .A2(
        DP_OP_422J2_124_3477_n2318), .Y(DP_OP_422J2_124_3477_n2279) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1517 ( .A1(DP_OP_422J2_124_3477_n2310), 
        .A2(DP_OP_422J2_124_3477_n2318), .Y(DP_OP_422J2_124_3477_n2278) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1497 ( .A1(DP_OP_422J2_124_3477_n2266), .A2(
        DP_OP_422J2_124_3477_n2277), .Y(DP_OP_422J2_124_3477_n2258) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1489 ( .A1(DP_OP_422J2_124_3477_n2266), .A2(
        DP_OP_422J2_124_3477_n2276), .Y(DP_OP_422J2_124_3477_n2250) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1481 ( .A1(DP_OP_422J2_124_3477_n2266), .A2(
        n1427), .Y(DP_OP_422J2_124_3477_n2242) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1480 ( .A1(DP_OP_424J2_126_3477_n2669), .A2(
        n1370), .Y(DP_OP_422J2_124_3477_n2241) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1479 ( .A1(DP_OP_425J2_127_3477_n2404), .A2(
        n1338), .Y(DP_OP_422J2_124_3477_n2240) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1478 ( .A1(DP_OP_425J2_127_3477_n2403), .A2(
        n1338), .Y(DP_OP_422J2_124_3477_n2239) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1477 ( .A1(DP_OP_422J2_124_3477_n2270), .A2(
        n1338), .Y(DP_OP_422J2_124_3477_n2238) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1476 ( .A1(DP_OP_422J2_124_3477_n2269), .A2(
        DP_OP_424J2_126_3477_n2274), .Y(DP_OP_422J2_124_3477_n2237) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1475 ( .A1(DP_OP_422J2_124_3477_n2268), .A2(
        n1338), .Y(DP_OP_422J2_124_3477_n2236) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1474 ( .A1(DP_OP_422J2_124_3477_n2267), .A2(
        n1370), .Y(DP_OP_422J2_124_3477_n2235) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1473 ( .A1(DP_OP_422J2_124_3477_n2266), 
        .A2(DP_OP_424J2_126_3477_n2274), .Y(DP_OP_422J2_124_3477_n2234) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1445 ( .A1(DP_OP_422J2_124_3477_n2222), .A2(
        n365), .Y(DP_OP_422J2_124_3477_n2206) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1432 ( .A1(DP_OP_422J2_124_3477_n2225), .A2(
        DP_OP_423J2_125_3477_n2230), .Y(DP_OP_422J2_124_3477_n2193) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1409 ( .A1(DP_OP_422J2_124_3477_n2178), .A2(
        DP_OP_422J2_124_3477_n2189), .Y(DP_OP_422J2_124_3477_n2170) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1401 ( .A1(DP_OP_422J2_124_3477_n2178), .A2(
        n1344), .Y(DP_OP_422J2_124_3477_n2162) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1394 ( .A1(DP_OP_422J2_124_3477_n2179), 
        .A2(n1339), .Y(DP_OP_422J2_124_3477_n2155) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1393 ( .A1(DP_OP_422J2_124_3477_n2178), .A2(
        n1339), .Y(DP_OP_422J2_124_3477_n2154) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1392 ( .A1(DP_OP_422J2_124_3477_n2185), .A2(
        DP_OP_422J2_124_3477_n2186), .Y(DP_OP_422J2_124_3477_n2153) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1391 ( .A1(DP_OP_424J2_126_3477_n2756), .A2(
        DP_OP_425J2_127_3477_n2186), .Y(DP_OP_422J2_124_3477_n2152) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1390 ( .A1(DP_OP_422J2_124_3477_n2183), .A2(
        DP_OP_424J2_126_3477_n2186), .Y(DP_OP_422J2_124_3477_n2151) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1389 ( .A1(DP_OP_424J2_126_3477_n2754), .A2(
        DP_OP_422J2_124_3477_n2186), .Y(DP_OP_422J2_124_3477_n2150) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1388 ( .A1(DP_OP_422J2_124_3477_n2181), .A2(
        DP_OP_425J2_127_3477_n2186), .Y(DP_OP_422J2_124_3477_n2149) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1387 ( .A1(DP_OP_424J2_126_3477_n2752), .A2(
        DP_OP_425J2_127_3477_n2186), .Y(DP_OP_422J2_124_3477_n2148) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1386 ( .A1(DP_OP_422J2_124_3477_n2179), .A2(
        DP_OP_422J2_124_3477_n2186), .Y(DP_OP_422J2_124_3477_n2147) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1385 ( .A1(DP_OP_422J2_124_3477_n2178), 
        .A2(DP_OP_425J2_127_3477_n2186), .Y(DP_OP_422J2_124_3477_n2146) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1365 ( .A1(DP_OP_422J2_124_3477_n2134), .A2(
        n1500), .Y(DP_OP_422J2_124_3477_n2126) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1358 ( .A1(DP_OP_422J2_124_3477_n2135), 
        .A2(DP_OP_424J2_126_3477_n2144), .Y(DP_OP_422J2_124_3477_n2119) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1357 ( .A1(DP_OP_422J2_124_3477_n2134), .A2(
        DP_OP_422J2_124_3477_n2144), .Y(DP_OP_422J2_124_3477_n2118) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1350 ( .A1(DP_OP_422J2_124_3477_n2135), 
        .A2(DP_OP_422J2_124_3477_n2143), .Y(DP_OP_422J2_124_3477_n2111) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1349 ( .A1(DP_OP_422J2_124_3477_n2134), .A2(
        DP_OP_422J2_124_3477_n2143), .Y(DP_OP_422J2_124_3477_n2110) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1348 ( .A1(DP_OP_423J2_125_3477_n2889), .A2(
        DP_OP_422J2_124_3477_n2142), .Y(DP_OP_422J2_124_3477_n2109) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1347 ( .A1(DP_OP_422J2_124_3477_n2140), .A2(
        DP_OP_422J2_124_3477_n2142), .Y(DP_OP_422J2_124_3477_n2108) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1346 ( .A1(DP_OP_424J2_126_3477_n2799), .A2(
        DP_OP_422J2_124_3477_n2142), .Y(DP_OP_422J2_124_3477_n2107) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1345 ( .A1(DP_OP_422J2_124_3477_n2138), .A2(
        DP_OP_422J2_124_3477_n2142), .Y(DP_OP_422J2_124_3477_n2106) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1344 ( .A1(DP_OP_422J2_124_3477_n2137), .A2(
        DP_OP_422J2_124_3477_n2142), .Y(DP_OP_422J2_124_3477_n2105) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1343 ( .A1(DP_OP_425J2_127_3477_n2268), .A2(
        DP_OP_422J2_124_3477_n2142), .Y(DP_OP_422J2_124_3477_n2104) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1342 ( .A1(DP_OP_422J2_124_3477_n2135), .A2(
        DP_OP_422J2_124_3477_n2142), .Y(DP_OP_422J2_124_3477_n2103) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1341 ( .A1(DP_OP_422J2_124_3477_n2134), 
        .A2(DP_OP_422J2_124_3477_n2142), .Y(DP_OP_422J2_124_3477_n2102) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1314 ( .A1(DP_OP_422J2_124_3477_n2091), 
        .A2(DP_OP_423J2_125_3477_n2100), .Y(DP_OP_422J2_124_3477_n2075) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1313 ( .A1(DP_OP_422J2_124_3477_n2090), .A2(
        DP_OP_422J2_124_3477_n2100), .Y(DP_OP_422J2_124_3477_n2074) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1306 ( .A1(DP_OP_422J2_124_3477_n2091), 
        .A2(DP_OP_424J2_126_3477_n2099), .Y(DP_OP_422J2_124_3477_n2067) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1305 ( .A1(DP_OP_422J2_124_3477_n2090), .A2(
        DP_OP_424J2_126_3477_n2099), .Y(DP_OP_422J2_124_3477_n2066) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1303 ( .A1(DP_OP_423J2_125_3477_n2932), .A2(
        DP_OP_423J2_125_3477_n2098), .Y(DP_OP_422J2_124_3477_n2064) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1301 ( .A1(DP_OP_425J2_127_3477_n2226), .A2(
        DP_OP_423J2_125_3477_n2098), .Y(DP_OP_422J2_124_3477_n2062) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1278 ( .A1(DP_OP_422J2_124_3477_n2047), 
        .A2(n1475), .Y(DP_OP_422J2_124_3477_n2039) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1277 ( .A1(DP_OP_422J2_124_3477_n2046), .A2(
        n1475), .Y(DP_OP_422J2_124_3477_n2038) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1269 ( .A1(DP_OP_422J2_124_3477_n2046), .A2(
        DP_OP_422J2_124_3477_n2056), .Y(DP_OP_422J2_124_3477_n2030) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1261 ( .A1(DP_OP_422J2_124_3477_n2046), .A2(
        DP_OP_422J2_124_3477_n2055), .Y(DP_OP_422J2_124_3477_n2022) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1259 ( .A1(DP_OP_425J2_127_3477_n2184), .A2(
        n30), .Y(DP_OP_422J2_124_3477_n2020) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1257 ( .A1(DP_OP_424J2_126_3477_n2886), .A2(
        n30), .Y(DP_OP_422J2_124_3477_n2018) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1255 ( .A1(DP_OP_422J2_124_3477_n2048), .A2(
        n30), .Y(DP_OP_422J2_124_3477_n2016) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1254 ( .A1(DP_OP_422J2_124_3477_n2047), .A2(
        n30), .Y(DP_OP_422J2_124_3477_n2015) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1233 ( .A1(DP_OP_422J2_124_3477_n2002), .A2(
        n1431), .Y(DP_OP_422J2_124_3477_n1994) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1226 ( .A1(DP_OP_422J2_124_3477_n2003), 
        .A2(n558), .Y(DP_OP_422J2_124_3477_n1987) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1225 ( .A1(DP_OP_422J2_124_3477_n2002), .A2(
        n558), .Y(DP_OP_422J2_124_3477_n1986) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1217 ( .A1(DP_OP_422J2_124_3477_n2002), .A2(
        DP_OP_422J2_124_3477_n2011), .Y(DP_OP_422J2_124_3477_n1978) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1216 ( .A1(DP_OP_424J2_126_3477_n2933), .A2(
        DP_OP_425J2_127_3477_n2010), .Y(DP_OP_422J2_124_3477_n1977) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1215 ( .A1(DP_OP_424J2_126_3477_n2932), .A2(
        DP_OP_424J2_126_3477_n2010), .Y(DP_OP_422J2_124_3477_n1976) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1214 ( .A1(DP_OP_422J2_124_3477_n2007), .A2(
        DP_OP_425J2_127_3477_n2010), .Y(DP_OP_422J2_124_3477_n1975) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1212 ( .A1(DP_OP_422J2_124_3477_n2005), .A2(
        DP_OP_423J2_125_3477_n2010), .Y(DP_OP_422J2_124_3477_n1973) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1211 ( .A1(DP_OP_422J2_124_3477_n2004), .A2(
        DP_OP_424J2_126_3477_n2010), .Y(DP_OP_422J2_124_3477_n1972) );
  OR2X1_HVT DP_OP_422J2_124_3477_U1210 ( .A1(DP_OP_422J2_124_3477_n2003), .A2(
        DP_OP_424J2_126_3477_n2010), .Y(DP_OP_422J2_124_3477_n1971) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1209 ( .A1(DP_OP_422J2_124_3477_n2002), 
        .A2(DP_OP_424J2_126_3477_n2010), .Y(DP_OP_422J2_124_3477_n1970) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1165 ( .A1(n1849), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_422J2_124_3477_n510) );
  HADDX1_HVT DP_OP_422J2_124_3477_U1143 ( .A0(DP_OP_422J2_124_3477_n1936), 
        .B0(DP_OP_422J2_124_3477_n2045), .C1(DP_OP_422J2_124_3477_n1920), .SO(
        DP_OP_422J2_124_3477_n1921) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1142 ( .A(DP_OP_422J2_124_3477_n2089), .B(
        DP_OP_422J2_124_3477_n2001), .CI(DP_OP_422J2_124_3477_n2133), .CO(
        DP_OP_422J2_124_3477_n1918), .S(DP_OP_422J2_124_3477_n1919) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1141 ( .A(DP_OP_422J2_124_3477_n2221), .B(
        DP_OP_422J2_124_3477_n2177), .CI(DP_OP_422J2_124_3477_n2265), .CO(
        DP_OP_422J2_124_3477_n1916), .S(DP_OP_422J2_124_3477_n1917) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1140 ( .A(DP_OP_422J2_124_3477_n2353), .B(
        DP_OP_422J2_124_3477_n2309), .CI(DP_OP_422J2_124_3477_n2397), .CO(
        DP_OP_422J2_124_3477_n1914), .S(DP_OP_422J2_124_3477_n1915) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1139 ( .A(DP_OP_422J2_124_3477_n2485), .B(
        DP_OP_422J2_124_3477_n2441), .CI(DP_OP_422J2_124_3477_n2529), .CO(
        DP_OP_422J2_124_3477_n1912), .S(DP_OP_422J2_124_3477_n1913) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1138 ( .A(DP_OP_422J2_124_3477_n2617), .B(
        DP_OP_422J2_124_3477_n2573), .CI(DP_OP_422J2_124_3477_n2661), .CO(
        DP_OP_422J2_124_3477_n1910), .S(DP_OP_422J2_124_3477_n1911) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1137 ( .A(DP_OP_422J2_124_3477_n2749), .B(
        DP_OP_422J2_124_3477_n2705), .CI(DP_OP_422J2_124_3477_n2793), .CO(
        DP_OP_422J2_124_3477_n1908), .S(DP_OP_422J2_124_3477_n1909) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1136 ( .A(DP_OP_422J2_124_3477_n3055), .B(
        DP_OP_422J2_124_3477_n2837), .CI(DP_OP_422J2_124_3477_n2881), .CO(
        DP_OP_422J2_124_3477_n1906), .S(DP_OP_422J2_124_3477_n1907) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1135 ( .A(DP_OP_422J2_124_3477_n3013), .B(
        DP_OP_422J2_124_3477_n2925), .CI(DP_OP_422J2_124_3477_n2969), .CO(
        DP_OP_422J2_124_3477_n1904), .S(DP_OP_422J2_124_3477_n1905) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1134 ( .A(DP_OP_422J2_124_3477_n1921), .B(
        DP_OP_422J2_124_3477_n1907), .CI(DP_OP_422J2_124_3477_n1909), .CO(
        DP_OP_422J2_124_3477_n1902), .S(DP_OP_422J2_124_3477_n1903) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1133 ( .A(DP_OP_422J2_124_3477_n1911), .B(
        DP_OP_422J2_124_3477_n1905), .CI(DP_OP_422J2_124_3477_n1913), .CO(
        DP_OP_422J2_124_3477_n1900), .S(DP_OP_422J2_124_3477_n1901) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1132 ( .A(DP_OP_422J2_124_3477_n1919), .B(
        DP_OP_422J2_124_3477_n1915), .CI(DP_OP_422J2_124_3477_n1917), .CO(
        DP_OP_422J2_124_3477_n1898), .S(DP_OP_422J2_124_3477_n1899) );
  HADDX1_HVT DP_OP_422J2_124_3477_U1131 ( .A0(DP_OP_422J2_124_3477_n1935), 
        .B0(DP_OP_422J2_124_3477_n2000), .C1(DP_OP_422J2_124_3477_n1896), .SO(
        DP_OP_422J2_124_3477_n1897) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1130 ( .A(DP_OP_422J2_124_3477_n2037), .B(
        DP_OP_422J2_124_3477_n1993), .CI(DP_OP_422J2_124_3477_n2044), .CO(
        DP_OP_422J2_124_3477_n1894), .S(DP_OP_422J2_124_3477_n1895) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1129 ( .A(DP_OP_422J2_124_3477_n2088), .B(
        DP_OP_422J2_124_3477_n2081), .CI(DP_OP_422J2_124_3477_n2125), .CO(
        DP_OP_422J2_124_3477_n1892), .S(DP_OP_422J2_124_3477_n1893) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1128 ( .A(DP_OP_422J2_124_3477_n2169), .B(
        DP_OP_422J2_124_3477_n2132), .CI(DP_OP_422J2_124_3477_n2176), .CO(
        DP_OP_422J2_124_3477_n1890), .S(DP_OP_422J2_124_3477_n1891) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1127 ( .A(DP_OP_422J2_124_3477_n2220), .B(
        DP_OP_422J2_124_3477_n2213), .CI(DP_OP_422J2_124_3477_n2257), .CO(
        DP_OP_422J2_124_3477_n1888), .S(DP_OP_422J2_124_3477_n1889) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1126 ( .A(DP_OP_422J2_124_3477_n2301), .B(
        DP_OP_422J2_124_3477_n2264), .CI(DP_OP_422J2_124_3477_n2308), .CO(
        DP_OP_422J2_124_3477_n1886), .S(DP_OP_422J2_124_3477_n1887) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1125 ( .A(DP_OP_422J2_124_3477_n2352), .B(
        DP_OP_422J2_124_3477_n2345), .CI(DP_OP_422J2_124_3477_n2389), .CO(
        DP_OP_422J2_124_3477_n1884), .S(DP_OP_422J2_124_3477_n1885) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1124 ( .A(DP_OP_422J2_124_3477_n2433), .B(
        DP_OP_422J2_124_3477_n2396), .CI(DP_OP_422J2_124_3477_n2440), .CO(
        DP_OP_422J2_124_3477_n1882), .S(DP_OP_422J2_124_3477_n1883) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1123 ( .A(DP_OP_422J2_124_3477_n2484), .B(
        DP_OP_422J2_124_3477_n2477), .CI(DP_OP_422J2_124_3477_n2521), .CO(
        DP_OP_422J2_124_3477_n1880), .S(DP_OP_422J2_124_3477_n1881) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1122 ( .A(DP_OP_422J2_124_3477_n2565), .B(
        DP_OP_422J2_124_3477_n2528), .CI(DP_OP_422J2_124_3477_n2572), .CO(
        DP_OP_422J2_124_3477_n1878), .S(DP_OP_422J2_124_3477_n1879) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1121 ( .A(DP_OP_422J2_124_3477_n3054), .B(
        DP_OP_422J2_124_3477_n2609), .CI(DP_OP_422J2_124_3477_n3047), .CO(
        DP_OP_422J2_124_3477_n1876), .S(DP_OP_422J2_124_3477_n1877) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1120 ( .A(DP_OP_422J2_124_3477_n2792), .B(
        DP_OP_422J2_124_3477_n2616), .CI(DP_OP_422J2_124_3477_n2653), .CO(
        DP_OP_422J2_124_3477_n1874), .S(DP_OP_422J2_124_3477_n1875) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1119 ( .A(DP_OP_422J2_124_3477_n2829), .B(
        DP_OP_422J2_124_3477_n3012), .CI(DP_OP_422J2_124_3477_n3005), .CO(
        DP_OP_422J2_124_3477_n1872), .S(DP_OP_422J2_124_3477_n1873) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1118 ( .A(DP_OP_422J2_124_3477_n2748), .B(
        DP_OP_422J2_124_3477_n2968), .CI(DP_OP_422J2_124_3477_n2961), .CO(
        DP_OP_422J2_124_3477_n1870), .S(DP_OP_422J2_124_3477_n1871) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1117 ( .A(DP_OP_422J2_124_3477_n2741), .B(
        DP_OP_422J2_124_3477_n2924), .CI(DP_OP_422J2_124_3477_n2660), .CO(
        DP_OP_422J2_124_3477_n1868), .S(DP_OP_422J2_124_3477_n1869) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1116 ( .A(DP_OP_422J2_124_3477_n2917), .B(
        DP_OP_422J2_124_3477_n2697), .CI(DP_OP_422J2_124_3477_n2704), .CO(
        DP_OP_422J2_124_3477_n1866), .S(DP_OP_422J2_124_3477_n1867) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1115 ( .A(DP_OP_422J2_124_3477_n2873), .B(
        DP_OP_422J2_124_3477_n2785), .CI(DP_OP_422J2_124_3477_n2836), .CO(
        DP_OP_422J2_124_3477_n1864), .S(DP_OP_422J2_124_3477_n1865) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1114 ( .A(DP_OP_422J2_124_3477_n2880), .B(
        DP_OP_422J2_124_3477_n1920), .CI(DP_OP_422J2_124_3477_n1897), .CO(
        DP_OP_422J2_124_3477_n1862), .S(DP_OP_422J2_124_3477_n1863) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1113 ( .A(DP_OP_422J2_124_3477_n1904), .B(
        DP_OP_422J2_124_3477_n1918), .CI(DP_OP_422J2_124_3477_n1916), .CO(
        DP_OP_422J2_124_3477_n1860), .S(DP_OP_422J2_124_3477_n1861) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1112 ( .A(DP_OP_422J2_124_3477_n1910), .B(
        DP_OP_422J2_124_3477_n1906), .CI(DP_OP_422J2_124_3477_n1914), .CO(
        DP_OP_422J2_124_3477_n1858), .S(DP_OP_422J2_124_3477_n1859) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1111 ( .A(DP_OP_422J2_124_3477_n1912), .B(
        DP_OP_422J2_124_3477_n1908), .CI(DP_OP_422J2_124_3477_n1865), .CO(
        DP_OP_422J2_124_3477_n1856), .S(DP_OP_422J2_124_3477_n1857) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1110 ( .A(DP_OP_422J2_124_3477_n1887), .B(
        DP_OP_422J2_124_3477_n1873), .CI(DP_OP_422J2_124_3477_n1871), .CO(
        DP_OP_422J2_124_3477_n1854), .S(DP_OP_422J2_124_3477_n1855) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1109 ( .A(DP_OP_422J2_124_3477_n1891), .B(
        DP_OP_422J2_124_3477_n1875), .CI(DP_OP_422J2_124_3477_n1879), .CO(
        DP_OP_422J2_124_3477_n1852), .S(DP_OP_422J2_124_3477_n1853) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1108 ( .A(DP_OP_422J2_124_3477_n1893), .B(
        DP_OP_422J2_124_3477_n1881), .CI(DP_OP_422J2_124_3477_n1877), .CO(
        DP_OP_422J2_124_3477_n1850), .S(DP_OP_422J2_124_3477_n1851) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1107 ( .A(DP_OP_422J2_124_3477_n1895), .B(
        DP_OP_422J2_124_3477_n1885), .CI(DP_OP_422J2_124_3477_n1869), .CO(
        DP_OP_422J2_124_3477_n1848), .S(DP_OP_422J2_124_3477_n1849) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1106 ( .A(DP_OP_422J2_124_3477_n1889), .B(
        DP_OP_422J2_124_3477_n1883), .CI(DP_OP_422J2_124_3477_n1867), .CO(
        DP_OP_422J2_124_3477_n1846), .S(DP_OP_422J2_124_3477_n1847) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1105 ( .A(DP_OP_422J2_124_3477_n1863), .B(
        DP_OP_422J2_124_3477_n1902), .CI(DP_OP_422J2_124_3477_n1900), .CO(
        DP_OP_422J2_124_3477_n1844), .S(DP_OP_422J2_124_3477_n1845) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1104 ( .A(DP_OP_422J2_124_3477_n1898), .B(
        DP_OP_422J2_124_3477_n1859), .CI(DP_OP_422J2_124_3477_n1861), .CO(
        DP_OP_422J2_124_3477_n1842), .S(DP_OP_422J2_124_3477_n1843) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1103 ( .A(DP_OP_422J2_124_3477_n1857), .B(
        DP_OP_422J2_124_3477_n1849), .CI(DP_OP_422J2_124_3477_n1851), .CO(
        DP_OP_422J2_124_3477_n1840), .S(DP_OP_422J2_124_3477_n1841) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1102 ( .A(DP_OP_422J2_124_3477_n1855), .B(
        DP_OP_422J2_124_3477_n1847), .CI(DP_OP_422J2_124_3477_n1853), .CO(
        DP_OP_422J2_124_3477_n1838), .S(DP_OP_422J2_124_3477_n1839) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1101 ( .A(DP_OP_422J2_124_3477_n1845), .B(
        DP_OP_422J2_124_3477_n1843), .CI(DP_OP_422J2_124_3477_n1841), .CO(
        DP_OP_422J2_124_3477_n1836), .S(DP_OP_422J2_124_3477_n1837) );
  HADDX1_HVT DP_OP_422J2_124_3477_U1100 ( .A0(DP_OP_422J2_124_3477_n1934), 
        .B0(DP_OP_422J2_124_3477_n1999), .C1(DP_OP_422J2_124_3477_n1834), .SO(
        DP_OP_422J2_124_3477_n1835) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1099 ( .A(DP_OP_422J2_124_3477_n2029), .B(
        DP_OP_422J2_124_3477_n1992), .CI(DP_OP_422J2_124_3477_n1985), .CO(
        DP_OP_422J2_124_3477_n1832), .S(DP_OP_422J2_124_3477_n1833) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1098 ( .A(DP_OP_422J2_124_3477_n2043), .B(
        DP_OP_422J2_124_3477_n2036), .CI(DP_OP_422J2_124_3477_n2073), .CO(
        DP_OP_422J2_124_3477_n1830), .S(DP_OP_422J2_124_3477_n1831) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1097 ( .A(DP_OP_422J2_124_3477_n2087), .B(
        DP_OP_422J2_124_3477_n2080), .CI(DP_OP_422J2_124_3477_n2117), .CO(
        DP_OP_422J2_124_3477_n1828), .S(DP_OP_422J2_124_3477_n1829) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1096 ( .A(DP_OP_422J2_124_3477_n2131), .B(
        DP_OP_422J2_124_3477_n2124), .CI(DP_OP_422J2_124_3477_n2161), .CO(
        DP_OP_422J2_124_3477_n1826), .S(DP_OP_422J2_124_3477_n1827) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1095 ( .A(DP_OP_422J2_124_3477_n2175), .B(
        DP_OP_422J2_124_3477_n2168), .CI(DP_OP_422J2_124_3477_n2205), .CO(
        DP_OP_422J2_124_3477_n1824), .S(DP_OP_422J2_124_3477_n1825) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1094 ( .A(DP_OP_422J2_124_3477_n2219), .B(
        DP_OP_422J2_124_3477_n2212), .CI(DP_OP_422J2_124_3477_n2249), .CO(
        DP_OP_422J2_124_3477_n1822), .S(DP_OP_422J2_124_3477_n1823) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1093 ( .A(DP_OP_422J2_124_3477_n2263), .B(
        DP_OP_422J2_124_3477_n2256), .CI(DP_OP_422J2_124_3477_n2293), .CO(
        DP_OP_422J2_124_3477_n1820), .S(DP_OP_422J2_124_3477_n1821) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1092 ( .A(DP_OP_422J2_124_3477_n2307), .B(
        DP_OP_422J2_124_3477_n2300), .CI(DP_OP_422J2_124_3477_n2337), .CO(
        DP_OP_422J2_124_3477_n1818), .S(DP_OP_422J2_124_3477_n1819) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1091 ( .A(DP_OP_422J2_124_3477_n2351), .B(
        DP_OP_422J2_124_3477_n2344), .CI(DP_OP_422J2_124_3477_n2381), .CO(
        DP_OP_422J2_124_3477_n1816), .S(DP_OP_422J2_124_3477_n1817) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1090 ( .A(DP_OP_422J2_124_3477_n2395), .B(
        DP_OP_422J2_124_3477_n2388), .CI(DP_OP_422J2_124_3477_n2425), .CO(
        DP_OP_422J2_124_3477_n1814), .S(DP_OP_422J2_124_3477_n1815) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1089 ( .A(DP_OP_422J2_124_3477_n2439), .B(
        DP_OP_422J2_124_3477_n2432), .CI(DP_OP_422J2_124_3477_n2469), .CO(
        DP_OP_422J2_124_3477_n1812), .S(DP_OP_422J2_124_3477_n1813) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1088 ( .A(DP_OP_422J2_124_3477_n2740), .B(
        DP_OP_422J2_124_3477_n3053), .CI(DP_OP_422J2_124_3477_n3046), .CO(
        DP_OP_422J2_124_3477_n1810), .S(DP_OP_422J2_124_3477_n1811) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1087 ( .A(DP_OP_422J2_124_3477_n2703), .B(
        DP_OP_422J2_124_3477_n2476), .CI(DP_OP_422J2_124_3477_n3039), .CO(
        DP_OP_422J2_124_3477_n1808), .S(DP_OP_422J2_124_3477_n1809) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1086 ( .A(DP_OP_422J2_124_3477_n2696), .B(
        DP_OP_422J2_124_3477_n3011), .CI(DP_OP_422J2_124_3477_n2483), .CO(
        DP_OP_422J2_124_3477_n1806), .S(DP_OP_422J2_124_3477_n1807) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1085 ( .A(DP_OP_422J2_124_3477_n2733), .B(
        DP_OP_422J2_124_3477_n2513), .CI(DP_OP_422J2_124_3477_n2520), .CO(
        DP_OP_422J2_124_3477_n1804), .S(DP_OP_422J2_124_3477_n1805) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1084 ( .A(DP_OP_422J2_124_3477_n2747), .B(
        DP_OP_422J2_124_3477_n2527), .CI(DP_OP_422J2_124_3477_n3004), .CO(
        DP_OP_422J2_124_3477_n1802), .S(DP_OP_422J2_124_3477_n1803) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1083 ( .A(DP_OP_422J2_124_3477_n2777), .B(
        DP_OP_422J2_124_3477_n2557), .CI(DP_OP_422J2_124_3477_n2997), .CO(
        DP_OP_422J2_124_3477_n1800), .S(DP_OP_422J2_124_3477_n1801) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1082 ( .A(DP_OP_422J2_124_3477_n2689), .B(
        DP_OP_422J2_124_3477_n2564), .CI(DP_OP_422J2_124_3477_n2967), .CO(
        DP_OP_422J2_124_3477_n1798), .S(DP_OP_422J2_124_3477_n1799) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1081 ( .A(DP_OP_422J2_124_3477_n2659), .B(
        DP_OP_422J2_124_3477_n2571), .CI(DP_OP_422J2_124_3477_n2960), .CO(
        DP_OP_422J2_124_3477_n1796), .S(DP_OP_422J2_124_3477_n1797) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1080 ( .A(DP_OP_422J2_124_3477_n2953), .B(
        DP_OP_422J2_124_3477_n2601), .CI(DP_OP_422J2_124_3477_n2608), .CO(
        DP_OP_422J2_124_3477_n1794), .S(DP_OP_422J2_124_3477_n1795) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1079 ( .A(DP_OP_422J2_124_3477_n2923), .B(
        DP_OP_422J2_124_3477_n2615), .CI(DP_OP_422J2_124_3477_n2645), .CO(
        DP_OP_422J2_124_3477_n1792), .S(DP_OP_422J2_124_3477_n1793) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1078 ( .A(DP_OP_422J2_124_3477_n2916), .B(
        DP_OP_422J2_124_3477_n2652), .CI(DP_OP_422J2_124_3477_n2784), .CO(
        DP_OP_422J2_124_3477_n1790), .S(DP_OP_422J2_124_3477_n1791) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1077 ( .A(DP_OP_422J2_124_3477_n2909), .B(
        DP_OP_422J2_124_3477_n2791), .CI(DP_OP_422J2_124_3477_n2821), .CO(
        DP_OP_422J2_124_3477_n1788), .S(DP_OP_422J2_124_3477_n1789) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1076 ( .A(DP_OP_422J2_124_3477_n2879), .B(
        DP_OP_422J2_124_3477_n2828), .CI(DP_OP_422J2_124_3477_n2835), .CO(
        DP_OP_422J2_124_3477_n1786), .S(DP_OP_422J2_124_3477_n1787) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1075 ( .A(DP_OP_422J2_124_3477_n2872), .B(
        DP_OP_422J2_124_3477_n2865), .CI(DP_OP_422J2_124_3477_n1896), .CO(
        DP_OP_422J2_124_3477_n1784), .S(DP_OP_422J2_124_3477_n1785) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1074 ( .A(DP_OP_422J2_124_3477_n1835), .B(
        DP_OP_422J2_124_3477_n1864), .CI(DP_OP_422J2_124_3477_n1866), .CO(
        DP_OP_422J2_124_3477_n1782), .S(DP_OP_422J2_124_3477_n1783) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1073 ( .A(DP_OP_422J2_124_3477_n1882), .B(
        DP_OP_422J2_124_3477_n1894), .CI(DP_OP_422J2_124_3477_n1868), .CO(
        DP_OP_422J2_124_3477_n1780), .S(DP_OP_422J2_124_3477_n1781) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1072 ( .A(DP_OP_422J2_124_3477_n1880), .B(
        DP_OP_422J2_124_3477_n1892), .CI(DP_OP_422J2_124_3477_n1870), .CO(
        DP_OP_422J2_124_3477_n1778), .S(DP_OP_422J2_124_3477_n1779) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1071 ( .A(DP_OP_422J2_124_3477_n1876), .B(
        DP_OP_422J2_124_3477_n1890), .CI(DP_OP_422J2_124_3477_n1872), .CO(
        DP_OP_422J2_124_3477_n1776), .S(DP_OP_422J2_124_3477_n1777) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1070 ( .A(DP_OP_422J2_124_3477_n1888), .B(
        DP_OP_422J2_124_3477_n1886), .CI(DP_OP_422J2_124_3477_n1884), .CO(
        DP_OP_422J2_124_3477_n1774), .S(DP_OP_422J2_124_3477_n1775) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1068 ( .A(DP_OP_422J2_124_3477_n1801), .B(
        DP_OP_422J2_124_3477_n1815), .CI(DP_OP_422J2_124_3477_n1819), .CO(
        DP_OP_422J2_124_3477_n1770), .S(DP_OP_422J2_124_3477_n1771) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1067 ( .A(DP_OP_422J2_124_3477_n1797), .B(
        DP_OP_422J2_124_3477_n1825), .CI(DP_OP_422J2_124_3477_n1827), .CO(
        DP_OP_422J2_124_3477_n1768), .S(DP_OP_422J2_124_3477_n1769) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1066 ( .A(DP_OP_422J2_124_3477_n1795), .B(
        DP_OP_422J2_124_3477_n1817), .CI(DP_OP_422J2_124_3477_n1831), .CO(
        DP_OP_422J2_124_3477_n1766), .S(DP_OP_422J2_124_3477_n1767) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1065 ( .A(DP_OP_422J2_124_3477_n1793), .B(
        DP_OP_422J2_124_3477_n1811), .CI(DP_OP_422J2_124_3477_n1829), .CO(
        DP_OP_422J2_124_3477_n1764), .S(DP_OP_422J2_124_3477_n1765) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1064 ( .A(DP_OP_422J2_124_3477_n1791), .B(
        DP_OP_422J2_124_3477_n1821), .CI(DP_OP_422J2_124_3477_n1809), .CO(
        DP_OP_422J2_124_3477_n1762), .S(DP_OP_422J2_124_3477_n1763) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1063 ( .A(DP_OP_422J2_124_3477_n1789), .B(
        DP_OP_422J2_124_3477_n1823), .CI(DP_OP_422J2_124_3477_n1833), .CO(
        DP_OP_422J2_124_3477_n1760), .S(DP_OP_422J2_124_3477_n1761) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1062 ( .A(DP_OP_422J2_124_3477_n1787), .B(
        DP_OP_422J2_124_3477_n1813), .CI(DP_OP_422J2_124_3477_n1799), .CO(
        DP_OP_422J2_124_3477_n1758), .S(DP_OP_422J2_124_3477_n1759) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1061 ( .A(DP_OP_422J2_124_3477_n1805), .B(
        DP_OP_422J2_124_3477_n1803), .CI(DP_OP_422J2_124_3477_n1862), .CO(
        DP_OP_422J2_124_3477_n1756), .S(DP_OP_422J2_124_3477_n1757) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1060 ( .A(DP_OP_422J2_124_3477_n1785), .B(
        DP_OP_422J2_124_3477_n1860), .CI(DP_OP_422J2_124_3477_n1858), .CO(
        DP_OP_422J2_124_3477_n1754), .S(DP_OP_422J2_124_3477_n1755) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1059 ( .A(DP_OP_422J2_124_3477_n1856), .B(
        DP_OP_422J2_124_3477_n1783), .CI(DP_OP_422J2_124_3477_n1850), .CO(
        DP_OP_422J2_124_3477_n1752), .S(DP_OP_422J2_124_3477_n1753) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1058 ( .A(DP_OP_422J2_124_3477_n1854), .B(
        DP_OP_422J2_124_3477_n1775), .CI(DP_OP_422J2_124_3477_n1781), .CO(
        DP_OP_422J2_124_3477_n1750), .S(DP_OP_422J2_124_3477_n1751) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1057 ( .A(DP_OP_422J2_124_3477_n1852), .B(
        DP_OP_422J2_124_3477_n1779), .CI(DP_OP_422J2_124_3477_n1777), .CO(
        DP_OP_422J2_124_3477_n1748), .S(DP_OP_422J2_124_3477_n1749) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1056 ( .A(DP_OP_422J2_124_3477_n1848), .B(
        DP_OP_422J2_124_3477_n1846), .CI(DP_OP_422J2_124_3477_n1773), .CO(
        DP_OP_422J2_124_3477_n1746), .S(DP_OP_422J2_124_3477_n1747) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1055 ( .A(DP_OP_422J2_124_3477_n1771), .B(
        DP_OP_422J2_124_3477_n1759), .CI(DP_OP_422J2_124_3477_n1757), .CO(
        DP_OP_422J2_124_3477_n1744), .S(DP_OP_422J2_124_3477_n1745) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1054 ( .A(DP_OP_422J2_124_3477_n1761), .B(
        DP_OP_422J2_124_3477_n1769), .CI(DP_OP_422J2_124_3477_n1767), .CO(
        DP_OP_422J2_124_3477_n1742), .S(DP_OP_422J2_124_3477_n1743) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1053 ( .A(DP_OP_422J2_124_3477_n1763), .B(
        DP_OP_422J2_124_3477_n1765), .CI(DP_OP_422J2_124_3477_n1844), .CO(
        DP_OP_422J2_124_3477_n1740), .S(DP_OP_422J2_124_3477_n1741) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1052 ( .A(DP_OP_422J2_124_3477_n1755), .B(
        DP_OP_422J2_124_3477_n1842), .CI(DP_OP_422J2_124_3477_n1753), .CO(
        DP_OP_422J2_124_3477_n1738), .S(DP_OP_422J2_124_3477_n1739) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1051 ( .A(DP_OP_422J2_124_3477_n1840), .B(
        DP_OP_422J2_124_3477_n1838), .CI(DP_OP_422J2_124_3477_n1749), .CO(
        DP_OP_422J2_124_3477_n1736), .S(DP_OP_422J2_124_3477_n1737) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1050 ( .A(DP_OP_422J2_124_3477_n1751), .B(
        DP_OP_422J2_124_3477_n1747), .CI(DP_OP_422J2_124_3477_n1745), .CO(
        DP_OP_422J2_124_3477_n1734), .S(DP_OP_422J2_124_3477_n1735) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1049 ( .A(DP_OP_422J2_124_3477_n1743), .B(
        DP_OP_422J2_124_3477_n1741), .CI(DP_OP_422J2_124_3477_n1739), .CO(
        DP_OP_422J2_124_3477_n1732), .S(DP_OP_422J2_124_3477_n1733) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1048 ( .A(DP_OP_422J2_124_3477_n1836), .B(
        DP_OP_422J2_124_3477_n1737), .CI(DP_OP_422J2_124_3477_n1735), .CO(
        DP_OP_422J2_124_3477_n1730), .S(DP_OP_422J2_124_3477_n1731) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1046 ( .A(DP_OP_422J2_124_3477_n2505), .B(
        DP_OP_422J2_124_3477_n1977), .CI(DP_OP_422J2_124_3477_n1933), .CO(
        DP_OP_422J2_124_3477_n1726), .S(DP_OP_422J2_124_3477_n1727) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1045 ( .A(DP_OP_422J2_124_3477_n2197), .B(
        DP_OP_422J2_124_3477_n2637), .CI(DP_OP_422J2_124_3477_n2417), .CO(
        DP_OP_422J2_124_3477_n1724), .S(DP_OP_422J2_124_3477_n1725) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1044 ( .A(DP_OP_422J2_124_3477_n2945), .B(
        DP_OP_422J2_124_3477_n2153), .CI(DP_OP_422J2_124_3477_n2373), .CO(
        DP_OP_422J2_124_3477_n1722), .S(DP_OP_422J2_124_3477_n1723) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1043 ( .A(DP_OP_422J2_124_3477_n2549), .B(
        DP_OP_422J2_124_3477_n2857), .CI(DP_OP_422J2_124_3477_n2461), .CO(
        DP_OP_422J2_124_3477_n1720), .S(DP_OP_422J2_124_3477_n1721) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1042 ( .A(DP_OP_422J2_124_3477_n2285), .B(
        DP_OP_422J2_124_3477_n2329), .CI(DP_OP_422J2_124_3477_n2109), .CO(
        DP_OP_422J2_124_3477_n1718), .S(DP_OP_422J2_124_3477_n1719) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1041 ( .A(DP_OP_422J2_124_3477_n2813), .B(
        DP_OP_422J2_124_3477_n2681), .CI(DP_OP_422J2_124_3477_n2725), .CO(
        DP_OP_422J2_124_3477_n1716), .S(DP_OP_422J2_124_3477_n1717) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1039 ( .A(DP_OP_422J2_124_3477_n2593), .B(
        DP_OP_422J2_124_3477_n2989), .CI(DP_OP_422J2_124_3477_n2241), .CO(
        DP_OP_422J2_124_3477_n1712), .S(DP_OP_422J2_124_3477_n1713) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1038 ( .A(DP_OP_422J2_124_3477_n2021), .B(
        DP_OP_422J2_124_3477_n1729), .CI(DP_OP_422J2_124_3477_n1998), .CO(
        DP_OP_422J2_124_3477_n1710), .S(DP_OP_422J2_124_3477_n1711) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1037 ( .A(DP_OP_422J2_124_3477_n2028), .B(
        DP_OP_422J2_124_3477_n1991), .CI(DP_OP_422J2_124_3477_n1984), .CO(
        DP_OP_422J2_124_3477_n1708), .S(DP_OP_422J2_124_3477_n1709) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1036 ( .A(DP_OP_422J2_124_3477_n2042), .B(
        DP_OP_422J2_124_3477_n2035), .CI(DP_OP_422J2_124_3477_n2072), .CO(
        DP_OP_422J2_124_3477_n1706), .S(DP_OP_422J2_124_3477_n1707) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1035 ( .A(DP_OP_422J2_124_3477_n2086), .B(
        DP_OP_422J2_124_3477_n2079), .CI(DP_OP_422J2_124_3477_n2116), .CO(
        DP_OP_422J2_124_3477_n1704), .S(DP_OP_422J2_124_3477_n1705) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1034 ( .A(DP_OP_422J2_124_3477_n3052), .B(
        DP_OP_422J2_124_3477_n2123), .CI(DP_OP_422J2_124_3477_n2130), .CO(
        DP_OP_422J2_124_3477_n1702), .S(DP_OP_422J2_124_3477_n1703) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1033 ( .A(DP_OP_422J2_124_3477_n2563), .B(
        DP_OP_422J2_124_3477_n3045), .CI(DP_OP_422J2_124_3477_n3038), .CO(
        DP_OP_422J2_124_3477_n1700), .S(DP_OP_422J2_124_3477_n1701) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1032 ( .A(DP_OP_422J2_124_3477_n2526), .B(
        DP_OP_422J2_124_3477_n2160), .CI(DP_OP_422J2_124_3477_n3010), .CO(
        DP_OP_422J2_124_3477_n1698), .S(DP_OP_422J2_124_3477_n1699) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1031 ( .A(DP_OP_422J2_124_3477_n2556), .B(
        DP_OP_422J2_124_3477_n2167), .CI(DP_OP_422J2_124_3477_n3003), .CO(
        DP_OP_422J2_124_3477_n1696), .S(DP_OP_422J2_124_3477_n1697) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1030 ( .A(DP_OP_422J2_124_3477_n2996), .B(
        DP_OP_422J2_124_3477_n2174), .CI(DP_OP_422J2_124_3477_n2204), .CO(
        DP_OP_422J2_124_3477_n1694), .S(DP_OP_422J2_124_3477_n1695) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1029 ( .A(DP_OP_422J2_124_3477_n2519), .B(
        DP_OP_422J2_124_3477_n2211), .CI(DP_OP_422J2_124_3477_n2218), .CO(
        DP_OP_422J2_124_3477_n1692), .S(DP_OP_422J2_124_3477_n1693) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1028 ( .A(DP_OP_422J2_124_3477_n2600), .B(
        DP_OP_422J2_124_3477_n2248), .CI(DP_OP_422J2_124_3477_n2255), .CO(
        DP_OP_422J2_124_3477_n1690), .S(DP_OP_422J2_124_3477_n1691) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1027 ( .A(DP_OP_422J2_124_3477_n2607), .B(
        DP_OP_422J2_124_3477_n2262), .CI(DP_OP_422J2_124_3477_n2292), .CO(
        DP_OP_422J2_124_3477_n1688), .S(DP_OP_422J2_124_3477_n1689) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1026 ( .A(DP_OP_422J2_124_3477_n2614), .B(
        DP_OP_422J2_124_3477_n2966), .CI(DP_OP_422J2_124_3477_n2299), .CO(
        DP_OP_422J2_124_3477_n1686), .S(DP_OP_422J2_124_3477_n1687) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1025 ( .A(DP_OP_422J2_124_3477_n2644), .B(
        DP_OP_422J2_124_3477_n2306), .CI(DP_OP_422J2_124_3477_n2959), .CO(
        DP_OP_422J2_124_3477_n1684), .S(DP_OP_422J2_124_3477_n1685) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1023 ( .A(DP_OP_422J2_124_3477_n2482), .B(
        DP_OP_422J2_124_3477_n2915), .CI(DP_OP_422J2_124_3477_n2336), .CO(
        DP_OP_422J2_124_3477_n1680), .S(DP_OP_422J2_124_3477_n1681) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1022 ( .A(DP_OP_422J2_124_3477_n2908), .B(
        DP_OP_422J2_124_3477_n2343), .CI(DP_OP_422J2_124_3477_n2878), .CO(
        DP_OP_422J2_124_3477_n1678), .S(DP_OP_422J2_124_3477_n1679) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1021 ( .A(DP_OP_422J2_124_3477_n2871), .B(
        DP_OP_422J2_124_3477_n2864), .CI(DP_OP_422J2_124_3477_n2350), .CO(
        DP_OP_422J2_124_3477_n1676), .S(DP_OP_422J2_124_3477_n1677) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1020 ( .A(DP_OP_422J2_124_3477_n2475), .B(
        DP_OP_422J2_124_3477_n2380), .CI(DP_OP_422J2_124_3477_n2834), .CO(
        DP_OP_422J2_124_3477_n1674), .S(DP_OP_422J2_124_3477_n1675) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1019 ( .A(DP_OP_422J2_124_3477_n2468), .B(
        DP_OP_422J2_124_3477_n2827), .CI(DP_OP_422J2_124_3477_n2820), .CO(
        DP_OP_422J2_124_3477_n1672), .S(DP_OP_422J2_124_3477_n1673) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1018 ( .A(DP_OP_422J2_124_3477_n2424), .B(
        DP_OP_422J2_124_3477_n2790), .CI(DP_OP_422J2_124_3477_n2783), .CO(
        DP_OP_422J2_124_3477_n1670), .S(DP_OP_422J2_124_3477_n1671) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1017 ( .A(DP_OP_422J2_124_3477_n2387), .B(
        DP_OP_422J2_124_3477_n2776), .CI(DP_OP_422J2_124_3477_n2746), .CO(
        DP_OP_422J2_124_3477_n1668), .S(DP_OP_422J2_124_3477_n1669) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1016 ( .A(DP_OP_422J2_124_3477_n2658), .B(
        DP_OP_422J2_124_3477_n2739), .CI(DP_OP_422J2_124_3477_n2394), .CO(
        DP_OP_422J2_124_3477_n1666), .S(DP_OP_422J2_124_3477_n1667) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1015 ( .A(DP_OP_422J2_124_3477_n2512), .B(
        DP_OP_422J2_124_3477_n2431), .CI(DP_OP_422J2_124_3477_n2732), .CO(
        DP_OP_422J2_124_3477_n1664), .S(DP_OP_422J2_124_3477_n1665) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1014 ( .A(DP_OP_422J2_124_3477_n2702), .B(
        DP_OP_422J2_124_3477_n2438), .CI(DP_OP_422J2_124_3477_n2651), .CO(
        DP_OP_422J2_124_3477_n1662), .S(DP_OP_422J2_124_3477_n1663) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1012 ( .A(DP_OP_422J2_124_3477_n1810), .B(
        DP_OP_422J2_124_3477_n1832), .CI(DP_OP_422J2_124_3477_n1786), .CO(
        DP_OP_422J2_124_3477_n1658), .S(DP_OP_422J2_124_3477_n1659) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1011 ( .A(DP_OP_422J2_124_3477_n1808), .B(
        DP_OP_422J2_124_3477_n1830), .CI(DP_OP_422J2_124_3477_n1828), .CO(
        DP_OP_422J2_124_3477_n1656), .S(DP_OP_422J2_124_3477_n1657) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1010 ( .A(DP_OP_422J2_124_3477_n1824), .B(
        DP_OP_422J2_124_3477_n1826), .CI(DP_OP_422J2_124_3477_n1802), .CO(
        DP_OP_422J2_124_3477_n1654), .S(DP_OP_422J2_124_3477_n1655) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1009 ( .A(DP_OP_422J2_124_3477_n1798), .B(
        DP_OP_422J2_124_3477_n1788), .CI(DP_OP_422J2_124_3477_n1790), .CO(
        DP_OP_422J2_124_3477_n1652), .S(DP_OP_422J2_124_3477_n1653) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1008 ( .A(DP_OP_422J2_124_3477_n1796), .B(
        DP_OP_422J2_124_3477_n1822), .CI(DP_OP_422J2_124_3477_n1792), .CO(
        DP_OP_422J2_124_3477_n1650), .S(DP_OP_422J2_124_3477_n1651) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1007 ( .A(DP_OP_422J2_124_3477_n1794), .B(
        DP_OP_422J2_124_3477_n1820), .CI(DP_OP_422J2_124_3477_n1818), .CO(
        DP_OP_422J2_124_3477_n1648), .S(DP_OP_422J2_124_3477_n1649) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1006 ( .A(DP_OP_422J2_124_3477_n1806), .B(
        DP_OP_422J2_124_3477_n1816), .CI(DP_OP_422J2_124_3477_n1800), .CO(
        DP_OP_422J2_124_3477_n1646), .S(DP_OP_422J2_124_3477_n1647) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1005 ( .A(DP_OP_422J2_124_3477_n1814), .B(
        DP_OP_422J2_124_3477_n1812), .CI(DP_OP_422J2_124_3477_n1804), .CO(
        DP_OP_422J2_124_3477_n1644), .S(DP_OP_422J2_124_3477_n1645) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1004 ( .A(DP_OP_422J2_124_3477_n1723), .B(
        DP_OP_422J2_124_3477_n1725), .CI(DP_OP_422J2_124_3477_n1711), .CO(
        DP_OP_422J2_124_3477_n1642), .S(DP_OP_422J2_124_3477_n1643) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1003 ( .A(DP_OP_422J2_124_3477_n1717), .B(
        DP_OP_422J2_124_3477_n1719), .CI(DP_OP_422J2_124_3477_n1784), .CO(
        DP_OP_422J2_124_3477_n1640), .S(DP_OP_422J2_124_3477_n1641) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1002 ( .A(DP_OP_422J2_124_3477_n1713), .B(
        DP_OP_422J2_124_3477_n1715), .CI(DP_OP_422J2_124_3477_n1721), .CO(
        DP_OP_422J2_124_3477_n1638), .S(DP_OP_422J2_124_3477_n1639) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1001 ( .A(DP_OP_422J2_124_3477_n1727), .B(
        DP_OP_422J2_124_3477_n1677), .CI(DP_OP_422J2_124_3477_n1675), .CO(
        DP_OP_422J2_124_3477_n1636), .S(DP_OP_422J2_124_3477_n1637) );
  FADDX1_HVT DP_OP_422J2_124_3477_U1000 ( .A(DP_OP_422J2_124_3477_n1679), .B(
        DP_OP_422J2_124_3477_n1695), .CI(DP_OP_422J2_124_3477_n1703), .CO(
        DP_OP_422J2_124_3477_n1634), .S(DP_OP_422J2_124_3477_n1635) );
  FADDX1_HVT DP_OP_422J2_124_3477_U999 ( .A(DP_OP_422J2_124_3477_n1671), .B(
        DP_OP_422J2_124_3477_n1691), .CI(DP_OP_422J2_124_3477_n1689), .CO(
        DP_OP_422J2_124_3477_n1632), .S(DP_OP_422J2_124_3477_n1633) );
  FADDX1_HVT DP_OP_422J2_124_3477_U998 ( .A(DP_OP_422J2_124_3477_n1669), .B(
        DP_OP_422J2_124_3477_n1705), .CI(DP_OP_422J2_124_3477_n1693), .CO(
        DP_OP_422J2_124_3477_n1630), .S(DP_OP_422J2_124_3477_n1631) );
  FADDX1_HVT DP_OP_422J2_124_3477_U997 ( .A(DP_OP_422J2_124_3477_n1667), .B(
        DP_OP_422J2_124_3477_n1699), .CI(DP_OP_422J2_124_3477_n1701), .CO(
        DP_OP_422J2_124_3477_n1628), .S(DP_OP_422J2_124_3477_n1629) );
  FADDX1_HVT DP_OP_422J2_124_3477_U996 ( .A(DP_OP_422J2_124_3477_n1665), .B(
        DP_OP_422J2_124_3477_n1697), .CI(DP_OP_422J2_124_3477_n1709), .CO(
        DP_OP_422J2_124_3477_n1626), .S(DP_OP_422J2_124_3477_n1627) );
  FADDX1_HVT DP_OP_422J2_124_3477_U995 ( .A(DP_OP_422J2_124_3477_n1687), .B(
        DP_OP_422J2_124_3477_n1707), .CI(DP_OP_422J2_124_3477_n1663), .CO(
        DP_OP_422J2_124_3477_n1624), .S(DP_OP_422J2_124_3477_n1625) );
  FADDX1_HVT DP_OP_422J2_124_3477_U994 ( .A(DP_OP_422J2_124_3477_n1673), .B(
        DP_OP_422J2_124_3477_n1683), .CI(DP_OP_422J2_124_3477_n1685), .CO(
        DP_OP_422J2_124_3477_n1622), .S(DP_OP_422J2_124_3477_n1623) );
  FADDX1_HVT DP_OP_422J2_124_3477_U993 ( .A(DP_OP_422J2_124_3477_n1681), .B(
        DP_OP_422J2_124_3477_n1661), .CI(DP_OP_422J2_124_3477_n1782), .CO(
        DP_OP_422J2_124_3477_n1620), .S(DP_OP_422J2_124_3477_n1621) );
  FADDX1_HVT DP_OP_422J2_124_3477_U992 ( .A(DP_OP_422J2_124_3477_n1780), .B(
        DP_OP_422J2_124_3477_n1778), .CI(DP_OP_422J2_124_3477_n1776), .CO(
        DP_OP_422J2_124_3477_n1618), .S(DP_OP_422J2_124_3477_n1619) );
  FADDX1_HVT DP_OP_422J2_124_3477_U991 ( .A(DP_OP_422J2_124_3477_n1774), .B(
        DP_OP_422J2_124_3477_n1772), .CI(DP_OP_422J2_124_3477_n1760), .CO(
        DP_OP_422J2_124_3477_n1616), .S(DP_OP_422J2_124_3477_n1617) );
  FADDX1_HVT DP_OP_422J2_124_3477_U990 ( .A(DP_OP_422J2_124_3477_n1758), .B(
        DP_OP_422J2_124_3477_n1659), .CI(DP_OP_422J2_124_3477_n1756), .CO(
        DP_OP_422J2_124_3477_n1614), .S(DP_OP_422J2_124_3477_n1615) );
  FADDX1_HVT DP_OP_422J2_124_3477_U989 ( .A(DP_OP_422J2_124_3477_n1657), .B(
        DP_OP_422J2_124_3477_n1649), .CI(DP_OP_422J2_124_3477_n1770), .CO(
        DP_OP_422J2_124_3477_n1612), .S(DP_OP_422J2_124_3477_n1613) );
  FADDX1_HVT DP_OP_422J2_124_3477_U988 ( .A(DP_OP_422J2_124_3477_n1768), .B(
        DP_OP_422J2_124_3477_n1647), .CI(DP_OP_422J2_124_3477_n1651), .CO(
        DP_OP_422J2_124_3477_n1610), .S(DP_OP_422J2_124_3477_n1611) );
  FADDX1_HVT DP_OP_422J2_124_3477_U987 ( .A(DP_OP_422J2_124_3477_n1764), .B(
        DP_OP_422J2_124_3477_n1653), .CI(DP_OP_422J2_124_3477_n1655), .CO(
        DP_OP_422J2_124_3477_n1608), .S(DP_OP_422J2_124_3477_n1609) );
  FADDX1_HVT DP_OP_422J2_124_3477_U986 ( .A(DP_OP_422J2_124_3477_n1762), .B(
        DP_OP_422J2_124_3477_n1766), .CI(DP_OP_422J2_124_3477_n1645), .CO(
        DP_OP_422J2_124_3477_n1606), .S(DP_OP_422J2_124_3477_n1607) );
  FADDX1_HVT DP_OP_422J2_124_3477_U985 ( .A(DP_OP_422J2_124_3477_n1641), .B(
        DP_OP_422J2_124_3477_n1643), .CI(DP_OP_422J2_124_3477_n1637), .CO(
        DP_OP_422J2_124_3477_n1604), .S(DP_OP_422J2_124_3477_n1605) );
  FADDX1_HVT DP_OP_422J2_124_3477_U984 ( .A(DP_OP_422J2_124_3477_n1639), .B(
        DP_OP_422J2_124_3477_n1625), .CI(DP_OP_422J2_124_3477_n1627), .CO(
        DP_OP_422J2_124_3477_n1602), .S(DP_OP_422J2_124_3477_n1603) );
  FADDX1_HVT DP_OP_422J2_124_3477_U983 ( .A(DP_OP_422J2_124_3477_n1633), .B(
        DP_OP_422J2_124_3477_n1631), .CI(DP_OP_422J2_124_3477_n1754), .CO(
        DP_OP_422J2_124_3477_n1600), .S(DP_OP_422J2_124_3477_n1601) );
  FADDX1_HVT DP_OP_422J2_124_3477_U982 ( .A(DP_OP_422J2_124_3477_n1629), .B(
        DP_OP_422J2_124_3477_n1623), .CI(DP_OP_422J2_124_3477_n1635), .CO(
        DP_OP_422J2_124_3477_n1598), .S(DP_OP_422J2_124_3477_n1599) );
  FADDX1_HVT DP_OP_422J2_124_3477_U981 ( .A(DP_OP_422J2_124_3477_n1621), .B(
        DP_OP_422J2_124_3477_n1752), .CI(DP_OP_422J2_124_3477_n1748), .CO(
        DP_OP_422J2_124_3477_n1596), .S(DP_OP_422J2_124_3477_n1597) );
  FADDX1_HVT DP_OP_422J2_124_3477_U980 ( .A(DP_OP_422J2_124_3477_n1750), .B(
        DP_OP_422J2_124_3477_n1619), .CI(DP_OP_422J2_124_3477_n1746), .CO(
        DP_OP_422J2_124_3477_n1594), .S(DP_OP_422J2_124_3477_n1595) );
  FADDX1_HVT DP_OP_422J2_124_3477_U979 ( .A(DP_OP_422J2_124_3477_n1617), .B(
        DP_OP_422J2_124_3477_n1607), .CI(DP_OP_422J2_124_3477_n1609), .CO(
        DP_OP_422J2_124_3477_n1592), .S(DP_OP_422J2_124_3477_n1593) );
  FADDX1_HVT DP_OP_422J2_124_3477_U978 ( .A(DP_OP_422J2_124_3477_n1611), .B(
        DP_OP_422J2_124_3477_n1744), .CI(DP_OP_422J2_124_3477_n1742), .CO(
        DP_OP_422J2_124_3477_n1590), .S(DP_OP_422J2_124_3477_n1591) );
  FADDX1_HVT DP_OP_422J2_124_3477_U977 ( .A(DP_OP_422J2_124_3477_n1615), .B(
        DP_OP_422J2_124_3477_n1613), .CI(DP_OP_422J2_124_3477_n1605), .CO(
        DP_OP_422J2_124_3477_n1588), .S(DP_OP_422J2_124_3477_n1589) );
  FADDX1_HVT DP_OP_422J2_124_3477_U976 ( .A(DP_OP_422J2_124_3477_n1740), .B(
        DP_OP_422J2_124_3477_n1603), .CI(DP_OP_422J2_124_3477_n1599), .CO(
        DP_OP_422J2_124_3477_n1586), .S(DP_OP_422J2_124_3477_n1587) );
  FADDX1_HVT DP_OP_422J2_124_3477_U975 ( .A(DP_OP_422J2_124_3477_n1601), .B(
        DP_OP_422J2_124_3477_n1738), .CI(DP_OP_422J2_124_3477_n1597), .CO(
        DP_OP_422J2_124_3477_n1584), .S(DP_OP_422J2_124_3477_n1585) );
  FADDX1_HVT DP_OP_422J2_124_3477_U974 ( .A(DP_OP_422J2_124_3477_n1736), .B(
        DP_OP_422J2_124_3477_n1595), .CI(DP_OP_422J2_124_3477_n1734), .CO(
        DP_OP_422J2_124_3477_n1582), .S(DP_OP_422J2_124_3477_n1583) );
  FADDX1_HVT DP_OP_422J2_124_3477_U973 ( .A(DP_OP_422J2_124_3477_n1593), .B(
        DP_OP_422J2_124_3477_n1591), .CI(DP_OP_422J2_124_3477_n1589), .CO(
        DP_OP_422J2_124_3477_n1580), .S(DP_OP_422J2_124_3477_n1581) );
  FADDX1_HVT DP_OP_422J2_124_3477_U972 ( .A(DP_OP_422J2_124_3477_n1587), .B(
        DP_OP_422J2_124_3477_n1732), .CI(DP_OP_422J2_124_3477_n1585), .CO(
        DP_OP_422J2_124_3477_n1578), .S(DP_OP_422J2_124_3477_n1579) );
  FADDX1_HVT DP_OP_422J2_124_3477_U971 ( .A(DP_OP_422J2_124_3477_n1730), .B(
        DP_OP_422J2_124_3477_n1583), .CI(DP_OP_422J2_124_3477_n1581), .CO(
        DP_OP_422J2_124_3477_n1576), .S(DP_OP_422J2_124_3477_n1577) );
  FADDX1_HVT DP_OP_422J2_124_3477_U970 ( .A(DP_OP_422J2_124_3477_n1728), .B(
        DP_OP_422J2_124_3477_n1976), .CI(DP_OP_422J2_124_3477_n1932), .CO(
        DP_OP_422J2_124_3477_n1574), .S(DP_OP_422J2_124_3477_n1575) );
  FADDX1_HVT DP_OP_422J2_124_3477_U969 ( .A(DP_OP_422J2_124_3477_n3031), .B(
        DP_OP_422J2_124_3477_n2548), .CI(DP_OP_422J2_124_3477_n2416), .CO(
        DP_OP_422J2_124_3477_n1572), .S(DP_OP_422J2_124_3477_n1573) );
  FADDX1_HVT DP_OP_422J2_124_3477_U968 ( .A(DP_OP_422J2_124_3477_n2944), .B(
        DP_OP_422J2_124_3477_n2680), .CI(DP_OP_422J2_124_3477_n2328), .CO(
        DP_OP_422J2_124_3477_n1570), .S(DP_OP_422J2_124_3477_n1571) );
  FADDX1_HVT DP_OP_422J2_124_3477_U967 ( .A(DP_OP_422J2_124_3477_n2108), .B(
        DP_OP_422J2_124_3477_n2636), .CI(DP_OP_422J2_124_3477_n2856), .CO(
        DP_OP_422J2_124_3477_n1568), .S(DP_OP_422J2_124_3477_n1569) );
  FADDX1_HVT DP_OP_422J2_124_3477_U966 ( .A(DP_OP_422J2_124_3477_n2196), .B(
        DP_OP_422J2_124_3477_n2372), .CI(DP_OP_422J2_124_3477_n2460), .CO(
        DP_OP_422J2_124_3477_n1566), .S(DP_OP_422J2_124_3477_n1567) );
  FADDX1_HVT DP_OP_422J2_124_3477_U965 ( .A(DP_OP_422J2_124_3477_n2812), .B(
        DP_OP_422J2_124_3477_n2284), .CI(DP_OP_422J2_124_3477_n2900), .CO(
        DP_OP_422J2_124_3477_n1564), .S(DP_OP_422J2_124_3477_n1565) );
  FADDX1_HVT DP_OP_422J2_124_3477_U964 ( .A(DP_OP_422J2_124_3477_n2152), .B(
        DP_OP_422J2_124_3477_n2504), .CI(DP_OP_422J2_124_3477_n2592), .CO(
        DP_OP_422J2_124_3477_n1562), .S(DP_OP_422J2_124_3477_n1563) );
  FADDX1_HVT DP_OP_422J2_124_3477_U963 ( .A(DP_OP_422J2_124_3477_n2988), .B(
        DP_OP_422J2_124_3477_n2724), .CI(DP_OP_422J2_124_3477_n2768), .CO(
        DP_OP_422J2_124_3477_n1560), .S(DP_OP_422J2_124_3477_n1561) );
  FADDX1_HVT DP_OP_422J2_124_3477_U962 ( .A(DP_OP_422J2_124_3477_n2064), .B(
        DP_OP_422J2_124_3477_n2240), .CI(DP_OP_422J2_124_3477_n2020), .CO(
        DP_OP_422J2_124_3477_n1558), .S(DP_OP_422J2_124_3477_n1559) );
  FADDX1_HVT DP_OP_422J2_124_3477_U961 ( .A(DP_OP_422J2_124_3477_n2555), .B(
        DP_OP_422J2_124_3477_n1990), .CI(DP_OP_422J2_124_3477_n1983), .CO(
        DP_OP_422J2_124_3477_n1556), .S(DP_OP_422J2_124_3477_n1557) );
  FADDX1_HVT DP_OP_422J2_124_3477_U960 ( .A(DP_OP_422J2_124_3477_n3051), .B(
        DP_OP_422J2_124_3477_n1997), .CI(DP_OP_422J2_124_3477_n2027), .CO(
        DP_OP_422J2_124_3477_n1554), .S(DP_OP_422J2_124_3477_n1555) );
  FADDX1_HVT DP_OP_422J2_124_3477_U959 ( .A(DP_OP_422J2_124_3477_n2437), .B(
        DP_OP_422J2_124_3477_n3044), .CI(DP_OP_422J2_124_3477_n2034), .CO(
        DP_OP_422J2_124_3477_n1552), .S(DP_OP_422J2_124_3477_n1553) );
  FADDX1_HVT DP_OP_422J2_124_3477_U958 ( .A(DP_OP_422J2_124_3477_n2430), .B(
        DP_OP_422J2_124_3477_n3037), .CI(DP_OP_422J2_124_3477_n2041), .CO(
        DP_OP_422J2_124_3477_n1550), .S(DP_OP_422J2_124_3477_n1551) );
  FADDX1_HVT DP_OP_422J2_124_3477_U957 ( .A(DP_OP_422J2_124_3477_n3009), .B(
        DP_OP_422J2_124_3477_n2071), .CI(DP_OP_422J2_124_3477_n2078), .CO(
        DP_OP_422J2_124_3477_n1548), .S(DP_OP_422J2_124_3477_n1549) );
  FADDX1_HVT DP_OP_422J2_124_3477_U956 ( .A(DP_OP_422J2_124_3477_n2467), .B(
        DP_OP_422J2_124_3477_n3002), .CI(DP_OP_422J2_124_3477_n2995), .CO(
        DP_OP_422J2_124_3477_n1546), .S(DP_OP_422J2_124_3477_n1547) );
  FADDX1_HVT DP_OP_422J2_124_3477_U955 ( .A(DP_OP_422J2_124_3477_n2393), .B(
        DP_OP_422J2_124_3477_n2965), .CI(DP_OP_422J2_124_3477_n2958), .CO(
        DP_OP_422J2_124_3477_n1544), .S(DP_OP_422J2_124_3477_n1545) );
  FADDX1_HVT DP_OP_422J2_124_3477_U954 ( .A(DP_OP_422J2_124_3477_n2386), .B(
        DP_OP_422J2_124_3477_n2951), .CI(DP_OP_422J2_124_3477_n2085), .CO(
        DP_OP_422J2_124_3477_n1542), .S(DP_OP_422J2_124_3477_n1543) );
  FADDX1_HVT DP_OP_422J2_124_3477_U953 ( .A(DP_OP_422J2_124_3477_n2379), .B(
        DP_OP_422J2_124_3477_n2921), .CI(DP_OP_422J2_124_3477_n2914), .CO(
        DP_OP_422J2_124_3477_n1540), .S(DP_OP_422J2_124_3477_n1541) );
  FADDX1_HVT DP_OP_422J2_124_3477_U952 ( .A(DP_OP_422J2_124_3477_n2349), .B(
        DP_OP_422J2_124_3477_n2907), .CI(DP_OP_422J2_124_3477_n2115), .CO(
        DP_OP_422J2_124_3477_n1538), .S(DP_OP_422J2_124_3477_n1539) );
  FADDX1_HVT DP_OP_422J2_124_3477_U951 ( .A(DP_OP_422J2_124_3477_n2342), .B(
        DP_OP_422J2_124_3477_n2122), .CI(DP_OP_422J2_124_3477_n2129), .CO(
        DP_OP_422J2_124_3477_n1536), .S(DP_OP_422J2_124_3477_n1537) );
  FADDX1_HVT DP_OP_422J2_124_3477_U950 ( .A(DP_OP_422J2_124_3477_n2423), .B(
        DP_OP_422J2_124_3477_n2159), .CI(DP_OP_422J2_124_3477_n2877), .CO(
        DP_OP_422J2_124_3477_n1534), .S(DP_OP_422J2_124_3477_n1535) );
  FADDX1_HVT DP_OP_422J2_124_3477_U949 ( .A(DP_OP_422J2_124_3477_n2474), .B(
        DP_OP_422J2_124_3477_n2870), .CI(DP_OP_422J2_124_3477_n2863), .CO(
        DP_OP_422J2_124_3477_n1532), .S(DP_OP_422J2_124_3477_n1533) );
  FADDX1_HVT DP_OP_422J2_124_3477_U948 ( .A(DP_OP_422J2_124_3477_n2833), .B(
        DP_OP_422J2_124_3477_n2166), .CI(DP_OP_422J2_124_3477_n2173), .CO(
        DP_OP_422J2_124_3477_n1530), .S(DP_OP_422J2_124_3477_n1531) );
  FADDX1_HVT DP_OP_422J2_124_3477_U947 ( .A(DP_OP_422J2_124_3477_n2606), .B(
        DP_OP_422J2_124_3477_n2203), .CI(DP_OP_422J2_124_3477_n2210), .CO(
        DP_OP_422J2_124_3477_n1528), .S(DP_OP_422J2_124_3477_n1529) );
  FADDX1_HVT DP_OP_422J2_124_3477_U946 ( .A(DP_OP_422J2_124_3477_n2826), .B(
        DP_OP_422J2_124_3477_n2217), .CI(DP_OP_422J2_124_3477_n2247), .CO(
        DP_OP_422J2_124_3477_n1526), .S(DP_OP_422J2_124_3477_n1527) );
  FADDX1_HVT DP_OP_422J2_124_3477_U945 ( .A(DP_OP_422J2_124_3477_n2819), .B(
        DP_OP_422J2_124_3477_n2254), .CI(DP_OP_422J2_124_3477_n2261), .CO(
        DP_OP_422J2_124_3477_n1524), .S(DP_OP_422J2_124_3477_n1525) );
  FADDX1_HVT DP_OP_422J2_124_3477_U944 ( .A(DP_OP_422J2_124_3477_n2789), .B(
        DP_OP_422J2_124_3477_n2291), .CI(DP_OP_422J2_124_3477_n2298), .CO(
        DP_OP_422J2_124_3477_n1522), .S(DP_OP_422J2_124_3477_n1523) );
  FADDX1_HVT DP_OP_422J2_124_3477_U943 ( .A(DP_OP_422J2_124_3477_n2782), .B(
        DP_OP_422J2_124_3477_n2305), .CI(DP_OP_422J2_124_3477_n2335), .CO(
        DP_OP_422J2_124_3477_n1520), .S(DP_OP_422J2_124_3477_n1521) );
  FADDX1_HVT DP_OP_422J2_124_3477_U942 ( .A(DP_OP_422J2_124_3477_n2775), .B(
        DP_OP_422J2_124_3477_n2481), .CI(DP_OP_422J2_124_3477_n2511), .CO(
        DP_OP_422J2_124_3477_n1518), .S(DP_OP_422J2_124_3477_n1519) );
  FADDX1_HVT DP_OP_422J2_124_3477_U941 ( .A(DP_OP_422J2_124_3477_n2745), .B(
        DP_OP_422J2_124_3477_n2518), .CI(DP_OP_422J2_124_3477_n2738), .CO(
        DP_OP_422J2_124_3477_n1516), .S(DP_OP_422J2_124_3477_n1517) );
  FADDX1_HVT DP_OP_422J2_124_3477_U940 ( .A(DP_OP_422J2_124_3477_n2643), .B(
        DP_OP_422J2_124_3477_n2525), .CI(DP_OP_422J2_124_3477_n2562), .CO(
        DP_OP_422J2_124_3477_n1514), .S(DP_OP_422J2_124_3477_n1515) );
  FADDX1_HVT DP_OP_422J2_124_3477_U939 ( .A(DP_OP_422J2_124_3477_n2613), .B(
        DP_OP_422J2_124_3477_n2569), .CI(DP_OP_422J2_124_3477_n2731), .CO(
        DP_OP_422J2_124_3477_n1512), .S(DP_OP_422J2_124_3477_n1513) );
  FADDX1_HVT DP_OP_422J2_124_3477_U938 ( .A(DP_OP_422J2_124_3477_n2687), .B(
        DP_OP_422J2_124_3477_n2599), .CI(DP_OP_422J2_124_3477_n2701), .CO(
        DP_OP_422J2_124_3477_n1510), .S(DP_OP_422J2_124_3477_n1511) );
  FADDX1_HVT DP_OP_422J2_124_3477_U937 ( .A(DP_OP_422J2_124_3477_n2650), .B(
        DP_OP_422J2_124_3477_n2657), .CI(DP_OP_422J2_124_3477_n2694), .CO(
        DP_OP_422J2_124_3477_n1508), .S(DP_OP_422J2_124_3477_n1509) );
  FADDX1_HVT DP_OP_422J2_124_3477_U936 ( .A(DP_OP_422J2_124_3477_n1716), .B(
        DP_OP_422J2_124_3477_n1712), .CI(DP_OP_422J2_124_3477_n1710), .CO(
        DP_OP_422J2_124_3477_n1506), .S(DP_OP_422J2_124_3477_n1507) );
  FADDX1_HVT DP_OP_422J2_124_3477_U935 ( .A(DP_OP_422J2_124_3477_n1714), .B(
        DP_OP_422J2_124_3477_n1718), .CI(DP_OP_422J2_124_3477_n1720), .CO(
        DP_OP_422J2_124_3477_n1504), .S(DP_OP_422J2_124_3477_n1505) );
  FADDX1_HVT DP_OP_422J2_124_3477_U934 ( .A(DP_OP_422J2_124_3477_n1722), .B(
        DP_OP_422J2_124_3477_n1724), .CI(DP_OP_422J2_124_3477_n1726), .CO(
        DP_OP_422J2_124_3477_n1502), .S(DP_OP_422J2_124_3477_n1503) );
  FADDX1_HVT DP_OP_422J2_124_3477_U933 ( .A(DP_OP_422J2_124_3477_n1686), .B(
        DP_OP_422J2_124_3477_n1708), .CI(DP_OP_422J2_124_3477_n1706), .CO(
        DP_OP_422J2_124_3477_n1500), .S(DP_OP_422J2_124_3477_n1501) );
  FADDX1_HVT DP_OP_422J2_124_3477_U932 ( .A(DP_OP_422J2_124_3477_n1682), .B(
        DP_OP_422J2_124_3477_n1704), .CI(DP_OP_422J2_124_3477_n1702), .CO(
        DP_OP_422J2_124_3477_n1498), .S(DP_OP_422J2_124_3477_n1499) );
  FADDX1_HVT DP_OP_422J2_124_3477_U931 ( .A(DP_OP_422J2_124_3477_n1676), .B(
        DP_OP_422J2_124_3477_n1700), .CI(DP_OP_422J2_124_3477_n1698), .CO(
        DP_OP_422J2_124_3477_n1496), .S(DP_OP_422J2_124_3477_n1497) );
  FADDX1_HVT DP_OP_422J2_124_3477_U929 ( .A(DP_OP_422J2_124_3477_n1668), .B(
        DP_OP_422J2_124_3477_n1694), .CI(DP_OP_422J2_124_3477_n1692), .CO(
        DP_OP_422J2_124_3477_n1492), .S(DP_OP_422J2_124_3477_n1493) );
  FADDX1_HVT DP_OP_422J2_124_3477_U928 ( .A(DP_OP_422J2_124_3477_n1678), .B(
        DP_OP_422J2_124_3477_n1690), .CI(DP_OP_422J2_124_3477_n1688), .CO(
        DP_OP_422J2_124_3477_n1490), .S(DP_OP_422J2_124_3477_n1491) );
  FADDX1_HVT DP_OP_422J2_124_3477_U927 ( .A(DP_OP_422J2_124_3477_n1670), .B(
        DP_OP_422J2_124_3477_n1684), .CI(DP_OP_422J2_124_3477_n1680), .CO(
        DP_OP_422J2_124_3477_n1488), .S(DP_OP_422J2_124_3477_n1489) );
  FADDX1_HVT DP_OP_422J2_124_3477_U926 ( .A(DP_OP_422J2_124_3477_n1666), .B(
        DP_OP_422J2_124_3477_n1674), .CI(DP_OP_422J2_124_3477_n1664), .CO(
        DP_OP_422J2_124_3477_n1486), .S(DP_OP_422J2_124_3477_n1487) );
  FADDX1_HVT DP_OP_422J2_124_3477_U925 ( .A(DP_OP_422J2_124_3477_n1575), .B(
        DP_OP_422J2_124_3477_n1559), .CI(DP_OP_422J2_124_3477_n1660), .CO(
        DP_OP_422J2_124_3477_n1484), .S(DP_OP_422J2_124_3477_n1485) );
  FADDX1_HVT DP_OP_422J2_124_3477_U924 ( .A(DP_OP_422J2_124_3477_n1573), .B(
        DP_OP_422J2_124_3477_n1561), .CI(DP_OP_422J2_124_3477_n1563), .CO(
        DP_OP_422J2_124_3477_n1482), .S(DP_OP_422J2_124_3477_n1483) );
  FADDX1_HVT DP_OP_422J2_124_3477_U923 ( .A(DP_OP_422J2_124_3477_n1569), .B(
        DP_OP_422J2_124_3477_n1567), .CI(DP_OP_422J2_124_3477_n1571), .CO(
        DP_OP_422J2_124_3477_n1480), .S(DP_OP_422J2_124_3477_n1481) );
  FADDX1_HVT DP_OP_422J2_124_3477_U922 ( .A(DP_OP_422J2_124_3477_n1565), .B(
        DP_OP_422J2_124_3477_n1545), .CI(DP_OP_422J2_124_3477_n1549), .CO(
        DP_OP_422J2_124_3477_n1478), .S(DP_OP_422J2_124_3477_n1479) );
  FADDX1_HVT DP_OP_422J2_124_3477_U921 ( .A(DP_OP_422J2_124_3477_n1547), .B(
        DP_OP_422J2_124_3477_n1555), .CI(DP_OP_422J2_124_3477_n1553), .CO(
        DP_OP_422J2_124_3477_n1476), .S(DP_OP_422J2_124_3477_n1477) );
  FADDX1_HVT DP_OP_422J2_124_3477_U920 ( .A(DP_OP_422J2_124_3477_n1557), .B(
        DP_OP_422J2_124_3477_n1535), .CI(DP_OP_422J2_124_3477_n1529), .CO(
        DP_OP_422J2_124_3477_n1474), .S(DP_OP_422J2_124_3477_n1475) );
  FADDX1_HVT DP_OP_422J2_124_3477_U919 ( .A(DP_OP_422J2_124_3477_n1537), .B(
        DP_OP_422J2_124_3477_n1533), .CI(DP_OP_422J2_124_3477_n1527), .CO(
        DP_OP_422J2_124_3477_n1472), .S(DP_OP_422J2_124_3477_n1473) );
  FADDX1_HVT DP_OP_422J2_124_3477_U918 ( .A(DP_OP_422J2_124_3477_n1539), .B(
        DP_OP_422J2_124_3477_n1513), .CI(DP_OP_422J2_124_3477_n1511), .CO(
        DP_OP_422J2_124_3477_n1470), .S(DP_OP_422J2_124_3477_n1471) );
  FADDX1_HVT DP_OP_422J2_124_3477_U917 ( .A(DP_OP_422J2_124_3477_n1525), .B(
        DP_OP_422J2_124_3477_n1521), .CI(DP_OP_422J2_124_3477_n1523), .CO(
        DP_OP_422J2_124_3477_n1468), .S(DP_OP_422J2_124_3477_n1469) );
  FADDX1_HVT DP_OP_422J2_124_3477_U916 ( .A(DP_OP_422J2_124_3477_n1531), .B(
        DP_OP_422J2_124_3477_n1509), .CI(DP_OP_422J2_124_3477_n1517), .CO(
        DP_OP_422J2_124_3477_n1466), .S(DP_OP_422J2_124_3477_n1467) );
  FADDX1_HVT DP_OP_422J2_124_3477_U915 ( .A(DP_OP_422J2_124_3477_n1519), .B(
        DP_OP_422J2_124_3477_n1543), .CI(DP_OP_422J2_124_3477_n1551), .CO(
        DP_OP_422J2_124_3477_n1464), .S(DP_OP_422J2_124_3477_n1465) );
  FADDX1_HVT DP_OP_422J2_124_3477_U914 ( .A(DP_OP_422J2_124_3477_n1515), .B(
        DP_OP_422J2_124_3477_n1541), .CI(DP_OP_422J2_124_3477_n1658), .CO(
        DP_OP_422J2_124_3477_n1462), .S(DP_OP_422J2_124_3477_n1463) );
  FADDX1_HVT DP_OP_422J2_124_3477_U912 ( .A(DP_OP_422J2_124_3477_n1644), .B(
        DP_OP_422J2_124_3477_n1650), .CI(DP_OP_422J2_124_3477_n1646), .CO(
        DP_OP_422J2_124_3477_n1458), .S(DP_OP_422J2_124_3477_n1459) );
  FADDX1_HVT DP_OP_422J2_124_3477_U911 ( .A(DP_OP_422J2_124_3477_n1648), .B(
        DP_OP_422J2_124_3477_n1642), .CI(DP_OP_422J2_124_3477_n1503), .CO(
        DP_OP_422J2_124_3477_n1456), .S(DP_OP_422J2_124_3477_n1457) );
  FADDX1_HVT DP_OP_422J2_124_3477_U910 ( .A(DP_OP_422J2_124_3477_n1505), .B(
        DP_OP_422J2_124_3477_n1640), .CI(DP_OP_422J2_124_3477_n1636), .CO(
        DP_OP_422J2_124_3477_n1454), .S(DP_OP_422J2_124_3477_n1455) );
  FADDX1_HVT DP_OP_422J2_124_3477_U909 ( .A(DP_OP_422J2_124_3477_n1507), .B(
        DP_OP_422J2_124_3477_n1638), .CI(DP_OP_422J2_124_3477_n1634), .CO(
        DP_OP_422J2_124_3477_n1452), .S(DP_OP_422J2_124_3477_n1453) );
  FADDX1_HVT DP_OP_422J2_124_3477_U908 ( .A(DP_OP_422J2_124_3477_n1624), .B(
        DP_OP_422J2_124_3477_n1487), .CI(DP_OP_422J2_124_3477_n1499), .CO(
        DP_OP_422J2_124_3477_n1450), .S(DP_OP_422J2_124_3477_n1451) );
  FADDX1_HVT DP_OP_422J2_124_3477_U907 ( .A(DP_OP_422J2_124_3477_n1632), .B(
        DP_OP_422J2_124_3477_n1501), .CI(DP_OP_422J2_124_3477_n1497), .CO(
        DP_OP_422J2_124_3477_n1448), .S(DP_OP_422J2_124_3477_n1449) );
  FADDX1_HVT DP_OP_422J2_124_3477_U906 ( .A(DP_OP_422J2_124_3477_n1630), .B(
        DP_OP_422J2_124_3477_n1489), .CI(DP_OP_422J2_124_3477_n1491), .CO(
        DP_OP_422J2_124_3477_n1446), .S(DP_OP_422J2_124_3477_n1447) );
  FADDX1_HVT DP_OP_422J2_124_3477_U905 ( .A(DP_OP_422J2_124_3477_n1628), .B(
        DP_OP_422J2_124_3477_n1495), .CI(DP_OP_422J2_124_3477_n1493), .CO(
        DP_OP_422J2_124_3477_n1444), .S(DP_OP_422J2_124_3477_n1445) );
  FADDX1_HVT DP_OP_422J2_124_3477_U904 ( .A(DP_OP_422J2_124_3477_n1626), .B(
        DP_OP_422J2_124_3477_n1622), .CI(DP_OP_422J2_124_3477_n1483), .CO(
        DP_OP_422J2_124_3477_n1442), .S(DP_OP_422J2_124_3477_n1443) );
  FADDX1_HVT DP_OP_422J2_124_3477_U903 ( .A(DP_OP_422J2_124_3477_n1485), .B(
        DP_OP_422J2_124_3477_n1481), .CI(DP_OP_422J2_124_3477_n1479), .CO(
        DP_OP_422J2_124_3477_n1440), .S(DP_OP_422J2_124_3477_n1441) );
  FADDX1_HVT DP_OP_422J2_124_3477_U902 ( .A(DP_OP_422J2_124_3477_n1620), .B(
        DP_OP_422J2_124_3477_n1471), .CI(DP_OP_422J2_124_3477_n1469), .CO(
        DP_OP_422J2_124_3477_n1438), .S(DP_OP_422J2_124_3477_n1439) );
  FADDX1_HVT DP_OP_422J2_124_3477_U901 ( .A(DP_OP_422J2_124_3477_n1475), .B(
        DP_OP_422J2_124_3477_n1465), .CI(DP_OP_422J2_124_3477_n1467), .CO(
        DP_OP_422J2_124_3477_n1436), .S(DP_OP_422J2_124_3477_n1437) );
  FADDX1_HVT DP_OP_422J2_124_3477_U900 ( .A(DP_OP_422J2_124_3477_n1473), .B(
        DP_OP_422J2_124_3477_n1477), .CI(DP_OP_422J2_124_3477_n1618), .CO(
        DP_OP_422J2_124_3477_n1434), .S(DP_OP_422J2_124_3477_n1435) );
  FADDX1_HVT DP_OP_422J2_124_3477_U899 ( .A(DP_OP_422J2_124_3477_n1616), .B(
        DP_OP_422J2_124_3477_n1463), .CI(DP_OP_422J2_124_3477_n1614), .CO(
        DP_OP_422J2_124_3477_n1432), .S(DP_OP_422J2_124_3477_n1433) );
  FADDX1_HVT DP_OP_422J2_124_3477_U898 ( .A(DP_OP_422J2_124_3477_n1461), .B(
        DP_OP_422J2_124_3477_n1459), .CI(DP_OP_422J2_124_3477_n1612), .CO(
        DP_OP_422J2_124_3477_n1430), .S(DP_OP_422J2_124_3477_n1431) );
  FADDX1_HVT DP_OP_422J2_124_3477_U897 ( .A(DP_OP_422J2_124_3477_n1610), .B(
        DP_OP_422J2_124_3477_n1606), .CI(DP_OP_422J2_124_3477_n1608), .CO(
        DP_OP_422J2_124_3477_n1428), .S(DP_OP_422J2_124_3477_n1429) );
  FADDX1_HVT DP_OP_422J2_124_3477_U896 ( .A(DP_OP_422J2_124_3477_n1457), .B(
        DP_OP_422J2_124_3477_n1604), .CI(DP_OP_422J2_124_3477_n1602), .CO(
        DP_OP_422J2_124_3477_n1426), .S(DP_OP_422J2_124_3477_n1427) );
  FADDX1_HVT DP_OP_422J2_124_3477_U895 ( .A(DP_OP_422J2_124_3477_n1455), .B(
        DP_OP_422J2_124_3477_n1453), .CI(DP_OP_422J2_124_3477_n1449), .CO(
        DP_OP_422J2_124_3477_n1424), .S(DP_OP_422J2_124_3477_n1425) );
  FADDX1_HVT DP_OP_422J2_124_3477_U894 ( .A(DP_OP_422J2_124_3477_n1451), .B(
        DP_OP_422J2_124_3477_n1447), .CI(DP_OP_422J2_124_3477_n1443), .CO(
        DP_OP_422J2_124_3477_n1422), .S(DP_OP_422J2_124_3477_n1423) );
  FADDX1_HVT DP_OP_422J2_124_3477_U893 ( .A(DP_OP_422J2_124_3477_n1600), .B(
        DP_OP_422J2_124_3477_n1445), .CI(DP_OP_422J2_124_3477_n1598), .CO(
        DP_OP_422J2_124_3477_n1420), .S(DP_OP_422J2_124_3477_n1421) );
  FADDX1_HVT DP_OP_422J2_124_3477_U892 ( .A(DP_OP_422J2_124_3477_n1441), .B(
        DP_OP_422J2_124_3477_n1439), .CI(DP_OP_422J2_124_3477_n1437), .CO(
        DP_OP_422J2_124_3477_n1418), .S(DP_OP_422J2_124_3477_n1419) );
  FADDX1_HVT DP_OP_422J2_124_3477_U891 ( .A(DP_OP_422J2_124_3477_n1596), .B(
        DP_OP_422J2_124_3477_n1435), .CI(DP_OP_422J2_124_3477_n1594), .CO(
        DP_OP_422J2_124_3477_n1416), .S(DP_OP_422J2_124_3477_n1417) );
  FADDX1_HVT DP_OP_422J2_124_3477_U889 ( .A(DP_OP_422J2_124_3477_n1429), .B(
        DP_OP_422J2_124_3477_n1431), .CI(DP_OP_422J2_124_3477_n1588), .CO(
        DP_OP_422J2_124_3477_n1412), .S(DP_OP_422J2_124_3477_n1413) );
  FADDX1_HVT DP_OP_422J2_124_3477_U888 ( .A(DP_OP_422J2_124_3477_n1427), .B(
        DP_OP_422J2_124_3477_n1425), .CI(DP_OP_422J2_124_3477_n1586), .CO(
        DP_OP_422J2_124_3477_n1410), .S(DP_OP_422J2_124_3477_n1411) );
  FADDX1_HVT DP_OP_422J2_124_3477_U887 ( .A(DP_OP_422J2_124_3477_n1421), .B(
        DP_OP_422J2_124_3477_n1423), .CI(DP_OP_422J2_124_3477_n1584), .CO(
        DP_OP_422J2_124_3477_n1408), .S(DP_OP_422J2_124_3477_n1409) );
  FADDX1_HVT DP_OP_422J2_124_3477_U886 ( .A(DP_OP_422J2_124_3477_n1419), .B(
        DP_OP_422J2_124_3477_n1417), .CI(DP_OP_422J2_124_3477_n1582), .CO(
        DP_OP_422J2_124_3477_n1406), .S(DP_OP_422J2_124_3477_n1407) );
  FADDX1_HVT DP_OP_422J2_124_3477_U885 ( .A(DP_OP_422J2_124_3477_n1415), .B(
        DP_OP_422J2_124_3477_n1580), .CI(DP_OP_422J2_124_3477_n1413), .CO(
        DP_OP_422J2_124_3477_n1404), .S(DP_OP_422J2_124_3477_n1405) );
  FADDX1_HVT DP_OP_422J2_124_3477_U884 ( .A(DP_OP_422J2_124_3477_n1411), .B(
        DP_OP_422J2_124_3477_n1578), .CI(DP_OP_422J2_124_3477_n1409), .CO(
        DP_OP_422J2_124_3477_n1402), .S(DP_OP_422J2_124_3477_n1403) );
  FADDX1_HVT DP_OP_422J2_124_3477_U883 ( .A(DP_OP_422J2_124_3477_n1407), .B(
        DP_OP_422J2_124_3477_n1576), .CI(DP_OP_422J2_124_3477_n1405), .CO(
        DP_OP_422J2_124_3477_n1400), .S(DP_OP_422J2_124_3477_n1401) );
  HADDX1_HVT DP_OP_422J2_124_3477_U882 ( .A0(DP_OP_422J2_124_3477_n3030), .B0(
        DP_OP_422J2_124_3477_n1975), .C1(DP_OP_422J2_124_3477_n1398), .SO(
        DP_OP_422J2_124_3477_n1399) );
  FADDX1_HVT DP_OP_422J2_124_3477_U881 ( .A(DP_OP_422J2_124_3477_n2503), .B(
        DP_OP_422J2_124_3477_n2415), .CI(DP_OP_422J2_124_3477_n1931), .CO(
        DP_OP_422J2_124_3477_n1396), .S(DP_OP_422J2_124_3477_n1397) );
  FADDX1_HVT DP_OP_422J2_124_3477_U880 ( .A(DP_OP_422J2_124_3477_n2547), .B(
        DP_OP_422J2_124_3477_n2327), .CI(DP_OP_422J2_124_3477_n2371), .CO(
        DP_OP_422J2_124_3477_n1394), .S(DP_OP_422J2_124_3477_n1395) );
  FADDX1_HVT DP_OP_422J2_124_3477_U879 ( .A(DP_OP_422J2_124_3477_n2855), .B(
        DP_OP_422J2_124_3477_n2019), .CI(DP_OP_422J2_124_3477_n2107), .CO(
        DP_OP_422J2_124_3477_n1392), .S(DP_OP_422J2_124_3477_n1393) );
  FADDX1_HVT DP_OP_422J2_124_3477_U878 ( .A(DP_OP_422J2_124_3477_n2591), .B(
        DP_OP_422J2_124_3477_n2151), .CI(DP_OP_422J2_124_3477_n2679), .CO(
        DP_OP_422J2_124_3477_n1390), .S(DP_OP_422J2_124_3477_n1391) );
  FADDX1_HVT DP_OP_422J2_124_3477_U877 ( .A(DP_OP_422J2_124_3477_n2063), .B(
        DP_OP_422J2_124_3477_n2899), .CI(DP_OP_422J2_124_3477_n2195), .CO(
        DP_OP_422J2_124_3477_n1388), .S(DP_OP_422J2_124_3477_n1389) );
  FADDX1_HVT DP_OP_422J2_124_3477_U876 ( .A(DP_OP_422J2_124_3477_n2459), .B(
        DP_OP_422J2_124_3477_n2943), .CI(DP_OP_422J2_124_3477_n2767), .CO(
        DP_OP_422J2_124_3477_n1386), .S(DP_OP_422J2_124_3477_n1387) );
  FADDX1_HVT DP_OP_422J2_124_3477_U875 ( .A(DP_OP_422J2_124_3477_n2283), .B(
        DP_OP_422J2_124_3477_n2239), .CI(DP_OP_422J2_124_3477_n2723), .CO(
        DP_OP_422J2_124_3477_n1384), .S(DP_OP_422J2_124_3477_n1385) );
  FADDX1_HVT DP_OP_422J2_124_3477_U874 ( .A(DP_OP_422J2_124_3477_n2987), .B(
        DP_OP_422J2_124_3477_n2635), .CI(DP_OP_422J2_124_3477_n2811), .CO(
        DP_OP_422J2_124_3477_n1382), .S(DP_OP_422J2_124_3477_n1383) );
  FADDX1_HVT DP_OP_422J2_124_3477_U873 ( .A(DP_OP_422J2_124_3477_n2429), .B(
        DP_OP_422J2_124_3477_n3050), .CI(DP_OP_422J2_124_3477_n1982), .CO(
        DP_OP_422J2_124_3477_n1380), .S(DP_OP_422J2_124_3477_n1381) );
  FADDX1_HVT DP_OP_422J2_124_3477_U872 ( .A(DP_OP_422J2_124_3477_n2422), .B(
        DP_OP_422J2_124_3477_n1989), .CI(DP_OP_422J2_124_3477_n1996), .CO(
        DP_OP_422J2_124_3477_n1378), .S(DP_OP_422J2_124_3477_n1379) );
  FADDX1_HVT DP_OP_422J2_124_3477_U871 ( .A(DP_OP_422J2_124_3477_n2436), .B(
        DP_OP_422J2_124_3477_n2026), .CI(DP_OP_422J2_124_3477_n3043), .CO(
        DP_OP_422J2_124_3477_n1376), .S(DP_OP_422J2_124_3477_n1377) );
  FADDX1_HVT DP_OP_422J2_124_3477_U870 ( .A(DP_OP_422J2_124_3477_n2392), .B(
        DP_OP_422J2_124_3477_n3036), .CI(DP_OP_422J2_124_3477_n3008), .CO(
        DP_OP_422J2_124_3477_n1374), .S(DP_OP_422J2_124_3477_n1375) );
  FADDX1_HVT DP_OP_422J2_124_3477_U869 ( .A(DP_OP_422J2_124_3477_n2385), .B(
        DP_OP_422J2_124_3477_n3001), .CI(DP_OP_422J2_124_3477_n2994), .CO(
        DP_OP_422J2_124_3477_n1372), .S(DP_OP_422J2_124_3477_n1373) );
  FADDX1_HVT DP_OP_422J2_124_3477_U868 ( .A(DP_OP_422J2_124_3477_n2348), .B(
        DP_OP_422J2_124_3477_n2964), .CI(DP_OP_422J2_124_3477_n2957), .CO(
        DP_OP_422J2_124_3477_n1370), .S(DP_OP_422J2_124_3477_n1371) );
  FADDX1_HVT DP_OP_422J2_124_3477_U867 ( .A(DP_OP_422J2_124_3477_n2341), .B(
        DP_OP_422J2_124_3477_n2033), .CI(DP_OP_422J2_124_3477_n2950), .CO(
        DP_OP_422J2_124_3477_n1368), .S(DP_OP_422J2_124_3477_n1369) );
  FADDX1_HVT DP_OP_422J2_124_3477_U866 ( .A(DP_OP_422J2_124_3477_n2334), .B(
        DP_OP_422J2_124_3477_n2920), .CI(DP_OP_422J2_124_3477_n2913), .CO(
        DP_OP_422J2_124_3477_n1366), .S(DP_OP_422J2_124_3477_n1367) );
  FADDX1_HVT DP_OP_422J2_124_3477_U865 ( .A(DP_OP_422J2_124_3477_n2304), .B(
        DP_OP_422J2_124_3477_n2906), .CI(DP_OP_422J2_124_3477_n2040), .CO(
        DP_OP_422J2_124_3477_n1364), .S(DP_OP_422J2_124_3477_n1365) );
  FADDX1_HVT DP_OP_422J2_124_3477_U864 ( .A(DP_OP_422J2_124_3477_n2297), .B(
        DP_OP_422J2_124_3477_n2070), .CI(DP_OP_422J2_124_3477_n2077), .CO(
        DP_OP_422J2_124_3477_n1362), .S(DP_OP_422J2_124_3477_n1363) );
  FADDX1_HVT DP_OP_422J2_124_3477_U863 ( .A(DP_OP_422J2_124_3477_n2378), .B(
        DP_OP_422J2_124_3477_n2084), .CI(DP_OP_422J2_124_3477_n2876), .CO(
        DP_OP_422J2_124_3477_n1360), .S(DP_OP_422J2_124_3477_n1361) );
  FADDX1_HVT DP_OP_422J2_124_3477_U862 ( .A(DP_OP_422J2_124_3477_n2466), .B(
        DP_OP_422J2_124_3477_n2869), .CI(DP_OP_422J2_124_3477_n2114), .CO(
        DP_OP_422J2_124_3477_n1358), .S(DP_OP_422J2_124_3477_n1359) );
  FADDX1_HVT DP_OP_422J2_124_3477_U861 ( .A(DP_OP_422J2_124_3477_n2862), .B(
        DP_OP_422J2_124_3477_n2121), .CI(DP_OP_422J2_124_3477_n2128), .CO(
        DP_OP_422J2_124_3477_n1356), .S(DP_OP_422J2_124_3477_n1357) );
  FADDX1_HVT DP_OP_422J2_124_3477_U860 ( .A(DP_OP_422J2_124_3477_n2832), .B(
        DP_OP_422J2_124_3477_n2158), .CI(DP_OP_422J2_124_3477_n2165), .CO(
        DP_OP_422J2_124_3477_n1354), .S(DP_OP_422J2_124_3477_n1355) );
  FADDX1_HVT DP_OP_422J2_124_3477_U859 ( .A(DP_OP_422J2_124_3477_n2825), .B(
        DP_OP_422J2_124_3477_n2172), .CI(DP_OP_422J2_124_3477_n2202), .CO(
        DP_OP_422J2_124_3477_n1352), .S(DP_OP_422J2_124_3477_n1353) );
  FADDX1_HVT DP_OP_422J2_124_3477_U858 ( .A(DP_OP_422J2_124_3477_n2818), .B(
        DP_OP_422J2_124_3477_n2209), .CI(DP_OP_422J2_124_3477_n2216), .CO(
        DP_OP_422J2_124_3477_n1350), .S(DP_OP_422J2_124_3477_n1351) );
  FADDX1_HVT DP_OP_422J2_124_3477_U857 ( .A(DP_OP_422J2_124_3477_n2788), .B(
        DP_OP_422J2_124_3477_n2246), .CI(DP_OP_422J2_124_3477_n2253), .CO(
        DP_OP_422J2_124_3477_n1348), .S(DP_OP_422J2_124_3477_n1349) );
  FADDX1_HVT DP_OP_422J2_124_3477_U856 ( .A(DP_OP_422J2_124_3477_n2781), .B(
        DP_OP_422J2_124_3477_n2260), .CI(DP_OP_422J2_124_3477_n2290), .CO(
        DP_OP_422J2_124_3477_n1346), .S(DP_OP_422J2_124_3477_n1347) );
  FADDX1_HVT DP_OP_422J2_124_3477_U855 ( .A(DP_OP_422J2_124_3477_n2774), .B(
        DP_OP_422J2_124_3477_n2473), .CI(DP_OP_422J2_124_3477_n2480), .CO(
        DP_OP_422J2_124_3477_n1344), .S(DP_OP_422J2_124_3477_n1345) );
  FADDX1_HVT DP_OP_422J2_124_3477_U854 ( .A(DP_OP_422J2_124_3477_n2744), .B(
        DP_OP_422J2_124_3477_n2510), .CI(DP_OP_422J2_124_3477_n2517), .CO(
        DP_OP_422J2_124_3477_n1342), .S(DP_OP_422J2_124_3477_n1343) );
  FADDX1_HVT DP_OP_422J2_124_3477_U853 ( .A(DP_OP_422J2_124_3477_n2737), .B(
        DP_OP_422J2_124_3477_n2524), .CI(DP_OP_422J2_124_3477_n2554), .CO(
        DP_OP_422J2_124_3477_n1340), .S(DP_OP_422J2_124_3477_n1341) );
  FADDX1_HVT DP_OP_422J2_124_3477_U852 ( .A(DP_OP_422J2_124_3477_n2730), .B(
        DP_OP_422J2_124_3477_n2561), .CI(DP_OP_422J2_124_3477_n2568), .CO(
        DP_OP_422J2_124_3477_n1338), .S(DP_OP_422J2_124_3477_n1339) );
  FADDX1_HVT DP_OP_422J2_124_3477_U851 ( .A(DP_OP_422J2_124_3477_n2700), .B(
        DP_OP_422J2_124_3477_n2693), .CI(DP_OP_422J2_124_3477_n2686), .CO(
        DP_OP_422J2_124_3477_n1336), .S(DP_OP_422J2_124_3477_n1337) );
  FADDX1_HVT DP_OP_422J2_124_3477_U850 ( .A(DP_OP_422J2_124_3477_n2642), .B(
        DP_OP_422J2_124_3477_n2656), .CI(DP_OP_422J2_124_3477_n2598), .CO(
        DP_OP_422J2_124_3477_n1334), .S(DP_OP_422J2_124_3477_n1335) );
  FADDX1_HVT DP_OP_422J2_124_3477_U848 ( .A(DP_OP_422J2_124_3477_n1399), .B(
        DP_OP_422J2_124_3477_n1574), .CI(DP_OP_422J2_124_3477_n1564), .CO(
        DP_OP_422J2_124_3477_n1330), .S(DP_OP_422J2_124_3477_n1331) );
  FADDX1_HVT DP_OP_422J2_124_3477_U847 ( .A(DP_OP_422J2_124_3477_n1572), .B(
        DP_OP_422J2_124_3477_n1570), .CI(DP_OP_422J2_124_3477_n1568), .CO(
        DP_OP_422J2_124_3477_n1328), .S(DP_OP_422J2_124_3477_n1329) );
  FADDX1_HVT DP_OP_422J2_124_3477_U846 ( .A(DP_OP_422J2_124_3477_n1566), .B(
        DP_OP_422J2_124_3477_n1562), .CI(DP_OP_422J2_124_3477_n1558), .CO(
        DP_OP_422J2_124_3477_n1326), .S(DP_OP_422J2_124_3477_n1327) );
  FADDX1_HVT DP_OP_422J2_124_3477_U845 ( .A(DP_OP_422J2_124_3477_n1560), .B(
        DP_OP_422J2_124_3477_n1534), .CI(DP_OP_422J2_124_3477_n1532), .CO(
        DP_OP_422J2_124_3477_n1324), .S(DP_OP_422J2_124_3477_n1325) );
  FADDX1_HVT DP_OP_422J2_124_3477_U844 ( .A(DP_OP_422J2_124_3477_n1536), .B(
        DP_OP_422J2_124_3477_n1508), .CI(DP_OP_422J2_124_3477_n1556), .CO(
        DP_OP_422J2_124_3477_n1322), .S(DP_OP_422J2_124_3477_n1323) );
  FADDX1_HVT DP_OP_422J2_124_3477_U843 ( .A(DP_OP_422J2_124_3477_n1528), .B(
        DP_OP_422J2_124_3477_n1554), .CI(DP_OP_422J2_124_3477_n1552), .CO(
        DP_OP_422J2_124_3477_n1320), .S(DP_OP_422J2_124_3477_n1321) );
  FADDX1_HVT DP_OP_422J2_124_3477_U842 ( .A(DP_OP_422J2_124_3477_n1548), .B(
        DP_OP_422J2_124_3477_n1524), .CI(DP_OP_422J2_124_3477_n1550), .CO(
        DP_OP_422J2_124_3477_n1318), .S(DP_OP_422J2_124_3477_n1319) );
  FADDX1_HVT DP_OP_422J2_124_3477_U841 ( .A(DP_OP_422J2_124_3477_n1518), .B(
        DP_OP_422J2_124_3477_n1510), .CI(DP_OP_422J2_124_3477_n1512), .CO(
        DP_OP_422J2_124_3477_n1316), .S(DP_OP_422J2_124_3477_n1317) );
  FADDX1_HVT DP_OP_422J2_124_3477_U840 ( .A(DP_OP_422J2_124_3477_n1516), .B(
        DP_OP_422J2_124_3477_n1546), .CI(DP_OP_422J2_124_3477_n1544), .CO(
        DP_OP_422J2_124_3477_n1314), .S(DP_OP_422J2_124_3477_n1315) );
  FADDX1_HVT DP_OP_422J2_124_3477_U839 ( .A(DP_OP_422J2_124_3477_n1526), .B(
        DP_OP_422J2_124_3477_n1542), .CI(DP_OP_422J2_124_3477_n1514), .CO(
        DP_OP_422J2_124_3477_n1312), .S(DP_OP_422J2_124_3477_n1313) );
  FADDX1_HVT DP_OP_422J2_124_3477_U838 ( .A(DP_OP_422J2_124_3477_n1522), .B(
        DP_OP_422J2_124_3477_n1540), .CI(DP_OP_422J2_124_3477_n1538), .CO(
        DP_OP_422J2_124_3477_n1310), .S(DP_OP_422J2_124_3477_n1311) );
  FADDX1_HVT DP_OP_422J2_124_3477_U837 ( .A(DP_OP_422J2_124_3477_n1520), .B(
        DP_OP_422J2_124_3477_n1530), .CI(DP_OP_422J2_124_3477_n1389), .CO(
        DP_OP_422J2_124_3477_n1308), .S(DP_OP_422J2_124_3477_n1309) );
  FADDX1_HVT DP_OP_422J2_124_3477_U836 ( .A(DP_OP_422J2_124_3477_n1391), .B(
        DP_OP_422J2_124_3477_n1383), .CI(DP_OP_422J2_124_3477_n1385), .CO(
        DP_OP_422J2_124_3477_n1306), .S(DP_OP_422J2_124_3477_n1307) );
  FADDX1_HVT DP_OP_422J2_124_3477_U835 ( .A(DP_OP_422J2_124_3477_n1395), .B(
        DP_OP_422J2_124_3477_n1393), .CI(DP_OP_422J2_124_3477_n1397), .CO(
        DP_OP_422J2_124_3477_n1304), .S(DP_OP_422J2_124_3477_n1305) );
  FADDX1_HVT DP_OP_422J2_124_3477_U834 ( .A(DP_OP_422J2_124_3477_n1387), .B(
        DP_OP_422J2_124_3477_n1339), .CI(DP_OP_422J2_124_3477_n1337), .CO(
        DP_OP_422J2_124_3477_n1302), .S(DP_OP_422J2_124_3477_n1303) );
  FADDX1_HVT DP_OP_422J2_124_3477_U833 ( .A(DP_OP_422J2_124_3477_n1333), .B(
        DP_OP_422J2_124_3477_n1381), .CI(DP_OP_422J2_124_3477_n1379), .CO(
        DP_OP_422J2_124_3477_n1300), .S(DP_OP_422J2_124_3477_n1301) );
  FADDX1_HVT DP_OP_422J2_124_3477_U832 ( .A(DP_OP_422J2_124_3477_n1369), .B(
        DP_OP_422J2_124_3477_n1359), .CI(DP_OP_422J2_124_3477_n1365), .CO(
        DP_OP_422J2_124_3477_n1298), .S(DP_OP_422J2_124_3477_n1299) );
  FADDX1_HVT DP_OP_422J2_124_3477_U831 ( .A(DP_OP_422J2_124_3477_n1363), .B(
        DP_OP_422J2_124_3477_n1361), .CI(DP_OP_422J2_124_3477_n1345), .CO(
        DP_OP_422J2_124_3477_n1296), .S(DP_OP_422J2_124_3477_n1297) );
  FADDX1_HVT DP_OP_422J2_124_3477_U830 ( .A(DP_OP_422J2_124_3477_n1367), .B(
        DP_OP_422J2_124_3477_n1341), .CI(DP_OP_422J2_124_3477_n1335), .CO(
        DP_OP_422J2_124_3477_n1294), .S(DP_OP_422J2_124_3477_n1295) );
  FADDX1_HVT DP_OP_422J2_124_3477_U829 ( .A(DP_OP_422J2_124_3477_n1371), .B(
        DP_OP_422J2_124_3477_n1353), .CI(DP_OP_422J2_124_3477_n1355), .CO(
        DP_OP_422J2_124_3477_n1292), .S(DP_OP_422J2_124_3477_n1293) );
  FADDX1_HVT DP_OP_422J2_124_3477_U828 ( .A(DP_OP_422J2_124_3477_n1351), .B(
        DP_OP_422J2_124_3477_n1349), .CI(DP_OP_422J2_124_3477_n1343), .CO(
        DP_OP_422J2_124_3477_n1290), .S(DP_OP_422J2_124_3477_n1291) );
  FADDX1_HVT DP_OP_422J2_124_3477_U827 ( .A(DP_OP_422J2_124_3477_n1347), .B(
        DP_OP_422J2_124_3477_n1377), .CI(DP_OP_422J2_124_3477_n1373), .CO(
        DP_OP_422J2_124_3477_n1288), .S(DP_OP_422J2_124_3477_n1289) );
  FADDX1_HVT DP_OP_422J2_124_3477_U826 ( .A(DP_OP_422J2_124_3477_n1375), .B(
        DP_OP_422J2_124_3477_n1357), .CI(DP_OP_422J2_124_3477_n1506), .CO(
        DP_OP_422J2_124_3477_n1286), .S(DP_OP_422J2_124_3477_n1287) );
  FADDX1_HVT DP_OP_422J2_124_3477_U825 ( .A(DP_OP_422J2_124_3477_n1504), .B(
        DP_OP_422J2_124_3477_n1502), .CI(DP_OP_422J2_124_3477_n1500), .CO(
        DP_OP_422J2_124_3477_n1284), .S(DP_OP_422J2_124_3477_n1285) );
  FADDX1_HVT DP_OP_422J2_124_3477_U823 ( .A(DP_OP_422J2_124_3477_n1492), .B(
        DP_OP_422J2_124_3477_n1496), .CI(DP_OP_422J2_124_3477_n1490), .CO(
        DP_OP_422J2_124_3477_n1280), .S(DP_OP_422J2_124_3477_n1281) );
  FADDX1_HVT DP_OP_422J2_124_3477_U822 ( .A(DP_OP_422J2_124_3477_n1494), .B(
        DP_OP_422J2_124_3477_n1331), .CI(DP_OP_422J2_124_3477_n1484), .CO(
        DP_OP_422J2_124_3477_n1278), .S(DP_OP_422J2_124_3477_n1279) );
  FADDX1_HVT DP_OP_422J2_124_3477_U821 ( .A(DP_OP_422J2_124_3477_n1329), .B(
        DP_OP_422J2_124_3477_n1327), .CI(DP_OP_422J2_124_3477_n1325), .CO(
        DP_OP_422J2_124_3477_n1276), .S(DP_OP_422J2_124_3477_n1277) );
  FADDX1_HVT DP_OP_422J2_124_3477_U820 ( .A(DP_OP_422J2_124_3477_n1482), .B(
        DP_OP_422J2_124_3477_n1480), .CI(DP_OP_422J2_124_3477_n1478), .CO(
        DP_OP_422J2_124_3477_n1274), .S(DP_OP_422J2_124_3477_n1275) );
  FADDX1_HVT DP_OP_422J2_124_3477_U819 ( .A(DP_OP_422J2_124_3477_n1466), .B(
        DP_OP_422J2_124_3477_n1311), .CI(DP_OP_422J2_124_3477_n1309), .CO(
        DP_OP_422J2_124_3477_n1272), .S(DP_OP_422J2_124_3477_n1273) );
  FADDX1_HVT DP_OP_422J2_124_3477_U818 ( .A(DP_OP_422J2_124_3477_n1476), .B(
        DP_OP_422J2_124_3477_n1321), .CI(DP_OP_422J2_124_3477_n1323), .CO(
        DP_OP_422J2_124_3477_n1270), .S(DP_OP_422J2_124_3477_n1271) );
  FADDX1_HVT DP_OP_422J2_124_3477_U817 ( .A(DP_OP_422J2_124_3477_n1474), .B(
        DP_OP_422J2_124_3477_n1317), .CI(DP_OP_422J2_124_3477_n1313), .CO(
        DP_OP_422J2_124_3477_n1268), .S(DP_OP_422J2_124_3477_n1269) );
  FADDX1_HVT DP_OP_422J2_124_3477_U816 ( .A(DP_OP_422J2_124_3477_n1472), .B(
        DP_OP_422J2_124_3477_n1319), .CI(DP_OP_422J2_124_3477_n1315), .CO(
        DP_OP_422J2_124_3477_n1266), .S(DP_OP_422J2_124_3477_n1267) );
  FADDX1_HVT DP_OP_422J2_124_3477_U815 ( .A(DP_OP_422J2_124_3477_n1470), .B(
        DP_OP_422J2_124_3477_n1464), .CI(DP_OP_422J2_124_3477_n1468), .CO(
        DP_OP_422J2_124_3477_n1264), .S(DP_OP_422J2_124_3477_n1265) );
  FADDX1_HVT DP_OP_422J2_124_3477_U814 ( .A(DP_OP_422J2_124_3477_n1305), .B(
        DP_OP_422J2_124_3477_n1307), .CI(DP_OP_422J2_124_3477_n1303), .CO(
        DP_OP_422J2_124_3477_n1262), .S(DP_OP_422J2_124_3477_n1263) );
  FADDX1_HVT DP_OP_422J2_124_3477_U813 ( .A(DP_OP_422J2_124_3477_n1295), .B(
        DP_OP_422J2_124_3477_n1297), .CI(DP_OP_422J2_124_3477_n1462), .CO(
        DP_OP_422J2_124_3477_n1260), .S(DP_OP_422J2_124_3477_n1261) );
  FADDX1_HVT DP_OP_422J2_124_3477_U812 ( .A(DP_OP_422J2_124_3477_n1293), .B(
        DP_OP_422J2_124_3477_n1301), .CI(DP_OP_422J2_124_3477_n1299), .CO(
        DP_OP_422J2_124_3477_n1258), .S(DP_OP_422J2_124_3477_n1259) );
  FADDX1_HVT DP_OP_422J2_124_3477_U810 ( .A(DP_OP_422J2_124_3477_n1287), .B(
        DP_OP_422J2_124_3477_n1460), .CI(DP_OP_422J2_124_3477_n1456), .CO(
        DP_OP_422J2_124_3477_n1254), .S(DP_OP_422J2_124_3477_n1255) );
  FADDX1_HVT DP_OP_422J2_124_3477_U809 ( .A(DP_OP_422J2_124_3477_n1285), .B(
        DP_OP_422J2_124_3477_n1452), .CI(DP_OP_422J2_124_3477_n1454), .CO(
        DP_OP_422J2_124_3477_n1252), .S(DP_OP_422J2_124_3477_n1253) );
  FADDX1_HVT DP_OP_422J2_124_3477_U808 ( .A(DP_OP_422J2_124_3477_n1450), .B(
        DP_OP_422J2_124_3477_n1442), .CI(DP_OP_422J2_124_3477_n1279), .CO(
        DP_OP_422J2_124_3477_n1250), .S(DP_OP_422J2_124_3477_n1251) );
  FADDX1_HVT DP_OP_422J2_124_3477_U806 ( .A(DP_OP_422J2_124_3477_n1446), .B(
        DP_OP_422J2_124_3477_n1444), .CI(DP_OP_422J2_124_3477_n1440), .CO(
        DP_OP_422J2_124_3477_n1246), .S(DP_OP_422J2_124_3477_n1247) );
  FADDX1_HVT DP_OP_422J2_124_3477_U805 ( .A(DP_OP_422J2_124_3477_n1275), .B(
        DP_OP_422J2_124_3477_n1277), .CI(DP_OP_422J2_124_3477_n1438), .CO(
        DP_OP_422J2_124_3477_n1244), .S(DP_OP_422J2_124_3477_n1245) );
  FADDX1_HVT DP_OP_422J2_124_3477_U804 ( .A(DP_OP_422J2_124_3477_n1436), .B(
        DP_OP_422J2_124_3477_n1269), .CI(DP_OP_422J2_124_3477_n1434), .CO(
        DP_OP_422J2_124_3477_n1242), .S(DP_OP_422J2_124_3477_n1243) );
  FADDX1_HVT DP_OP_422J2_124_3477_U803 ( .A(DP_OP_422J2_124_3477_n1267), .B(
        DP_OP_422J2_124_3477_n1273), .CI(DP_OP_422J2_124_3477_n1271), .CO(
        DP_OP_422J2_124_3477_n1240), .S(DP_OP_422J2_124_3477_n1241) );
  FADDX1_HVT DP_OP_422J2_124_3477_U802 ( .A(DP_OP_422J2_124_3477_n1265), .B(
        DP_OP_422J2_124_3477_n1263), .CI(DP_OP_422J2_124_3477_n1259), .CO(
        DP_OP_422J2_124_3477_n1238), .S(DP_OP_422J2_124_3477_n1239) );
  FADDX1_HVT DP_OP_422J2_124_3477_U801 ( .A(DP_OP_422J2_124_3477_n1261), .B(
        DP_OP_422J2_124_3477_n1432), .CI(DP_OP_422J2_124_3477_n1257), .CO(
        DP_OP_422J2_124_3477_n1236), .S(DP_OP_422J2_124_3477_n1237) );
  FADDX1_HVT DP_OP_422J2_124_3477_U800 ( .A(DP_OP_422J2_124_3477_n1430), .B(
        DP_OP_422J2_124_3477_n1428), .CI(DP_OP_422J2_124_3477_n1255), .CO(
        DP_OP_422J2_124_3477_n1234), .S(DP_OP_422J2_124_3477_n1235) );
  FADDX1_HVT DP_OP_422J2_124_3477_U799 ( .A(DP_OP_422J2_124_3477_n1426), .B(
        DP_OP_422J2_124_3477_n1424), .CI(DP_OP_422J2_124_3477_n1253), .CO(
        DP_OP_422J2_124_3477_n1232), .S(DP_OP_422J2_124_3477_n1233) );
  FADDX1_HVT DP_OP_422J2_124_3477_U798 ( .A(DP_OP_422J2_124_3477_n1422), .B(
        DP_OP_422J2_124_3477_n1249), .CI(DP_OP_422J2_124_3477_n1247), .CO(
        DP_OP_422J2_124_3477_n1230), .S(DP_OP_422J2_124_3477_n1231) );
  FADDX1_HVT DP_OP_422J2_124_3477_U797 ( .A(DP_OP_422J2_124_3477_n1420), .B(
        DP_OP_422J2_124_3477_n1251), .CI(DP_OP_422J2_124_3477_n1245), .CO(
        DP_OP_422J2_124_3477_n1228), .S(DP_OP_422J2_124_3477_n1229) );
  FADDX1_HVT DP_OP_422J2_124_3477_U796 ( .A(DP_OP_422J2_124_3477_n1418), .B(
        DP_OP_422J2_124_3477_n1241), .CI(DP_OP_422J2_124_3477_n1416), .CO(
        DP_OP_422J2_124_3477_n1226), .S(DP_OP_422J2_124_3477_n1227) );
  FADDX1_HVT DP_OP_422J2_124_3477_U795 ( .A(DP_OP_422J2_124_3477_n1243), .B(
        DP_OP_422J2_124_3477_n1239), .CI(DP_OP_422J2_124_3477_n1237), .CO(
        DP_OP_422J2_124_3477_n1224), .S(DP_OP_422J2_124_3477_n1225) );
  FADDX1_HVT DP_OP_422J2_124_3477_U794 ( .A(DP_OP_422J2_124_3477_n1414), .B(
        DP_OP_422J2_124_3477_n1235), .CI(DP_OP_422J2_124_3477_n1412), .CO(
        DP_OP_422J2_124_3477_n1222), .S(DP_OP_422J2_124_3477_n1223) );
  FADDX1_HVT DP_OP_422J2_124_3477_U793 ( .A(DP_OP_422J2_124_3477_n1410), .B(
        DP_OP_422J2_124_3477_n1233), .CI(DP_OP_422J2_124_3477_n1231), .CO(
        DP_OP_422J2_124_3477_n1220), .S(DP_OP_422J2_124_3477_n1221) );
  FADDX1_HVT DP_OP_422J2_124_3477_U792 ( .A(DP_OP_422J2_124_3477_n1229), .B(
        DP_OP_422J2_124_3477_n1408), .CI(DP_OP_422J2_124_3477_n1227), .CO(
        DP_OP_422J2_124_3477_n1218), .S(DP_OP_422J2_124_3477_n1219) );
  FADDX1_HVT DP_OP_422J2_124_3477_U791 ( .A(DP_OP_422J2_124_3477_n1406), .B(n5), .CI(DP_OP_422J2_124_3477_n1404), .CO(DP_OP_422J2_124_3477_n1216), .S(
        DP_OP_422J2_124_3477_n1217) );
  FADDX1_HVT DP_OP_422J2_124_3477_U790 ( .A(DP_OP_422J2_124_3477_n1223), .B(
        DP_OP_422J2_124_3477_n1221), .CI(DP_OP_422J2_124_3477_n1402), .CO(
        DP_OP_422J2_124_3477_n1214), .S(DP_OP_422J2_124_3477_n1215) );
  FADDX1_HVT DP_OP_422J2_124_3477_U786 ( .A(DP_OP_422J2_124_3477_n2194), .B(
        DP_OP_422J2_124_3477_n1974), .CI(DP_OP_422J2_124_3477_n1930), .CO(
        DP_OP_422J2_124_3477_n1208), .S(DP_OP_422J2_124_3477_n1209) );
  FADDX1_HVT DP_OP_422J2_124_3477_U785 ( .A(DP_OP_422J2_124_3477_n2634), .B(
        DP_OP_422J2_124_3477_n2062), .CI(DP_OP_422J2_124_3477_n2414), .CO(
        DP_OP_422J2_124_3477_n1206), .S(DP_OP_422J2_124_3477_n1207) );
  FADDX1_HVT DP_OP_422J2_124_3477_U784 ( .A(DP_OP_422J2_124_3477_n2854), .B(
        DP_OP_422J2_124_3477_n2678), .CI(DP_OP_422J2_124_3477_n2238), .CO(
        DP_OP_422J2_124_3477_n1204), .S(DP_OP_422J2_124_3477_n1205) );
  FADDX1_HVT DP_OP_422J2_124_3477_U783 ( .A(DP_OP_422J2_124_3477_n2326), .B(
        DP_OP_422J2_124_3477_n2150), .CI(DP_OP_422J2_124_3477_n2898), .CO(
        DP_OP_422J2_124_3477_n1202), .S(DP_OP_422J2_124_3477_n1203) );
  FADDX1_HVT DP_OP_422J2_124_3477_U782 ( .A(DP_OP_422J2_124_3477_n2458), .B(
        DP_OP_422J2_124_3477_n2722), .CI(DP_OP_422J2_124_3477_n2942), .CO(
        DP_OP_422J2_124_3477_n1200), .S(DP_OP_422J2_124_3477_n1201) );
  FADDX1_HVT DP_OP_422J2_124_3477_U781 ( .A(DP_OP_422J2_124_3477_n2546), .B(
        DP_OP_422J2_124_3477_n2766), .CI(DP_OP_422J2_124_3477_n2590), .CO(
        DP_OP_422J2_124_3477_n1198), .S(DP_OP_422J2_124_3477_n1199) );
  FADDX1_HVT DP_OP_422J2_124_3477_U780 ( .A(DP_OP_422J2_124_3477_n2282), .B(
        DP_OP_422J2_124_3477_n2106), .CI(DP_OP_422J2_124_3477_n2986), .CO(
        DP_OP_422J2_124_3477_n1196), .S(DP_OP_422J2_124_3477_n1197) );
  FADDX1_HVT DP_OP_422J2_124_3477_U779 ( .A(DP_OP_422J2_124_3477_n2810), .B(
        DP_OP_422J2_124_3477_n2018), .CI(DP_OP_422J2_124_3477_n2370), .CO(
        DP_OP_422J2_124_3477_n1194), .S(DP_OP_422J2_124_3477_n1195) );
  FADDX1_HVT DP_OP_422J2_124_3477_U778 ( .A(DP_OP_422J2_124_3477_n2421), .B(
        DP_OP_422J2_124_3477_n3049), .CI(DP_OP_422J2_124_3477_n1981), .CO(
        DP_OP_422J2_124_3477_n1192), .S(DP_OP_422J2_124_3477_n1193) );
  FADDX1_HVT DP_OP_422J2_124_3477_U777 ( .A(DP_OP_422J2_124_3477_n2428), .B(
        DP_OP_422J2_124_3477_n3042), .CI(DP_OP_422J2_124_3477_n3035), .CO(
        DP_OP_422J2_124_3477_n1190), .S(DP_OP_422J2_124_3477_n1191) );
  FADDX1_HVT DP_OP_422J2_124_3477_U776 ( .A(DP_OP_422J2_124_3477_n2384), .B(
        DP_OP_422J2_124_3477_n3007), .CI(DP_OP_422J2_124_3477_n3000), .CO(
        DP_OP_422J2_124_3477_n1188), .S(DP_OP_422J2_124_3477_n1189) );
  FADDX1_HVT DP_OP_422J2_124_3477_U775 ( .A(DP_OP_422J2_124_3477_n2347), .B(
        DP_OP_422J2_124_3477_n2993), .CI(DP_OP_422J2_124_3477_n2963), .CO(
        DP_OP_422J2_124_3477_n1186), .S(DP_OP_422J2_124_3477_n1187) );
  FADDX1_HVT DP_OP_422J2_124_3477_U774 ( .A(DP_OP_422J2_124_3477_n2340), .B(
        DP_OP_422J2_124_3477_n1988), .CI(DP_OP_422J2_124_3477_n2956), .CO(
        DP_OP_422J2_124_3477_n1184), .S(DP_OP_422J2_124_3477_n1185) );
  FADDX1_HVT DP_OP_422J2_124_3477_U773 ( .A(DP_OP_422J2_124_3477_n2377), .B(
        DP_OP_422J2_124_3477_n2949), .CI(DP_OP_422J2_124_3477_n1995), .CO(
        DP_OP_422J2_124_3477_n1182), .S(DP_OP_422J2_124_3477_n1183) );
  FADDX1_HVT DP_OP_422J2_124_3477_U772 ( .A(DP_OP_422J2_124_3477_n2333), .B(
        DP_OP_422J2_124_3477_n2919), .CI(DP_OP_422J2_124_3477_n2025), .CO(
        DP_OP_422J2_124_3477_n1180), .S(DP_OP_422J2_124_3477_n1181) );
  FADDX1_HVT DP_OP_422J2_124_3477_U771 ( .A(DP_OP_422J2_124_3477_n2303), .B(
        DP_OP_422J2_124_3477_n2912), .CI(DP_OP_422J2_124_3477_n2905), .CO(
        DP_OP_422J2_124_3477_n1178), .S(DP_OP_422J2_124_3477_n1179) );
  FADDX1_HVT DP_OP_422J2_124_3477_U770 ( .A(DP_OP_422J2_124_3477_n2296), .B(
        DP_OP_422J2_124_3477_n2032), .CI(DP_OP_422J2_124_3477_n2875), .CO(
        DP_OP_422J2_124_3477_n1176), .S(DP_OP_422J2_124_3477_n1177) );
  FADDX1_HVT DP_OP_422J2_124_3477_U769 ( .A(DP_OP_422J2_124_3477_n2289), .B(
        DP_OP_422J2_124_3477_n2039), .CI(DP_OP_422J2_124_3477_n2868), .CO(
        DP_OP_422J2_124_3477_n1174), .S(DP_OP_422J2_124_3477_n1175) );
  FADDX1_HVT DP_OP_422J2_124_3477_U768 ( .A(DP_OP_422J2_124_3477_n2069), .B(
        DP_OP_422J2_124_3477_n2076), .CI(DP_OP_422J2_124_3477_n2083), .CO(
        DP_OP_422J2_124_3477_n1172), .S(DP_OP_422J2_124_3477_n1173) );
  FADDX1_HVT DP_OP_422J2_124_3477_U767 ( .A(DP_OP_422J2_124_3477_n2861), .B(
        DP_OP_422J2_124_3477_n2113), .CI(DP_OP_422J2_124_3477_n2120), .CO(
        DP_OP_422J2_124_3477_n1170), .S(DP_OP_422J2_124_3477_n1171) );
  FADDX1_HVT DP_OP_422J2_124_3477_U766 ( .A(DP_OP_422J2_124_3477_n2831), .B(
        DP_OP_422J2_124_3477_n2127), .CI(DP_OP_422J2_124_3477_n2157), .CO(
        DP_OP_422J2_124_3477_n1168), .S(DP_OP_422J2_124_3477_n1169) );
  FADDX1_HVT DP_OP_422J2_124_3477_U765 ( .A(DP_OP_422J2_124_3477_n2824), .B(
        DP_OP_422J2_124_3477_n2164), .CI(DP_OP_422J2_124_3477_n2171), .CO(
        DP_OP_422J2_124_3477_n1166), .S(DP_OP_422J2_124_3477_n1167) );
  FADDX1_HVT DP_OP_422J2_124_3477_U764 ( .A(DP_OP_422J2_124_3477_n2817), .B(
        DP_OP_422J2_124_3477_n2201), .CI(DP_OP_422J2_124_3477_n2208), .CO(
        DP_OP_422J2_124_3477_n1164), .S(DP_OP_422J2_124_3477_n1165) );
  FADDX1_HVT DP_OP_422J2_124_3477_U763 ( .A(DP_OP_422J2_124_3477_n2787), .B(
        DP_OP_422J2_124_3477_n2215), .CI(DP_OP_422J2_124_3477_n2245), .CO(
        DP_OP_422J2_124_3477_n1162), .S(DP_OP_422J2_124_3477_n1163) );
  FADDX1_HVT DP_OP_422J2_124_3477_U762 ( .A(DP_OP_422J2_124_3477_n2780), .B(
        DP_OP_422J2_124_3477_n2252), .CI(DP_OP_422J2_124_3477_n2259), .CO(
        DP_OP_422J2_124_3477_n1160), .S(DP_OP_422J2_124_3477_n1161) );
  FADDX1_HVT DP_OP_422J2_124_3477_U761 ( .A(DP_OP_422J2_124_3477_n2773), .B(
        DP_OP_422J2_124_3477_n2391), .CI(DP_OP_422J2_124_3477_n2435), .CO(
        DP_OP_422J2_124_3477_n1158), .S(DP_OP_422J2_124_3477_n1159) );
  FADDX1_HVT DP_OP_422J2_124_3477_U760 ( .A(DP_OP_422J2_124_3477_n2743), .B(
        DP_OP_422J2_124_3477_n2465), .CI(DP_OP_422J2_124_3477_n2472), .CO(
        DP_OP_422J2_124_3477_n1156), .S(DP_OP_422J2_124_3477_n1157) );
  FADDX1_HVT DP_OP_422J2_124_3477_U759 ( .A(DP_OP_422J2_124_3477_n2736), .B(
        DP_OP_422J2_124_3477_n2479), .CI(DP_OP_422J2_124_3477_n2509), .CO(
        DP_OP_422J2_124_3477_n1154), .S(DP_OP_422J2_124_3477_n1155) );
  FADDX1_HVT DP_OP_422J2_124_3477_U758 ( .A(DP_OP_422J2_124_3477_n2729), .B(
        DP_OP_422J2_124_3477_n2516), .CI(DP_OP_422J2_124_3477_n2523), .CO(
        DP_OP_422J2_124_3477_n1152), .S(DP_OP_422J2_124_3477_n1153) );
  FADDX1_HVT DP_OP_422J2_124_3477_U757 ( .A(DP_OP_422J2_124_3477_n2699), .B(
        DP_OP_422J2_124_3477_n2553), .CI(DP_OP_422J2_124_3477_n2560), .CO(
        DP_OP_422J2_124_3477_n1150), .S(DP_OP_422J2_124_3477_n1151) );
  FADDX1_HVT DP_OP_422J2_124_3477_U756 ( .A(DP_OP_422J2_124_3477_n2692), .B(
        DP_OP_422J2_124_3477_n2567), .CI(DP_OP_422J2_124_3477_n2597), .CO(
        DP_OP_422J2_124_3477_n1148), .S(DP_OP_422J2_124_3477_n1149) );
  FADDX1_HVT DP_OP_422J2_124_3477_U755 ( .A(DP_OP_422J2_124_3477_n2685), .B(
        DP_OP_422J2_124_3477_n2604), .CI(DP_OP_422J2_124_3477_n2611), .CO(
        DP_OP_422J2_124_3477_n1146), .S(DP_OP_422J2_124_3477_n1147) );
  FADDX1_HVT DP_OP_422J2_124_3477_U754 ( .A(DP_OP_422J2_124_3477_n2641), .B(
        DP_OP_422J2_124_3477_n2648), .CI(DP_OP_422J2_124_3477_n2655), .CO(
        DP_OP_422J2_124_3477_n1144), .S(DP_OP_422J2_124_3477_n1145) );
  FADDX1_HVT DP_OP_422J2_124_3477_U753 ( .A(DP_OP_422J2_124_3477_n1398), .B(
        DP_OP_422J2_124_3477_n1386), .CI(DP_OP_422J2_124_3477_n1384), .CO(
        DP_OP_422J2_124_3477_n1142), .S(DP_OP_422J2_124_3477_n1143) );
  FADDX1_HVT DP_OP_422J2_124_3477_U752 ( .A(DP_OP_422J2_124_3477_n1382), .B(
        DP_OP_422J2_124_3477_n1388), .CI(DP_OP_422J2_124_3477_n1211), .CO(
        DP_OP_422J2_124_3477_n1140), .S(DP_OP_422J2_124_3477_n1141) );
  FADDX1_HVT DP_OP_422J2_124_3477_U751 ( .A(DP_OP_422J2_124_3477_n1392), .B(
        DP_OP_422J2_124_3477_n1396), .CI(DP_OP_422J2_124_3477_n1390), .CO(
        DP_OP_422J2_124_3477_n1138), .S(DP_OP_422J2_124_3477_n1139) );
  FADDX1_HVT DP_OP_422J2_124_3477_U750 ( .A(DP_OP_422J2_124_3477_n1394), .B(
        DP_OP_422J2_124_3477_n1358), .CI(DP_OP_422J2_124_3477_n1356), .CO(
        DP_OP_422J2_124_3477_n1136), .S(DP_OP_422J2_124_3477_n1137) );
  FADDX1_HVT DP_OP_422J2_124_3477_U749 ( .A(DP_OP_422J2_124_3477_n1360), .B(
        DP_OP_422J2_124_3477_n1332), .CI(DP_OP_422J2_124_3477_n1380), .CO(
        DP_OP_422J2_124_3477_n1134), .S(DP_OP_422J2_124_3477_n1135) );
  FADDX1_HVT DP_OP_422J2_124_3477_U748 ( .A(DP_OP_422J2_124_3477_n1352), .B(
        DP_OP_422J2_124_3477_n1334), .CI(DP_OP_422J2_124_3477_n1378), .CO(
        DP_OP_422J2_124_3477_n1132), .S(DP_OP_422J2_124_3477_n1133) );
  FADDX1_HVT DP_OP_422J2_124_3477_U747 ( .A(DP_OP_422J2_124_3477_n1350), .B(
        DP_OP_422J2_124_3477_n1336), .CI(DP_OP_422J2_124_3477_n1376), .CO(
        DP_OP_422J2_124_3477_n1130), .S(DP_OP_422J2_124_3477_n1131) );
  FADDX1_HVT DP_OP_422J2_124_3477_U746 ( .A(DP_OP_422J2_124_3477_n1346), .B(
        DP_OP_422J2_124_3477_n1374), .CI(DP_OP_422J2_124_3477_n1372), .CO(
        DP_OP_422J2_124_3477_n1128), .S(DP_OP_422J2_124_3477_n1129) );
  FADDX1_HVT DP_OP_422J2_124_3477_U745 ( .A(DP_OP_422J2_124_3477_n1340), .B(
        DP_OP_422J2_124_3477_n1370), .CI(DP_OP_422J2_124_3477_n1368), .CO(
        DP_OP_422J2_124_3477_n1126), .S(DP_OP_422J2_124_3477_n1127) );
  FADDX1_HVT DP_OP_422J2_124_3477_U744 ( .A(DP_OP_422J2_124_3477_n1348), .B(
        DP_OP_422J2_124_3477_n1366), .CI(DP_OP_422J2_124_3477_n1364), .CO(
        DP_OP_422J2_124_3477_n1124), .S(DP_OP_422J2_124_3477_n1125) );
  FADDX1_HVT DP_OP_422J2_124_3477_U743 ( .A(DP_OP_422J2_124_3477_n1342), .B(
        DP_OP_422J2_124_3477_n1362), .CI(DP_OP_422J2_124_3477_n1354), .CO(
        DP_OP_422J2_124_3477_n1122), .S(DP_OP_422J2_124_3477_n1123) );
  FADDX1_HVT DP_OP_422J2_124_3477_U742 ( .A(DP_OP_422J2_124_3477_n1344), .B(
        DP_OP_422J2_124_3477_n1338), .CI(DP_OP_422J2_124_3477_n1201), .CO(
        DP_OP_422J2_124_3477_n1120), .S(DP_OP_422J2_124_3477_n1121) );
  FADDX1_HVT DP_OP_422J2_124_3477_U741 ( .A(DP_OP_422J2_124_3477_n1197), .B(
        DP_OP_422J2_124_3477_n1195), .CI(DP_OP_422J2_124_3477_n1199), .CO(
        DP_OP_422J2_124_3477_n1118), .S(DP_OP_422J2_124_3477_n1119) );
  FADDX1_HVT DP_OP_422J2_124_3477_U740 ( .A(DP_OP_422J2_124_3477_n1207), .B(
        DP_OP_422J2_124_3477_n1205), .CI(DP_OP_422J2_124_3477_n1209), .CO(
        DP_OP_422J2_124_3477_n1116), .S(DP_OP_422J2_124_3477_n1117) );
  FADDX1_HVT DP_OP_422J2_124_3477_U739 ( .A(DP_OP_422J2_124_3477_n1203), .B(
        DP_OP_422J2_124_3477_n1151), .CI(DP_OP_422J2_124_3477_n1153), .CO(
        DP_OP_422J2_124_3477_n1114), .S(DP_OP_422J2_124_3477_n1115) );
  FADDX1_HVT DP_OP_422J2_124_3477_U738 ( .A(DP_OP_422J2_124_3477_n1149), .B(
        DP_OP_422J2_124_3477_n1185), .CI(DP_OP_422J2_124_3477_n1181), .CO(
        DP_OP_422J2_124_3477_n1112), .S(DP_OP_422J2_124_3477_n1113) );
  FADDX1_HVT DP_OP_422J2_124_3477_U737 ( .A(DP_OP_422J2_124_3477_n1187), .B(
        DP_OP_422J2_124_3477_n1171), .CI(DP_OP_422J2_124_3477_n1177), .CO(
        DP_OP_422J2_124_3477_n1110), .S(DP_OP_422J2_124_3477_n1111) );
  FADDX1_HVT DP_OP_422J2_124_3477_U736 ( .A(DP_OP_422J2_124_3477_n1175), .B(
        DP_OP_422J2_124_3477_n1173), .CI(DP_OP_422J2_124_3477_n1157), .CO(
        DP_OP_422J2_124_3477_n1108), .S(DP_OP_422J2_124_3477_n1109) );
  FADDX1_HVT DP_OP_422J2_124_3477_U735 ( .A(DP_OP_422J2_124_3477_n1179), .B(
        DP_OP_422J2_124_3477_n1147), .CI(DP_OP_422J2_124_3477_n1145), .CO(
        DP_OP_422J2_124_3477_n1106), .S(DP_OP_422J2_124_3477_n1107) );
  FADDX1_HVT DP_OP_422J2_124_3477_U734 ( .A(DP_OP_422J2_124_3477_n1183), .B(
        DP_OP_422J2_124_3477_n1165), .CI(DP_OP_422J2_124_3477_n1167), .CO(
        DP_OP_422J2_124_3477_n1104), .S(DP_OP_422J2_124_3477_n1105) );
  FADDX1_HVT DP_OP_422J2_124_3477_U733 ( .A(DP_OP_422J2_124_3477_n1163), .B(
        DP_OP_422J2_124_3477_n1161), .CI(DP_OP_422J2_124_3477_n1155), .CO(
        DP_OP_422J2_124_3477_n1102), .S(DP_OP_422J2_124_3477_n1103) );
  FADDX1_HVT DP_OP_422J2_124_3477_U732 ( .A(DP_OP_422J2_124_3477_n1159), .B(
        DP_OP_422J2_124_3477_n1193), .CI(DP_OP_422J2_124_3477_n1191), .CO(
        DP_OP_422J2_124_3477_n1100), .S(DP_OP_422J2_124_3477_n1101) );
  FADDX1_HVT DP_OP_422J2_124_3477_U731 ( .A(DP_OP_422J2_124_3477_n1189), .B(
        DP_OP_422J2_124_3477_n1169), .CI(DP_OP_422J2_124_3477_n1330), .CO(
        DP_OP_422J2_124_3477_n1098), .S(DP_OP_422J2_124_3477_n1099) );
  FADDX1_HVT DP_OP_422J2_124_3477_U730 ( .A(DP_OP_422J2_124_3477_n1328), .B(
        DP_OP_422J2_124_3477_n1326), .CI(DP_OP_422J2_124_3477_n1324), .CO(
        DP_OP_422J2_124_3477_n1096), .S(DP_OP_422J2_124_3477_n1097) );
  FADDX1_HVT DP_OP_422J2_124_3477_U729 ( .A(DP_OP_422J2_124_3477_n1310), .B(
        DP_OP_422J2_124_3477_n1322), .CI(DP_OP_422J2_124_3477_n1308), .CO(
        DP_OP_422J2_124_3477_n1094), .S(DP_OP_422J2_124_3477_n1095) );
  FADDX1_HVT DP_OP_422J2_124_3477_U728 ( .A(DP_OP_422J2_124_3477_n1312), .B(
        DP_OP_422J2_124_3477_n1314), .CI(DP_OP_422J2_124_3477_n1320), .CO(
        DP_OP_422J2_124_3477_n1092), .S(DP_OP_422J2_124_3477_n1093) );
  FADDX1_HVT DP_OP_422J2_124_3477_U727 ( .A(DP_OP_422J2_124_3477_n1318), .B(
        DP_OP_422J2_124_3477_n1316), .CI(DP_OP_422J2_124_3477_n1143), .CO(
        DP_OP_422J2_124_3477_n1090), .S(DP_OP_422J2_124_3477_n1091) );
  FADDX1_HVT DP_OP_422J2_124_3477_U726 ( .A(DP_OP_422J2_124_3477_n1306), .B(
        DP_OP_422J2_124_3477_n1137), .CI(DP_OP_422J2_124_3477_n1304), .CO(
        DP_OP_422J2_124_3477_n1088), .S(DP_OP_422J2_124_3477_n1089) );
  FADDX1_HVT DP_OP_422J2_124_3477_U725 ( .A(DP_OP_422J2_124_3477_n1141), .B(
        DP_OP_422J2_124_3477_n1139), .CI(DP_OP_422J2_124_3477_n1302), .CO(
        DP_OP_422J2_124_3477_n1086), .S(DP_OP_422J2_124_3477_n1087) );
  FADDX1_HVT DP_OP_422J2_124_3477_U724 ( .A(DP_OP_422J2_124_3477_n1290), .B(
        DP_OP_422J2_124_3477_n1121), .CI(DP_OP_422J2_124_3477_n1135), .CO(
        DP_OP_422J2_124_3477_n1084), .S(DP_OP_422J2_124_3477_n1085) );
  FADDX1_HVT DP_OP_422J2_124_3477_U723 ( .A(DP_OP_422J2_124_3477_n1288), .B(
        DP_OP_422J2_124_3477_n1131), .CI(DP_OP_422J2_124_3477_n1133), .CO(
        DP_OP_422J2_124_3477_n1082), .S(DP_OP_422J2_124_3477_n1083) );
  FADDX1_HVT DP_OP_422J2_124_3477_U722 ( .A(DP_OP_422J2_124_3477_n1292), .B(
        DP_OP_422J2_124_3477_n1129), .CI(DP_OP_422J2_124_3477_n1127), .CO(
        DP_OP_422J2_124_3477_n1080), .S(DP_OP_422J2_124_3477_n1081) );
  FADDX1_HVT DP_OP_422J2_124_3477_U721 ( .A(DP_OP_422J2_124_3477_n1300), .B(
        DP_OP_422J2_124_3477_n1123), .CI(DP_OP_422J2_124_3477_n1125), .CO(
        DP_OP_422J2_124_3477_n1078), .S(DP_OP_422J2_124_3477_n1079) );
  FADDX1_HVT DP_OP_422J2_124_3477_U720 ( .A(DP_OP_422J2_124_3477_n1298), .B(
        DP_OP_422J2_124_3477_n1294), .CI(DP_OP_422J2_124_3477_n1296), .CO(
        DP_OP_422J2_124_3477_n1076), .S(DP_OP_422J2_124_3477_n1077) );
  FADDX1_HVT DP_OP_422J2_124_3477_U719 ( .A(DP_OP_422J2_124_3477_n1117), .B(
        DP_OP_422J2_124_3477_n1286), .CI(DP_OP_422J2_124_3477_n1115), .CO(
        DP_OP_422J2_124_3477_n1074), .S(DP_OP_422J2_124_3477_n1075) );
  FADDX1_HVT DP_OP_422J2_124_3477_U718 ( .A(DP_OP_422J2_124_3477_n1119), .B(
        DP_OP_422J2_124_3477_n1109), .CI(DP_OP_422J2_124_3477_n1111), .CO(
        DP_OP_422J2_124_3477_n1072), .S(DP_OP_422J2_124_3477_n1073) );
  FADDX1_HVT DP_OP_422J2_124_3477_U717 ( .A(DP_OP_422J2_124_3477_n1107), .B(
        DP_OP_422J2_124_3477_n1101), .CI(DP_OP_422J2_124_3477_n1284), .CO(
        DP_OP_422J2_124_3477_n1070), .S(DP_OP_422J2_124_3477_n1071) );
  FADDX1_HVT DP_OP_422J2_124_3477_U716 ( .A(DP_OP_422J2_124_3477_n1103), .B(
        DP_OP_422J2_124_3477_n1113), .CI(DP_OP_422J2_124_3477_n1105), .CO(
        DP_OP_422J2_124_3477_n1068), .S(DP_OP_422J2_124_3477_n1069) );
  FADDX1_HVT DP_OP_422J2_124_3477_U715 ( .A(DP_OP_422J2_124_3477_n1099), .B(
        DP_OP_422J2_124_3477_n1282), .CI(DP_OP_422J2_124_3477_n1278), .CO(
        DP_OP_422J2_124_3477_n1066), .S(DP_OP_422J2_124_3477_n1067) );
  FADDX1_HVT DP_OP_422J2_124_3477_U714 ( .A(DP_OP_422J2_124_3477_n1280), .B(
        DP_OP_422J2_124_3477_n1276), .CI(DP_OP_422J2_124_3477_n1274), .CO(
        DP_OP_422J2_124_3477_n1064), .S(DP_OP_422J2_124_3477_n1065) );
  FADDX1_HVT DP_OP_422J2_124_3477_U713 ( .A(DP_OP_422J2_124_3477_n1097), .B(
        DP_OP_422J2_124_3477_n1272), .CI(DP_OP_422J2_124_3477_n1270), .CO(
        DP_OP_422J2_124_3477_n1062), .S(DP_OP_422J2_124_3477_n1063) );
  FADDX1_HVT DP_OP_422J2_124_3477_U712 ( .A(DP_OP_422J2_124_3477_n1268), .B(
        DP_OP_422J2_124_3477_n1093), .CI(DP_OP_422J2_124_3477_n1091), .CO(
        DP_OP_422J2_124_3477_n1060), .S(DP_OP_422J2_124_3477_n1061) );
  FADDX1_HVT DP_OP_422J2_124_3477_U711 ( .A(DP_OP_422J2_124_3477_n1266), .B(
        DP_OP_422J2_124_3477_n1264), .CI(DP_OP_422J2_124_3477_n1095), .CO(
        DP_OP_422J2_124_3477_n1058), .S(DP_OP_422J2_124_3477_n1059) );
  FADDX1_HVT DP_OP_422J2_124_3477_U710 ( .A(DP_OP_422J2_124_3477_n1087), .B(
        DP_OP_422J2_124_3477_n1262), .CI(DP_OP_422J2_124_3477_n1089), .CO(
        DP_OP_422J2_124_3477_n1056), .S(DP_OP_422J2_124_3477_n1057) );
  FADDX1_HVT DP_OP_422J2_124_3477_U709 ( .A(DP_OP_422J2_124_3477_n1081), .B(
        DP_OP_422J2_124_3477_n1085), .CI(DP_OP_422J2_124_3477_n1256), .CO(
        DP_OP_422J2_124_3477_n1054), .S(DP_OP_422J2_124_3477_n1055) );
  FADDX1_HVT DP_OP_422J2_124_3477_U708 ( .A(DP_OP_422J2_124_3477_n1260), .B(
        DP_OP_422J2_124_3477_n1079), .CI(DP_OP_422J2_124_3477_n1083), .CO(
        DP_OP_422J2_124_3477_n1052), .S(DP_OP_422J2_124_3477_n1053) );
  FADDX1_HVT DP_OP_422J2_124_3477_U706 ( .A(DP_OP_422J2_124_3477_n1075), .B(
        DP_OP_422J2_124_3477_n1073), .CI(DP_OP_422J2_124_3477_n1071), .CO(
        DP_OP_422J2_124_3477_n1048), .S(DP_OP_422J2_124_3477_n1049) );
  FADDX1_HVT DP_OP_422J2_124_3477_U705 ( .A(DP_OP_422J2_124_3477_n1069), .B(
        DP_OP_422J2_124_3477_n1252), .CI(DP_OP_422J2_124_3477_n1067), .CO(
        DP_OP_422J2_124_3477_n1046), .S(DP_OP_422J2_124_3477_n1047) );
  FADDX1_HVT DP_OP_422J2_124_3477_U703 ( .A(DP_OP_422J2_124_3477_n1065), .B(
        DP_OP_422J2_124_3477_n1244), .CI(DP_OP_422J2_124_3477_n1063), .CO(
        DP_OP_422J2_124_3477_n1042), .S(DP_OP_422J2_124_3477_n1043) );
  FADDX1_HVT DP_OP_422J2_124_3477_U702 ( .A(DP_OP_422J2_124_3477_n1059), .B(
        DP_OP_422J2_124_3477_n1242), .CI(DP_OP_422J2_124_3477_n1061), .CO(
        DP_OP_422J2_124_3477_n1040), .S(DP_OP_422J2_124_3477_n1041) );
  FADDX1_HVT DP_OP_422J2_124_3477_U701 ( .A(DP_OP_422J2_124_3477_n1240), .B(
        DP_OP_422J2_124_3477_n1238), .CI(DP_OP_422J2_124_3477_n1057), .CO(
        DP_OP_422J2_124_3477_n1038), .S(DP_OP_422J2_124_3477_n1039) );
  FADDX1_HVT DP_OP_422J2_124_3477_U700 ( .A(DP_OP_422J2_124_3477_n1236), .B(
        DP_OP_422J2_124_3477_n1053), .CI(DP_OP_422J2_124_3477_n1051), .CO(
        DP_OP_422J2_124_3477_n1036), .S(DP_OP_422J2_124_3477_n1037) );
  FADDX1_HVT DP_OP_422J2_124_3477_U699 ( .A(DP_OP_422J2_124_3477_n1055), .B(
        DP_OP_422J2_124_3477_n1234), .CI(DP_OP_422J2_124_3477_n1049), .CO(
        DP_OP_422J2_124_3477_n1034), .S(DP_OP_422J2_124_3477_n1035) );
  FADDX1_HVT DP_OP_422J2_124_3477_U698 ( .A(DP_OP_422J2_124_3477_n1232), .B(
        DP_OP_422J2_124_3477_n1047), .CI(DP_OP_422J2_124_3477_n1230), .CO(
        DP_OP_422J2_124_3477_n1032), .S(DP_OP_422J2_124_3477_n1033) );
  FADDX1_HVT DP_OP_422J2_124_3477_U697 ( .A(DP_OP_422J2_124_3477_n1045), .B(
        DP_OP_422J2_124_3477_n1228), .CI(DP_OP_422J2_124_3477_n1043), .CO(
        DP_OP_422J2_124_3477_n1030), .S(DP_OP_422J2_124_3477_n1031) );
  FADDX1_HVT DP_OP_422J2_124_3477_U696 ( .A(DP_OP_422J2_124_3477_n1226), .B(
        DP_OP_422J2_124_3477_n1041), .CI(DP_OP_422J2_124_3477_n1039), .CO(
        DP_OP_422J2_124_3477_n1028), .S(DP_OP_422J2_124_3477_n1029) );
  FADDX1_HVT DP_OP_422J2_124_3477_U695 ( .A(DP_OP_422J2_124_3477_n1224), .B(
        DP_OP_422J2_124_3477_n1037), .CI(DP_OP_422J2_124_3477_n1222), .CO(
        DP_OP_422J2_124_3477_n1026), .S(DP_OP_422J2_124_3477_n1027) );
  FADDX1_HVT DP_OP_422J2_124_3477_U694 ( .A(DP_OP_422J2_124_3477_n1035), .B(
        DP_OP_422J2_124_3477_n1220), .CI(DP_OP_422J2_124_3477_n1033), .CO(
        DP_OP_422J2_124_3477_n1024), .S(DP_OP_422J2_124_3477_n1025) );
  FADDX1_HVT DP_OP_422J2_124_3477_U693 ( .A(DP_OP_422J2_124_3477_n1031), .B(
        DP_OP_422J2_124_3477_n1218), .CI(DP_OP_422J2_124_3477_n1029), .CO(
        DP_OP_422J2_124_3477_n1022), .S(DP_OP_422J2_124_3477_n1023) );
  FADDX1_HVT DP_OP_422J2_124_3477_U692 ( .A(DP_OP_422J2_124_3477_n1216), .B(
        DP_OP_422J2_124_3477_n1027), .CI(DP_OP_422J2_124_3477_n1025), .CO(
        DP_OP_422J2_124_3477_n1020), .S(DP_OP_422J2_124_3477_n1021) );
  FADDX1_HVT DP_OP_422J2_124_3477_U691 ( .A(DP_OP_422J2_124_3477_n1214), .B(
        DP_OP_422J2_124_3477_n1023), .CI(DP_OP_422J2_124_3477_n1212), .CO(
        DP_OP_422J2_124_3477_n1018), .S(DP_OP_422J2_124_3477_n1019) );
  FADDX1_HVT DP_OP_422J2_124_3477_U690 ( .A(DP_OP_422J2_124_3477_n3028), .B(
        DP_OP_422J2_124_3477_n1973), .CI(DP_OP_422J2_124_3477_n1929), .CO(
        DP_OP_422J2_124_3477_n1016), .S(DP_OP_422J2_124_3477_n1017) );
  FADDX1_HVT DP_OP_422J2_124_3477_U689 ( .A(DP_OP_422J2_124_3477_n2853), .B(
        DP_OP_422J2_124_3477_n2170), .CI(DP_OP_422J2_124_3477_n2434), .CO(
        DP_OP_422J2_124_3477_n1014), .S(DP_OP_422J2_124_3477_n1015) );
  FADDX1_HVT DP_OP_422J2_124_3477_U688 ( .A(DP_OP_422J2_124_3477_n2061), .B(
        DP_OP_422J2_124_3477_n2478), .CI(DP_OP_422J2_124_3477_n2038), .CO(
        DP_OP_422J2_124_3477_n1012), .S(DP_OP_422J2_124_3477_n1013) );
  FADDX1_HVT DP_OP_422J2_124_3477_U687 ( .A(DP_OP_422J2_124_3477_n2369), .B(
        DP_OP_422J2_124_3477_n1994), .CI(DP_OP_422J2_124_3477_n2962), .CO(
        DP_OP_422J2_124_3477_n1010), .S(DP_OP_422J2_124_3477_n1011) );
  FADDX1_HVT DP_OP_422J2_124_3477_U686 ( .A(DP_OP_422J2_124_3477_n2325), .B(
        DP_OP_422J2_124_3477_n2302), .CI(DP_OP_422J2_124_3477_n2654), .CO(
        DP_OP_422J2_124_3477_n1008), .S(DP_OP_422J2_124_3477_n1009) );
  FADDX1_HVT DP_OP_422J2_124_3477_U685 ( .A(DP_OP_422J2_124_3477_n2237), .B(
        DP_OP_422J2_124_3477_n2346), .CI(DP_OP_422J2_124_3477_n3006), .CO(
        DP_OP_422J2_124_3477_n1006), .S(DP_OP_422J2_124_3477_n1007) );
  FADDX1_HVT DP_OP_422J2_124_3477_U684 ( .A(DP_OP_422J2_124_3477_n2017), .B(
        DP_OP_422J2_124_3477_n2082), .CI(DP_OP_422J2_124_3477_n2522), .CO(
        DP_OP_422J2_124_3477_n1004), .S(DP_OP_422J2_124_3477_n1005) );
  FADDX1_HVT DP_OP_422J2_124_3477_U683 ( .A(DP_OP_422J2_124_3477_n2105), .B(
        DP_OP_422J2_124_3477_n2786), .CI(DP_OP_422J2_124_3477_n2830), .CO(
        DP_OP_422J2_124_3477_n1002), .S(DP_OP_422J2_124_3477_n1003) );
  FADDX1_HVT DP_OP_422J2_124_3477_U682 ( .A(DP_OP_422J2_124_3477_n2193), .B(
        DP_OP_422J2_124_3477_n2742), .CI(DP_OP_422J2_124_3477_n2610), .CO(
        DP_OP_422J2_124_3477_n1000), .S(DP_OP_422J2_124_3477_n1001) );
  FADDX1_HVT DP_OP_422J2_124_3477_U681 ( .A(DP_OP_422J2_124_3477_n2545), .B(
        DP_OP_422J2_124_3477_n2390), .CI(DP_OP_422J2_124_3477_n2874), .CO(
        DP_OP_422J2_124_3477_n998), .S(DP_OP_422J2_124_3477_n999) );
  FADDX1_HVT DP_OP_422J2_124_3477_U680 ( .A(DP_OP_422J2_124_3477_n2941), .B(
        DP_OP_422J2_124_3477_n2214), .CI(DP_OP_422J2_124_3477_n2126), .CO(
        DP_OP_422J2_124_3477_n996), .S(DP_OP_422J2_124_3477_n997) );
  FADDX1_HVT DP_OP_422J2_124_3477_U679 ( .A(DP_OP_422J2_124_3477_n2677), .B(
        DP_OP_422J2_124_3477_n2918), .CI(DP_OP_422J2_124_3477_n2566), .CO(
        DP_OP_422J2_124_3477_n994), .S(DP_OP_422J2_124_3477_n995) );
  FADDX1_HVT DP_OP_422J2_124_3477_U678 ( .A(DP_OP_422J2_124_3477_n2457), .B(
        DP_OP_422J2_124_3477_n3048), .CI(DP_OP_422J2_124_3477_n2258), .CO(
        DP_OP_422J2_124_3477_n992), .S(DP_OP_422J2_124_3477_n993) );
  FADDX1_HVT DP_OP_422J2_124_3477_U677 ( .A(DP_OP_422J2_124_3477_n2149), .B(
        DP_OP_422J2_124_3477_n2413), .CI(DP_OP_422J2_124_3477_n2698), .CO(
        DP_OP_422J2_124_3477_n990), .S(DP_OP_422J2_124_3477_n991) );
  FADDX1_HVT DP_OP_422J2_124_3477_U676 ( .A(DP_OP_422J2_124_3477_n2765), .B(
        DP_OP_422J2_124_3477_n2809), .CI(DP_OP_422J2_124_3477_n2897), .CO(
        DP_OP_422J2_124_3477_n988), .S(DP_OP_422J2_124_3477_n989) );
  FADDX1_HVT DP_OP_422J2_124_3477_U675 ( .A(DP_OP_422J2_124_3477_n2501), .B(
        DP_OP_422J2_124_3477_n2589), .CI(DP_OP_422J2_124_3477_n2985), .CO(
        DP_OP_422J2_124_3477_n986), .S(DP_OP_422J2_124_3477_n987) );
  FADDX1_HVT DP_OP_422J2_124_3477_U674 ( .A(DP_OP_422J2_124_3477_n2633), .B(
        DP_OP_422J2_124_3477_n2281), .CI(DP_OP_422J2_124_3477_n2721), .CO(
        DP_OP_422J2_124_3477_n984), .S(DP_OP_422J2_124_3477_n985) );
  FADDX1_HVT DP_OP_422J2_124_3477_U673 ( .A(DP_OP_422J2_124_3477_n3041), .B(
        DP_OP_422J2_124_3477_n1987), .CI(DP_OP_422J2_124_3477_n1980), .CO(
        DP_OP_422J2_124_3477_n982), .S(DP_OP_422J2_124_3477_n983) );
  FADDX1_HVT DP_OP_422J2_124_3477_U672 ( .A(DP_OP_422J2_124_3477_n3034), .B(
        DP_OP_422J2_124_3477_n2999), .CI(DP_OP_422J2_124_3477_n2992), .CO(
        DP_OP_422J2_124_3477_n980), .S(DP_OP_422J2_124_3477_n981) );
  FADDX1_HVT DP_OP_422J2_124_3477_U671 ( .A(DP_OP_422J2_124_3477_n2515), .B(
        DP_OP_422J2_124_3477_n2955), .CI(DP_OP_422J2_124_3477_n2948), .CO(
        DP_OP_422J2_124_3477_n978), .S(DP_OP_422J2_124_3477_n979) );
  FADDX1_HVT DP_OP_422J2_124_3477_U670 ( .A(DP_OP_422J2_124_3477_n2911), .B(
        DP_OP_422J2_124_3477_n2024), .CI(DP_OP_422J2_124_3477_n2031), .CO(
        DP_OP_422J2_124_3477_n976), .S(DP_OP_422J2_124_3477_n977) );
  FADDX1_HVT DP_OP_422J2_124_3477_U669 ( .A(DP_OP_422J2_124_3477_n2904), .B(
        DP_OP_422J2_124_3477_n2068), .CI(DP_OP_422J2_124_3477_n2075), .CO(
        DP_OP_422J2_124_3477_n974), .S(DP_OP_422J2_124_3477_n975) );
  FADDX1_HVT DP_OP_422J2_124_3477_U668 ( .A(DP_OP_422J2_124_3477_n2867), .B(
        DP_OP_422J2_124_3477_n2112), .CI(DP_OP_422J2_124_3477_n2119), .CO(
        DP_OP_422J2_124_3477_n972), .S(DP_OP_422J2_124_3477_n973) );
  FADDX1_HVT DP_OP_422J2_124_3477_U666 ( .A(DP_OP_422J2_124_3477_n2823), .B(
        DP_OP_422J2_124_3477_n2200), .CI(DP_OP_422J2_124_3477_n2207), .CO(
        DP_OP_422J2_124_3477_n968), .S(DP_OP_422J2_124_3477_n969) );
  FADDX1_HVT DP_OP_422J2_124_3477_U665 ( .A(DP_OP_422J2_124_3477_n2816), .B(
        DP_OP_422J2_124_3477_n2244), .CI(DP_OP_422J2_124_3477_n2251), .CO(
        DP_OP_422J2_124_3477_n966), .S(DP_OP_422J2_124_3477_n967) );
  FADDX1_HVT DP_OP_422J2_124_3477_U664 ( .A(DP_OP_422J2_124_3477_n2779), .B(
        DP_OP_422J2_124_3477_n2288), .CI(DP_OP_422J2_124_3477_n2295), .CO(
        DP_OP_422J2_124_3477_n964), .S(DP_OP_422J2_124_3477_n965) );
  FADDX1_HVT DP_OP_422J2_124_3477_U663 ( .A(DP_OP_422J2_124_3477_n2772), .B(
        DP_OP_422J2_124_3477_n2339), .CI(DP_OP_422J2_124_3477_n2332), .CO(
        DP_OP_422J2_124_3477_n962), .S(DP_OP_422J2_124_3477_n963) );
  FADDX1_HVT DP_OP_422J2_124_3477_U662 ( .A(DP_OP_422J2_124_3477_n2735), .B(
        DP_OP_422J2_124_3477_n2376), .CI(DP_OP_422J2_124_3477_n2383), .CO(
        DP_OP_422J2_124_3477_n960), .S(DP_OP_422J2_124_3477_n961) );
  FADDX1_HVT DP_OP_422J2_124_3477_U661 ( .A(DP_OP_422J2_124_3477_n2728), .B(
        DP_OP_422J2_124_3477_n2420), .CI(DP_OP_422J2_124_3477_n2427), .CO(
        DP_OP_422J2_124_3477_n958), .S(DP_OP_422J2_124_3477_n959) );
  FADDX1_HVT DP_OP_422J2_124_3477_U660 ( .A(DP_OP_422J2_124_3477_n2691), .B(
        DP_OP_422J2_124_3477_n2464), .CI(DP_OP_422J2_124_3477_n2471), .CO(
        DP_OP_422J2_124_3477_n956), .S(DP_OP_422J2_124_3477_n957) );
  FADDX1_HVT DP_OP_422J2_124_3477_U659 ( .A(DP_OP_422J2_124_3477_n2684), .B(
        DP_OP_422J2_124_3477_n2508), .CI(DP_OP_422J2_124_3477_n2552), .CO(
        DP_OP_422J2_124_3477_n954), .S(DP_OP_422J2_124_3477_n955) );
  FADDX1_HVT DP_OP_422J2_124_3477_U658 ( .A(DP_OP_422J2_124_3477_n2647), .B(
        DP_OP_422J2_124_3477_n2559), .CI(DP_OP_422J2_124_3477_n2596), .CO(
        DP_OP_422J2_124_3477_n952), .S(DP_OP_422J2_124_3477_n953) );
  FADDX1_HVT DP_OP_422J2_124_3477_U657 ( .A(DP_OP_422J2_124_3477_n2640), .B(
        DP_OP_422J2_124_3477_n2603), .CI(DP_OP_422J2_124_3477_n1210), .CO(
        DP_OP_422J2_124_3477_n950), .S(DP_OP_422J2_124_3477_n951) );
  FADDX1_HVT DP_OP_422J2_124_3477_U656 ( .A(DP_OP_422J2_124_3477_n1198), .B(
        DP_OP_422J2_124_3477_n1194), .CI(DP_OP_422J2_124_3477_n1208), .CO(
        DP_OP_422J2_124_3477_n948), .S(DP_OP_422J2_124_3477_n949) );
  FADDX1_HVT DP_OP_422J2_124_3477_U655 ( .A(DP_OP_422J2_124_3477_n1206), .B(
        DP_OP_422J2_124_3477_n1196), .CI(DP_OP_422J2_124_3477_n1204), .CO(
        DP_OP_422J2_124_3477_n946), .S(DP_OP_422J2_124_3477_n947) );
  FADDX1_HVT DP_OP_422J2_124_3477_U654 ( .A(DP_OP_422J2_124_3477_n1202), .B(
        DP_OP_422J2_124_3477_n1200), .CI(DP_OP_422J2_124_3477_n1170), .CO(
        DP_OP_422J2_124_3477_n944), .S(DP_OP_422J2_124_3477_n945) );
  FADDX1_HVT DP_OP_422J2_124_3477_U653 ( .A(DP_OP_422J2_124_3477_n1168), .B(
        DP_OP_422J2_124_3477_n1144), .CI(DP_OP_422J2_124_3477_n1192), .CO(
        DP_OP_422J2_124_3477_n942), .S(DP_OP_422J2_124_3477_n943) );
  FADDX1_HVT DP_OP_422J2_124_3477_U652 ( .A(DP_OP_422J2_124_3477_n1166), .B(
        DP_OP_422J2_124_3477_n1190), .CI(DP_OP_422J2_124_3477_n1188), .CO(
        DP_OP_422J2_124_3477_n940), .S(DP_OP_422J2_124_3477_n941) );
  FADDX1_HVT DP_OP_422J2_124_3477_U651 ( .A(DP_OP_422J2_124_3477_n1160), .B(
        DP_OP_422J2_124_3477_n1186), .CI(DP_OP_422J2_124_3477_n1184), .CO(
        DP_OP_422J2_124_3477_n938), .S(DP_OP_422J2_124_3477_n939) );
  FADDX1_HVT DP_OP_422J2_124_3477_U650 ( .A(DP_OP_422J2_124_3477_n1182), .B(
        DP_OP_422J2_124_3477_n1180), .CI(DP_OP_422J2_124_3477_n1178), .CO(
        DP_OP_422J2_124_3477_n936), .S(DP_OP_422J2_124_3477_n937) );
  FADDX1_HVT DP_OP_422J2_124_3477_U649 ( .A(DP_OP_422J2_124_3477_n1150), .B(
        DP_OP_422J2_124_3477_n1176), .CI(DP_OP_422J2_124_3477_n1174), .CO(
        DP_OP_422J2_124_3477_n934), .S(DP_OP_422J2_124_3477_n935) );
  FADDX1_HVT DP_OP_422J2_124_3477_U648 ( .A(DP_OP_422J2_124_3477_n1156), .B(
        DP_OP_422J2_124_3477_n1172), .CI(DP_OP_422J2_124_3477_n1164), .CO(
        DP_OP_422J2_124_3477_n932), .S(DP_OP_422J2_124_3477_n933) );
  FADDX1_HVT DP_OP_422J2_124_3477_U647 ( .A(DP_OP_422J2_124_3477_n1148), .B(
        DP_OP_422J2_124_3477_n1162), .CI(DP_OP_422J2_124_3477_n1158), .CO(
        DP_OP_422J2_124_3477_n930), .S(DP_OP_422J2_124_3477_n931) );
  FADDX1_HVT DP_OP_422J2_124_3477_U646 ( .A(DP_OP_422J2_124_3477_n1152), .B(
        DP_OP_422J2_124_3477_n1146), .CI(DP_OP_422J2_124_3477_n1154), .CO(
        DP_OP_422J2_124_3477_n928), .S(DP_OP_422J2_124_3477_n929) );
  FADDX1_HVT DP_OP_422J2_124_3477_U645 ( .A(DP_OP_422J2_124_3477_n1017), .B(
        DP_OP_422J2_124_3477_n1003), .CI(DP_OP_422J2_124_3477_n1005), .CO(
        DP_OP_422J2_124_3477_n926), .S(DP_OP_422J2_124_3477_n927) );
  FADDX1_HVT DP_OP_422J2_124_3477_U644 ( .A(DP_OP_422J2_124_3477_n1009), .B(
        DP_OP_422J2_124_3477_n987), .CI(DP_OP_422J2_124_3477_n985), .CO(
        DP_OP_422J2_124_3477_n924), .S(DP_OP_422J2_124_3477_n925) );
  FADDX1_HVT DP_OP_422J2_124_3477_U643 ( .A(DP_OP_422J2_124_3477_n1001), .B(
        DP_OP_422J2_124_3477_n999), .CI(DP_OP_422J2_124_3477_n995), .CO(
        DP_OP_422J2_124_3477_n922), .S(DP_OP_422J2_124_3477_n923) );
  FADDX1_HVT DP_OP_422J2_124_3477_U642 ( .A(DP_OP_422J2_124_3477_n1007), .B(
        DP_OP_422J2_124_3477_n989), .CI(DP_OP_422J2_124_3477_n993), .CO(
        DP_OP_422J2_124_3477_n920), .S(DP_OP_422J2_124_3477_n921) );
  FADDX1_HVT DP_OP_422J2_124_3477_U641 ( .A(DP_OP_422J2_124_3477_n997), .B(
        DP_OP_422J2_124_3477_n1015), .CI(DP_OP_422J2_124_3477_n1011), .CO(
        DP_OP_422J2_124_3477_n918), .S(DP_OP_422J2_124_3477_n919) );
  FADDX1_HVT DP_OP_422J2_124_3477_U640 ( .A(DP_OP_422J2_124_3477_n991), .B(
        DP_OP_422J2_124_3477_n1013), .CI(DP_OP_422J2_124_3477_n973), .CO(
        DP_OP_422J2_124_3477_n916), .S(DP_OP_422J2_124_3477_n917) );
  FADDX1_HVT DP_OP_422J2_124_3477_U639 ( .A(DP_OP_422J2_124_3477_n975), .B(
        DP_OP_422J2_124_3477_n957), .CI(DP_OP_422J2_124_3477_n951), .CO(
        DP_OP_422J2_124_3477_n914), .S(DP_OP_422J2_124_3477_n915) );
  FADDX1_HVT DP_OP_422J2_124_3477_U638 ( .A(DP_OP_422J2_124_3477_n977), .B(
        DP_OP_422J2_124_3477_n953), .CI(DP_OP_422J2_124_3477_n969), .CO(
        DP_OP_422J2_124_3477_n912), .S(DP_OP_422J2_124_3477_n913) );
  FADDX1_HVT DP_OP_422J2_124_3477_U637 ( .A(DP_OP_422J2_124_3477_n967), .B(
        DP_OP_422J2_124_3477_n965), .CI(DP_OP_422J2_124_3477_n955), .CO(
        DP_OP_422J2_124_3477_n910), .S(DP_OP_422J2_124_3477_n911) );
  FADDX1_HVT DP_OP_422J2_124_3477_U636 ( .A(DP_OP_422J2_124_3477_n961), .B(
        DP_OP_422J2_124_3477_n959), .CI(DP_OP_422J2_124_3477_n971), .CO(
        DP_OP_422J2_124_3477_n908), .S(DP_OP_422J2_124_3477_n909) );
  FADDX1_HVT DP_OP_422J2_124_3477_U635 ( .A(DP_OP_422J2_124_3477_n979), .B(
        DP_OP_422J2_124_3477_n983), .CI(DP_OP_422J2_124_3477_n981), .CO(
        DP_OP_422J2_124_3477_n906), .S(DP_OP_422J2_124_3477_n907) );
  FADDX1_HVT DP_OP_422J2_124_3477_U634 ( .A(DP_OP_422J2_124_3477_n963), .B(
        DP_OP_422J2_124_3477_n1142), .CI(DP_OP_422J2_124_3477_n1140), .CO(
        DP_OP_422J2_124_3477_n904), .S(DP_OP_422J2_124_3477_n905) );
  FADDX1_HVT DP_OP_422J2_124_3477_U633 ( .A(DP_OP_422J2_124_3477_n1138), .B(
        DP_OP_422J2_124_3477_n1136), .CI(DP_OP_422J2_124_3477_n1122), .CO(
        DP_OP_422J2_124_3477_n902), .S(DP_OP_422J2_124_3477_n903) );
  FADDX1_HVT DP_OP_422J2_124_3477_U631 ( .A(DP_OP_422J2_124_3477_n1130), .B(
        DP_OP_422J2_124_3477_n1124), .CI(DP_OP_422J2_124_3477_n1126), .CO(
        DP_OP_422J2_124_3477_n898), .S(DP_OP_422J2_124_3477_n899) );
  FADDX1_HVT DP_OP_422J2_124_3477_U630 ( .A(DP_OP_422J2_124_3477_n1128), .B(
        DP_OP_422J2_124_3477_n1118), .CI(DP_OP_422J2_124_3477_n1116), .CO(
        DP_OP_422J2_124_3477_n896), .S(DP_OP_422J2_124_3477_n897) );
  FADDX1_HVT DP_OP_422J2_124_3477_U629 ( .A(DP_OP_422J2_124_3477_n949), .B(
        DP_OP_422J2_124_3477_n945), .CI(DP_OP_422J2_124_3477_n1114), .CO(
        DP_OP_422J2_124_3477_n894), .S(DP_OP_422J2_124_3477_n895) );
  FADDX1_HVT DP_OP_422J2_124_3477_U628 ( .A(DP_OP_422J2_124_3477_n947), .B(
        DP_OP_422J2_124_3477_n1102), .CI(DP_OP_422J2_124_3477_n1100), .CO(
        DP_OP_422J2_124_3477_n892), .S(DP_OP_422J2_124_3477_n893) );
  FADDX1_HVT DP_OP_422J2_124_3477_U626 ( .A(DP_OP_422J2_124_3477_n929), .B(
        DP_OP_422J2_124_3477_n939), .CI(DP_OP_422J2_124_3477_n1106), .CO(
        DP_OP_422J2_124_3477_n888), .S(DP_OP_422J2_124_3477_n889) );
  FADDX1_HVT DP_OP_422J2_124_3477_U625 ( .A(DP_OP_422J2_124_3477_n1112), .B(
        DP_OP_422J2_124_3477_n935), .CI(DP_OP_422J2_124_3477_n937), .CO(
        DP_OP_422J2_124_3477_n886), .S(DP_OP_422J2_124_3477_n887) );
  FADDX1_HVT DP_OP_422J2_124_3477_U624 ( .A(DP_OP_422J2_124_3477_n1110), .B(
        DP_OP_422J2_124_3477_n931), .CI(DP_OP_422J2_124_3477_n933), .CO(
        DP_OP_422J2_124_3477_n884), .S(DP_OP_422J2_124_3477_n885) );
  FADDX1_HVT DP_OP_422J2_124_3477_U623 ( .A(DP_OP_422J2_124_3477_n1104), .B(
        DP_OP_422J2_124_3477_n941), .CI(DP_OP_422J2_124_3477_n927), .CO(
        DP_OP_422J2_124_3477_n882), .S(DP_OP_422J2_124_3477_n883) );
  FADDX1_HVT DP_OP_422J2_124_3477_U622 ( .A(DP_OP_422J2_124_3477_n921), .B(
        DP_OP_422J2_124_3477_n925), .CI(DP_OP_422J2_124_3477_n917), .CO(
        DP_OP_422J2_124_3477_n880), .S(DP_OP_422J2_124_3477_n881) );
  FADDX1_HVT DP_OP_422J2_124_3477_U621 ( .A(DP_OP_422J2_124_3477_n919), .B(
        DP_OP_422J2_124_3477_n923), .CI(DP_OP_422J2_124_3477_n911), .CO(
        DP_OP_422J2_124_3477_n878), .S(DP_OP_422J2_124_3477_n879) );
  FADDX1_HVT DP_OP_422J2_124_3477_U620 ( .A(DP_OP_422J2_124_3477_n909), .B(
        DP_OP_422J2_124_3477_n915), .CI(DP_OP_422J2_124_3477_n1096), .CO(
        DP_OP_422J2_124_3477_n876), .S(DP_OP_422J2_124_3477_n877) );
  FADDX1_HVT DP_OP_422J2_124_3477_U619 ( .A(DP_OP_422J2_124_3477_n907), .B(
        DP_OP_422J2_124_3477_n913), .CI(DP_OP_422J2_124_3477_n1092), .CO(
        DP_OP_422J2_124_3477_n874), .S(DP_OP_422J2_124_3477_n875) );
  FADDX1_HVT DP_OP_422J2_124_3477_U618 ( .A(DP_OP_422J2_124_3477_n905), .B(
        DP_OP_422J2_124_3477_n1090), .CI(DP_OP_422J2_124_3477_n1094), .CO(
        DP_OP_422J2_124_3477_n872), .S(DP_OP_422J2_124_3477_n873) );
  FADDX1_HVT DP_OP_422J2_124_3477_U617 ( .A(DP_OP_422J2_124_3477_n1088), .B(
        DP_OP_422J2_124_3477_n1086), .CI(DP_OP_422J2_124_3477_n903), .CO(
        DP_OP_422J2_124_3477_n870), .S(DP_OP_422J2_124_3477_n871) );
  FADDX1_HVT DP_OP_422J2_124_3477_U616 ( .A(DP_OP_422J2_124_3477_n1084), .B(
        DP_OP_422J2_124_3477_n901), .CI(DP_OP_422J2_124_3477_n899), .CO(
        DP_OP_422J2_124_3477_n868), .S(DP_OP_422J2_124_3477_n869) );
  FADDX1_HVT DP_OP_422J2_124_3477_U615 ( .A(DP_OP_422J2_124_3477_n1082), .B(
        DP_OP_422J2_124_3477_n1076), .CI(DP_OP_422J2_124_3477_n1078), .CO(
        DP_OP_422J2_124_3477_n866), .S(DP_OP_422J2_124_3477_n867) );
  FADDX1_HVT DP_OP_422J2_124_3477_U614 ( .A(DP_OP_422J2_124_3477_n1080), .B(
        DP_OP_422J2_124_3477_n897), .CI(DP_OP_422J2_124_3477_n1074), .CO(
        DP_OP_422J2_124_3477_n864), .S(DP_OP_422J2_124_3477_n865) );
  FADDX1_HVT DP_OP_422J2_124_3477_U613 ( .A(DP_OP_422J2_124_3477_n895), .B(
        DP_OP_422J2_124_3477_n1072), .CI(DP_OP_422J2_124_3477_n893), .CO(
        DP_OP_422J2_124_3477_n862), .S(DP_OP_422J2_124_3477_n863) );
  FADDX1_HVT DP_OP_422J2_124_3477_U612 ( .A(DP_OP_422J2_124_3477_n1070), .B(
        DP_OP_422J2_124_3477_n887), .CI(DP_OP_422J2_124_3477_n883), .CO(
        DP_OP_422J2_124_3477_n860), .S(DP_OP_422J2_124_3477_n861) );
  FADDX1_HVT DP_OP_422J2_124_3477_U611 ( .A(DP_OP_422J2_124_3477_n1068), .B(
        DP_OP_422J2_124_3477_n891), .CI(DP_OP_422J2_124_3477_n889), .CO(
        DP_OP_422J2_124_3477_n858), .S(DP_OP_422J2_124_3477_n859) );
  FADDX1_HVT DP_OP_422J2_124_3477_U610 ( .A(DP_OP_422J2_124_3477_n885), .B(
        DP_OP_422J2_124_3477_n881), .CI(DP_OP_422J2_124_3477_n1066), .CO(
        DP_OP_422J2_124_3477_n856), .S(DP_OP_422J2_124_3477_n857) );
  FADDX1_HVT DP_OP_422J2_124_3477_U609 ( .A(DP_OP_422J2_124_3477_n879), .B(
        DP_OP_422J2_124_3477_n1064), .CI(DP_OP_422J2_124_3477_n877), .CO(
        DP_OP_422J2_124_3477_n854), .S(DP_OP_422J2_124_3477_n855) );
  FADDX1_HVT DP_OP_422J2_124_3477_U608 ( .A(DP_OP_422J2_124_3477_n875), .B(
        DP_OP_422J2_124_3477_n1062), .CI(DP_OP_422J2_124_3477_n1058), .CO(
        DP_OP_422J2_124_3477_n852), .S(DP_OP_422J2_124_3477_n853) );
  FADDX1_HVT DP_OP_422J2_124_3477_U607 ( .A(DP_OP_422J2_124_3477_n1060), .B(
        DP_OP_422J2_124_3477_n873), .CI(DP_OP_422J2_124_3477_n1056), .CO(
        DP_OP_422J2_124_3477_n850), .S(DP_OP_422J2_124_3477_n851) );
  FADDX1_HVT DP_OP_422J2_124_3477_U606 ( .A(DP_OP_422J2_124_3477_n871), .B(
        DP_OP_422J2_124_3477_n1054), .CI(DP_OP_422J2_124_3477_n1052), .CO(
        DP_OP_422J2_124_3477_n848), .S(DP_OP_422J2_124_3477_n849) );
  FADDX1_HVT DP_OP_422J2_124_3477_U605 ( .A(DP_OP_422J2_124_3477_n869), .B(
        DP_OP_422J2_124_3477_n1050), .CI(DP_OP_422J2_124_3477_n865), .CO(
        DP_OP_422J2_124_3477_n846), .S(DP_OP_422J2_124_3477_n847) );
  FADDX1_HVT DP_OP_422J2_124_3477_U604 ( .A(DP_OP_422J2_124_3477_n867), .B(
        DP_OP_422J2_124_3477_n1048), .CI(DP_OP_422J2_124_3477_n863), .CO(
        DP_OP_422J2_124_3477_n844), .S(DP_OP_422J2_124_3477_n845) );
  FADDX1_HVT DP_OP_422J2_124_3477_U603 ( .A(DP_OP_422J2_124_3477_n861), .B(
        DP_OP_422J2_124_3477_n1046), .CI(DP_OP_422J2_124_3477_n857), .CO(
        DP_OP_422J2_124_3477_n842), .S(DP_OP_422J2_124_3477_n843) );
  FADDX1_HVT DP_OP_422J2_124_3477_U602 ( .A(DP_OP_422J2_124_3477_n859), .B(
        DP_OP_422J2_124_3477_n1044), .CI(DP_OP_422J2_124_3477_n855), .CO(
        DP_OP_422J2_124_3477_n840), .S(DP_OP_422J2_124_3477_n841) );
  FADDX1_HVT DP_OP_422J2_124_3477_U601 ( .A(DP_OP_422J2_124_3477_n1042), .B(
        DP_OP_422J2_124_3477_n853), .CI(DP_OP_422J2_124_3477_n1040), .CO(
        DP_OP_422J2_124_3477_n838), .S(DP_OP_422J2_124_3477_n839) );
  FADDX1_HVT DP_OP_422J2_124_3477_U600 ( .A(DP_OP_422J2_124_3477_n851), .B(
        DP_OP_422J2_124_3477_n849), .CI(DP_OP_422J2_124_3477_n1038), .CO(
        DP_OP_422J2_124_3477_n836), .S(DP_OP_422J2_124_3477_n837) );
  FADDX1_HVT DP_OP_422J2_124_3477_U599 ( .A(DP_OP_422J2_124_3477_n1036), .B(
        DP_OP_422J2_124_3477_n847), .CI(DP_OP_422J2_124_3477_n1034), .CO(
        DP_OP_422J2_124_3477_n834), .S(DP_OP_422J2_124_3477_n835) );
  FADDX1_HVT DP_OP_422J2_124_3477_U598 ( .A(DP_OP_422J2_124_3477_n845), .B(
        DP_OP_422J2_124_3477_n843), .CI(DP_OP_422J2_124_3477_n1032), .CO(
        DP_OP_422J2_124_3477_n832), .S(DP_OP_422J2_124_3477_n833) );
  FADDX1_HVT DP_OP_422J2_124_3477_U597 ( .A(DP_OP_422J2_124_3477_n841), .B(
        DP_OP_422J2_124_3477_n1030), .CI(DP_OP_422J2_124_3477_n839), .CO(
        DP_OP_422J2_124_3477_n830), .S(DP_OP_422J2_124_3477_n831) );
  FADDX1_HVT DP_OP_422J2_124_3477_U596 ( .A(DP_OP_422J2_124_3477_n1028), .B(
        DP_OP_422J2_124_3477_n837), .CI(DP_OP_422J2_124_3477_n1026), .CO(
        DP_OP_422J2_124_3477_n828), .S(DP_OP_422J2_124_3477_n829) );
  FADDX1_HVT DP_OP_422J2_124_3477_U595 ( .A(DP_OP_422J2_124_3477_n835), .B(
        DP_OP_422J2_124_3477_n1024), .CI(DP_OP_422J2_124_3477_n833), .CO(
        DP_OP_422J2_124_3477_n826), .S(DP_OP_422J2_124_3477_n827) );
  FADDX1_HVT DP_OP_422J2_124_3477_U594 ( .A(DP_OP_422J2_124_3477_n831), .B(
        DP_OP_422J2_124_3477_n1022), .CI(DP_OP_422J2_124_3477_n829), .CO(
        DP_OP_422J2_124_3477_n824), .S(DP_OP_422J2_124_3477_n825) );
  FADDX1_HVT DP_OP_422J2_124_3477_U593 ( .A(DP_OP_422J2_124_3477_n1020), .B(
        DP_OP_422J2_124_3477_n827), .CI(DP_OP_422J2_124_3477_n825), .CO(
        DP_OP_422J2_124_3477_n822), .S(DP_OP_422J2_124_3477_n823) );
  FADDX1_HVT DP_OP_422J2_124_3477_U591 ( .A(DP_OP_422J2_124_3477_n2236), .B(
        DP_OP_422J2_124_3477_n1972), .CI(DP_OP_422J2_124_3477_n1928), .CO(
        DP_OP_422J2_124_3477_n818), .S(DP_OP_422J2_124_3477_n819) );
  FADDX1_HVT DP_OP_422J2_124_3477_U590 ( .A(DP_OP_422J2_124_3477_n2808), .B(
        DP_OP_422J2_124_3477_n2030), .CI(DP_OP_422J2_124_3477_n2294), .CO(
        DP_OP_422J2_124_3477_n816), .S(DP_OP_422J2_124_3477_n817) );
  FADDX1_HVT DP_OP_422J2_124_3477_U589 ( .A(DP_OP_422J2_124_3477_n2280), .B(
        DP_OP_422J2_124_3477_n3040), .CI(DP_OP_422J2_124_3477_n2690), .CO(
        DP_OP_422J2_124_3477_n814), .S(DP_OP_422J2_124_3477_n815) );
  FADDX1_HVT DP_OP_422J2_124_3477_U588 ( .A(DP_OP_422J2_124_3477_n2500), .B(
        DP_OP_422J2_124_3477_n2074), .CI(DP_OP_422J2_124_3477_n2118), .CO(
        DP_OP_422J2_124_3477_n812), .S(DP_OP_422J2_124_3477_n813) );
  FADDX1_HVT DP_OP_422J2_124_3477_U587 ( .A(DP_OP_422J2_124_3477_n2060), .B(
        DP_OP_422J2_124_3477_n2162), .CI(DP_OP_422J2_124_3477_n2206), .CO(
        DP_OP_422J2_124_3477_n810), .S(DP_OP_422J2_124_3477_n811) );
  FADDX1_HVT DP_OP_422J2_124_3477_U586 ( .A(DP_OP_422J2_124_3477_n2764), .B(
        DP_OP_422J2_124_3477_n2866), .CI(DP_OP_422J2_124_3477_n2910), .CO(
        DP_OP_422J2_124_3477_n808), .S(DP_OP_422J2_124_3477_n809) );
  FADDX1_HVT DP_OP_422J2_124_3477_U585 ( .A(DP_OP_422J2_124_3477_n2104), .B(
        DP_OP_422J2_124_3477_n2822), .CI(DP_OP_422J2_124_3477_n2646), .CO(
        DP_OP_422J2_124_3477_n806), .S(DP_OP_422J2_124_3477_n807) );
  FADDX1_HVT DP_OP_422J2_124_3477_U584 ( .A(DP_OP_422J2_124_3477_n2192), .B(
        DP_OP_422J2_124_3477_n2470), .CI(DP_OP_422J2_124_3477_n2998), .CO(
        DP_OP_422J2_124_3477_n804), .S(DP_OP_422J2_124_3477_n805) );
  FADDX1_HVT DP_OP_422J2_124_3477_U583 ( .A(DP_OP_422J2_124_3477_n2720), .B(
        DP_OP_422J2_124_3477_n2954), .CI(DP_OP_422J2_124_3477_n2514), .CO(
        DP_OP_422J2_124_3477_n802), .S(DP_OP_422J2_124_3477_n803) );
  FADDX1_HVT DP_OP_422J2_124_3477_U582 ( .A(DP_OP_422J2_124_3477_n2676), .B(
        DP_OP_422J2_124_3477_n2426), .CI(DP_OP_422J2_124_3477_n2778), .CO(
        DP_OP_422J2_124_3477_n800), .S(DP_OP_422J2_124_3477_n801) );
  FADDX1_HVT DP_OP_422J2_124_3477_U581 ( .A(DP_OP_422J2_124_3477_n2896), .B(
        DP_OP_422J2_124_3477_n2558), .CI(DP_OP_422J2_124_3477_n2382), .CO(
        DP_OP_422J2_124_3477_n798), .S(DP_OP_422J2_124_3477_n799) );
  FADDX1_HVT DP_OP_422J2_124_3477_U580 ( .A(DP_OP_422J2_124_3477_n2368), .B(
        DP_OP_422J2_124_3477_n2338), .CI(DP_OP_422J2_124_3477_n1986), .CO(
        DP_OP_422J2_124_3477_n796), .S(DP_OP_422J2_124_3477_n797) );
  FADDX1_HVT DP_OP_422J2_124_3477_U579 ( .A(DP_OP_422J2_124_3477_n2588), .B(
        DP_OP_422J2_124_3477_n2250), .CI(DP_OP_422J2_124_3477_n2602), .CO(
        DP_OP_422J2_124_3477_n794), .S(DP_OP_422J2_124_3477_n795) );
  FADDX1_HVT DP_OP_422J2_124_3477_U578 ( .A(DP_OP_422J2_124_3477_n2544), .B(
        DP_OP_422J2_124_3477_n2412), .CI(DP_OP_422J2_124_3477_n2734), .CO(
        DP_OP_422J2_124_3477_n792), .S(DP_OP_422J2_124_3477_n793) );
  FADDX1_HVT DP_OP_422J2_124_3477_U577 ( .A(DP_OP_422J2_124_3477_n2852), .B(
        DP_OP_422J2_124_3477_n2148), .CI(DP_OP_422J2_124_3477_n2324), .CO(
        DP_OP_422J2_124_3477_n790), .S(DP_OP_422J2_124_3477_n791) );
  FADDX1_HVT DP_OP_422J2_124_3477_U576 ( .A(DP_OP_422J2_124_3477_n2016), .B(
        DP_OP_422J2_124_3477_n2632), .CI(DP_OP_422J2_124_3477_n2984), .CO(
        DP_OP_422J2_124_3477_n788), .S(DP_OP_422J2_124_3477_n789) );
  FADDX1_HVT DP_OP_422J2_124_3477_U575 ( .A(DP_OP_422J2_124_3477_n2940), .B(
        DP_OP_422J2_124_3477_n2456), .CI(DP_OP_422J2_124_3477_n821), .CO(
        DP_OP_422J2_124_3477_n786), .S(DP_OP_422J2_124_3477_n787) );
  FADDX1_HVT DP_OP_422J2_124_3477_U574 ( .A(DP_OP_422J2_124_3477_n2287), .B(
        DP_OP_422J2_124_3477_n2023), .CI(DP_OP_422J2_124_3477_n1979), .CO(
        DP_OP_422J2_124_3477_n784), .S(DP_OP_422J2_124_3477_n785) );
  FADDX1_HVT DP_OP_422J2_124_3477_U573 ( .A(DP_OP_422J2_124_3477_n3033), .B(
        DP_OP_422J2_124_3477_n2067), .CI(DP_OP_422J2_124_3477_n2111), .CO(
        DP_OP_422J2_124_3477_n782), .S(DP_OP_422J2_124_3477_n783) );
  FADDX1_HVT DP_OP_422J2_124_3477_U572 ( .A(DP_OP_422J2_124_3477_n2991), .B(
        DP_OP_422J2_124_3477_n2155), .CI(DP_OP_422J2_124_3477_n2199), .CO(
        DP_OP_422J2_124_3477_n780), .S(DP_OP_422J2_124_3477_n781) );
  FADDX1_HVT DP_OP_422J2_124_3477_U571 ( .A(DP_OP_422J2_124_3477_n2947), .B(
        DP_OP_422J2_124_3477_n2243), .CI(DP_OP_422J2_124_3477_n2331), .CO(
        DP_OP_422J2_124_3477_n778), .S(DP_OP_422J2_124_3477_n779) );
  FADDX1_HVT DP_OP_422J2_124_3477_U570 ( .A(DP_OP_422J2_124_3477_n2903), .B(
        DP_OP_422J2_124_3477_n2375), .CI(DP_OP_422J2_124_3477_n2419), .CO(
        DP_OP_422J2_124_3477_n776), .S(DP_OP_422J2_124_3477_n777) );
  FADDX1_HVT DP_OP_422J2_124_3477_U569 ( .A(DP_OP_422J2_124_3477_n2859), .B(
        DP_OP_422J2_124_3477_n2463), .CI(DP_OP_422J2_124_3477_n2507), .CO(
        DP_OP_422J2_124_3477_n774), .S(DP_OP_422J2_124_3477_n775) );
  FADDX1_HVT DP_OP_422J2_124_3477_U568 ( .A(DP_OP_422J2_124_3477_n2815), .B(
        DP_OP_422J2_124_3477_n2551), .CI(DP_OP_422J2_124_3477_n2595), .CO(
        DP_OP_422J2_124_3477_n772), .S(DP_OP_422J2_124_3477_n773) );
  FADDX1_HVT DP_OP_422J2_124_3477_U567 ( .A(DP_OP_422J2_124_3477_n2771), .B(
        DP_OP_422J2_124_3477_n2639), .CI(DP_OP_422J2_124_3477_n2683), .CO(
        DP_OP_422J2_124_3477_n770), .S(DP_OP_422J2_124_3477_n771) );
  FADDX1_HVT DP_OP_422J2_124_3477_U566 ( .A(DP_OP_422J2_124_3477_n2727), .B(
        DP_OP_422J2_124_3477_n1016), .CI(DP_OP_422J2_124_3477_n1014), .CO(
        DP_OP_422J2_124_3477_n768), .S(DP_OP_422J2_124_3477_n769) );
  FADDX1_HVT DP_OP_422J2_124_3477_U565 ( .A(DP_OP_422J2_124_3477_n1012), .B(
        DP_OP_422J2_124_3477_n984), .CI(DP_OP_422J2_124_3477_n986), .CO(
        DP_OP_422J2_124_3477_n766), .S(DP_OP_422J2_124_3477_n767) );
  FADDX1_HVT DP_OP_422J2_124_3477_U564 ( .A(DP_OP_422J2_124_3477_n1010), .B(
        DP_OP_422J2_124_3477_n988), .CI(DP_OP_422J2_124_3477_n990), .CO(
        DP_OP_422J2_124_3477_n764), .S(DP_OP_422J2_124_3477_n765) );
  FADDX1_HVT DP_OP_422J2_124_3477_U563 ( .A(DP_OP_422J2_124_3477_n1008), .B(
        DP_OP_422J2_124_3477_n992), .CI(DP_OP_422J2_124_3477_n994), .CO(
        DP_OP_422J2_124_3477_n762), .S(DP_OP_422J2_124_3477_n763) );
  FADDX1_HVT DP_OP_422J2_124_3477_U562 ( .A(DP_OP_422J2_124_3477_n1000), .B(
        DP_OP_422J2_124_3477_n1006), .CI(DP_OP_422J2_124_3477_n996), .CO(
        DP_OP_422J2_124_3477_n760), .S(DP_OP_422J2_124_3477_n761) );
  FADDX1_HVT DP_OP_422J2_124_3477_U561 ( .A(DP_OP_422J2_124_3477_n998), .B(
        DP_OP_422J2_124_3477_n1002), .CI(DP_OP_422J2_124_3477_n1004), .CO(
        DP_OP_422J2_124_3477_n758), .S(DP_OP_422J2_124_3477_n759) );
  FADDX1_HVT DP_OP_422J2_124_3477_U560 ( .A(DP_OP_422J2_124_3477_n950), .B(
        DP_OP_422J2_124_3477_n980), .CI(DP_OP_422J2_124_3477_n982), .CO(
        DP_OP_422J2_124_3477_n756), .S(DP_OP_422J2_124_3477_n757) );
  FADDX1_HVT DP_OP_422J2_124_3477_U559 ( .A(DP_OP_422J2_124_3477_n964), .B(
        DP_OP_422J2_124_3477_n952), .CI(DP_OP_422J2_124_3477_n954), .CO(
        DP_OP_422J2_124_3477_n754), .S(DP_OP_422J2_124_3477_n755) );
  FADDX1_HVT DP_OP_422J2_124_3477_U557 ( .A(DP_OP_422J2_124_3477_n960), .B(
        DP_OP_422J2_124_3477_n978), .CI(DP_OP_422J2_124_3477_n976), .CO(
        DP_OP_422J2_124_3477_n750), .S(DP_OP_422J2_124_3477_n751) );
  FADDX1_HVT DP_OP_422J2_124_3477_U556 ( .A(DP_OP_422J2_124_3477_n970), .B(
        DP_OP_422J2_124_3477_n966), .CI(DP_OP_422J2_124_3477_n968), .CO(
        DP_OP_422J2_124_3477_n748), .S(DP_OP_422J2_124_3477_n749) );
  FADDX1_HVT DP_OP_422J2_124_3477_U555 ( .A(DP_OP_422J2_124_3477_n974), .B(
        DP_OP_422J2_124_3477_n972), .CI(DP_OP_422J2_124_3477_n813), .CO(
        DP_OP_422J2_124_3477_n746), .S(DP_OP_422J2_124_3477_n747) );
  FADDX1_HVT DP_OP_422J2_124_3477_U554 ( .A(DP_OP_422J2_124_3477_n809), .B(
        DP_OP_422J2_124_3477_n805), .CI(DP_OP_422J2_124_3477_n787), .CO(
        DP_OP_422J2_124_3477_n744), .S(DP_OP_422J2_124_3477_n745) );
  FADDX1_HVT DP_OP_422J2_124_3477_U553 ( .A(DP_OP_422J2_124_3477_n811), .B(
        DP_OP_422J2_124_3477_n793), .CI(DP_OP_422J2_124_3477_n791), .CO(
        DP_OP_422J2_124_3477_n742), .S(DP_OP_422J2_124_3477_n743) );
  FADDX1_HVT DP_OP_422J2_124_3477_U552 ( .A(DP_OP_422J2_124_3477_n803), .B(
        DP_OP_422J2_124_3477_n807), .CI(DP_OP_422J2_124_3477_n799), .CO(
        DP_OP_422J2_124_3477_n740), .S(DP_OP_422J2_124_3477_n741) );
  FADDX1_HVT DP_OP_422J2_124_3477_U551 ( .A(DP_OP_422J2_124_3477_n815), .B(
        DP_OP_422J2_124_3477_n795), .CI(DP_OP_422J2_124_3477_n789), .CO(
        DP_OP_422J2_124_3477_n738), .S(DP_OP_422J2_124_3477_n739) );
  FADDX1_HVT DP_OP_422J2_124_3477_U550 ( .A(DP_OP_422J2_124_3477_n797), .B(
        DP_OP_422J2_124_3477_n819), .CI(DP_OP_422J2_124_3477_n817), .CO(
        DP_OP_422J2_124_3477_n736), .S(DP_OP_422J2_124_3477_n737) );
  FADDX1_HVT DP_OP_422J2_124_3477_U549 ( .A(DP_OP_422J2_124_3477_n801), .B(
        DP_OP_422J2_124_3477_n781), .CI(DP_OP_422J2_124_3477_n777), .CO(
        DP_OP_422J2_124_3477_n734), .S(DP_OP_422J2_124_3477_n735) );
  FADDX1_HVT DP_OP_422J2_124_3477_U548 ( .A(DP_OP_422J2_124_3477_n773), .B(
        DP_OP_422J2_124_3477_n771), .CI(DP_OP_422J2_124_3477_n783), .CO(
        DP_OP_422J2_124_3477_n732), .S(DP_OP_422J2_124_3477_n733) );
  FADDX1_HVT DP_OP_422J2_124_3477_U547 ( .A(DP_OP_422J2_124_3477_n779), .B(
        DP_OP_422J2_124_3477_n775), .CI(DP_OP_422J2_124_3477_n785), .CO(
        DP_OP_422J2_124_3477_n730), .S(DP_OP_422J2_124_3477_n731) );
  FADDX1_HVT DP_OP_422J2_124_3477_U546 ( .A(DP_OP_422J2_124_3477_n948), .B(
        DP_OP_422J2_124_3477_n944), .CI(DP_OP_422J2_124_3477_n946), .CO(
        DP_OP_422J2_124_3477_n728), .S(DP_OP_422J2_124_3477_n729) );
  FADDX1_HVT DP_OP_422J2_124_3477_U545 ( .A(DP_OP_422J2_124_3477_n942), .B(
        DP_OP_422J2_124_3477_n928), .CI(DP_OP_422J2_124_3477_n930), .CO(
        DP_OP_422J2_124_3477_n726), .S(DP_OP_422J2_124_3477_n727) );
  FADDX1_HVT DP_OP_422J2_124_3477_U544 ( .A(DP_OP_422J2_124_3477_n940), .B(
        DP_OP_422J2_124_3477_n932), .CI(DP_OP_422J2_124_3477_n938), .CO(
        DP_OP_422J2_124_3477_n724), .S(DP_OP_422J2_124_3477_n725) );
  FADDX1_HVT DP_OP_422J2_124_3477_U543 ( .A(DP_OP_422J2_124_3477_n936), .B(
        DP_OP_422J2_124_3477_n934), .CI(DP_OP_422J2_124_3477_n769), .CO(
        DP_OP_422J2_124_3477_n722), .S(DP_OP_422J2_124_3477_n723) );
  FADDX1_HVT DP_OP_422J2_124_3477_U542 ( .A(DP_OP_422J2_124_3477_n926), .B(
        DP_OP_422J2_124_3477_n767), .CI(DP_OP_422J2_124_3477_n765), .CO(
        DP_OP_422J2_124_3477_n720), .S(DP_OP_422J2_124_3477_n721) );
  FADDX1_HVT DP_OP_422J2_124_3477_U541 ( .A(DP_OP_422J2_124_3477_n924), .B(
        DP_OP_422J2_124_3477_n761), .CI(DP_OP_422J2_124_3477_n763), .CO(
        DP_OP_422J2_124_3477_n718), .S(DP_OP_422J2_124_3477_n719) );
  FADDX1_HVT DP_OP_422J2_124_3477_U540 ( .A(DP_OP_422J2_124_3477_n922), .B(
        DP_OP_422J2_124_3477_n759), .CI(DP_OP_422J2_124_3477_n916), .CO(
        DP_OP_422J2_124_3477_n716), .S(DP_OP_422J2_124_3477_n717) );
  FADDX1_HVT DP_OP_422J2_124_3477_U539 ( .A(DP_OP_422J2_124_3477_n920), .B(
        DP_OP_422J2_124_3477_n918), .CI(DP_OP_422J2_124_3477_n906), .CO(
        DP_OP_422J2_124_3477_n714), .S(DP_OP_422J2_124_3477_n715) );
  FADDX1_HVT DP_OP_422J2_124_3477_U538 ( .A(DP_OP_422J2_124_3477_n914), .B(
        DP_OP_422J2_124_3477_n757), .CI(DP_OP_422J2_124_3477_n747), .CO(
        DP_OP_422J2_124_3477_n712), .S(DP_OP_422J2_124_3477_n713) );
  FADDX1_HVT DP_OP_422J2_124_3477_U537 ( .A(DP_OP_422J2_124_3477_n912), .B(
        DP_OP_422J2_124_3477_n753), .CI(DP_OP_422J2_124_3477_n749), .CO(
        DP_OP_422J2_124_3477_n710), .S(DP_OP_422J2_124_3477_n711) );
  FADDX1_HVT DP_OP_422J2_124_3477_U536 ( .A(DP_OP_422J2_124_3477_n910), .B(
        DP_OP_422J2_124_3477_n755), .CI(DP_OP_422J2_124_3477_n751), .CO(
        DP_OP_422J2_124_3477_n708), .S(DP_OP_422J2_124_3477_n709) );
  FADDX1_HVT DP_OP_422J2_124_3477_U535 ( .A(DP_OP_422J2_124_3477_n908), .B(
        DP_OP_422J2_124_3477_n743), .CI(DP_OP_422J2_124_3477_n739), .CO(
        DP_OP_422J2_124_3477_n706), .S(DP_OP_422J2_124_3477_n707) );
  FADDX1_HVT DP_OP_422J2_124_3477_U534 ( .A(DP_OP_422J2_124_3477_n741), .B(
        DP_OP_422J2_124_3477_n735), .CI(DP_OP_422J2_124_3477_n904), .CO(
        DP_OP_422J2_124_3477_n704), .S(DP_OP_422J2_124_3477_n705) );
  FADDX1_HVT DP_OP_422J2_124_3477_U533 ( .A(DP_OP_422J2_124_3477_n737), .B(
        DP_OP_422J2_124_3477_n745), .CI(DP_OP_422J2_124_3477_n731), .CO(
        DP_OP_422J2_124_3477_n702), .S(DP_OP_422J2_124_3477_n703) );
  FADDX1_HVT DP_OP_422J2_124_3477_U532 ( .A(DP_OP_422J2_124_3477_n733), .B(
        DP_OP_422J2_124_3477_n902), .CI(DP_OP_422J2_124_3477_n900), .CO(
        DP_OP_422J2_124_3477_n700), .S(DP_OP_422J2_124_3477_n701) );
  FADDX1_HVT DP_OP_422J2_124_3477_U531 ( .A(DP_OP_422J2_124_3477_n729), .B(
        DP_OP_422J2_124_3477_n898), .CI(DP_OP_422J2_124_3477_n896), .CO(
        DP_OP_422J2_124_3477_n698), .S(DP_OP_422J2_124_3477_n699) );
  FADDX1_HVT DP_OP_422J2_124_3477_U530 ( .A(DP_OP_422J2_124_3477_n894), .B(
        DP_OP_422J2_124_3477_n892), .CI(DP_OP_422J2_124_3477_n890), .CO(
        DP_OP_422J2_124_3477_n696), .S(DP_OP_422J2_124_3477_n697) );
  FADDX1_HVT DP_OP_422J2_124_3477_U529 ( .A(DP_OP_422J2_124_3477_n888), .B(
        DP_OP_422J2_124_3477_n723), .CI(DP_OP_422J2_124_3477_n882), .CO(
        DP_OP_422J2_124_3477_n694), .S(DP_OP_422J2_124_3477_n695) );
  FADDX1_HVT DP_OP_422J2_124_3477_U528 ( .A(DP_OP_422J2_124_3477_n886), .B(
        DP_OP_422J2_124_3477_n725), .CI(DP_OP_422J2_124_3477_n727), .CO(
        DP_OP_422J2_124_3477_n692), .S(DP_OP_422J2_124_3477_n693) );
  FADDX1_HVT DP_OP_422J2_124_3477_U527 ( .A(DP_OP_422J2_124_3477_n884), .B(
        DP_OP_422J2_124_3477_n721), .CI(DP_OP_422J2_124_3477_n717), .CO(
        DP_OP_422J2_124_3477_n690), .S(DP_OP_422J2_124_3477_n691) );
  FADDX1_HVT DP_OP_422J2_124_3477_U526 ( .A(DP_OP_422J2_124_3477_n880), .B(
        DP_OP_422J2_124_3477_n719), .CI(DP_OP_422J2_124_3477_n715), .CO(
        DP_OP_422J2_124_3477_n688), .S(DP_OP_422J2_124_3477_n689) );
  FADDX1_HVT DP_OP_422J2_124_3477_U525 ( .A(DP_OP_422J2_124_3477_n878), .B(
        DP_OP_422J2_124_3477_n711), .CI(DP_OP_422J2_124_3477_n876), .CO(
        DP_OP_422J2_124_3477_n686), .S(DP_OP_422J2_124_3477_n687) );
  FADDX1_HVT DP_OP_422J2_124_3477_U524 ( .A(DP_OP_422J2_124_3477_n709), .B(
        DP_OP_422J2_124_3477_n713), .CI(DP_OP_422J2_124_3477_n874), .CO(
        DP_OP_422J2_124_3477_n684), .S(DP_OP_422J2_124_3477_n685) );
  FADDX1_HVT DP_OP_422J2_124_3477_U523 ( .A(DP_OP_422J2_124_3477_n707), .B(
        DP_OP_422J2_124_3477_n872), .CI(DP_OP_422J2_124_3477_n703), .CO(
        DP_OP_422J2_124_3477_n682), .S(DP_OP_422J2_124_3477_n683) );
  FADDX1_HVT DP_OP_422J2_124_3477_U522 ( .A(DP_OP_422J2_124_3477_n705), .B(
        DP_OP_422J2_124_3477_n870), .CI(DP_OP_422J2_124_3477_n701), .CO(
        DP_OP_422J2_124_3477_n680), .S(DP_OP_422J2_124_3477_n681) );
  FADDX1_HVT DP_OP_422J2_124_3477_U521 ( .A(DP_OP_422J2_124_3477_n868), .B(
        DP_OP_422J2_124_3477_n866), .CI(DP_OP_422J2_124_3477_n699), .CO(
        DP_OP_422J2_124_3477_n678), .S(DP_OP_422J2_124_3477_n679) );
  FADDX1_HVT DP_OP_422J2_124_3477_U520 ( .A(DP_OP_422J2_124_3477_n864), .B(
        DP_OP_422J2_124_3477_n862), .CI(DP_OP_422J2_124_3477_n697), .CO(
        DP_OP_422J2_124_3477_n676), .S(DP_OP_422J2_124_3477_n677) );
  FADDX1_HVT DP_OP_422J2_124_3477_U519 ( .A(DP_OP_422J2_124_3477_n860), .B(
        DP_OP_422J2_124_3477_n693), .CI(DP_OP_422J2_124_3477_n856), .CO(
        DP_OP_422J2_124_3477_n674), .S(DP_OP_422J2_124_3477_n675) );
  FADDX1_HVT DP_OP_422J2_124_3477_U518 ( .A(DP_OP_422J2_124_3477_n858), .B(
        DP_OP_422J2_124_3477_n695), .CI(DP_OP_422J2_124_3477_n691), .CO(
        DP_OP_422J2_124_3477_n672), .S(DP_OP_422J2_124_3477_n673) );
  FADDX1_HVT DP_OP_422J2_124_3477_U516 ( .A(DP_OP_422J2_124_3477_n685), .B(
        DP_OP_422J2_124_3477_n852), .CI(DP_OP_422J2_124_3477_n683), .CO(
        DP_OP_422J2_124_3477_n668), .S(DP_OP_422J2_124_3477_n669) );
  FADDX1_HVT DP_OP_422J2_124_3477_U515 ( .A(DP_OP_422J2_124_3477_n850), .B(
        DP_OP_422J2_124_3477_n681), .CI(DP_OP_422J2_124_3477_n848), .CO(
        DP_OP_422J2_124_3477_n666), .S(DP_OP_422J2_124_3477_n667) );
  FADDX1_HVT DP_OP_422J2_124_3477_U514 ( .A(DP_OP_422J2_124_3477_n679), .B(
        DP_OP_422J2_124_3477_n846), .CI(DP_OP_422J2_124_3477_n844), .CO(
        DP_OP_422J2_124_3477_n664), .S(DP_OP_422J2_124_3477_n665) );
  FADDX1_HVT DP_OP_422J2_124_3477_U513 ( .A(DP_OP_422J2_124_3477_n677), .B(
        DP_OP_422J2_124_3477_n842), .CI(DP_OP_422J2_124_3477_n675), .CO(
        DP_OP_422J2_124_3477_n662), .S(DP_OP_422J2_124_3477_n663) );
  FADDX1_HVT DP_OP_422J2_124_3477_U512 ( .A(DP_OP_422J2_124_3477_n673), .B(
        DP_OP_422J2_124_3477_n840), .CI(DP_OP_422J2_124_3477_n671), .CO(
        DP_OP_422J2_124_3477_n660), .S(DP_OP_422J2_124_3477_n661) );
  FADDX1_HVT DP_OP_422J2_124_3477_U511 ( .A(DP_OP_422J2_124_3477_n838), .B(
        DP_OP_422J2_124_3477_n669), .CI(DP_OP_422J2_124_3477_n836), .CO(
        DP_OP_422J2_124_3477_n658), .S(DP_OP_422J2_124_3477_n659) );
  FADDX1_HVT DP_OP_422J2_124_3477_U509 ( .A(DP_OP_422J2_124_3477_n832), .B(
        DP_OP_422J2_124_3477_n663), .CI(DP_OP_422J2_124_3477_n661), .CO(
        DP_OP_422J2_124_3477_n654), .S(DP_OP_422J2_124_3477_n655) );
  FADDX1_HVT DP_OP_422J2_124_3477_U508 ( .A(DP_OP_422J2_124_3477_n830), .B(
        DP_OP_422J2_124_3477_n659), .CI(DP_OP_422J2_124_3477_n828), .CO(
        DP_OP_422J2_124_3477_n652), .S(DP_OP_422J2_124_3477_n653) );
  FADDX1_HVT DP_OP_422J2_124_3477_U507 ( .A(DP_OP_422J2_124_3477_n657), .B(
        DP_OP_422J2_124_3477_n826), .CI(DP_OP_422J2_124_3477_n655), .CO(
        DP_OP_422J2_124_3477_n650), .S(DP_OP_422J2_124_3477_n651) );
  FADDX1_HVT DP_OP_422J2_124_3477_U506 ( .A(DP_OP_422J2_124_3477_n824), .B(
        DP_OP_422J2_124_3477_n653), .CI(DP_OP_422J2_124_3477_n651), .CO(
        DP_OP_422J2_124_3477_n648), .S(DP_OP_422J2_124_3477_n649) );
  FADDX1_HVT DP_OP_422J2_124_3477_U505 ( .A(DP_OP_422J2_124_3477_n3027), .B(
        DP_OP_422J2_124_3477_n1971), .CI(DP_OP_422J2_124_3477_n1927), .CO(
        DP_OP_422J2_124_3477_n646), .S(DP_OP_422J2_124_3477_n647) );
  FADDX1_HVT DP_OP_422J2_124_3477_U504 ( .A(DP_OP_422J2_124_3477_n820), .B(
        DP_OP_422J2_124_3477_n2286), .CI(DP_OP_422J2_124_3477_n1978), .CO(
        DP_OP_422J2_124_3477_n644), .S(DP_OP_422J2_124_3477_n645) );
  FADDX1_HVT DP_OP_422J2_124_3477_U503 ( .A(DP_OP_422J2_124_3477_n2367), .B(
        DP_OP_422J2_124_3477_n3032), .CI(DP_OP_422J2_124_3477_n2682), .CO(
        DP_OP_422J2_124_3477_n642), .S(DP_OP_422J2_124_3477_n643) );
  FADDX1_HVT DP_OP_422J2_124_3477_U502 ( .A(DP_OP_422J2_124_3477_n2059), .B(
        DP_OP_422J2_124_3477_n2594), .CI(DP_OP_422J2_124_3477_n2814), .CO(
        DP_OP_422J2_124_3477_n640), .S(DP_OP_422J2_124_3477_n641) );
  FADDX1_HVT DP_OP_422J2_124_3477_U501 ( .A(DP_OP_422J2_124_3477_n2279), .B(
        DP_OP_422J2_124_3477_n2374), .CI(DP_OP_422J2_124_3477_n2990), .CO(
        DP_OP_422J2_124_3477_n638), .S(DP_OP_422J2_124_3477_n639) );
  FADDX1_HVT DP_OP_422J2_124_3477_U500 ( .A(DP_OP_422J2_124_3477_n2015), .B(
        DP_OP_422J2_124_3477_n2902), .CI(DP_OP_422J2_124_3477_n2066), .CO(
        DP_OP_422J2_124_3477_n636), .S(DP_OP_422J2_124_3477_n637) );
  FADDX1_HVT DP_OP_422J2_124_3477_U499 ( .A(DP_OP_422J2_124_3477_n2147), .B(
        DP_OP_422J2_124_3477_n2022), .CI(DP_OP_422J2_124_3477_n2858), .CO(
        DP_OP_422J2_124_3477_n634), .S(DP_OP_422J2_124_3477_n635) );
  FADDX1_HVT DP_OP_422J2_124_3477_U498 ( .A(DP_OP_422J2_124_3477_n2983), .B(
        DP_OP_422J2_124_3477_n2418), .CI(DP_OP_422J2_124_3477_n2506), .CO(
        DP_OP_422J2_124_3477_n632), .S(DP_OP_422J2_124_3477_n633) );
  FADDX1_HVT DP_OP_422J2_124_3477_U497 ( .A(DP_OP_422J2_124_3477_n2499), .B(
        DP_OP_422J2_124_3477_n2550), .CI(DP_OP_422J2_124_3477_n2946), .CO(
        DP_OP_422J2_124_3477_n630), .S(DP_OP_422J2_124_3477_n631) );
  FADDX1_HVT DP_OP_422J2_124_3477_U496 ( .A(DP_OP_422J2_124_3477_n2763), .B(
        DP_OP_422J2_124_3477_n2242), .CI(DP_OP_422J2_124_3477_n2770), .CO(
        DP_OP_422J2_124_3477_n628), .S(DP_OP_422J2_124_3477_n629) );
  FADDX1_HVT DP_OP_422J2_124_3477_U495 ( .A(DP_OP_422J2_124_3477_n2939), .B(
        DP_OP_422J2_124_3477_n2462), .CI(DP_OP_422J2_124_3477_n2638), .CO(
        DP_OP_422J2_124_3477_n626), .S(DP_OP_422J2_124_3477_n627) );
  FADDX1_HVT DP_OP_422J2_124_3477_U494 ( .A(DP_OP_422J2_124_3477_n2235), .B(
        DP_OP_422J2_124_3477_n2110), .CI(DP_OP_422J2_124_3477_n2726), .CO(
        DP_OP_422J2_124_3477_n624), .S(DP_OP_422J2_124_3477_n625) );
  FADDX1_HVT DP_OP_422J2_124_3477_U493 ( .A(DP_OP_422J2_124_3477_n2191), .B(
        DP_OP_422J2_124_3477_n2330), .CI(DP_OP_422J2_124_3477_n2198), .CO(
        DP_OP_422J2_124_3477_n622), .S(DP_OP_422J2_124_3477_n623) );
  FADDX1_HVT DP_OP_422J2_124_3477_U492 ( .A(DP_OP_422J2_124_3477_n2587), .B(
        DP_OP_422J2_124_3477_n2411), .CI(DP_OP_422J2_124_3477_n2154), .CO(
        DP_OP_422J2_124_3477_n620), .S(DP_OP_422J2_124_3477_n621) );
  FADDX1_HVT DP_OP_422J2_124_3477_U491 ( .A(DP_OP_422J2_124_3477_n2895), .B(
        DP_OP_422J2_124_3477_n2103), .CI(DP_OP_422J2_124_3477_n2323), .CO(
        DP_OP_422J2_124_3477_n618), .S(DP_OP_422J2_124_3477_n619) );
  FADDX1_HVT DP_OP_422J2_124_3477_U490 ( .A(DP_OP_422J2_124_3477_n2851), .B(
        DP_OP_422J2_124_3477_n2455), .CI(DP_OP_422J2_124_3477_n2543), .CO(
        DP_OP_422J2_124_3477_n616), .S(DP_OP_422J2_124_3477_n617) );
  FADDX1_HVT DP_OP_422J2_124_3477_U489 ( .A(DP_OP_422J2_124_3477_n2807), .B(
        DP_OP_422J2_124_3477_n2631), .CI(DP_OP_422J2_124_3477_n2675), .CO(
        DP_OP_422J2_124_3477_n614), .S(DP_OP_422J2_124_3477_n615) );
  FADDX1_HVT DP_OP_422J2_124_3477_U488 ( .A(DP_OP_422J2_124_3477_n2719), .B(
        DP_OP_422J2_124_3477_n818), .CI(DP_OP_422J2_124_3477_n816), .CO(
        DP_OP_422J2_124_3477_n612), .S(DP_OP_422J2_124_3477_n613) );
  FADDX1_HVT DP_OP_422J2_124_3477_U487 ( .A(DP_OP_422J2_124_3477_n786), .B(
        DP_OP_422J2_124_3477_n814), .CI(DP_OP_422J2_124_3477_n788), .CO(
        DP_OP_422J2_124_3477_n610), .S(DP_OP_422J2_124_3477_n611) );
  FADDX1_HVT DP_OP_422J2_124_3477_U486 ( .A(DP_OP_422J2_124_3477_n812), .B(
        DP_OP_422J2_124_3477_n790), .CI(DP_OP_422J2_124_3477_n792), .CO(
        DP_OP_422J2_124_3477_n608), .S(DP_OP_422J2_124_3477_n609) );
  FADDX1_HVT DP_OP_422J2_124_3477_U485 ( .A(DP_OP_422J2_124_3477_n810), .B(
        DP_OP_422J2_124_3477_n794), .CI(DP_OP_422J2_124_3477_n796), .CO(
        DP_OP_422J2_124_3477_n606), .S(DP_OP_422J2_124_3477_n607) );
  FADDX1_HVT DP_OP_422J2_124_3477_U484 ( .A(DP_OP_422J2_124_3477_n808), .B(
        DP_OP_422J2_124_3477_n798), .CI(DP_OP_422J2_124_3477_n800), .CO(
        DP_OP_422J2_124_3477_n604), .S(DP_OP_422J2_124_3477_n605) );
  FADDX1_HVT DP_OP_422J2_124_3477_U483 ( .A(DP_OP_422J2_124_3477_n806), .B(
        DP_OP_422J2_124_3477_n802), .CI(DP_OP_422J2_124_3477_n804), .CO(
        DP_OP_422J2_124_3477_n602), .S(DP_OP_422J2_124_3477_n603) );
  FADDX1_HVT DP_OP_422J2_124_3477_U482 ( .A(DP_OP_422J2_124_3477_n784), .B(
        DP_OP_422J2_124_3477_n770), .CI(DP_OP_422J2_124_3477_n782), .CO(
        DP_OP_422J2_124_3477_n600), .S(DP_OP_422J2_124_3477_n601) );
  FADDX1_HVT DP_OP_422J2_124_3477_U481 ( .A(DP_OP_422J2_124_3477_n776), .B(
        DP_OP_422J2_124_3477_n772), .CI(DP_OP_422J2_124_3477_n774), .CO(
        DP_OP_422J2_124_3477_n598), .S(DP_OP_422J2_124_3477_n599) );
  FADDX1_HVT DP_OP_422J2_124_3477_U480 ( .A(DP_OP_422J2_124_3477_n780), .B(
        DP_OP_422J2_124_3477_n778), .CI(DP_OP_422J2_124_3477_n645), .CO(
        DP_OP_422J2_124_3477_n596), .S(DP_OP_422J2_124_3477_n597) );
  FADDX1_HVT DP_OP_422J2_124_3477_U479 ( .A(DP_OP_422J2_124_3477_n647), .B(
        DP_OP_422J2_124_3477_n633), .CI(DP_OP_422J2_124_3477_n639), .CO(
        DP_OP_422J2_124_3477_n594), .S(DP_OP_422J2_124_3477_n595) );
  FADDX1_HVT DP_OP_422J2_124_3477_U478 ( .A(DP_OP_422J2_124_3477_n615), .B(
        DP_OP_422J2_124_3477_n637), .CI(DP_OP_422J2_124_3477_n635), .CO(
        DP_OP_422J2_124_3477_n592), .S(DP_OP_422J2_124_3477_n593) );
  FADDX1_HVT DP_OP_422J2_124_3477_U477 ( .A(DP_OP_422J2_124_3477_n641), .B(
        DP_OP_422J2_124_3477_n623), .CI(DP_OP_422J2_124_3477_n625), .CO(
        DP_OP_422J2_124_3477_n590), .S(DP_OP_422J2_124_3477_n591) );
  FADDX1_HVT DP_OP_422J2_124_3477_U476 ( .A(DP_OP_422J2_124_3477_n627), .B(
        DP_OP_422J2_124_3477_n617), .CI(DP_OP_422J2_124_3477_n619), .CO(
        DP_OP_422J2_124_3477_n588), .S(DP_OP_422J2_124_3477_n589) );
  FADDX1_HVT DP_OP_422J2_124_3477_U475 ( .A(DP_OP_422J2_124_3477_n621), .B(
        DP_OP_422J2_124_3477_n643), .CI(DP_OP_422J2_124_3477_n631), .CO(
        DP_OP_422J2_124_3477_n586), .S(DP_OP_422J2_124_3477_n587) );
  FADDX1_HVT DP_OP_422J2_124_3477_U474 ( .A(DP_OP_422J2_124_3477_n629), .B(
        DP_OP_422J2_124_3477_n768), .CI(DP_OP_422J2_124_3477_n766), .CO(
        DP_OP_422J2_124_3477_n584), .S(DP_OP_422J2_124_3477_n585) );
  FADDX1_HVT DP_OP_422J2_124_3477_U473 ( .A(DP_OP_422J2_124_3477_n764), .B(
        DP_OP_422J2_124_3477_n758), .CI(DP_OP_422J2_124_3477_n760), .CO(
        DP_OP_422J2_124_3477_n582), .S(DP_OP_422J2_124_3477_n583) );
  FADDX1_HVT DP_OP_422J2_124_3477_U472 ( .A(DP_OP_422J2_124_3477_n762), .B(
        DP_OP_422J2_124_3477_n756), .CI(DP_OP_422J2_124_3477_n754), .CO(
        DP_OP_422J2_124_3477_n580), .S(DP_OP_422J2_124_3477_n581) );
  FADDX1_HVT DP_OP_422J2_124_3477_U471 ( .A(DP_OP_422J2_124_3477_n752), .B(
        DP_OP_422J2_124_3477_n748), .CI(DP_OP_422J2_124_3477_n746), .CO(
        DP_OP_422J2_124_3477_n578), .S(DP_OP_422J2_124_3477_n579) );
  FADDX1_HVT DP_OP_422J2_124_3477_U470 ( .A(DP_OP_422J2_124_3477_n750), .B(
        DP_OP_422J2_124_3477_n613), .CI(DP_OP_422J2_124_3477_n607), .CO(
        DP_OP_422J2_124_3477_n576), .S(DP_OP_422J2_124_3477_n577) );
  FADDX1_HVT DP_OP_422J2_124_3477_U469 ( .A(DP_OP_422J2_124_3477_n609), .B(
        DP_OP_422J2_124_3477_n603), .CI(DP_OP_422J2_124_3477_n734), .CO(
        DP_OP_422J2_124_3477_n574), .S(DP_OP_422J2_124_3477_n575) );
  FADDX1_HVT DP_OP_422J2_124_3477_U468 ( .A(DP_OP_422J2_124_3477_n744), .B(
        DP_OP_422J2_124_3477_n611), .CI(DP_OP_422J2_124_3477_n605), .CO(
        DP_OP_422J2_124_3477_n572), .S(DP_OP_422J2_124_3477_n573) );
  FADDX1_HVT DP_OP_422J2_124_3477_U467 ( .A(DP_OP_422J2_124_3477_n738), .B(
        DP_OP_422J2_124_3477_n742), .CI(DP_OP_422J2_124_3477_n736), .CO(
        DP_OP_422J2_124_3477_n570), .S(DP_OP_422J2_124_3477_n571) );
  FADDX1_HVT DP_OP_422J2_124_3477_U466 ( .A(DP_OP_422J2_124_3477_n740), .B(
        DP_OP_422J2_124_3477_n732), .CI(DP_OP_422J2_124_3477_n730), .CO(
        DP_OP_422J2_124_3477_n568), .S(DP_OP_422J2_124_3477_n569) );
  FADDX1_HVT DP_OP_422J2_124_3477_U465 ( .A(DP_OP_422J2_124_3477_n599), .B(
        DP_OP_422J2_124_3477_n601), .CI(DP_OP_422J2_124_3477_n597), .CO(
        DP_OP_422J2_124_3477_n566), .S(DP_OP_422J2_124_3477_n567) );
  FADDX1_HVT DP_OP_422J2_124_3477_U464 ( .A(DP_OP_422J2_124_3477_n595), .B(
        DP_OP_422J2_124_3477_n589), .CI(DP_OP_422J2_124_3477_n593), .CO(
        DP_OP_422J2_124_3477_n564), .S(DP_OP_422J2_124_3477_n565) );
  FADDX1_HVT DP_OP_422J2_124_3477_U463 ( .A(DP_OP_422J2_124_3477_n587), .B(
        DP_OP_422J2_124_3477_n591), .CI(DP_OP_422J2_124_3477_n728), .CO(
        DP_OP_422J2_124_3477_n562), .S(DP_OP_422J2_124_3477_n563) );
  FADDX1_HVT DP_OP_422J2_124_3477_U462 ( .A(DP_OP_422J2_124_3477_n726), .B(
        DP_OP_422J2_124_3477_n722), .CI(DP_OP_422J2_124_3477_n585), .CO(
        DP_OP_422J2_124_3477_n560), .S(DP_OP_422J2_124_3477_n561) );
  FADDX1_HVT DP_OP_422J2_124_3477_U461 ( .A(DP_OP_422J2_124_3477_n724), .B(
        DP_OP_422J2_124_3477_n720), .CI(DP_OP_422J2_124_3477_n718), .CO(
        DP_OP_422J2_124_3477_n558), .S(DP_OP_422J2_124_3477_n559) );
  FADDX1_HVT DP_OP_422J2_124_3477_U460 ( .A(DP_OP_422J2_124_3477_n716), .B(
        DP_OP_422J2_124_3477_n583), .CI(DP_OP_422J2_124_3477_n581), .CO(
        DP_OP_422J2_124_3477_n556), .S(DP_OP_422J2_124_3477_n557) );
  FADDX1_HVT DP_OP_422J2_124_3477_U459 ( .A(DP_OP_422J2_124_3477_n714), .B(
        DP_OP_422J2_124_3477_n712), .CI(DP_OP_422J2_124_3477_n710), .CO(
        DP_OP_422J2_124_3477_n554), .S(DP_OP_422J2_124_3477_n555) );
  FADDX1_HVT DP_OP_422J2_124_3477_U458 ( .A(DP_OP_422J2_124_3477_n708), .B(
        DP_OP_422J2_124_3477_n579), .CI(DP_OP_422J2_124_3477_n706), .CO(
        DP_OP_422J2_124_3477_n552), .S(DP_OP_422J2_124_3477_n553) );
  FADDX1_HVT DP_OP_422J2_124_3477_U457 ( .A(DP_OP_422J2_124_3477_n577), .B(
        DP_OP_422J2_124_3477_n575), .CI(DP_OP_422J2_124_3477_n704), .CO(
        DP_OP_422J2_124_3477_n550), .S(DP_OP_422J2_124_3477_n551) );
  FADDX1_HVT DP_OP_422J2_124_3477_U456 ( .A(DP_OP_422J2_124_3477_n702), .B(
        DP_OP_422J2_124_3477_n571), .CI(DP_OP_422J2_124_3477_n569), .CO(
        DP_OP_422J2_124_3477_n548), .S(DP_OP_422J2_124_3477_n549) );
  FADDX1_HVT DP_OP_422J2_124_3477_U455 ( .A(DP_OP_422J2_124_3477_n573), .B(
        DP_OP_422J2_124_3477_n567), .CI(DP_OP_422J2_124_3477_n700), .CO(
        DP_OP_422J2_124_3477_n546), .S(DP_OP_422J2_124_3477_n547) );
  FADDX1_HVT DP_OP_422J2_124_3477_U454 ( .A(DP_OP_422J2_124_3477_n565), .B(
        DP_OP_422J2_124_3477_n698), .CI(DP_OP_422J2_124_3477_n563), .CO(
        DP_OP_422J2_124_3477_n544), .S(DP_OP_422J2_124_3477_n545) );
  FADDX1_HVT DP_OP_422J2_124_3477_U453 ( .A(DP_OP_422J2_124_3477_n696), .B(
        DP_OP_422J2_124_3477_n694), .CI(DP_OP_422J2_124_3477_n692), .CO(
        DP_OP_422J2_124_3477_n542), .S(DP_OP_422J2_124_3477_n543) );
  FADDX1_HVT DP_OP_422J2_124_3477_U452 ( .A(DP_OP_422J2_124_3477_n561), .B(
        DP_OP_422J2_124_3477_n690), .CI(DP_OP_422J2_124_3477_n559), .CO(
        DP_OP_422J2_124_3477_n540), .S(DP_OP_422J2_124_3477_n541) );
  FADDX1_HVT DP_OP_422J2_124_3477_U451 ( .A(DP_OP_422J2_124_3477_n688), .B(
        DP_OP_422J2_124_3477_n557), .CI(DP_OP_422J2_124_3477_n555), .CO(
        DP_OP_422J2_124_3477_n538), .S(DP_OP_422J2_124_3477_n539) );
  FADDX1_HVT DP_OP_422J2_124_3477_U450 ( .A(DP_OP_422J2_124_3477_n686), .B(
        DP_OP_422J2_124_3477_n684), .CI(DP_OP_422J2_124_3477_n553), .CO(
        DP_OP_422J2_124_3477_n536), .S(DP_OP_422J2_124_3477_n537) );
  FADDX1_HVT DP_OP_422J2_124_3477_U449 ( .A(DP_OP_422J2_124_3477_n682), .B(
        DP_OP_422J2_124_3477_n551), .CI(DP_OP_422J2_124_3477_n549), .CO(
        DP_OP_422J2_124_3477_n534), .S(DP_OP_422J2_124_3477_n535) );
  FADDX1_HVT DP_OP_422J2_124_3477_U447 ( .A(DP_OP_422J2_124_3477_n545), .B(
        DP_OP_422J2_124_3477_n676), .CI(DP_OP_422J2_124_3477_n543), .CO(
        DP_OP_422J2_124_3477_n530), .S(DP_OP_422J2_124_3477_n531) );
  FADDX1_HVT DP_OP_422J2_124_3477_U446 ( .A(DP_OP_422J2_124_3477_n674), .B(
        DP_OP_422J2_124_3477_n672), .CI(DP_OP_422J2_124_3477_n541), .CO(
        DP_OP_422J2_124_3477_n528), .S(DP_OP_422J2_124_3477_n529) );
  FADDX1_HVT DP_OP_422J2_124_3477_U445 ( .A(DP_OP_422J2_124_3477_n670), .B(
        DP_OP_422J2_124_3477_n539), .CI(DP_OP_422J2_124_3477_n537), .CO(
        DP_OP_422J2_124_3477_n526), .S(DP_OP_422J2_124_3477_n527) );
  FADDX1_HVT DP_OP_422J2_124_3477_U444 ( .A(DP_OP_422J2_124_3477_n668), .B(
        DP_OP_422J2_124_3477_n535), .CI(DP_OP_422J2_124_3477_n666), .CO(
        DP_OP_422J2_124_3477_n524), .S(DP_OP_422J2_124_3477_n525) );
  FADDX1_HVT DP_OP_422J2_124_3477_U443 ( .A(DP_OP_422J2_124_3477_n533), .B(
        DP_OP_422J2_124_3477_n664), .CI(DP_OP_422J2_124_3477_n531), .CO(
        DP_OP_422J2_124_3477_n522), .S(DP_OP_422J2_124_3477_n523) );
  FADDX1_HVT DP_OP_422J2_124_3477_U442 ( .A(DP_OP_422J2_124_3477_n662), .B(
        DP_OP_422J2_124_3477_n529), .CI(DP_OP_422J2_124_3477_n660), .CO(
        DP_OP_422J2_124_3477_n520), .S(DP_OP_422J2_124_3477_n521) );
  FADDX1_HVT DP_OP_422J2_124_3477_U441 ( .A(DP_OP_422J2_124_3477_n527), .B(
        DP_OP_422J2_124_3477_n525), .CI(DP_OP_422J2_124_3477_n658), .CO(
        DP_OP_422J2_124_3477_n518), .S(DP_OP_422J2_124_3477_n519) );
  FADDX1_HVT DP_OP_422J2_124_3477_U439 ( .A(DP_OP_422J2_124_3477_n521), .B(
        DP_OP_422J2_124_3477_n519), .CI(DP_OP_422J2_124_3477_n652), .CO(
        DP_OP_422J2_124_3477_n514), .S(DP_OP_422J2_124_3477_n515) );
  FADDX1_HVT DP_OP_422J2_124_3477_U436 ( .A(DP_OP_422J2_124_3477_n3026), .B(
        DP_OP_422J2_124_3477_n1970), .CI(DP_OP_422J2_124_3477_n511), .CO(
        DP_OP_422J2_124_3477_n508), .S(DP_OP_422J2_124_3477_n509) );
  FADDX1_HVT DP_OP_422J2_124_3477_U435 ( .A(DP_OP_422J2_124_3477_n2058), .B(
        DP_OP_422J2_124_3477_n2982), .CI(DP_OP_422J2_124_3477_n2410), .CO(
        DP_OP_422J2_124_3477_n506), .S(DP_OP_422J2_124_3477_n507) );
  FADDX1_HVT DP_OP_422J2_124_3477_U434 ( .A(DP_OP_422J2_124_3477_n2542), .B(
        DP_OP_422J2_124_3477_n2938), .CI(DP_OP_422J2_124_3477_n2894), .CO(
        DP_OP_422J2_124_3477_n504), .S(DP_OP_422J2_124_3477_n505) );
  FADDX1_HVT DP_OP_422J2_124_3477_U433 ( .A(DP_OP_422J2_124_3477_n2366), .B(
        DP_OP_422J2_124_3477_n2850), .CI(DP_OP_422J2_124_3477_n2806), .CO(
        DP_OP_422J2_124_3477_n502), .S(DP_OP_422J2_124_3477_n503) );
  FADDX1_HVT DP_OP_422J2_124_3477_U432 ( .A(DP_OP_422J2_124_3477_n2234), .B(
        DP_OP_422J2_124_3477_n2014), .CI(DP_OP_422J2_124_3477_n2762), .CO(
        DP_OP_422J2_124_3477_n500), .S(DP_OP_422J2_124_3477_n501) );
  FADDX1_HVT DP_OP_422J2_124_3477_U431 ( .A(DP_OP_422J2_124_3477_n2718), .B(
        DP_OP_422J2_124_3477_n2674), .CI(DP_OP_422J2_124_3477_n2630), .CO(
        DP_OP_422J2_124_3477_n498), .S(DP_OP_422J2_124_3477_n499) );
  FADDX1_HVT DP_OP_422J2_124_3477_U430 ( .A(DP_OP_422J2_124_3477_n2278), .B(
        DP_OP_422J2_124_3477_n2102), .CI(DP_OP_422J2_124_3477_n2146), .CO(
        DP_OP_422J2_124_3477_n496), .S(DP_OP_422J2_124_3477_n497) );
  FADDX1_HVT DP_OP_422J2_124_3477_U429 ( .A(DP_OP_422J2_124_3477_n2190), .B(
        DP_OP_422J2_124_3477_n2586), .CI(DP_OP_422J2_124_3477_n2498), .CO(
        DP_OP_422J2_124_3477_n494), .S(DP_OP_422J2_124_3477_n495) );
  FADDX1_HVT DP_OP_422J2_124_3477_U428 ( .A(DP_OP_422J2_124_3477_n2322), .B(
        DP_OP_422J2_124_3477_n2454), .CI(DP_OP_422J2_124_3477_n646), .CO(
        DP_OP_422J2_124_3477_n492), .S(DP_OP_422J2_124_3477_n493) );
  FADDX1_HVT DP_OP_422J2_124_3477_U427 ( .A(DP_OP_422J2_124_3477_n644), .B(
        DP_OP_422J2_124_3477_n614), .CI(DP_OP_422J2_124_3477_n642), .CO(
        DP_OP_422J2_124_3477_n490), .S(DP_OP_422J2_124_3477_n491) );
  FADDX1_HVT DP_OP_422J2_124_3477_U426 ( .A(DP_OP_422J2_124_3477_n640), .B(
        DP_OP_422J2_124_3477_n616), .CI(DP_OP_422J2_124_3477_n618), .CO(
        DP_OP_422J2_124_3477_n488), .S(DP_OP_422J2_124_3477_n489) );
  FADDX1_HVT DP_OP_422J2_124_3477_U425 ( .A(DP_OP_422J2_124_3477_n638), .B(
        DP_OP_422J2_124_3477_n620), .CI(DP_OP_422J2_124_3477_n622), .CO(
        DP_OP_422J2_124_3477_n486), .S(DP_OP_422J2_124_3477_n487) );
  FADDX1_HVT DP_OP_422J2_124_3477_U424 ( .A(DP_OP_422J2_124_3477_n636), .B(
        DP_OP_422J2_124_3477_n624), .CI(DP_OP_422J2_124_3477_n626), .CO(
        DP_OP_422J2_124_3477_n484), .S(DP_OP_422J2_124_3477_n485) );
  FADDX1_HVT DP_OP_422J2_124_3477_U423 ( .A(DP_OP_422J2_124_3477_n634), .B(
        DP_OP_422J2_124_3477_n628), .CI(DP_OP_422J2_124_3477_n630), .CO(
        DP_OP_422J2_124_3477_n482), .S(DP_OP_422J2_124_3477_n483) );
  FADDX1_HVT DP_OP_422J2_124_3477_U422 ( .A(DP_OP_422J2_124_3477_n632), .B(
        DP_OP_422J2_124_3477_n509), .CI(DP_OP_422J2_124_3477_n505), .CO(
        DP_OP_422J2_124_3477_n480), .S(DP_OP_422J2_124_3477_n481) );
  FADDX1_HVT DP_OP_422J2_124_3477_U421 ( .A(DP_OP_422J2_124_3477_n501), .B(
        DP_OP_422J2_124_3477_n495), .CI(DP_OP_422J2_124_3477_n497), .CO(
        DP_OP_422J2_124_3477_n478), .S(DP_OP_422J2_124_3477_n479) );
  FADDX1_HVT DP_OP_422J2_124_3477_U420 ( .A(DP_OP_422J2_124_3477_n499), .B(
        DP_OP_422J2_124_3477_n507), .CI(DP_OP_422J2_124_3477_n503), .CO(
        DP_OP_422J2_124_3477_n476), .S(DP_OP_422J2_124_3477_n477) );
  FADDX1_HVT DP_OP_422J2_124_3477_U419 ( .A(DP_OP_422J2_124_3477_n612), .B(
        DP_OP_422J2_124_3477_n610), .CI(DP_OP_422J2_124_3477_n602), .CO(
        DP_OP_422J2_124_3477_n474), .S(DP_OP_422J2_124_3477_n475) );
  FADDX1_HVT DP_OP_422J2_124_3477_U418 ( .A(DP_OP_422J2_124_3477_n608), .B(
        DP_OP_422J2_124_3477_n604), .CI(DP_OP_422J2_124_3477_n606), .CO(
        DP_OP_422J2_124_3477_n472), .S(DP_OP_422J2_124_3477_n473) );
  FADDX1_HVT DP_OP_422J2_124_3477_U417 ( .A(DP_OP_422J2_124_3477_n600), .B(
        DP_OP_422J2_124_3477_n596), .CI(DP_OP_422J2_124_3477_n493), .CO(
        DP_OP_422J2_124_3477_n470), .S(DP_OP_422J2_124_3477_n471) );
  FADDX1_HVT DP_OP_422J2_124_3477_U416 ( .A(DP_OP_422J2_124_3477_n598), .B(
        DP_OP_422J2_124_3477_n594), .CI(DP_OP_422J2_124_3477_n491), .CO(
        DP_OP_422J2_124_3477_n468), .S(DP_OP_422J2_124_3477_n469) );
  FADDX1_HVT DP_OP_422J2_124_3477_U415 ( .A(DP_OP_422J2_124_3477_n592), .B(
        DP_OP_422J2_124_3477_n485), .CI(DP_OP_422J2_124_3477_n487), .CO(
        DP_OP_422J2_124_3477_n466), .S(DP_OP_422J2_124_3477_n467) );
  FADDX1_HVT DP_OP_422J2_124_3477_U414 ( .A(DP_OP_422J2_124_3477_n590), .B(
        DP_OP_422J2_124_3477_n489), .CI(DP_OP_422J2_124_3477_n483), .CO(
        DP_OP_422J2_124_3477_n464), .S(DP_OP_422J2_124_3477_n465) );
  FADDX1_HVT DP_OP_422J2_124_3477_U413 ( .A(DP_OP_422J2_124_3477_n588), .B(
        DP_OP_422J2_124_3477_n586), .CI(DP_OP_422J2_124_3477_n584), .CO(
        DP_OP_422J2_124_3477_n462), .S(DP_OP_422J2_124_3477_n463) );
  FADDX1_HVT DP_OP_422J2_124_3477_U412 ( .A(DP_OP_422J2_124_3477_n481), .B(
        DP_OP_422J2_124_3477_n477), .CI(DP_OP_422J2_124_3477_n582), .CO(
        DP_OP_422J2_124_3477_n460), .S(DP_OP_422J2_124_3477_n461) );
  FADDX1_HVT DP_OP_422J2_124_3477_U411 ( .A(DP_OP_422J2_124_3477_n479), .B(
        DP_OP_422J2_124_3477_n580), .CI(DP_OP_422J2_124_3477_n578), .CO(
        DP_OP_422J2_124_3477_n458), .S(DP_OP_422J2_124_3477_n459) );
  FADDX1_HVT DP_OP_422J2_124_3477_U410 ( .A(DP_OP_422J2_124_3477_n576), .B(
        DP_OP_422J2_124_3477_n475), .CI(DP_OP_422J2_124_3477_n473), .CO(
        DP_OP_422J2_124_3477_n456), .S(DP_OP_422J2_124_3477_n457) );
  FADDX1_HVT DP_OP_422J2_124_3477_U409 ( .A(DP_OP_422J2_124_3477_n574), .B(
        DP_OP_422J2_124_3477_n570), .CI(DP_OP_422J2_124_3477_n568), .CO(
        DP_OP_422J2_124_3477_n454), .S(DP_OP_422J2_124_3477_n455) );
  FADDX1_HVT DP_OP_422J2_124_3477_U408 ( .A(DP_OP_422J2_124_3477_n572), .B(
        DP_OP_422J2_124_3477_n566), .CI(DP_OP_422J2_124_3477_n471), .CO(
        DP_OP_422J2_124_3477_n452), .S(DP_OP_422J2_124_3477_n453) );
  FADDX1_HVT DP_OP_422J2_124_3477_U407 ( .A(DP_OP_422J2_124_3477_n469), .B(
        DP_OP_422J2_124_3477_n564), .CI(DP_OP_422J2_124_3477_n562), .CO(
        DP_OP_422J2_124_3477_n450), .S(DP_OP_422J2_124_3477_n451) );
  FADDX1_HVT DP_OP_422J2_124_3477_U406 ( .A(DP_OP_422J2_124_3477_n467), .B(
        DP_OP_422J2_124_3477_n465), .CI(DP_OP_422J2_124_3477_n463), .CO(
        DP_OP_422J2_124_3477_n448), .S(DP_OP_422J2_124_3477_n449) );
  FADDX1_HVT DP_OP_422J2_124_3477_U405 ( .A(DP_OP_422J2_124_3477_n558), .B(
        DP_OP_422J2_124_3477_n560), .CI(DP_OP_422J2_124_3477_n461), .CO(
        DP_OP_422J2_124_3477_n446), .S(DP_OP_422J2_124_3477_n447) );
  FADDX1_HVT DP_OP_422J2_124_3477_U404 ( .A(DP_OP_422J2_124_3477_n556), .B(
        DP_OP_422J2_124_3477_n459), .CI(DP_OP_422J2_124_3477_n554), .CO(
        DP_OP_422J2_124_3477_n444), .S(DP_OP_422J2_124_3477_n445) );
  FADDX1_HVT DP_OP_422J2_124_3477_U403 ( .A(DP_OP_422J2_124_3477_n552), .B(
        DP_OP_422J2_124_3477_n457), .CI(DP_OP_422J2_124_3477_n550), .CO(
        DP_OP_422J2_124_3477_n442), .S(DP_OP_422J2_124_3477_n443) );
  FADDX1_HVT DP_OP_422J2_124_3477_U402 ( .A(DP_OP_422J2_124_3477_n548), .B(
        DP_OP_422J2_124_3477_n455), .CI(DP_OP_422J2_124_3477_n453), .CO(
        DP_OP_422J2_124_3477_n440), .S(DP_OP_422J2_124_3477_n441) );
  FADDX1_HVT DP_OP_422J2_124_3477_U401 ( .A(DP_OP_422J2_124_3477_n546), .B(
        DP_OP_422J2_124_3477_n451), .CI(DP_OP_422J2_124_3477_n544), .CO(
        DP_OP_422J2_124_3477_n438), .S(DP_OP_422J2_124_3477_n439) );
  FADDX1_HVT DP_OP_422J2_124_3477_U400 ( .A(DP_OP_422J2_124_3477_n449), .B(
        DP_OP_422J2_124_3477_n542), .CI(DP_OP_422J2_124_3477_n540), .CO(
        DP_OP_422J2_124_3477_n436), .S(DP_OP_422J2_124_3477_n437) );
  FADDX1_HVT DP_OP_422J2_124_3477_U399 ( .A(DP_OP_422J2_124_3477_n447), .B(
        DP_OP_422J2_124_3477_n538), .CI(DP_OP_422J2_124_3477_n445), .CO(
        DP_OP_422J2_124_3477_n434), .S(DP_OP_422J2_124_3477_n435) );
  FADDX1_HVT DP_OP_422J2_124_3477_U398 ( .A(DP_OP_422J2_124_3477_n536), .B(
        DP_OP_422J2_124_3477_n443), .CI(DP_OP_422J2_124_3477_n534), .CO(
        DP_OP_422J2_124_3477_n432), .S(DP_OP_422J2_124_3477_n433) );
  FADDX1_HVT DP_OP_422J2_124_3477_U397 ( .A(DP_OP_422J2_124_3477_n441), .B(
        DP_OP_422J2_124_3477_n532), .CI(DP_OP_422J2_124_3477_n439), .CO(
        DP_OP_422J2_124_3477_n430), .S(DP_OP_422J2_124_3477_n431) );
  FADDX1_HVT DP_OP_422J2_124_3477_U396 ( .A(DP_OP_422J2_124_3477_n530), .B(
        DP_OP_422J2_124_3477_n437), .CI(DP_OP_422J2_124_3477_n528), .CO(
        DP_OP_422J2_124_3477_n428), .S(DP_OP_422J2_124_3477_n429) );
  FADDX1_HVT DP_OP_422J2_124_3477_U395 ( .A(DP_OP_422J2_124_3477_n435), .B(
        DP_OP_422J2_124_3477_n526), .CI(DP_OP_422J2_124_3477_n433), .CO(
        DP_OP_422J2_124_3477_n426), .S(DP_OP_422J2_124_3477_n427) );
  FADDX1_HVT DP_OP_422J2_124_3477_U394 ( .A(DP_OP_422J2_124_3477_n524), .B(
        DP_OP_422J2_124_3477_n431), .CI(DP_OP_422J2_124_3477_n522), .CO(
        DP_OP_422J2_124_3477_n424), .S(DP_OP_422J2_124_3477_n425) );
  FADDX1_HVT DP_OP_422J2_124_3477_U393 ( .A(DP_OP_422J2_124_3477_n429), .B(
        DP_OP_422J2_124_3477_n520), .CI(DP_OP_422J2_124_3477_n427), .CO(
        DP_OP_422J2_124_3477_n422), .S(DP_OP_422J2_124_3477_n423) );
  FADDX1_HVT DP_OP_422J2_124_3477_U391 ( .A(DP_OP_422J2_124_3477_n423), .B(
        DP_OP_422J2_124_3477_n514), .CI(DP_OP_422J2_124_3477_n421), .CO(
        DP_OP_422J2_124_3477_n418), .S(DP_OP_422J2_124_3477_n419) );
  FADDX1_HVT DP_OP_422J2_124_3477_U390 ( .A(DP_OP_422J2_124_3477_n1926), .B(
        DP_OP_422J2_124_3477_n510), .CI(DP_OP_422J2_124_3477_n508), .CO(
        DP_OP_422J2_124_3477_n416), .S(DP_OP_422J2_124_3477_n417) );
  FADDX1_HVT DP_OP_422J2_124_3477_U389 ( .A(DP_OP_422J2_124_3477_n498), .B(
        DP_OP_422J2_124_3477_n494), .CI(DP_OP_422J2_124_3477_n506), .CO(
        DP_OP_422J2_124_3477_n414), .S(DP_OP_422J2_124_3477_n415) );
  FADDX1_HVT DP_OP_422J2_124_3477_U388 ( .A(DP_OP_422J2_124_3477_n504), .B(
        DP_OP_422J2_124_3477_n502), .CI(DP_OP_422J2_124_3477_n500), .CO(
        DP_OP_422J2_124_3477_n412), .S(DP_OP_422J2_124_3477_n413) );
  FADDX1_HVT DP_OP_422J2_124_3477_U387 ( .A(DP_OP_422J2_124_3477_n496), .B(
        DP_OP_422J2_124_3477_n492), .CI(DP_OP_422J2_124_3477_n490), .CO(
        DP_OP_422J2_124_3477_n410), .S(DP_OP_422J2_124_3477_n411) );
  FADDX1_HVT DP_OP_422J2_124_3477_U386 ( .A(DP_OP_422J2_124_3477_n488), .B(
        DP_OP_422J2_124_3477_n486), .CI(DP_OP_422J2_124_3477_n484), .CO(
        DP_OP_422J2_124_3477_n408), .S(DP_OP_422J2_124_3477_n409) );
  FADDX1_HVT DP_OP_422J2_124_3477_U385 ( .A(DP_OP_422J2_124_3477_n482), .B(
        DP_OP_422J2_124_3477_n417), .CI(DP_OP_422J2_124_3477_n480), .CO(
        DP_OP_422J2_124_3477_n406), .S(DP_OP_422J2_124_3477_n407) );
  FADDX1_HVT DP_OP_422J2_124_3477_U384 ( .A(DP_OP_422J2_124_3477_n478), .B(
        DP_OP_422J2_124_3477_n413), .CI(DP_OP_422J2_124_3477_n415), .CO(
        DP_OP_422J2_124_3477_n404), .S(DP_OP_422J2_124_3477_n405) );
  FADDX1_HVT DP_OP_422J2_124_3477_U383 ( .A(DP_OP_422J2_124_3477_n476), .B(
        DP_OP_422J2_124_3477_n474), .CI(DP_OP_422J2_124_3477_n472), .CO(
        DP_OP_422J2_124_3477_n402), .S(DP_OP_422J2_124_3477_n403) );
  FADDX1_HVT DP_OP_422J2_124_3477_U382 ( .A(DP_OP_422J2_124_3477_n470), .B(
        DP_OP_422J2_124_3477_n411), .CI(DP_OP_422J2_124_3477_n468), .CO(
        DP_OP_422J2_124_3477_n400), .S(DP_OP_422J2_124_3477_n401) );
  FADDX1_HVT DP_OP_422J2_124_3477_U381 ( .A(DP_OP_422J2_124_3477_n466), .B(
        DP_OP_422J2_124_3477_n409), .CI(DP_OP_422J2_124_3477_n464), .CO(
        DP_OP_422J2_124_3477_n398), .S(DP_OP_422J2_124_3477_n399) );
  FADDX1_HVT DP_OP_422J2_124_3477_U380 ( .A(DP_OP_422J2_124_3477_n462), .B(
        DP_OP_422J2_124_3477_n407), .CI(DP_OP_422J2_124_3477_n460), .CO(
        DP_OP_422J2_124_3477_n396), .S(DP_OP_422J2_124_3477_n397) );
  FADDX1_HVT DP_OP_422J2_124_3477_U379 ( .A(DP_OP_422J2_124_3477_n405), .B(
        DP_OP_422J2_124_3477_n458), .CI(DP_OP_422J2_124_3477_n456), .CO(
        DP_OP_422J2_124_3477_n394), .S(DP_OP_422J2_124_3477_n395) );
  FADDX1_HVT DP_OP_422J2_124_3477_U378 ( .A(DP_OP_422J2_124_3477_n403), .B(
        DP_OP_422J2_124_3477_n454), .CI(DP_OP_422J2_124_3477_n452), .CO(
        DP_OP_422J2_124_3477_n392), .S(DP_OP_422J2_124_3477_n393) );
  FADDX1_HVT DP_OP_422J2_124_3477_U377 ( .A(DP_OP_422J2_124_3477_n401), .B(
        DP_OP_422J2_124_3477_n450), .CI(DP_OP_422J2_124_3477_n399), .CO(
        DP_OP_422J2_124_3477_n390), .S(DP_OP_422J2_124_3477_n391) );
  FADDX1_HVT DP_OP_422J2_124_3477_U376 ( .A(DP_OP_422J2_124_3477_n448), .B(
        DP_OP_422J2_124_3477_n397), .CI(DP_OP_422J2_124_3477_n446), .CO(
        DP_OP_422J2_124_3477_n388), .S(DP_OP_422J2_124_3477_n389) );
  FADDX1_HVT DP_OP_422J2_124_3477_U375 ( .A(DP_OP_422J2_124_3477_n444), .B(
        DP_OP_422J2_124_3477_n395), .CI(DP_OP_422J2_124_3477_n442), .CO(
        DP_OP_422J2_124_3477_n386), .S(DP_OP_422J2_124_3477_n387) );
  FADDX1_HVT DP_OP_422J2_124_3477_U374 ( .A(DP_OP_422J2_124_3477_n393), .B(
        DP_OP_422J2_124_3477_n440), .CI(DP_OP_422J2_124_3477_n438), .CO(
        DP_OP_422J2_124_3477_n384), .S(DP_OP_422J2_124_3477_n385) );
  FADDX1_HVT DP_OP_422J2_124_3477_U373 ( .A(DP_OP_422J2_124_3477_n391), .B(
        DP_OP_422J2_124_3477_n436), .CI(DP_OP_422J2_124_3477_n389), .CO(
        DP_OP_422J2_124_3477_n382), .S(DP_OP_422J2_124_3477_n383) );
  FADDX1_HVT DP_OP_422J2_124_3477_U372 ( .A(DP_OP_422J2_124_3477_n434), .B(
        DP_OP_422J2_124_3477_n387), .CI(DP_OP_422J2_124_3477_n432), .CO(
        DP_OP_422J2_124_3477_n380), .S(DP_OP_422J2_124_3477_n381) );
  FADDX1_HVT DP_OP_422J2_124_3477_U371 ( .A(DP_OP_422J2_124_3477_n430), .B(
        DP_OP_422J2_124_3477_n385), .CI(DP_OP_422J2_124_3477_n383), .CO(
        DP_OP_422J2_124_3477_n378), .S(DP_OP_422J2_124_3477_n379) );
  FADDX1_HVT DP_OP_422J2_124_3477_U370 ( .A(DP_OP_422J2_124_3477_n428), .B(
        DP_OP_422J2_124_3477_n381), .CI(DP_OP_422J2_124_3477_n426), .CO(
        DP_OP_422J2_124_3477_n376), .S(DP_OP_422J2_124_3477_n377) );
  FADDX1_HVT DP_OP_422J2_124_3477_U367 ( .A(DP_OP_422J2_124_3477_n1925), .B(
        DP_OP_422J2_124_3477_n416), .CI(DP_OP_422J2_124_3477_n414), .CO(
        DP_OP_422J2_124_3477_n370), .S(DP_OP_422J2_124_3477_n371) );
  FADDX1_HVT DP_OP_422J2_124_3477_U366 ( .A(DP_OP_422J2_124_3477_n412), .B(
        DP_OP_422J2_124_3477_n410), .CI(DP_OP_422J2_124_3477_n408), .CO(
        DP_OP_422J2_124_3477_n368), .S(DP_OP_422J2_124_3477_n369) );
  FADDX1_HVT DP_OP_422J2_124_3477_U365 ( .A(DP_OP_422J2_124_3477_n406), .B(
        DP_OP_422J2_124_3477_n371), .CI(DP_OP_422J2_124_3477_n404), .CO(
        DP_OP_422J2_124_3477_n366), .S(DP_OP_422J2_124_3477_n367) );
  FADDX1_HVT DP_OP_422J2_124_3477_U364 ( .A(DP_OP_422J2_124_3477_n402), .B(
        DP_OP_422J2_124_3477_n400), .CI(DP_OP_422J2_124_3477_n369), .CO(
        DP_OP_422J2_124_3477_n364), .S(DP_OP_422J2_124_3477_n365) );
  FADDX1_HVT DP_OP_422J2_124_3477_U363 ( .A(DP_OP_422J2_124_3477_n398), .B(
        DP_OP_422J2_124_3477_n396), .CI(DP_OP_422J2_124_3477_n367), .CO(
        DP_OP_422J2_124_3477_n362), .S(DP_OP_422J2_124_3477_n363) );
  FADDX1_HVT DP_OP_422J2_124_3477_U362 ( .A(DP_OP_422J2_124_3477_n394), .B(
        DP_OP_422J2_124_3477_n392), .CI(DP_OP_422J2_124_3477_n365), .CO(
        DP_OP_422J2_124_3477_n360), .S(DP_OP_422J2_124_3477_n361) );
  FADDX1_HVT DP_OP_422J2_124_3477_U361 ( .A(DP_OP_422J2_124_3477_n390), .B(
        DP_OP_422J2_124_3477_n363), .CI(DP_OP_422J2_124_3477_n388), .CO(
        DP_OP_422J2_124_3477_n358), .S(DP_OP_422J2_124_3477_n359) );
  FADDX1_HVT DP_OP_422J2_124_3477_U360 ( .A(DP_OP_422J2_124_3477_n386), .B(
        DP_OP_422J2_124_3477_n361), .CI(DP_OP_422J2_124_3477_n384), .CO(
        DP_OP_422J2_124_3477_n356), .S(DP_OP_422J2_124_3477_n357) );
  FADDX1_HVT DP_OP_422J2_124_3477_U358 ( .A(DP_OP_422J2_124_3477_n357), .B(
        DP_OP_422J2_124_3477_n378), .CI(DP_OP_422J2_124_3477_n355), .CO(
        DP_OP_422J2_124_3477_n352), .S(DP_OP_422J2_124_3477_n353) );
  FADDX1_HVT DP_OP_422J2_124_3477_U357 ( .A(DP_OP_422J2_124_3477_n376), .B(
        DP_OP_422J2_124_3477_n374), .CI(DP_OP_422J2_124_3477_n353), .CO(
        DP_OP_422J2_124_3477_n350), .S(DP_OP_422J2_124_3477_n351) );
  FADDX1_HVT DP_OP_422J2_124_3477_U356 ( .A(DP_OP_422J2_124_3477_n1924), .B(
        DP_OP_422J2_124_3477_n370), .CI(DP_OP_422J2_124_3477_n368), .CO(
        DP_OP_422J2_124_3477_n348), .S(DP_OP_422J2_124_3477_n349) );
  FADDX1_HVT DP_OP_422J2_124_3477_U355 ( .A(DP_OP_422J2_124_3477_n366), .B(
        DP_OP_422J2_124_3477_n349), .CI(DP_OP_422J2_124_3477_n364), .CO(
        DP_OP_422J2_124_3477_n346), .S(DP_OP_422J2_124_3477_n347) );
  FADDX1_HVT DP_OP_422J2_124_3477_U354 ( .A(DP_OP_422J2_124_3477_n362), .B(
        DP_OP_422J2_124_3477_n360), .CI(DP_OP_422J2_124_3477_n347), .CO(
        DP_OP_422J2_124_3477_n344), .S(DP_OP_422J2_124_3477_n345) );
  FADDX1_HVT DP_OP_422J2_124_3477_U353 ( .A(DP_OP_422J2_124_3477_n358), .B(
        DP_OP_422J2_124_3477_n345), .CI(DP_OP_422J2_124_3477_n356), .CO(
        DP_OP_422J2_124_3477_n342), .S(DP_OP_422J2_124_3477_n343) );
  FADDX1_HVT DP_OP_422J2_124_3477_U352 ( .A(DP_OP_422J2_124_3477_n354), .B(
        DP_OP_422J2_124_3477_n343), .CI(DP_OP_422J2_124_3477_n352), .CO(
        DP_OP_422J2_124_3477_n340), .S(DP_OP_422J2_124_3477_n341) );
  FADDX1_HVT DP_OP_422J2_124_3477_U350 ( .A(DP_OP_422J2_124_3477_n339), .B(
        DP_OP_422J2_124_3477_n348), .CI(DP_OP_422J2_124_3477_n346), .CO(
        DP_OP_422J2_124_3477_n336), .S(DP_OP_422J2_124_3477_n337) );
  FADDX1_HVT DP_OP_422J2_124_3477_U349 ( .A(DP_OP_422J2_124_3477_n337), .B(
        DP_OP_422J2_124_3477_n344), .CI(DP_OP_422J2_124_3477_n342), .CO(
        DP_OP_422J2_124_3477_n334), .S(DP_OP_422J2_124_3477_n335) );
  FADDX1_HVT DP_OP_422J2_124_3477_U348 ( .A(DP_OP_422J2_124_3477_n1923), .B(
        DP_OP_422J2_124_3477_n338), .CI(DP_OP_422J2_124_3477_n336), .CO(
        DP_OP_422J2_124_3477_n332), .S(DP_OP_422J2_124_3477_n333) );
  FADDX1_HVT DP_OP_422J2_124_3477_U331 ( .A(DP_OP_422J2_124_3477_n1903), .B(
        DP_OP_422J2_124_3477_n1901), .CI(DP_OP_422J2_124_3477_n1899), .CO(
        DP_OP_422J2_124_3477_n269), .S(n_conv2_sum_a[0]) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U330 ( .A1(DP_OP_422J2_124_3477_n1837), 
        .A2(DP_OP_422J2_124_3477_n1839), .Y(DP_OP_422J2_124_3477_n268) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U329 ( .A1(DP_OP_422J2_124_3477_n1839), .A2(
        DP_OP_422J2_124_3477_n1837), .Y(DP_OP_422J2_124_3477_n267) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U323 ( .A1(DP_OP_422J2_124_3477_n1731), 
        .A2(DP_OP_422J2_124_3477_n1733), .Y(DP_OP_422J2_124_3477_n265) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U315 ( .A1(DP_OP_422J2_124_3477_n1577), 
        .A2(DP_OP_422J2_124_3477_n1579), .Y(DP_OP_422J2_124_3477_n260) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U314 ( .A1(DP_OP_422J2_124_3477_n1579), .A2(
        DP_OP_422J2_124_3477_n1577), .Y(DP_OP_422J2_124_3477_n259) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U309 ( .A1(DP_OP_422J2_124_3477_n1401), 
        .A2(DP_OP_422J2_124_3477_n1403), .Y(DP_OP_422J2_124_3477_n257) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U295 ( .A1(DP_OP_422J2_124_3477_n1019), 
        .A2(DP_OP_422J2_124_3477_n1021), .Y(DP_OP_422J2_124_3477_n249) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U294 ( .A1(DP_OP_422J2_124_3477_n1021), .A2(
        DP_OP_422J2_124_3477_n1019), .Y(DP_OP_422J2_124_3477_n248) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U287 ( .A1(DP_OP_422J2_124_3477_n823), .A2(
        DP_OP_422J2_124_3477_n1018), .Y(DP_OP_422J2_124_3477_n244) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U274 ( .A1(DP_OP_422J2_124_3477_n648), .A2(
        DP_OP_422J2_124_3477_n513), .Y(DP_OP_422J2_124_3477_n237) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U257 ( .A1(DP_OP_422J2_124_3477_n418), .A2(
        DP_OP_422J2_124_3477_n373), .Y(DP_OP_422J2_124_3477_n226) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U235 ( .A1(DP_OP_422J2_124_3477_n350), .A2(
        DP_OP_422J2_124_3477_n341), .Y(DP_OP_422J2_124_3477_n210) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U234 ( .A1(DP_OP_422J2_124_3477_n341), .A2(
        DP_OP_422J2_124_3477_n350), .Y(DP_OP_422J2_124_3477_n209) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U217 ( .A1(DP_OP_422J2_124_3477_n334), .A2(
        DP_OP_422J2_124_3477_n333), .Y(DP_OP_422J2_124_3477_n198) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U216 ( .A1(DP_OP_422J2_124_3477_n333), .A2(
        DP_OP_422J2_124_3477_n334), .Y(DP_OP_422J2_124_3477_n197) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U214 ( .A1(DP_OP_422J2_124_3477_n286), .A2(
        DP_OP_422J2_124_3477_n198), .Y(DP_OP_422J2_124_3477_n22) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U210 ( .A1(n1592), .A2(
        DP_OP_422J2_124_3477_n286), .Y(DP_OP_422J2_124_3477_n189) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U201 ( .A1(DP_OP_422J2_124_3477_n332), .A2(
        DP_OP_422J2_124_3477_n331), .Y(DP_OP_422J2_124_3477_n185) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U200 ( .A1(DP_OP_422J2_124_3477_n331), .A2(
        DP_OP_422J2_124_3477_n332), .Y(DP_OP_422J2_124_3477_n182) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U194 ( .A1(DP_OP_422J2_124_3477_n182), .A2(
        DP_OP_422J2_124_3477_n189), .Y(DP_OP_422J2_124_3477_n176) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U187 ( .A1(DP_OP_422J2_124_3477_n329), .A2(
        DP_OP_422J2_124_3477_n330), .Y(DP_OP_422J2_124_3477_n174) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U186 ( .A1(DP_OP_422J2_124_3477_n330), .A2(
        DP_OP_422J2_124_3477_n329), .Y(DP_OP_422J2_124_3477_n171) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U177 ( .A1(DP_OP_422J2_124_3477_n327), .A2(
        DP_OP_422J2_124_3477_n328), .Y(DP_OP_422J2_124_3477_n167) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U176 ( .A1(DP_OP_422J2_124_3477_n328), .A2(
        DP_OP_422J2_124_3477_n327), .Y(DP_OP_422J2_124_3477_n166) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U172 ( .A1(DP_OP_422J2_124_3477_n166), .A2(
        DP_OP_422J2_124_3477_n171), .Y(DP_OP_422J2_124_3477_n162) );
  AOI21X1_HVT DP_OP_422J2_124_3477_U169 ( .A1(DP_OP_422J2_124_3477_n177), .A2(
        DP_OP_422J2_124_3477_n162), .A3(DP_OP_422J2_124_3477_n165), .Y(
        DP_OP_422J2_124_3477_n161) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U168 ( .A1(DP_OP_422J2_124_3477_n176), .A2(
        DP_OP_422J2_124_3477_n162), .Y(DP_OP_422J2_124_3477_n160) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U163 ( .A1(DP_OP_422J2_124_3477_n325), .A2(
        DP_OP_422J2_124_3477_n326), .Y(DP_OP_422J2_124_3477_n156) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U162 ( .A1(DP_OP_422J2_124_3477_n326), .A2(
        DP_OP_422J2_124_3477_n325), .Y(DP_OP_422J2_124_3477_n153) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U153 ( .A1(DP_OP_422J2_124_3477_n323), .A2(
        DP_OP_422J2_124_3477_n324), .Y(DP_OP_422J2_124_3477_n149) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U152 ( .A1(DP_OP_422J2_124_3477_n324), .A2(
        DP_OP_422J2_124_3477_n323), .Y(DP_OP_422J2_124_3477_n148) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U148 ( .A1(DP_OP_422J2_124_3477_n148), .A2(
        DP_OP_422J2_124_3477_n153), .Y(DP_OP_422J2_124_3477_n146) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U146 ( .A1(DP_OP_422J2_124_3477_n162), .A2(
        DP_OP_422J2_124_3477_n146), .Y(DP_OP_422J2_124_3477_n144) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U142 ( .A1(DP_OP_422J2_124_3477_n176), .A2(
        DP_OP_422J2_124_3477_n142), .Y(DP_OP_422J2_124_3477_n140) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U137 ( .A1(DP_OP_422J2_124_3477_n321), .A2(
        DP_OP_422J2_124_3477_n322), .Y(DP_OP_422J2_124_3477_n136) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U136 ( .A1(DP_OP_422J2_124_3477_n322), .A2(
        DP_OP_422J2_124_3477_n321), .Y(DP_OP_422J2_124_3477_n133) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U127 ( .A1(DP_OP_422J2_124_3477_n319), .A2(
        DP_OP_422J2_124_3477_n320), .Y(DP_OP_422J2_124_3477_n129) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U126 ( .A1(DP_OP_422J2_124_3477_n320), .A2(
        DP_OP_422J2_124_3477_n319), .Y(DP_OP_422J2_124_3477_n128) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U122 ( .A1(DP_OP_422J2_124_3477_n128), .A2(
        DP_OP_422J2_124_3477_n133), .Y(DP_OP_422J2_124_3477_n126) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U115 ( .A1(DP_OP_422J2_124_3477_n317), .A2(
        DP_OP_422J2_124_3477_n318), .Y(DP_OP_422J2_124_3477_n120) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U108 ( .A1(DP_OP_422J2_124_3477_n126), .A2(
        n1588), .Y(DP_OP_422J2_124_3477_n115) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U106 ( .A1(DP_OP_422J2_124_3477_n115), .A2(
        DP_OP_422J2_124_3477_n144), .Y(DP_OP_422J2_124_3477_n111) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U102 ( .A1(DP_OP_422J2_124_3477_n176), .A2(
        DP_OP_422J2_124_3477_n111), .Y(DP_OP_422J2_124_3477_n109) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U97 ( .A1(DP_OP_422J2_124_3477_n315), .A2(
        DP_OP_422J2_124_3477_n316), .Y(DP_OP_422J2_124_3477_n105) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U96 ( .A1(DP_OP_422J2_124_3477_n316), .A2(
        DP_OP_422J2_124_3477_n315), .Y(DP_OP_422J2_124_3477_n102) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U87 ( .A1(DP_OP_422J2_124_3477_n313), .A2(
        DP_OP_422J2_124_3477_n314), .Y(DP_OP_422J2_124_3477_n98) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U86 ( .A1(DP_OP_422J2_124_3477_n314), .A2(
        DP_OP_422J2_124_3477_n313), .Y(DP_OP_422J2_124_3477_n97) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U82 ( .A1(DP_OP_422J2_124_3477_n97), .A2(
        DP_OP_422J2_124_3477_n102), .Y(DP_OP_422J2_124_3477_n95) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U75 ( .A1(DP_OP_422J2_124_3477_n311), .A2(
        DP_OP_422J2_124_3477_n312), .Y(DP_OP_422J2_124_3477_n89) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U68 ( .A1(DP_OP_422J2_124_3477_n95), .A2(
        n1587), .Y(DP_OP_422J2_124_3477_n82) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U61 ( .A1(DP_OP_422J2_124_3477_n309), .A2(
        DP_OP_422J2_124_3477_n310), .Y(DP_OP_422J2_124_3477_n78) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U60 ( .A1(DP_OP_422J2_124_3477_n310), .A2(
        DP_OP_422J2_124_3477_n309), .Y(DP_OP_422J2_124_3477_n77) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U54 ( .A1(DP_OP_422J2_124_3477_n111), .A2(
        DP_OP_422J2_124_3477_n75), .Y(DP_OP_422J2_124_3477_n73) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U45 ( .A1(n1383), .A2(
        DP_OP_422J2_124_3477_n308), .Y(DP_OP_422J2_124_3477_n65) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U38 ( .A1(DP_OP_422J2_124_3477_n71), .A2(
        n1586), .Y(DP_OP_422J2_124_3477_n60) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U34 ( .A1(n1592), .A2(
        DP_OP_422J2_124_3477_n58), .Y(DP_OP_422J2_124_3477_n56) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U29 ( .A1(DP_OP_422J2_124_3477_n305), .A2(
        DP_OP_422J2_124_3477_n306), .Y(DP_OP_422J2_124_3477_n52) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U28 ( .A1(DP_OP_422J2_124_3477_n306), .A2(
        DP_OP_422J2_124_3477_n305), .Y(DP_OP_422J2_124_3477_n51) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U21 ( .A1(DP_OP_422J2_124_3477_n303), .A2(
        DP_OP_422J2_124_3477_n304), .Y(DP_OP_422J2_124_3477_n47) );
  NAND2X0_HVT DP_OP_422J2_124_3477_U9 ( .A1(n1584), .A2(
        DP_OP_422J2_124_3477_n302), .Y(DP_OP_422J2_124_3477_n38) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2192 ( .A1(DP_OP_424J2_126_3477_n2977), 
        .A2(DP_OP_424J2_126_3477_n2979), .Y(DP_OP_424J2_126_3477_n2953) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2189 ( .A1(DP_OP_425J2_127_3477_n2182), 
        .A2(DP_OP_424J2_126_3477_n2979), .Y(DP_OP_423J2_125_3477_n2950) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2187 ( .A1(DP_OP_424J2_126_3477_n2972), 
        .A2(DP_OP_424J2_126_3477_n2979), .Y(DP_OP_424J2_126_3477_n2948) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2190 ( .A1(DP_OP_424J2_126_3477_n2975), 
        .A2(DP_OP_424J2_126_3477_n2979), .Y(DP_OP_424J2_126_3477_n2951) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2189 ( .A1(DP_OP_424J2_126_3477_n2974), 
        .A2(DP_OP_424J2_126_3477_n2979), .Y(DP_OP_424J2_126_3477_n2950) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2188 ( .A1(DP_OP_424J2_126_3477_n2973), 
        .A2(DP_OP_424J2_126_3477_n2979), .Y(DP_OP_424J2_126_3477_n2949) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2188 ( .A1(DP_OP_423J2_125_3477_n2973), 
        .A2(DP_OP_424J2_126_3477_n2979), .Y(DP_OP_423J2_125_3477_n2949) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1942 ( .A1(DP_OP_424J2_126_3477_n2315), 
        .A2(n597), .Y(DP_OP_425J2_127_3477_n2703) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1493 ( .A1(DP_OP_423J2_125_3477_n2886), 
        .A2(DP_OP_423J2_125_3477_n2276), .Y(DP_OP_425J2_127_3477_n2254) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1309 ( .A1(DP_OP_423J2_125_3477_n2006), 
        .A2(DP_OP_424J2_126_3477_n2099), .Y(DP_OP_424J2_126_3477_n2070) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1359 ( .A1(DP_OP_422J2_124_3477_n2004), 
        .A2(DP_OP_424J2_126_3477_n2144), .Y(DP_OP_425J2_127_3477_n2120) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1851 ( .A1(DP_OP_425J2_127_3477_n2620), 
        .A2(DP_OP_424J2_126_3477_n2629), .Y(DP_OP_425J2_127_3477_n2612) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1228 ( .A1(DP_OP_424J2_126_3477_n3059), 
        .A2(n558), .Y(DP_OP_425J2_127_3477_n1989) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1625 ( .A1(DP_OP_424J2_126_3477_n2534), 
        .A2(DP_OP_424J2_126_3477_n2408), .Y(DP_OP_422J2_124_3477_n2386) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2280 ( .A1(DP_OP_425J2_127_3477_n3063), 
        .A2(DP_OP_425J2_127_3477_n3065), .Y(DP_OP_425J2_127_3477_n3039) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1942 ( .A1(DP_OP_425J2_127_3477_n2447), 
        .A2(n596), .Y(DP_OP_423J2_125_3477_n2703) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1543 ( .A1(DP_OP_422J2_124_3477_n2312), 
        .A2(DP_OP_422J2_124_3477_n2321), .Y(DP_OP_422J2_124_3477_n2304) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1933 ( .A1(DP_OP_425J2_127_3477_n2710), 
        .A2(n1341), .Y(DP_OP_425J2_127_3477_n2694) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1837 ( .A1(DP_OP_425J2_127_3477_n2622), 
        .A2(DP_OP_423J2_125_3477_n2627), .Y(DP_OP_425J2_127_3477_n2598) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1500 ( .A1(DP_OP_425J2_127_3477_n2269), 
        .A2(DP_OP_424J2_126_3477_n2277), .Y(DP_OP_425J2_127_3477_n2261) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1799 ( .A1(DP_OP_422J2_124_3477_n2444), 
        .A2(n186), .Y(DP_OP_423J2_125_3477_n2560) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1312 ( .A1(DP_OP_423J2_125_3477_n3063), 
        .A2(DP_OP_425J2_127_3477_n2099), .Y(DP_OP_425J2_127_3477_n2073) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1500 ( .A1(DP_OP_422J2_124_3477_n2269), 
        .A2(DP_OP_422J2_124_3477_n2277), .Y(DP_OP_422J2_124_3477_n2261) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1939 ( .A1(DP_OP_422J2_124_3477_n2708), 
        .A2(n596), .Y(DP_OP_422J2_124_3477_n2700) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1985 ( .A1(DP_OP_423J2_125_3477_n2754), 
        .A2(n66), .Y(DP_OP_423J2_125_3477_n2746) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1221 ( .A1(DP_OP_424J2_126_3477_n3060), 
        .A2(DP_OP_425J2_127_3477_n2011), .Y(DP_OP_425J2_127_3477_n1982) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1502 ( .A1(DP_OP_423J2_125_3477_n2271), 
        .A2(DP_OP_423J2_125_3477_n2277), .Y(DP_OP_423J2_125_3477_n2263) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1221 ( .A1(DP_OP_422J2_124_3477_n2006), 
        .A2(DP_OP_422J2_124_3477_n2011), .Y(DP_OP_422J2_124_3477_n1982) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2278 ( .A1(DP_OP_425J2_127_3477_n3061), 
        .A2(DP_OP_425J2_127_3477_n3065), .Y(DP_OP_425J2_127_3477_n3037) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1493 ( .A1(DP_OP_422J2_124_3477_n2270), 
        .A2(DP_OP_422J2_124_3477_n2276), .Y(DP_OP_422J2_124_3477_n2254) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2064 ( .A1(DP_OP_425J2_127_3477_n2841), 
        .A2(DP_OP_425J2_127_3477_n2848), .Y(DP_OP_425J2_127_3477_n2825) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2280 ( .A1(DP_OP_423J2_125_3477_n3063), 
        .A2(DP_OP_423J2_125_3477_n3065), .Y(DP_OP_423J2_125_3477_n3039) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1360 ( .A1(DP_OP_425J2_127_3477_n2885), 
        .A2(DP_OP_424J2_126_3477_n2144), .Y(DP_OP_424J2_126_3477_n2121) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1984 ( .A1(DP_OP_424J2_126_3477_n2269), 
        .A2(n66), .Y(DP_OP_425J2_127_3477_n2745) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2116 ( .A1(DP_OP_422J2_124_3477_n2885), 
        .A2(DP_OP_422J2_124_3477_n2893), .Y(DP_OP_422J2_124_3477_n2877) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1977 ( .A1(DP_OP_425J2_127_3477_n2754), 
        .A2(DP_OP_425J2_127_3477_n2760), .Y(DP_OP_425J2_127_3477_n2738) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1451 ( .A1(DP_OP_423J2_125_3477_n2228), 
        .A2(n364), .Y(DP_OP_423J2_125_3477_n2212) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1935 ( .A1(DP_OP_423J2_125_3477_n2712), 
        .A2(DP_OP_424J2_126_3477_n2716), .Y(DP_OP_423J2_125_3477_n2696) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1492 ( .A1(DP_OP_422J2_124_3477_n2269), 
        .A2(DP_OP_422J2_124_3477_n2276), .Y(DP_OP_422J2_124_3477_n2253) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2250 ( .A1(DP_OP_423J2_125_3477_n3019), 
        .A2(DP_OP_423J2_125_3477_n3025), .Y(DP_OP_423J2_125_3477_n3011) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2119 ( .A1(DP_OP_425J2_127_3477_n2888), 
        .A2(DP_OP_425J2_127_3477_n2893), .Y(DP_OP_425J2_127_3477_n2880) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1396 ( .A1(DP_OP_423J2_125_3477_n2973), 
        .A2(n1339), .Y(DP_OP_425J2_127_3477_n2157) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1934 ( .A1(DP_OP_425J2_127_3477_n2447), 
        .A2(n1342), .Y(DP_OP_423J2_125_3477_n2695) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1449 ( .A1(DP_OP_425J2_127_3477_n2226), 
        .A2(n365), .Y(DP_OP_425J2_127_3477_n2210) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2016 ( .A1(DP_OP_423J2_125_3477_n2801), 
        .A2(DP_OP_423J2_125_3477_n2803), .Y(DP_OP_423J2_125_3477_n2777) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1986 ( .A1(DP_OP_425J2_127_3477_n2755), 
        .A2(n66), .Y(DP_OP_425J2_127_3477_n2747) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2292 ( .A1(DP_OP_425J2_127_3477_n3059), 
        .A2(n691), .Y(DP_OP_425J2_127_3477_n3051) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1838 ( .A1(DP_OP_423J2_125_3477_n2447), 
        .A2(DP_OP_422J2_124_3477_n2627), .Y(DP_OP_422J2_124_3477_n2599) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1309 ( .A1(DP_OP_425J2_127_3477_n2226), 
        .A2(DP_OP_424J2_126_3477_n2099), .Y(DP_OP_422J2_124_3477_n2070) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1360 ( .A1(DP_OP_424J2_126_3477_n2929), 
        .A2(DP_OP_425J2_127_3477_n2144), .Y(DP_OP_425J2_127_3477_n2121) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1266 ( .A1(DP_OP_424J2_126_3477_n3019), 
        .A2(DP_OP_425J2_127_3477_n2055), .Y(DP_OP_425J2_127_3477_n2027) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1265 ( .A1(DP_OP_425J2_127_3477_n2182), 
        .A2(DP_OP_422J2_124_3477_n2055), .Y(DP_OP_422J2_124_3477_n2026) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1676 ( .A1(DP_OP_425J2_127_3477_n2445), 
        .A2(DP_OP_425J2_127_3477_n2453), .Y(DP_OP_425J2_127_3477_n2437) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2067 ( .A1(DP_OP_423J2_125_3477_n2096), 
        .A2(DP_OP_425J2_127_3477_n2848), .Y(DP_OP_425J2_127_3477_n2828) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1620 ( .A1(DP_OP_423J2_125_3477_n2405), 
        .A2(n799), .Y(DP_OP_423J2_125_3477_n2381) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2118 ( .A1(DP_OP_423J2_125_3477_n2051), 
        .A2(DP_OP_425J2_127_3477_n2893), .Y(DP_OP_425J2_127_3477_n2879) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1361 ( .A1(DP_OP_425J2_127_3477_n2138), 
        .A2(DP_OP_422J2_124_3477_n2144), .Y(DP_OP_425J2_127_3477_n2122) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1224 ( .A1(DP_OP_424J2_126_3477_n3063), 
        .A2(DP_OP_425J2_127_3477_n2011), .Y(DP_OP_425J2_127_3477_n1985) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1231 ( .A1(DP_OP_425J2_127_3477_n2008), 
        .A2(n557), .Y(DP_OP_425J2_127_3477_n1992) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1263 ( .A1(DP_OP_425J2_127_3477_n2972), 
        .A2(DP_OP_424J2_126_3477_n2055), .Y(DP_OP_424J2_126_3477_n2024) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1268 ( .A1(DP_OP_425J2_127_3477_n2053), 
        .A2(DP_OP_425J2_127_3477_n2055), .Y(DP_OP_425J2_127_3477_n2029) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2278 ( .A1(DP_OP_423J2_125_3477_n2007), 
        .A2(DP_OP_425J2_127_3477_n3065), .Y(DP_OP_422J2_124_3477_n3037) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1626 ( .A1(DP_OP_422J2_124_3477_n2667), 
        .A2(DP_OP_424J2_126_3477_n2408), .Y(DP_OP_423J2_125_3477_n2387) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1504 ( .A1(DP_OP_424J2_126_3477_n2801), 
        .A2(DP_OP_422J2_124_3477_n2277), .Y(DP_OP_425J2_127_3477_n2265) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1546 ( .A1(DP_OP_423J2_125_3477_n2843), 
        .A2(DP_OP_425J2_127_3477_n2321), .Y(DP_OP_425J2_127_3477_n2307) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2065 ( .A1(DP_OP_423J2_125_3477_n2094), 
        .A2(DP_OP_425J2_127_3477_n2848), .Y(DP_OP_425J2_127_3477_n2826) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1450 ( .A1(DP_OP_423J2_125_3477_n2227), 
        .A2(n365), .Y(DP_OP_423J2_125_3477_n2211) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2115 ( .A1(DP_OP_423J2_125_3477_n2048), 
        .A2(DP_OP_425J2_127_3477_n2893), .Y(DP_OP_425J2_127_3477_n2876) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1835 ( .A1(DP_OP_423J2_125_3477_n2620), 
        .A2(DP_OP_423J2_125_3477_n2627), .Y(DP_OP_423J2_125_3477_n2596) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1495 ( .A1(DP_OP_425J2_127_3477_n2272), 
        .A2(DP_OP_423J2_125_3477_n2276), .Y(DP_OP_425J2_127_3477_n2256) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1617 ( .A1(DP_OP_423J2_125_3477_n2754), 
        .A2(n799), .Y(DP_OP_425J2_127_3477_n2378) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1502 ( .A1(DP_OP_424J2_126_3477_n2799), 
        .A2(DP_OP_423J2_125_3477_n2277), .Y(DP_OP_425J2_127_3477_n2263) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1840 ( .A1(DP_OP_423J2_125_3477_n2625), 
        .A2(DP_OP_423J2_125_3477_n2627), .Y(DP_OP_423J2_125_3477_n2601) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1932 ( .A1(DP_OP_422J2_124_3477_n2709), 
        .A2(n1340), .Y(DP_OP_422J2_124_3477_n2693) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1840 ( .A1(DP_OP_423J2_125_3477_n2317), 
        .A2(DP_OP_423J2_125_3477_n2627), .Y(DP_OP_425J2_127_3477_n2601) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1404 ( .A1(DP_OP_423J2_125_3477_n2973), 
        .A2(n1343), .Y(DP_OP_425J2_127_3477_n2165) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1404 ( .A1(DP_OP_422J2_124_3477_n2181), 
        .A2(n1345), .Y(DP_OP_422J2_124_3477_n2165) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2162 ( .A1(DP_OP_423J2_125_3477_n2931), 
        .A2(n445), .Y(DP_OP_423J2_125_3477_n2923) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1359 ( .A1(DP_OP_424J2_126_3477_n2136), 
        .A2(DP_OP_425J2_127_3477_n2144), .Y(DP_OP_424J2_126_3477_n2120) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1397 ( .A1(DP_OP_425J2_127_3477_n2182), 
        .A2(n1339), .Y(DP_OP_425J2_127_3477_n2158) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1627 ( .A1(DP_OP_425J2_127_3477_n2404), 
        .A2(n1333), .Y(DP_OP_425J2_127_3477_n2388) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1397 ( .A1(DP_OP_424J2_126_3477_n2754), 
        .A2(n1339), .Y(DP_OP_422J2_124_3477_n2158) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1835 ( .A1(DP_OP_425J2_127_3477_n2620), 
        .A2(DP_OP_423J2_125_3477_n2627), .Y(DP_OP_425J2_127_3477_n2596) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2016 ( .A1(DP_OP_425J2_127_3477_n2801), 
        .A2(n1444), .Y(DP_OP_425J2_127_3477_n2777) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1801 ( .A1(DP_OP_425J2_127_3477_n2578), 
        .A2(n186), .Y(DP_OP_425J2_127_3477_n2562) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1309 ( .A1(DP_OP_423J2_125_3477_n3060), 
        .A2(DP_OP_425J2_127_3477_n2099), .Y(DP_OP_425J2_127_3477_n2070) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2118 ( .A1(DP_OP_423J2_125_3477_n2887), 
        .A2(DP_OP_425J2_127_3477_n2893), .Y(DP_OP_423J2_125_3477_n2879) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1266 ( .A1(DP_OP_422J2_124_3477_n2051), 
        .A2(DP_OP_422J2_124_3477_n2055), .Y(DP_OP_422J2_124_3477_n2027) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1492 ( .A1(DP_OP_424J2_126_3477_n2269), 
        .A2(DP_OP_424J2_126_3477_n2276), .Y(DP_OP_424J2_126_3477_n2253) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2030 ( .A1(DP_OP_423J2_125_3477_n2799), 
        .A2(DP_OP_423J2_125_3477_n2805), .Y(DP_OP_423J2_125_3477_n2791) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1838 ( .A1(DP_OP_423J2_125_3477_n2315), 
        .A2(DP_OP_424J2_126_3477_n2627), .Y(DP_OP_425J2_127_3477_n2599) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2027 ( .A1(DP_OP_424J2_126_3477_n2796), 
        .A2(DP_OP_424J2_126_3477_n2805), .Y(DP_OP_424J2_126_3477_n2788) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1222 ( .A1(DP_OP_425J2_127_3477_n2007), 
        .A2(DP_OP_425J2_127_3477_n2011), .Y(DP_OP_425J2_127_3477_n1983) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2117 ( .A1(DP_OP_423J2_125_3477_n2886), 
        .A2(DP_OP_422J2_124_3477_n2893), .Y(DP_OP_423J2_125_3477_n2878) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1588 ( .A1(DP_OP_425J2_127_3477_n2357), 
        .A2(DP_OP_425J2_127_3477_n2365), .Y(DP_OP_425J2_127_3477_n2349) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2277 ( .A1(DP_OP_424J2_126_3477_n3060), 
        .A2(DP_OP_424J2_126_3477_n3065), .Y(DP_OP_424J2_126_3477_n3036) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1265 ( .A1(DP_OP_425J2_127_3477_n2974), 
        .A2(DP_OP_424J2_126_3477_n2055), .Y(DP_OP_424J2_126_3477_n2026) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1219 ( .A1(DP_OP_422J2_124_3477_n3058), 
        .A2(DP_OP_422J2_124_3477_n2011), .Y(DP_OP_423J2_125_3477_n1980) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1492 ( .A1(DP_OP_425J2_127_3477_n2269), 
        .A2(DP_OP_423J2_125_3477_n2276), .Y(DP_OP_425J2_127_3477_n2253) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2296 ( .A1(DP_OP_422J2_124_3477_n3063), 
        .A2(n32), .Y(DP_OP_422J2_124_3477_n3055) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2275 ( .A1(DP_OP_425J2_127_3477_n2092), 
        .A2(DP_OP_423J2_125_3477_n3065), .Y(DP_OP_423J2_125_3477_n3034) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1932 ( .A1(DP_OP_425J2_127_3477_n2357), 
        .A2(n1342), .Y(DP_OP_424J2_126_3477_n2693) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1231 ( .A1(DP_OP_423J2_125_3477_n2008), 
        .A2(n558), .Y(DP_OP_423J2_125_3477_n1992) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1984 ( .A1(DP_OP_425J2_127_3477_n2401), 
        .A2(n66), .Y(DP_OP_423J2_125_3477_n2745) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2116 ( .A1(DP_OP_425J2_127_3477_n2269), 
        .A2(DP_OP_422J2_124_3477_n2893), .Y(DP_OP_423J2_125_3477_n2877) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2247 ( .A1(DP_OP_425J2_127_3477_n2048), 
        .A2(DP_OP_424J2_126_3477_n3025), .Y(DP_OP_424J2_126_3477_n3008) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2027 ( .A1(DP_OP_425J2_127_3477_n2796), 
        .A2(DP_OP_423J2_125_3477_n2805), .Y(DP_OP_425J2_127_3477_n2788) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1448 ( .A1(DP_OP_425J2_127_3477_n2797), 
        .A2(n365), .Y(DP_OP_424J2_126_3477_n2209) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1624 ( .A1(DP_OP_422J2_124_3477_n2753), 
        .A2(n1333), .Y(DP_OP_424J2_126_3477_n2385) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1803 ( .A1(DP_OP_422J2_124_3477_n2448), 
        .A2(n186), .Y(DP_OP_423J2_125_3477_n2564) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1265 ( .A1(DP_OP_425J2_127_3477_n2050), 
        .A2(DP_OP_425J2_127_3477_n2055), .Y(DP_OP_425J2_127_3477_n2026) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1988 ( .A1(DP_OP_424J2_126_3477_n2405), 
        .A2(n66), .Y(DP_OP_422J2_124_3477_n2749) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2249 ( .A1(DP_OP_425J2_127_3477_n2138), 
        .A2(DP_OP_423J2_125_3477_n3025), .Y(DP_OP_423J2_125_3477_n3010) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1944 ( .A1(DP_OP_423J2_125_3477_n2361), 
        .A2(n597), .Y(DP_OP_422J2_124_3477_n2705) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1616 ( .A1(DP_OP_423J2_125_3477_n2401), 
        .A2(n798), .Y(DP_OP_423J2_125_3477_n2377) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1675 ( .A1(DP_OP_422J2_124_3477_n2312), 
        .A2(DP_OP_425J2_127_3477_n2453), .Y(DP_OP_425J2_127_3477_n2436) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2155 ( .A1(DP_OP_423J2_125_3477_n2932), 
        .A2(DP_OP_423J2_125_3477_n2936), .Y(DP_OP_423J2_125_3477_n2916) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1398 ( .A1(DP_OP_425J2_127_3477_n2755), 
        .A2(n1339), .Y(DP_OP_423J2_125_3477_n2159) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1548 ( .A1(DP_OP_423J2_125_3477_n2713), 
        .A2(DP_OP_422J2_124_3477_n2321), .Y(DP_OP_422J2_124_3477_n2309) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2028 ( .A1(DP_OP_425J2_127_3477_n2797), 
        .A2(DP_OP_424J2_126_3477_n2805), .Y(DP_OP_425J2_127_3477_n2789) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1501 ( .A1(DP_OP_424J2_126_3477_n2358), 
        .A2(DP_OP_423J2_125_3477_n2277), .Y(DP_OP_423J2_125_3477_n2262) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1407 ( .A1(DP_OP_422J2_124_3477_n2888), 
        .A2(n1343), .Y(DP_OP_423J2_125_3477_n2168) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1592 ( .A1(DP_OP_425J2_127_3477_n2493), 
        .A2(DP_OP_425J2_127_3477_n2365), .Y(DP_OP_422J2_124_3477_n2353) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1852 ( .A1(DP_OP_425J2_127_3477_n2621), 
        .A2(DP_OP_423J2_125_3477_n2629), .Y(DP_OP_425J2_127_3477_n2613) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1263 ( .A1(DP_OP_425J2_127_3477_n2048), 
        .A2(DP_OP_425J2_127_3477_n2055), .Y(DP_OP_425J2_127_3477_n2024) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2067 ( .A1(DP_OP_423J2_125_3477_n2844), 
        .A2(DP_OP_425J2_127_3477_n2848), .Y(DP_OP_423J2_125_3477_n2828) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2120 ( .A1(DP_OP_422J2_124_3477_n2889), 
        .A2(DP_OP_422J2_124_3477_n2893), .Y(DP_OP_422J2_124_3477_n2881) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1618 ( .A1(DP_OP_425J2_127_3477_n2403), 
        .A2(n792), .Y(DP_OP_425J2_127_3477_n2379) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1940 ( .A1(DP_OP_423J2_125_3477_n2225), 
        .A2(n597), .Y(DP_OP_425J2_127_3477_n2701) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1494 ( .A1(DP_OP_423J2_125_3477_n2271), 
        .A2(DP_OP_423J2_125_3477_n2276), .Y(DP_OP_423J2_125_3477_n2255) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1224 ( .A1(DP_OP_425J2_127_3477_n2933), 
        .A2(DP_OP_425J2_127_3477_n2011), .Y(DP_OP_423J2_125_3477_n1985) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2160 ( .A1(DP_OP_423J2_125_3477_n2005), 
        .A2(n446), .Y(DP_OP_425J2_127_3477_n2921) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1976 ( .A1(DP_OP_424J2_126_3477_n2269), 
        .A2(DP_OP_425J2_127_3477_n2760), .Y(DP_OP_425J2_127_3477_n2737) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1543 ( .A1(DP_OP_425J2_127_3477_n2708), 
        .A2(DP_OP_422J2_124_3477_n2321), .Y(DP_OP_424J2_126_3477_n2304) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2152 ( .A1(DP_OP_424J2_126_3477_n2929), 
        .A2(DP_OP_424J2_126_3477_n2936), .Y(DP_OP_424J2_126_3477_n2913) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1839 ( .A1(DP_OP_423J2_125_3477_n2624), 
        .A2(DP_OP_423J2_125_3477_n2627), .Y(DP_OP_423J2_125_3477_n2600) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1543 ( .A1(DP_OP_425J2_127_3477_n2312), 
        .A2(DP_OP_425J2_127_3477_n2321), .Y(DP_OP_425J2_127_3477_n2304) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1800 ( .A1(DP_OP_422J2_124_3477_n2577), 
        .A2(n186), .Y(DP_OP_422J2_124_3477_n2561) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1615 ( .A1(DP_OP_425J2_127_3477_n2400), 
        .A2(n799), .Y(DP_OP_425J2_127_3477_n2376) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1617 ( .A1(DP_OP_424J2_126_3477_n2534), 
        .A2(n798), .Y(DP_OP_422J2_124_3477_n2378) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2115 ( .A1(DP_OP_422J2_124_3477_n2884), 
        .A2(DP_OP_422J2_124_3477_n2893), .Y(DP_OP_422J2_124_3477_n2876) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1363 ( .A1(DP_OP_423J2_125_3477_n2140), 
        .A2(DP_OP_422J2_124_3477_n2144), .Y(DP_OP_423J2_125_3477_n2124) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2277 ( .A1(DP_OP_422J2_124_3477_n3060), 
        .A2(DP_OP_425J2_127_3477_n3065), .Y(DP_OP_422J2_124_3477_n3036) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1264 ( .A1(DP_OP_422J2_124_3477_n3017), 
        .A2(DP_OP_424J2_126_3477_n2055), .Y(DP_OP_423J2_125_3477_n2025) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1398 ( .A1(DP_OP_422J2_124_3477_n2183), 
        .A2(n1339), .Y(DP_OP_422J2_124_3477_n2159) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1267 ( .A1(DP_OP_425J2_127_3477_n2184), 
        .A2(DP_OP_422J2_124_3477_n2055), .Y(DP_OP_422J2_124_3477_n2028) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1221 ( .A1(DP_OP_424J2_126_3477_n2006), 
        .A2(DP_OP_424J2_126_3477_n2011), .Y(DP_OP_424J2_126_3477_n1982) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2151 ( .A1(DP_OP_422J2_124_3477_n2092), 
        .A2(DP_OP_423J2_125_3477_n2936), .Y(DP_OP_423J2_125_3477_n2912) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2294 ( .A1(DP_OP_423J2_125_3477_n3061), 
        .A2(n34), .Y(DP_OP_423J2_125_3477_n3053) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1678 ( .A1(DP_OP_423J2_125_3477_n2447), 
        .A2(DP_OP_425J2_127_3477_n2453), .Y(DP_OP_423J2_125_3477_n2439) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1228 ( .A1(DP_OP_422J2_124_3477_n2005), 
        .A2(n558), .Y(DP_OP_422J2_124_3477_n1989) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1499 ( .A1(DP_OP_422J2_124_3477_n2268), 
        .A2(DP_OP_422J2_124_3477_n2277), .Y(DP_OP_422J2_124_3477_n2260) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1851 ( .A1(DP_OP_422J2_124_3477_n2312), 
        .A2(DP_OP_424J2_126_3477_n2629), .Y(DP_OP_424J2_126_3477_n2612) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2164 ( .A1(DP_OP_425J2_127_3477_n2801), 
        .A2(n446), .Y(DP_OP_422J2_124_3477_n2925) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1448 ( .A1(DP_OP_422J2_124_3477_n2225), 
        .A2(DP_OP_423J2_125_3477_n2232), .Y(DP_OP_422J2_124_3477_n2209) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1802 ( .A1(DP_OP_423J2_125_3477_n2579), 
        .A2(n186), .Y(DP_OP_423J2_125_3477_n2563) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2115 ( .A1(DP_OP_425J2_127_3477_n2180), 
        .A2(DP_OP_424J2_126_3477_n2893), .Y(DP_OP_424J2_126_3477_n2876) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1310 ( .A1(DP_OP_423J2_125_3477_n3061), 
        .A2(DP_OP_425J2_127_3477_n2099), .Y(DP_OP_425J2_127_3477_n2071) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1617 ( .A1(DP_OP_422J2_124_3477_n2754), 
        .A2(DP_OP_422J2_124_3477_n2407), .Y(DP_OP_424J2_126_3477_n2378) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2252 ( .A1(DP_OP_422J2_124_3477_n3021), 
        .A2(n846), .Y(DP_OP_422J2_124_3477_n3013) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1800 ( .A1(DP_OP_425J2_127_3477_n2577), 
        .A2(n186), .Y(DP_OP_425J2_127_3477_n2561) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2116 ( .A1(DP_OP_425J2_127_3477_n2885), 
        .A2(DP_OP_425J2_127_3477_n2893), .Y(DP_OP_425J2_127_3477_n2877) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1853 ( .A1(DP_OP_422J2_124_3477_n2622), 
        .A2(DP_OP_422J2_124_3477_n2629), .Y(DP_OP_422J2_124_3477_n2614) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1404 ( .A1(DP_OP_422J2_124_3477_n2973), 
        .A2(n1344), .Y(DP_OP_424J2_126_3477_n2165) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1397 ( .A1(DP_OP_422J2_124_3477_n2974), 
        .A2(n1339), .Y(DP_OP_424J2_126_3477_n2158) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2248 ( .A1(DP_OP_424J2_126_3477_n2005), 
        .A2(DP_OP_425J2_127_3477_n3025), .Y(DP_OP_425J2_127_3477_n3009) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1837 ( .A1(DP_OP_422J2_124_3477_n2622), 
        .A2(DP_OP_422J2_124_3477_n2627), .Y(DP_OP_422J2_124_3477_n2598) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1395 ( .A1(DP_OP_425J2_127_3477_n2180), 
        .A2(n1339), .Y(DP_OP_425J2_127_3477_n2156) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1932 ( .A1(DP_OP_422J2_124_3477_n2841), 
        .A2(n1340), .Y(DP_OP_425J2_127_3477_n2693) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1800 ( .A1(DP_OP_423J2_125_3477_n2665), 
        .A2(DP_OP_424J2_126_3477_n2584), .Y(DP_OP_424J2_126_3477_n2561) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1399 ( .A1(DP_OP_422J2_124_3477_n2888), 
        .A2(n1339), .Y(DP_OP_423J2_125_3477_n2160) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1400 ( .A1(DP_OP_423J2_125_3477_n2185), 
        .A2(n1339), .Y(DP_OP_423J2_125_3477_n2161) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1939 ( .A1(DP_OP_425J2_127_3477_n2708), 
        .A2(n597), .Y(DP_OP_425J2_127_3477_n2700) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2277 ( .A1(DP_OP_425J2_127_3477_n3060), 
        .A2(DP_OP_425J2_127_3477_n3065), .Y(DP_OP_425J2_127_3477_n3036) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1359 ( .A1(DP_OP_425J2_127_3477_n2268), 
        .A2(DP_OP_424J2_126_3477_n2144), .Y(DP_OP_422J2_124_3477_n2120) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1268 ( .A1(DP_OP_423J2_125_3477_n2053), 
        .A2(DP_OP_425J2_127_3477_n2055), .Y(DP_OP_423J2_125_3477_n2029) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1544 ( .A1(DP_OP_423J2_125_3477_n2841), 
        .A2(DP_OP_425J2_127_3477_n2321), .Y(DP_OP_425J2_127_3477_n2305) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1307 ( .A1(DP_OP_425J2_127_3477_n2092), 
        .A2(DP_OP_425J2_127_3477_n2099), .Y(DP_OP_425J2_127_3477_n2068) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1449 ( .A1(DP_OP_423J2_125_3477_n2798), 
        .A2(n365), .Y(DP_OP_422J2_124_3477_n2210) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1504 ( .A1(DP_OP_423J2_125_3477_n2757), 
        .A2(DP_OP_422J2_124_3477_n2277), .Y(DP_OP_422J2_124_3477_n2265) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1448 ( .A1(DP_OP_422J2_124_3477_n2093), 
        .A2(n365), .Y(DP_OP_425J2_127_3477_n2209) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2247 ( .A1(DP_OP_424J2_126_3477_n2004), 
        .A2(DP_OP_425J2_127_3477_n3025), .Y(DP_OP_425J2_127_3477_n3008) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1495 ( .A1(DP_OP_423J2_125_3477_n2272), 
        .A2(DP_OP_423J2_125_3477_n2276), .Y(DP_OP_423J2_125_3477_n2256) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1229 ( .A1(DP_OP_424J2_126_3477_n3060), 
        .A2(n558), .Y(DP_OP_425J2_127_3477_n1990) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1624 ( .A1(DP_OP_422J2_124_3477_n2401), 
        .A2(n1346), .Y(DP_OP_422J2_124_3477_n2385) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1228 ( .A1(DP_OP_424J2_126_3477_n2005), 
        .A2(n558), .Y(DP_OP_424J2_126_3477_n1989) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2248 ( .A1(DP_OP_422J2_124_3477_n3017), 
        .A2(DP_OP_425J2_127_3477_n3025), .Y(DP_OP_422J2_124_3477_n3009) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2279 ( .A1(DP_OP_423J2_125_3477_n3062), 
        .A2(DP_OP_423J2_125_3477_n3065), .Y(DP_OP_423J2_125_3477_n3038) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1624 ( .A1(DP_OP_425J2_127_3477_n2401), 
        .A2(DP_OP_424J2_126_3477_n2408), .Y(DP_OP_425J2_127_3477_n2385) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1837 ( .A1(DP_OP_424J2_126_3477_n2622), 
        .A2(DP_OP_424J2_126_3477_n2627), .Y(DP_OP_424J2_126_3477_n2598) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1627 ( .A1(DP_OP_423J2_125_3477_n2404), 
        .A2(n1346), .Y(DP_OP_423J2_125_3477_n2388) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1801 ( .A1(DP_OP_422J2_124_3477_n2578), 
        .A2(n186), .Y(DP_OP_422J2_124_3477_n2562) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1223 ( .A1(DP_OP_424J2_126_3477_n2932), 
        .A2(DP_OP_422J2_124_3477_n2011), .Y(DP_OP_422J2_124_3477_n1984) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2247 ( .A1(DP_OP_424J2_126_3477_n2136), 
        .A2(DP_OP_423J2_125_3477_n3025), .Y(DP_OP_422J2_124_3477_n3008) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1446 ( .A1(DP_OP_422J2_124_3477_n2091), 
        .A2(n365), .Y(DP_OP_425J2_127_3477_n2207) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1230 ( .A1(DP_OP_422J2_124_3477_n2007), 
        .A2(n558), .Y(DP_OP_422J2_124_3477_n1991) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1405 ( .A1(DP_OP_425J2_127_3477_n2182), 
        .A2(n1345), .Y(DP_OP_425J2_127_3477_n2166) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1627 ( .A1(DP_OP_422J2_124_3477_n2404), 
        .A2(DP_OP_424J2_126_3477_n2408), .Y(DP_OP_422J2_124_3477_n2388) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1359 ( .A1(DP_OP_425J2_127_3477_n2796), 
        .A2(DP_OP_422J2_124_3477_n2144), .Y(DP_OP_423J2_125_3477_n2120) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2032 ( .A1(DP_OP_425J2_127_3477_n2801), 
        .A2(DP_OP_423J2_125_3477_n2805), .Y(DP_OP_425J2_127_3477_n2793) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1944 ( .A1(DP_OP_423J2_125_3477_n2229), 
        .A2(n597), .Y(DP_OP_425J2_127_3477_n2705) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1988 ( .A1(DP_OP_422J2_124_3477_n2889), 
        .A2(n66), .Y(DP_OP_425J2_127_3477_n2749) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1680 ( .A1(DP_OP_425J2_127_3477_n2449), 
        .A2(DP_OP_425J2_127_3477_n2453), .Y(DP_OP_425J2_127_3477_n2441) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1361 ( .A1(DP_OP_422J2_124_3477_n2930), 
        .A2(DP_OP_425J2_127_3477_n2144), .Y(DP_OP_423J2_125_3477_n2122) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1501 ( .A1(DP_OP_423J2_125_3477_n2182), 
        .A2(DP_OP_424J2_126_3477_n2277), .Y(DP_OP_424J2_126_3477_n2262) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1396 ( .A1(DP_OP_424J2_126_3477_n2269), 
        .A2(n1339), .Y(DP_OP_423J2_125_3477_n2157) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1494 ( .A1(DP_OP_425J2_127_3477_n2755), 
        .A2(DP_OP_424J2_126_3477_n2276), .Y(DP_OP_424J2_126_3477_n2255) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1839 ( .A1(DP_OP_423J2_125_3477_n2712), 
        .A2(DP_OP_424J2_126_3477_n2627), .Y(DP_OP_424J2_126_3477_n2600) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2117 ( .A1(DP_OP_424J2_126_3477_n2886), 
        .A2(DP_OP_424J2_126_3477_n2893), .Y(DP_OP_424J2_126_3477_n2878) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1220 ( .A1(DP_OP_422J2_124_3477_n2005), 
        .A2(DP_OP_422J2_124_3477_n2011), .Y(DP_OP_422J2_124_3477_n1981) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1308 ( .A1(DP_OP_423J2_125_3477_n3059), 
        .A2(DP_OP_425J2_127_3477_n2099), .Y(DP_OP_425J2_127_3477_n2069) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2249 ( .A1(DP_OP_425J2_127_3477_n2050), 
        .A2(DP_OP_424J2_126_3477_n3025), .Y(DP_OP_424J2_126_3477_n3010) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1934 ( .A1(DP_OP_424J2_126_3477_n2315), 
        .A2(n1342), .Y(DP_OP_425J2_127_3477_n2695) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1399 ( .A1(DP_OP_424J2_126_3477_n2184), 
        .A2(n1339), .Y(DP_OP_424J2_126_3477_n2160) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2279 ( .A1(DP_OP_425J2_127_3477_n2008), 
        .A2(DP_OP_424J2_126_3477_n3065), .Y(DP_OP_424J2_126_3477_n3038) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1802 ( .A1(DP_OP_424J2_126_3477_n2579), 
        .A2(n186), .Y(DP_OP_424J2_126_3477_n2563) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1589 ( .A1(DP_OP_424J2_126_3477_n2358), 
        .A2(DP_OP_424J2_126_3477_n2365), .Y(DP_OP_424J2_126_3477_n2350) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2276 ( .A1(DP_OP_423J2_125_3477_n3059), 
        .A2(DP_OP_423J2_125_3477_n3065), .Y(DP_OP_423J2_125_3477_n3035) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1450 ( .A1(DP_OP_425J2_127_3477_n2799), 
        .A2(n365), .Y(DP_OP_424J2_126_3477_n2211) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1985 ( .A1(DP_OP_424J2_126_3477_n2754), 
        .A2(n66), .Y(DP_OP_424J2_126_3477_n2746) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1626 ( .A1(DP_OP_424J2_126_3477_n2403), 
        .A2(n1346), .Y(DP_OP_424J2_126_3477_n2387) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1934 ( .A1(DP_OP_425J2_127_3477_n2359), 
        .A2(n1341), .Y(DP_OP_424J2_126_3477_n2695) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1941 ( .A1(DP_OP_423J2_125_3477_n2798), 
        .A2(n597), .Y(DP_OP_424J2_126_3477_n2702) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1406 ( .A1(DP_OP_422J2_124_3477_n2975), 
        .A2(n1345), .Y(DP_OP_424J2_126_3477_n2167) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1978 ( .A1(DP_OP_422J2_124_3477_n2183), 
        .A2(DP_OP_425J2_127_3477_n2760), .Y(DP_OP_424J2_126_3477_n2739) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2154 ( .A1(DP_OP_422J2_124_3477_n2007), 
        .A2(DP_OP_424J2_126_3477_n2936), .Y(DP_OP_424J2_126_3477_n2915) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1545 ( .A1(DP_OP_425J2_127_3477_n2710), 
        .A2(DP_OP_423J2_125_3477_n2321), .Y(DP_OP_424J2_126_3477_n2306) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2029 ( .A1(DP_OP_422J2_124_3477_n2138), 
        .A2(DP_OP_424J2_126_3477_n2805), .Y(DP_OP_424J2_126_3477_n2790) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2247 ( .A1(DP_OP_422J2_124_3477_n2004), 
        .A2(DP_OP_423J2_125_3477_n3025), .Y(DP_OP_423J2_125_3477_n3008) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2277 ( .A1(DP_OP_423J2_125_3477_n3060), 
        .A2(DP_OP_423J2_125_3477_n3065), .Y(DP_OP_423J2_125_3477_n3036) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1619 ( .A1(DP_OP_422J2_124_3477_n2756), 
        .A2(n799), .Y(DP_OP_424J2_126_3477_n2380) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1499 ( .A1(DP_OP_423J2_125_3477_n2268), 
        .A2(DP_OP_423J2_125_3477_n2277), .Y(DP_OP_423J2_125_3477_n2260) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1362 ( .A1(DP_OP_423J2_125_3477_n2051), 
        .A2(DP_OP_424J2_126_3477_n2144), .Y(DP_OP_424J2_126_3477_n2123) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2293 ( .A1(DP_OP_424J2_126_3477_n3060), 
        .A2(n693), .Y(DP_OP_424J2_126_3477_n3052) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2161 ( .A1(DP_OP_425J2_127_3477_n2138), 
        .A2(n446), .Y(DP_OP_424J2_126_3477_n2922) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1311 ( .A1(DP_OP_423J2_125_3477_n2008), 
        .A2(DP_OP_424J2_126_3477_n2099), .Y(DP_OP_424J2_126_3477_n2072) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1223 ( .A1(DP_OP_425J2_127_3477_n3020), 
        .A2(DP_OP_424J2_126_3477_n2011), .Y(DP_OP_424J2_126_3477_n1984) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1618 ( .A1(DP_OP_424J2_126_3477_n2403), 
        .A2(n799), .Y(DP_OP_424J2_126_3477_n2379) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2278 ( .A1(DP_OP_423J2_125_3477_n3061), 
        .A2(DP_OP_423J2_125_3477_n3065), .Y(DP_OP_423J2_125_3477_n3037) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1616 ( .A1(DP_OP_422J2_124_3477_n2401), 
        .A2(n797), .Y(DP_OP_422J2_124_3477_n2377) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2028 ( .A1(DP_OP_425J2_127_3477_n2269), 
        .A2(DP_OP_424J2_126_3477_n2805), .Y(DP_OP_424J2_126_3477_n2789) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1222 ( .A1(DP_OP_425J2_127_3477_n3019), 
        .A2(DP_OP_424J2_126_3477_n2011), .Y(DP_OP_424J2_126_3477_n1983) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1229 ( .A1(DP_OP_424J2_126_3477_n2006), 
        .A2(DP_OP_423J2_125_3477_n2012), .Y(DP_OP_424J2_126_3477_n1990) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1944 ( .A1(DP_OP_423J2_125_3477_n2713), 
        .A2(n597), .Y(DP_OP_423J2_125_3477_n2705) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1933 ( .A1(DP_OP_423J2_125_3477_n2798), 
        .A2(n1342), .Y(DP_OP_424J2_126_3477_n2694) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1988 ( .A1(DP_OP_423J2_125_3477_n2757), 
        .A2(n66), .Y(DP_OP_423J2_125_3477_n2749) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1361 ( .A1(DP_OP_424J2_126_3477_n2138), 
        .A2(DP_OP_425J2_127_3477_n2144), .Y(DP_OP_424J2_126_3477_n2122) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1220 ( .A1(DP_OP_423J2_125_3477_n2005), 
        .A2(DP_OP_422J2_124_3477_n2011), .Y(DP_OP_423J2_125_3477_n1981) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1852 ( .A1(DP_OP_425J2_127_3477_n2445), 
        .A2(DP_OP_424J2_126_3477_n2629), .Y(DP_OP_424J2_126_3477_n2613) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1838 ( .A1(DP_OP_424J2_126_3477_n2623), 
        .A2(DP_OP_424J2_126_3477_n2627), .Y(DP_OP_424J2_126_3477_n2599) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2014 ( .A1(DP_OP_424J2_126_3477_n2799), 
        .A2(DP_OP_423J2_125_3477_n2803), .Y(DP_OP_424J2_126_3477_n2775) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2120 ( .A1(DP_OP_423J2_125_3477_n2889), 
        .A2(DP_OP_422J2_124_3477_n2893), .Y(DP_OP_423J2_125_3477_n2881) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1310 ( .A1(DP_OP_424J2_126_3477_n2095), 
        .A2(DP_OP_424J2_126_3477_n2099), .Y(DP_OP_424J2_126_3477_n2071) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2248 ( .A1(DP_OP_425J2_127_3477_n2049), 
        .A2(DP_OP_424J2_126_3477_n3025), .Y(DP_OP_424J2_126_3477_n3009) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2278 ( .A1(DP_OP_425J2_127_3477_n2007), 
        .A2(DP_OP_424J2_126_3477_n3065), .Y(DP_OP_424J2_126_3477_n3037) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1504 ( .A1(DP_OP_423J2_125_3477_n2273), 
        .A2(DP_OP_423J2_125_3477_n2277), .Y(DP_OP_423J2_125_3477_n2265) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1500 ( .A1(DP_OP_424J2_126_3477_n2269), 
        .A2(DP_OP_424J2_126_3477_n2277), .Y(DP_OP_424J2_126_3477_n2261) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1493 ( .A1(DP_OP_423J2_125_3477_n2182), 
        .A2(DP_OP_424J2_126_3477_n2276), .Y(DP_OP_424J2_126_3477_n2254) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1452 ( .A1(DP_OP_423J2_125_3477_n2801), 
        .A2(n365), .Y(DP_OP_422J2_124_3477_n2213) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2162 ( .A1(DP_OP_425J2_127_3477_n2799), 
        .A2(n445), .Y(DP_OP_422J2_124_3477_n2923) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1403 ( .A1(DP_OP_425J2_127_3477_n2180), 
        .A2(n1344), .Y(DP_OP_425J2_127_3477_n2164) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1496 ( .A1(DP_OP_424J2_126_3477_n2669), 
        .A2(DP_OP_422J2_124_3477_n2276), .Y(DP_OP_422J2_124_3477_n2257) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1266 ( .A1(DP_OP_424J2_126_3477_n2051), 
        .A2(DP_OP_424J2_126_3477_n2055), .Y(DP_OP_424J2_126_3477_n2027) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2164 ( .A1(DP_OP_424J2_126_3477_n2845), 
        .A2(n446), .Y(DP_OP_423J2_125_3477_n2925) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2292 ( .A1(DP_OP_424J2_126_3477_n3059), 
        .A2(n694), .Y(DP_OP_424J2_126_3477_n3051) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1449 ( .A1(DP_OP_422J2_124_3477_n2930), 
        .A2(n364), .Y(DP_OP_424J2_126_3477_n2210) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2252 ( .A1(DP_OP_423J2_125_3477_n3021), 
        .A2(DP_OP_423J2_125_3477_n3025), .Y(DP_OP_423J2_125_3477_n3013) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2248 ( .A1(DP_OP_424J2_126_3477_n2929), 
        .A2(DP_OP_423J2_125_3477_n3025), .Y(DP_OP_423J2_125_3477_n3009) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1836 ( .A1(DP_OP_422J2_124_3477_n2621), 
        .A2(DP_OP_422J2_124_3477_n2627), .Y(DP_OP_422J2_124_3477_n2597) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1503 ( .A1(DP_OP_425J2_127_3477_n2404), 
        .A2(DP_OP_422J2_124_3477_n2277), .Y(DP_OP_422J2_124_3477_n2264) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1801 ( .A1(DP_OP_423J2_125_3477_n2666), 
        .A2(n186), .Y(DP_OP_424J2_126_3477_n2562) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1931 ( .A1(DP_OP_422J2_124_3477_n2708), 
        .A2(DP_OP_424J2_126_3477_n2716), .Y(DP_OP_422J2_124_3477_n2692) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1451 ( .A1(DP_OP_424J2_126_3477_n2712), 
        .A2(n364), .Y(DP_OP_422J2_124_3477_n2212) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1547 ( .A1(DP_OP_425J2_127_3477_n2448), 
        .A2(DP_OP_422J2_124_3477_n2321), .Y(DP_OP_422J2_124_3477_n2308) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1591 ( .A1(DP_OP_424J2_126_3477_n2580), 
        .A2(DP_OP_425J2_127_3477_n2365), .Y(DP_OP_422J2_124_3477_n2352) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1628 ( .A1(DP_OP_422J2_124_3477_n2405), 
        .A2(n1346), .Y(DP_OP_422J2_124_3477_n2389) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1984 ( .A1(DP_OP_422J2_124_3477_n2181), 
        .A2(DP_OP_425J2_127_3477_n2761), .Y(DP_OP_424J2_126_3477_n2745) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2276 ( .A1(DP_OP_425J2_127_3477_n3059), 
        .A2(DP_OP_425J2_127_3477_n3065), .Y(DP_OP_425J2_127_3477_n3035) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2116 ( .A1(DP_OP_423J2_125_3477_n2973), 
        .A2(DP_OP_424J2_126_3477_n2893), .Y(DP_OP_424J2_126_3477_n2877) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1398 ( .A1(DP_OP_422J2_124_3477_n2975), 
        .A2(n1339), .Y(DP_OP_424J2_126_3477_n2159) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1447 ( .A1(DP_OP_422J2_124_3477_n2840), 
        .A2(n365), .Y(DP_OP_423J2_125_3477_n2208) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1804 ( .A1(DP_OP_423J2_125_3477_n2493), 
        .A2(DP_OP_424J2_126_3477_n2584), .Y(DP_OP_422J2_124_3477_n2565) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1835 ( .A1(DP_OP_422J2_124_3477_n2620), 
        .A2(DP_OP_422J2_124_3477_n2627), .Y(DP_OP_422J2_124_3477_n2596) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2031 ( .A1(DP_OP_422J2_124_3477_n2800), 
        .A2(DP_OP_422J2_124_3477_n2805), .Y(DP_OP_422J2_124_3477_n2792) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1623 ( .A1(DP_OP_425J2_127_3477_n2400), 
        .A2(DP_OP_424J2_126_3477_n2408), .Y(DP_OP_425J2_127_3477_n2384) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1943 ( .A1(DP_OP_425J2_127_3477_n2712), 
        .A2(n597), .Y(DP_OP_425J2_127_3477_n2704) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1936 ( .A1(DP_OP_424J2_126_3477_n2317), 
        .A2(n1341), .Y(DP_OP_425J2_127_3477_n2697) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2119 ( .A1(DP_OP_422J2_124_3477_n2888), 
        .A2(DP_OP_422J2_124_3477_n2893), .Y(DP_OP_422J2_124_3477_n2880) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1230 ( .A1(DP_OP_425J2_127_3477_n3019), 
        .A2(n558), .Y(DP_OP_424J2_126_3477_n1991) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2276 ( .A1(DP_OP_422J2_124_3477_n3059), 
        .A2(DP_OP_425J2_127_3477_n3065), .Y(DP_OP_422J2_124_3477_n3035) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1618 ( .A1(DP_OP_424J2_126_3477_n2491), 
        .A2(n794), .Y(DP_OP_423J2_125_3477_n2379) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1227 ( .A1(DP_OP_422J2_124_3477_n2004), 
        .A2(n556), .Y(DP_OP_422J2_124_3477_n1988) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2294 ( .A1(DP_OP_425J2_127_3477_n2007), 
        .A2(n694), .Y(DP_OP_424J2_126_3477_n3053) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2066 ( .A1(DP_OP_425J2_127_3477_n2843), 
        .A2(DP_OP_425J2_127_3477_n2848), .Y(DP_OP_425J2_127_3477_n2827) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1501 ( .A1(DP_OP_422J2_124_3477_n2270), 
        .A2(DP_OP_422J2_124_3477_n2277), .Y(DP_OP_422J2_124_3477_n2262) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1854 ( .A1(DP_OP_424J2_126_3477_n2623), 
        .A2(DP_OP_424J2_126_3477_n2629), .Y(DP_OP_424J2_126_3477_n2615) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2162 ( .A1(DP_OP_423J2_125_3477_n3019), 
        .A2(n445), .Y(DP_OP_424J2_126_3477_n2923) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2161 ( .A1(DP_OP_422J2_124_3477_n2930), 
        .A2(n446), .Y(DP_OP_422J2_124_3477_n2922) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1545 ( .A1(DP_OP_423J2_125_3477_n2842), 
        .A2(DP_OP_425J2_127_3477_n2321), .Y(DP_OP_425J2_127_3477_n2306) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1620 ( .A1(DP_OP_424J2_126_3477_n2405), 
        .A2(n799), .Y(DP_OP_424J2_126_3477_n2381) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1590 ( .A1(DP_OP_422J2_124_3477_n2799), 
        .A2(DP_OP_425J2_127_3477_n2365), .Y(DP_OP_424J2_126_3477_n2351) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1494 ( .A1(DP_OP_425J2_127_3477_n2403), 
        .A2(DP_OP_422J2_124_3477_n2276), .Y(DP_OP_422J2_124_3477_n2255) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1545 ( .A1(DP_OP_422J2_124_3477_n2314), 
        .A2(DP_OP_422J2_124_3477_n2321), .Y(DP_OP_422J2_124_3477_n2306) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2161 ( .A1(DP_OP_423J2_125_3477_n2006), 
        .A2(n446), .Y(DP_OP_425J2_127_3477_n2922) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2156 ( .A1(DP_OP_424J2_126_3477_n2933), 
        .A2(DP_OP_424J2_126_3477_n2936), .Y(DP_OP_424J2_126_3477_n2917) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1936 ( .A1(DP_OP_423J2_125_3477_n2801), 
        .A2(n1341), .Y(DP_OP_424J2_126_3477_n2697) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1627 ( .A1(DP_OP_422J2_124_3477_n2756), 
        .A2(n1333), .Y(DP_OP_424J2_126_3477_n2388) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1839 ( .A1(DP_OP_423J2_125_3477_n2448), 
        .A2(DP_OP_422J2_124_3477_n2627), .Y(DP_OP_422J2_124_3477_n2600) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1800 ( .A1(DP_OP_422J2_124_3477_n2445), 
        .A2(n186), .Y(DP_OP_423J2_125_3477_n2561) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1941 ( .A1(DP_OP_422J2_124_3477_n2710), 
        .A2(n597), .Y(DP_OP_422J2_124_3477_n2702) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1223 ( .A1(DP_OP_425J2_127_3477_n2008), 
        .A2(DP_OP_425J2_127_3477_n2011), .Y(DP_OP_425J2_127_3477_n1984) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2117 ( .A1(DP_OP_423J2_125_3477_n2182), 
        .A2(DP_OP_422J2_124_3477_n2893), .Y(DP_OP_422J2_124_3477_n2878) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1230 ( .A1(DP_OP_425J2_127_3477_n2007), 
        .A2(n558), .Y(DP_OP_425J2_127_3477_n1991) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1267 ( .A1(DP_OP_424J2_126_3477_n3020), 
        .A2(DP_OP_425J2_127_3477_n2055), .Y(DP_OP_425J2_127_3477_n2028) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1451 ( .A1(DP_OP_425J2_127_3477_n2800), 
        .A2(DP_OP_423J2_125_3477_n2232), .Y(DP_OP_424J2_126_3477_n2212) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1221 ( .A1(DP_OP_423J2_125_3477_n2006), 
        .A2(DP_OP_424J2_126_3477_n2011), .Y(DP_OP_423J2_125_3477_n1982) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2249 ( .A1(DP_OP_424J2_126_3477_n2138), 
        .A2(DP_OP_423J2_125_3477_n3025), .Y(DP_OP_422J2_124_3477_n3010) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1232 ( .A1(DP_OP_425J2_127_3477_n3021), 
        .A2(n558), .Y(DP_OP_424J2_126_3477_n1993) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1406 ( .A1(DP_OP_422J2_124_3477_n2183), 
        .A2(n1344), .Y(DP_OP_422J2_124_3477_n2167) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2016 ( .A1(DP_OP_424J2_126_3477_n2801), 
        .A2(DP_OP_423J2_125_3477_n2803), .Y(DP_OP_424J2_126_3477_n2777) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1399 ( .A1(DP_OP_424J2_126_3477_n2756), 
        .A2(n1339), .Y(DP_OP_422J2_124_3477_n2160) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1362 ( .A1(DP_OP_422J2_124_3477_n2007), 
        .A2(DP_OP_425J2_127_3477_n2144), .Y(DP_OP_425J2_127_3477_n2123) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2293 ( .A1(DP_OP_425J2_127_3477_n3060), 
        .A2(n693), .Y(DP_OP_425J2_127_3477_n3052) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2163 ( .A1(DP_OP_424J2_126_3477_n2932), 
        .A2(n446), .Y(DP_OP_424J2_126_3477_n2924) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2250 ( .A1(DP_OP_424J2_126_3477_n3019), 
        .A2(DP_OP_424J2_126_3477_n3025), .Y(DP_OP_424J2_126_3477_n3011) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1935 ( .A1(DP_OP_424J2_126_3477_n2712), 
        .A2(DP_OP_424J2_126_3477_n2716), .Y(DP_OP_424J2_126_3477_n2696) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1307 ( .A1(DP_OP_422J2_124_3477_n2092), 
        .A2(DP_OP_424J2_126_3477_n2099), .Y(DP_OP_422J2_124_3477_n2068) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2279 ( .A1(DP_OP_423J2_125_3477_n2008), 
        .A2(DP_OP_423J2_125_3477_n3065), .Y(DP_OP_422J2_124_3477_n3038) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1626 ( .A1(DP_OP_424J2_126_3477_n2535), 
        .A2(n1346), .Y(DP_OP_422J2_124_3477_n2387) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1802 ( .A1(DP_OP_422J2_124_3477_n2579), 
        .A2(n185), .Y(DP_OP_422J2_124_3477_n2563) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2118 ( .A1(DP_OP_424J2_126_3477_n2887), 
        .A2(DP_OP_424J2_126_3477_n2893), .Y(DP_OP_424J2_126_3477_n2879) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1364 ( .A1(DP_OP_422J2_124_3477_n3021), 
        .A2(DP_OP_424J2_126_3477_n2144), .Y(DP_OP_424J2_126_3477_n2125) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1224 ( .A1(DP_OP_425J2_127_3477_n3021), 
        .A2(DP_OP_424J2_126_3477_n2011), .Y(DP_OP_424J2_126_3477_n1985) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1978 ( .A1(DP_OP_425J2_127_3477_n2755), 
        .A2(DP_OP_425J2_127_3477_n2760), .Y(DP_OP_425J2_127_3477_n2739) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1987 ( .A1(DP_OP_424J2_126_3477_n2756), 
        .A2(n66), .Y(DP_OP_424J2_126_3477_n2748) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1231 ( .A1(DP_OP_425J2_127_3477_n3020), 
        .A2(n557), .Y(DP_OP_424J2_126_3477_n1992) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1308 ( .A1(DP_OP_422J2_124_3477_n2093), 
        .A2(DP_OP_425J2_127_3477_n2099), .Y(DP_OP_422J2_124_3477_n2069) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1268 ( .A1(DP_OP_425J2_127_3477_n2977), 
        .A2(DP_OP_424J2_126_3477_n2055), .Y(DP_OP_424J2_126_3477_n2029) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2295 ( .A1(DP_OP_425J2_127_3477_n2008), 
        .A2(n34), .Y(DP_OP_424J2_126_3477_n3054) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1311 ( .A1(DP_OP_423J2_125_3477_n3062), 
        .A2(DP_OP_425J2_127_3477_n2099), .Y(DP_OP_425J2_127_3477_n2072) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1589 ( .A1(DP_OP_422J2_124_3477_n2358), 
        .A2(DP_OP_425J2_127_3477_n2365), .Y(DP_OP_422J2_124_3477_n2350) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2119 ( .A1(DP_OP_425J2_127_3477_n2184), 
        .A2(DP_OP_424J2_126_3477_n2893), .Y(DP_OP_424J2_126_3477_n2880) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1408 ( .A1(DP_OP_424J2_126_3477_n2185), 
        .A2(DP_OP_425J2_127_3477_n2188), .Y(DP_OP_424J2_126_3477_n2169) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1853 ( .A1(DP_OP_425J2_127_3477_n2622), 
        .A2(DP_OP_424J2_126_3477_n2629), .Y(DP_OP_425J2_127_3477_n2614) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2251 ( .A1(DP_OP_424J2_126_3477_n3020), 
        .A2(DP_OP_424J2_126_3477_n3025), .Y(DP_OP_424J2_126_3477_n3012) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1855 ( .A1(DP_OP_425J2_127_3477_n2448), 
        .A2(DP_OP_424J2_126_3477_n2629), .Y(DP_OP_424J2_126_3477_n2616) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2031 ( .A1(DP_OP_422J2_124_3477_n2140), 
        .A2(DP_OP_424J2_126_3477_n2805), .Y(DP_OP_424J2_126_3477_n2792) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1804 ( .A1(DP_OP_425J2_127_3477_n2493), 
        .A2(n186), .Y(DP_OP_424J2_126_3477_n2565) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2160 ( .A1(DP_OP_422J2_124_3477_n2093), 
        .A2(n446), .Y(DP_OP_423J2_125_3477_n2921) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1934 ( .A1(DP_OP_424J2_126_3477_n2447), 
        .A2(n1340), .Y(DP_OP_422J2_124_3477_n2695) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1591 ( .A1(DP_OP_423J2_125_3477_n2272), 
        .A2(DP_OP_425J2_127_3477_n2365), .Y(DP_OP_424J2_126_3477_n2352) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1228 ( .A1(DP_OP_423J2_125_3477_n2005), 
        .A2(n558), .Y(DP_OP_423J2_125_3477_n1989) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1547 ( .A1(DP_OP_423J2_125_3477_n2228), 
        .A2(DP_OP_422J2_124_3477_n2321), .Y(DP_OP_424J2_126_3477_n2308) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1450 ( .A1(DP_OP_423J2_125_3477_n2799), 
        .A2(n365), .Y(DP_OP_422J2_124_3477_n2211) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1503 ( .A1(DP_OP_425J2_127_3477_n2756), 
        .A2(DP_OP_424J2_126_3477_n2277), .Y(DP_OP_424J2_126_3477_n2264) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1496 ( .A1(DP_OP_422J2_124_3477_n2889), 
        .A2(DP_OP_424J2_126_3477_n2276), .Y(DP_OP_424J2_126_3477_n2257) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1452 ( .A1(DP_OP_425J2_127_3477_n2801), 
        .A2(n365), .Y(DP_OP_424J2_126_3477_n2213) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2029 ( .A1(DP_OP_425J2_127_3477_n2798), 
        .A2(DP_OP_424J2_126_3477_n2805), .Y(DP_OP_425J2_127_3477_n2790) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1837 ( .A1(DP_OP_423J2_125_3477_n2622), 
        .A2(DP_OP_423J2_125_3477_n2627), .Y(DP_OP_423J2_125_3477_n2598) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1548 ( .A1(DP_OP_423J2_125_3477_n2845), 
        .A2(DP_OP_425J2_127_3477_n2321), .Y(DP_OP_425J2_127_3477_n2309) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2120 ( .A1(DP_OP_422J2_124_3477_n3021), 
        .A2(DP_OP_425J2_127_3477_n2893), .Y(DP_OP_425J2_127_3477_n2881) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2296 ( .A1(DP_OP_425J2_127_3477_n3063), 
        .A2(n34), .Y(DP_OP_425J2_127_3477_n3055) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1446 ( .A1(DP_OP_422J2_124_3477_n2223), 
        .A2(n365), .Y(DP_OP_422J2_124_3477_n2207) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1985 ( .A1(DP_OP_422J2_124_3477_n2754), 
        .A2(n66), .Y(DP_OP_422J2_124_3477_n2746) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2252 ( .A1(DP_OP_425J2_127_3477_n3021), 
        .A2(DP_OP_425J2_127_3477_n3025), .Y(DP_OP_425J2_127_3477_n3013) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1856 ( .A1(DP_OP_423J2_125_3477_n2317), 
        .A2(DP_OP_423J2_125_3477_n2629), .Y(DP_OP_425J2_127_3477_n2617) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2015 ( .A1(DP_OP_422J2_124_3477_n2800), 
        .A2(DP_OP_422J2_124_3477_n2803), .Y(DP_OP_422J2_124_3477_n2776) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2164 ( .A1(DP_OP_425J2_127_3477_n2933), 
        .A2(n446), .Y(DP_OP_425J2_127_3477_n2925) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2153 ( .A1(DP_OP_425J2_127_3477_n2226), 
        .A2(DP_OP_423J2_125_3477_n2936), .Y(DP_OP_423J2_125_3477_n2914) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1447 ( .A1(DP_OP_422J2_124_3477_n2224), 
        .A2(n364), .Y(DP_OP_422J2_124_3477_n2208) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1267 ( .A1(DP_OP_425J2_127_3477_n2976), 
        .A2(DP_OP_424J2_126_3477_n2055), .Y(DP_OP_424J2_126_3477_n2028) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1853 ( .A1(DP_OP_424J2_126_3477_n2622), 
        .A2(DP_OP_424J2_126_3477_n2629), .Y(DP_OP_424J2_126_3477_n2614) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1396 ( .A1(DP_OP_422J2_124_3477_n2181), 
        .A2(n1339), .Y(DP_OP_422J2_124_3477_n2157) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2252 ( .A1(DP_OP_425J2_127_3477_n2053), 
        .A2(DP_OP_424J2_126_3477_n3025), .Y(DP_OP_424J2_126_3477_n3013) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2164 ( .A1(DP_OP_424J2_126_3477_n2933), 
        .A2(n445), .Y(DP_OP_424J2_126_3477_n2925) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1263 ( .A1(DP_OP_422J2_124_3477_n2048), 
        .A2(DP_OP_422J2_124_3477_n2055), .Y(DP_OP_422J2_124_3477_n2024) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1360 ( .A1(DP_OP_425J2_127_3477_n2797), 
        .A2(DP_OP_424J2_126_3477_n2144), .Y(DP_OP_423J2_125_3477_n2121) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1405 ( .A1(DP_OP_423J2_125_3477_n2182), 
        .A2(n1343), .Y(DP_OP_423J2_125_3477_n2166) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1491 ( .A1(DP_OP_425J2_127_3477_n2268), 
        .A2(DP_OP_422J2_124_3477_n2276), .Y(DP_OP_425J2_127_3477_n2252) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1504 ( .A1(DP_OP_422J2_124_3477_n2889), 
        .A2(DP_OP_424J2_126_3477_n2277), .Y(DP_OP_424J2_126_3477_n2265) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1856 ( .A1(DP_OP_425J2_127_3477_n2449), 
        .A2(DP_OP_424J2_126_3477_n2629), .Y(DP_OP_424J2_126_3477_n2617) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2296 ( .A1(DP_OP_424J2_126_3477_n3063), 
        .A2(n693), .Y(DP_OP_424J2_126_3477_n3055) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1501 ( .A1(DP_OP_423J2_125_3477_n2886), 
        .A2(DP_OP_424J2_126_3477_n2277), .Y(DP_OP_425J2_127_3477_n2262) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2120 ( .A1(DP_OP_424J2_126_3477_n2889), 
        .A2(DP_OP_424J2_126_3477_n2893), .Y(DP_OP_424J2_126_3477_n2881) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2152 ( .A1(DP_OP_422J2_124_3477_n2093), 
        .A2(DP_OP_423J2_125_3477_n2936), .Y(DP_OP_423J2_125_3477_n2913) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1592 ( .A1(DP_OP_423J2_125_3477_n2273), 
        .A2(DP_OP_425J2_127_3477_n2365), .Y(DP_OP_424J2_126_3477_n2353) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1494 ( .A1(DP_OP_424J2_126_3477_n2799), 
        .A2(DP_OP_422J2_124_3477_n2276), .Y(DP_OP_425J2_127_3477_n2255) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1548 ( .A1(DP_OP_424J2_126_3477_n2317), 
        .A2(DP_OP_422J2_124_3477_n2321), .Y(DP_OP_424J2_126_3477_n2309) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1933 ( .A1(DP_OP_422J2_124_3477_n2314), 
        .A2(n1340), .Y(DP_OP_423J2_125_3477_n2694) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1839 ( .A1(DP_OP_423J2_125_3477_n2316), 
        .A2(DP_OP_424J2_126_3477_n2627), .Y(DP_OP_425J2_127_3477_n2600) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2117 ( .A1(DP_OP_425J2_127_3477_n2886), 
        .A2(DP_OP_425J2_127_3477_n2893), .Y(DP_OP_425J2_127_3477_n2878) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1229 ( .A1(DP_OP_423J2_125_3477_n2006), 
        .A2(n558), .Y(DP_OP_423J2_125_3477_n1990) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2249 ( .A1(DP_OP_424J2_126_3477_n2006), 
        .A2(DP_OP_425J2_127_3477_n3025), .Y(DP_OP_425J2_127_3477_n3010) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1265 ( .A1(DP_OP_424J2_126_3477_n2138), 
        .A2(DP_OP_422J2_124_3477_n2055), .Y(DP_OP_423J2_125_3477_n2026) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1399 ( .A1(DP_OP_425J2_127_3477_n2184), 
        .A2(n1339), .Y(DP_OP_425J2_127_3477_n2160) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1546 ( .A1(DP_OP_424J2_126_3477_n2315), 
        .A2(DP_OP_425J2_127_3477_n2321), .Y(DP_OP_424J2_126_3477_n2307) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1406 ( .A1(DP_OP_422J2_124_3477_n2051), 
        .A2(n1345), .Y(DP_OP_425J2_127_3477_n2167) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1988 ( .A1(DP_OP_422J2_124_3477_n2185), 
        .A2(n66), .Y(DP_OP_424J2_126_3477_n2749) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1495 ( .A1(DP_OP_422J2_124_3477_n2888), 
        .A2(DP_OP_424J2_126_3477_n2276), .Y(DP_OP_424J2_126_3477_n2256) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2279 ( .A1(DP_OP_425J2_127_3477_n3062), 
        .A2(DP_OP_425J2_127_3477_n3065), .Y(DP_OP_425J2_127_3477_n3038) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1502 ( .A1(DP_OP_425J2_127_3477_n2755), 
        .A2(DP_OP_424J2_126_3477_n2277), .Y(DP_OP_424J2_126_3477_n2263) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2032 ( .A1(DP_OP_424J2_126_3477_n2801), 
        .A2(DP_OP_424J2_126_3477_n2805), .Y(DP_OP_424J2_126_3477_n2793) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1840 ( .A1(DP_OP_425J2_127_3477_n2449), 
        .A2(DP_OP_424J2_126_3477_n2627), .Y(DP_OP_424J2_126_3477_n2601) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1222 ( .A1(DP_OP_423J2_125_3477_n2007), 
        .A2(DP_OP_422J2_124_3477_n2011), .Y(DP_OP_423J2_125_3477_n1983) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1802 ( .A1(DP_OP_425J2_127_3477_n2579), 
        .A2(n186), .Y(DP_OP_425J2_127_3477_n2563) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1619 ( .A1(DP_OP_422J2_124_3477_n2404), 
        .A2(n799), .Y(DP_OP_422J2_124_3477_n2380) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1397 ( .A1(DP_OP_423J2_125_3477_n2182), 
        .A2(n1339), .Y(DP_OP_423J2_125_3477_n2158) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1450 ( .A1(DP_OP_423J2_125_3477_n2931), 
        .A2(n365), .Y(DP_OP_425J2_127_3477_n2211) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1404 ( .A1(DP_OP_424J2_126_3477_n2269), 
        .A2(n1345), .Y(DP_OP_423J2_125_3477_n2165) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1932 ( .A1(DP_OP_425J2_127_3477_n2445), 
        .A2(n1341), .Y(DP_OP_423J2_125_3477_n2693) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1939 ( .A1(DP_OP_423J2_125_3477_n2708), 
        .A2(n597), .Y(DP_OP_423J2_125_3477_n2700) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1403 ( .A1(DP_OP_424J2_126_3477_n2752), 
        .A2(DP_OP_425J2_127_3477_n2188), .Y(DP_OP_422J2_124_3477_n2164) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2293 ( .A1(DP_OP_422J2_124_3477_n3060), 
        .A2(n34), .Y(DP_OP_422J2_124_3477_n3052) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1362 ( .A1(DP_OP_424J2_126_3477_n2799), 
        .A2(DP_OP_425J2_127_3477_n2144), .Y(DP_OP_422J2_124_3477_n2123) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1227 ( .A1(DP_OP_424J2_126_3477_n3058), 
        .A2(n558), .Y(DP_OP_425J2_127_3477_n1988) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1985 ( .A1(DP_OP_425J2_127_3477_n2754), 
        .A2(n66), .Y(DP_OP_425J2_127_3477_n2746) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2115 ( .A1(DP_OP_425J2_127_3477_n2268), 
        .A2(DP_OP_424J2_126_3477_n2893), .Y(DP_OP_423J2_125_3477_n2876) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1312 ( .A1(DP_OP_422J2_124_3477_n3063), 
        .A2(DP_OP_424J2_126_3477_n2099), .Y(DP_OP_424J2_126_3477_n2073) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2280 ( .A1(DP_OP_424J2_126_3477_n3063), 
        .A2(DP_OP_424J2_126_3477_n3065), .Y(DP_OP_424J2_126_3477_n3039) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1448 ( .A1(DP_OP_423J2_125_3477_n2225), 
        .A2(n365), .Y(DP_OP_423J2_125_3477_n2209) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1626 ( .A1(DP_OP_425J2_127_3477_n2403), 
        .A2(n1333), .Y(DP_OP_425J2_127_3477_n2387) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1942 ( .A1(DP_OP_425J2_127_3477_n2359), 
        .A2(n596), .Y(DP_OP_424J2_126_3477_n2703) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1407 ( .A1(DP_OP_424J2_126_3477_n2184), 
        .A2(n1344), .Y(DP_OP_424J2_126_3477_n2168) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1400 ( .A1(DP_OP_424J2_126_3477_n2185), 
        .A2(n1339), .Y(DP_OP_424J2_126_3477_n2161) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1363 ( .A1(DP_OP_423J2_125_3477_n2052), 
        .A2(DP_OP_424J2_126_3477_n2144), .Y(DP_OP_424J2_126_3477_n2124) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1615 ( .A1(DP_OP_424J2_126_3477_n2532), 
        .A2(n799), .Y(DP_OP_422J2_124_3477_n2376) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1986 ( .A1(DP_OP_422J2_124_3477_n2183), 
        .A2(DP_OP_425J2_127_3477_n2761), .Y(DP_OP_424J2_126_3477_n2747) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2155 ( .A1(DP_OP_424J2_126_3477_n2932), 
        .A2(DP_OP_424J2_126_3477_n2936), .Y(DP_OP_424J2_126_3477_n2916) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2030 ( .A1(DP_OP_424J2_126_3477_n2799), 
        .A2(DP_OP_424J2_126_3477_n2805), .Y(DP_OP_424J2_126_3477_n2791) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1677 ( .A1(DP_OP_424J2_126_3477_n2622), 
        .A2(DP_OP_425J2_127_3477_n2453), .Y(DP_OP_425J2_127_3477_n2438) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1803 ( .A1(DP_OP_424J2_126_3477_n2580), 
        .A2(DP_OP_424J2_126_3477_n2584), .Y(DP_OP_424J2_126_3477_n2564) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1941 ( .A1(DP_OP_425J2_127_3477_n2710), 
        .A2(n597), .Y(DP_OP_425J2_127_3477_n2702) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2294 ( .A1(DP_OP_425J2_127_3477_n3061), 
        .A2(n34), .Y(DP_OP_425J2_127_3477_n3053) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1935 ( .A1(DP_OP_425J2_127_3477_n2712), 
        .A2(DP_OP_424J2_126_3477_n2716), .Y(DP_OP_425J2_127_3477_n2696) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1931 ( .A1(DP_OP_425J2_127_3477_n2708), 
        .A2(n1340), .Y(DP_OP_425J2_127_3477_n2692) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1618 ( .A1(DP_OP_424J2_126_3477_n2535), 
        .A2(n799), .Y(DP_OP_422J2_124_3477_n2379) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1625 ( .A1(DP_OP_425J2_127_3477_n2534), 
        .A2(DP_OP_424J2_126_3477_n2408), .Y(DP_OP_423J2_125_3477_n2386) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1836 ( .A1(DP_OP_425J2_127_3477_n2621), 
        .A2(DP_OP_423J2_125_3477_n2627), .Y(DP_OP_425J2_127_3477_n2597) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1232 ( .A1(DP_OP_423J2_125_3477_n3021), 
        .A2(n557), .Y(DP_OP_422J2_124_3477_n1993) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1803 ( .A1(DP_OP_422J2_124_3477_n2580), 
        .A2(n185), .Y(DP_OP_422J2_124_3477_n2564) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1588 ( .A1(DP_OP_422J2_124_3477_n2357), 
        .A2(DP_OP_425J2_127_3477_n2365), .Y(DP_OP_422J2_124_3477_n2349) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1801 ( .A1(DP_OP_422J2_124_3477_n2446), 
        .A2(n186), .Y(DP_OP_423J2_125_3477_n2562) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2163 ( .A1(DP_OP_425J2_127_3477_n2800), 
        .A2(n445), .Y(DP_OP_422J2_124_3477_n2924) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1449 ( .A1(DP_OP_425J2_127_3477_n2710), 
        .A2(n365), .Y(DP_OP_423J2_125_3477_n2210) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2292 ( .A1(DP_OP_423J2_125_3477_n3059), 
        .A2(n34), .Y(DP_OP_423J2_125_3477_n3051) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1362 ( .A1(DP_OP_425J2_127_3477_n2799), 
        .A2(DP_OP_422J2_124_3477_n2144), .Y(DP_OP_423J2_125_3477_n2123) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2293 ( .A1(DP_OP_423J2_125_3477_n3060), 
        .A2(n34), .Y(DP_OP_423J2_125_3477_n3052) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2280 ( .A1(DP_OP_422J2_124_3477_n3063), 
        .A2(DP_OP_424J2_126_3477_n3065), .Y(DP_OP_422J2_124_3477_n3039) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2161 ( .A1(DP_OP_425J2_127_3477_n2226), 
        .A2(n446), .Y(DP_OP_423J2_125_3477_n2922) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1855 ( .A1(DP_OP_423J2_125_3477_n2316), 
        .A2(DP_OP_424J2_126_3477_n2629), .Y(DP_OP_425J2_127_3477_n2616) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1942 ( .A1(DP_OP_425J2_127_3477_n2579), 
        .A2(n596), .Y(DP_OP_422J2_124_3477_n2703) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2031 ( .A1(DP_OP_425J2_127_3477_n2800), 
        .A2(DP_OP_424J2_126_3477_n2805), .Y(DP_OP_425J2_127_3477_n2792) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1619 ( .A1(DP_OP_423J2_125_3477_n2404), 
        .A2(n799), .Y(DP_OP_423J2_125_3477_n2380) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1804 ( .A1(DP_OP_425J2_127_3477_n2581), 
        .A2(n186), .Y(DP_OP_425J2_127_3477_n2565) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1364 ( .A1(DP_OP_423J2_125_3477_n2889), 
        .A2(DP_OP_422J2_124_3477_n2144), .Y(DP_OP_422J2_124_3477_n2125) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1361 ( .A1(DP_OP_422J2_124_3477_n2138), 
        .A2(DP_OP_422J2_124_3477_n2144), .Y(DP_OP_422J2_124_3477_n2122) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1407 ( .A1(DP_OP_424J2_126_3477_n2756), 
        .A2(DP_OP_425J2_127_3477_n2188), .Y(DP_OP_422J2_124_3477_n2168) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1616 ( .A1(DP_OP_425J2_127_3477_n2401), 
        .A2(n799), .Y(DP_OP_425J2_127_3477_n2377) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1547 ( .A1(DP_OP_423J2_125_3477_n2844), 
        .A2(DP_OP_425J2_127_3477_n2321), .Y(DP_OP_425J2_127_3477_n2308) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1503 ( .A1(DP_OP_425J2_127_3477_n2272), 
        .A2(DP_OP_422J2_124_3477_n2277), .Y(DP_OP_425J2_127_3477_n2264) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1266 ( .A1(DP_OP_423J2_125_3477_n2051), 
        .A2(DP_OP_422J2_124_3477_n2055), .Y(DP_OP_423J2_125_3477_n2027) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1400 ( .A1(DP_OP_422J2_124_3477_n2185), 
        .A2(n1339), .Y(DP_OP_422J2_124_3477_n2161) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1987 ( .A1(DP_OP_422J2_124_3477_n2756), 
        .A2(n66), .Y(DP_OP_422J2_124_3477_n2748) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1496 ( .A1(DP_OP_424J2_126_3477_n2801), 
        .A2(DP_OP_423J2_125_3477_n2276), .Y(DP_OP_425J2_127_3477_n2257) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1363 ( .A1(DP_OP_422J2_124_3477_n2140), 
        .A2(DP_OP_425J2_127_3477_n2144), .Y(DP_OP_422J2_124_3477_n2124) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1452 ( .A1(DP_OP_424J2_126_3477_n2845), 
        .A2(n365), .Y(DP_OP_425J2_127_3477_n2213) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1219 ( .A1(DP_OP_422J2_124_3477_n2004), 
        .A2(DP_OP_422J2_124_3477_n2011), .Y(DP_OP_422J2_124_3477_n1980) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1676 ( .A1(DP_OP_422J2_124_3477_n2621), 
        .A2(DP_OP_425J2_127_3477_n2453), .Y(DP_OP_423J2_125_3477_n2437) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2295 ( .A1(DP_OP_423J2_125_3477_n2008), 
        .A2(n34), .Y(DP_OP_422J2_124_3477_n3054) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2250 ( .A1(DP_OP_425J2_127_3477_n3019), 
        .A2(DP_OP_425J2_127_3477_n3025), .Y(DP_OP_425J2_127_3477_n3011) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1979 ( .A1(DP_OP_425J2_127_3477_n2756), 
        .A2(DP_OP_425J2_127_3477_n2760), .Y(DP_OP_425J2_127_3477_n2740) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1677 ( .A1(DP_OP_422J2_124_3477_n2622), 
        .A2(DP_OP_425J2_127_3477_n2453), .Y(DP_OP_423J2_125_3477_n2438) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2275 ( .A1(DP_OP_422J2_124_3477_n3058), 
        .A2(DP_OP_425J2_127_3477_n3065), .Y(DP_OP_422J2_124_3477_n3034) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1803 ( .A1(DP_OP_425J2_127_3477_n2580), 
        .A2(n186), .Y(DP_OP_425J2_127_3477_n2564) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1220 ( .A1(DP_OP_424J2_126_3477_n3059), 
        .A2(DP_OP_425J2_127_3477_n2011), .Y(DP_OP_425J2_127_3477_n1981) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1615 ( .A1(DP_OP_424J2_126_3477_n2400), 
        .A2(n799), .Y(DP_OP_424J2_126_3477_n2376) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1941 ( .A1(DP_OP_424J2_126_3477_n2622), 
        .A2(n597), .Y(DP_OP_423J2_125_3477_n2702) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1678 ( .A1(DP_OP_425J2_127_3477_n2447), 
        .A2(DP_OP_425J2_127_3477_n2453), .Y(DP_OP_425J2_127_3477_n2439) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1983 ( .A1(DP_OP_424J2_126_3477_n2400), 
        .A2(DP_OP_425J2_127_3477_n2761), .Y(DP_OP_422J2_124_3477_n2744) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1307 ( .A1(DP_OP_424J2_126_3477_n2092), 
        .A2(DP_OP_424J2_126_3477_n2099), .Y(DP_OP_424J2_126_3477_n2068) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2275 ( .A1(DP_OP_425J2_127_3477_n3058), 
        .A2(DP_OP_425J2_127_3477_n3065), .Y(DP_OP_425J2_127_3477_n3034) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1407 ( .A1(DP_OP_425J2_127_3477_n2184), 
        .A2(n1344), .Y(DP_OP_425J2_127_3477_n2168) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1406 ( .A1(DP_OP_422J2_124_3477_n2887), 
        .A2(n1345), .Y(DP_OP_423J2_125_3477_n2167) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1400 ( .A1(DP_OP_425J2_127_3477_n2185), 
        .A2(n1339), .Y(DP_OP_425J2_127_3477_n2161) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1395 ( .A1(DP_OP_422J2_124_3477_n2972), 
        .A2(n1339), .Y(DP_OP_424J2_126_3477_n2156) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1219 ( .A1(DP_OP_424J2_126_3477_n3058), 
        .A2(DP_OP_425J2_127_3477_n2011), .Y(DP_OP_425J2_127_3477_n1980) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1836 ( .A1(DP_OP_423J2_125_3477_n2621), 
        .A2(DP_OP_423J2_125_3477_n2627), .Y(DP_OP_423J2_125_3477_n2597) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1931 ( .A1(DP_OP_423J2_125_3477_n2708), 
        .A2(DP_OP_424J2_126_3477_n2716), .Y(DP_OP_423J2_125_3477_n2692) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1546 ( .A1(DP_OP_424J2_126_3477_n2623), 
        .A2(DP_OP_422J2_124_3477_n2321), .Y(DP_OP_422J2_124_3477_n2307) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2030 ( .A1(DP_OP_425J2_127_3477_n2799), 
        .A2(DP_OP_424J2_126_3477_n2805), .Y(DP_OP_425J2_127_3477_n2791) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1835 ( .A1(DP_OP_422J2_124_3477_n2312), 
        .A2(DP_OP_424J2_126_3477_n2627), .Y(DP_OP_424J2_126_3477_n2596) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1403 ( .A1(DP_OP_424J2_126_3477_n2268), 
        .A2(n1345), .Y(DP_OP_423J2_125_3477_n2164) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1360 ( .A1(DP_OP_422J2_124_3477_n2137), 
        .A2(DP_OP_424J2_126_3477_n2144), .Y(DP_OP_422J2_124_3477_n2121) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1936 ( .A1(DP_OP_425J2_127_3477_n2581), 
        .A2(n1341), .Y(DP_OP_422J2_124_3477_n2697) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1943 ( .A1(DP_OP_422J2_124_3477_n2712), 
        .A2(n597), .Y(DP_OP_422J2_124_3477_n2704) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1495 ( .A1(DP_OP_423J2_125_3477_n2756), 
        .A2(DP_OP_422J2_124_3477_n2276), .Y(DP_OP_422J2_124_3477_n2256) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1854 ( .A1(DP_OP_423J2_125_3477_n2315), 
        .A2(DP_OP_424J2_126_3477_n2629), .Y(DP_OP_425J2_127_3477_n2615) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2275 ( .A1(DP_OP_424J2_126_3477_n3058), 
        .A2(DP_OP_424J2_126_3477_n3065), .Y(DP_OP_424J2_126_3477_n3034) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1219 ( .A1(DP_OP_424J2_126_3477_n2004), 
        .A2(DP_OP_424J2_126_3477_n2011), .Y(DP_OP_424J2_126_3477_n1980) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2162 ( .A1(DP_OP_424J2_126_3477_n2095), 
        .A2(n445), .Y(DP_OP_425J2_127_3477_n2923) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1502 ( .A1(DP_OP_425J2_127_3477_n2403), 
        .A2(DP_OP_422J2_124_3477_n2277), .Y(DP_OP_422J2_124_3477_n2263) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1451 ( .A1(DP_OP_423J2_125_3477_n2932), 
        .A2(n365), .Y(DP_OP_425J2_127_3477_n2212) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1975 ( .A1(DP_OP_424J2_126_3477_n2268), 
        .A2(DP_OP_425J2_127_3477_n2760), .Y(DP_OP_425J2_127_3477_n2736) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2154 ( .A1(DP_OP_423J2_125_3477_n2931), 
        .A2(DP_OP_423J2_125_3477_n2936), .Y(DP_OP_423J2_125_3477_n2915) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1840 ( .A1(DP_OP_422J2_124_3477_n2625), 
        .A2(DP_OP_422J2_124_3477_n2627), .Y(DP_OP_422J2_124_3477_n2601) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1620 ( .A1(DP_OP_424J2_126_3477_n2669), 
        .A2(n799), .Y(DP_OP_425J2_127_3477_n2381) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1395 ( .A1(DP_OP_424J2_126_3477_n2268), 
        .A2(n1339), .Y(DP_OP_423J2_125_3477_n2156) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1622 ( .A1(DP_OP_423J2_125_3477_n2399), 
        .A2(n1346), .Y(DP_OP_423J2_125_3477_n2383) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1232 ( .A1(DP_OP_424J2_126_3477_n3063), 
        .A2(n558), .Y(DP_OP_425J2_127_3477_n1993) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1590 ( .A1(DP_OP_423J2_125_3477_n2667), 
        .A2(DP_OP_425J2_127_3477_n2365), .Y(DP_OP_422J2_124_3477_n2351) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1943 ( .A1(DP_OP_423J2_125_3477_n2712), 
        .A2(n597), .Y(DP_OP_423J2_125_3477_n2704) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1264 ( .A1(DP_OP_422J2_124_3477_n2049), 
        .A2(DP_OP_422J2_124_3477_n2055), .Y(DP_OP_422J2_124_3477_n2025) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2118 ( .A1(DP_OP_422J2_124_3477_n2887), 
        .A2(DP_OP_422J2_124_3477_n2893), .Y(DP_OP_422J2_124_3477_n2879) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2276 ( .A1(DP_OP_424J2_126_3477_n3059), 
        .A2(DP_OP_424J2_126_3477_n3065), .Y(DP_OP_424J2_126_3477_n3035) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1503 ( .A1(DP_OP_423J2_125_3477_n2272), 
        .A2(DP_OP_423J2_125_3477_n2277), .Y(DP_OP_423J2_125_3477_n2264) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1496 ( .A1(DP_OP_423J2_125_3477_n2273), 
        .A2(DP_OP_423J2_125_3477_n2276), .Y(DP_OP_423J2_125_3477_n2257) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1980 ( .A1(DP_OP_423J2_125_3477_n2185), 
        .A2(DP_OP_425J2_127_3477_n2760), .Y(DP_OP_425J2_127_3477_n2741) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1403 ( .A1(DP_OP_422J2_124_3477_n2972), 
        .A2(n1344), .Y(DP_OP_424J2_126_3477_n2164) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1452 ( .A1(DP_OP_423J2_125_3477_n2229), 
        .A2(n365), .Y(DP_OP_423J2_125_3477_n2213) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1224 ( .A1(DP_OP_424J2_126_3477_n2933), 
        .A2(DP_OP_422J2_124_3477_n2011), .Y(DP_OP_422J2_124_3477_n1985) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1396 ( .A1(DP_OP_422J2_124_3477_n2973), 
        .A2(n1339), .Y(DP_OP_424J2_126_3477_n2157) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1232 ( .A1(DP_OP_425J2_127_3477_n2933), 
        .A2(n558), .Y(DP_OP_423J2_125_3477_n1993) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2163 ( .A1(DP_OP_423J2_125_3477_n2008), 
        .A2(n446), .Y(DP_OP_425J2_127_3477_n2924) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2251 ( .A1(DP_OP_424J2_126_3477_n2932), 
        .A2(DP_OP_423J2_125_3477_n3025), .Y(DP_OP_423J2_125_3477_n3012) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1231 ( .A1(DP_OP_424J2_126_3477_n2932), 
        .A2(n557), .Y(DP_OP_422J2_124_3477_n1992) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1220 ( .A1(DP_OP_424J2_126_3477_n2005), 
        .A2(DP_OP_424J2_126_3477_n2011), .Y(DP_OP_424J2_126_3477_n1981) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1620 ( .A1(DP_OP_422J2_124_3477_n2405), 
        .A2(n798), .Y(DP_OP_422J2_124_3477_n2381) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2163 ( .A1(DP_OP_423J2_125_3477_n2932), 
        .A2(n446), .Y(DP_OP_423J2_125_3477_n2924) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1799 ( .A1(DP_OP_424J2_126_3477_n2576), 
        .A2(n186), .Y(DP_OP_424J2_126_3477_n2560) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1268 ( .A1(DP_OP_424J2_126_3477_n2889), 
        .A2(DP_OP_422J2_124_3477_n2055), .Y(DP_OP_422J2_124_3477_n2029) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2251 ( .A1(DP_OP_425J2_127_3477_n3020), 
        .A2(DP_OP_425J2_127_3477_n3025), .Y(DP_OP_425J2_127_3477_n3012) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2151 ( .A1(DP_OP_424J2_126_3477_n2928), 
        .A2(DP_OP_424J2_126_3477_n2936), .Y(DP_OP_424J2_126_3477_n2912) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1493 ( .A1(DP_OP_422J2_124_3477_n2798), 
        .A2(DP_OP_423J2_125_3477_n2276), .Y(DP_OP_423J2_125_3477_n2254) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2068 ( .A1(DP_OP_423J2_125_3477_n2097), 
        .A2(DP_OP_425J2_127_3477_n2848), .Y(DP_OP_425J2_127_3477_n2829) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1229 ( .A1(DP_OP_422J2_124_3477_n2006), 
        .A2(n558), .Y(DP_OP_422J2_124_3477_n1990) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2294 ( .A1(DP_OP_424J2_126_3477_n2095), 
        .A2(n693), .Y(DP_OP_422J2_124_3477_n3053) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1975 ( .A1(DP_OP_424J2_126_3477_n2752), 
        .A2(DP_OP_425J2_127_3477_n2760), .Y(DP_OP_424J2_126_3477_n2736) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1408 ( .A1(DP_OP_423J2_125_3477_n2185), 
        .A2(n1345), .Y(DP_OP_423J2_125_3477_n2169) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1853 ( .A1(DP_OP_423J2_125_3477_n2622), 
        .A2(DP_OP_423J2_125_3477_n2629), .Y(DP_OP_423J2_125_3477_n2614) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1364 ( .A1(DP_OP_425J2_127_3477_n2801), 
        .A2(DP_OP_425J2_127_3477_n2144), .Y(DP_OP_423J2_125_3477_n2125) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1931 ( .A1(DP_OP_422J2_124_3477_n2224), 
        .A2(n1340), .Y(DP_OP_424J2_126_3477_n2692) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1799 ( .A1(DP_OP_425J2_127_3477_n2576), 
        .A2(n186), .Y(DP_OP_425J2_127_3477_n2560) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1544 ( .A1(DP_OP_422J2_124_3477_n2313), 
        .A2(DP_OP_422J2_124_3477_n2321), .Y(DP_OP_422J2_124_3477_n2305) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1408 ( .A1(DP_OP_425J2_127_3477_n2185), 
        .A2(DP_OP_425J2_127_3477_n2188), .Y(DP_OP_425J2_127_3477_n2169) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1500 ( .A1(DP_OP_423J2_125_3477_n2269), 
        .A2(DP_OP_423J2_125_3477_n2277), .Y(DP_OP_423J2_125_3477_n2261) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1222 ( .A1(DP_OP_422J2_124_3477_n2007), 
        .A2(DP_OP_422J2_124_3477_n2011), .Y(DP_OP_422J2_124_3477_n1983) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2295 ( .A1(DP_OP_423J2_125_3477_n3062), 
        .A2(n692), .Y(DP_OP_423J2_125_3477_n3054) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1616 ( .A1(DP_OP_422J2_124_3477_n2753), 
        .A2(n799), .Y(DP_OP_424J2_126_3477_n2377) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2295 ( .A1(DP_OP_425J2_127_3477_n3062), 
        .A2(n33), .Y(DP_OP_425J2_127_3477_n3054) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1364 ( .A1(DP_OP_423J2_125_3477_n3021), 
        .A2(DP_OP_424J2_126_3477_n2144), .Y(DP_OP_425J2_127_3477_n2125) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1799 ( .A1(DP_OP_422J2_124_3477_n2576), 
        .A2(DP_OP_424J2_126_3477_n2584), .Y(DP_OP_422J2_124_3477_n2560) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2012 ( .A1(DP_OP_422J2_124_3477_n2137), 
        .A2(DP_OP_422J2_124_3477_n2803), .Y(DP_OP_424J2_126_3477_n2773) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1987 ( .A1(DP_OP_423J2_125_3477_n2756), 
        .A2(n66), .Y(DP_OP_423J2_125_3477_n2748) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1836 ( .A1(DP_OP_422J2_124_3477_n2313), 
        .A2(DP_OP_424J2_126_3477_n2627), .Y(DP_OP_424J2_126_3477_n2597) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1987 ( .A1(DP_OP_425J2_127_3477_n2756), 
        .A2(n66), .Y(DP_OP_425J2_127_3477_n2748) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1308 ( .A1(DP_OP_423J2_125_3477_n2005), 
        .A2(DP_OP_424J2_126_3477_n2099), .Y(DP_OP_424J2_126_3477_n2069) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1544 ( .A1(DP_OP_423J2_125_3477_n2225), 
        .A2(DP_OP_425J2_127_3477_n2321), .Y(DP_OP_424J2_126_3477_n2305) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1230 ( .A1(DP_OP_423J2_125_3477_n2007), 
        .A2(n558), .Y(DP_OP_423J2_125_3477_n1991) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2119 ( .A1(DP_OP_422J2_124_3477_n2140), 
        .A2(DP_OP_425J2_127_3477_n2893), .Y(DP_OP_423J2_125_3477_n2880) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1264 ( .A1(DP_OP_425J2_127_3477_n2049), 
        .A2(DP_OP_425J2_127_3477_n2055), .Y(DP_OP_425J2_127_3477_n2025) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2251 ( .A1(DP_OP_423J2_125_3477_n2052), 
        .A2(n846), .Y(DP_OP_422J2_124_3477_n3012) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1227 ( .A1(DP_OP_422J2_124_3477_n3058), 
        .A2(n558), .Y(DP_OP_423J2_125_3477_n1988) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2156 ( .A1(DP_OP_424J2_126_3477_n2845), 
        .A2(DP_OP_423J2_125_3477_n2936), .Y(DP_OP_423J2_125_3477_n2917) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1408 ( .A1(DP_OP_422J2_124_3477_n2185), 
        .A2(DP_OP_425J2_127_3477_n2188), .Y(DP_OP_422J2_124_3477_n2169) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1227 ( .A1(DP_OP_424J2_126_3477_n2004), 
        .A2(n558), .Y(DP_OP_424J2_126_3477_n1988) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1223 ( .A1(DP_OP_423J2_125_3477_n2008), 
        .A2(DP_OP_425J2_127_3477_n2011), .Y(DP_OP_423J2_125_3477_n1984) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1933 ( .A1(DP_OP_422J2_124_3477_n2710), 
        .A2(n1341), .Y(DP_OP_422J2_124_3477_n2694) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2153 ( .A1(DP_OP_422J2_124_3477_n2006), 
        .A2(DP_OP_424J2_126_3477_n2936), .Y(DP_OP_424J2_126_3477_n2914) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1405 ( .A1(DP_OP_424J2_126_3477_n2754), 
        .A2(n1343), .Y(DP_OP_422J2_124_3477_n2166) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2250 ( .A1(DP_OP_422J2_124_3477_n3019), 
        .A2(DP_OP_423J2_125_3477_n3025), .Y(DP_OP_422J2_124_3477_n3011) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1936 ( .A1(DP_OP_423J2_125_3477_n2713), 
        .A2(n1341), .Y(DP_OP_423J2_125_3477_n2697) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1838 ( .A1(DP_OP_423J2_125_3477_n2623), 
        .A2(DP_OP_423J2_125_3477_n2627), .Y(DP_OP_423J2_125_3477_n2599) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1679 ( .A1(DP_OP_425J2_127_3477_n2448), 
        .A2(DP_OP_425J2_127_3477_n2453), .Y(DP_OP_425J2_127_3477_n2440) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1986 ( .A1(DP_OP_424J2_126_3477_n2403), 
        .A2(n66), .Y(DP_OP_422J2_124_3477_n2747) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1615 ( .A1(DP_OP_423J2_125_3477_n2400), 
        .A2(n799), .Y(DP_OP_423J2_125_3477_n2376) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1491 ( .A1(DP_OP_424J2_126_3477_n2268), 
        .A2(DP_OP_424J2_126_3477_n2276), .Y(DP_OP_424J2_126_3477_n2252) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1267 ( .A1(DP_OP_423J2_125_3477_n2052), 
        .A2(DP_OP_425J2_127_3477_n2055), .Y(DP_OP_423J2_125_3477_n2028) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1804 ( .A1(DP_OP_423J2_125_3477_n2581), 
        .A2(n186), .Y(DP_OP_423J2_125_3477_n2565) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1498 ( .A1(DP_OP_424J2_126_3477_n2267), 
        .A2(DP_OP_424J2_126_3477_n2277), .Y(DP_OP_424J2_126_3477_n2259) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2160 ( .A1(DP_OP_424J2_126_3477_n2929), 
        .A2(n446), .Y(DP_OP_424J2_126_3477_n2921) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1263 ( .A1(DP_OP_423J2_125_3477_n2048), 
        .A2(DP_OP_422J2_124_3477_n2055), .Y(DP_OP_423J2_125_3477_n2024) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1935 ( .A1(DP_OP_422J2_124_3477_n2712), 
        .A2(DP_OP_424J2_126_3477_n2716), .Y(DP_OP_422J2_124_3477_n2696) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1628 ( .A1(DP_OP_423J2_125_3477_n2405), 
        .A2(DP_OP_424J2_126_3477_n2408), .Y(DP_OP_423J2_125_3477_n2389) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1447 ( .A1(DP_OP_422J2_124_3477_n2928), 
        .A2(n365), .Y(DP_OP_424J2_126_3477_n2208) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1238 ( .A1(DP_OP_422J2_124_3477_n2007), 
        .A2(DP_OP_422J2_124_3477_n2013), .Y(DP_OP_422J2_124_3477_n1999) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1173 ( .A1(n1867), .A2(n1508), .Y(
        DP_OP_422J2_124_3477_n1934) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1659 ( .A1(DP_OP_422J2_124_3477_n2444), 
        .A2(n789), .Y(DP_OP_422J2_124_3477_n2420) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1763 ( .A1(DP_OP_422J2_124_3477_n2532), 
        .A2(DP_OP_422J2_124_3477_n2541), .Y(DP_OP_422J2_124_3477_n2524) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1272 ( .A1(DP_OP_425J2_127_3477_n2885), 
        .A2(DP_OP_424J2_126_3477_n2056), .Y(DP_OP_423J2_125_3477_n2033) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2145 ( .A1(DP_OP_422J2_124_3477_n2930), 
        .A2(DP_OP_425J2_127_3477_n2935), .Y(DP_OP_422J2_124_3477_n2906) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1274 ( .A1(DP_OP_424J2_126_3477_n2051), 
        .A2(DP_OP_424J2_126_3477_n2056), .Y(DP_OP_424J2_126_3477_n2035) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1767 ( .A1(DP_OP_422J2_124_3477_n2404), 
        .A2(DP_OP_424J2_126_3477_n2541), .Y(DP_OP_424J2_126_3477_n2528) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1881 ( .A1(DP_OP_423J2_125_3477_n2666), 
        .A2(DP_OP_424J2_126_3477_n2671), .Y(DP_OP_423J2_125_3477_n2642) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1663 ( .A1(DP_OP_425J2_127_3477_n2448), 
        .A2(n789), .Y(DP_OP_425J2_127_3477_n2424) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2208 ( .A1(DP_OP_425J2_127_3477_n2977), 
        .A2(n677), .Y(DP_OP_425J2_127_3477_n2969) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1483 ( .A1(DP_OP_422J2_124_3477_n2268), 
        .A2(DP_OP_422J2_124_3477_n2275), .Y(DP_OP_422J2_124_3477_n2244) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1485 ( .A1(DP_OP_422J2_124_3477_n2270), 
        .A2(DP_OP_424J2_126_3477_n2275), .Y(DP_OP_422J2_124_3477_n2246) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2205 ( .A1(DP_OP_424J2_126_3477_n2974), 
        .A2(n676), .Y(DP_OP_424J2_126_3477_n2966) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2143 ( .A1(DP_OP_422J2_124_3477_n2928), 
        .A2(DP_OP_425J2_127_3477_n2935), .Y(DP_OP_422J2_124_3477_n2904) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1488 ( .A1(DP_OP_423J2_125_3477_n2185), 
        .A2(DP_OP_422J2_124_3477_n2275), .Y(DP_OP_424J2_126_3477_n2249) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1661 ( .A1(DP_OP_422J2_124_3477_n2446), 
        .A2(n789), .Y(DP_OP_422J2_124_3477_n2422) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1411 ( .A1(DP_OP_424J2_126_3477_n2752), 
        .A2(DP_OP_422J2_124_3477_n2189), .Y(DP_OP_422J2_124_3477_n2172) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2073 ( .A1(DP_OP_422J2_124_3477_n2842), 
        .A2(DP_OP_424J2_126_3477_n2849), .Y(DP_OP_422J2_124_3477_n2834) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1275 ( .A1(DP_OP_425J2_127_3477_n2976), 
        .A2(DP_OP_424J2_126_3477_n2056), .Y(DP_OP_424J2_126_3477_n2036) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1414 ( .A1(DP_OP_422J2_124_3477_n2975), 
        .A2(DP_OP_424J2_126_3477_n2189), .Y(DP_OP_424J2_126_3477_n2175) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2243 ( .A1(DP_OP_424J2_126_3477_n3020), 
        .A2(n704), .Y(DP_OP_424J2_126_3477_n3004) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2101 ( .A1(DP_OP_423J2_125_3477_n2182), 
        .A2(DP_OP_423J2_125_3477_n2891), .Y(DP_OP_422J2_124_3477_n2862) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1766 ( .A1(DP_OP_424J2_126_3477_n2535), 
        .A2(DP_OP_424J2_126_3477_n2541), .Y(DP_OP_424J2_126_3477_n2527) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1151 ( .A1(n1296), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_423J2_125_3477_n314) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1971 ( .A1(DP_OP_422J2_124_3477_n2756), 
        .A2(DP_OP_422J2_124_3477_n2759), .Y(DP_OP_422J2_124_3477_n2732) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2206 ( .A1(DP_OP_424J2_126_3477_n2975), 
        .A2(n676), .Y(DP_OP_424J2_126_3477_n2967) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2195 ( .A1(DP_OP_422J2_124_3477_n2972), 
        .A2(DP_OP_425J2_127_3477_n2980), .Y(DP_OP_422J2_124_3477_n2956) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1967 ( .A1(DP_OP_424J2_126_3477_n2400), 
        .A2(DP_OP_422J2_124_3477_n2759), .Y(DP_OP_422J2_124_3477_n2728) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1703 ( .A1(DP_OP_422J2_124_3477_n2488), 
        .A2(DP_OP_422J2_124_3477_n2495), .Y(DP_OP_422J2_124_3477_n2464) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1171 ( .A1(n1287), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_423J2_125_3477_n1932) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1571 ( .A1(DP_OP_422J2_124_3477_n2356), 
        .A2(n874), .Y(DP_OP_422J2_124_3477_n2332) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2074 ( .A1(DP_OP_423J2_125_3477_n2931), 
        .A2(DP_OP_424J2_126_3477_n2849), .Y(DP_OP_424J2_126_3477_n2835) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1573 ( .A1(DP_OP_422J2_124_3477_n2710), 
        .A2(n874), .Y(DP_OP_423J2_125_3477_n2334) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1157 ( .A1(n1892), .A2(n1508), .Y(
        DP_OP_424J2_126_3477_n326) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1707 ( .A1(DP_OP_423J2_125_3477_n2536), 
        .A2(DP_OP_422J2_124_3477_n2495), .Y(DP_OP_422J2_124_3477_n2468) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1239 ( .A1(DP_OP_425J2_127_3477_n3020), 
        .A2(DP_OP_423J2_125_3477_n2013), .Y(DP_OP_424J2_126_3477_n2000) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1721 ( .A1(DP_OP_422J2_124_3477_n2490), 
        .A2(DP_OP_425J2_127_3477_n2497), .Y(DP_OP_422J2_124_3477_n2482) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2104 ( .A1(DP_OP_424J2_126_3477_n2889), 
        .A2(DP_OP_425J2_127_3477_n2891), .Y(DP_OP_424J2_126_3477_n2865) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1722 ( .A1(DP_OP_424J2_126_3477_n2491), 
        .A2(DP_OP_422J2_124_3477_n2497), .Y(DP_OP_424J2_126_3477_n2483) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1576 ( .A1(DP_OP_423J2_125_3477_n2361), 
        .A2(n876), .Y(DP_OP_423J2_125_3477_n2337) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2111 ( .A1(DP_OP_423J2_125_3477_n2976), 
        .A2(DP_OP_423J2_125_3477_n2892), .Y(DP_OP_424J2_126_3477_n2872) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1719 ( .A1(DP_OP_422J2_124_3477_n2488), 
        .A2(DP_OP_424J2_126_3477_n2497), .Y(DP_OP_422J2_124_3477_n2480) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1274 ( .A1(DP_OP_423J2_125_3477_n2051), 
        .A2(DP_OP_425J2_127_3477_n2056), .Y(DP_OP_423J2_125_3477_n2035) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2199 ( .A1(DP_OP_424J2_126_3477_n2976), 
        .A2(DP_OP_424J2_126_3477_n2980), .Y(DP_OP_424J2_126_3477_n2960) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1576 ( .A1(DP_OP_423J2_125_3477_n2273), 
        .A2(n875), .Y(DP_OP_424J2_126_3477_n2337) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1235 ( .A1(DP_OP_422J2_124_3477_n2004), 
        .A2(DP_OP_423J2_125_3477_n2013), .Y(DP_OP_422J2_124_3477_n1996) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2241 ( .A1(DP_OP_425J2_127_3477_n2138), 
        .A2(n704), .Y(DP_OP_423J2_125_3477_n3002) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1415 ( .A1(DP_OP_424J2_126_3477_n2756), 
        .A2(DP_OP_422J2_124_3477_n2189), .Y(DP_OP_422J2_124_3477_n2176) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1706 ( .A1(DP_OP_422J2_124_3477_n2579), 
        .A2(DP_OP_422J2_124_3477_n2495), .Y(DP_OP_423J2_125_3477_n2467) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1273 ( .A1(DP_OP_425J2_127_3477_n2886), 
        .A2(DP_OP_424J2_126_3477_n2056), .Y(DP_OP_423J2_125_3477_n2034) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2071 ( .A1(DP_OP_422J2_124_3477_n2092), 
        .A2(DP_OP_423J2_125_3477_n2849), .Y(DP_OP_424J2_126_3477_n2832) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2195 ( .A1(DP_OP_424J2_126_3477_n2972), 
        .A2(DP_OP_425J2_127_3477_n2980), .Y(DP_OP_424J2_126_3477_n2956) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1767 ( .A1(DP_OP_423J2_125_3477_n2536), 
        .A2(DP_OP_422J2_124_3477_n2541), .Y(DP_OP_423J2_125_3477_n2528) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2239 ( .A1(DP_OP_425J2_127_3477_n2048), 
        .A2(n704), .Y(DP_OP_424J2_126_3477_n3000) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1410 ( .A1(DP_OP_422J2_124_3477_n2971), 
        .A2(DP_OP_424J2_126_3477_n2189), .Y(DP_OP_424J2_126_3477_n2171) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1459 ( .A1(DP_OP_423J2_125_3477_n2228), 
        .A2(DP_OP_423J2_125_3477_n2233), .Y(DP_OP_423J2_125_3477_n2220) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1411 ( .A1(DP_OP_422J2_124_3477_n2972), 
        .A2(DP_OP_424J2_126_3477_n2189), .Y(DP_OP_424J2_126_3477_n2172) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2107 ( .A1(DP_OP_425J2_127_3477_n2180), 
        .A2(DP_OP_423J2_125_3477_n2892), .Y(DP_OP_424J2_126_3477_n2868) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1271 ( .A1(DP_OP_425J2_127_3477_n2972), 
        .A2(DP_OP_424J2_126_3477_n2056), .Y(DP_OP_424J2_126_3477_n2032) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2244 ( .A1(DP_OP_423J2_125_3477_n3021), 
        .A2(n704), .Y(DP_OP_423J2_125_3477_n3005) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1271 ( .A1(DP_OP_422J2_124_3477_n2048), 
        .A2(DP_OP_422J2_124_3477_n2056), .Y(DP_OP_422J2_124_3477_n2032) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1765 ( .A1(DP_OP_422J2_124_3477_n2490), 
        .A2(DP_OP_424J2_126_3477_n2541), .Y(DP_OP_423J2_125_3477_n2526) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1484 ( .A1(DP_OP_424J2_126_3477_n2269), 
        .A2(DP_OP_422J2_124_3477_n2275), .Y(DP_OP_424J2_126_3477_n2245) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1719 ( .A1(DP_OP_422J2_124_3477_n2664), 
        .A2(DP_OP_424J2_126_3477_n2497), .Y(DP_OP_424J2_126_3477_n2480) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1762 ( .A1(DP_OP_422J2_124_3477_n2399), 
        .A2(DP_OP_424J2_126_3477_n2541), .Y(DP_OP_424J2_126_3477_n2523) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2144 ( .A1(DP_OP_422J2_124_3477_n2929), 
        .A2(DP_OP_422J2_124_3477_n2935), .Y(DP_OP_422J2_124_3477_n2905) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1768 ( .A1(DP_OP_422J2_124_3477_n2537), 
        .A2(DP_OP_422J2_124_3477_n2541), .Y(DP_OP_422J2_124_3477_n2529) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1276 ( .A1(DP_OP_423J2_125_3477_n2053), 
        .A2(DP_OP_425J2_127_3477_n2056), .Y(DP_OP_423J2_125_3477_n2037) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1455 ( .A1(DP_OP_422J2_124_3477_n2928), 
        .A2(DP_OP_423J2_125_3477_n2233), .Y(DP_OP_424J2_126_3477_n2216) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1724 ( .A1(DP_OP_423J2_125_3477_n2537), 
        .A2(DP_OP_424J2_126_3477_n2497), .Y(DP_OP_422J2_124_3477_n2485) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1412 ( .A1(DP_OP_422J2_124_3477_n2973), 
        .A2(DP_OP_424J2_126_3477_n2189), .Y(DP_OP_424J2_126_3477_n2173) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2072 ( .A1(DP_OP_422J2_124_3477_n2093), 
        .A2(DP_OP_423J2_125_3477_n2849), .Y(DP_OP_424J2_126_3477_n2833) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1574 ( .A1(DP_OP_423J2_125_3477_n2271), 
        .A2(n874), .Y(DP_OP_424J2_126_3477_n2335) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2112 ( .A1(DP_OP_423J2_125_3477_n2889), 
        .A2(DP_OP_423J2_125_3477_n2892), .Y(DP_OP_423J2_125_3477_n2873) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1485 ( .A1(DP_OP_425J2_127_3477_n2754), 
        .A2(n1427), .Y(DP_OP_424J2_126_3477_n2246) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1570 ( .A1(DP_OP_424J2_126_3477_n2443), 
        .A2(n876), .Y(DP_OP_423J2_125_3477_n2331) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1530 ( .A1(DP_OP_424J2_126_3477_n2315), 
        .A2(DP_OP_425J2_127_3477_n2319), .Y(DP_OP_424J2_126_3477_n2291) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1768 ( .A1(DP_OP_423J2_125_3477_n2537), 
        .A2(DP_OP_422J2_124_3477_n2541), .Y(DP_OP_423J2_125_3477_n2529) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1763 ( .A1(DP_OP_424J2_126_3477_n2532), 
        .A2(DP_OP_424J2_126_3477_n2541), .Y(DP_OP_424J2_126_3477_n2524) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1720 ( .A1(DP_OP_423J2_125_3477_n2401), 
        .A2(DP_OP_424J2_126_3477_n2497), .Y(DP_OP_424J2_126_3477_n2481) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2203 ( .A1(DP_OP_424J2_126_3477_n2972), 
        .A2(DP_OP_425J2_127_3477_n2981), .Y(DP_OP_424J2_126_3477_n2964) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2099 ( .A1(DP_OP_422J2_124_3477_n2048), 
        .A2(DP_OP_424J2_126_3477_n2891), .Y(DP_OP_424J2_126_3477_n2860) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2242 ( .A1(DP_OP_423J2_125_3477_n3019), 
        .A2(n704), .Y(DP_OP_423J2_125_3477_n3003) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2106 ( .A1(DP_OP_424J2_126_3477_n2883), 
        .A2(DP_OP_423J2_125_3477_n2892), .Y(DP_OP_424J2_126_3477_n2867) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2075 ( .A1(DP_OP_425J2_127_3477_n2712), 
        .A2(n1428), .Y(DP_OP_422J2_124_3477_n2836) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2194 ( .A1(DP_OP_424J2_126_3477_n2971), 
        .A2(DP_OP_422J2_124_3477_n2980), .Y(DP_OP_424J2_126_3477_n2955) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1456 ( .A1(DP_OP_423J2_125_3477_n2225), 
        .A2(DP_OP_423J2_125_3477_n2233), .Y(DP_OP_423J2_125_3477_n2217) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1173 ( .A1(n1866), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_423J2_125_3477_n1934) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1764 ( .A1(DP_OP_422J2_124_3477_n2489), 
        .A2(DP_OP_425J2_127_3477_n2541), .Y(DP_OP_423J2_125_3477_n2525) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1276 ( .A1(DP_OP_424J2_126_3477_n2889), 
        .A2(DP_OP_422J2_124_3477_n2056), .Y(DP_OP_422J2_124_3477_n2037) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1658 ( .A1(DP_OP_422J2_124_3477_n2443), 
        .A2(n789), .Y(DP_OP_422J2_124_3477_n2419) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1723 ( .A1(DP_OP_423J2_125_3477_n2536), 
        .A2(DP_OP_424J2_126_3477_n2497), .Y(DP_OP_422J2_124_3477_n2484) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1457 ( .A1(DP_OP_425J2_127_3477_n2710), 
        .A2(DP_OP_423J2_125_3477_n2233), .Y(DP_OP_423J2_125_3477_n2218) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1482 ( .A1(DP_OP_422J2_124_3477_n2267), 
        .A2(DP_OP_422J2_124_3477_n2275), .Y(DP_OP_422J2_124_3477_n2243) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2108 ( .A1(DP_OP_423J2_125_3477_n2973), 
        .A2(DP_OP_423J2_125_3477_n2892), .Y(DP_OP_424J2_126_3477_n2869) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2101 ( .A1(DP_OP_424J2_126_3477_n2886), 
        .A2(DP_OP_424J2_126_3477_n2891), .Y(DP_OP_424J2_126_3477_n2862) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2207 ( .A1(DP_OP_424J2_126_3477_n2184), 
        .A2(n677), .Y(DP_OP_422J2_124_3477_n2968) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2100 ( .A1(DP_OP_422J2_124_3477_n2885), 
        .A2(DP_OP_423J2_125_3477_n2891), .Y(DP_OP_422J2_124_3477_n2861) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1487 ( .A1(DP_OP_425J2_127_3477_n2756), 
        .A2(n1427), .Y(DP_OP_424J2_126_3477_n2248) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2147 ( .A1(DP_OP_424J2_126_3477_n2932), 
        .A2(n1432), .Y(DP_OP_424J2_126_3477_n2908) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1765 ( .A1(DP_OP_424J2_126_3477_n2534), 
        .A2(DP_OP_424J2_126_3477_n2541), .Y(DP_OP_424J2_126_3477_n2526) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2110 ( .A1(DP_OP_424J2_126_3477_n2887), 
        .A2(DP_OP_423J2_125_3477_n2892), .Y(DP_OP_424J2_126_3477_n2871) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1413 ( .A1(DP_OP_422J2_124_3477_n2974), 
        .A2(DP_OP_424J2_126_3477_n2189), .Y(DP_OP_424J2_126_3477_n2174) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1238 ( .A1(DP_OP_425J2_127_3477_n3019), 
        .A2(DP_OP_422J2_124_3477_n2013), .Y(DP_OP_424J2_126_3477_n1999) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2104 ( .A1(DP_OP_422J2_124_3477_n2889), 
        .A2(DP_OP_424J2_126_3477_n2891), .Y(DP_OP_422J2_124_3477_n2865) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2242 ( .A1(DP_OP_424J2_126_3477_n3019), 
        .A2(n704), .Y(DP_OP_424J2_126_3477_n3003) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1721 ( .A1(DP_OP_425J2_127_3477_n2534), 
        .A2(DP_OP_424J2_126_3477_n2497), .Y(DP_OP_424J2_126_3477_n2482) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1275 ( .A1(DP_OP_423J2_125_3477_n2052), 
        .A2(DP_OP_424J2_126_3477_n2056), .Y(DP_OP_423J2_125_3477_n2036) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2198 ( .A1(DP_OP_424J2_126_3477_n2975), 
        .A2(DP_OP_422J2_124_3477_n2980), .Y(DP_OP_424J2_126_3477_n2959) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2240 ( .A1(DP_OP_424J2_126_3477_n2929), 
        .A2(n704), .Y(DP_OP_423J2_125_3477_n3001) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1272 ( .A1(DP_OP_422J2_124_3477_n2049), 
        .A2(DP_OP_422J2_124_3477_n2056), .Y(DP_OP_422J2_124_3477_n2033) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2073 ( .A1(DP_OP_425J2_127_3477_n2226), 
        .A2(DP_OP_424J2_126_3477_n2849), .Y(DP_OP_424J2_126_3477_n2834) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1484 ( .A1(DP_OP_422J2_124_3477_n2269), 
        .A2(n1427), .Y(DP_OP_422J2_124_3477_n2245) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2196 ( .A1(DP_OP_424J2_126_3477_n2973), 
        .A2(DP_OP_425J2_127_3477_n2980), .Y(DP_OP_424J2_126_3477_n2957) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1272 ( .A1(DP_OP_425J2_127_3477_n2973), 
        .A2(DP_OP_424J2_126_3477_n2056), .Y(DP_OP_424J2_126_3477_n2033) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1460 ( .A1(DP_OP_423J2_125_3477_n2229), 
        .A2(DP_OP_423J2_125_3477_n2233), .Y(DP_OP_423J2_125_3477_n2221) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1273 ( .A1(DP_OP_425J2_127_3477_n2974), 
        .A2(DP_OP_424J2_126_3477_n2056), .Y(DP_OP_424J2_126_3477_n2034) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1764 ( .A1(DP_OP_422J2_124_3477_n2401), 
        .A2(DP_OP_424J2_126_3477_n2541), .Y(DP_OP_424J2_126_3477_n2525) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1486 ( .A1(DP_OP_425J2_127_3477_n2755), 
        .A2(DP_OP_422J2_124_3477_n2275), .Y(DP_OP_424J2_126_3477_n2247) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1456 ( .A1(DP_OP_422J2_124_3477_n2929), 
        .A2(DP_OP_423J2_125_3477_n2233), .Y(DP_OP_424J2_126_3477_n2217) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2240 ( .A1(DP_OP_425J2_127_3477_n2049), 
        .A2(n703), .Y(DP_OP_424J2_126_3477_n3001) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2197 ( .A1(DP_OP_424J2_126_3477_n2974), 
        .A2(DP_OP_425J2_127_3477_n2980), .Y(DP_OP_424J2_126_3477_n2958) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2204 ( .A1(DP_OP_424J2_126_3477_n2973), 
        .A2(n677), .Y(DP_OP_424J2_126_3477_n2965) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2241 ( .A1(DP_OP_425J2_127_3477_n2050), 
        .A2(DP_OP_425J2_127_3477_n3024), .Y(DP_OP_424J2_126_3477_n3002) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2102 ( .A1(DP_OP_424J2_126_3477_n2887), 
        .A2(DP_OP_423J2_125_3477_n2891), .Y(DP_OP_424J2_126_3477_n2863) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2109 ( .A1(DP_OP_424J2_126_3477_n2886), 
        .A2(DP_OP_423J2_125_3477_n2892), .Y(DP_OP_424J2_126_3477_n2870) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1416 ( .A1(DP_OP_422J2_124_3477_n2185), 
        .A2(DP_OP_422J2_124_3477_n2189), .Y(DP_OP_422J2_124_3477_n2177) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1767 ( .A1(DP_OP_422J2_124_3477_n2536), 
        .A2(DP_OP_422J2_124_3477_n2541), .Y(DP_OP_422J2_124_3477_n2528) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1240 ( .A1(DP_OP_424J2_126_3477_n2933), 
        .A2(DP_OP_423J2_125_3477_n2013), .Y(DP_OP_422J2_124_3477_n2001) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2208 ( .A1(DP_OP_424J2_126_3477_n2185), 
        .A2(n677), .Y(DP_OP_422J2_124_3477_n2969) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1708 ( .A1(DP_OP_423J2_125_3477_n2493), 
        .A2(DP_OP_425J2_127_3477_n2495), .Y(DP_OP_423J2_125_3477_n2469) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1458 ( .A1(DP_OP_423J2_125_3477_n2227), 
        .A2(DP_OP_423J2_125_3477_n2233), .Y(DP_OP_423J2_125_3477_n2219) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2100 ( .A1(DP_OP_423J2_125_3477_n2973), 
        .A2(DP_OP_424J2_126_3477_n2891), .Y(DP_OP_424J2_126_3477_n2861) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1762 ( .A1(DP_OP_422J2_124_3477_n2531), 
        .A2(DP_OP_422J2_124_3477_n2541), .Y(DP_OP_422J2_124_3477_n2523) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1723 ( .A1(DP_OP_424J2_126_3477_n2580), 
        .A2(DP_OP_424J2_126_3477_n2497), .Y(DP_OP_425J2_127_3477_n2484) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1574 ( .A1(DP_OP_424J2_126_3477_n2579), 
        .A2(n874), .Y(DP_OP_422J2_124_3477_n2335) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2102 ( .A1(DP_OP_422J2_124_3477_n2887), 
        .A2(DP_OP_425J2_127_3477_n2891), .Y(DP_OP_422J2_124_3477_n2863) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1720 ( .A1(DP_OP_423J2_125_3477_n2665), 
        .A2(DP_OP_425J2_127_3477_n2497), .Y(DP_OP_425J2_127_3477_n2481) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2207 ( .A1(DP_OP_425J2_127_3477_n2976), 
        .A2(n677), .Y(DP_OP_425J2_127_3477_n2968) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2200 ( .A1(DP_OP_425J2_127_3477_n2977), 
        .A2(DP_OP_422J2_124_3477_n2980), .Y(DP_OP_425J2_127_3477_n2961) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1271 ( .A1(DP_OP_423J2_125_3477_n2048), 
        .A2(DP_OP_425J2_127_3477_n2056), .Y(DP_OP_423J2_125_3477_n2032) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1415 ( .A1(DP_OP_425J2_127_3477_n2184), 
        .A2(DP_OP_425J2_127_3477_n2189), .Y(DP_OP_425J2_127_3477_n2176) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2244 ( .A1(DP_OP_425J2_127_3477_n3021), 
        .A2(n704), .Y(DP_OP_425J2_127_3477_n3005) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1273 ( .A1(DP_OP_425J2_127_3477_n2050), 
        .A2(DP_OP_425J2_127_3477_n2056), .Y(DP_OP_425J2_127_3477_n2034) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2074 ( .A1(DP_OP_423J2_125_3477_n2227), 
        .A2(DP_OP_424J2_126_3477_n2849), .Y(DP_OP_422J2_124_3477_n2835) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2108 ( .A1(DP_OP_425J2_127_3477_n2885), 
        .A2(DP_OP_423J2_125_3477_n2892), .Y(DP_OP_425J2_127_3477_n2869) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2101 ( .A1(DP_OP_425J2_127_3477_n2886), 
        .A2(DP_OP_425J2_127_3477_n2891), .Y(DP_OP_425J2_127_3477_n2862) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1486 ( .A1(DP_OP_424J2_126_3477_n2667), 
        .A2(n1427), .Y(DP_OP_422J2_124_3477_n2247) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1764 ( .A1(DP_OP_422J2_124_3477_n2665), 
        .A2(DP_OP_425J2_127_3477_n2541), .Y(DP_OP_425J2_127_3477_n2525) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2206 ( .A1(DP_OP_422J2_124_3477_n2975), 
        .A2(n676), .Y(DP_OP_422J2_124_3477_n2967) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1766 ( .A1(DP_OP_422J2_124_3477_n2535), 
        .A2(DP_OP_422J2_124_3477_n2541), .Y(DP_OP_422J2_124_3477_n2527) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2243 ( .A1(DP_OP_425J2_127_3477_n2888), 
        .A2(n703), .Y(DP_OP_422J2_124_3477_n3004) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2071 ( .A1(DP_OP_425J2_127_3477_n2840), 
        .A2(n1428), .Y(DP_OP_425J2_127_3477_n2832) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1486 ( .A1(DP_OP_424J2_126_3477_n2799), 
        .A2(DP_OP_422J2_124_3477_n2275), .Y(DP_OP_425J2_127_3477_n2247) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2197 ( .A1(DP_OP_425J2_127_3477_n2974), 
        .A2(DP_OP_422J2_124_3477_n2980), .Y(DP_OP_425J2_127_3477_n2958) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2204 ( .A1(DP_OP_425J2_127_3477_n2973), 
        .A2(n677), .Y(DP_OP_425J2_127_3477_n2965) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1414 ( .A1(DP_OP_422J2_124_3477_n2183), 
        .A2(DP_OP_422J2_124_3477_n2189), .Y(DP_OP_422J2_124_3477_n2175) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2241 ( .A1(DP_OP_424J2_126_3477_n2006), 
        .A2(n704), .Y(DP_OP_425J2_127_3477_n3002) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1411 ( .A1(DP_OP_425J2_127_3477_n2180), 
        .A2(DP_OP_425J2_127_3477_n2189), .Y(DP_OP_425J2_127_3477_n2172) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1881 ( .A1(DP_OP_424J2_126_3477_n2358), 
        .A2(DP_OP_425J2_127_3477_n2671), .Y(DP_OP_425J2_127_3477_n2642) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1275 ( .A1(DP_OP_425J2_127_3477_n2184), 
        .A2(DP_OP_422J2_124_3477_n2056), .Y(DP_OP_422J2_124_3477_n2036) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1661 ( .A1(DP_OP_424J2_126_3477_n2622), 
        .A2(n789), .Y(DP_OP_425J2_127_3477_n2422) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2102 ( .A1(DP_OP_423J2_125_3477_n2051), 
        .A2(DP_OP_424J2_126_3477_n2891), .Y(DP_OP_425J2_127_3477_n2863) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1153 ( .A1(n1309), .A2(n1508), .Y(
        DP_OP_425J2_127_3477_n318) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2109 ( .A1(DP_OP_425J2_127_3477_n2886), 
        .A2(DP_OP_423J2_125_3477_n2892), .Y(DP_OP_425J2_127_3477_n2870) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2146 ( .A1(DP_OP_425J2_127_3477_n2799), 
        .A2(n1432), .Y(DP_OP_422J2_124_3477_n2907) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1662 ( .A1(DP_OP_425J2_127_3477_n2447), 
        .A2(n789), .Y(DP_OP_425J2_127_3477_n2423) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1155 ( .A1(n1310), .A2(n1508), .Y(
        DP_OP_425J2_127_3477_n322) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1764 ( .A1(DP_OP_422J2_124_3477_n2533), 
        .A2(DP_OP_422J2_124_3477_n2541), .Y(DP_OP_422J2_124_3477_n2525) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1719 ( .A1(DP_OP_424J2_126_3477_n2576), 
        .A2(DP_OP_422J2_124_3477_n2497), .Y(DP_OP_425J2_127_3477_n2480) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1660 ( .A1(DP_OP_425J2_127_3477_n2445), 
        .A2(n789), .Y(DP_OP_425J2_127_3477_n2421) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1721 ( .A1(DP_OP_422J2_124_3477_n2358), 
        .A2(DP_OP_422J2_124_3477_n2497), .Y(DP_OP_425J2_127_3477_n2482) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1527 ( .A1(DP_OP_425J2_127_3477_n2312), 
        .A2(DP_OP_425J2_127_3477_n2319), .Y(DP_OP_425J2_127_3477_n2288) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1724 ( .A1(DP_OP_425J2_127_3477_n2493), 
        .A2(DP_OP_425J2_127_3477_n2497), .Y(DP_OP_425J2_127_3477_n2485) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1768 ( .A1(DP_OP_422J2_124_3477_n2669), 
        .A2(DP_OP_425J2_127_3477_n2541), .Y(DP_OP_425J2_127_3477_n2529) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1238 ( .A1(DP_OP_425J2_127_3477_n2007), 
        .A2(n1431), .Y(DP_OP_425J2_127_3477_n1999) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2075 ( .A1(DP_OP_423J2_125_3477_n2096), 
        .A2(n1428), .Y(DP_OP_425J2_127_3477_n2836) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1967 ( .A1(DP_OP_424J2_126_3477_n2268), 
        .A2(DP_OP_422J2_124_3477_n2759), .Y(DP_OP_425J2_127_3477_n2728) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1659 ( .A1(DP_OP_423J2_125_3477_n2708), 
        .A2(n789), .Y(DP_OP_425J2_127_3477_n2420) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1483 ( .A1(DP_OP_425J2_127_3477_n2268), 
        .A2(n1427), .Y(DP_OP_425J2_127_3477_n2244) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1412 ( .A1(DP_OP_423J2_125_3477_n2973), 
        .A2(DP_OP_425J2_127_3477_n2189), .Y(DP_OP_425J2_127_3477_n2173) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1708 ( .A1(DP_OP_423J2_125_3477_n2537), 
        .A2(DP_OP_422J2_124_3477_n2495), .Y(DP_OP_422J2_124_3477_n2469) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2072 ( .A1(DP_OP_425J2_127_3477_n2841), 
        .A2(DP_OP_423J2_125_3477_n2849), .Y(DP_OP_425J2_127_3477_n2833) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1972 ( .A1(DP_OP_424J2_126_3477_n2405), 
        .A2(DP_OP_422J2_124_3477_n2759), .Y(DP_OP_422J2_124_3477_n2733) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2106 ( .A1(DP_OP_425J2_127_3477_n2883), 
        .A2(DP_OP_423J2_125_3477_n2892), .Y(DP_OP_425J2_127_3477_n2867) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2146 ( .A1(DP_OP_424J2_126_3477_n2095), 
        .A2(n1432), .Y(DP_OP_425J2_127_3477_n2907) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1662 ( .A1(DP_OP_423J2_125_3477_n2579), 
        .A2(n789), .Y(DP_OP_422J2_124_3477_n2423) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2194 ( .A1(DP_OP_425J2_127_3477_n2971), 
        .A2(DP_OP_425J2_127_3477_n2980), .Y(DP_OP_425J2_127_3477_n2955) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1488 ( .A1(DP_OP_424J2_126_3477_n2669), 
        .A2(n1427), .Y(DP_OP_422J2_124_3477_n2249) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1530 ( .A1(DP_OP_423J2_125_3477_n2843), 
        .A2(DP_OP_425J2_127_3477_n2319), .Y(DP_OP_425J2_127_3477_n2291) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1412 ( .A1(DP_OP_422J2_124_3477_n2181), 
        .A2(DP_OP_422J2_124_3477_n2189), .Y(DP_OP_422J2_124_3477_n2173) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1722 ( .A1(DP_OP_422J2_124_3477_n2491), 
        .A2(DP_OP_425J2_127_3477_n2497), .Y(DP_OP_422J2_124_3477_n2483) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1276 ( .A1(DP_OP_425J2_127_3477_n2053), 
        .A2(DP_OP_425J2_127_3477_n2056), .Y(DP_OP_425J2_127_3477_n2037) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1766 ( .A1(DP_OP_422J2_124_3477_n2667), 
        .A2(DP_OP_425J2_127_3477_n2541), .Y(DP_OP_425J2_127_3477_n2527) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2243 ( .A1(DP_OP_425J2_127_3477_n3020), 
        .A2(n703), .Y(DP_OP_425J2_127_3477_n3004) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2100 ( .A1(DP_OP_425J2_127_3477_n2885), 
        .A2(DP_OP_425J2_127_3477_n2891), .Y(DP_OP_425J2_127_3477_n2861) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2197 ( .A1(DP_OP_422J2_124_3477_n2974), 
        .A2(DP_OP_422J2_124_3477_n2980), .Y(DP_OP_422J2_124_3477_n2958) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1720 ( .A1(DP_OP_422J2_124_3477_n2489), 
        .A2(DP_OP_425J2_127_3477_n2497), .Y(DP_OP_422J2_124_3477_n2481) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1664 ( .A1(DP_OP_425J2_127_3477_n2449), 
        .A2(n789), .Y(DP_OP_425J2_127_3477_n2425) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1658 ( .A1(DP_OP_424J2_126_3477_n2619), 
        .A2(n261), .Y(DP_OP_425J2_127_3477_n2419) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1532 ( .A1(DP_OP_423J2_125_3477_n2845), 
        .A2(DP_OP_425J2_127_3477_n2319), .Y(DP_OP_425J2_127_3477_n2293) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1482 ( .A1(DP_OP_424J2_126_3477_n2795), 
        .A2(DP_OP_424J2_126_3477_n2275), .Y(DP_OP_425J2_127_3477_n2243) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1576 ( .A1(DP_OP_423J2_125_3477_n2801), 
        .A2(n874), .Y(DP_OP_425J2_127_3477_n2337) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1236 ( .A1(DP_OP_422J2_124_3477_n2005), 
        .A2(DP_OP_422J2_124_3477_n2013), .Y(DP_OP_422J2_124_3477_n1997) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1237 ( .A1(DP_OP_422J2_124_3477_n2006), 
        .A2(DP_OP_422J2_124_3477_n2013), .Y(DP_OP_422J2_124_3477_n1998) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1275 ( .A1(DP_OP_424J2_126_3477_n3020), 
        .A2(DP_OP_425J2_127_3477_n2056), .Y(DP_OP_425J2_127_3477_n2036) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1572 ( .A1(DP_OP_425J2_127_3477_n2577), 
        .A2(n876), .Y(DP_OP_423J2_125_3477_n2333) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1273 ( .A1(DP_OP_425J2_127_3477_n2182), 
        .A2(DP_OP_422J2_124_3477_n2056), .Y(DP_OP_422J2_124_3477_n2034) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1172 ( .A1(n1872), .A2(n1508), .Y(
        DP_OP_422J2_124_3477_n1933) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2111 ( .A1(DP_OP_425J2_127_3477_n2888), 
        .A2(DP_OP_423J2_125_3477_n2892), .Y(DP_OP_425J2_127_3477_n2872) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2104 ( .A1(DP_OP_422J2_124_3477_n3021), 
        .A2(DP_OP_423J2_125_3477_n2891), .Y(DP_OP_425J2_127_3477_n2865) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1239 ( .A1(DP_OP_425J2_127_3477_n2008), 
        .A2(n1431), .Y(DP_OP_425J2_127_3477_n2000) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2205 ( .A1(DP_OP_422J2_124_3477_n2974), 
        .A2(n677), .Y(DP_OP_422J2_124_3477_n2966) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2073 ( .A1(DP_OP_423J2_125_3477_n2094), 
        .A2(n1428), .Y(DP_OP_425J2_127_3477_n2834) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1274 ( .A1(DP_OP_422J2_124_3477_n2051), 
        .A2(DP_OP_422J2_124_3477_n2056), .Y(DP_OP_422J2_124_3477_n2035) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2148 ( .A1(DP_OP_425J2_127_3477_n2801), 
        .A2(DP_OP_425J2_127_3477_n2935), .Y(DP_OP_422J2_124_3477_n2909) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1722 ( .A1(DP_OP_423J2_125_3477_n2667), 
        .A2(DP_OP_425J2_127_3477_n2497), .Y(DP_OP_425J2_127_3477_n2483) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1485 ( .A1(DP_OP_423J2_125_3477_n2886), 
        .A2(DP_OP_424J2_126_3477_n2275), .Y(DP_OP_425J2_127_3477_n2246) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2199 ( .A1(DP_OP_425J2_127_3477_n2976), 
        .A2(DP_OP_424J2_126_3477_n2980), .Y(DP_OP_425J2_127_3477_n2960) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1488 ( .A1(DP_OP_424J2_126_3477_n2801), 
        .A2(DP_OP_422J2_124_3477_n2275), .Y(DP_OP_425J2_127_3477_n2249) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2148 ( .A1(DP_OP_425J2_127_3477_n2933), 
        .A2(n1432), .Y(DP_OP_425J2_127_3477_n2909) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1763 ( .A1(DP_OP_422J2_124_3477_n2664), 
        .A2(DP_OP_425J2_127_3477_n2541), .Y(DP_OP_425J2_127_3477_n2524) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2203 ( .A1(DP_OP_425J2_127_3477_n2972), 
        .A2(n677), .Y(DP_OP_425J2_127_3477_n2964) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2196 ( .A1(DP_OP_425J2_127_3477_n2973), 
        .A2(DP_OP_422J2_124_3477_n2980), .Y(DP_OP_425J2_127_3477_n2957) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1272 ( .A1(DP_OP_425J2_127_3477_n2049), 
        .A2(DP_OP_425J2_127_3477_n2056), .Y(DP_OP_425J2_127_3477_n2033) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1529 ( .A1(DP_OP_423J2_125_3477_n2842), 
        .A2(DP_OP_425J2_127_3477_n2319), .Y(DP_OP_425J2_127_3477_n2290) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2240 ( .A1(DP_OP_424J2_126_3477_n2005), 
        .A2(n704), .Y(DP_OP_425J2_127_3477_n3001) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1414 ( .A1(DP_OP_422J2_124_3477_n2051), 
        .A2(DP_OP_425J2_127_3477_n2189), .Y(DP_OP_425J2_127_3477_n2175) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1706 ( .A1(DP_OP_422J2_124_3477_n2491), 
        .A2(DP_OP_422J2_124_3477_n2495), .Y(DP_OP_422J2_124_3477_n2467) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2206 ( .A1(DP_OP_424J2_126_3477_n2051), 
        .A2(n677), .Y(DP_OP_425J2_127_3477_n2967) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1571 ( .A1(DP_OP_425J2_127_3477_n2576), 
        .A2(n875), .Y(DP_OP_423J2_125_3477_n2332) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2074 ( .A1(DP_OP_425J2_127_3477_n2843), 
        .A2(n1428), .Y(DP_OP_425J2_127_3477_n2835) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2204 ( .A1(DP_OP_422J2_124_3477_n2973), 
        .A2(n677), .Y(DP_OP_422J2_124_3477_n2965) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1972 ( .A1(DP_OP_422J2_124_3477_n2889), 
        .A2(DP_OP_422J2_124_3477_n2759), .Y(DP_OP_425J2_127_3477_n2733) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1415 ( .A1(DP_OP_424J2_126_3477_n2184), 
        .A2(DP_OP_424J2_126_3477_n2189), .Y(DP_OP_424J2_126_3477_n2176) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2075 ( .A1(DP_OP_423J2_125_3477_n2932), 
        .A2(DP_OP_423J2_125_3477_n2849), .Y(DP_OP_424J2_126_3477_n2836) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2144 ( .A1(DP_OP_423J2_125_3477_n2005), 
        .A2(DP_OP_422J2_124_3477_n2935), .Y(DP_OP_425J2_127_3477_n2905) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1416 ( .A1(DP_OP_424J2_126_3477_n2185), 
        .A2(DP_OP_424J2_126_3477_n2189), .Y(DP_OP_424J2_126_3477_n2177) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1413 ( .A1(DP_OP_424J2_126_3477_n2754), 
        .A2(DP_OP_422J2_124_3477_n2189), .Y(DP_OP_422J2_124_3477_n2174) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1487 ( .A1(DP_OP_425J2_127_3477_n2404), 
        .A2(n1427), .Y(DP_OP_422J2_124_3477_n2248) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1704 ( .A1(DP_OP_422J2_124_3477_n2489), 
        .A2(DP_OP_422J2_124_3477_n2495), .Y(DP_OP_422J2_124_3477_n2465) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2205 ( .A1(DP_OP_425J2_127_3477_n2974), 
        .A2(n676), .Y(DP_OP_425J2_127_3477_n2966) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1723 ( .A1(DP_OP_425J2_127_3477_n2536), 
        .A2(DP_OP_422J2_124_3477_n2497), .Y(DP_OP_424J2_126_3477_n2484) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1528 ( .A1(DP_OP_423J2_125_3477_n2841), 
        .A2(DP_OP_425J2_127_3477_n2319), .Y(DP_OP_425J2_127_3477_n2289) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2103 ( .A1(DP_OP_422J2_124_3477_n2888), 
        .A2(DP_OP_425J2_127_3477_n2891), .Y(DP_OP_422J2_124_3477_n2864) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1168 ( .A1(n1278), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_423J2_125_3477_n1929) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1531 ( .A1(DP_OP_423J2_125_3477_n2844), 
        .A2(DP_OP_425J2_127_3477_n2319), .Y(DP_OP_425J2_127_3477_n2292) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1484 ( .A1(DP_OP_425J2_127_3477_n2269), 
        .A2(DP_OP_424J2_126_3477_n2275), .Y(DP_OP_425J2_127_3477_n2245) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1768 ( .A1(DP_OP_422J2_124_3477_n2405), 
        .A2(DP_OP_424J2_126_3477_n2541), .Y(DP_OP_424J2_126_3477_n2529) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1271 ( .A1(DP_OP_425J2_127_3477_n2048), 
        .A2(DP_OP_425J2_127_3477_n2056), .Y(DP_OP_425J2_127_3477_n2032) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1724 ( .A1(DP_OP_423J2_125_3477_n2405), 
        .A2(DP_OP_425J2_127_3477_n2497), .Y(DP_OP_424J2_126_3477_n2485) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2147 ( .A1(DP_OP_425J2_127_3477_n2800), 
        .A2(DP_OP_422J2_124_3477_n2935), .Y(DP_OP_422J2_124_3477_n2908) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2239 ( .A1(DP_OP_424J2_126_3477_n2004), 
        .A2(n704), .Y(DP_OP_425J2_127_3477_n3000) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2202 ( .A1(DP_OP_425J2_127_3477_n2971), 
        .A2(n677), .Y(DP_OP_425J2_127_3477_n2963) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2076 ( .A1(DP_OP_424J2_126_3477_n2845), 
        .A2(DP_OP_423J2_125_3477_n2849), .Y(DP_OP_424J2_126_3477_n2837) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1487 ( .A1(DP_OP_425J2_127_3477_n2272), 
        .A2(n1427), .Y(DP_OP_425J2_127_3477_n2248) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2239 ( .A1(DP_OP_424J2_126_3477_n2928), 
        .A2(n704), .Y(DP_OP_423J2_125_3477_n3000) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1765 ( .A1(DP_OP_422J2_124_3477_n2534), 
        .A2(DP_OP_422J2_124_3477_n2541), .Y(DP_OP_422J2_124_3477_n2526) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2244 ( .A1(DP_OP_425J2_127_3477_n2053), 
        .A2(n703), .Y(DP_OP_424J2_126_3477_n3005) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2195 ( .A1(DP_OP_425J2_127_3477_n2972), 
        .A2(DP_OP_424J2_126_3477_n2980), .Y(DP_OP_425J2_127_3477_n2956) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2147 ( .A1(DP_OP_423J2_125_3477_n2008), 
        .A2(n1432), .Y(DP_OP_425J2_127_3477_n2908) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1276 ( .A1(DP_OP_425J2_127_3477_n2977), 
        .A2(DP_OP_424J2_126_3477_n2056), .Y(DP_OP_424J2_126_3477_n2037) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2110 ( .A1(DP_OP_422J2_124_3477_n2887), 
        .A2(DP_OP_423J2_125_3477_n2892), .Y(DP_OP_422J2_124_3477_n2871) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1410 ( .A1(DP_OP_422J2_124_3477_n2179), 
        .A2(DP_OP_422J2_124_3477_n2189), .Y(DP_OP_422J2_124_3477_n2171) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2242 ( .A1(DP_OP_425J2_127_3477_n3019), 
        .A2(n704), .Y(DP_OP_425J2_127_3477_n3003) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2198 ( .A1(DP_OP_424J2_126_3477_n2051), 
        .A2(DP_OP_425J2_127_3477_n2980), .Y(DP_OP_425J2_127_3477_n2959) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1705 ( .A1(DP_OP_422J2_124_3477_n2578), 
        .A2(DP_OP_422J2_124_3477_n2495), .Y(DP_OP_423J2_125_3477_n2466) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2107 ( .A1(DP_OP_423J2_125_3477_n2048), 
        .A2(DP_OP_423J2_125_3477_n2892), .Y(DP_OP_425J2_127_3477_n2868) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2200 ( .A1(DP_OP_424J2_126_3477_n2977), 
        .A2(DP_OP_424J2_126_3477_n2980), .Y(DP_OP_424J2_126_3477_n2961) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2207 ( .A1(DP_OP_424J2_126_3477_n2976), 
        .A2(n677), .Y(DP_OP_424J2_126_3477_n2968) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2112 ( .A1(DP_OP_424J2_126_3477_n2889), 
        .A2(DP_OP_423J2_125_3477_n2892), .Y(DP_OP_424J2_126_3477_n2873) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2208 ( .A1(DP_OP_424J2_126_3477_n2977), 
        .A2(n677), .Y(DP_OP_424J2_126_3477_n2969) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1704 ( .A1(DP_OP_422J2_124_3477_n2577), 
        .A2(DP_OP_422J2_124_3477_n2495), .Y(DP_OP_423J2_125_3477_n2465) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1274 ( .A1(DP_OP_424J2_126_3477_n3019), 
        .A2(DP_OP_425J2_127_3477_n2056), .Y(DP_OP_425J2_127_3477_n2035) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1966 ( .A1(DP_OP_422J2_124_3477_n2883), 
        .A2(DP_OP_422J2_124_3477_n2759), .Y(DP_OP_425J2_127_3477_n2727) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1416 ( .A1(DP_OP_425J2_127_3477_n2185), 
        .A2(DP_OP_425J2_127_3477_n2189), .Y(DP_OP_425J2_127_3477_n2177) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1413 ( .A1(DP_OP_425J2_127_3477_n2182), 
        .A2(DP_OP_425J2_127_3477_n2189), .Y(DP_OP_425J2_127_3477_n2174) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1326 ( .A1(DP_OP_423J2_125_3477_n2931), 
        .A2(n621), .Y(DP_OP_422J2_124_3477_n2087) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1354 ( .A1(DP_OP_425J2_127_3477_n2799), 
        .A2(DP_OP_425J2_127_3477_n2143), .Y(DP_OP_423J2_125_3477_n2115) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1807 ( .A1(DP_OP_422J2_124_3477_n2444), 
        .A2(DP_OP_423J2_125_3477_n2585), .Y(DP_OP_423J2_125_3477_n2568) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1890 ( .A1(DP_OP_422J2_124_3477_n2667), 
        .A2(n279), .Y(DP_OP_422J2_124_3477_n2651) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1582 ( .A1(DP_OP_423J2_125_3477_n2667), 
        .A2(n1386), .Y(DP_OP_422J2_124_3477_n2343) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1440 ( .A1(DP_OP_423J2_125_3477_n2225), 
        .A2(DP_OP_422J2_124_3477_n2231), .Y(DP_OP_423J2_125_3477_n2201) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1320 ( .A1(DP_OP_424J2_126_3477_n2845), 
        .A2(DP_OP_424J2_126_3477_n2100), .Y(DP_OP_422J2_124_3477_n2081) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1352 ( .A1(DP_OP_425J2_127_3477_n2797), 
        .A2(DP_OP_425J2_127_3477_n2143), .Y(DP_OP_423J2_125_3477_n2113) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1319 ( .A1(DP_OP_423J2_125_3477_n2932), 
        .A2(DP_OP_424J2_126_3477_n2100), .Y(DP_OP_422J2_124_3477_n2080) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1755 ( .A1(DP_OP_422J2_124_3477_n2532), 
        .A2(n1486), .Y(DP_OP_422J2_124_3477_n2516) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1792 ( .A1(DP_OP_422J2_124_3477_n2445), 
        .A2(n671), .Y(DP_OP_423J2_125_3477_n2553) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1442 ( .A1(DP_OP_423J2_125_3477_n2227), 
        .A2(DP_OP_424J2_126_3477_n2231), .Y(DP_OP_423J2_125_3477_n2203) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1888 ( .A1(DP_OP_423J2_125_3477_n2665), 
        .A2(n279), .Y(DP_OP_423J2_125_3477_n2649) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2019 ( .A1(DP_OP_422J2_124_3477_n2224), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_423J2_125_3477_n2780) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1748 ( .A1(DP_OP_422J2_124_3477_n2533), 
        .A2(n771), .Y(DP_OP_422J2_124_3477_n2509) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2287 ( .A1(DP_OP_423J2_125_3477_n2008), 
        .A2(DP_OP_425J2_127_3477_n3066), .Y(DP_OP_422J2_124_3477_n3046) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1900 ( .A1(DP_OP_422J2_124_3477_n2669), 
        .A2(DP_OP_424J2_126_3477_n2673), .Y(DP_OP_422J2_124_3477_n2661) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1327 ( .A1(DP_OP_423J2_125_3477_n2932), 
        .A2(n621), .Y(DP_OP_422J2_124_3477_n2088) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1812 ( .A1(DP_OP_423J2_125_3477_n2493), 
        .A2(DP_OP_424J2_126_3477_n2585), .Y(DP_OP_422J2_124_3477_n2573) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1356 ( .A1(DP_OP_423J2_125_3477_n2889), 
        .A2(DP_OP_422J2_124_3477_n2143), .Y(DP_OP_422J2_124_3477_n2117) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1444 ( .A1(DP_OP_423J2_125_3477_n2801), 
        .A2(DP_OP_424J2_126_3477_n2231), .Y(DP_OP_422J2_124_3477_n2205) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1324 ( .A1(DP_OP_422J2_124_3477_n2093), 
        .A2(n621), .Y(DP_OP_422J2_124_3477_n2085) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1317 ( .A1(DP_OP_423J2_125_3477_n2094), 
        .A2(DP_OP_424J2_126_3477_n2100), .Y(DP_OP_423J2_125_3477_n2078) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1440 ( .A1(DP_OP_422J2_124_3477_n2225), 
        .A2(DP_OP_424J2_126_3477_n2231), .Y(DP_OP_422J2_124_3477_n2201) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1281 ( .A1(DP_OP_424J2_126_3477_n2886), 
        .A2(n1475), .Y(DP_OP_422J2_124_3477_n2042) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2235 ( .A1(DP_OP_423J2_125_3477_n2052), 
        .A2(DP_OP_424J2_126_3477_n3023), .Y(DP_OP_422J2_124_3477_n2996) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2056 ( .A1(DP_OP_422J2_124_3477_n2841), 
        .A2(DP_OP_422J2_124_3477_n2847), .Y(DP_OP_422J2_124_3477_n2817) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1895 ( .A1(DP_OP_424J2_126_3477_n2576), 
        .A2(DP_OP_422J2_124_3477_n2673), .Y(DP_OP_423J2_125_3477_n2656) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1758 ( .A1(DP_OP_422J2_124_3477_n2535), 
        .A2(n1487), .Y(DP_OP_422J2_124_3477_n2519) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2024 ( .A1(DP_OP_422J2_124_3477_n2801), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_422J2_124_3477_n2785) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1538 ( .A1(DP_OP_425J2_127_3477_n2447), 
        .A2(DP_OP_425J2_127_3477_n2320), .Y(DP_OP_422J2_124_3477_n2299) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1811 ( .A1(DP_OP_422J2_124_3477_n2580), 
        .A2(DP_OP_424J2_126_3477_n2585), .Y(DP_OP_422J2_124_3477_n2572) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1368 ( .A1(DP_OP_422J2_124_3477_n2137), 
        .A2(n1500), .Y(DP_OP_422J2_124_3477_n2129) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1666 ( .A1(DP_OP_422J2_124_3477_n2443), 
        .A2(n1489), .Y(DP_OP_422J2_124_3477_n2427) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1927 ( .A1(DP_OP_422J2_124_3477_n2712), 
        .A2(DP_OP_422J2_124_3477_n2715), .Y(DP_OP_422J2_124_3477_n2688) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1317 ( .A1(DP_OP_425J2_127_3477_n2226), 
        .A2(DP_OP_422J2_124_3477_n2100), .Y(DP_OP_422J2_124_3477_n2078) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2232 ( .A1(DP_OP_422J2_124_3477_n3017), 
        .A2(DP_OP_425J2_127_3477_n3023), .Y(DP_OP_422J2_124_3477_n2993) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1889 ( .A1(DP_OP_425J2_127_3477_n2534), 
        .A2(n279), .Y(DP_OP_422J2_124_3477_n2650) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1672 ( .A1(DP_OP_423J2_125_3477_n2581), 
        .A2(DP_OP_423J2_125_3477_n2452), .Y(DP_OP_422J2_124_3477_n2433) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1578 ( .A1(DP_OP_422J2_124_3477_n2355), 
        .A2(DP_OP_423J2_125_3477_n2364), .Y(DP_OP_422J2_124_3477_n2339) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1282 ( .A1(DP_OP_422J2_124_3477_n2051), 
        .A2(DP_OP_425J2_127_3477_n2057), .Y(DP_OP_422J2_124_3477_n2043) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1896 ( .A1(DP_OP_422J2_124_3477_n2665), 
        .A2(DP_OP_425J2_127_3477_n2673), .Y(DP_OP_422J2_124_3477_n2657) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1315 ( .A1(DP_OP_422J2_124_3477_n2092), 
        .A2(DP_OP_424J2_126_3477_n2100), .Y(DP_OP_422J2_124_3477_n2076) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2059 ( .A1(DP_OP_423J2_125_3477_n2228), 
        .A2(DP_OP_425J2_127_3477_n2847), .Y(DP_OP_422J2_124_3477_n2820) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1284 ( .A1(DP_OP_424J2_126_3477_n2889), 
        .A2(DP_OP_424J2_126_3477_n2057), .Y(DP_OP_422J2_124_3477_n2045) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1324 ( .A1(DP_OP_425J2_127_3477_n2841), 
        .A2(n621), .Y(DP_OP_423J2_125_3477_n2085) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1791 ( .A1(DP_OP_422J2_124_3477_n2576), 
        .A2(n671), .Y(DP_OP_422J2_124_3477_n2552) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1711 ( .A1(DP_OP_422J2_124_3477_n2488), 
        .A2(n1491), .Y(DP_OP_422J2_124_3477_n2472) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2286 ( .A1(DP_OP_423J2_125_3477_n2007), 
        .A2(DP_OP_424J2_126_3477_n3066), .Y(DP_OP_422J2_124_3477_n3045) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1354 ( .A1(DP_OP_424J2_126_3477_n2799), 
        .A2(DP_OP_422J2_124_3477_n2143), .Y(DP_OP_422J2_124_3477_n2115) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1747 ( .A1(DP_OP_422J2_124_3477_n2532), 
        .A2(n772), .Y(DP_OP_422J2_124_3477_n2508) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1372 ( .A1(DP_OP_423J2_125_3477_n2889), 
        .A2(n1501), .Y(DP_OP_422J2_124_3477_n2133) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1351 ( .A1(DP_OP_425J2_127_3477_n2796), 
        .A2(DP_OP_424J2_126_3477_n2143), .Y(DP_OP_423J2_125_3477_n2112) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1283 ( .A1(DP_OP_425J2_127_3477_n2184), 
        .A2(DP_OP_424J2_126_3477_n2057), .Y(DP_OP_422J2_124_3477_n2044) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1794 ( .A1(DP_OP_422J2_124_3477_n2579), 
        .A2(n671), .Y(DP_OP_422J2_124_3477_n2555) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1795 ( .A1(DP_OP_422J2_124_3477_n2580), 
        .A2(n671), .Y(DP_OP_422J2_124_3477_n2556) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1886 ( .A1(DP_OP_422J2_124_3477_n2663), 
        .A2(n279), .Y(DP_OP_422J2_124_3477_n2647) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1899 ( .A1(DP_OP_423J2_125_3477_n2404), 
        .A2(DP_OP_424J2_126_3477_n2673), .Y(DP_OP_422J2_124_3477_n2660) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1900 ( .A1(DP_OP_422J2_124_3477_n2801), 
        .A2(n1), .Y(DP_OP_425J2_127_3477_n2661) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1794 ( .A1(DP_OP_423J2_125_3477_n2579), 
        .A2(n671), .Y(DP_OP_423J2_125_3477_n2555) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1755 ( .A1(DP_OP_422J2_124_3477_n2488), 
        .A2(n1486), .Y(DP_OP_423J2_125_3477_n2516) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1280 ( .A1(DP_OP_425J2_127_3477_n2885), 
        .A2(DP_OP_424J2_126_3477_n2057), .Y(DP_OP_423J2_125_3477_n2041) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1808 ( .A1(DP_OP_422J2_124_3477_n2445), 
        .A2(DP_OP_424J2_126_3477_n2585), .Y(DP_OP_423J2_125_3477_n2569) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1757 ( .A1(DP_OP_422J2_124_3477_n2490), 
        .A2(DP_OP_424J2_126_3477_n2540), .Y(DP_OP_423J2_125_3477_n2518) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2234 ( .A1(DP_OP_422J2_124_3477_n3019), 
        .A2(DP_OP_424J2_126_3477_n3023), .Y(DP_OP_422J2_124_3477_n2995) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1537 ( .A1(DP_OP_422J2_124_3477_n2314), 
        .A2(DP_OP_423J2_125_3477_n2320), .Y(DP_OP_422J2_124_3477_n2298) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1896 ( .A1(DP_OP_423J2_125_3477_n2665), 
        .A2(DP_OP_422J2_124_3477_n2673), .Y(DP_OP_423J2_125_3477_n2657) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1889 ( .A1(DP_OP_423J2_125_3477_n2666), 
        .A2(n279), .Y(DP_OP_423J2_125_3477_n2650) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1887 ( .A1(DP_OP_422J2_124_3477_n2664), 
        .A2(n279), .Y(DP_OP_422J2_124_3477_n2648) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1366 ( .A1(DP_OP_422J2_124_3477_n2135), 
        .A2(n1501), .Y(DP_OP_422J2_124_3477_n2127) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1793 ( .A1(DP_OP_422J2_124_3477_n2446), 
        .A2(n671), .Y(DP_OP_423J2_125_3477_n2554) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1535 ( .A1(DP_OP_422J2_124_3477_n2312), 
        .A2(DP_OP_422J2_124_3477_n2320), .Y(DP_OP_422J2_124_3477_n2296) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1808 ( .A1(DP_OP_422J2_124_3477_n2577), 
        .A2(DP_OP_422J2_124_3477_n2585), .Y(DP_OP_422J2_124_3477_n2569) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1666 ( .A1(DP_OP_422J2_124_3477_n2619), 
        .A2(DP_OP_423J2_125_3477_n2452), .Y(DP_OP_423J2_125_3477_n2427) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1634 ( .A1(DP_OP_424J2_126_3477_n2535), 
        .A2(DP_OP_423J2_125_3477_n2409), .Y(DP_OP_422J2_124_3477_n2395) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1810 ( .A1(DP_OP_422J2_124_3477_n2579), 
        .A2(DP_OP_423J2_125_3477_n2585), .Y(DP_OP_422J2_124_3477_n2571) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1898 ( .A1(DP_OP_422J2_124_3477_n2667), 
        .A2(DP_OP_425J2_127_3477_n2673), .Y(DP_OP_422J2_124_3477_n2659) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1671 ( .A1(DP_OP_422J2_124_3477_n2448), 
        .A2(n1488), .Y(DP_OP_422J2_124_3477_n2432) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2233 ( .A1(DP_OP_422J2_124_3477_n2006), 
        .A2(DP_OP_424J2_126_3477_n3023), .Y(DP_OP_423J2_125_3477_n2994) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1757 ( .A1(DP_OP_422J2_124_3477_n2534), 
        .A2(n1486), .Y(DP_OP_422J2_124_3477_n2518) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1759 ( .A1(DP_OP_422J2_124_3477_n2536), 
        .A2(n1487), .Y(DP_OP_422J2_124_3477_n2520) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1539 ( .A1(DP_OP_425J2_127_3477_n2448), 
        .A2(DP_OP_423J2_125_3477_n2320), .Y(DP_OP_422J2_124_3477_n2300) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1752 ( .A1(DP_OP_422J2_124_3477_n2537), 
        .A2(n771), .Y(DP_OP_422J2_124_3477_n2513) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1669 ( .A1(DP_OP_422J2_124_3477_n2622), 
        .A2(n1489), .Y(DP_OP_423J2_125_3477_n2430) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1928 ( .A1(DP_OP_423J2_125_3477_n2361), 
        .A2(n1497), .Y(DP_OP_422J2_124_3477_n2689) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1540 ( .A1(DP_OP_425J2_127_3477_n2449), 
        .A2(DP_OP_422J2_124_3477_n2320), .Y(DP_OP_422J2_124_3477_n2301) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2282 ( .A1(DP_OP_422J2_124_3477_n3057), 
        .A2(DP_OP_423J2_125_3477_n3066), .Y(DP_OP_422J2_124_3477_n3041) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1667 ( .A1(DP_OP_422J2_124_3477_n2620), 
        .A2(DP_OP_423J2_125_3477_n2452), .Y(DP_OP_423J2_125_3477_n2428) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2232 ( .A1(DP_OP_424J2_126_3477_n2929), 
        .A2(DP_OP_422J2_124_3477_n3023), .Y(DP_OP_423J2_125_3477_n2993) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1713 ( .A1(DP_OP_422J2_124_3477_n2578), 
        .A2(DP_OP_423J2_125_3477_n2496), .Y(DP_OP_423J2_125_3477_n2474) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1537 ( .A1(DP_OP_425J2_127_3477_n2622), 
        .A2(DP_OP_422J2_124_3477_n2320), .Y(DP_OP_423J2_125_3477_n2298) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2231 ( .A1(DP_OP_423J2_125_3477_n2048), 
        .A2(DP_OP_425J2_127_3477_n3023), .Y(DP_OP_422J2_124_3477_n2992) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1923 ( .A1(DP_OP_423J2_125_3477_n2708), 
        .A2(DP_OP_422J2_124_3477_n2715), .Y(DP_OP_423J2_125_3477_n2684) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1670 ( .A1(DP_OP_423J2_125_3477_n2579), 
        .A2(DP_OP_423J2_125_3477_n2452), .Y(DP_OP_422J2_124_3477_n2431) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1323 ( .A1(DP_OP_425J2_127_3477_n2840), 
        .A2(n621), .Y(DP_OP_423J2_125_3477_n2084) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1579 ( .A1(DP_OP_425J2_127_3477_n2576), 
        .A2(n1386), .Y(DP_OP_423J2_125_3477_n2340) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2021 ( .A1(DP_OP_423J2_125_3477_n2798), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_423J2_125_3477_n2782) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1751 ( .A1(DP_OP_422J2_124_3477_n2536), 
        .A2(n772), .Y(DP_OP_422J2_124_3477_n2512) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1924 ( .A1(DP_OP_422J2_124_3477_n2313), 
        .A2(n1497), .Y(DP_OP_423J2_125_3477_n2685) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2021 ( .A1(DP_OP_422J2_124_3477_n2798), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_422J2_124_3477_n2782) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1442 ( .A1(DP_OP_425J2_127_3477_n2359), 
        .A2(DP_OP_424J2_126_3477_n2231), .Y(DP_OP_422J2_124_3477_n2203) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1369 ( .A1(DP_OP_422J2_124_3477_n2138), 
        .A2(n1501), .Y(DP_OP_422J2_124_3477_n2130) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2236 ( .A1(DP_OP_422J2_124_3477_n3021), 
        .A2(DP_OP_422J2_124_3477_n3023), .Y(DP_OP_422J2_124_3477_n2997) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1355 ( .A1(DP_OP_422J2_124_3477_n2140), 
        .A2(DP_OP_422J2_124_3477_n2143), .Y(DP_OP_422J2_124_3477_n2116) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1318 ( .A1(DP_OP_423J2_125_3477_n2931), 
        .A2(DP_OP_422J2_124_3477_n2100), .Y(DP_OP_422J2_124_3477_n2079) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1325 ( .A1(DP_OP_425J2_127_3477_n2226), 
        .A2(n621), .Y(DP_OP_422J2_124_3477_n2086) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1316 ( .A1(DP_OP_425J2_127_3477_n2841), 
        .A2(DP_OP_423J2_125_3477_n2100), .Y(DP_OP_423J2_125_3477_n2077) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1925 ( .A1(DP_OP_422J2_124_3477_n2314), 
        .A2(DP_OP_422J2_124_3477_n2715), .Y(DP_OP_423J2_125_3477_n2686) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1796 ( .A1(DP_OP_423J2_125_3477_n2493), 
        .A2(n670), .Y(DP_OP_422J2_124_3477_n2557) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1842 ( .A1(DP_OP_422J2_124_3477_n2619), 
        .A2(n1499), .Y(DP_OP_422J2_124_3477_n2603) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1371 ( .A1(DP_OP_422J2_124_3477_n2140), 
        .A2(n1501), .Y(DP_OP_422J2_124_3477_n2132) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1714 ( .A1(DP_OP_422J2_124_3477_n2491), 
        .A2(n1491), .Y(DP_OP_422J2_124_3477_n2475) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1756 ( .A1(DP_OP_422J2_124_3477_n2489), 
        .A2(DP_OP_424J2_126_3477_n2540), .Y(DP_OP_423J2_125_3477_n2517) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1633 ( .A1(DP_OP_424J2_126_3477_n2534), 
        .A2(DP_OP_424J2_126_3477_n2409), .Y(DP_OP_422J2_124_3477_n2394) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1897 ( .A1(DP_OP_425J2_127_3477_n2534), 
        .A2(DP_OP_425J2_127_3477_n2673), .Y(DP_OP_422J2_124_3477_n2658) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2284 ( .A1(DP_OP_423J2_125_3477_n3059), 
        .A2(DP_OP_423J2_125_3477_n3066), .Y(DP_OP_423J2_125_3477_n3043) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1750 ( .A1(DP_OP_422J2_124_3477_n2535), 
        .A2(n772), .Y(DP_OP_422J2_124_3477_n2511) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1891 ( .A1(DP_OP_425J2_127_3477_n2536), 
        .A2(n278), .Y(DP_OP_422J2_124_3477_n2652) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1926 ( .A1(DP_OP_424J2_126_3477_n2623), 
        .A2(DP_OP_422J2_124_3477_n2715), .Y(DP_OP_423J2_125_3477_n2687) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2022 ( .A1(DP_OP_422J2_124_3477_n2799), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_422J2_124_3477_n2783) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1353 ( .A1(DP_OP_425J2_127_3477_n2798), 
        .A2(DP_OP_424J2_126_3477_n2143), .Y(DP_OP_423J2_125_3477_n2114) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1926 ( .A1(DP_OP_425J2_127_3477_n2579), 
        .A2(n1497), .Y(DP_OP_422J2_124_3477_n2687) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1316 ( .A1(DP_OP_423J2_125_3477_n2005), 
        .A2(DP_OP_423J2_125_3477_n2100), .Y(DP_OP_424J2_126_3477_n2077) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1756 ( .A1(DP_OP_422J2_124_3477_n2401), 
        .A2(n1486), .Y(DP_OP_424J2_126_3477_n2517) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1749 ( .A1(DP_OP_424J2_126_3477_n2534), 
        .A2(DP_OP_425J2_127_3477_n2539), .Y(DP_OP_424J2_126_3477_n2510) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1353 ( .A1(DP_OP_424J2_126_3477_n2138), 
        .A2(DP_OP_424J2_126_3477_n2143), .Y(DP_OP_424J2_126_3477_n2114) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1372 ( .A1(DP_OP_423J2_125_3477_n3021), 
        .A2(n1500), .Y(DP_OP_425J2_127_3477_n2133) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1812 ( .A1(DP_OP_425J2_127_3477_n2581), 
        .A2(DP_OP_424J2_126_3477_n2585), .Y(DP_OP_425J2_127_3477_n2573) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1538 ( .A1(DP_OP_423J2_125_3477_n2843), 
        .A2(DP_OP_422J2_124_3477_n2320), .Y(DP_OP_425J2_127_3477_n2299) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1281 ( .A1(DP_OP_425J2_127_3477_n2050), 
        .A2(DP_OP_425J2_127_3477_n2057), .Y(DP_OP_425J2_127_3477_n2042) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1897 ( .A1(DP_OP_422J2_124_3477_n2798), 
        .A2(n1), .Y(DP_OP_425J2_127_3477_n2658) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1633 ( .A1(DP_OP_423J2_125_3477_n2754), 
        .A2(DP_OP_425J2_127_3477_n2409), .Y(DP_OP_425J2_127_3477_n2394) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1325 ( .A1(DP_OP_423J2_125_3477_n3060), 
        .A2(n621), .Y(DP_OP_425J2_127_3477_n2086) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1318 ( .A1(DP_OP_423J2_125_3477_n3061), 
        .A2(DP_OP_422J2_124_3477_n2100), .Y(DP_OP_425J2_127_3477_n2079) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1355 ( .A1(DP_OP_424J2_126_3477_n2932), 
        .A2(DP_OP_425J2_127_3477_n2143), .Y(DP_OP_425J2_127_3477_n2116) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1369 ( .A1(DP_OP_425J2_127_3477_n2138), 
        .A2(n1501), .Y(DP_OP_425J2_127_3477_n2130) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1751 ( .A1(DP_OP_425J2_127_3477_n2536), 
        .A2(n771), .Y(DP_OP_425J2_127_3477_n2512) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1670 ( .A1(DP_OP_425J2_127_3477_n2447), 
        .A2(DP_OP_423J2_125_3477_n2452), .Y(DP_OP_425J2_127_3477_n2431) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2059 ( .A1(DP_OP_423J2_125_3477_n2096), 
        .A2(DP_OP_425J2_127_3477_n2847), .Y(DP_OP_425J2_127_3477_n2820) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1539 ( .A1(DP_OP_423J2_125_3477_n2228), 
        .A2(DP_OP_425J2_127_3477_n2320), .Y(DP_OP_424J2_126_3477_n2300) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1795 ( .A1(DP_OP_425J2_127_3477_n2580), 
        .A2(n671), .Y(DP_OP_425J2_127_3477_n2556) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1890 ( .A1(DP_OP_422J2_124_3477_n2799), 
        .A2(n279), .Y(DP_OP_425J2_127_3477_n2651) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1351 ( .A1(DP_OP_424J2_126_3477_n2136), 
        .A2(DP_OP_424J2_126_3477_n2143), .Y(DP_OP_424J2_126_3477_n2112) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1314 ( .A1(DP_OP_423J2_125_3477_n2003), 
        .A2(DP_OP_423J2_125_3477_n2100), .Y(DP_OP_424J2_126_3477_n2075) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2235 ( .A1(DP_OP_425J2_127_3477_n3020), 
        .A2(DP_OP_425J2_127_3477_n3023), .Y(DP_OP_425J2_127_3477_n2996) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1540 ( .A1(DP_OP_424J2_126_3477_n2317), 
        .A2(DP_OP_425J2_127_3477_n2320), .Y(DP_OP_424J2_126_3477_n2301) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1443 ( .A1(DP_OP_423J2_125_3477_n2932), 
        .A2(DP_OP_425J2_127_3477_n2231), .Y(DP_OP_425J2_127_3477_n2204) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1439 ( .A1(DP_OP_425J2_127_3477_n2796), 
        .A2(DP_OP_424J2_126_3477_n2231), .Y(DP_OP_424J2_126_3477_n2200) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1758 ( .A1(DP_OP_422J2_124_3477_n2667), 
        .A2(n1487), .Y(DP_OP_425J2_127_3477_n2519) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2019 ( .A1(DP_OP_425J2_127_3477_n2796), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_425J2_127_3477_n2780) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2284 ( .A1(DP_OP_425J2_127_3477_n3059), 
        .A2(DP_OP_424J2_126_3477_n3066), .Y(DP_OP_425J2_127_3477_n3043) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2286 ( .A1(DP_OP_425J2_127_3477_n3061), 
        .A2(DP_OP_424J2_126_3477_n3066), .Y(DP_OP_425J2_127_3477_n3045) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1666 ( .A1(DP_OP_424J2_126_3477_n2443), 
        .A2(n1489), .Y(DP_OP_424J2_126_3477_n2427) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1582 ( .A1(DP_OP_425J2_127_3477_n2359), 
        .A2(n1386), .Y(DP_OP_425J2_127_3477_n2343) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1710 ( .A1(DP_OP_423J2_125_3477_n2399), 
        .A2(n1491), .Y(DP_OP_424J2_126_3477_n2471) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1578 ( .A1(DP_OP_423J2_125_3477_n2267), 
        .A2(n1386), .Y(DP_OP_424J2_126_3477_n2339) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1747 ( .A1(DP_OP_424J2_126_3477_n2532), 
        .A2(n772), .Y(DP_OP_424J2_126_3477_n2508) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1886 ( .A1(DP_OP_423J2_125_3477_n2751), 
        .A2(n279), .Y(DP_OP_424J2_126_3477_n2647) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1892 ( .A1(DP_OP_424J2_126_3477_n2669), 
        .A2(n279), .Y(DP_OP_424J2_126_3477_n2653) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2024 ( .A1(DP_OP_425J2_127_3477_n2801), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_425J2_127_3477_n2785) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1534 ( .A1(DP_OP_424J2_126_3477_n2311), 
        .A2(DP_OP_423J2_125_3477_n2320), .Y(DP_OP_424J2_126_3477_n2295) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2018 ( .A1(DP_OP_424J2_126_3477_n2795), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_424J2_126_3477_n2779) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1315 ( .A1(DP_OP_425J2_127_3477_n2092), 
        .A2(DP_OP_423J2_125_3477_n2100), .Y(DP_OP_425J2_127_3477_n2076) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1327 ( .A1(DP_OP_423J2_125_3477_n2096), 
        .A2(n621), .Y(DP_OP_423J2_125_3477_n2088) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1760 ( .A1(DP_OP_423J2_125_3477_n2537), 
        .A2(n1487), .Y(DP_OP_423J2_125_3477_n2521) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1716 ( .A1(DP_OP_423J2_125_3477_n2493), 
        .A2(n1491), .Y(DP_OP_423J2_125_3477_n2477) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2024 ( .A1(DP_OP_424J2_126_3477_n2801), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_424J2_126_3477_n2785) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1283 ( .A1(DP_OP_423J2_125_3477_n2052), 
        .A2(DP_OP_424J2_126_3477_n2057), .Y(DP_OP_423J2_125_3477_n2044) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1635 ( .A1(DP_OP_423J2_125_3477_n2404), 
        .A2(DP_OP_423J2_125_3477_n2409), .Y(DP_OP_423J2_125_3477_n2396) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1672 ( .A1(DP_OP_422J2_124_3477_n2625), 
        .A2(n1488), .Y(DP_OP_423J2_125_3477_n2433) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2024 ( .A1(DP_OP_423J2_125_3477_n2801), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_423J2_125_3477_n2785) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1672 ( .A1(DP_OP_423J2_125_3477_n2361), 
        .A2(DP_OP_423J2_125_3477_n2452), .Y(DP_OP_424J2_126_3477_n2433) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1636 ( .A1(DP_OP_423J2_125_3477_n2405), 
        .A2(DP_OP_424J2_126_3477_n2409), .Y(DP_OP_423J2_125_3477_n2397) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1635 ( .A1(DP_OP_422J2_124_3477_n2756), 
        .A2(DP_OP_424J2_126_3477_n2409), .Y(DP_OP_424J2_126_3477_n2396) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1900 ( .A1(DP_OP_423J2_125_3477_n2669), 
        .A2(DP_OP_424J2_126_3477_n2673), .Y(DP_OP_423J2_125_3477_n2661) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1793 ( .A1(DP_OP_423J2_125_3477_n2666), 
        .A2(DP_OP_422J2_124_3477_n2583), .Y(DP_OP_424J2_126_3477_n2554) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1812 ( .A1(DP_OP_423J2_125_3477_n2581), 
        .A2(DP_OP_422J2_124_3477_n2585), .Y(DP_OP_423J2_125_3477_n2573) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1790 ( .A1(DP_OP_424J2_126_3477_n2443), 
        .A2(n671), .Y(DP_OP_425J2_127_3477_n2551) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2057 ( .A1(DP_OP_425J2_127_3477_n2226), 
        .A2(DP_OP_425J2_127_3477_n2847), .Y(DP_OP_424J2_126_3477_n2818) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1320 ( .A1(DP_OP_425J2_127_3477_n2933), 
        .A2(DP_OP_422J2_124_3477_n2100), .Y(DP_OP_424J2_126_3477_n2081) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1712 ( .A1(DP_OP_423J2_125_3477_n2401), 
        .A2(DP_OP_423J2_125_3477_n2496), .Y(DP_OP_424J2_126_3477_n2473) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1371 ( .A1(DP_OP_423J2_125_3477_n2052), 
        .A2(n1500), .Y(DP_OP_424J2_126_3477_n2132) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1441 ( .A1(DP_OP_422J2_124_3477_n2930), 
        .A2(DP_OP_424J2_126_3477_n2231), .Y(DP_OP_424J2_126_3477_n2202) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1668 ( .A1(DP_OP_425J2_127_3477_n2577), 
        .A2(DP_OP_423J2_125_3477_n2452), .Y(DP_OP_424J2_126_3477_n2429) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1888 ( .A1(DP_OP_422J2_124_3477_n2269), 
        .A2(n278), .Y(DP_OP_424J2_126_3477_n2649) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1323 ( .A1(DP_OP_424J2_126_3477_n2092), 
        .A2(DP_OP_423J2_125_3477_n2101), .Y(DP_OP_424J2_126_3477_n2084) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2019 ( .A1(DP_OP_424J2_126_3477_n2796), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_424J2_126_3477_n2780) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1671 ( .A1(DP_OP_425J2_127_3477_n2580), 
        .A2(n1488), .Y(DP_OP_424J2_126_3477_n2432) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1440 ( .A1(DP_OP_425J2_127_3477_n2797), 
        .A2(DP_OP_422J2_124_3477_n2231), .Y(DP_OP_424J2_126_3477_n2201) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1714 ( .A1(DP_OP_423J2_125_3477_n2667), 
        .A2(DP_OP_423J2_125_3477_n2496), .Y(DP_OP_425J2_127_3477_n2475) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1315 ( .A1(DP_OP_424J2_126_3477_n2092), 
        .A2(DP_OP_424J2_126_3477_n2100), .Y(DP_OP_424J2_126_3477_n2076) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1583 ( .A1(DP_OP_422J2_124_3477_n2800), 
        .A2(n825), .Y(DP_OP_424J2_126_3477_n2344) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1748 ( .A1(DP_OP_423J2_125_3477_n2401), 
        .A2(n772), .Y(DP_OP_425J2_127_3477_n2509) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1667 ( .A1(DP_OP_425J2_127_3477_n2576), 
        .A2(n1488), .Y(DP_OP_424J2_126_3477_n2428) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1535 ( .A1(DP_OP_422J2_124_3477_n2840), 
        .A2(DP_OP_425J2_127_3477_n2320), .Y(DP_OP_424J2_126_3477_n2296) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2287 ( .A1(DP_OP_425J2_127_3477_n2008), 
        .A2(DP_OP_425J2_127_3477_n3066), .Y(DP_OP_424J2_126_3477_n3046) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1630 ( .A1(DP_OP_422J2_124_3477_n2751), 
        .A2(DP_OP_422J2_124_3477_n2409), .Y(DP_OP_424J2_126_3477_n2391) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1748 ( .A1(DP_OP_422J2_124_3477_n2401), 
        .A2(n772), .Y(DP_OP_424J2_126_3477_n2509) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1924 ( .A1(DP_OP_422J2_124_3477_n2225), 
        .A2(DP_OP_422J2_124_3477_n2715), .Y(DP_OP_424J2_126_3477_n2685) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1891 ( .A1(DP_OP_425J2_127_3477_n2404), 
        .A2(n278), .Y(DP_OP_424J2_126_3477_n2652) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1887 ( .A1(DP_OP_422J2_124_3477_n2268), 
        .A2(n279), .Y(DP_OP_424J2_126_3477_n2648) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2023 ( .A1(DP_OP_425J2_127_3477_n2272), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_424J2_126_3477_n2784) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1352 ( .A1(DP_OP_424J2_126_3477_n2929), 
        .A2(DP_OP_425J2_127_3477_n2143), .Y(DP_OP_425J2_127_3477_n2113) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1887 ( .A1(DP_OP_423J2_125_3477_n2268), 
        .A2(n279), .Y(DP_OP_425J2_127_3477_n2648) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2021 ( .A1(DP_OP_422J2_124_3477_n2138), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_424J2_126_3477_n2782) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1354 ( .A1(DP_OP_422J2_124_3477_n3019), 
        .A2(DP_OP_424J2_126_3477_n2143), .Y(DP_OP_424J2_126_3477_n2115) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1370 ( .A1(DP_OP_423J2_125_3477_n2051), 
        .A2(n1500), .Y(DP_OP_424J2_126_3477_n2131) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1537 ( .A1(DP_OP_425J2_127_3477_n2710), 
        .A2(DP_OP_423J2_125_3477_n2320), .Y(DP_OP_424J2_126_3477_n2298) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1794 ( .A1(DP_OP_424J2_126_3477_n2579), 
        .A2(DP_OP_422J2_124_3477_n2583), .Y(DP_OP_424J2_126_3477_n2555) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1713 ( .A1(DP_OP_423J2_125_3477_n2666), 
        .A2(n1491), .Y(DP_OP_425J2_127_3477_n2474) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1889 ( .A1(DP_OP_422J2_124_3477_n2270), 
        .A2(n278), .Y(DP_OP_424J2_126_3477_n2650) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1366 ( .A1(DP_OP_424J2_126_3477_n2927), 
        .A2(n1501), .Y(DP_OP_425J2_127_3477_n2127) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1757 ( .A1(DP_OP_425J2_127_3477_n2534), 
        .A2(n1487), .Y(DP_OP_425J2_127_3477_n2518) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1368 ( .A1(DP_OP_425J2_127_3477_n2885), 
        .A2(n1500), .Y(DP_OP_424J2_126_3477_n2129) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1444 ( .A1(DP_OP_425J2_127_3477_n2801), 
        .A2(DP_OP_422J2_124_3477_n2231), .Y(DP_OP_424J2_126_3477_n2205) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1442 ( .A1(DP_OP_423J2_125_3477_n2931), 
        .A2(DP_OP_425J2_127_3477_n2231), .Y(DP_OP_425J2_127_3477_n2203) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1750 ( .A1(DP_OP_424J2_126_3477_n2535), 
        .A2(n772), .Y(DP_OP_424J2_126_3477_n2511) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1317 ( .A1(DP_OP_423J2_125_3477_n2006), 
        .A2(DP_OP_422J2_124_3477_n2100), .Y(DP_OP_424J2_126_3477_n2078) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2058 ( .A1(DP_OP_425J2_127_3477_n2843), 
        .A2(DP_OP_422J2_124_3477_n2847), .Y(DP_OP_425J2_127_3477_n2819) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1669 ( .A1(DP_OP_422J2_124_3477_n2710), 
        .A2(n1488), .Y(DP_OP_424J2_126_3477_n2430) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1669 ( .A1(DP_OP_422J2_124_3477_n2314), 
        .A2(n1488), .Y(DP_OP_425J2_127_3477_n2430) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2058 ( .A1(DP_OP_423J2_125_3477_n2931), 
        .A2(DP_OP_422J2_124_3477_n2847), .Y(DP_OP_424J2_126_3477_n2819) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2285 ( .A1(DP_OP_424J2_126_3477_n3060), 
        .A2(DP_OP_425J2_127_3477_n3066), .Y(DP_OP_424J2_126_3477_n3044) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1317 ( .A1(DP_OP_423J2_125_3477_n3060), 
        .A2(DP_OP_423J2_125_3477_n2100), .Y(DP_OP_425J2_127_3477_n2078) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1750 ( .A1(DP_OP_422J2_124_3477_n2667), 
        .A2(n772), .Y(DP_OP_425J2_127_3477_n2511) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1319 ( .A1(DP_OP_423J2_125_3477_n2008), 
        .A2(DP_OP_423J2_125_3477_n2100), .Y(DP_OP_424J2_126_3477_n2080) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1713 ( .A1(DP_OP_425J2_127_3477_n2534), 
        .A2(n1491), .Y(DP_OP_424J2_126_3477_n2474) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1356 ( .A1(DP_OP_422J2_124_3477_n3021), 
        .A2(DP_OP_424J2_126_3477_n2143), .Y(DP_OP_424J2_126_3477_n2117) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1442 ( .A1(DP_OP_425J2_127_3477_n2799), 
        .A2(DP_OP_422J2_124_3477_n2231), .Y(DP_OP_424J2_126_3477_n2203) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1368 ( .A1(DP_OP_424J2_126_3477_n2929), 
        .A2(n1501), .Y(DP_OP_425J2_127_3477_n2129) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1889 ( .A1(DP_OP_422J2_124_3477_n2798), 
        .A2(n279), .Y(DP_OP_425J2_127_3477_n2650) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1896 ( .A1(DP_OP_422J2_124_3477_n2797), 
        .A2(DP_OP_424J2_126_3477_n2673), .Y(DP_OP_425J2_127_3477_n2657) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1794 ( .A1(DP_OP_425J2_127_3477_n2579), 
        .A2(n671), .Y(DP_OP_425J2_127_3477_n2555) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1757 ( .A1(DP_OP_424J2_126_3477_n2534), 
        .A2(DP_OP_424J2_126_3477_n2540), .Y(DP_OP_424J2_126_3477_n2518) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1537 ( .A1(DP_OP_423J2_125_3477_n2842), 
        .A2(DP_OP_422J2_124_3477_n2320), .Y(DP_OP_425J2_127_3477_n2298) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1354 ( .A1(DP_OP_423J2_125_3477_n3019), 
        .A2(DP_OP_425J2_127_3477_n2143), .Y(DP_OP_425J2_127_3477_n2115) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1632 ( .A1(DP_OP_422J2_124_3477_n2753), 
        .A2(DP_OP_422J2_124_3477_n2409), .Y(DP_OP_424J2_126_3477_n2393) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1672 ( .A1(DP_OP_425J2_127_3477_n2449), 
        .A2(n1488), .Y(DP_OP_425J2_127_3477_n2433) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1635 ( .A1(DP_OP_425J2_127_3477_n2404), 
        .A2(DP_OP_425J2_127_3477_n2409), .Y(DP_OP_425J2_127_3477_n2396) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1899 ( .A1(DP_OP_423J2_125_3477_n2272), 
        .A2(n1), .Y(DP_OP_425J2_127_3477_n2660) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1716 ( .A1(DP_OP_425J2_127_3477_n2493), 
        .A2(n1491), .Y(DP_OP_425J2_127_3477_n2477) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2283 ( .A1(DP_OP_425J2_127_3477_n3058), 
        .A2(DP_OP_425J2_127_3477_n3066), .Y(DP_OP_425J2_127_3477_n3042) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1320 ( .A1(DP_OP_423J2_125_3477_n3063), 
        .A2(DP_OP_422J2_124_3477_n2100), .Y(DP_OP_425J2_127_3477_n2081) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1667 ( .A1(DP_OP_423J2_125_3477_n2708), 
        .A2(n1488), .Y(DP_OP_425J2_127_3477_n2428) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1371 ( .A1(DP_OP_424J2_126_3477_n2932), 
        .A2(n1500), .Y(DP_OP_425J2_127_3477_n2132) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1540 ( .A1(DP_OP_423J2_125_3477_n2845), 
        .A2(DP_OP_423J2_125_3477_n2320), .Y(DP_OP_425J2_127_3477_n2301) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1535 ( .A1(DP_OP_425J2_127_3477_n2312), 
        .A2(DP_OP_425J2_127_3477_n2320), .Y(DP_OP_425J2_127_3477_n2296) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1892 ( .A1(DP_OP_423J2_125_3477_n2273), 
        .A2(n279), .Y(DP_OP_425J2_127_3477_n2653) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1796 ( .A1(DP_OP_425J2_127_3477_n2493), 
        .A2(n670), .Y(DP_OP_424J2_126_3477_n2557) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2236 ( .A1(DP_OP_425J2_127_3477_n2053), 
        .A2(DP_OP_424J2_126_3477_n3023), .Y(DP_OP_424J2_126_3477_n2997) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1583 ( .A1(DP_OP_424J2_126_3477_n2712), 
        .A2(n1386), .Y(DP_OP_425J2_127_3477_n2344) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1898 ( .A1(DP_OP_423J2_125_3477_n2271), 
        .A2(DP_OP_424J2_126_3477_n2673), .Y(DP_OP_425J2_127_3477_n2659) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1810 ( .A1(DP_OP_424J2_126_3477_n2579), 
        .A2(DP_OP_423J2_125_3477_n2585), .Y(DP_OP_424J2_126_3477_n2571) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1810 ( .A1(DP_OP_425J2_127_3477_n2579), 
        .A2(DP_OP_423J2_125_3477_n2585), .Y(DP_OP_425J2_127_3477_n2571) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1891 ( .A1(DP_OP_422J2_124_3477_n2800), 
        .A2(n279), .Y(DP_OP_425J2_127_3477_n2652) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2023 ( .A1(DP_OP_425J2_127_3477_n2800), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_425J2_127_3477_n2784) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1671 ( .A1(DP_OP_425J2_127_3477_n2448), 
        .A2(n1489), .Y(DP_OP_425J2_127_3477_n2432) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2287 ( .A1(DP_OP_425J2_127_3477_n3062), 
        .A2(DP_OP_424J2_126_3477_n3066), .Y(DP_OP_425J2_127_3477_n3046) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1752 ( .A1(DP_OP_422J2_124_3477_n2669), 
        .A2(n772), .Y(DP_OP_425J2_127_3477_n2513) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1759 ( .A1(DP_OP_425J2_127_3477_n2536), 
        .A2(n1486), .Y(DP_OP_425J2_127_3477_n2520) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1796 ( .A1(DP_OP_425J2_127_3477_n2581), 
        .A2(n671), .Y(DP_OP_425J2_127_3477_n2557) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2236 ( .A1(DP_OP_425J2_127_3477_n3021), 
        .A2(DP_OP_422J2_124_3477_n3023), .Y(DP_OP_425J2_127_3477_n2997) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1634 ( .A1(DP_OP_425J2_127_3477_n2403), 
        .A2(DP_OP_423J2_125_3477_n2409), .Y(DP_OP_425J2_127_3477_n2395) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1634 ( .A1(DP_OP_424J2_126_3477_n2403), 
        .A2(DP_OP_423J2_125_3477_n2409), .Y(DP_OP_424J2_126_3477_n2395) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1539 ( .A1(DP_OP_423J2_125_3477_n2844), 
        .A2(DP_OP_422J2_124_3477_n2320), .Y(DP_OP_425J2_127_3477_n2300) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1793 ( .A1(DP_OP_425J2_127_3477_n2578), 
        .A2(n671), .Y(DP_OP_425J2_127_3477_n2554) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1319 ( .A1(DP_OP_423J2_125_3477_n3062), 
        .A2(DP_OP_424J2_126_3477_n2100), .Y(DP_OP_425J2_127_3477_n2080) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1356 ( .A1(DP_OP_424J2_126_3477_n2933), 
        .A2(DP_OP_425J2_127_3477_n2143), .Y(DP_OP_425J2_127_3477_n2117) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1752 ( .A1(DP_OP_422J2_124_3477_n2405), 
        .A2(DP_OP_425J2_127_3477_n2539), .Y(DP_OP_424J2_126_3477_n2513) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1759 ( .A1(DP_OP_422J2_124_3477_n2404), 
        .A2(n1487), .Y(DP_OP_424J2_126_3477_n2520) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1444 ( .A1(DP_OP_423J2_125_3477_n2229), 
        .A2(DP_OP_425J2_127_3477_n2231), .Y(DP_OP_423J2_125_3477_n2205) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1756 ( .A1(DP_OP_423J2_125_3477_n2401), 
        .A2(n1486), .Y(DP_OP_425J2_127_3477_n2517) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1318 ( .A1(DP_OP_424J2_126_3477_n2095), 
        .A2(DP_OP_422J2_124_3477_n2100), .Y(DP_OP_424J2_126_3477_n2079) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1925 ( .A1(DP_OP_422J2_124_3477_n2710), 
        .A2(n1497), .Y(DP_OP_422J2_124_3477_n2686) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1666 ( .A1(DP_OP_424J2_126_3477_n2619), 
        .A2(n1488), .Y(DP_OP_425J2_127_3477_n2427) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1355 ( .A1(DP_OP_425J2_127_3477_n2888), 
        .A2(DP_OP_424J2_126_3477_n2143), .Y(DP_OP_424J2_126_3477_n2116) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1279 ( .A1(DP_OP_422J2_124_3477_n2048), 
        .A2(DP_OP_424J2_126_3477_n2057), .Y(DP_OP_422J2_124_3477_n2040) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1536 ( .A1(DP_OP_423J2_125_3477_n2841), 
        .A2(DP_OP_422J2_124_3477_n2320), .Y(DP_OP_425J2_127_3477_n2297) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1715 ( .A1(DP_OP_422J2_124_3477_n2580), 
        .A2(DP_OP_423J2_125_3477_n2496), .Y(DP_OP_423J2_125_3477_n2476) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2020 ( .A1(DP_OP_422J2_124_3477_n2797), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_422J2_124_3477_n2781) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1282 ( .A1(DP_OP_423J2_125_3477_n2051), 
        .A2(DP_OP_425J2_127_3477_n2057), .Y(DP_OP_423J2_125_3477_n2043) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1356 ( .A1(DP_OP_425J2_127_3477_n2801), 
        .A2(DP_OP_422J2_124_3477_n2143), .Y(DP_OP_423J2_125_3477_n2117) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2233 ( .A1(DP_OP_424J2_126_3477_n2138), 
        .A2(DP_OP_425J2_127_3477_n3023), .Y(DP_OP_422J2_124_3477_n2994) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1319 ( .A1(DP_OP_423J2_125_3477_n2096), 
        .A2(DP_OP_424J2_126_3477_n2100), .Y(DP_OP_423J2_125_3477_n2080) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2023 ( .A1(DP_OP_423J2_125_3477_n2800), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_423J2_125_3477_n2784) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1891 ( .A1(DP_OP_423J2_125_3477_n2668), 
        .A2(n278), .Y(DP_OP_423J2_125_3477_n2652) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1928 ( .A1(DP_OP_423J2_125_3477_n2713), 
        .A2(DP_OP_422J2_124_3477_n2715), .Y(DP_OP_423J2_125_3477_n2689) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1316 ( .A1(DP_OP_423J2_125_3477_n3059), 
        .A2(DP_OP_422J2_124_3477_n2100), .Y(DP_OP_425J2_127_3477_n2077) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1747 ( .A1(DP_OP_423J2_125_3477_n2400), 
        .A2(n772), .Y(DP_OP_425J2_127_3477_n2508) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1320 ( .A1(DP_OP_423J2_125_3477_n2097), 
        .A2(DP_OP_423J2_125_3477_n2100), .Y(DP_OP_423J2_125_3477_n2081) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1352 ( .A1(DP_OP_422J2_124_3477_n2137), 
        .A2(DP_OP_422J2_124_3477_n2143), .Y(DP_OP_422J2_124_3477_n2113) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2287 ( .A1(DP_OP_423J2_125_3477_n3062), 
        .A2(DP_OP_423J2_125_3477_n3066), .Y(DP_OP_423J2_125_3477_n3046) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1790 ( .A1(DP_OP_424J2_126_3477_n2575), 
        .A2(n670), .Y(DP_OP_424J2_126_3477_n2551) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1886 ( .A1(DP_OP_423J2_125_3477_n2267), 
        .A2(n279), .Y(DP_OP_425J2_127_3477_n2647) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2236 ( .A1(DP_OP_423J2_125_3477_n3021), 
        .A2(DP_OP_424J2_126_3477_n3023), .Y(DP_OP_423J2_125_3477_n2997) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1796 ( .A1(DP_OP_423J2_125_3477_n2581), 
        .A2(n670), .Y(DP_OP_423J2_125_3477_n2557) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2018 ( .A1(DP_OP_423J2_125_3477_n2135), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_425J2_127_3477_n2779) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1810 ( .A1(DP_OP_423J2_125_3477_n2579), 
        .A2(DP_OP_423J2_125_3477_n2585), .Y(DP_OP_423J2_125_3477_n2571) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1898 ( .A1(DP_OP_423J2_125_3477_n2667), 
        .A2(n1), .Y(DP_OP_423J2_125_3477_n2659) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1671 ( .A1(DP_OP_423J2_125_3477_n2448), 
        .A2(n1489), .Y(DP_OP_423J2_125_3477_n2432) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1633 ( .A1(DP_OP_422J2_124_3477_n2754), 
        .A2(DP_OP_424J2_126_3477_n2409), .Y(DP_OP_424J2_126_3477_n2394) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1351 ( .A1(DP_OP_424J2_126_3477_n2796), 
        .A2(DP_OP_422J2_124_3477_n2143), .Y(DP_OP_422J2_124_3477_n2112) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1538 ( .A1(DP_OP_424J2_126_3477_n2315), 
        .A2(DP_OP_423J2_125_3477_n2320), .Y(DP_OP_424J2_126_3477_n2299) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1281 ( .A1(DP_OP_425J2_127_3477_n2974), 
        .A2(DP_OP_424J2_126_3477_n2057), .Y(DP_OP_424J2_126_3477_n2042) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1281 ( .A1(DP_OP_424J2_126_3477_n2138), 
        .A2(DP_OP_425J2_127_3477_n2057), .Y(DP_OP_423J2_125_3477_n2042) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1668 ( .A1(DP_OP_422J2_124_3477_n2445), 
        .A2(n1489), .Y(DP_OP_422J2_124_3477_n2429) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1538 ( .A1(DP_OP_423J2_125_3477_n2315), 
        .A2(DP_OP_422J2_124_3477_n2320), .Y(DP_OP_423J2_125_3477_n2299) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1369 ( .A1(DP_OP_424J2_126_3477_n2138), 
        .A2(n1501), .Y(DP_OP_424J2_126_3477_n2130) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1353 ( .A1(DP_OP_425J2_127_3477_n2138), 
        .A2(DP_OP_425J2_127_3477_n2143), .Y(DP_OP_425J2_127_3477_n2114) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1353 ( .A1(DP_OP_422J2_124_3477_n2138), 
        .A2(DP_OP_422J2_124_3477_n2143), .Y(DP_OP_422J2_124_3477_n2114) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1367 ( .A1(DP_OP_425J2_127_3477_n2268), 
        .A2(n1500), .Y(DP_OP_422J2_124_3477_n2128) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1351 ( .A1(DP_OP_422J2_124_3477_n2004), 
        .A2(DP_OP_425J2_127_3477_n2143), .Y(DP_OP_425J2_127_3477_n2112) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1749 ( .A1(DP_OP_422J2_124_3477_n2534), 
        .A2(DP_OP_425J2_127_3477_n2539), .Y(DP_OP_422J2_124_3477_n2510) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1756 ( .A1(DP_OP_422J2_124_3477_n2533), 
        .A2(n1487), .Y(DP_OP_422J2_124_3477_n2517) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1536 ( .A1(DP_OP_422J2_124_3477_n2313), 
        .A2(DP_OP_423J2_125_3477_n2320), .Y(DP_OP_422J2_124_3477_n2297) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1316 ( .A1(DP_OP_422J2_124_3477_n2093), 
        .A2(DP_OP_423J2_125_3477_n2100), .Y(DP_OP_422J2_124_3477_n2077) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1441 ( .A1(DP_OP_423J2_125_3477_n2798), 
        .A2(DP_OP_422J2_124_3477_n2231), .Y(DP_OP_422J2_124_3477_n2202) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1367 ( .A1(DP_OP_424J2_126_3477_n2928), 
        .A2(n1500), .Y(DP_OP_425J2_127_3477_n2128) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1895 ( .A1(DP_OP_422J2_124_3477_n2664), 
        .A2(n1), .Y(DP_OP_422J2_124_3477_n2656) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1751 ( .A1(DP_OP_422J2_124_3477_n2404), 
        .A2(n772), .Y(DP_OP_424J2_126_3477_n2512) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1670 ( .A1(DP_OP_424J2_126_3477_n2447), 
        .A2(DP_OP_423J2_125_3477_n2452), .Y(DP_OP_424J2_126_3477_n2431) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1539 ( .A1(DP_OP_423J2_125_3477_n2316), 
        .A2(DP_OP_423J2_125_3477_n2320), .Y(DP_OP_423J2_125_3477_n2300) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1807 ( .A1(DP_OP_422J2_124_3477_n2576), 
        .A2(DP_OP_422J2_124_3477_n2585), .Y(DP_OP_422J2_124_3477_n2568) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1749 ( .A1(DP_OP_425J2_127_3477_n2534), 
        .A2(n772), .Y(DP_OP_425J2_127_3477_n2510) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1323 ( .A1(DP_OP_422J2_124_3477_n2092), 
        .A2(n621), .Y(DP_OP_422J2_124_3477_n2084) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1888 ( .A1(DP_OP_422J2_124_3477_n2665), 
        .A2(n278), .Y(DP_OP_422J2_124_3477_n2649) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1844 ( .A1(DP_OP_422J2_124_3477_n2621), 
        .A2(n1498), .Y(DP_OP_422J2_124_3477_n2605) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1441 ( .A1(DP_OP_425J2_127_3477_n2226), 
        .A2(DP_OP_425J2_127_3477_n2231), .Y(DP_OP_425J2_127_3477_n2202) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1443 ( .A1(DP_OP_425J2_127_3477_n2800), 
        .A2(DP_OP_425J2_127_3477_n2231), .Y(DP_OP_424J2_126_3477_n2204) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1897 ( .A1(DP_OP_423J2_125_3477_n2666), 
        .A2(n1), .Y(DP_OP_423J2_125_3477_n2658) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1895 ( .A1(DP_OP_423J2_125_3477_n2268), 
        .A2(DP_OP_422J2_124_3477_n2673), .Y(DP_OP_425J2_127_3477_n2656) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1758 ( .A1(DP_OP_424J2_126_3477_n2535), 
        .A2(n1486), .Y(DP_OP_424J2_126_3477_n2519) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1355 ( .A1(DP_OP_423J2_125_3477_n2140), 
        .A2(DP_OP_424J2_126_3477_n2143), .Y(DP_OP_423J2_125_3477_n2116) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1318 ( .A1(DP_OP_425J2_127_3477_n2843), 
        .A2(DP_OP_422J2_124_3477_n2100), .Y(DP_OP_423J2_125_3477_n2079) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1325 ( .A1(DP_OP_423J2_125_3477_n2094), 
        .A2(n621), .Y(DP_OP_423J2_125_3477_n2086) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1369 ( .A1(DP_OP_425J2_127_3477_n2798), 
        .A2(n1500), .Y(DP_OP_423J2_125_3477_n2130) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1809 ( .A1(DP_OP_422J2_124_3477_n2446), 
        .A2(DP_OP_423J2_125_3477_n2585), .Y(DP_OP_423J2_125_3477_n2570) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1670 ( .A1(DP_OP_423J2_125_3477_n2447), 
        .A2(n1488), .Y(DP_OP_423J2_125_3477_n2431) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1751 ( .A1(DP_OP_423J2_125_3477_n2536), 
        .A2(n772), .Y(DP_OP_423J2_125_3477_n2512) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1714 ( .A1(DP_OP_422J2_124_3477_n2579), 
        .A2(DP_OP_423J2_125_3477_n2496), .Y(DP_OP_423J2_125_3477_n2475) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2286 ( .A1(DP_OP_425J2_127_3477_n2007), 
        .A2(DP_OP_423J2_125_3477_n3066), .Y(DP_OP_424J2_126_3477_n3045) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1582 ( .A1(DP_OP_422J2_124_3477_n2799), 
        .A2(n1386), .Y(DP_OP_424J2_126_3477_n2343) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1892 ( .A1(DP_OP_423J2_125_3477_n2669), 
        .A2(n279), .Y(DP_OP_423J2_125_3477_n2653) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1352 ( .A1(DP_OP_425J2_127_3477_n2885), 
        .A2(DP_OP_424J2_126_3477_n2143), .Y(DP_OP_424J2_126_3477_n2113) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1811 ( .A1(DP_OP_422J2_124_3477_n2448), 
        .A2(DP_OP_424J2_126_3477_n2585), .Y(DP_OP_423J2_125_3477_n2572) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1712 ( .A1(DP_OP_423J2_125_3477_n2665), 
        .A2(n1491), .Y(DP_OP_425J2_127_3477_n2473) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2059 ( .A1(DP_OP_423J2_125_3477_n2932), 
        .A2(DP_OP_422J2_124_3477_n2847), .Y(DP_OP_424J2_126_3477_n2820) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1323 ( .A1(DP_OP_425J2_127_3477_n2092), 
        .A2(n621), .Y(DP_OP_425J2_127_3477_n2084) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1795 ( .A1(DP_OP_424J2_126_3477_n2580), 
        .A2(n671), .Y(DP_OP_424J2_126_3477_n2556) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2286 ( .A1(DP_OP_423J2_125_3477_n3061), 
        .A2(DP_OP_425J2_127_3477_n3066), .Y(DP_OP_423J2_125_3477_n3045) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1890 ( .A1(DP_OP_424J2_126_3477_n2667), 
        .A2(n279), .Y(DP_OP_424J2_126_3477_n2651) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1443 ( .A1(DP_OP_423J2_125_3477_n2228), 
        .A2(DP_OP_422J2_124_3477_n2231), .Y(DP_OP_423J2_125_3477_n2204) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1812 ( .A1(DP_OP_425J2_127_3477_n2493), 
        .A2(DP_OP_424J2_126_3477_n2585), .Y(DP_OP_424J2_126_3477_n2573) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2235 ( .A1(DP_OP_424J2_126_3477_n2932), 
        .A2(DP_OP_422J2_124_3477_n3023), .Y(DP_OP_423J2_125_3477_n2996) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1890 ( .A1(DP_OP_423J2_125_3477_n2667), 
        .A2(n279), .Y(DP_OP_423J2_125_3477_n2651) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1922 ( .A1(DP_OP_422J2_124_3477_n2707), 
        .A2(DP_OP_422J2_124_3477_n2715), .Y(DP_OP_422J2_124_3477_n2683) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1758 ( .A1(DP_OP_422J2_124_3477_n2491), 
        .A2(DP_OP_424J2_126_3477_n2540), .Y(DP_OP_423J2_125_3477_n2519) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2230 ( .A1(DP_OP_422J2_124_3477_n3015), 
        .A2(DP_OP_425J2_127_3477_n3023), .Y(DP_OP_422J2_124_3477_n2991) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1790 ( .A1(DP_OP_422J2_124_3477_n2575), 
        .A2(n671), .Y(DP_OP_422J2_124_3477_n2551) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1888 ( .A1(DP_OP_423J2_125_3477_n2269), 
        .A2(n279), .Y(DP_OP_425J2_127_3477_n2649) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1795 ( .A1(DP_OP_422J2_124_3477_n2448), 
        .A2(n671), .Y(DP_OP_423J2_125_3477_n2556) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1438 ( .A1(DP_OP_422J2_124_3477_n2223), 
        .A2(DP_OP_424J2_126_3477_n2231), .Y(DP_OP_422J2_124_3477_n2199) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1668 ( .A1(DP_OP_425J2_127_3477_n2445), 
        .A2(DP_OP_423J2_125_3477_n2452), .Y(DP_OP_425J2_127_3477_n2429) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1147 ( .A1(n1328), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_423J2_125_3477_n306) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1175 ( .A1(n1293), .A2(n1508), .Y(
        DP_OP_423J2_125_3477_n1936) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1922 ( .A1(DP_OP_424J2_126_3477_n2619), 
        .A2(DP_OP_422J2_124_3477_n2715), .Y(DP_OP_423J2_125_3477_n2683) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1175 ( .A1(n1869), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_422J2_124_3477_n1936) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1145 ( .A1(n1912), .A2(n1508), .Y(
        DP_OP_422J2_124_3477_n302) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1153 ( .A1(n1887), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_422J2_124_3477_n318) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1152 ( .A1(n1902), .A2(
        DP_OP_422J2_124_3477_n2), .Y(DP_OP_422J2_124_3477_n316) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1149 ( .A1(n1889), .A2(n1508), .Y(
        DP_OP_422J2_124_3477_n310) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1157 ( .A1(n1885), .A2(n1508), .Y(
        DP_OP_422J2_124_3477_n326) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1164 ( .A1(n1973), .A2(n1508), .Y(
        DP_OP_422J2_124_3477_n1926) );
  AND2X1_HVT DP_OP_423J2_125_3477_U184 ( .A1(DP_OP_423J2_125_3477_n284), .A2(
        DP_OP_423J2_125_3477_n174), .Y(DP_OP_423J2_125_3477_n20) );
  AND2X1_HVT DP_OP_423J2_125_3477_U160 ( .A1(DP_OP_423J2_125_3477_n282), .A2(
        DP_OP_423J2_125_3477_n156), .Y(DP_OP_423J2_125_3477_n18) );
  AND2X1_HVT DP_OP_423J2_125_3477_U134 ( .A1(DP_OP_423J2_125_3477_n280), .A2(
        DP_OP_423J2_125_3477_n136), .Y(DP_OP_423J2_125_3477_n16) );
  AND2X1_HVT DP_OP_423J2_125_3477_U94 ( .A1(DP_OP_423J2_125_3477_n277), .A2(
        DP_OP_423J2_125_3477_n105), .Y(DP_OP_423J2_125_3477_n13) );
  AND2X1_HVT DP_OP_423J2_125_3477_U18 ( .A1(n1670), .A2(
        DP_OP_423J2_125_3477_n47), .Y(DP_OP_423J2_125_3477_n7) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U56 ( .A1(DP_OP_424J2_126_3477_n77), .A2(
        DP_OP_424J2_126_3477_n82), .Y(DP_OP_424J2_126_3477_n75) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U56 ( .A1(DP_OP_423J2_125_3477_n77), .A2(
        DP_OP_423J2_125_3477_n82), .Y(DP_OP_423J2_125_3477_n75) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U106 ( .A1(DP_OP_425J2_127_3477_n115), .A2(
        DP_OP_425J2_127_3477_n144), .Y(DP_OP_425J2_127_3477_n111) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U56 ( .A1(DP_OP_425J2_127_3477_n77), .A2(
        DP_OP_425J2_127_3477_n82), .Y(DP_OP_425J2_127_3477_n75) );
  AND2X1_HVT DP_OP_423J2_125_3477_U26 ( .A1(DP_OP_423J2_125_3477_n272), .A2(
        DP_OP_423J2_125_3477_n52), .Y(DP_OP_423J2_125_3477_n8) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U56 ( .A1(DP_OP_422J2_124_3477_n77), .A2(
        DP_OP_422J2_124_3477_n82), .Y(DP_OP_422J2_124_3477_n75) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U52 ( .A1(DP_OP_424J2_126_3477_n73), .A2(
        DP_OP_424J2_126_3477_n182), .Y(DP_OP_424J2_126_3477_n71) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U52 ( .A1(DP_OP_423J2_125_3477_n73), .A2(
        DP_OP_423J2_125_3477_n182), .Y(DP_OP_423J2_125_3477_n71) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U52 ( .A1(DP_OP_425J2_127_3477_n73), .A2(
        DP_OP_425J2_127_3477_n182), .Y(DP_OP_425J2_127_3477_n71) );
  AND2X1_HVT DP_OP_423J2_125_3477_U198 ( .A1(DP_OP_423J2_125_3477_n285), .A2(
        DP_OP_423J2_125_3477_n185), .Y(DP_OP_423J2_125_3477_n21) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U224 ( .A1(DP_OP_424J2_126_3477_n335), .A2(
        DP_OP_424J2_126_3477_n340), .Y(DP_OP_424J2_126_3477_n202) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U36 ( .A1(DP_OP_424J2_126_3477_n60), .A2(
        DP_OP_424J2_126_3477_n197), .Y(DP_OP_424J2_126_3477_n58) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U36 ( .A1(DP_OP_423J2_125_3477_n60), .A2(
        DP_OP_423J2_125_3477_n197), .Y(DP_OP_423J2_125_3477_n58) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U36 ( .A1(DP_OP_425J2_127_3477_n60), .A2(
        DP_OP_425J2_127_3477_n197), .Y(DP_OP_425J2_127_3477_n58) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U224 ( .A1(DP_OP_425J2_127_3477_n335), .A2(
        DP_OP_425J2_127_3477_n340), .Y(DP_OP_425J2_127_3477_n202) );
  AND2X1_HVT DP_OP_423J2_125_3477_U214 ( .A1(DP_OP_423J2_125_3477_n286), .A2(
        DP_OP_423J2_125_3477_n198), .Y(DP_OP_423J2_125_3477_n22) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U36 ( .A1(DP_OP_422J2_124_3477_n60), .A2(
        DP_OP_422J2_124_3477_n197), .Y(DP_OP_422J2_124_3477_n58) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U195 ( .A1(DP_OP_423J2_125_3477_n182), .A2(
        DP_OP_423J2_125_3477_n190), .A3(DP_OP_423J2_125_3477_n185), .Y(
        DP_OP_423J2_125_3477_n177) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U48 ( .A1(DP_OP_423J2_125_3477_n69), .A2(
        DP_OP_423J2_125_3477_n189), .Y(DP_OP_423J2_125_3477_n67) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U25 ( .A1(DP_OP_423J2_125_3477_n51), .A2(
        DP_OP_423J2_125_3477_n57), .A3(DP_OP_423J2_125_3477_n52), .Y(
        DP_OP_423J2_125_3477_n50) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U24 ( .A1(DP_OP_423J2_125_3477_n51), .A2(
        DP_OP_423J2_125_3477_n56), .Y(DP_OP_423J2_125_3477_n49) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U24 ( .A1(DP_OP_425J2_127_3477_n51), .A2(
        DP_OP_425J2_127_3477_n56), .Y(DP_OP_425J2_127_3477_n49) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U25 ( .A1(DP_OP_425J2_127_3477_n51), .A2(
        DP_OP_425J2_127_3477_n57), .A3(DP_OP_425J2_127_3477_n52), .Y(
        DP_OP_425J2_127_3477_n50) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U48 ( .A1(DP_OP_425J2_127_3477_n69), .A2(
        DP_OP_425J2_127_3477_n189), .Y(DP_OP_425J2_127_3477_n67) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U24 ( .A1(DP_OP_424J2_126_3477_n51), .A2(
        DP_OP_424J2_126_3477_n56), .Y(DP_OP_424J2_126_3477_n49) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U48 ( .A1(DP_OP_424J2_126_3477_n69), .A2(
        DP_OP_424J2_126_3477_n189), .Y(DP_OP_424J2_126_3477_n67) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U25 ( .A1(DP_OP_424J2_126_3477_n51), .A2(
        DP_OP_424J2_126_3477_n57), .A3(DP_OP_424J2_126_3477_n52), .Y(
        DP_OP_424J2_126_3477_n50) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U195 ( .A1(DP_OP_422J2_124_3477_n182), .A2(
        DP_OP_422J2_124_3477_n190), .A3(DP_OP_422J2_124_3477_n185), .Y(
        DP_OP_422J2_124_3477_n177) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U25 ( .A1(DP_OP_422J2_124_3477_n51), .A2(
        DP_OP_422J2_124_3477_n57), .A3(DP_OP_422J2_124_3477_n52), .Y(
        DP_OP_422J2_124_3477_n50) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U24 ( .A1(DP_OP_422J2_124_3477_n51), .A2(
        DP_OP_422J2_124_3477_n56), .Y(DP_OP_422J2_124_3477_n49) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U48 ( .A1(DP_OP_422J2_124_3477_n69), .A2(
        DP_OP_422J2_124_3477_n189), .Y(DP_OP_422J2_124_3477_n67) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U65 ( .A1(DP_OP_423J2_125_3477_n82), .A2(
        DP_OP_423J2_125_3477_n110), .A3(DP_OP_423J2_125_3477_n85), .Y(
        DP_OP_423J2_125_3477_n81) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U156 ( .A1(DP_OP_423J2_125_3477_n153), .A2(
        DP_OP_423J2_125_3477_n160), .Y(DP_OP_423J2_125_3477_n151) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U64 ( .A1(DP_OP_423J2_125_3477_n82), .A2(
        DP_OP_423J2_125_3477_n109), .Y(DP_OP_423J2_125_3477_n80) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U91 ( .A1(DP_OP_423J2_125_3477_n102), .A2(
        DP_OP_423J2_125_3477_n110), .A3(DP_OP_423J2_125_3477_n105), .Y(
        DP_OP_423J2_125_3477_n101) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U90 ( .A1(DP_OP_423J2_125_3477_n102), .A2(
        DP_OP_423J2_125_3477_n109), .Y(DP_OP_423J2_125_3477_n100) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U78 ( .A1(DP_OP_423J2_125_3477_n93), .A2(
        DP_OP_423J2_125_3477_n109), .Y(DP_OP_423J2_125_3477_n91) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U79 ( .A1(DP_OP_423J2_125_3477_n93), .A2(
        DP_OP_423J2_125_3477_n110), .A3(DP_OP_423J2_125_3477_n94), .Y(
        DP_OP_423J2_125_3477_n92) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U118 ( .A1(DP_OP_423J2_125_3477_n124), .A2(
        DP_OP_423J2_125_3477_n140), .Y(DP_OP_423J2_125_3477_n122) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U130 ( .A1(DP_OP_423J2_125_3477_n133), .A2(
        DP_OP_423J2_125_3477_n140), .Y(DP_OP_423J2_125_3477_n131) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U78 ( .A1(DP_OP_422J2_124_3477_n93), .A2(
        DP_OP_422J2_124_3477_n109), .Y(DP_OP_422J2_124_3477_n91) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U118 ( .A1(DP_OP_422J2_124_3477_n124), .A2(
        DP_OP_422J2_124_3477_n140), .Y(DP_OP_422J2_124_3477_n122) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U156 ( .A1(DP_OP_424J2_126_3477_n153), .A2(
        DP_OP_424J2_126_3477_n160), .Y(DP_OP_424J2_126_3477_n151) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U130 ( .A1(DP_OP_422J2_124_3477_n133), .A2(
        DP_OP_422J2_124_3477_n140), .Y(DP_OP_422J2_124_3477_n131) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U90 ( .A1(DP_OP_422J2_124_3477_n102), .A2(
        DP_OP_422J2_124_3477_n109), .Y(DP_OP_422J2_124_3477_n100) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U157 ( .A1(DP_OP_422J2_124_3477_n153), .A2(
        DP_OP_422J2_124_3477_n161), .A3(DP_OP_422J2_124_3477_n156), .Y(
        DP_OP_422J2_124_3477_n152) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U64 ( .A1(DP_OP_422J2_124_3477_n82), .A2(
        DP_OP_422J2_124_3477_n109), .Y(DP_OP_422J2_124_3477_n80) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U130 ( .A1(DP_OP_424J2_126_3477_n133), .A2(
        DP_OP_424J2_126_3477_n140), .Y(DP_OP_424J2_126_3477_n131) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U156 ( .A1(DP_OP_422J2_124_3477_n153), .A2(
        DP_OP_422J2_124_3477_n160), .Y(DP_OP_422J2_124_3477_n151) );
  OAI21X1_HVT DP_OP_422J2_124_3477_U181 ( .A1(DP_OP_422J2_124_3477_n171), .A2(
        DP_OP_422J2_124_3477_n179), .A3(DP_OP_422J2_124_3477_n174), .Y(
        DP_OP_422J2_124_3477_n170) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U64 ( .A1(DP_OP_425J2_127_3477_n82), .A2(
        DP_OP_425J2_127_3477_n109), .Y(DP_OP_425J2_127_3477_n80) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U78 ( .A1(DP_OP_425J2_127_3477_n93), .A2(
        DP_OP_425J2_127_3477_n109), .Y(DP_OP_425J2_127_3477_n91) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U156 ( .A1(DP_OP_425J2_127_3477_n153), .A2(
        DP_OP_425J2_127_3477_n160), .Y(DP_OP_425J2_127_3477_n151) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U90 ( .A1(DP_OP_425J2_127_3477_n102), .A2(
        DP_OP_425J2_127_3477_n109), .Y(DP_OP_425J2_127_3477_n100) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U130 ( .A1(DP_OP_425J2_127_3477_n133), .A2(
        DP_OP_425J2_127_3477_n140), .Y(DP_OP_425J2_127_3477_n131) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U118 ( .A1(DP_OP_425J2_127_3477_n124), .A2(
        DP_OP_425J2_127_3477_n140), .Y(DP_OP_425J2_127_3477_n122) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U78 ( .A1(DP_OP_424J2_126_3477_n93), .A2(
        DP_OP_424J2_126_3477_n109), .Y(DP_OP_424J2_126_3477_n91) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U90 ( .A1(DP_OP_424J2_126_3477_n102), .A2(
        DP_OP_424J2_126_3477_n109), .Y(DP_OP_424J2_126_3477_n100) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U118 ( .A1(DP_OP_424J2_126_3477_n124), .A2(
        DP_OP_424J2_126_3477_n140), .Y(DP_OP_424J2_126_3477_n122) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U64 ( .A1(DP_OP_424J2_126_3477_n82), .A2(
        DP_OP_424J2_126_3477_n109), .Y(DP_OP_424J2_126_3477_n80) );
  OAI21X1_HVT DP_OP_424J2_126_3477_U131 ( .A1(DP_OP_424J2_126_3477_n133), .A2(
        DP_OP_424J2_126_3477_n141), .A3(DP_OP_424J2_126_3477_n136), .Y(
        DP_OP_424J2_126_3477_n132) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U238 ( .A1(DP_OP_423J2_125_3477_n214), .A2(
        n1522), .Y(DP_OP_423J2_125_3477_n212) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U131 ( .A1(DP_OP_425J2_127_3477_n133), .A2(
        DP_OP_425J2_127_3477_n141), .A3(DP_OP_425J2_127_3477_n136), .Y(
        DP_OP_425J2_127_3477_n132) );
  OAI21X1_HVT DP_OP_425J2_127_3477_U91 ( .A1(DP_OP_425J2_127_3477_n102), .A2(
        DP_OP_425J2_127_3477_n110), .A3(DP_OP_425J2_127_3477_n105), .Y(
        DP_OP_425J2_127_3477_n101) );
  OAI21X1_HVT DP_OP_423J2_125_3477_U239 ( .A1(DP_OP_423J2_125_3477_n214), .A2(
        DP_OP_423J2_125_3477_n222), .A3(DP_OP_423J2_125_3477_n217), .Y(
        DP_OP_423J2_125_3477_n213) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2015 ( .A1(DP_OP_425J2_127_3477_n2272), 
        .A2(n1444), .Y(DP_OP_424J2_126_3477_n2776) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1983 ( .A1(DP_OP_424J2_126_3477_n2268), 
        .A2(n66), .Y(DP_OP_425J2_127_3477_n2744) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2274 ( .A1(DP_OP_422J2_124_3477_n3057), 
        .A2(DP_OP_424J2_126_3477_n3065), .Y(DP_OP_422J2_124_3477_n3033) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1218 ( .A1(DP_OP_422J2_124_3477_n2003), 
        .A2(DP_OP_422J2_124_3477_n2011), .Y(DP_OP_422J2_124_3477_n1979) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1262 ( .A1(DP_OP_422J2_124_3477_n2047), 
        .A2(DP_OP_422J2_124_3477_n2055), .Y(DP_OP_422J2_124_3477_n2023) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2011 ( .A1(DP_OP_422J2_124_3477_n2224), 
        .A2(DP_OP_422J2_124_3477_n2803), .Y(DP_OP_423J2_125_3477_n2772) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1402 ( .A1(DP_OP_424J2_126_3477_n2883), 
        .A2(DP_OP_425J2_127_3477_n2188), .Y(DP_OP_425J2_127_3477_n2163) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1490 ( .A1(DP_OP_422J2_124_3477_n2135), 
        .A2(DP_OP_422J2_124_3477_n2276), .Y(DP_OP_425J2_127_3477_n2251) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1402 ( .A1(DP_OP_422J2_124_3477_n2883), 
        .A2(n1343), .Y(DP_OP_423J2_125_3477_n2163) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1446 ( .A1(DP_OP_424J2_126_3477_n2311), 
        .A2(n364), .Y(DP_OP_423J2_125_3477_n2207) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2015 ( .A1(DP_OP_425J2_127_3477_n2800), 
        .A2(DP_OP_422J2_124_3477_n2803), .Y(DP_OP_425J2_127_3477_n2776) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1226 ( .A1(DP_OP_424J2_126_3477_n3057), 
        .A2(n558), .Y(DP_OP_425J2_127_3477_n1987) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2274 ( .A1(DP_OP_424J2_126_3477_n3057), 
        .A2(DP_OP_424J2_126_3477_n3065), .Y(DP_OP_424J2_126_3477_n3033) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1218 ( .A1(DP_OP_424J2_126_3477_n2003), 
        .A2(DP_OP_424J2_126_3477_n2011), .Y(DP_OP_424J2_126_3477_n1979) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2029 ( .A1(DP_OP_423J2_125_3477_n2798), 
        .A2(DP_OP_423J2_125_3477_n2805), .Y(DP_OP_423J2_125_3477_n2790) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2012 ( .A1(DP_OP_422J2_124_3477_n2225), 
        .A2(DP_OP_423J2_125_3477_n2803), .Y(DP_OP_423J2_125_3477_n2773) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2246 ( .A1(DP_OP_424J2_126_3477_n2003), 
        .A2(DP_OP_425J2_127_3477_n3025), .Y(DP_OP_425J2_127_3477_n3007) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1447 ( .A1(DP_OP_422J2_124_3477_n2092), 
        .A2(n365), .Y(DP_OP_425J2_127_3477_n2208) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1498 ( .A1(DP_OP_424J2_126_3477_n2795), 
        .A2(DP_OP_423J2_125_3477_n2277), .Y(DP_OP_425J2_127_3477_n2259) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U2246 ( .A1(DP_OP_424J2_126_3477_n2927), 
        .A2(DP_OP_423J2_125_3477_n3025), .Y(DP_OP_423J2_125_3477_n3007) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1491 ( .A1(DP_OP_423J2_125_3477_n2268), 
        .A2(DP_OP_423J2_125_3477_n2276), .Y(DP_OP_423J2_125_3477_n2252) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2014 ( .A1(DP_OP_423J2_125_3477_n2799), 
        .A2(DP_OP_423J2_125_3477_n2803), .Y(DP_OP_423J2_125_3477_n2775) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2031 ( .A1(DP_OP_423J2_125_3477_n2800), 
        .A2(DP_OP_423J2_125_3477_n2805), .Y(DP_OP_423J2_125_3477_n2792) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1850 ( .A1(DP_OP_423J2_125_3477_n2311), 
        .A2(DP_OP_422J2_124_3477_n2629), .Y(DP_OP_425J2_127_3477_n2611) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2028 ( .A1(DP_OP_425J2_127_3477_n2357), 
        .A2(DP_OP_423J2_125_3477_n2805), .Y(DP_OP_423J2_125_3477_n2789) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1938 ( .A1(DP_OP_422J2_124_3477_n2839), 
        .A2(n597), .Y(DP_OP_425J2_127_3477_n2699) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2032 ( .A1(DP_OP_423J2_125_3477_n2801), 
        .A2(DP_OP_423J2_125_3477_n2805), .Y(DP_OP_423J2_125_3477_n2793) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U2114 ( .A1(DP_OP_425J2_127_3477_n2883), 
        .A2(DP_OP_425J2_127_3477_n2893), .Y(DP_OP_425J2_127_3477_n2875) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2063 ( .A1(DP_OP_425J2_127_3477_n2840), 
        .A2(DP_OP_425J2_127_3477_n2848), .Y(DP_OP_425J2_127_3477_n2824) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1984 ( .A1(DP_OP_422J2_124_3477_n2753), 
        .A2(n66), .Y(DP_OP_422J2_124_3477_n2745) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1218 ( .A1(DP_OP_423J2_125_3477_n2003), 
        .A2(DP_OP_425J2_127_3477_n2011), .Y(DP_OP_423J2_125_3477_n1979) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1834 ( .A1(DP_OP_423J2_125_3477_n2619), 
        .A2(DP_OP_423J2_125_3477_n2627), .Y(DP_OP_423J2_125_3477_n2595) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U2150 ( .A1(DP_OP_424J2_126_3477_n2927), 
        .A2(DP_OP_424J2_126_3477_n2936), .Y(DP_OP_424J2_126_3477_n2911) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2014 ( .A1(DP_OP_422J2_124_3477_n2799), 
        .A2(n1444), .Y(DP_OP_422J2_124_3477_n2775) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1974 ( .A1(DP_OP_422J2_124_3477_n2179), 
        .A2(DP_OP_425J2_127_3477_n2760), .Y(DP_OP_424J2_126_3477_n2735) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1798 ( .A1(DP_OP_422J2_124_3477_n2575), 
        .A2(n186), .Y(DP_OP_422J2_124_3477_n2559) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2028 ( .A1(DP_OP_422J2_124_3477_n2797), 
        .A2(DP_OP_422J2_124_3477_n2805), .Y(DP_OP_422J2_124_3477_n2789) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1491 ( .A1(DP_OP_422J2_124_3477_n2268), 
        .A2(DP_OP_422J2_124_3477_n2276), .Y(DP_OP_422J2_124_3477_n2252) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1498 ( .A1(DP_OP_422J2_124_3477_n2267), 
        .A2(DP_OP_422J2_124_3477_n2277), .Y(DP_OP_422J2_124_3477_n2259) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1226 ( .A1(DP_OP_424J2_126_3477_n2003), 
        .A2(n558), .Y(DP_OP_424J2_126_3477_n1987) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2026 ( .A1(DP_OP_422J2_124_3477_n2795), 
        .A2(DP_OP_422J2_124_3477_n2805), .Y(DP_OP_422J2_124_3477_n2787) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1542 ( .A1(DP_OP_422J2_124_3477_n2311), 
        .A2(DP_OP_422J2_124_3477_n2321), .Y(DP_OP_422J2_124_3477_n2303) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2032 ( .A1(DP_OP_422J2_124_3477_n2801), 
        .A2(DP_OP_422J2_124_3477_n2805), .Y(DP_OP_422J2_124_3477_n2793) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2160 ( .A1(DP_OP_422J2_124_3477_n2929), 
        .A2(n446), .Y(DP_OP_422J2_124_3477_n2921) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1446 ( .A1(DP_OP_422J2_124_3477_n2927), 
        .A2(n365), .Y(DP_OP_424J2_126_3477_n2207) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1218 ( .A1(DP_OP_424J2_126_3477_n3057), 
        .A2(DP_OP_425J2_127_3477_n2011), .Y(DP_OP_425J2_127_3477_n1979) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1490 ( .A1(DP_OP_424J2_126_3477_n2267), 
        .A2(DP_OP_424J2_126_3477_n2276), .Y(DP_OP_424J2_126_3477_n2251) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2274 ( .A1(DP_OP_425J2_127_3477_n3057), 
        .A2(DP_OP_425J2_127_3477_n3065), .Y(DP_OP_425J2_127_3477_n3033) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1402 ( .A1(DP_OP_422J2_124_3477_n2971), 
        .A2(n1344), .Y(DP_OP_424J2_126_3477_n2163) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1834 ( .A1(DP_OP_423J2_125_3477_n2311), 
        .A2(DP_OP_424J2_126_3477_n2627), .Y(DP_OP_425J2_127_3477_n2595) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2029 ( .A1(DP_OP_422J2_124_3477_n2798), 
        .A2(DP_OP_422J2_124_3477_n2805), .Y(DP_OP_422J2_124_3477_n2790) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1623 ( .A1(DP_OP_424J2_126_3477_n2532), 
        .A2(n1333), .Y(DP_OP_422J2_124_3477_n2384) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1798 ( .A1(DP_OP_424J2_126_3477_n2575), 
        .A2(n186), .Y(DP_OP_424J2_126_3477_n2559) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2159 ( .A1(DP_OP_422J2_124_3477_n2928), 
        .A2(n445), .Y(DP_OP_422J2_124_3477_n2920) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2159 ( .A1(DP_OP_424J2_126_3477_n2928), 
        .A2(n444), .Y(DP_OP_424J2_126_3477_n2920) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2027 ( .A1(DP_OP_422J2_124_3477_n2796), 
        .A2(DP_OP_422J2_124_3477_n2805), .Y(DP_OP_422J2_124_3477_n2788) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2016 ( .A1(DP_OP_422J2_124_3477_n2801), 
        .A2(DP_OP_423J2_125_3477_n2803), .Y(DP_OP_422J2_124_3477_n2777) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2159 ( .A1(DP_OP_424J2_126_3477_n2092), 
        .A2(n445), .Y(DP_OP_425J2_127_3477_n2920) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2030 ( .A1(DP_OP_422J2_124_3477_n2799), 
        .A2(DP_OP_422J2_124_3477_n2805), .Y(DP_OP_422J2_124_3477_n2791) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2027 ( .A1(DP_OP_422J2_124_3477_n2224), 
        .A2(DP_OP_423J2_125_3477_n2805), .Y(DP_OP_423J2_125_3477_n2788) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2159 ( .A1(DP_OP_422J2_124_3477_n2092), 
        .A2(n445), .Y(DP_OP_423J2_125_3477_n2920) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1623 ( .A1(DP_OP_424J2_126_3477_n2400), 
        .A2(n1346), .Y(DP_OP_424J2_126_3477_n2384) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1492 ( .A1(DP_OP_423J2_125_3477_n2269), 
        .A2(DP_OP_423J2_125_3477_n2276), .Y(DP_OP_423J2_125_3477_n2253) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1807 ( .A1(DP_OP_425J2_127_3477_n2576), 
        .A2(DP_OP_424J2_126_3477_n2585), .Y(DP_OP_425J2_127_3477_n2568) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1632 ( .A1(DP_OP_422J2_124_3477_n2401), 
        .A2(DP_OP_425J2_127_3477_n2409), .Y(DP_OP_422J2_124_3477_n2393) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1807 ( .A1(DP_OP_424J2_126_3477_n2576), 
        .A2(DP_OP_424J2_126_3477_n2585), .Y(DP_OP_424J2_126_3477_n2568) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1718 ( .A1(DP_OP_423J2_125_3477_n2399), 
        .A2(DP_OP_425J2_127_3477_n2497), .Y(DP_OP_424J2_126_3477_n2479) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2057 ( .A1(DP_OP_423J2_125_3477_n2094), 
        .A2(n1438), .Y(DP_OP_425J2_127_3477_n2818) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2202 ( .A1(DP_OP_424J2_126_3477_n2971), 
        .A2(n677), .Y(DP_OP_424J2_126_3477_n2963) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2055 ( .A1(DP_OP_425J2_127_3477_n2840), 
        .A2(n1438), .Y(DP_OP_425J2_127_3477_n2816) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2283 ( .A1(DP_OP_424J2_126_3477_n3058), 
        .A2(DP_OP_425J2_127_3477_n3066), .Y(DP_OP_424J2_126_3477_n3042) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1270 ( .A1(DP_OP_424J2_126_3477_n3015), 
        .A2(DP_OP_425J2_127_3477_n2056), .Y(DP_OP_425J2_127_3477_n2031) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1712 ( .A1(DP_OP_422J2_124_3477_n2577), 
        .A2(DP_OP_423J2_125_3477_n2496), .Y(DP_OP_423J2_125_3477_n2473) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1455 ( .A1(DP_OP_425J2_127_3477_n2708), 
        .A2(DP_OP_423J2_125_3477_n2233), .Y(DP_OP_423J2_125_3477_n2216) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1844 ( .A1(DP_OP_425J2_127_3477_n2621), 
        .A2(n1441), .Y(DP_OP_425J2_127_3477_n2605) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1847 ( .A1(DP_OP_423J2_125_3477_n2448), 
        .A2(n1441), .Y(DP_OP_422J2_124_3477_n2608) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2023 ( .A1(DP_OP_422J2_124_3477_n2800), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_422J2_124_3477_n2784) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2060 ( .A1(DP_OP_424J2_126_3477_n2317), 
        .A2(n1438), .Y(DP_OP_422J2_124_3477_n2821) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1844 ( .A1(DP_OP_423J2_125_3477_n2621), 
        .A2(n1441), .Y(DP_OP_423J2_125_3477_n2605) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1668 ( .A1(DP_OP_422J2_124_3477_n2621), 
        .A2(n1489), .Y(DP_OP_423J2_125_3477_n2429) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1370 ( .A1(DP_OP_424J2_126_3477_n2799), 
        .A2(n1442), .Y(DP_OP_422J2_124_3477_n2131) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1441 ( .A1(DP_OP_425J2_127_3477_n2710), 
        .A2(DP_OP_425J2_127_3477_n2231), .Y(DP_OP_423J2_125_3477_n2202) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1270 ( .A1(DP_OP_425J2_127_3477_n2971), 
        .A2(DP_OP_424J2_126_3477_n2056), .Y(DP_OP_424J2_126_3477_n2031) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2107 ( .A1(DP_OP_422J2_124_3477_n2884), 
        .A2(DP_OP_423J2_125_3477_n2892), .Y(DP_OP_422J2_124_3477_n2868) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1534 ( .A1(DP_OP_422J2_124_3477_n2311), 
        .A2(DP_OP_422J2_124_3477_n2320), .Y(DP_OP_422J2_124_3477_n2295) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1270 ( .A1(DP_OP_422J2_124_3477_n2047), 
        .A2(DP_OP_422J2_124_3477_n2056), .Y(DP_OP_422J2_124_3477_n2031) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1234 ( .A1(DP_OP_422J2_124_3477_n2003), 
        .A2(DP_OP_422J2_124_3477_n2013), .Y(DP_OP_422J2_124_3477_n1995) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2282 ( .A1(DP_OP_424J2_126_3477_n3057), 
        .A2(DP_OP_423J2_125_3477_n3066), .Y(DP_OP_424J2_126_3477_n3041) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1483 ( .A1(DP_OP_424J2_126_3477_n2268), 
        .A2(n1427), .Y(DP_OP_424J2_126_3477_n2244) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1570 ( .A1(DP_OP_423J2_125_3477_n2795), 
        .A2(n875), .Y(DP_OP_425J2_127_3477_n2331) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2057 ( .A1(DP_OP_422J2_124_3477_n2842), 
        .A2(n1438), .Y(DP_OP_422J2_124_3477_n2818) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1844 ( .A1(DP_OP_425J2_127_3477_n2445), 
        .A2(n1441), .Y(DP_OP_424J2_126_3477_n2605) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U2203 ( .A1(DP_OP_422J2_124_3477_n2972), 
        .A2(n676), .Y(DP_OP_422J2_124_3477_n2964) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2058 ( .A1(DP_OP_424J2_126_3477_n2315), 
        .A2(n1438), .Y(DP_OP_422J2_124_3477_n2819) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1669 ( .A1(DP_OP_422J2_124_3477_n2446), 
        .A2(n1489), .Y(DP_OP_422J2_124_3477_n2430) );
  NOR2X0_HVT DP_OP_422J2_124_3477_U1667 ( .A1(DP_OP_422J2_124_3477_n2444), 
        .A2(n1489), .Y(DP_OP_422J2_124_3477_n2428) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U2283 ( .A1(DP_OP_422J2_124_3477_n3058), 
        .A2(DP_OP_424J2_126_3477_n3066), .Y(DP_OP_422J2_124_3477_n3042) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1663 ( .A1(DP_OP_423J2_125_3477_n2448), 
        .A2(n789), .Y(DP_OP_423J2_125_3477_n2424) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2022 ( .A1(DP_OP_423J2_125_3477_n2799), 
        .A2(DP_OP_423J2_125_3477_n2804), .Y(DP_OP_423J2_125_3477_n2783) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U2059 ( .A1(DP_OP_423J2_125_3477_n2844), 
        .A2(n1438), .Y(DP_OP_423J2_125_3477_n2820) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1927 ( .A1(DP_OP_423J2_125_3477_n2712), 
        .A2(n1440), .Y(DP_OP_423J2_125_3477_n2688) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U2060 ( .A1(DP_OP_424J2_126_3477_n2845), 
        .A2(n1438), .Y(DP_OP_424J2_126_3477_n2821) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1371 ( .A1(DP_OP_423J2_125_3477_n2140), 
        .A2(n1442), .Y(DP_OP_423J2_125_3477_n2132) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1924 ( .A1(DP_OP_423J2_125_3477_n2225), 
        .A2(n1440), .Y(DP_OP_425J2_127_3477_n2685) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1368 ( .A1(DP_OP_422J2_124_3477_n2929), 
        .A2(n1442), .Y(DP_OP_423J2_125_3477_n2129) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1843 ( .A1(DP_OP_425J2_127_3477_n2620), 
        .A2(n1441), .Y(DP_OP_425J2_127_3477_n2604) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1806 ( .A1(DP_OP_424J2_126_3477_n2443), 
        .A2(DP_OP_422J2_124_3477_n2585), .Y(DP_OP_425J2_127_3477_n2567) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1928 ( .A1(DP_OP_423J2_125_3477_n2801), 
        .A2(n1440), .Y(DP_OP_424J2_126_3477_n2689) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1370 ( .A1(DP_OP_425J2_127_3477_n2799), 
        .A2(n1442), .Y(DP_OP_423J2_125_3477_n2131) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1847 ( .A1(DP_OP_423J2_125_3477_n2624), 
        .A2(n1441), .Y(DP_OP_423J2_125_3477_n2608) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1746 ( .A1(DP_OP_422J2_124_3477_n2399), 
        .A2(n772), .Y(DP_OP_424J2_126_3477_n2507) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1570 ( .A1(DP_OP_423J2_125_3477_n2267), 
        .A2(n875), .Y(DP_OP_424J2_126_3477_n2331) );
  NOR2X1_HVT DP_OP_424J2_126_3477_U1482 ( .A1(DP_OP_424J2_126_3477_n2267), 
        .A2(DP_OP_424J2_126_3477_n2275), .Y(DP_OP_424J2_126_3477_n2243) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1350 ( .A1(DP_OP_425J2_127_3477_n2883), 
        .A2(DP_OP_424J2_126_3477_n2143), .Y(DP_OP_424J2_126_3477_n2111) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1878 ( .A1(DP_OP_423J2_125_3477_n2751), 
        .A2(n1400), .Y(DP_OP_424J2_126_3477_n2639) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1928 ( .A1(DP_OP_423J2_125_3477_n2229), 
        .A2(n1440), .Y(DP_OP_425J2_127_3477_n2689) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U2060 ( .A1(DP_OP_423J2_125_3477_n2097), 
        .A2(n1438), .Y(DP_OP_425J2_127_3477_n2821) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1370 ( .A1(DP_OP_422J2_124_3477_n2007), 
        .A2(n1442), .Y(DP_OP_425J2_127_3477_n2131) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1410 ( .A1(DP_OP_424J2_126_3477_n2883), 
        .A2(DP_OP_425J2_127_3477_n2189), .Y(DP_OP_425J2_127_3477_n2171) );
  NOR2X1_HVT DP_OP_425J2_127_3477_U1534 ( .A1(DP_OP_425J2_127_3477_n2311), 
        .A2(DP_OP_423J2_125_3477_n2320), .Y(DP_OP_425J2_127_3477_n2295) );
  NOR2X0_HVT DP_OP_423J2_125_3477_U1535 ( .A1(DP_OP_425J2_127_3477_n2620), 
        .A2(DP_OP_425J2_127_3477_n2320), .Y(DP_OP_423J2_125_3477_n2296) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U1570 ( .A1(DP_OP_422J2_124_3477_n2355), 
        .A2(n876), .Y(DP_OP_422J2_124_3477_n2331) );
  NOR2X1_HVT DP_OP_423J2_125_3477_U1887 ( .A1(DP_OP_424J2_126_3477_n2576), 
        .A2(n279), .Y(DP_OP_423J2_125_3477_n2648) );
  NOR2X0_HVT DP_OP_425J2_127_3477_U1894 ( .A1(DP_OP_422J2_124_3477_n2795), 
        .A2(DP_OP_425J2_127_3477_n2673), .Y(DP_OP_425J2_127_3477_n2655) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U1894 ( .A1(DP_OP_422J2_124_3477_n2267), 
        .A2(DP_OP_425J2_127_3477_n2673), .Y(DP_OP_424J2_126_3477_n2655) );
  NOR2X0_HVT DP_OP_424J2_126_3477_U106 ( .A1(DP_OP_424J2_126_3477_n115), .A2(
        DP_OP_424J2_126_3477_n144), .Y(DP_OP_424J2_126_3477_n111) );
  NOR2X1_HVT DP_OP_422J2_124_3477_U52 ( .A1(DP_OP_422J2_124_3477_n73), .A2(
        DP_OP_422J2_124_3477_n182), .Y(DP_OP_422J2_124_3477_n71) );
  DFFSSRX1_HVT conv2_sum_c_reg_3_ ( .D(1'b0), .SETB(n1495), .RSTB(
        n_conv2_sum_c[3]), .CLK(clk), .Q(conv2_sum_c[3]), .QN(n1988) );
  DFFSSRX2_HVT conv2_sum_a_reg_9_ ( .D(1'b0), .SETB(n1434), .RSTB(
        n_conv2_sum_a[9]), .CLK(clk), .Q(conv2_sum_a[9]), .QN(n1874) );
  AO221X1_HVT U3 ( .A1(1'b1), .A2(n2141), .A3(n980), .A4(n983), .A5(n984), .Y(
        n1932) );
  OA221X1_HVT U4 ( .A1(1'b0), .A2(DP_OP_423J2_125_3477_n149), .A3(
        DP_OP_423J2_125_3477_n148), .A4(DP_OP_423J2_125_3477_n156), .A5(n1196), 
        .Y(DP_OP_423J2_125_3477_n145) );
  OA221X1_HVT U5 ( .A1(1'b0), .A2(DP_OP_423J2_125_3477_n78), .A3(
        DP_OP_423J2_125_3477_n77), .A4(DP_OP_423J2_125_3477_n85), .A5(n1157), 
        .Y(n1159) );
  OA221X1_HVT U6 ( .A1(1'b0), .A2(DP_OP_425J2_127_3477_n78), .A3(
        DP_OP_425J2_127_3477_n77), .A4(DP_OP_425J2_127_3477_n85), .A5(n1123), 
        .Y(n1124) );
  OA221X1_HVT U7 ( .A1(1'b0), .A2(DP_OP_422J2_124_3477_n65), .A3(
        DP_OP_422J2_124_3477_n60), .A4(DP_OP_422J2_124_3477_n198), .A5(n1120), 
        .Y(DP_OP_422J2_124_3477_n57) );
  OAI22X1_HVT U8 ( .A1(n2039), .A2(1'b0), .A3(conv2_sum_a[16]), .A4(n1883), 
        .Y(n1039) );
  OA221X1_HVT U9 ( .A1(1'b0), .A2(DP_OP_424J2_126_3477_n78), .A3(
        DP_OP_424J2_126_3477_n77), .A4(DP_OP_424J2_126_3477_n85), .A5(n1074), 
        .Y(n1075) );
  OA221X1_HVT U10 ( .A1(1'b0), .A2(DP_OP_422J2_124_3477_n78), .A3(
        DP_OP_422J2_124_3477_n77), .A4(DP_OP_422J2_124_3477_n85), .A5(n1071), 
        .Y(n1072) );
  OA221X1_HVT U11 ( .A1(1'b0), .A2(DP_OP_423J2_125_3477_n65), .A3(
        DP_OP_423J2_125_3477_n60), .A4(DP_OP_423J2_125_3477_n198), .A5(n1069), 
        .Y(DP_OP_423J2_125_3477_n57) );
  OA221X1_HVT U12 ( .A1(1'b0), .A2(DP_OP_425J2_127_3477_n65), .A3(
        DP_OP_425J2_127_3477_n60), .A4(DP_OP_425J2_127_3477_n198), .A5(n1044), 
        .Y(DP_OP_425J2_127_3477_n57) );
  OA221X1_HVT U13 ( .A1(1'b0), .A2(DP_OP_422J2_124_3477_n149), .A3(
        DP_OP_422J2_124_3477_n148), .A4(DP_OP_422J2_124_3477_n156), .A5(n1024), 
        .Y(DP_OP_422J2_124_3477_n145) );
  OA221X1_HVT U14 ( .A1(1'b0), .A2(DP_OP_424J2_126_3477_n65), .A3(
        DP_OP_424J2_126_3477_n60), .A4(DP_OP_424J2_126_3477_n198), .A5(n1013), 
        .Y(DP_OP_424J2_126_3477_n57) );
  OA221X1_HVT U15 ( .A1(1'b0), .A2(DP_OP_424J2_126_3477_n149), .A3(
        DP_OP_424J2_126_3477_n148), .A4(DP_OP_424J2_126_3477_n156), .A5(n1011), 
        .Y(DP_OP_424J2_126_3477_n145) );
  OA221X1_HVT U16 ( .A1(1'b0), .A2(DP_OP_425J2_127_3477_n149), .A3(
        DP_OP_425J2_127_3477_n148), .A4(DP_OP_425J2_127_3477_n156), .A5(n977), 
        .Y(DP_OP_425J2_127_3477_n145) );
  OA221X1_HVT U17 ( .A1(1'b0), .A2(n2136), .A3(tmp_big1[8]), .A4(n973), .A5(
        n974), .Y(n1951) );
  NOR2X4_HVT U18 ( .A1(DP_OP_424J2_126_3477_n2932), .A2(
        DP_OP_422J2_124_3477_n2144), .Y(DP_OP_425J2_127_3477_n2124) );
  NOR2X4_HVT U19 ( .A1(DP_OP_425J2_127_3477_n2843), .A2(
        DP_OP_423J2_125_3477_n2099), .Y(DP_OP_423J2_125_3477_n2071) );
  NOR2X4_HVT U20 ( .A1(DP_OP_425J2_127_3477_n2840), .A2(
        DP_OP_423J2_125_3477_n2099), .Y(DP_OP_423J2_125_3477_n2068) );
  NOR2X2_HVT U21 ( .A1(DP_OP_423J2_125_3477_n2097), .A2(
        DP_OP_423J2_125_3477_n2099), .Y(DP_OP_423J2_125_3477_n2073) );
  OR2X2_HVT U22 ( .A1(DP_OP_423J2_125_3477_n2090), .A2(
        DP_OP_423J2_125_3477_n2099), .Y(DP_OP_423J2_125_3477_n2066) );
  NOR2X2_HVT U23 ( .A1(DP_OP_423J2_125_3477_n2096), .A2(
        DP_OP_423J2_125_3477_n2099), .Y(DP_OP_423J2_125_3477_n2072) );
  NOR2X2_HVT U24 ( .A1(DP_OP_423J2_125_3477_n2094), .A2(
        DP_OP_423J2_125_3477_n2099), .Y(DP_OP_423J2_125_3477_n2070) );
  NOR2X2_HVT U25 ( .A1(DP_OP_424J2_126_3477_n2845), .A2(
        DP_OP_423J2_125_3477_n2099), .Y(DP_OP_422J2_124_3477_n2073) );
  NOR2X0_HVT U26 ( .A1(DP_OP_425J2_127_3477_n2841), .A2(
        DP_OP_423J2_125_3477_n2099), .Y(DP_OP_423J2_125_3477_n2069) );
  INVX1_HVT U27 ( .A(conv_weight_box[49]), .Y(n1) );
  NOR2X4_HVT U28 ( .A1(DP_OP_423J2_125_3477_n2931), .A2(
        DP_OP_423J2_125_3477_n2099), .Y(DP_OP_422J2_124_3477_n2071) );
  NOR2X4_HVT U29 ( .A1(DP_OP_423J2_125_3477_n2932), .A2(
        DP_OP_423J2_125_3477_n2099), .Y(DP_OP_422J2_124_3477_n2072) );
  MUX21X2_HVT U30 ( .A1(conv1_sram_rdata_weight[40]), .A2(
        conv2_sram_rdata_weight[40]), .S0(n1515), .Y(conv_weight_box[26]) );
  NOR2X4_HVT U31 ( .A1(DP_OP_422J2_124_3477_n2091), .A2(n1428), .Y(
        DP_OP_424J2_126_3477_n2831) );
  MUX21X2_HVT U32 ( .A1(conv2_sram_rdata_weight[80]), .A2(
        conv1_sram_rdata_weight[80]), .S0(n345), .Y(conv_weight_box[53]) );
  NOR2X4_HVT U33 ( .A1(DP_OP_425J2_127_3477_n2404), .A2(
        DP_OP_424J2_126_3477_n2673), .Y(DP_OP_424J2_126_3477_n2660) );
  NOR2X4_HVT U34 ( .A1(DP_OP_425J2_127_3477_n2401), .A2(
        DP_OP_424J2_126_3477_n2673), .Y(DP_OP_424J2_126_3477_n2657) );
  NOR2X4_HVT U35 ( .A1(DP_OP_423J2_125_3477_n2668), .A2(
        DP_OP_422J2_124_3477_n2673), .Y(DP_OP_423J2_125_3477_n2660) );
  NOR2X4_HVT U36 ( .A1(DP_OP_424J2_126_3477_n2669), .A2(n1), .Y(
        DP_OP_424J2_126_3477_n2661) );
  NOR2X4_HVT U37 ( .A1(DP_OP_423J2_125_3477_n2754), .A2(
        DP_OP_425J2_127_3477_n2673), .Y(DP_OP_424J2_126_3477_n2658) );
  NOR2X4_HVT U38 ( .A1(DP_OP_422J2_124_3477_n2268), .A2(
        DP_OP_422J2_124_3477_n2673), .Y(DP_OP_424J2_126_3477_n2656) );
  OR2X4_HVT U39 ( .A1(DP_OP_425J2_127_3477_n2049), .A2(n1506), .Y(
        DP_OP_424J2_126_3477_n2985) );
  OR2X2_HVT U40 ( .A1(DP_OP_425J2_127_3477_n2053), .A2(n1506), .Y(
        DP_OP_424J2_126_3477_n2989) );
  OR2X2_HVT U41 ( .A1(DP_OP_422J2_124_3477_n3017), .A2(n1506), .Y(
        DP_OP_422J2_124_3477_n2985) );
  OR2X2_HVT U42 ( .A1(DP_OP_424J2_126_3477_n2138), .A2(n1506), .Y(
        DP_OP_422J2_124_3477_n2986) );
  OR2X2_HVT U43 ( .A1(DP_OP_424J2_126_3477_n3015), .A2(n1506), .Y(
        DP_OP_424J2_126_3477_n2983) );
  OR2X2_HVT U44 ( .A1(DP_OP_424J2_126_3477_n2003), .A2(n1506), .Y(
        DP_OP_425J2_127_3477_n2983) );
  OR2X2_HVT U45 ( .A1(DP_OP_424J2_126_3477_n2929), .A2(n1506), .Y(
        DP_OP_423J2_125_3477_n2985) );
  OR2X2_HVT U46 ( .A1(DP_OP_422J2_124_3477_n2003), .A2(n1506), .Y(
        DP_OP_423J2_125_3477_n2983) );
  OR2X2_HVT U47 ( .A1(DP_OP_424J2_126_3477_n2006), .A2(n1506), .Y(
        DP_OP_425J2_127_3477_n2986) );
  OR2X2_HVT U48 ( .A1(DP_OP_425J2_127_3477_n3021), .A2(n1506), .Y(
        DP_OP_425J2_127_3477_n2989) );
  OA21X2_HVT U49 ( .A1(DP_OP_422J2_124_3477_n241), .A2(n1255), .A3(
        DP_OP_422J2_124_3477_n240), .Y(n1256) );
  NOR2X0_HVT U50 ( .A1(DP_OP_424J2_126_3477_n2667), .A2(
        DP_OP_425J2_127_3477_n2673), .Y(DP_OP_424J2_126_3477_n2659) );
  OR2X4_HVT U51 ( .A1(DP_OP_423J2_125_3477_n2750), .A2(
        DP_OP_422J2_124_3477_n2673), .Y(DP_OP_424J2_126_3477_n2654) );
  OR2X2_HVT U52 ( .A1(DP_OP_422J2_124_3477_n2975), .A2(
        DP_OP_424J2_126_3477_n2186), .Y(DP_OP_424J2_126_3477_n2151) );
  OR2X4_HVT U53 ( .A1(DP_OP_424J2_126_3477_n2268), .A2(
        DP_OP_425J2_127_3477_n2186), .Y(DP_OP_423J2_125_3477_n2148) );
  NOR2X0_HVT U54 ( .A1(DP_OP_422J2_124_3477_n2974), .A2(n1344), .Y(
        DP_OP_424J2_126_3477_n2166) );
  INVX2_HVT U55 ( .A(conv_weight_box[8]), .Y(DP_OP_425J2_127_3477_n2057) );
  NBUFFX8_HVT U56 ( .A(n1332), .Y(n1366) );
  INVX1_HVT U57 ( .A(DP_OP_424J2_126_3477_n666), .Y(n2) );
  INVX2_HVT U58 ( .A(n2), .Y(n3) );
  INVX2_HVT U59 ( .A(n182), .Y(n1001) );
  INVX2_HVT U60 ( .A(conv_weight_box[12]), .Y(DP_OP_424J2_126_3477_n2979) );
  INVX2_HVT U61 ( .A(conv_weight_box[46]), .Y(DP_OP_425J2_127_3477_n2714) );
  OR2X1_HVT U62 ( .A1(DP_OP_425J2_127_3477_n2445), .A2(
        DP_OP_425J2_127_3477_n2714), .Y(DP_OP_423J2_125_3477_n2677) );
  OR2X1_HVT U63 ( .A1(DP_OP_424J2_126_3477_n2623), .A2(
        DP_OP_425J2_127_3477_n2714), .Y(DP_OP_423J2_125_3477_n2679) );
  NOR2X0_HVT U64 ( .A1(DP_OP_423J2_125_3477_n2706), .A2(
        DP_OP_425J2_127_3477_n2714), .Y(DP_OP_423J2_125_3477_n2674) );
  OR2X4_HVT U65 ( .A1(DP_OP_425J2_127_3477_n2710), .A2(
        DP_OP_425J2_127_3477_n2714), .Y(DP_OP_425J2_127_3477_n2678) );
  OR2X4_HVT U66 ( .A1(mode[0]), .A2(n951), .Y(n4) );
  FADDX1_HVT U67 ( .A(DP_OP_422J2_124_3477_n1243), .B(
        DP_OP_422J2_124_3477_n1239), .CI(DP_OP_422J2_124_3477_n1237), .S(n5)
         );
  AND2X1_HVT U68 ( .A1(DP_OP_422J2_124_3477_n419), .A2(
        DP_OP_422J2_124_3477_n512), .Y(n6) );
  INVX1_HVT U69 ( .A(n286), .Y(n285) );
  NBUFFX8_HVT U70 ( .A(DP_OP_423J2_125_3477_n2101), .Y(n621) );
  INVX1_HVT U71 ( .A(DP_OP_423J2_125_3477_n2101), .Y(n620) );
  INVX1_HVT U72 ( .A(DP_OP_423J2_125_3477_n2101), .Y(n622) );
  NAND2X0_HVT U73 ( .A1(DP_OP_423J2_125_3477_n220), .A2(n1394), .Y(n1392) );
  NAND2X0_HVT U74 ( .A1(n7010), .A2(DP_OP_423J2_125_3477_n226), .Y(
        DP_OP_423J2_125_3477_n220) );
  NAND2X0_HVT U75 ( .A1(n1610), .A2(n1609), .Y(n7010) );
  OR2X1_HVT U76 ( .A1(DP_OP_423J2_125_3477_n418), .A2(
        DP_OP_423J2_125_3477_n373), .Y(n1609) );
  AND2X1_HVT U77 ( .A1(DP_OP_423J2_125_3477_n419), .A2(
        DP_OP_423J2_125_3477_n512), .Y(n1610) );
  NBUFFX2_HVT U78 ( .A(conv_weight_box[46]), .Y(n8) );
  NAND2X0_HVT U79 ( .A1(conv_weight_box[46]), .A2(n9010), .Y(
        DP_OP_424J2_126_3477_n2679) );
  INVX2_HVT U80 ( .A(DP_OP_425J2_127_3477_n2359), .Y(n9010) );
  NAND2X0_HVT U81 ( .A1(conv_weight_box[46]), .A2(n10), .Y(
        DP_OP_424J2_126_3477_n2681) );
  INVX2_HVT U82 ( .A(DP_OP_423J2_125_3477_n2801), .Y(n10) );
  NAND2X0_HVT U83 ( .A1(n8), .A2(n11), .Y(DP_OP_423J2_125_3477_n2678) );
  INVX2_HVT U84 ( .A(DP_OP_422J2_124_3477_n2314), .Y(n11) );
  NAND2X0_HVT U85 ( .A1(n8), .A2(n12), .Y(DP_OP_424J2_126_3477_n2676) );
  INVX2_HVT U86 ( .A(DP_OP_422J2_124_3477_n2224), .Y(n12) );
  NAND2X0_HVT U87 ( .A1(n8), .A2(n13), .Y(DP_OP_424J2_126_3477_n2677) );
  INVX2_HVT U88 ( .A(DP_OP_422J2_124_3477_n2225), .Y(n13) );
  NAND2X0_HVT U89 ( .A1(n8), .A2(n14), .Y(DP_OP_424J2_126_3477_n2680) );
  INVX2_HVT U90 ( .A(DP_OP_424J2_126_3477_n2712), .Y(n14) );
  NAND2X0_HVT U91 ( .A1(n8), .A2(n15), .Y(DP_OP_423J2_125_3477_n2680) );
  INVX2_HVT U92 ( .A(DP_OP_423J2_125_3477_n2712), .Y(n15) );
  NAND2X0_HVT U93 ( .A1(n8), .A2(n16), .Y(DP_OP_423J2_125_3477_n2675) );
  INVX2_HVT U94 ( .A(DP_OP_424J2_126_3477_n2619), .Y(n16) );
  NAND2X0_HVT U95 ( .A1(n8), .A2(n17), .Y(DP_OP_424J2_126_3477_n2678) );
  INVX2_HVT U96 ( .A(DP_OP_423J2_125_3477_n2798), .Y(n17) );
  NAND2X0_HVT U97 ( .A1(n8), .A2(n18), .Y(DP_OP_423J2_125_3477_n2676) );
  INVX2_HVT U98 ( .A(DP_OP_423J2_125_3477_n2708), .Y(n18) );
  NAND2X0_HVT U99 ( .A1(n8), .A2(n19), .Y(DP_OP_424J2_126_3477_n2675) );
  INVX2_HVT U100 ( .A(DP_OP_422J2_124_3477_n2223), .Y(n19) );
  AND2X4_HVT U101 ( .A1(n8), .A2(n20), .Y(DP_OP_424J2_126_3477_n2674) );
  INVX2_HVT U102 ( .A(DP_OP_423J2_125_3477_n2794), .Y(n20) );
  NAND2X0_HVT U103 ( .A1(n778), .A2(n21), .Y(DP_OP_422J2_124_3477_n2017) );
  INVX2_HVT U104 ( .A(DP_OP_422J2_124_3477_n2049), .Y(n21) );
  NAND2X0_HVT U105 ( .A1(n778), .A2(n22), .Y(DP_OP_424J2_126_3477_n2021) );
  INVX2_HVT U106 ( .A(DP_OP_425J2_127_3477_n2977), .Y(n22) );
  NAND2X0_HVT U107 ( .A1(n778), .A2(n23), .Y(DP_OP_422J2_124_3477_n2019) );
  INVX2_HVT U108 ( .A(DP_OP_422J2_124_3477_n2051), .Y(n23) );
  NAND2X0_HVT U109 ( .A1(n778), .A2(n24), .Y(DP_OP_422J2_124_3477_n2021) );
  INVX2_HVT U110 ( .A(DP_OP_424J2_126_3477_n2889), .Y(n24) );
  AND2X1_HVT U111 ( .A1(n778), .A2(n25), .Y(DP_OP_422J2_124_3477_n2014) );
  INVX2_HVT U112 ( .A(DP_OP_422J2_124_3477_n2046), .Y(n25) );
  AO22X1_HVT U113 ( .A1(n619), .A2(conv1_sram_rdata_weight[52]), .A3(n26), 
        .A4(conv2_sram_rdata_weight[52]), .Y(conv_weight_box[36]) );
  INVX4_HVT U114 ( .A(n619), .Y(n26) );
  NAND3X0_HVT U115 ( .A1(n1465), .A2(n1466), .A3(n1467), .Y(
        DP_OP_423J2_125_3477_n512) );
  NBUFFX8_HVT U116 ( .A(n1518), .Y(n27) );
  INVX4_HVT U117 ( .A(n29), .Y(n1518) );
  AO21X2_HVT U118 ( .A1(n182), .A2(n1766), .A3(n28), .Y(n_conv2_sum_c[24]) );
  AO22X1_HVT U119 ( .A1(n29), .A2(n1151), .A3(n1750), .A4(n1751), .Y(n28) );
  OA21X1_HVT U120 ( .A1(n806), .A2(n805), .A3(n802), .Y(n29) );
  NBUFFX8_HVT U121 ( .A(n779), .Y(n30) );
  IBUFFX8_HVT U122 ( .A(n31), .Y(DP_OP_425J2_127_3477_n2014) );
  OR2X2_HVT U123 ( .A1(DP_OP_425J2_127_3477_n2046), .A2(n779), .Y(n31) );
  OA21X2_HVT U124 ( .A1(n711), .A2(n781), .A3(n780), .Y(n779) );
  NBUFFX2_HVT U125 ( .A(n694), .Y(n32) );
  NBUFFX2_HVT U126 ( .A(n34), .Y(n33) );
  NBUFFX16_HVT U127 ( .A(n694), .Y(n34) );
  NOR2X0_HVT U128 ( .A1(DP_OP_422J2_124_3477_n3059), .A2(n32), .Y(
        DP_OP_422J2_124_3477_n3051) );
  OA21X2_HVT U129 ( .A1(n843), .A2(n697), .A3(n696), .Y(n694) );
  NBUFFX8_HVT U130 ( .A(n601), .Y(n35) );
  INVX2_HVT U131 ( .A(n1485), .Y(n329) );
  MUX21X2_HVT U132 ( .A1(n606), .A2(n178), .S0(n1485), .Y(n601) );
  NBUFFX2_HVT U133 ( .A(n585), .Y(n36) );
  AO22X1_HVT U134 ( .A1(n769), .A2(n784), .A3(n785), .A4(n38), .Y(n585) );
  NBUFFX2_HVT U135 ( .A(n585), .Y(n37) );
  INVX2_HVT U136 ( .A(n769), .Y(n38) );
  INVX2_HVT U137 ( .A(conv_weight_box[23]), .Y(DP_OP_422J2_124_3477_n2890) );
  AO22X1_HVT U138 ( .A1(n92), .A2(conv1_sram_rdata_weight[35]), .A3(
        conv2_sram_rdata_weight[35]), .A4(n41), .Y(conv_weight_box[23]) );
  XOR3X1_HVT U139 ( .A1(DP_OP_424J2_126_3477_n2019), .A2(n39), .A3(n42), .Y(
        DP_OP_424J2_126_3477_n1393) );
  NAND2X2_HVT U140 ( .A1(n585), .A2(n586), .Y(n42) );
  NAND2X2_HVT U141 ( .A1(conv_weight_box[23]), .A2(n40), .Y(n39) );
  FADDX2_HVT U142 ( .A(n42), .B(n39), .CI(DP_OP_424J2_126_3477_n2019), .CO(
        DP_OP_424J2_126_3477_n1392) );
  INVX4_HVT U143 ( .A(DP_OP_424J2_126_3477_n2887), .Y(n40) );
  INVX1_HVT U144 ( .A(n92), .Y(n41) );
  NBUFFX2_HVT U145 ( .A(n1425), .Y(n43) );
  AND2X1_HVT U146 ( .A1(n1425), .A2(n44), .Y(DP_OP_422J2_124_3477_n1927) );
  INVX2_HVT U147 ( .A(n1874), .Y(n44) );
  AND2X1_HVT U148 ( .A1(n1425), .A2(n45), .Y(DP_OP_424J2_126_3477_n1929) );
  INVX2_HVT U149 ( .A(n1855), .Y(n45) );
  AND2X1_HVT U150 ( .A1(n43), .A2(n46), .Y(DP_OP_424J2_126_3477_n1933) );
  INVX2_HVT U151 ( .A(n1988), .Y(n46) );
  AND2X1_HVT U152 ( .A1(n43), .A2(n47), .Y(DP_OP_425J2_127_3477_n510) );
  INVX2_HVT U153 ( .A(n1288), .Y(n47) );
  AND2X1_HVT U154 ( .A1(n43), .A2(n48), .Y(DP_OP_424J2_126_3477_n1927) );
  INVX2_HVT U155 ( .A(n1993), .Y(n48) );
  AND2X1_HVT U156 ( .A1(n43), .A2(n49), .Y(DP_OP_425J2_127_3477_n1936) );
  INVX2_HVT U157 ( .A(n1294), .Y(n49) );
  AND2X1_HVT U158 ( .A1(n43), .A2(n50), .Y(DP_OP_423J2_125_3477_n328) );
  INVX2_HVT U159 ( .A(n1322), .Y(n50) );
  AND2X1_HVT U160 ( .A1(n43), .A2(n51), .Y(DP_OP_423J2_125_3477_n326) );
  INVX2_HVT U161 ( .A(n1316), .Y(n51) );
  AND2X1_HVT U162 ( .A1(n43), .A2(n52), .Y(DP_OP_423J2_125_3477_n320) );
  INVX2_HVT U163 ( .A(n1315), .Y(n52) );
  AND2X1_HVT U164 ( .A1(n43), .A2(n53), .Y(DP_OP_425J2_127_3477_n312) );
  INVX2_HVT U165 ( .A(n1314), .Y(n53) );
  AND2X1_HVT U166 ( .A1(n43), .A2(n54), .Y(DP_OP_425J2_127_3477_n310) );
  INVX2_HVT U167 ( .A(n1304), .Y(n54) );
  AND2X4_HVT U168 ( .A1(n43), .A2(n55), .Y(DP_OP_425J2_127_3477_n306) );
  INVX2_HVT U169 ( .A(n1327), .Y(n55) );
  NBUFFX2_HVT U170 ( .A(conv_weight_box[57]), .Y(n56) );
  NAND2X0_HVT U171 ( .A1(conv_weight_box[57]), .A2(n57), .Y(
        DP_OP_422J2_124_3477_n2434) );
  INVX2_HVT U172 ( .A(DP_OP_422J2_124_3477_n2442), .Y(n57) );
  AND2X1_HVT U173 ( .A1(conv_weight_box[57]), .A2(n58), .Y(
        DP_OP_422J2_124_3477_n2439) );
  INVX2_HVT U174 ( .A(DP_OP_423J2_125_3477_n2579), .Y(n58) );
  AND2X1_HVT U175 ( .A1(n56), .A2(n59), .Y(DP_OP_422J2_124_3477_n2436) );
  INVX2_HVT U176 ( .A(DP_OP_422J2_124_3477_n2444), .Y(n59) );
  AND2X1_HVT U177 ( .A1(n56), .A2(n60), .Y(DP_OP_422J2_124_3477_n2435) );
  INVX2_HVT U178 ( .A(DP_OP_422J2_124_3477_n2443), .Y(n60) );
  AND2X1_HVT U179 ( .A1(n56), .A2(n61), .Y(DP_OP_422J2_124_3477_n2438) );
  INVX2_HVT U180 ( .A(DP_OP_422J2_124_3477_n2446), .Y(n61) );
  AND2X1_HVT U181 ( .A1(n56), .A2(n62), .Y(DP_OP_422J2_124_3477_n2441) );
  INVX2_HVT U182 ( .A(DP_OP_423J2_125_3477_n2581), .Y(n62) );
  AND2X1_HVT U183 ( .A1(n56), .A2(n63), .Y(DP_OP_422J2_124_3477_n2440) );
  INVX2_HVT U184 ( .A(DP_OP_422J2_124_3477_n2448), .Y(n63) );
  AND2X1_HVT U185 ( .A1(n56), .A2(n64), .Y(DP_OP_422J2_124_3477_n2437) );
  INVX2_HVT U186 ( .A(DP_OP_422J2_124_3477_n2445), .Y(n64) );
  AND2X4_HVT U187 ( .A1(n56), .A2(n65), .Y(DP_OP_423J2_125_3477_n2440) );
  INVX2_HVT U188 ( .A(DP_OP_423J2_125_3477_n2448), .Y(n65) );
  NBUFFX8_HVT U189 ( .A(DP_OP_425J2_127_3477_n2761), .Y(n66) );
  OR2X1_HVT U190 ( .A1(n67), .A2(DP_OP_425J2_127_3477_n2761), .Y(n1646) );
  INVX2_HVT U191 ( .A(src_window[178]), .Y(n67) );
  AND2X1_HVT U192 ( .A1(n68), .A2(n669), .Y(DP_OP_424J2_126_3477_n2744) );
  INVX2_HVT U193 ( .A(DP_OP_425J2_127_3477_n2761), .Y(n68) );
  OA21X1_HVT U194 ( .A1(n858), .A2(n7000), .A3(n69), .Y(
        DP_OP_425J2_127_3477_n2761) );
  NAND2X0_HVT U195 ( .A1(n858), .A2(conv2_sram_rdata_weight[56]), .Y(n69) );
  INVX2_HVT U196 ( .A(conv1_sram_rdata_weight[56]), .Y(n7000) );
  INVX2_HVT U197 ( .A(n72), .Y(DP_OP_423J2_125_3477_n241) );
  AO21X1_HVT U198 ( .A1(n1666), .A2(n1665), .A3(n139), .Y(n72) );
  NBUFFX2_HVT U199 ( .A(DP_OP_423J2_125_3477_n241), .Y(n71) );
  AO21X1_HVT U200 ( .A1(n72), .A2(n892), .A3(n1391), .Y(n1390) );
  XOR3X2_HVT U201 ( .A1(DP_OP_424J2_126_3477_n1317), .A2(
        DP_OP_424J2_126_3477_n1474), .A3(DP_OP_424J2_126_3477_n1313), .Y(
        DP_OP_424J2_126_3477_n1269) );
  NBUFFX2_HVT U202 ( .A(n74), .Y(n73) );
  NBUFFX2_HVT U203 ( .A(conv_weight_box[57]), .Y(n74) );
  AND2X1_HVT U204 ( .A1(conv_weight_box[57]), .A2(n75), .Y(
        DP_OP_424J2_126_3477_n2439) );
  INVX2_HVT U205 ( .A(DP_OP_424J2_126_3477_n2447), .Y(n75) );
  NAND2X0_HVT U206 ( .A1(n74), .A2(n76), .Y(DP_OP_424J2_126_3477_n2434) );
  INVX2_HVT U207 ( .A(DP_OP_425J2_127_3477_n2574), .Y(n76) );
  AND2X1_HVT U208 ( .A1(conv_weight_box[57]), .A2(n77), .Y(
        DP_OP_424J2_126_3477_n2437) );
  INVX2_HVT U209 ( .A(DP_OP_422J2_124_3477_n2709), .Y(n77) );
  AND2X1_HVT U210 ( .A1(n74), .A2(n78), .Y(DP_OP_424J2_126_3477_n2436) );
  INVX2_HVT U211 ( .A(DP_OP_425J2_127_3477_n2576), .Y(n78) );
  AND2X1_HVT U212 ( .A1(n74), .A2(n79), .Y(DP_OP_423J2_125_3477_n2435) );
  INVX2_HVT U213 ( .A(DP_OP_422J2_124_3477_n2619), .Y(n79) );
  AND2X1_HVT U214 ( .A1(n74), .A2(n80), .Y(DP_OP_423J2_125_3477_n2436) );
  INVX2_HVT U215 ( .A(DP_OP_422J2_124_3477_n2620), .Y(n80) );
  AND2X1_HVT U216 ( .A1(n73), .A2(n81), .Y(DP_OP_424J2_126_3477_n2435) );
  INVX2_HVT U217 ( .A(DP_OP_424J2_126_3477_n2443), .Y(n81) );
  AND2X1_HVT U218 ( .A1(n74), .A2(n82), .Y(DP_OP_424J2_126_3477_n2440) );
  INVX2_HVT U219 ( .A(DP_OP_425J2_127_3477_n2580), .Y(n82) );
  AND2X1_HVT U220 ( .A1(n73), .A2(n83), .Y(DP_OP_424J2_126_3477_n2438) );
  INVX2_HVT U221 ( .A(DP_OP_425J2_127_3477_n2578), .Y(n83) );
  AND2X1_HVT U222 ( .A1(n73), .A2(n84), .Y(DP_OP_424J2_126_3477_n2441) );
  INVX2_HVT U223 ( .A(DP_OP_425J2_127_3477_n2581), .Y(n84) );
  AND2X4_HVT U224 ( .A1(n74), .A2(n85), .Y(DP_OP_423J2_125_3477_n2441) );
  INVX2_HVT U225 ( .A(DP_OP_422J2_124_3477_n2625), .Y(n85) );
  NBUFFX8_HVT U226 ( .A(DP_OP_422J2_124_3477_n2670), .Y(n86) );
  NBUFFX2_HVT U227 ( .A(n755), .Y(n87) );
  NBUFFX2_HVT U228 ( .A(n755), .Y(n88) );
  INVX2_HVT U229 ( .A(n755), .Y(DP_OP_422J2_124_3477_n2670) );
  NAND2X0_HVT U230 ( .A1(n87), .A2(n756), .Y(DP_OP_424J2_126_3477_n2635) );
  NAND2X0_HVT U231 ( .A1(n88), .A2(n757), .Y(DP_OP_424J2_126_3477_n2637) );
  AO21X1_HVT U232 ( .A1(n9000), .A2(conv1_sram_rdata_weight[75]), .A3(n89), 
        .Y(n755) );
  AND2X1_HVT U233 ( .A1(n425), .A2(conv2_sram_rdata_weight[75]), .Y(n89) );
  INVX2_HVT U234 ( .A(n425), .Y(n9000) );
  INVX4_HVT U235 ( .A(n91), .Y(n423) );
  NBUFFX8_HVT U236 ( .A(n423), .Y(n92) );
  MUX21X2_HVT U237 ( .A1(conv2_sram_rdata_weight[50]), .A2(
        conv1_sram_rdata_weight[50]), .S0(n92), .Y(conv_weight_box[34]) );
  AND2X1_HVT U238 ( .A1(n1516), .A2(mode[1]), .Y(n91) );
  INVX2_HVT U239 ( .A(n93), .Y(conv_weight_box[48]) );
  AO21X1_HVT U240 ( .A1(n687), .A2(n689), .A3(n686), .Y(n93) );
  NAND2X0_HVT U241 ( .A1(conv_weight_box[48]), .A2(n94), .Y(
        DP_OP_424J2_126_3477_n2327) );
  INVX2_HVT U242 ( .A(DP_OP_423J2_125_3477_n2271), .Y(n94) );
  NAND2X0_HVT U243 ( .A1(conv_weight_box[48]), .A2(n95), .Y(
        DP_OP_424J2_126_3477_n2325) );
  INVX2_HVT U244 ( .A(DP_OP_423J2_125_3477_n2269), .Y(n95) );
  NAND2X0_HVT U245 ( .A1(conv_weight_box[48]), .A2(n96), .Y(
        DP_OP_424J2_126_3477_n2329) );
  INVX2_HVT U246 ( .A(DP_OP_422J2_124_3477_n2801), .Y(n96) );
  NAND2X0_HVT U247 ( .A1(conv_weight_box[48]), .A2(n97), .Y(
        DP_OP_425J2_127_3477_n2325) );
  INVX2_HVT U248 ( .A(DP_OP_425J2_127_3477_n2357), .Y(n97) );
  NAND2X0_HVT U249 ( .A1(conv_weight_box[48]), .A2(n98), .Y(
        DP_OP_425J2_127_3477_n2329) );
  INVX2_HVT U250 ( .A(DP_OP_423J2_125_3477_n2801), .Y(n98) );
  NAND2X0_HVT U251 ( .A1(conv_weight_box[48]), .A2(n99), .Y(
        DP_OP_424J2_126_3477_n2324) );
  INVX2_HVT U252 ( .A(DP_OP_423J2_125_3477_n2268), .Y(n99) );
  NAND2X0_HVT U253 ( .A1(conv_weight_box[48]), .A2(n100), .Y(
        DP_OP_424J2_126_3477_n2326) );
  INVX2_HVT U254 ( .A(DP_OP_424J2_126_3477_n2358), .Y(n100) );
  NAND2X0_HVT U255 ( .A1(conv_weight_box[48]), .A2(n101), .Y(
        DP_OP_425J2_127_3477_n2327) );
  INVX2_HVT U256 ( .A(DP_OP_425J2_127_3477_n2359), .Y(n101) );
  NAND2X0_HVT U257 ( .A1(conv_weight_box[48]), .A2(n102), .Y(
        DP_OP_425J2_127_3477_n2324) );
  INVX2_HVT U258 ( .A(DP_OP_425J2_127_3477_n2356), .Y(n102) );
  NAND2X0_HVT U259 ( .A1(conv_weight_box[48]), .A2(n103), .Y(
        DP_OP_424J2_126_3477_n2328) );
  INVX2_HVT U260 ( .A(DP_OP_422J2_124_3477_n2800), .Y(n103) );
  NAND2X0_HVT U261 ( .A1(conv_weight_box[48]), .A2(n104), .Y(
        DP_OP_424J2_126_3477_n2323) );
  INVX2_HVT U262 ( .A(DP_OP_422J2_124_3477_n2795), .Y(n104) );
  AND2X1_HVT U263 ( .A1(conv_weight_box[48]), .A2(n105), .Y(
        DP_OP_424J2_126_3477_n2322) );
  INVX2_HVT U264 ( .A(DP_OP_424J2_126_3477_n2354), .Y(n105) );
  AND2X4_HVT U265 ( .A1(conv_weight_box[48]), .A2(n106), .Y(
        DP_OP_425J2_127_3477_n2322) );
  INVX2_HVT U266 ( .A(DP_OP_423J2_125_3477_n2794), .Y(n106) );
  INVX4_HVT U267 ( .A(n858), .Y(n857) );
  OA22X2_HVT U268 ( .A1(n107), .A2(n858), .A3(n665), .A4(n857), .Y(n254) );
  INVX2_HVT U269 ( .A(conv1_sram_rdata_weight[19]), .Y(n107) );
  INVX4_HVT U270 ( .A(n109), .Y(n1339) );
  AO22X1_HVT U271 ( .A1(n843), .A2(conv1_sram_rdata_weight[38]), .A3(n1154), 
        .A4(conv2_sram_rdata_weight[38]), .Y(n109) );
  NBUFFX2_HVT U272 ( .A(n109), .Y(n108) );
  AND2X1_HVT U273 ( .A1(n108), .A2(n782), .Y(DP_OP_422J2_124_3477_n2156) );
  AND2X4_HVT U274 ( .A1(n108), .A2(n783), .Y(DP_OP_425J2_127_3477_n2159) );
  OA21X1_HVT U275 ( .A1(n1545), .A2(DP_OP_422J2_124_3477_n233), .A3(n1570), 
        .Y(n110) );
  INVX2_HVT U276 ( .A(n110), .Y(n1517) );
  INVX2_HVT U277 ( .A(n1517), .Y(n1580) );
  XOR2X2_HVT U278 ( .A1(n111), .A2(n945), .Y(n_conv2_sum_a[28]) );
  AO21X1_HVT U279 ( .A1(n1517), .A2(DP_OP_422J2_124_3477_n67), .A3(
        DP_OP_422J2_124_3477_n68), .Y(n111) );
  FADDX1_HVT U280 ( .A(DP_OP_425J2_127_3477_n1119), .B(
        DP_OP_425J2_127_3477_n1111), .CI(DP_OP_425J2_127_3477_n1109), .CO(
        DP_OP_425J2_127_3477_n1072) );
  XOR3X2_HVT U281 ( .A1(DP_OP_425J2_127_3477_n1119), .A2(
        DP_OP_425J2_127_3477_n1111), .A3(DP_OP_425J2_127_3477_n1109), .Y(
        DP_OP_425J2_127_3477_n1073) );
  AO22X1_HVT U282 ( .A1(DP_OP_425J2_127_3477_n653), .A2(n114), .A3(
        DP_OP_425J2_127_3477_n651), .A4(n112), .Y(DP_OP_425J2_127_3477_n648)
         );
  NAND2X0_HVT U283 ( .A1(n116), .A2(n113), .Y(n112) );
  INVX2_HVT U284 ( .A(DP_OP_425J2_127_3477_n653), .Y(n113) );
  INVX2_HVT U285 ( .A(n116), .Y(n114) );
  XOR3X2_HVT U286 ( .A1(n116), .A2(DP_OP_425J2_127_3477_n653), .A3(n115), .Y(
        DP_OP_425J2_127_3477_n649) );
  INVX2_HVT U287 ( .A(DP_OP_425J2_127_3477_n651), .Y(n115) );
  AND3X1_HVT U288 ( .A1(n1451), .A2(n1450), .A3(n1452), .Y(n116) );
  NAND2X0_HVT U289 ( .A1(n119), .A2(n1740), .Y(n626) );
  NAND2X0_HVT U290 ( .A1(n119), .A2(n117), .Y(n1033) );
  AND2X1_HVT U291 ( .A1(n1740), .A2(n118), .Y(n117) );
  INVX2_HVT U292 ( .A(n625), .Y(n118) );
  NAND2X0_HVT U293 ( .A1(n1518), .A2(DP_OP_424J2_126_3477_n176), .Y(n119) );
  NBUFFX8_HVT U294 ( .A(n254), .Y(n120) );
  OR2X1_HVT U295 ( .A1(DP_OP_423J2_125_3477_n2973), .A2(n254), .Y(
        DP_OP_423J2_125_3477_n2941) );
  OR2X1_HVT U296 ( .A1(DP_OP_424J2_126_3477_n2051), .A2(n120), .Y(
        DP_OP_425J2_127_3477_n2943) );
  OR2X1_HVT U297 ( .A1(DP_OP_422J2_124_3477_n2971), .A2(n120), .Y(
        DP_OP_422J2_124_3477_n2939) );
  OR2X1_HVT U298 ( .A1(DP_OP_425J2_127_3477_n2974), .A2(n120), .Y(
        DP_OP_425J2_127_3477_n2942) );
  OR2X1_HVT U299 ( .A1(DP_OP_424J2_126_3477_n2973), .A2(n120), .Y(
        DP_OP_424J2_126_3477_n2941) );
  OR2X1_HVT U300 ( .A1(DP_OP_425J2_127_3477_n2973), .A2(n120), .Y(
        DP_OP_425J2_127_3477_n2941) );
  OR2X1_HVT U301 ( .A1(DP_OP_425J2_127_3477_n2182), .A2(n120), .Y(
        DP_OP_423J2_125_3477_n2942) );
  OR2X1_HVT U302 ( .A1(DP_OP_422J2_124_3477_n2975), .A2(n120), .Y(
        DP_OP_422J2_124_3477_n2943) );
  OR2X1_HVT U303 ( .A1(DP_OP_424J2_126_3477_n2883), .A2(n120), .Y(
        DP_OP_423J2_125_3477_n2939) );
  OR2X1_HVT U304 ( .A1(DP_OP_422J2_124_3477_n2051), .A2(n120), .Y(
        DP_OP_423J2_125_3477_n2943) );
  OR2X1_HVT U305 ( .A1(DP_OP_425J2_127_3477_n2971), .A2(n120), .Y(
        DP_OP_425J2_127_3477_n2939) );
  OR2X1_HVT U306 ( .A1(DP_OP_424J2_126_3477_n2972), .A2(n120), .Y(
        DP_OP_424J2_126_3477_n2940) );
  OR2X1_HVT U307 ( .A1(DP_OP_422J2_124_3477_n2972), .A2(n120), .Y(
        DP_OP_422J2_124_3477_n2940) );
  OR2X1_HVT U308 ( .A1(DP_OP_425J2_127_3477_n2972), .A2(n120), .Y(
        DP_OP_425J2_127_3477_n2940) );
  OR2X1_HVT U309 ( .A1(DP_OP_425J2_127_3477_n2976), .A2(n120), .Y(
        DP_OP_425J2_127_3477_n2944) );
  OR2X4_HVT U310 ( .A1(DP_OP_424J2_126_3477_n2971), .A2(n120), .Y(
        DP_OP_424J2_126_3477_n2939) );
  OR2X1_HVT U311 ( .A1(DP_OP_422J2_124_3477_n2048), .A2(n120), .Y(
        DP_OP_423J2_125_3477_n2940) );
  AND2X1_HVT U312 ( .A1(n257), .A2(n121), .Y(DP_OP_425J2_127_3477_n2938) );
  INVX2_HVT U313 ( .A(DP_OP_425J2_127_3477_n2970), .Y(n121) );
  INVX2_HVT U314 ( .A(n120), .Y(n257) );
  INVX2_HVT U315 ( .A(n124), .Y(DP_OP_424J2_126_3477_n245) );
  AO21X1_HVT U316 ( .A1(DP_OP_424J2_126_3477_n295), .A2(
        DP_OP_424J2_126_3477_n250), .A3(n122), .Y(n124) );
  INVX2_HVT U317 ( .A(DP_OP_424J2_126_3477_n249), .Y(n122) );
  IBUFFX8_HVT U318 ( .A(n1042), .Y(n1519) );
  AO21X1_HVT U319 ( .A1(n124), .A2(n1734), .A3(n123), .Y(n1042) );
  INVX2_HVT U320 ( .A(DP_OP_424J2_126_3477_n244), .Y(n123) );
  NAND2X0_HVT U321 ( .A1(DP_OP_424J2_126_3477_n823), .A2(
        DP_OP_424J2_126_3477_n1018), .Y(DP_OP_424J2_126_3477_n244) );
  OR2X1_HVT U322 ( .A1(DP_OP_424J2_126_3477_n1018), .A2(
        DP_OP_424J2_126_3477_n823), .Y(n1734) );
  NAND2X0_HVT U323 ( .A1(DP_OP_424J2_126_3477_n1019), .A2(
        DP_OP_424J2_126_3477_n1021), .Y(DP_OP_424J2_126_3477_n249) );
  NBUFFX2_HVT U324 ( .A(conv_weight_box[43]), .Y(n125) );
  NAND2X0_HVT U325 ( .A1(conv_weight_box[43]), .A2(n415), .Y(
        DP_OP_423J2_125_3477_n2286) );
  AND2X1_HVT U326 ( .A1(conv_weight_box[43]), .A2(n412), .Y(
        DP_OP_424J2_126_3477_n2289) );
  AND2X1_HVT U327 ( .A1(conv_weight_box[43]), .A2(n413), .Y(
        DP_OP_424J2_126_3477_n2288) );
  AND2X1_HVT U328 ( .A1(conv_weight_box[43]), .A2(n416), .Y(
        DP_OP_424J2_126_3477_n2287) );
  AND2X1_HVT U329 ( .A1(n125), .A2(n417), .Y(DP_OP_423J2_125_3477_n2290) );
  AND2X1_HVT U330 ( .A1(n125), .A2(n418), .Y(DP_OP_423J2_125_3477_n2288) );
  AND2X1_HVT U331 ( .A1(conv_weight_box[43]), .A2(n419), .Y(
        DP_OP_423J2_125_3477_n2287) );
  AND2X1_HVT U332 ( .A1(n125), .A2(n420), .Y(DP_OP_424J2_126_3477_n2292) );
  AND2X1_HVT U333 ( .A1(n125), .A2(n421), .Y(DP_OP_423J2_125_3477_n2291) );
  AND2X4_HVT U334 ( .A1(n125), .A2(n422), .Y(DP_OP_423J2_125_3477_n2292) );
  AND2X1_HVT U335 ( .A1(n1484), .A2(n126), .Y(DP_OP_424J2_126_3477_n1928) );
  INVX2_HVT U336 ( .A(n1286), .Y(n126) );
  AND2X1_HVT U337 ( .A1(n1484), .A2(n127), .Y(DP_OP_423J2_125_3477_n1933) );
  INVX2_HVT U338 ( .A(n1981), .Y(n127) );
  AND2X1_HVT U339 ( .A1(n1484), .A2(n129), .Y(DP_OP_425J2_127_3477_n1928) );
  INVX2_HVT U340 ( .A(n1856), .Y(n129) );
  AND2X1_HVT U341 ( .A1(n1484), .A2(n130), .Y(DP_OP_424J2_126_3477_n1936) );
  INVX2_HVT U342 ( .A(n1292), .Y(n130) );
  AND2X1_HVT U343 ( .A1(n1484), .A2(n131), .Y(DP_OP_424J2_126_3477_n1930) );
  INVX2_HVT U344 ( .A(n1862), .Y(n131) );
  AND2X1_HVT U345 ( .A1(n1484), .A2(n132), .Y(DP_OP_424J2_126_3477_n1924) );
  INVX2_HVT U346 ( .A(n1904), .Y(n132) );
  AND2X1_HVT U347 ( .A1(n1484), .A2(n133), .Y(DP_OP_425J2_127_3477_n328) );
  INVX2_HVT U348 ( .A(n1321), .Y(n133) );
  AND2X1_HVT U349 ( .A1(n1484), .A2(n134), .Y(DP_OP_423J2_125_3477_n330) );
  INVX2_HVT U350 ( .A(n1883), .Y(n134) );
  AND2X1_HVT U351 ( .A1(n1484), .A2(n135), .Y(DP_OP_425J2_127_3477_n320) );
  INVX2_HVT U352 ( .A(n1313), .Y(n135) );
  AND2X1_HVT U353 ( .A1(n1484), .A2(n136), .Y(DP_OP_423J2_125_3477_n316) );
  INVX2_HVT U354 ( .A(n1298), .Y(n136) );
  AND2X1_HVT U355 ( .A1(n1484), .A2(n137), .Y(DP_OP_424J2_126_3477_n306) );
  INVX2_HVT U356 ( .A(n1897), .Y(n137) );
  AND2X1_HVT U357 ( .A1(n1484), .A2(n138), .Y(DP_OP_422J2_124_3477_n304) );
  INVX2_HVT U358 ( .A(n1916), .Y(n138) );
  INVX2_HVT U359 ( .A(DP_OP_423J2_125_3477_n244), .Y(n139) );
  INVX2_HVT U360 ( .A(conv_weight_box[63]), .Y(n1491) );
  AND2X1_HVT U361 ( .A1(conv_weight_box[63]), .A2(n140), .Y(
        DP_OP_422J2_124_3477_n2473) );
  INVX2_HVT U362 ( .A(DP_OP_422J2_124_3477_n2489), .Y(n140) );
  OA22X1_HVT U363 ( .A1(n141), .A2(n4), .A3(n237), .A4(n1515), .Y(
        conv_weight_box[63]) );
  INVX2_HVT U364 ( .A(n768), .Y(n1515) );
  INVX2_HVT U365 ( .A(n855), .Y(n141) );
  NBUFFX2_HVT U366 ( .A(conv_weight_box[12]), .Y(n142) );
  NAND2X0_HVT U367 ( .A1(conv_weight_box[12]), .A2(n143), .Y(n1779) );
  INVX2_HVT U368 ( .A(DP_OP_425J2_127_3477_n2976), .Y(n143) );
  AND2X1_HVT U369 ( .A1(conv_weight_box[12]), .A2(n144), .Y(
        DP_OP_423J2_125_3477_n2953) );
  INVX2_HVT U370 ( .A(DP_OP_424J2_126_3477_n2889), .Y(n144) );
  AND2X1_HVT U371 ( .A1(n142), .A2(n145), .Y(DP_OP_425J2_127_3477_n2953) );
  INVX2_HVT U372 ( .A(DP_OP_425J2_127_3477_n2977), .Y(n145) );
  AND2X1_HVT U373 ( .A1(n142), .A2(n146), .Y(DP_OP_425J2_127_3477_n2947) );
  INVX2_HVT U374 ( .A(DP_OP_425J2_127_3477_n2971), .Y(n146) );
  AND2X1_HVT U375 ( .A1(n142), .A2(n147), .Y(DP_OP_425J2_127_3477_n2950) );
  INVX2_HVT U376 ( .A(DP_OP_425J2_127_3477_n2974), .Y(n147) );
  AND2X1_HVT U377 ( .A1(n142), .A2(n148), .Y(DP_OP_425J2_127_3477_n2949) );
  INVX2_HVT U378 ( .A(DP_OP_425J2_127_3477_n2973), .Y(n148) );
  AND2X1_HVT U379 ( .A1(n142), .A2(n149), .Y(DP_OP_423J2_125_3477_n2952) );
  INVX2_HVT U380 ( .A(DP_OP_423J2_125_3477_n2976), .Y(n149) );
  NAND2X0_HVT U381 ( .A1(n142), .A2(n150), .Y(DP_OP_425J2_127_3477_n2946) );
  INVX2_HVT U382 ( .A(DP_OP_425J2_127_3477_n2970), .Y(n150) );
  AND2X1_HVT U383 ( .A1(n142), .A2(n151), .Y(DP_OP_425J2_127_3477_n2948) );
  INVX2_HVT U384 ( .A(DP_OP_425J2_127_3477_n2972), .Y(n151) );
  AND2X1_HVT U385 ( .A1(n142), .A2(n152), .Y(DP_OP_423J2_125_3477_n2948) );
  INVX2_HVT U386 ( .A(DP_OP_422J2_124_3477_n2048), .Y(n152) );
  AND2X1_HVT U387 ( .A1(n142), .A2(n153), .Y(DP_OP_423J2_125_3477_n2951) );
  INVX2_HVT U388 ( .A(DP_OP_424J2_126_3477_n2887), .Y(n153) );
  AND2X4_HVT U389 ( .A1(n142), .A2(n154), .Y(DP_OP_425J2_127_3477_n2951) );
  INVX2_HVT U390 ( .A(DP_OP_424J2_126_3477_n2051), .Y(n154) );
  NAND2X0_HVT U391 ( .A1(n182), .A2(n163), .Y(n161) );
  AO21X1_HVT U392 ( .A1(n158), .A2(n1769), .A3(n155), .Y(n1275) );
  NAND2X0_HVT U393 ( .A1(n156), .A2(n162), .Y(n155) );
  NAND2X0_HVT U394 ( .A1(n1769), .A2(n157), .Y(n156) );
  INVX2_HVT U395 ( .A(n163), .Y(n157) );
  INVX2_HVT U396 ( .A(n27), .Y(n158) );
  NAND2X0_HVT U397 ( .A1(n161), .A2(n159), .Y(n1276) );
  AND2X1_HVT U398 ( .A1(n1769), .A2(n160), .Y(n159) );
  INVX2_HVT U399 ( .A(n162), .Y(n160) );
  NAND2X0_HVT U400 ( .A1(n1756), .A2(DP_OP_424J2_126_3477_n38), .Y(n162) );
  INVX2_HVT U401 ( .A(n164), .Y(n163) );
  NAND2X0_HVT U402 ( .A1(DP_OP_424J2_126_3477_n49), .A2(n1758), .Y(n164) );
  NBUFFX2_HVT U403 ( .A(conv_weight_box[30]), .Y(n165) );
  NBUFFX2_HVT U404 ( .A(conv_weight_box[30]), .Y(n166) );
  NAND2X0_HVT U405 ( .A1(n165), .A2(n167), .Y(DP_OP_422J2_124_3477_n2214) );
  INVX2_HVT U406 ( .A(DP_OP_422J2_124_3477_n2222), .Y(n167) );
  AND2X1_HVT U407 ( .A1(n166), .A2(n168), .Y(DP_OP_422J2_124_3477_n2216) );
  INVX2_HVT U408 ( .A(DP_OP_422J2_124_3477_n2224), .Y(n168) );
  AND2X1_HVT U409 ( .A1(n166), .A2(n169), .Y(DP_OP_422J2_124_3477_n2219) );
  INVX2_HVT U410 ( .A(DP_OP_425J2_127_3477_n2359), .Y(n169) );
  AND2X1_HVT U411 ( .A1(n165), .A2(n170), .Y(DP_OP_422J2_124_3477_n2215) );
  INVX2_HVT U412 ( .A(DP_OP_422J2_124_3477_n2223), .Y(n170) );
  AND2X1_HVT U413 ( .A1(n166), .A2(n171), .Y(DP_OP_424J2_126_3477_n2220) );
  INVX2_HVT U414 ( .A(DP_OP_423J2_125_3477_n2140), .Y(n171) );
  AND2X1_HVT U415 ( .A1(n166), .A2(n172), .Y(DP_OP_422J2_124_3477_n2220) );
  INVX2_HVT U416 ( .A(DP_OP_424J2_126_3477_n2712), .Y(n172) );
  AND2X1_HVT U417 ( .A1(n166), .A2(n173), .Y(DP_OP_422J2_124_3477_n2218) );
  INVX2_HVT U418 ( .A(DP_OP_423J2_125_3477_n2798), .Y(n173) );
  AND2X1_HVT U419 ( .A1(n166), .A2(n174), .Y(DP_OP_422J2_124_3477_n2217) );
  INVX2_HVT U420 ( .A(DP_OP_422J2_124_3477_n2225), .Y(n174) );
  AND2X1_HVT U421 ( .A1(n166), .A2(n175), .Y(DP_OP_424J2_126_3477_n2218) );
  INVX2_HVT U422 ( .A(DP_OP_422J2_124_3477_n2930), .Y(n175) );
  AND2X1_HVT U423 ( .A1(n166), .A2(n176), .Y(DP_OP_424J2_126_3477_n2221) );
  INVX2_HVT U424 ( .A(DP_OP_425J2_127_3477_n2801), .Y(n176) );
  AND2X4_HVT U425 ( .A1(n166), .A2(n177), .Y(DP_OP_422J2_124_3477_n2221) );
  INVX2_HVT U426 ( .A(DP_OP_423J2_125_3477_n2801), .Y(n177) );
  INVX4_HVT U427 ( .A(n1396), .Y(n1485) );
  INVX2_HVT U428 ( .A(conv1_sram_rdata_weight[27]), .Y(n178) );
  INVX4_HVT U429 ( .A(n179), .Y(DP_OP_423J2_125_3477_n2804) );
  AO22X1_HVT U430 ( .A1(n857), .A2(conv1_sram_rdata_weight[49]), .A3(n324), 
        .A4(conv2_sram_rdata_weight[49]), .Y(n179) );
  NAND2X0_HVT U431 ( .A1(n179), .A2(n323), .Y(n322) );
  NBUFFX2_HVT U432 ( .A(n181), .Y(n180) );
  OR2X1_HVT U433 ( .A1(n181), .A2(n808), .Y(n1792) );
  OA21X1_HVT U434 ( .A1(n180), .A2(n1098), .A3(DP_OP_425J2_127_3477_n240), .Y(
        n1099) );
  XOR2X1_HVT U435 ( .A1(n1179), .A2(n180), .Y(n_conv2_sum_d[8]) );
  OA21X1_HVT U436 ( .A1(n810), .A2(DP_OP_425J2_127_3477_n245), .A3(
        DP_OP_425J2_127_3477_n244), .Y(n181) );
  NBUFFX4_HVT U437 ( .A(n1518), .Y(n182) );
  NAND2X0_HVT U438 ( .A1(n1722), .A2(n183), .Y(n1112) );
  INVX2_HVT U439 ( .A(n1754), .Y(n183) );
  XOR3X2_HVT U440 ( .A1(DP_OP_423J2_125_3477_n359), .A2(
        DP_OP_423J2_125_3477_n382), .A3(DP_OP_423J2_125_3477_n380), .Y(
        DP_OP_423J2_125_3477_n355) );
  INVX2_HVT U441 ( .A(conv_weight_box[59]), .Y(DP_OP_422J2_124_3477_n2450) );
  NAND2X0_HVT U442 ( .A1(conv_weight_box[59]), .A2(n184), .Y(
        DP_OP_422J2_124_3477_n2416) );
  INVX2_HVT U443 ( .A(DP_OP_422J2_124_3477_n2448), .Y(n184) );
  MUX21X1_HVT U444 ( .A1(conv1_sram_rdata_weight[87]), .A2(
        conv2_sram_rdata_weight[87]), .S0(n1396), .Y(conv_weight_box[59]) );
  NBUFFX2_HVT U445 ( .A(DP_OP_424J2_126_3477_n2584), .Y(n185) );
  NBUFFX16_HVT U446 ( .A(DP_OP_424J2_126_3477_n2584), .Y(n186) );
  OA21X2_HVT U447 ( .A1(n857), .A2(n188), .A3(n187), .Y(
        DP_OP_424J2_126_3477_n2584) );
  NAND2X0_HVT U448 ( .A1(n857), .A2(conv1_sram_rdata_weight[89]), .Y(n187) );
  INVX2_HVT U449 ( .A(conv2_sram_rdata_weight[89]), .Y(n188) );
  NAND3X1_HVT U450 ( .A1(n190), .A2(n189), .A3(n2045), .Y(n488) );
  NAND2X0_HVT U451 ( .A1(n490), .A2(n489), .Y(n189) );
  NAND4X0_HVT U452 ( .A1(n1955), .A2(n1954), .A3(n1876), .A4(n1965), .Y(n190)
         );
  OR2X1_HVT U453 ( .A1(DP_OP_423J2_125_3477_n1018), .A2(
        DP_OP_423J2_125_3477_n823), .Y(n1665) );
  XOR3X2_HVT U454 ( .A1(DP_OP_423J2_125_3477_n827), .A2(
        DP_OP_423J2_125_3477_n1020), .A3(DP_OP_423J2_125_3477_n825), .Y(
        DP_OP_423J2_125_3477_n823) );
  AO21X1_HVT U455 ( .A1(DP_OP_423J2_125_3477_n250), .A2(
        DP_OP_423J2_125_3477_n295), .A3(n191), .Y(n1666) );
  INVX2_HVT U456 ( .A(DP_OP_423J2_125_3477_n249), .Y(n191) );
  NAND2X0_HVT U457 ( .A1(DP_OP_423J2_125_3477_n1019), .A2(
        DP_OP_423J2_125_3477_n1021), .Y(DP_OP_423J2_125_3477_n249) );
  OR2X1_HVT U458 ( .A1(DP_OP_423J2_125_3477_n1021), .A2(
        DP_OP_423J2_125_3477_n1019), .Y(DP_OP_423J2_125_3477_n295) );
  AO21X1_HVT U459 ( .A1(n1635), .A2(n1636), .A3(n192), .Y(
        DP_OP_423J2_125_3477_n250) );
  INVX2_HVT U460 ( .A(DP_OP_423J2_125_3477_n252), .Y(n192) );
  INVX2_HVT U461 ( .A(n1961), .Y(N7) );
  MUX21X1_HVT U462 ( .A1(conv2_sum_c[9]), .A2(conv2_sum_d[9]), .S0(n1961), .Y(
        tmp_big2[9]) );
  AND2X1_HVT U463 ( .A1(n194), .A2(n193), .Y(n1961) );
  OA21X1_HVT U464 ( .A1(n1920), .A2(n1962), .A3(n2104), .Y(n193) );
  NAND3X0_HVT U465 ( .A1(n1921), .A2(n1963), .A3(n1922), .Y(n194) );
  INVX2_HVT U466 ( .A(mode[0]), .Y(n1516) );
  INVX4_HVT U467 ( .A(n196), .Y(DP_OP_423J2_125_3477_n2892) );
  AO21X1_HVT U468 ( .A1(n335), .A2(conv1_sram_rdata_weight[33]), .A3(n334), 
        .Y(n196) );
  NBUFFX2_HVT U469 ( .A(n196), .Y(n195) );
  AND2X1_HVT U470 ( .A1(n195), .A2(src_window[72]), .Y(
        DP_OP_425J2_127_3477_n2873) );
  AND2X4_HVT U471 ( .A1(n195), .A2(n333), .Y(n1116) );
  NBUFFX2_HVT U472 ( .A(n1484), .Y(n197) );
  AND2X4_HVT U473 ( .A1(n1484), .A2(n198), .Y(DP_OP_425J2_127_3477_n1930) );
  INVX4_HVT U474 ( .A(n1284), .Y(n198) );
  AND2X1_HVT U475 ( .A1(n1484), .A2(n199), .Y(DP_OP_424J2_126_3477_n510) );
  INVX2_HVT U476 ( .A(n1860), .Y(n199) );
  AND2X1_HVT U477 ( .A1(n197), .A2(n200), .Y(DP_OP_423J2_125_3477_n1925) );
  INVX2_HVT U478 ( .A(n1857), .Y(n200) );
  AND2X1_HVT U479 ( .A1(n197), .A2(n201), .Y(DP_OP_424J2_126_3477_n328) );
  INVX2_HVT U480 ( .A(n1906), .Y(n201) );
  AND2X1_HVT U481 ( .A1(n197), .A2(n202), .Y(DP_OP_422J2_124_3477_n328) );
  INVX2_HVT U482 ( .A(n1899), .Y(n202) );
  AND2X1_HVT U483 ( .A1(n197), .A2(n203), .Y(DP_OP_425J2_127_3477_n326) );
  INVX2_HVT U484 ( .A(n1306), .Y(n203) );
  AND2X1_HVT U485 ( .A1(n197), .A2(n204), .Y(DP_OP_422J2_124_3477_n312) );
  INVX2_HVT U486 ( .A(n1903), .Y(n204) );
  AND2X1_HVT U487 ( .A1(n197), .A2(n205), .Y(DP_OP_425J2_127_3477_n316) );
  INVX2_HVT U488 ( .A(n1297), .Y(n205) );
  AND2X1_HVT U489 ( .A1(n197), .A2(n206), .Y(DP_OP_424J2_126_3477_n310) );
  INVX2_HVT U490 ( .A(n1896), .Y(n206) );
  AND2X1_HVT U491 ( .A1(n197), .A2(n207), .Y(DP_OP_422J2_124_3477_n308) );
  INVX2_HVT U492 ( .A(n1882), .Y(n207) );
  NAND2X0_HVT U493 ( .A1(n197), .A2(n208), .Y(n1383) );
  INVX2_HVT U494 ( .A(n1890), .Y(n208) );
  NAND2X0_HVT U495 ( .A1(n197), .A2(n209), .Y(n1834) );
  INVX2_HVT U496 ( .A(n1915), .Y(n209) );
  NBUFFX2_HVT U497 ( .A(n215), .Y(n210) );
  NBUFFX2_HVT U498 ( .A(n215), .Y(n211) );
  NBUFFX2_HVT U499 ( .A(n215), .Y(n212) );
  NBUFFX8_HVT U500 ( .A(n215), .Y(n213) );
  NBUFFX2_HVT U501 ( .A(DP_OP_422J2_124_3477_n3064), .Y(n214) );
  NBUFFX16_HVT U502 ( .A(DP_OP_422J2_124_3477_n3064), .Y(n215) );
  NAND2X0_HVT U503 ( .A1(n4), .A2(conv1_sram_rdata_weight[3]), .Y(n217) );
  NAND2X1_HVT U504 ( .A1(n216), .A2(n849), .Y(DP_OP_424J2_126_3477_n1728) );
  NAND2X0_HVT U505 ( .A1(n216), .A2(src_window[51]), .Y(
        DP_OP_423J2_125_3477_n3029) );
  INVX4_HVT U506 ( .A(DP_OP_422J2_124_3477_n3064), .Y(n216) );
  OA21X2_HVT U507 ( .A1(n4), .A2(n218), .A3(n217), .Y(
        DP_OP_422J2_124_3477_n3064) );
  INVX4_HVT U508 ( .A(conv2_sram_rdata_weight[3]), .Y(n218) );
  OR2X1_HVT U509 ( .A1(n219), .A2(n220), .Y(n1153) );
  NAND2X0_HVT U510 ( .A1(n220), .A2(n219), .Y(n1152) );
  NAND2X0_HVT U511 ( .A1(n1759), .A2(DP_OP_424J2_126_3477_n65), .Y(n219) );
  NAND2X0_HVT U512 ( .A1(n221), .A2(n1761), .Y(n220) );
  NAND2X0_HVT U513 ( .A1(n1518), .A2(DP_OP_424J2_126_3477_n67), .Y(n221) );
  OR2X1_HVT U514 ( .A1(n222), .A2(n223), .Y(n1094) );
  NAND2X0_HVT U515 ( .A1(n223), .A2(n222), .Y(n1093) );
  NAND2X0_HVT U516 ( .A1(n1764), .A2(DP_OP_424J2_126_3477_n120), .Y(n222) );
  NAND2X0_HVT U517 ( .A1(n224), .A2(n1741), .Y(n223) );
  NAND2X0_HVT U518 ( .A1(n1518), .A2(DP_OP_424J2_126_3477_n122), .Y(n224) );
  XOR3X2_HVT U519 ( .A1(DP_OP_423J2_125_3477_n876), .A2(
        DP_OP_423J2_125_3477_n878), .A3(DP_OP_423J2_125_3477_n711), .Y(
        DP_OP_423J2_125_3477_n687) );
  XOR3X2_HVT U520 ( .A1(DP_OP_423J2_125_3477_n749), .A2(n832), .A3(n831), .Y(
        DP_OP_423J2_125_3477_n711) );
  AND3X1_HVT U521 ( .A1(n1230), .A2(n1708), .A3(n1707), .Y(n832) );
  AND2X1_HVT U522 ( .A1(conv_weight_box[63]), .A2(n225), .Y(
        DP_OP_424J2_126_3477_n2475) );
  INVX2_HVT U523 ( .A(DP_OP_424J2_126_3477_n2491), .Y(n225) );
  AND2X1_HVT U524 ( .A1(conv_weight_box[63]), .A2(n226), .Y(
        DP_OP_422J2_124_3477_n2476) );
  INVX2_HVT U525 ( .A(DP_OP_423J2_125_3477_n2536), .Y(n226) );
  AND2X1_HVT U526 ( .A1(conv_weight_box[63]), .A2(n227), .Y(
        DP_OP_424J2_126_3477_n2476) );
  INVX2_HVT U527 ( .A(DP_OP_423J2_125_3477_n2404), .Y(n227) );
  AND2X1_HVT U528 ( .A1(conv_weight_box[63]), .A2(n228), .Y(
        DP_OP_423J2_125_3477_n2472) );
  INVX2_HVT U529 ( .A(DP_OP_422J2_124_3477_n2576), .Y(n228) );
  AND2X1_HVT U530 ( .A1(conv_weight_box[63]), .A2(n229), .Y(
        DP_OP_422J2_124_3477_n2474) );
  INVX2_HVT U531 ( .A(DP_OP_422J2_124_3477_n2490), .Y(n229) );
  AND2X1_HVT U532 ( .A1(conv_weight_box[63]), .A2(n230), .Y(
        DP_OP_422J2_124_3477_n2471) );
  INVX2_HVT U533 ( .A(DP_OP_423J2_125_3477_n2531), .Y(n230) );
  AND2X1_HVT U534 ( .A1(conv_weight_box[63]), .A2(n231), .Y(
        DP_OP_425J2_127_3477_n2476) );
  INVX2_HVT U535 ( .A(DP_OP_424J2_126_3477_n2580), .Y(n231) );
  AND2X1_HVT U536 ( .A1(conv_weight_box[63]), .A2(n232), .Y(
        DP_OP_424J2_126_3477_n2477) );
  INVX2_HVT U537 ( .A(DP_OP_422J2_124_3477_n2669), .Y(n232) );
  AND2X1_HVT U538 ( .A1(conv_weight_box[63]), .A2(n233), .Y(
        DP_OP_425J2_127_3477_n2472) );
  INVX2_HVT U539 ( .A(DP_OP_424J2_126_3477_n2576), .Y(n233) );
  AND2X1_HVT U540 ( .A1(conv_weight_box[63]), .A2(n234), .Y(
        DP_OP_422J2_124_3477_n2477) );
  INVX2_HVT U541 ( .A(DP_OP_423J2_125_3477_n2537), .Y(n234) );
  AND2X1_HVT U542 ( .A1(conv_weight_box[63]), .A2(n235), .Y(
        DP_OP_424J2_126_3477_n2472) );
  INVX2_HVT U543 ( .A(DP_OP_423J2_125_3477_n2400), .Y(n235) );
  AND2X1_HVT U544 ( .A1(conv_weight_box[63]), .A2(n236), .Y(
        DP_OP_425J2_127_3477_n2471) );
  INVX2_HVT U545 ( .A(DP_OP_424J2_126_3477_n2575), .Y(n236) );
  INVX2_HVT U546 ( .A(n856), .Y(n237) );
  NAND2X0_HVT U547 ( .A1(n1351), .A2(n238), .Y(n1114) );
  AND2X1_HVT U548 ( .A1(n1352), .A2(n239), .Y(n238) );
  AND2X1_HVT U549 ( .A1(DP_OP_424J2_126_3477_n274), .A2(
        DP_OP_424J2_126_3477_n78), .Y(n239) );
  NAND2X0_HVT U550 ( .A1(n1518), .A2(DP_OP_424J2_126_3477_n80), .Y(n1351) );
  OR2X2_HVT U551 ( .A1(mode[0]), .A2(n951), .Y(n768) );
  NBUFFX2_HVT U552 ( .A(n768), .Y(n240) );
  NBUFFX16_HVT U553 ( .A(n768), .Y(n241) );
  FADDX1_HVT U554 ( .A(DP_OP_425J2_127_3477_n867), .B(
        DP_OP_425J2_127_3477_n863), .CI(DP_OP_425J2_127_3477_n1048), .CO(
        DP_OP_425J2_127_3477_n844) );
  XOR3X2_HVT U555 ( .A1(DP_OP_425J2_127_3477_n863), .A2(
        DP_OP_425J2_127_3477_n867), .A3(DP_OP_425J2_127_3477_n1048), .Y(
        DP_OP_425J2_127_3477_n845) );
  NBUFFX2_HVT U556 ( .A(n1518), .Y(n242) );
  NAND2X0_HVT U557 ( .A1(n1349), .A2(n243), .Y(n1227) );
  AND2X1_HVT U558 ( .A1(n1348), .A2(n244), .Y(n243) );
  INVX2_HVT U559 ( .A(n245), .Y(n244) );
  NAND2X0_HVT U560 ( .A1(DP_OP_424J2_126_3477_n276), .A2(
        DP_OP_424J2_126_3477_n98), .Y(n245) );
  NAND2X0_HVT U561 ( .A1(n1518), .A2(DP_OP_424J2_126_3477_n100), .Y(n1349) );
  INVX2_HVT U562 ( .A(n246), .Y(n1204) );
  AO21X1_HVT U563 ( .A1(n1203), .A2(n1291), .A3(n1523), .Y(n246) );
  NAND2X0_HVT U564 ( .A1(n247), .A2(n890), .Y(n1291) );
  NAND2X0_HVT U565 ( .A1(n248), .A2(n892), .Y(n247) );
  AND2X1_HVT U566 ( .A1(n1611), .A2(n1612), .Y(n892) );
  INVX2_HVT U567 ( .A(n71), .Y(n248) );
  NAND2X0_HVT U568 ( .A1(n620), .A2(n249), .Y(DP_OP_422J2_124_3477_n2082) );
  INVX2_HVT U569 ( .A(DP_OP_422J2_124_3477_n2090), .Y(n249) );
  AND2X1_HVT U570 ( .A1(n620), .A2(n250), .Y(DP_OP_422J2_124_3477_n2083) );
  INVX2_HVT U571 ( .A(DP_OP_422J2_124_3477_n2091), .Y(n250) );
  AND2X1_HVT U572 ( .A1(n620), .A2(n251), .Y(DP_OP_424J2_126_3477_n2087) );
  INVX2_HVT U573 ( .A(DP_OP_424J2_126_3477_n2095), .Y(n251) );
  AND2X1_HVT U574 ( .A1(n620), .A2(n252), .Y(DP_OP_424J2_126_3477_n2086) );
  INVX2_HVT U575 ( .A(DP_OP_422J2_124_3477_n3060), .Y(n252) );
  AND2X1_HVT U576 ( .A1(n620), .A2(n253), .Y(DP_OP_424J2_126_3477_n2088) );
  INVX2_HVT U577 ( .A(DP_OP_423J2_125_3477_n2008), .Y(n253) );
  OR2X1_HVT U578 ( .A1(DP_OP_422J2_124_3477_n2973), .A2(n254), .Y(
        DP_OP_422J2_124_3477_n2941) );
  OR2X1_HVT U579 ( .A1(DP_OP_424J2_126_3477_n2185), .A2(n254), .Y(
        DP_OP_422J2_124_3477_n2945) );
  OR2X1_HVT U580 ( .A1(DP_OP_422J2_124_3477_n2974), .A2(n254), .Y(
        DP_OP_422J2_124_3477_n2942) );
  OR2X1_HVT U581 ( .A1(DP_OP_424J2_126_3477_n2184), .A2(n254), .Y(
        DP_OP_422J2_124_3477_n2944) );
  OR2X4_HVT U582 ( .A1(DP_OP_424J2_126_3477_n2976), .A2(n254), .Y(
        DP_OP_424J2_126_3477_n2944) );
  AND2X1_HVT U583 ( .A1(n257), .A2(n255), .Y(DP_OP_422J2_124_3477_n2938) );
  INVX2_HVT U584 ( .A(DP_OP_422J2_124_3477_n2970), .Y(n255) );
  AND2X1_HVT U585 ( .A1(n257), .A2(n256), .Y(DP_OP_424J2_126_3477_n2938) );
  INVX2_HVT U586 ( .A(DP_OP_424J2_126_3477_n2970), .Y(n256) );
  FADDX1_HVT U587 ( .A(DP_OP_425J2_127_3477_n2834), .B(n258), .CI(
        DP_OP_425J2_127_3477_n2475), .CO(DP_OP_425J2_127_3477_n1674) );
  INVX2_HVT U588 ( .A(n260), .Y(n258) );
  XOR3X2_HVT U589 ( .A1(n260), .A2(DP_OP_425J2_127_3477_n2834), .A3(n259), .Y(
        DP_OP_425J2_127_3477_n1675) );
  INVX2_HVT U590 ( .A(DP_OP_425J2_127_3477_n2475), .Y(n259) );
  OR2X1_HVT U591 ( .A1(DP_OP_425J2_127_3477_n2404), .A2(n798), .Y(n260) );
  NBUFFX2_HVT U592 ( .A(n789), .Y(n261) );
  NBUFFX2_HVT U593 ( .A(n346), .Y(n262) );
  NBUFFX2_HVT U594 ( .A(n346), .Y(n263) );
  INVX2_HVT U595 ( .A(n346), .Y(n789) );
  AND2X1_HVT U596 ( .A1(n263), .A2(n349), .Y(DP_OP_422J2_124_3477_n2425) );
  AND2X1_HVT U597 ( .A1(n263), .A2(n751), .Y(DP_OP_422J2_124_3477_n2424) );
  AND2X4_HVT U598 ( .A1(n263), .A2(n752), .Y(DP_OP_423J2_125_3477_n2419) );
  OA21X1_HVT U599 ( .A1(n769), .A2(n754), .A3(n753), .Y(n346) );
  NBUFFX2_HVT U600 ( .A(n1425), .Y(n264) );
  NBUFFX2_HVT U601 ( .A(n1425), .Y(n265) );
  AND2X1_HVT U602 ( .A1(n264), .A2(n266), .Y(DP_OP_425J2_127_3477_n1935) );
  INVX2_HVT U603 ( .A(DP_OP_425J2_127_3477_n1968), .Y(n266) );
  AND2X1_HVT U604 ( .A1(n264), .A2(n267), .Y(DP_OP_422J2_124_3477_n1935) );
  INVX2_HVT U605 ( .A(n1975), .Y(n267) );
  AND2X1_HVT U606 ( .A1(n265), .A2(n268), .Y(DP_OP_424J2_126_3477_n1932) );
  INVX2_HVT U607 ( .A(n1859), .Y(n268) );
  AND2X1_HVT U608 ( .A1(n265), .A2(n269), .Y(DP_OP_422J2_124_3477_n1930) );
  INVX2_HVT U609 ( .A(n1861), .Y(n269) );
  AND2X1_HVT U610 ( .A1(n265), .A2(n270), .Y(DP_OP_424J2_126_3477_n1934) );
  INVX2_HVT U611 ( .A(n1865), .Y(n270) );
  AND2X1_HVT U612 ( .A1(n265), .A2(n271), .Y(DP_OP_423J2_125_3477_n1931) );
  INVX2_HVT U613 ( .A(n1851), .Y(n271) );
  AND2X1_HVT U614 ( .A1(n265), .A2(n272), .Y(DP_OP_422J2_124_3477_n314) );
  INVX2_HVT U615 ( .A(n1888), .Y(n272) );
  AND2X1_HVT U616 ( .A1(n265), .A2(n273), .Y(DP_OP_425J2_127_3477_n314) );
  INVX2_HVT U617 ( .A(n1311), .Y(n273) );
  AND2X1_HVT U618 ( .A1(n265), .A2(n274), .Y(DP_OP_424J2_126_3477_n312) );
  INVX2_HVT U619 ( .A(n1910), .Y(n274) );
  AND2X1_HVT U620 ( .A1(n265), .A2(n275), .Y(DP_OP_424J2_126_3477_n338) );
  INVX2_HVT U621 ( .A(n1891), .Y(n275) );
  AND2X1_HVT U622 ( .A1(n265), .A2(n276), .Y(DP_OP_424J2_126_3477_n304) );
  INVX2_HVT U623 ( .A(n1917), .Y(n276) );
  AND2X4_HVT U624 ( .A1(n265), .A2(n277), .Y(DP_OP_423J2_125_3477_n302) );
  INVX2_HVT U625 ( .A(n1326), .Y(n277) );
  NBUFFX8_HVT U626 ( .A(n1490), .Y(n278) );
  NBUFFX16_HVT U627 ( .A(n1490), .Y(n279) );
  OA21X2_HVT U628 ( .A1(n857), .A2(n281), .A3(n280), .Y(n1490) );
  NAND2X0_HVT U629 ( .A1(n857), .A2(conv1_sram_rdata_weight[73]), .Y(n280) );
  INVX2_HVT U630 ( .A(conv2_sram_rdata_weight[73]), .Y(n281) );
  AND2X1_HVT U631 ( .A1(n282), .A2(n1589), .Y(n1570) );
  NAND3X0_HVT U632 ( .A1(n1574), .A2(n285), .A3(n1576), .Y(n282) );
  AND2X1_HVT U633 ( .A1(n284), .A2(n283), .Y(DP_OP_422J2_124_3477_n233) );
  OA21X1_HVT U634 ( .A1(DP_OP_422J2_124_3477_n240), .A2(
        DP_OP_422J2_124_3477_n236), .A3(DP_OP_422J2_124_3477_n237), .Y(n283)
         );
  NAND2X0_HVT U635 ( .A1(n1593), .A2(DP_OP_422J2_124_3477_n242), .Y(n284) );
  NAND2X0_HVT U636 ( .A1(DP_OP_422J2_124_3477_n219), .A2(n285), .Y(n1545) );
  OR2X1_HVT U637 ( .A1(DP_OP_422J2_124_3477_n209), .A2(
        DP_OP_422J2_124_3477_n214), .Y(n286) );
  AND2X1_HVT U638 ( .A1(n1544), .A2(n1534), .Y(DP_OP_422J2_124_3477_n219) );
  FADDX1_HVT U639 ( .A(DP_OP_424J2_126_3477_n1509), .B(
        DP_OP_424J2_126_3477_n1517), .CI(DP_OP_424J2_126_3477_n1531), .CO(
        DP_OP_424J2_126_3477_n1466) );
  XOR3X2_HVT U640 ( .A1(DP_OP_424J2_126_3477_n1531), .A2(
        DP_OP_424J2_126_3477_n1517), .A3(DP_OP_424J2_126_3477_n1509), .Y(
        DP_OP_424J2_126_3477_n1467) );
  INVX2_HVT U641 ( .A(n1832), .Y(n1781) );
  OR2X1_HVT U642 ( .A1(n289), .A2(DP_OP_425J2_127_3477_n168), .Y(n1455) );
  AND2X1_HVT U643 ( .A1(n287), .A2(n1845), .Y(DP_OP_425J2_127_3477_n168) );
  NAND2X0_HVT U644 ( .A1(n1832), .A2(n288), .Y(n287) );
  INVX2_HVT U645 ( .A(n1837), .Y(n288) );
  INVX2_HVT U646 ( .A(DP_OP_425J2_127_3477_n19), .Y(n289) );
  INVX4_HVT U647 ( .A(conv_weight_box[43]), .Y(DP_OP_425J2_127_3477_n2319) );
  AO22X2_HVT U648 ( .A1(n1485), .A2(conv1_sram_rdata_weight[62]), .A3(n329), 
        .A4(conv2_sram_rdata_weight[62]), .Y(conv_weight_box[43]) );
  AND2X4_HVT U649 ( .A1(conv_weight_box[43]), .A2(n290), .Y(
        DP_OP_424J2_126_3477_n2293) );
  INVX2_HVT U650 ( .A(DP_OP_424J2_126_3477_n2317), .Y(n290) );
  XOR3X2_HVT U651 ( .A1(DP_OP_424J2_126_3477_n827), .A2(
        DP_OP_424J2_126_3477_n1020), .A3(DP_OP_424J2_126_3477_n825), .Y(
        DP_OP_424J2_126_3477_n823) );
  INVX4_HVT U652 ( .A(n342), .Y(DP_OP_423J2_125_3477_n4) );
  XOR2X2_HVT U653 ( .A1(n292), .A2(n291), .Y(n_conv2_sum_b[31]) );
  NAND2X0_HVT U654 ( .A1(n1668), .A2(DP_OP_423J2_125_3477_n38), .Y(n291) );
  OA21X1_HVT U655 ( .A1(n293), .A2(n342), .A3(n1680), .Y(n292) );
  INVX2_HVT U656 ( .A(n1682), .Y(n293) );
  OR2X1_HVT U657 ( .A1(n294), .A2(n295), .Y(n1229) );
  NAND2X0_HVT U658 ( .A1(n295), .A2(n294), .Y(n1228) );
  NAND2X0_HVT U659 ( .A1(n1758), .A2(DP_OP_424J2_126_3477_n47), .Y(n294) );
  NAND2X0_HVT U660 ( .A1(n296), .A2(n1739), .Y(n295) );
  NAND2X0_HVT U661 ( .A1(n1518), .A2(DP_OP_424J2_126_3477_n49), .Y(n296) );
  NBUFFX2_HVT U662 ( .A(conv_weight_box[59]), .Y(n297) );
  NAND2X0_HVT U663 ( .A1(conv_weight_box[59]), .A2(n298), .Y(
        DP_OP_423J2_125_3477_n2414) );
  INVX2_HVT U664 ( .A(DP_OP_422J2_124_3477_n2622), .Y(n298) );
  NAND2X0_HVT U665 ( .A1(n297), .A2(n299), .Y(DP_OP_425J2_127_3477_n2416) );
  INVX2_HVT U666 ( .A(DP_OP_425J2_127_3477_n2448), .Y(n299) );
  NAND2X0_HVT U667 ( .A1(conv_weight_box[59]), .A2(n300), .Y(
        DP_OP_423J2_125_3477_n2416) );
  INVX2_HVT U668 ( .A(DP_OP_423J2_125_3477_n2448), .Y(n300) );
  NAND2X0_HVT U669 ( .A1(n297), .A2(n301), .Y(DP_OP_423J2_125_3477_n2417) );
  INVX2_HVT U670 ( .A(DP_OP_422J2_124_3477_n2625), .Y(n301) );
  NAND2X0_HVT U671 ( .A1(n297), .A2(n302), .Y(DP_OP_425J2_127_3477_n2417) );
  INVX2_HVT U672 ( .A(DP_OP_425J2_127_3477_n2449), .Y(n302) );
  NAND2X0_HVT U673 ( .A1(n297), .A2(n303), .Y(DP_OP_425J2_127_3477_n2412) );
  INVX2_HVT U674 ( .A(DP_OP_423J2_125_3477_n2708), .Y(n303) );
  NAND2X0_HVT U675 ( .A1(n297), .A2(n304), .Y(DP_OP_423J2_125_3477_n2415) );
  INVX2_HVT U676 ( .A(DP_OP_423J2_125_3477_n2447), .Y(n304) );
  NAND2X0_HVT U677 ( .A1(n297), .A2(n305), .Y(DP_OP_423J2_125_3477_n2411) );
  INVX2_HVT U678 ( .A(DP_OP_422J2_124_3477_n2619), .Y(n305) );
  NAND2X0_HVT U679 ( .A1(n297), .A2(n306), .Y(DP_OP_425J2_127_3477_n2411) );
  INVX2_HVT U680 ( .A(DP_OP_424J2_126_3477_n2619), .Y(n306) );
  NAND2X0_HVT U681 ( .A1(n297), .A2(n307), .Y(DP_OP_423J2_125_3477_n2413) );
  INVX2_HVT U682 ( .A(DP_OP_422J2_124_3477_n2621), .Y(n307) );
  NAND2X0_HVT U683 ( .A1(n297), .A2(n308), .Y(DP_OP_423J2_125_3477_n2412) );
  INVX2_HVT U684 ( .A(DP_OP_422J2_124_3477_n2620), .Y(n308) );
  AND2X4_HVT U685 ( .A1(n297), .A2(n309), .Y(DP_OP_423J2_125_3477_n2410) );
  INVX2_HVT U686 ( .A(DP_OP_422J2_124_3477_n2618), .Y(n309) );
  XOR3X2_HVT U687 ( .A1(DP_OP_422J2_124_3477_n1246), .A2(
        DP_OP_422J2_124_3477_n1248), .A3(DP_OP_422J2_124_3477_n1250), .Y(
        DP_OP_422J2_124_3477_n1045) );
  AO22X1_HVT U688 ( .A1(DP_OP_422J2_124_3477_n1448), .A2(
        DP_OP_422J2_124_3477_n1281), .A3(n310), .A4(n1232), .Y(
        DP_OP_422J2_124_3477_n1248) );
  OR2X1_HVT U689 ( .A1(DP_OP_422J2_124_3477_n1448), .A2(
        DP_OP_422J2_124_3477_n1281), .Y(n310) );
  INVX2_HVT U690 ( .A(conv_weight_box[47]), .Y(DP_OP_425J2_127_3477_n2365) );
  INVX2_HVT U691 ( .A(n1363), .Y(n1337) );
  FADDX1_HVT U692 ( .A(n1233), .B(DP_OP_425J2_127_3477_n1727), .CI(
        DP_OP_425J2_127_3477_n1675), .CO(DP_OP_425J2_127_3477_n1636) );
  XOR3X2_HVT U693 ( .A1(DP_OP_425J2_127_3477_n2864), .A2(
        DP_OP_425J2_127_3477_n2350), .A3(DP_OP_425J2_127_3477_n2871), .Y(n1233) );
  AND2X1_HVT U694 ( .A1(conv_weight_box[47]), .A2(n311), .Y(
        DP_OP_425J2_127_3477_n2350) );
  INVX2_HVT U695 ( .A(DP_OP_425J2_127_3477_n2358), .Y(n311) );
  XOR3X2_HVT U696 ( .A1(n571), .A2(DP_OP_425J2_127_3477_n2505), .A3(n570), .Y(
        DP_OP_425J2_127_3477_n1727) );
  NAND2X0_HVT U697 ( .A1(n1363), .A2(n312), .Y(DP_OP_425J2_127_3477_n2505) );
  INVX2_HVT U698 ( .A(DP_OP_423J2_125_3477_n2405), .Y(n312) );
  OA21X1_HVT U699 ( .A1(n315), .A2(n314), .A3(n313), .Y(n327) );
  NAND3X0_HVT U700 ( .A1(n1485), .A2(conv1_sram_rdata_weight[62]), .A3(n328), 
        .Y(n313) );
  INVX2_HVT U701 ( .A(n329), .Y(n314) );
  NAND2X0_HVT U702 ( .A1(n328), .A2(conv2_sram_rdata_weight[62]), .Y(n315) );
  NBUFFX2_HVT U703 ( .A(DP_OP_425J2_127_3477_n2319), .Y(n316) );
  NBUFFX2_HVT U704 ( .A(DP_OP_425J2_127_3477_n2319), .Y(n317) );
  INVX2_HVT U705 ( .A(conv_weight_box[36]), .Y(DP_OP_424J2_126_3477_n2277) );
  AO22X1_HVT U706 ( .A1(n321), .A2(n325), .A3(n320), .A4(n318), .Y(
        DP_OP_424J2_126_3477_n1346) );
  NAND2X0_HVT U707 ( .A1(n319), .A2(n322), .Y(n318) );
  INVX2_HVT U708 ( .A(n325), .Y(n319) );
  INVX2_HVT U709 ( .A(n327), .Y(n320) );
  INVX2_HVT U710 ( .A(n322), .Y(n321) );
  XOR3X1_HVT U711 ( .A1(n327), .A2(n325), .A3(n322), .Y(
        DP_OP_424J2_126_3477_n1347) );
  INVX4_HVT U712 ( .A(DP_OP_425J2_127_3477_n2269), .Y(n323) );
  INVX1_HVT U713 ( .A(n857), .Y(n324) );
  AND2X2_HVT U714 ( .A1(conv_weight_box[36]), .A2(n326), .Y(n325) );
  INVX4_HVT U715 ( .A(DP_OP_424J2_126_3477_n2268), .Y(n326) );
  INVX4_HVT U716 ( .A(DP_OP_425J2_127_3477_n2710), .Y(n328) );
  NAND2X0_HVT U717 ( .A1(n726), .A2(n739), .Y(n737) );
  AND2X1_HVT U718 ( .A1(n726), .A2(n740), .Y(DP_OP_422J2_124_3477_n2729) );
  INVX2_HVT U719 ( .A(conv_weight_box[22]), .Y(DP_OP_423J2_125_3477_n2891) );
  AO22X1_HVT U720 ( .A1(n1116), .A2(n1115), .A3(n1117), .A4(n330), .Y(
        DP_OP_423J2_125_3477_n1784) );
  OR2X1_HVT U721 ( .A1(n1116), .A2(n1115), .Y(n330) );
  AND2X1_HVT U722 ( .A1(conv_weight_box[22]), .A2(n331), .Y(n1115) );
  INVX2_HVT U723 ( .A(DP_OP_423J2_125_3477_n2889), .Y(n331) );
  AO21X1_HVT U724 ( .A1(conv1_sram_rdata_weight[34]), .A2(n335), .A3(n332), 
        .Y(conv_weight_box[22]) );
  AND2X1_HVT U725 ( .A1(n1396), .A2(conv2_sram_rdata_weight[34]), .Y(n332) );
  INVX2_HVT U726 ( .A(DP_OP_422J2_124_3477_n2140), .Y(n333) );
  AND2X1_HVT U727 ( .A1(n1396), .A2(conv2_sram_rdata_weight[33]), .Y(n334) );
  INVX2_HVT U728 ( .A(n1396), .Y(n335) );
  NAND2X0_HVT U729 ( .A1(n1374), .A2(n336), .Y(n1274) );
  AND2X1_HVT U730 ( .A1(n1744), .A2(n337), .Y(n336) );
  INVX2_HVT U731 ( .A(n338), .Y(n337) );
  NAND2X0_HVT U732 ( .A1(n1763), .A2(DP_OP_424J2_126_3477_n89), .Y(n338) );
  NAND2X0_HVT U733 ( .A1(n1518), .A2(DP_OP_424J2_126_3477_n91), .Y(n1374) );
  OR2X1_HVT U734 ( .A1(n339), .A2(n340), .Y(n1190) );
  NAND2X0_HVT U735 ( .A1(n340), .A2(n339), .Y(n1189) );
  NAND2X0_HVT U736 ( .A1(DP_OP_424J2_126_3477_n272), .A2(
        DP_OP_424J2_126_3477_n52), .Y(n339) );
  NAND2X0_HVT U737 ( .A1(n341), .A2(DP_OP_424J2_126_3477_n57), .Y(n340) );
  NAND2X0_HVT U738 ( .A1(n1518), .A2(DP_OP_424J2_126_3477_n54), .Y(n341) );
  NAND3X0_HVT U739 ( .A1(n1657), .A2(n1658), .A3(n343), .Y(n1251) );
  AND2X2_HVT U740 ( .A1(DP_OP_423J2_125_3477_n279), .A2(
        DP_OP_423J2_125_3477_n129), .Y(n343) );
  NAND2X0_HVT U741 ( .A1(DP_OP_423J2_125_3477_n4), .A2(
        DP_OP_423J2_125_3477_n131), .Y(n1657) );
  AND3X1_HVT U742 ( .A1(n1393), .A2(n1392), .A3(n1675), .Y(n342) );
  INVX4_HVT U743 ( .A(n344), .Y(n345) );
  INVX2_HVT U744 ( .A(n423), .Y(n344) );
  MUX21X2_HVT U745 ( .A1(conv2_sram_rdata_weight[60]), .A2(
        conv1_sram_rdata_weight[60]), .S0(n345), .Y(conv_weight_box[41]) );
  AND2X1_HVT U746 ( .A1(n262), .A2(n347), .Y(DP_OP_424J2_126_3477_n2423) );
  INVX2_HVT U747 ( .A(DP_OP_424J2_126_3477_n2447), .Y(n347) );
  AND2X1_HVT U748 ( .A1(n262), .A2(n348), .Y(DP_OP_424J2_126_3477_n2425) );
  INVX2_HVT U749 ( .A(DP_OP_423J2_125_3477_n2361), .Y(n348) );
  INVX4_HVT U750 ( .A(DP_OP_423J2_125_3477_n2581), .Y(n349) );
  AND2X1_HVT U751 ( .A1(n263), .A2(n350), .Y(DP_OP_424J2_126_3477_n2420) );
  INVX2_HVT U752 ( .A(DP_OP_425J2_127_3477_n2576), .Y(n350) );
  AND2X1_HVT U753 ( .A1(n263), .A2(n351), .Y(DP_OP_422J2_124_3477_n2421) );
  INVX2_HVT U754 ( .A(DP_OP_422J2_124_3477_n2445), .Y(n351) );
  AND2X1_HVT U755 ( .A1(n263), .A2(n352), .Y(DP_OP_424J2_126_3477_n2424) );
  INVX2_HVT U756 ( .A(DP_OP_422J2_124_3477_n2712), .Y(n352) );
  AND2X1_HVT U757 ( .A1(n263), .A2(n353), .Y(DP_OP_424J2_126_3477_n2421) );
  INVX2_HVT U758 ( .A(DP_OP_422J2_124_3477_n2709), .Y(n353) );
  AND2X1_HVT U759 ( .A1(n263), .A2(n354), .Y(DP_OP_424J2_126_3477_n2422) );
  INVX2_HVT U760 ( .A(DP_OP_422J2_124_3477_n2710), .Y(n354) );
  AND2X1_HVT U761 ( .A1(n263), .A2(n355), .Y(DP_OP_424J2_126_3477_n2419) );
  INVX2_HVT U762 ( .A(DP_OP_424J2_126_3477_n2443), .Y(n355) );
  NAND2X0_HVT U763 ( .A1(n263), .A2(n356), .Y(DP_OP_424J2_126_3477_n2418) );
  INVX2_HVT U764 ( .A(DP_OP_425J2_127_3477_n2574), .Y(n356) );
  INVX2_HVT U765 ( .A(n359), .Y(DP_OP_422J2_124_3477_n4) );
  XNOR2X2_HVT U766 ( .A1(n357), .A2(n928), .Y(n_conv2_sum_a[29]) );
  OA21X1_HVT U767 ( .A1(n360), .A2(n359), .A3(n358), .Y(n357) );
  INVX2_HVT U768 ( .A(DP_OP_422J2_124_3477_n55), .Y(n358) );
  OA21X1_HVT U769 ( .A1(n1545), .A2(DP_OP_422J2_124_3477_n233), .A3(n1570), 
        .Y(n359) );
  INVX2_HVT U770 ( .A(DP_OP_422J2_124_3477_n54), .Y(n360) );
  NAND2X0_HVT U771 ( .A1(n361), .A2(DP_OP_422J2_124_3477_n217), .Y(
        DP_OP_422J2_124_3477_n213) );
  NAND2X0_HVT U772 ( .A1(DP_OP_422J2_124_3477_n220), .A2(n362), .Y(n361) );
  INVX2_HVT U773 ( .A(n914), .Y(n362) );
  NAND2X0_HVT U774 ( .A1(n363), .A2(DP_OP_422J2_124_3477_n226), .Y(
        DP_OP_422J2_124_3477_n220) );
  NAND2X0_HVT U775 ( .A1(n6), .A2(n1534), .Y(n363) );
  NBUFFX2_HVT U776 ( .A(DP_OP_423J2_125_3477_n2232), .Y(n364) );
  NBUFFX16_HVT U777 ( .A(DP_OP_423J2_125_3477_n2232), .Y(n365) );
  OA21X2_HVT U778 ( .A1(n345), .A2(n367), .A3(n366), .Y(
        DP_OP_423J2_125_3477_n2232) );
  NAND2X0_HVT U779 ( .A1(n345), .A2(conv1_sram_rdata_weight[45]), .Y(n366) );
  INVX2_HVT U780 ( .A(conv2_sram_rdata_weight[45]), .Y(n367) );
  AND2X1_HVT U781 ( .A1(n1484), .A2(n368), .Y(DP_OP_424J2_126_3477_n1931) );
  INVX2_HVT U782 ( .A(n1854), .Y(n368) );
  AND2X1_HVT U783 ( .A1(n1484), .A2(n369), .Y(DP_OP_422J2_124_3477_n1932) );
  INVX2_HVT U784 ( .A(n1863), .Y(n369) );
  AND2X1_HVT U785 ( .A1(n1484), .A2(n370), .Y(DP_OP_423J2_125_3477_n1927) );
  INVX2_HVT U786 ( .A(n1984), .Y(n370) );
  AND2X1_HVT U787 ( .A1(n1484), .A2(n371), .Y(DP_OP_425J2_127_3477_n1926) );
  INVX2_HVT U788 ( .A(n1986), .Y(n371) );
  NAND2X0_HVT U789 ( .A1(n1484), .A2(n372), .Y(n1381) );
  INVX2_HVT U790 ( .A(n1884), .Y(n372) );
  AND2X1_HVT U791 ( .A1(n1484), .A2(n373), .Y(DP_OP_424J2_126_3477_n324) );
  INVX2_HVT U792 ( .A(n1907), .Y(n373) );
  AND2X1_HVT U793 ( .A1(n1484), .A2(n374), .Y(DP_OP_424J2_126_3477_n330) );
  INVX2_HVT U794 ( .A(n1319), .Y(n374) );
  AND2X1_HVT U795 ( .A1(n1484), .A2(n375), .Y(DP_OP_424J2_126_3477_n314) );
  INVX2_HVT U796 ( .A(n1895), .Y(n375) );
  AND2X1_HVT U797 ( .A1(n1484), .A2(n376), .Y(DP_OP_425J2_127_3477_n338) );
  INVX2_HVT U798 ( .A(n1317), .Y(n376) );
  AND2X1_HVT U799 ( .A1(n1484), .A2(n377), .Y(DP_OP_423J2_125_3477_n310) );
  INVX2_HVT U800 ( .A(n1305), .Y(n377) );
  AND2X1_HVT U801 ( .A1(n1484), .A2(n378), .Y(DP_OP_424J2_126_3477_n308) );
  INVX2_HVT U802 ( .A(n1911), .Y(n378) );
  AND2X1_HVT U803 ( .A1(n1484), .A2(n379), .Y(DP_OP_424J2_126_3477_n302) );
  INVX2_HVT U804 ( .A(n1913), .Y(n379) );
  OR2X1_HVT U805 ( .A1(n380), .A2(n381), .Y(n1050) );
  NAND2X0_HVT U806 ( .A1(n381), .A2(n380), .Y(n1049) );
  NAND2X0_HVT U807 ( .A1(DP_OP_424J2_126_3477_n282), .A2(
        DP_OP_424J2_126_3477_n156), .Y(n380) );
  NAND2X0_HVT U808 ( .A1(n382), .A2(n1748), .Y(n381) );
  NAND2X0_HVT U809 ( .A1(n1518), .A2(n1058), .Y(n382) );
  NBUFFX2_HVT U810 ( .A(n1484), .Y(n383) );
  AND2X1_HVT U811 ( .A1(n1484), .A2(n384), .Y(DP_OP_425J2_127_3477_n1932) );
  INVX2_HVT U812 ( .A(n1283), .Y(n384) );
  AND2X1_HVT U813 ( .A1(n383), .A2(n385), .Y(DP_OP_422J2_124_3477_n1931) );
  INVX2_HVT U814 ( .A(n1852), .Y(n385) );
  AND2X1_HVT U815 ( .A1(n383), .A2(n386), .Y(DP_OP_423J2_125_3477_n1926) );
  INVX2_HVT U816 ( .A(n1524), .Y(n386) );
  AND2X1_HVT U817 ( .A1(n383), .A2(n387), .Y(DP_OP_424J2_126_3477_n1926) );
  INVX2_HVT U818 ( .A(n1982), .Y(n387) );
  AND2X1_HVT U819 ( .A1(n383), .A2(n388), .Y(DP_OP_422J2_124_3477_n324) );
  INVX2_HVT U820 ( .A(n1900), .Y(n388) );
  AND2X1_HVT U821 ( .A1(n383), .A2(n389), .Y(DP_OP_424J2_126_3477_n322) );
  INVX2_HVT U822 ( .A(n1893), .Y(n389) );
  AND2X1_HVT U823 ( .A1(n383), .A2(n390), .Y(DP_OP_422J2_124_3477_n322) );
  INVX2_HVT U824 ( .A(n1886), .Y(n390) );
  AND2X1_HVT U825 ( .A1(n383), .A2(n391), .Y(DP_OP_422J2_124_3477_n338) );
  INVX2_HVT U826 ( .A(n1978), .Y(n391) );
  AND2X1_HVT U827 ( .A1(n383), .A2(n392), .Y(DP_OP_422J2_124_3477_n1923) );
  INVX2_HVT U828 ( .A(n1898), .Y(n392) );
  AND2X4_HVT U829 ( .A1(n383), .A2(n393), .Y(DP_OP_425J2_127_3477_n302) );
  INVX2_HVT U830 ( .A(n1325), .Y(n393) );
  INVX8_HVT U831 ( .A(n423), .Y(n1928) );
  INVX2_HVT U832 ( .A(DP_OP_424J2_126_3477_n2716), .Y(n1378) );
  MUX21X1_HVT U833 ( .A1(n395), .A2(n394), .S0(n423), .Y(
        DP_OP_424J2_126_3477_n2716) );
  INVX2_HVT U834 ( .A(conv1_sram_rdata_weight[65]), .Y(n394) );
  INVX2_HVT U835 ( .A(conv2_sram_rdata_weight[65]), .Y(n395) );
  NBUFFX2_HVT U836 ( .A(conv_weight_box[59]), .Y(n396) );
  NAND2X0_HVT U837 ( .A1(conv_weight_box[59]), .A2(n397), .Y(
        DP_OP_424J2_126_3477_n2415) );
  INVX2_HVT U838 ( .A(DP_OP_424J2_126_3477_n2447), .Y(n397) );
  NAND2X0_HVT U839 ( .A1(n396), .A2(n398), .Y(DP_OP_424J2_126_3477_n2417) );
  INVX2_HVT U840 ( .A(DP_OP_423J2_125_3477_n2361), .Y(n398) );
  NAND2X0_HVT U841 ( .A1(conv_weight_box[59]), .A2(n399), .Y(
        DP_OP_424J2_126_3477_n2416) );
  INVX2_HVT U842 ( .A(DP_OP_425J2_127_3477_n2580), .Y(n399) );
  NAND2X0_HVT U843 ( .A1(n396), .A2(n400), .Y(DP_OP_424J2_126_3477_n2412) );
  INVX2_HVT U844 ( .A(DP_OP_425J2_127_3477_n2576), .Y(n400) );
  NAND2X0_HVT U845 ( .A1(n396), .A2(n401), .Y(DP_OP_424J2_126_3477_n2413) );
  INVX2_HVT U846 ( .A(DP_OP_425J2_127_3477_n2577), .Y(n401) );
  NAND2X0_HVT U847 ( .A1(n396), .A2(n402), .Y(DP_OP_425J2_127_3477_n2414) );
  INVX2_HVT U848 ( .A(DP_OP_424J2_126_3477_n2622), .Y(n402) );
  NAND2X0_HVT U849 ( .A1(n396), .A2(n403), .Y(DP_OP_424J2_126_3477_n2414) );
  INVX2_HVT U850 ( .A(DP_OP_422J2_124_3477_n2710), .Y(n403) );
  NAND2X0_HVT U851 ( .A1(n396), .A2(n404), .Y(DP_OP_425J2_127_3477_n2413) );
  INVX2_HVT U852 ( .A(DP_OP_425J2_127_3477_n2445), .Y(n404) );
  NAND2X0_HVT U853 ( .A1(n396), .A2(n405), .Y(DP_OP_425J2_127_3477_n2415) );
  INVX2_HVT U854 ( .A(DP_OP_425J2_127_3477_n2447), .Y(n405) );
  NAND2X0_HVT U855 ( .A1(n396), .A2(n406), .Y(DP_OP_424J2_126_3477_n2411) );
  INVX2_HVT U856 ( .A(DP_OP_424J2_126_3477_n2443), .Y(n406) );
  AND2X1_HVT U857 ( .A1(n396), .A2(n407), .Y(DP_OP_424J2_126_3477_n2410) );
  INVX2_HVT U858 ( .A(DP_OP_423J2_125_3477_n2354), .Y(n407) );
  AND2X4_HVT U859 ( .A1(n396), .A2(n408), .Y(DP_OP_425J2_127_3477_n2410) );
  INVX2_HVT U860 ( .A(DP_OP_423J2_125_3477_n2706), .Y(n408) );
  NAND2X0_HVT U861 ( .A1(n409), .A2(n1449), .Y(DP_OP_424J2_126_3477_n418) );
  NAND2X0_HVT U862 ( .A1(DP_OP_424J2_126_3477_n421), .A2(n410), .Y(n409) );
  OR2X1_HVT U863 ( .A1(DP_OP_424J2_126_3477_n514), .A2(
        DP_OP_424J2_126_3477_n423), .Y(n410) );
  INVX2_HVT U864 ( .A(DP_OP_424J2_126_3477_n226), .Y(n1067) );
  NAND2X0_HVT U865 ( .A1(DP_OP_424J2_126_3477_n373), .A2(
        DP_OP_424J2_126_3477_n418), .Y(DP_OP_424J2_126_3477_n226) );
  AND2X1_HVT U866 ( .A1(conv_weight_box[43]), .A2(n411), .Y(
        DP_OP_423J2_125_3477_n2289) );
  INVX2_HVT U867 ( .A(DP_OP_425J2_127_3477_n2621), .Y(n411) );
  INVX2_HVT U868 ( .A(DP_OP_423J2_125_3477_n2225), .Y(n412) );
  INVX2_HVT U869 ( .A(DP_OP_425J2_127_3477_n2708), .Y(n413) );
  AND2X1_HVT U870 ( .A1(conv_weight_box[43]), .A2(n414), .Y(
        DP_OP_423J2_125_3477_n2293) );
  INVX2_HVT U871 ( .A(DP_OP_423J2_125_3477_n2317), .Y(n414) );
  INVX2_HVT U872 ( .A(DP_OP_423J2_125_3477_n2310), .Y(n415) );
  INVX2_HVT U873 ( .A(DP_OP_424J2_126_3477_n2311), .Y(n416) );
  INVX2_HVT U874 ( .A(DP_OP_425J2_127_3477_n2622), .Y(n417) );
  INVX2_HVT U875 ( .A(DP_OP_425J2_127_3477_n2620), .Y(n418) );
  INVX2_HVT U876 ( .A(DP_OP_423J2_125_3477_n2311), .Y(n419) );
  INVX2_HVT U877 ( .A(DP_OP_423J2_125_3477_n2228), .Y(n420) );
  INVX2_HVT U878 ( .A(DP_OP_423J2_125_3477_n2315), .Y(n421) );
  INVX2_HVT U879 ( .A(DP_OP_423J2_125_3477_n2316), .Y(n422) );
  NBUFFX2_HVT U880 ( .A(DP_OP_424J2_126_3477_n2582), .Y(n424) );
  NBUFFX2_HVT U881 ( .A(n1928), .Y(n425) );
  INVX2_HVT U882 ( .A(DP_OP_424J2_126_3477_n2582), .Y(conv_weight_box[61]) );
  MUX21X1_HVT U883 ( .A1(n427), .A2(n426), .S0(n423), .Y(
        DP_OP_424J2_126_3477_n2582) );
  INVX2_HVT U884 ( .A(conv1_sram_rdata_weight[91]), .Y(n426) );
  INVX2_HVT U885 ( .A(conv2_sram_rdata_weight[91]), .Y(n427) );
  AND2X1_HVT U886 ( .A1(n1484), .A2(n428), .Y(DP_OP_424J2_126_3477_n1935) );
  INVX2_HVT U887 ( .A(n1980), .Y(n428) );
  AND2X1_HVT U888 ( .A1(n1484), .A2(n429), .Y(DP_OP_423J2_125_3477_n1930) );
  INVX2_HVT U889 ( .A(n1281), .Y(n429) );
  AND2X1_HVT U890 ( .A1(n1484), .A2(n430), .Y(DP_OP_425J2_127_3477_n1927) );
  INVX2_HVT U891 ( .A(n1983), .Y(n430) );
  AND2X1_HVT U892 ( .A1(n1484), .A2(n431), .Y(DP_OP_425J2_127_3477_n1931) );
  INVX2_HVT U893 ( .A(n1280), .Y(n431) );
  AND2X1_HVT U894 ( .A1(n1484), .A2(n432), .Y(DP_OP_424J2_126_3477_n1925) );
  INVX2_HVT U895 ( .A(n1868), .Y(n432) );
  AND2X1_HVT U896 ( .A1(n1484), .A2(n433), .Y(DP_OP_422J2_124_3477_n1924) );
  INVX2_HVT U897 ( .A(n1879), .Y(n433) );
  AND2X1_HVT U898 ( .A1(n1484), .A2(n434), .Y(DP_OP_425J2_127_3477_n1924) );
  INVX2_HVT U899 ( .A(n1320), .Y(n434) );
  AND2X1_HVT U900 ( .A1(n1484), .A2(n435), .Y(DP_OP_425J2_127_3477_n324) );
  INVX2_HVT U901 ( .A(n1300), .Y(n435) );
  AND2X1_HVT U902 ( .A1(n1484), .A2(n436), .Y(DP_OP_423J2_125_3477_n318) );
  INVX2_HVT U903 ( .A(n1308), .Y(n436) );
  AND2X1_HVT U904 ( .A1(n1484), .A2(n437), .Y(DP_OP_424J2_126_3477_n316) );
  INVX2_HVT U905 ( .A(n1909), .Y(n437) );
  AND2X1_HVT U906 ( .A1(n1484), .A2(n438), .Y(DP_OP_425J2_127_3477_n1923) );
  INVX2_HVT U907 ( .A(n1302), .Y(n438) );
  AND2X1_HVT U908 ( .A1(n1484), .A2(n439), .Y(DP_OP_425J2_127_3477_n304) );
  INVX2_HVT U909 ( .A(n1330), .Y(n439) );
  OA21X1_HVT U910 ( .A1(DP_OP_422J2_124_3477_n251), .A2(
        DP_OP_422J2_124_3477_n253), .A3(DP_OP_422J2_124_3477_n252), .Y(n1577)
         );
  OR2X1_HVT U911 ( .A1(n440), .A2(n441), .Y(DP_OP_422J2_124_3477_n252) );
  AND2X1_HVT U912 ( .A1(n441), .A2(n440), .Y(DP_OP_422J2_124_3477_n251) );
  INVX2_HVT U913 ( .A(DP_OP_422J2_124_3477_n1215), .Y(n440) );
  XOR3X2_HVT U914 ( .A1(n889), .A2(DP_OP_422J2_124_3477_n1219), .A3(n442), .Y(
        n441) );
  INVX2_HVT U915 ( .A(DP_OP_422J2_124_3477_n1400), .Y(n442) );
  XOR3X2_HVT U916 ( .A1(DP_OP_422J2_124_3477_n1225), .A2(
        DP_OP_422J2_124_3477_n1406), .A3(DP_OP_422J2_124_3477_n1404), .Y(n889)
         );
  INVX2_HVT U917 ( .A(n443), .Y(n444) );
  INVX2_HVT U918 ( .A(DP_OP_422J2_124_3477_n2937), .Y(n443) );
  NBUFFX8_HVT U919 ( .A(DP_OP_422J2_124_3477_n2937), .Y(n445) );
  NBUFFX8_HVT U920 ( .A(n444), .Y(n446) );
  NAND2X0_HVT U921 ( .A1(n843), .A2(conv1_sram_rdata_weight[24]), .Y(n448) );
  AND2X4_HVT U922 ( .A1(n447), .A2(n685), .Y(DP_OP_424J2_126_3477_n2919) );
  INVX4_HVT U923 ( .A(n445), .Y(n447) );
  OA21X2_HVT U924 ( .A1(n843), .A2(n449), .A3(n448), .Y(
        DP_OP_422J2_124_3477_n2937) );
  INVX4_HVT U925 ( .A(conv2_sram_rdata_weight[24]), .Y(n449) );
  NBUFFX2_HVT U926 ( .A(n1484), .Y(n450) );
  NAND2X0_HVT U927 ( .A1(n1484), .A2(n451), .Y(n571) );
  INVX2_HVT U928 ( .A(n1987), .Y(n451) );
  AND2X4_HVT U929 ( .A1(n1484), .A2(n452), .Y(DP_OP_423J2_125_3477_n1928) );
  INVX4_HVT U930 ( .A(n1858), .Y(n452) );
  AND2X1_HVT U931 ( .A1(n450), .A2(n453), .Y(DP_OP_425J2_127_3477_n1925) );
  INVX2_HVT U932 ( .A(n1289), .Y(n453) );
  AND2X1_HVT U933 ( .A1(n450), .A2(n454), .Y(DP_OP_423J2_125_3477_n1924) );
  INVX2_HVT U934 ( .A(n1880), .Y(n454) );
  AND2X1_HVT U935 ( .A1(n450), .A2(n455), .Y(DP_OP_422J2_124_3477_n330) );
  INVX2_HVT U936 ( .A(n1318), .Y(n455) );
  AND2X1_HVT U937 ( .A1(n450), .A2(n456), .Y(DP_OP_423J2_125_3477_n322) );
  INVX2_HVT U938 ( .A(n1312), .Y(n456) );
  NAND2X0_HVT U939 ( .A1(n450), .A2(n457), .Y(n1380) );
  INVX2_HVT U940 ( .A(n1908), .Y(n457) );
  AND2X1_HVT U941 ( .A1(n450), .A2(n458), .Y(DP_OP_424J2_126_3477_n318) );
  INVX2_HVT U942 ( .A(n1894), .Y(n458) );
  AND2X1_HVT U943 ( .A1(n450), .A2(n459), .Y(DP_OP_423J2_125_3477_n308) );
  INVX2_HVT U944 ( .A(n1881), .Y(n459) );
  AND2X1_HVT U945 ( .A1(n450), .A2(n460), .Y(DP_OP_424J2_126_3477_n1923) );
  INVX2_HVT U946 ( .A(n1905), .Y(n460) );
  AND2X1_HVT U947 ( .A1(n450), .A2(n461), .Y(DP_OP_423J2_125_3477_n304) );
  INVX2_HVT U948 ( .A(n1329), .Y(n461) );
  NAND2X0_HVT U949 ( .A1(n450), .A2(n462), .Y(n1584) );
  INVX2_HVT U950 ( .A(n1323), .Y(n462) );
  INVX4_HVT U951 ( .A(n463), .Y(n464) );
  INVX2_HVT U952 ( .A(conv_weight_box[65]), .Y(n463) );
  NAND2X0_HVT U953 ( .A1(conv_weight_box[65]), .A2(n465), .Y(
        DP_OP_424J2_126_3477_n2459) );
  INVX2_HVT U954 ( .A(DP_OP_424J2_126_3477_n2491), .Y(n465) );
  NAND2X0_HVT U955 ( .A1(conv_weight_box[65]), .A2(n466), .Y(
        DP_OP_423J2_125_3477_n2458) );
  INVX2_HVT U956 ( .A(DP_OP_422J2_124_3477_n2578), .Y(n466) );
  NAND2X0_HVT U957 ( .A1(conv_weight_box[65]), .A2(n467), .Y(
        DP_OP_422J2_124_3477_n2459) );
  INVX2_HVT U958 ( .A(DP_OP_422J2_124_3477_n2491), .Y(n467) );
  NAND2X0_HVT U959 ( .A1(conv_weight_box[65]), .A2(n468), .Y(
        DP_OP_423J2_125_3477_n2459) );
  INVX2_HVT U960 ( .A(DP_OP_422J2_124_3477_n2579), .Y(n468) );
  NAND2X0_HVT U961 ( .A1(n464), .A2(n469), .Y(DP_OP_422J2_124_3477_n2460) );
  INVX2_HVT U962 ( .A(DP_OP_423J2_125_3477_n2536), .Y(n469) );
  NAND2X0_HVT U963 ( .A1(n464), .A2(n470), .Y(DP_OP_424J2_126_3477_n2460) );
  INVX2_HVT U964 ( .A(DP_OP_425J2_127_3477_n2536), .Y(n470) );
  NAND2X0_HVT U965 ( .A1(n464), .A2(n471), .Y(DP_OP_423J2_125_3477_n2457) );
  INVX2_HVT U966 ( .A(DP_OP_422J2_124_3477_n2577), .Y(n471) );
  NAND2X0_HVT U967 ( .A1(n464), .A2(n472), .Y(DP_OP_422J2_124_3477_n2455) );
  INVX2_HVT U968 ( .A(DP_OP_423J2_125_3477_n2531), .Y(n472) );
  NAND2X0_HVT U969 ( .A1(n464), .A2(n473), .Y(DP_OP_424J2_126_3477_n2456) );
  INVX2_HVT U970 ( .A(DP_OP_423J2_125_3477_n2400), .Y(n473) );
  NAND2X0_HVT U971 ( .A1(n464), .A2(n474), .Y(DP_OP_423J2_125_3477_n2461) );
  INVX2_HVT U972 ( .A(DP_OP_423J2_125_3477_n2493), .Y(n474) );
  NAND2X0_HVT U973 ( .A1(n464), .A2(n475), .Y(DP_OP_422J2_124_3477_n2456) );
  INVX2_HVT U974 ( .A(DP_OP_422J2_124_3477_n2488), .Y(n475) );
  NAND2X0_HVT U975 ( .A1(n464), .A2(n476), .Y(DP_OP_422J2_124_3477_n2461) );
  INVX2_HVT U976 ( .A(DP_OP_423J2_125_3477_n2537), .Y(n476) );
  AND2X4_HVT U977 ( .A1(n464), .A2(n477), .Y(DP_OP_423J2_125_3477_n2454) );
  INVX2_HVT U978 ( .A(DP_OP_422J2_124_3477_n2574), .Y(n477) );
  AND2X1_HVT U979 ( .A1(n1484), .A2(n478), .Y(DP_OP_422J2_124_3477_n1928) );
  INVX2_HVT U980 ( .A(n1285), .Y(n478) );
  AND2X1_HVT U981 ( .A1(n1484), .A2(n479), .Y(DP_OP_425J2_127_3477_n1934) );
  INVX2_HVT U982 ( .A(n1282), .Y(n479) );
  AND2X1_HVT U983 ( .A1(n1484), .A2(n480), .Y(DP_OP_422J2_124_3477_n1925) );
  INVX2_HVT U984 ( .A(n1864), .Y(n480) );
  AND2X1_HVT U985 ( .A1(n1484), .A2(n481), .Y(DP_OP_423J2_125_3477_n324) );
  INVX2_HVT U986 ( .A(n1303), .Y(n481) );
  AND2X1_HVT U987 ( .A1(n1484), .A2(n482), .Y(DP_OP_422J2_124_3477_n320) );
  INVX2_HVT U988 ( .A(n1901), .Y(n482) );
  NAND2X0_HVT U989 ( .A1(n1484), .A2(n483), .Y(n1382) );
  INVX2_HVT U990 ( .A(n1307), .Y(n483) );
  AND2X1_HVT U991 ( .A1(n1484), .A2(n484), .Y(DP_OP_425J2_127_3477_n308) );
  INVX2_HVT U992 ( .A(n1299), .Y(n484) );
  AND2X1_HVT U993 ( .A1(n1484), .A2(n485), .Y(DP_OP_423J2_125_3477_n1923) );
  INVX2_HVT U994 ( .A(n1301), .Y(n485) );
  NAND2X0_HVT U995 ( .A1(n1484), .A2(n486), .Y(n1669) );
  INVX2_HVT U996 ( .A(n1914), .Y(n486) );
  NAND2X0_HVT U997 ( .A1(n1484), .A2(n487), .Y(n1757) );
  INVX2_HVT U998 ( .A(n1324), .Y(n487) );
  NAND3X0_HVT U999 ( .A1(n1958), .A2(n2037), .A3(n1956), .Y(n1955) );
  INVX2_HVT U1000 ( .A(n2043), .Y(n489) );
  OA21X1_HVT U1001 ( .A1(n2040), .A2(n2020), .A3(n491), .Y(n2043) );
  INVX2_HVT U1002 ( .A(n1966), .Y(n1965) );
  NAND2X0_HVT U1003 ( .A1(n1958), .A2(n993), .Y(n1954) );
  NBUFFX2_HVT U1004 ( .A(n1965), .Y(n490) );
  AND2X1_HVT U1005 ( .A1(n488), .A2(conv2_sum_a[9]), .Y(n2173) );
  OA21X1_HVT U1006 ( .A1(n2022), .A2(n2021), .A3(n2019), .Y(n491) );
  NBUFFX2_HVT U1007 ( .A(conv_weight_box[65]), .Y(n492) );
  NAND2X0_HVT U1008 ( .A1(conv_weight_box[65]), .A2(n493), .Y(
        DP_OP_422J2_124_3477_n2458) );
  INVX2_HVT U1009 ( .A(DP_OP_422J2_124_3477_n2490), .Y(n493) );
  NAND2X0_HVT U1010 ( .A1(conv_weight_box[65]), .A2(n494), .Y(
        DP_OP_424J2_126_3477_n2458) );
  INVX2_HVT U1011 ( .A(DP_OP_425J2_127_3477_n2534), .Y(n494) );
  NAND2X0_HVT U1012 ( .A1(conv_weight_box[65]), .A2(n495), .Y(
        DP_OP_424J2_126_3477_n2457) );
  INVX2_HVT U1013 ( .A(DP_OP_423J2_125_3477_n2401), .Y(n495) );
  NAND2X0_HVT U1014 ( .A1(conv_weight_box[65]), .A2(n496), .Y(
        DP_OP_422J2_124_3477_n2457) );
  INVX2_HVT U1015 ( .A(DP_OP_422J2_124_3477_n2489), .Y(n496) );
  NAND2X0_HVT U1016 ( .A1(n492), .A2(n497), .Y(DP_OP_424J2_126_3477_n2461) );
  INVX2_HVT U1017 ( .A(DP_OP_423J2_125_3477_n2405), .Y(n497) );
  NAND2X0_HVT U1018 ( .A1(n492), .A2(n498), .Y(DP_OP_423J2_125_3477_n2460) );
  INVX2_HVT U1019 ( .A(DP_OP_422J2_124_3477_n2580), .Y(n498) );
  NAND2X0_HVT U1020 ( .A1(n492), .A2(n499), .Y(DP_OP_423J2_125_3477_n2455) );
  INVX2_HVT U1021 ( .A(DP_OP_422J2_124_3477_n2575), .Y(n499) );
  NAND2X0_HVT U1022 ( .A1(n492), .A2(n500), .Y(DP_OP_424J2_126_3477_n2455) );
  INVX2_HVT U1023 ( .A(DP_OP_422J2_124_3477_n2663), .Y(n500) );
  NAND2X0_HVT U1024 ( .A1(n492), .A2(n501), .Y(DP_OP_423J2_125_3477_n2456) );
  INVX2_HVT U1025 ( .A(DP_OP_422J2_124_3477_n2576), .Y(n501) );
  AND2X1_HVT U1026 ( .A1(n492), .A2(n502), .Y(DP_OP_422J2_124_3477_n2454) );
  INVX2_HVT U1027 ( .A(DP_OP_422J2_124_3477_n2486), .Y(n502) );
  AND2X4_HVT U1028 ( .A1(n492), .A2(n503), .Y(DP_OP_424J2_126_3477_n2454) );
  INVX2_HVT U1029 ( .A(DP_OP_424J2_126_3477_n2486), .Y(n503) );
  NBUFFX2_HVT U1030 ( .A(conv_weight_box[27]), .Y(n504) );
  AND2X1_HVT U1031 ( .A1(conv_weight_box[27]), .A2(n505), .Y(
        DP_OP_422J2_124_3477_n2825) );
  INVX2_HVT U1032 ( .A(DP_OP_422J2_124_3477_n2841), .Y(n505) );
  AND2X1_HVT U1033 ( .A1(conv_weight_box[27]), .A2(n506), .Y(
        DP_OP_422J2_124_3477_n2824) );
  INVX2_HVT U1034 ( .A(DP_OP_422J2_124_3477_n2840), .Y(n506) );
  AND2X1_HVT U1035 ( .A1(n504), .A2(n507), .Y(DP_OP_422J2_124_3477_n2828) );
  INVX2_HVT U1036 ( .A(DP_OP_425J2_127_3477_n2712), .Y(n507) );
  AND2X1_HVT U1037 ( .A1(n504), .A2(n508), .Y(DP_OP_423J2_125_3477_n2825) );
  INVX2_HVT U1038 ( .A(DP_OP_423J2_125_3477_n2841), .Y(n508) );
  NAND2X0_HVT U1039 ( .A1(n504), .A2(n509), .Y(DP_OP_422J2_124_3477_n2822) );
  INVX2_HVT U1040 ( .A(DP_OP_422J2_124_3477_n2838), .Y(n509) );
  AND2X1_HVT U1041 ( .A1(n504), .A2(n510), .Y(DP_OP_422J2_124_3477_n2829) );
  INVX2_HVT U1042 ( .A(DP_OP_423J2_125_3477_n2229), .Y(n510) );
  AND2X1_HVT U1043 ( .A1(n504), .A2(n511), .Y(DP_OP_422J2_124_3477_n2826) );
  INVX2_HVT U1044 ( .A(DP_OP_422J2_124_3477_n2842), .Y(n511) );
  AND2X1_HVT U1045 ( .A1(n504), .A2(n512), .Y(DP_OP_423J2_125_3477_n2826) );
  INVX2_HVT U1046 ( .A(DP_OP_423J2_125_3477_n2842), .Y(n512) );
  AND2X1_HVT U1047 ( .A1(n504), .A2(n513), .Y(DP_OP_423J2_125_3477_n2827) );
  INVX2_HVT U1048 ( .A(DP_OP_423J2_125_3477_n2843), .Y(n513) );
  AND2X1_HVT U1049 ( .A1(n504), .A2(n514), .Y(DP_OP_422J2_124_3477_n2823) );
  INVX2_HVT U1050 ( .A(DP_OP_422J2_124_3477_n2839), .Y(n514) );
  AND2X4_HVT U1051 ( .A1(n504), .A2(n515), .Y(DP_OP_422J2_124_3477_n2827) );
  INVX2_HVT U1052 ( .A(DP_OP_423J2_125_3477_n2227), .Y(n515) );
  NAND2X0_HVT U1053 ( .A1(n517), .A2(n516), .Y(DP_OP_423J2_125_3477_n340) );
  NAND2X0_HVT U1054 ( .A1(DP_OP_423J2_125_3477_n343), .A2(
        DP_OP_423J2_125_3477_n354), .Y(n516) );
  NAND2X0_HVT U1055 ( .A1(DP_OP_423J2_125_3477_n352), .A2(n518), .Y(n517) );
  OR2X1_HVT U1056 ( .A1(DP_OP_423J2_125_3477_n354), .A2(
        DP_OP_423J2_125_3477_n343), .Y(n518) );
  XOR3X2_HVT U1057 ( .A1(DP_OP_423J2_125_3477_n343), .A2(
        DP_OP_423J2_125_3477_n354), .A3(DP_OP_423J2_125_3477_n352), .Y(
        DP_OP_423J2_125_3477_n341) );
  NAND3X0_HVT U1058 ( .A1(n527), .A2(n522), .A3(n519), .Y(n_conv2_sum_c[22])
         );
  NAND2X0_HVT U1059 ( .A1(n182), .A2(n520), .Y(n519) );
  INVX2_HVT U1060 ( .A(n521), .Y(n520) );
  NAND2X0_HVT U1061 ( .A1(DP_OP_424J2_126_3477_n131), .A2(
        DP_OP_424J2_126_3477_n15), .Y(n521) );
  NAND2X0_HVT U1062 ( .A1(n524), .A2(n523), .Y(n522) );
  NAND2X0_HVT U1063 ( .A1(DP_OP_424J2_126_3477_n132), .A2(n526), .Y(n523) );
  AO21X1_HVT U1064 ( .A1(n526), .A2(n525), .A3(DP_OP_424J2_126_3477_n132), .Y(
        n524) );
  INVX2_HVT U1065 ( .A(DP_OP_424J2_126_3477_n131), .Y(n525) );
  INVX2_HVT U1066 ( .A(DP_OP_424J2_126_3477_n15), .Y(n526) );
  OR3X1_HVT U1067 ( .A1(DP_OP_424J2_126_3477_n15), .A2(n242), .A3(
        DP_OP_424J2_126_3477_n132), .Y(n527) );
  AO22X1_HVT U1068 ( .A1(n531), .A2(n530), .A3(n529), .A4(n528), .Y(n536) );
  OR2X1_HVT U1069 ( .A1(n1981), .A2(conv2_sum_a[3]), .Y(n528) );
  AND2X1_HVT U1070 ( .A1(conv2_sum_a[2]), .A2(n1866), .Y(n529) );
  INVX2_HVT U1071 ( .A(n1872), .Y(n530) );
  INVX2_HVT U1072 ( .A(conv2_sum_b[3]), .Y(n531) );
  NAND3X0_HVT U1073 ( .A1(n534), .A2(n2038), .A3(n532), .Y(n1957) );
  NAND3X0_HVT U1074 ( .A1(n535), .A2(n533), .A3(n539), .Y(n532) );
  AND2X1_HVT U1075 ( .A1(n538), .A2(n537), .Y(n533) );
  NAND2X0_HVT U1076 ( .A1(n536), .A2(n535), .Y(n534) );
  INVX2_HVT U1077 ( .A(n2034), .Y(n535) );
  NAND2X0_HVT U1078 ( .A1(conv2_sum_b[3]), .A2(n1872), .Y(n537) );
  NAND3X0_HVT U1079 ( .A1(n996), .A2(n1869), .A3(conv2_sum_b[0]), .Y(n538) );
  OA21X1_HVT U1080 ( .A1(n1989), .A2(conv2_sum_a[1]), .A3(n540), .Y(n539) );
  NAND2X0_HVT U1081 ( .A1(conv2_sum_b[2]), .A2(n1867), .Y(n540) );
  INVX2_HVT U1082 ( .A(conv_weight_box[37]), .Y(DP_OP_423J2_125_3477_n2276) );
  FADDX1_HVT U1083 ( .A(n1191), .B(DP_OP_423J2_125_3477_n970), .CI(
        DP_OP_423J2_125_3477_n968), .CO(DP_OP_423J2_125_3477_n748) );
  AO22X1_HVT U1084 ( .A1(DP_OP_423J2_125_3477_n2816), .A2(
        DP_OP_423J2_125_3477_n2251), .A3(DP_OP_423J2_125_3477_n2244), .A4(n541), .Y(n1191) );
  NAND2X0_HVT U1085 ( .A1(n543), .A2(n542), .Y(n541) );
  INVX2_HVT U1086 ( .A(DP_OP_423J2_125_3477_n2816), .Y(n542) );
  INVX2_HVT U1087 ( .A(DP_OP_423J2_125_3477_n2251), .Y(n543) );
  AND2X1_HVT U1088 ( .A1(conv_weight_box[37]), .A2(n544), .Y(
        DP_OP_423J2_125_3477_n2251) );
  INVX2_HVT U1089 ( .A(DP_OP_423J2_125_3477_n2267), .Y(n544) );
  INVX2_HVT U1090 ( .A(n545), .Y(DP_OP_425J2_127_3477_n259) );
  OR2X1_HVT U1091 ( .A1(DP_OP_425J2_127_3477_n1579), .A2(
        DP_OP_425J2_127_3477_n1577), .Y(n545) );
  XOR3X2_HVT U1092 ( .A1(DP_OP_425J2_127_3477_n1583), .A2(
        DP_OP_425J2_127_3477_n1730), .A3(DP_OP_425J2_127_3477_n1581), .Y(
        DP_OP_425J2_127_3477_n1577) );
  NBUFFX2_HVT U1093 ( .A(n585), .Y(n546) );
  NAND2X0_HVT U1094 ( .A1(n585), .A2(n547), .Y(DP_OP_423J2_125_3477_n2105) );
  INVX2_HVT U1095 ( .A(DP_OP_425J2_127_3477_n2797), .Y(n547) );
  NAND2X0_HVT U1096 ( .A1(n36), .A2(n548), .Y(DP_OP_423J2_125_3477_n2106) );
  INVX2_HVT U1097 ( .A(DP_OP_425J2_127_3477_n2798), .Y(n548) );
  NAND2X0_HVT U1098 ( .A1(n546), .A2(n549), .Y(DP_OP_423J2_125_3477_n2109) );
  INVX2_HVT U1099 ( .A(DP_OP_425J2_127_3477_n2801), .Y(n549) );
  NAND2X0_HVT U1100 ( .A1(n546), .A2(n550), .Y(DP_OP_423J2_125_3477_n2108) );
  INVX2_HVT U1101 ( .A(DP_OP_423J2_125_3477_n2140), .Y(n550) );
  NAND2X0_HVT U1102 ( .A1(n546), .A2(n551), .Y(DP_OP_423J2_125_3477_n2107) );
  INVX2_HVT U1103 ( .A(DP_OP_425J2_127_3477_n2799), .Y(n551) );
  NAND2X0_HVT U1104 ( .A1(n546), .A2(n552), .Y(DP_OP_423J2_125_3477_n2104) );
  INVX2_HVT U1105 ( .A(DP_OP_425J2_127_3477_n2796), .Y(n552) );
  AND2X1_HVT U1106 ( .A1(n546), .A2(n553), .Y(DP_OP_423J2_125_3477_n2102) );
  INVX2_HVT U1107 ( .A(DP_OP_422J2_124_3477_n2926), .Y(n553) );
  NAND2X0_HVT U1108 ( .A1(n546), .A2(n554), .Y(DP_OP_423J2_125_3477_n2103) );
  INVX2_HVT U1109 ( .A(DP_OP_423J2_125_3477_n2135), .Y(n554) );
  AND2X4_HVT U1110 ( .A1(n546), .A2(n555), .Y(DP_OP_425J2_127_3477_n2102) );
  INVX2_HVT U1111 ( .A(DP_OP_423J2_125_3477_n3014), .Y(n555) );
  NBUFFX2_HVT U1112 ( .A(DP_OP_423J2_125_3477_n2012), .Y(n556) );
  NBUFFX8_HVT U1113 ( .A(DP_OP_423J2_125_3477_n2012), .Y(n557) );
  NBUFFX16_HVT U1114 ( .A(DP_OP_423J2_125_3477_n2012), .Y(n558) );
  OA21X2_HVT U1115 ( .A1(n843), .A2(n560), .A3(n559), .Y(
        DP_OP_423J2_125_3477_n2012) );
  NAND2X0_HVT U1116 ( .A1(n843), .A2(conv1_sram_rdata_weight[5]), .Y(n559) );
  INVX2_HVT U1117 ( .A(conv2_sram_rdata_weight[5]), .Y(n560) );
  AND2X1_HVT U1118 ( .A1(n1387), .A2(n561), .Y(DP_OP_424J2_126_3477_n2342) );
  INVX2_HVT U1119 ( .A(DP_OP_424J2_126_3477_n2358), .Y(n561) );
  NAND2X0_HVT U1120 ( .A1(n1387), .A2(n562), .Y(DP_OP_422J2_124_3477_n2338) );
  INVX2_HVT U1121 ( .A(DP_OP_422J2_124_3477_n2354), .Y(n562) );
  AND2X1_HVT U1122 ( .A1(n1387), .A2(n563), .Y(DP_OP_425J2_127_3477_n2342) );
  INVX2_HVT U1123 ( .A(DP_OP_425J2_127_3477_n2358), .Y(n563) );
  AND2X1_HVT U1124 ( .A1(n1387), .A2(n564), .Y(DP_OP_423J2_125_3477_n2344) );
  INVX2_HVT U1125 ( .A(DP_OP_422J2_124_3477_n2712), .Y(n564) );
  AND2X1_HVT U1126 ( .A1(n1387), .A2(n565), .Y(DP_OP_422J2_124_3477_n2342) );
  INVX2_HVT U1127 ( .A(DP_OP_422J2_124_3477_n2358), .Y(n565) );
  AND2X1_HVT U1128 ( .A1(n1387), .A2(n566), .Y(DP_OP_425J2_127_3477_n2340) );
  INVX2_HVT U1129 ( .A(DP_OP_425J2_127_3477_n2356), .Y(n566) );
  AND2X1_HVT U1130 ( .A1(n1387), .A2(n567), .Y(DP_OP_423J2_125_3477_n2343) );
  INVX2_HVT U1131 ( .A(DP_OP_424J2_126_3477_n2447), .Y(n567) );
  AND2X1_HVT U1132 ( .A1(n1387), .A2(n568), .Y(DP_OP_423J2_125_3477_n2345) );
  INVX2_HVT U1133 ( .A(DP_OP_423J2_125_3477_n2361), .Y(n568) );
  FADDX1_HVT U1134 ( .A(DP_OP_425J2_127_3477_n2505), .B(n569), .CI(
        DP_OP_425J2_127_3477_n1977), .CO(DP_OP_425J2_127_3477_n1726) );
  INVX2_HVT U1135 ( .A(n571), .Y(n569) );
  INVX2_HVT U1136 ( .A(DP_OP_425J2_127_3477_n1977), .Y(n570) );
  NBUFFX2_HVT U1137 ( .A(conv_weight_box[27]), .Y(n572) );
  AND2X1_HVT U1138 ( .A1(n572), .A2(n573), .Y(DP_OP_424J2_126_3477_n2826) );
  INVX2_HVT U1139 ( .A(DP_OP_425J2_127_3477_n2226), .Y(n573) );
  NAND2X0_HVT U1140 ( .A1(n572), .A2(n574), .Y(DP_OP_424J2_126_3477_n2822) );
  INVX2_HVT U1141 ( .A(DP_OP_422J2_124_3477_n2090), .Y(n574) );
  AND2X1_HVT U1142 ( .A1(n572), .A2(n575), .Y(DP_OP_424J2_126_3477_n2828) );
  INVX2_HVT U1143 ( .A(DP_OP_423J2_125_3477_n2932), .Y(n575) );
  AND2X1_HVT U1144 ( .A1(conv_weight_box[27]), .A2(n576), .Y(
        DP_OP_424J2_126_3477_n2825) );
  INVX2_HVT U1145 ( .A(DP_OP_422J2_124_3477_n2093), .Y(n576) );
  AND2X1_HVT U1146 ( .A1(n572), .A2(n577), .Y(DP_OP_423J2_125_3477_n2823) );
  INVX2_HVT U1147 ( .A(DP_OP_425J2_127_3477_n2311), .Y(n577) );
  AND2X1_HVT U1148 ( .A1(conv_weight_box[27]), .A2(n578), .Y(
        DP_OP_423J2_125_3477_n2824) );
  INVX2_HVT U1149 ( .A(DP_OP_425J2_127_3477_n2312), .Y(n578) );
  AND2X1_HVT U1150 ( .A1(n572), .A2(n579), .Y(DP_OP_424J2_126_3477_n2829) );
  INVX2_HVT U1151 ( .A(DP_OP_424J2_126_3477_n2845), .Y(n579) );
  AND2X1_HVT U1152 ( .A1(n572), .A2(n580), .Y(DP_OP_424J2_126_3477_n2824) );
  INVX2_HVT U1153 ( .A(DP_OP_422J2_124_3477_n2092), .Y(n580) );
  AND2X1_HVT U1154 ( .A1(n572), .A2(n581), .Y(DP_OP_424J2_126_3477_n2827) );
  INVX2_HVT U1155 ( .A(DP_OP_423J2_125_3477_n2931), .Y(n581) );
  AND2X1_HVT U1156 ( .A1(n572), .A2(n582), .Y(DP_OP_424J2_126_3477_n2823) );
  INVX2_HVT U1157 ( .A(DP_OP_422J2_124_3477_n2091), .Y(n582) );
  NAND2X0_HVT U1158 ( .A1(n572), .A2(n583), .Y(DP_OP_423J2_125_3477_n2822) );
  INVX2_HVT U1159 ( .A(DP_OP_425J2_127_3477_n2310), .Y(n583) );
  AND2X4_HVT U1160 ( .A1(n572), .A2(n584), .Y(DP_OP_423J2_125_3477_n2829) );
  INVX2_HVT U1161 ( .A(DP_OP_423J2_125_3477_n2845), .Y(n584) );
  INVX2_HVT U1162 ( .A(DP_OP_422J2_124_3477_n3019), .Y(n586) );
  NAND2X0_HVT U1163 ( .A1(n36), .A2(n587), .Y(DP_OP_424J2_126_3477_n2108) );
  INVX2_HVT U1164 ( .A(DP_OP_423J2_125_3477_n2052), .Y(n587) );
  NAND2X0_HVT U1165 ( .A1(n37), .A2(n588), .Y(DP_OP_424J2_126_3477_n2109) );
  INVX2_HVT U1166 ( .A(DP_OP_422J2_124_3477_n3021), .Y(n588) );
  NAND2X0_HVT U1167 ( .A1(n36), .A2(n589), .Y(DP_OP_424J2_126_3477_n2104) );
  INVX2_HVT U1168 ( .A(DP_OP_424J2_126_3477_n2136), .Y(n589) );
  NAND2X0_HVT U1169 ( .A1(n37), .A2(n590), .Y(DP_OP_424J2_126_3477_n2105) );
  INVX2_HVT U1170 ( .A(DP_OP_425J2_127_3477_n2885), .Y(n590) );
  NAND2X0_HVT U1171 ( .A1(n37), .A2(n591), .Y(DP_OP_424J2_126_3477_n2106) );
  INVX2_HVT U1172 ( .A(DP_OP_424J2_126_3477_n2138), .Y(n591) );
  NAND2X0_HVT U1173 ( .A1(n37), .A2(n592), .Y(DP_OP_425J2_127_3477_n2108) );
  INVX2_HVT U1174 ( .A(DP_OP_424J2_126_3477_n2932), .Y(n592) );
  NAND2X0_HVT U1175 ( .A1(n37), .A2(n593), .Y(DP_OP_425J2_127_3477_n2104) );
  INVX2_HVT U1176 ( .A(DP_OP_424J2_126_3477_n2928), .Y(n593) );
  NAND2X0_HVT U1177 ( .A1(n37), .A2(n594), .Y(DP_OP_424J2_126_3477_n2103) );
  INVX2_HVT U1178 ( .A(DP_OP_422J2_124_3477_n3015), .Y(n594) );
  AND2X4_HVT U1179 ( .A1(n37), .A2(n595), .Y(DP_OP_424J2_126_3477_n2102) );
  INVX2_HVT U1180 ( .A(DP_OP_425J2_127_3477_n2882), .Y(n595) );
  NBUFFX8_HVT U1181 ( .A(DP_OP_422J2_124_3477_n2717), .Y(n596) );
  NBUFFX16_HVT U1182 ( .A(DP_OP_422J2_124_3477_n2717), .Y(n597) );
  OA21X2_HVT U1183 ( .A1(n843), .A2(n599), .A3(n598), .Y(
        DP_OP_422J2_124_3477_n2717) );
  NAND2X0_HVT U1184 ( .A1(n843), .A2(conv1_sram_rdata_weight[64]), .Y(n598) );
  INVX2_HVT U1185 ( .A(conv2_sram_rdata_weight[64]), .Y(n599) );
  NBUFFX2_HVT U1186 ( .A(n35), .Y(n600) );
  NBUFFX2_HVT U1187 ( .A(n35), .Y(n602) );
  NBUFFX2_HVT U1188 ( .A(n35), .Y(n603) );
  NBUFFX2_HVT U1189 ( .A(n601), .Y(n604) );
  AND2X4_HVT U1190 ( .A1(n605), .A2(src_window[104]), .Y(n1641) );
  AND2X1_HVT U1191 ( .A1(n605), .A2(src_window[112]), .Y(n1546) );
  INVX4_HVT U1192 ( .A(n601), .Y(n605) );
  INVX4_HVT U1193 ( .A(conv2_sram_rdata_weight[27]), .Y(n606) );
  NBUFFX2_HVT U1194 ( .A(conv_weight_box[39]), .Y(n607) );
  AND2X1_HVT U1195 ( .A1(conv_weight_box[39]), .A2(n608), .Y(
        DP_OP_424J2_126_3477_n2740) );
  INVX2_HVT U1196 ( .A(DP_OP_424J2_126_3477_n2756), .Y(n608) );
  AND2X1_HVT U1197 ( .A1(n607), .A2(n609), .Y(DP_OP_422J2_124_3477_n2737) );
  INVX2_HVT U1198 ( .A(DP_OP_422J2_124_3477_n2753), .Y(n609) );
  AND2X1_HVT U1199 ( .A1(n607), .A2(n610), .Y(DP_OP_422J2_124_3477_n2735) );
  INVX2_HVT U1200 ( .A(DP_OP_422J2_124_3477_n2751), .Y(n610) );
  AND2X1_HVT U1201 ( .A1(n607), .A2(n611), .Y(DP_OP_422J2_124_3477_n2740) );
  INVX2_HVT U1202 ( .A(DP_OP_422J2_124_3477_n2756), .Y(n611) );
  AND2X1_HVT U1203 ( .A1(n607), .A2(n612), .Y(DP_OP_424J2_126_3477_n2738) );
  INVX2_HVT U1204 ( .A(DP_OP_424J2_126_3477_n2754), .Y(n612) );
  AND2X1_HVT U1205 ( .A1(n607), .A2(n613), .Y(DP_OP_422J2_124_3477_n2736) );
  INVX2_HVT U1206 ( .A(DP_OP_424J2_126_3477_n2400), .Y(n613) );
  NAND2X0_HVT U1207 ( .A1(n607), .A2(n614), .Y(DP_OP_422J2_124_3477_n2734) );
  INVX2_HVT U1208 ( .A(DP_OP_422J2_124_3477_n2750), .Y(n614) );
  AND2X1_HVT U1209 ( .A1(n607), .A2(n615), .Y(DP_OP_422J2_124_3477_n2739) );
  INVX2_HVT U1210 ( .A(DP_OP_424J2_126_3477_n2403), .Y(n615) );
  AND2X1_HVT U1211 ( .A1(n607), .A2(n616), .Y(DP_OP_422J2_124_3477_n2741) );
  INVX2_HVT U1212 ( .A(DP_OP_424J2_126_3477_n2405), .Y(n616) );
  AND2X4_HVT U1213 ( .A1(n607), .A2(n617), .Y(DP_OP_422J2_124_3477_n2738) );
  INVX2_HVT U1214 ( .A(DP_OP_422J2_124_3477_n2754), .Y(n617) );
  INVX4_HVT U1215 ( .A(n618), .Y(n619) );
  INVX2_HVT U1216 ( .A(n423), .Y(n618) );
  NAND2X0_HVT U1217 ( .A1(n711), .A2(conv1_sram_rdata_weight[20]), .Y(n623) );
  AND2X4_HVT U1218 ( .A1(n622), .A2(src_window[98]), .Y(
        DP_OP_423J2_125_3477_n2087) );
  OA21X2_HVT U1219 ( .A1(n711), .A2(n624), .A3(n623), .Y(
        DP_OP_423J2_125_3477_n2101) );
  INVX4_HVT U1220 ( .A(conv2_sram_rdata_weight[20]), .Y(n624) );
  NAND2X0_HVT U1221 ( .A1(n626), .A2(n625), .Y(n1032) );
  NAND2X0_HVT U1222 ( .A1(DP_OP_424J2_126_3477_n284), .A2(
        DP_OP_424J2_126_3477_n174), .Y(n625) );
  OR2X1_HVT U1223 ( .A1(n627), .A2(n628), .Y(n1065) );
  NAND2X0_HVT U1224 ( .A1(n628), .A2(n627), .Y(n1064) );
  NAND2X0_HVT U1225 ( .A1(DP_OP_424J2_126_3477_n280), .A2(
        DP_OP_424J2_126_3477_n136), .Y(n627) );
  NAND2X0_HVT U1226 ( .A1(n629), .A2(DP_OP_424J2_126_3477_n141), .Y(n628) );
  NAND2X0_HVT U1227 ( .A1(n1518), .A2(DP_OP_424J2_126_3477_n138), .Y(n629) );
  NAND3X0_HVT U1228 ( .A1(n635), .A2(n633), .A3(n630), .Y(n_conv2_sum_c[18])
         );
  AO22X1_HVT U1229 ( .A1(n632), .A2(n1767), .A3(n637), .A4(n631), .Y(n630) );
  INVX2_HVT U1230 ( .A(n1767), .Y(n631) );
  NAND2X0_HVT U1231 ( .A1(n1760), .A2(n1477), .Y(n632) );
  NAND2X0_HVT U1232 ( .A1(n1722), .A2(n634), .Y(n633) );
  AND2X1_HVT U1233 ( .A1(n1767), .A2(n1477), .Y(n634) );
  OR2X1_HVT U1234 ( .A1(n636), .A2(n1722), .Y(n635) );
  OR2X1_HVT U1235 ( .A1(n637), .A2(n1760), .Y(n636) );
  INVX2_HVT U1236 ( .A(DP_OP_424J2_126_3477_n19), .Y(n637) );
  OA21X1_HVT U1237 ( .A1(n2033), .A2(n642), .A3(n638), .Y(n2029) );
  OA22X1_HVT U1238 ( .A1(conv2_sum_b[11]), .A2(n1973), .A3(n640), .A4(n639), 
        .Y(n638) );
  INVX2_HVT U1239 ( .A(n2025), .Y(n639) );
  NAND2X0_HVT U1240 ( .A1(n641), .A2(conv2_sum_a[10]), .Y(n640) );
  INVX2_HVT U1241 ( .A(conv2_sum_b[10]), .Y(n641) );
  AND2X1_HVT U1242 ( .A1(n644), .A2(n643), .Y(n642) );
  OR2X1_HVT U1243 ( .A1(n1874), .A2(conv2_sum_b[9]), .Y(n643) );
  NAND3X0_HVT U1244 ( .A1(n2031), .A2(conv2_sum_a[8]), .A3(n645), .Y(n644) );
  INVX2_HVT U1245 ( .A(conv2_sum_b[8]), .Y(n645) );
  AO21X1_HVT U1246 ( .A1(n650), .A2(n646), .A3(n2086), .Y(n2095) );
  OA22X1_HVT U1247 ( .A1(n1988), .A2(conv2_sum_d[3]), .A3(n648), .A4(n647), 
        .Y(n646) );
  AND2X1_HVT U1248 ( .A1(conv2_sum_d[3]), .A2(n1988), .Y(n647) );
  NAND2X0_HVT U1249 ( .A1(n649), .A2(conv2_sum_c[2]), .Y(n648) );
  INVX2_HVT U1250 ( .A(conv2_sum_d[2]), .Y(n649) );
  NAND3X0_HVT U1251 ( .A1(n655), .A2(n654), .A3(n651), .Y(n650) );
  NAND3X0_HVT U1252 ( .A1(n653), .A2(conv2_sum_d[0]), .A3(n652), .Y(n651) );
  INVX2_HVT U1253 ( .A(conv2_sum_c[0]), .Y(n652) );
  OR2X1_HVT U1254 ( .A1(n1980), .A2(conv2_sum_d[1]), .Y(n653) );
  OR2X1_HVT U1255 ( .A1(conv2_sum_c[1]), .A2(DP_OP_425J2_127_3477_n1968), .Y(
        n654) );
  INVX2_HVT U1256 ( .A(n2087), .Y(n655) );
  INVX2_HVT U1257 ( .A(mode[1]), .Y(n951) );
  INVX0_HVT U1258 ( .A(tmp_big1[17]), .Y(n656) );
  AO22X1_HVT U1259 ( .A1(n659), .A2(tmp_big1[17]), .A3(n2142), .A4(n657), .Y(
        n1946) );
  AND2X1_HVT U1260 ( .A1(tmp_big1[16]), .A2(n658), .Y(n657) );
  INVX2_HVT U1261 ( .A(tmp_big2[16]), .Y(n658) );
  NAND2X0_HVT U1262 ( .A1(tmp_big2[17]), .A2(n656), .Y(n2142) );
  INVX2_HVT U1263 ( .A(tmp_big2[17]), .Y(n659) );
  NAND2X0_HVT U1264 ( .A1(n661), .A2(n660), .Y(tmp_big2[17]) );
  NAND2X0_HVT U1265 ( .A1(n1532), .A2(conv2_sum_c[17]), .Y(n660) );
  NAND2X0_HVT U1266 ( .A1(n662), .A2(conv2_sum_d[17]), .Y(n661) );
  INVX2_HVT U1267 ( .A(n1532), .Y(n662) );
  NBUFFX2_HVT U1268 ( .A(n254), .Y(n663) );
  NAND2X1_HVT U1269 ( .A1(n664), .A2(src_window[80]), .Y(
        DP_OP_423J2_125_3477_n2945) );
  INVX4_HVT U1270 ( .A(n254), .Y(n664) );
  INVX4_HVT U1271 ( .A(conv2_sram_rdata_weight[19]), .Y(n665) );
  AO22X1_HVT U1272 ( .A1(DP_OP_424J2_126_3477_n3026), .A2(
        DP_OP_424J2_126_3477_n1970), .A3(n667), .A4(n666), .Y(
        DP_OP_424J2_126_3477_n508) );
  OR2X1_HVT U1273 ( .A1(DP_OP_424J2_126_3477_n3026), .A2(
        DP_OP_424J2_126_3477_n1970), .Y(n666) );
  XOR3X2_HVT U1274 ( .A1(DP_OP_424J2_126_3477_n1970), .A2(
        DP_OP_424J2_126_3477_n3026), .A3(n667), .Y(DP_OP_424J2_126_3477_n509)
         );
  INVX2_HVT U1275 ( .A(DP_OP_424J2_126_3477_n510), .Y(n667) );
  AO22X1_HVT U1276 ( .A1(DP_OP_422J2_124_3477_n1219), .A2(n889), .A3(n668), 
        .A4(DP_OP_422J2_124_3477_n1400), .Y(DP_OP_422J2_124_3477_n1212) );
  OR2X1_HVT U1277 ( .A1(DP_OP_422J2_124_3477_n1219), .A2(
        DP_OP_422J2_124_3477_n1217), .Y(n668) );
  INVX2_HVT U1278 ( .A(DP_OP_424J2_126_3477_n2752), .Y(n669) );
  NBUFFX8_HVT U1279 ( .A(DP_OP_422J2_124_3477_n2583), .Y(n670) );
  NBUFFX16_HVT U1280 ( .A(DP_OP_422J2_124_3477_n2583), .Y(n671) );
  OA21X2_HVT U1281 ( .A1(n711), .A2(n673), .A3(n672), .Y(
        DP_OP_422J2_124_3477_n2583) );
  NAND2X0_HVT U1282 ( .A1(n711), .A2(conv1_sram_rdata_weight[90]), .Y(n672) );
  INVX2_HVT U1283 ( .A(conv2_sram_rdata_weight[90]), .Y(n673) );
  NBUFFX2_HVT U1284 ( .A(n677), .Y(n674) );
  NBUFFX2_HVT U1285 ( .A(DP_OP_425J2_127_3477_n2981), .Y(n675) );
  NBUFFX8_HVT U1286 ( .A(DP_OP_425J2_127_3477_n2981), .Y(n676) );
  NBUFFX16_HVT U1287 ( .A(DP_OP_425J2_127_3477_n2981), .Y(n677) );
  OA21X2_HVT U1288 ( .A1(n711), .A2(n679), .A3(n678), .Y(
        DP_OP_425J2_127_3477_n2981) );
  NAND2X0_HVT U1289 ( .A1(n711), .A2(conv1_sram_rdata_weight[16]), .Y(n678) );
  INVX2_HVT U1290 ( .A(conv2_sram_rdata_weight[16]), .Y(n679) );
  INVX1_HVT U1291 ( .A(n680), .Y(n726) );
  AND2X4_HVT U1292 ( .A1(n726), .A2(n728), .Y(DP_OP_424J2_126_3477_n2733) );
  AND2X1_HVT U1293 ( .A1(n682), .A2(n681), .Y(n680) );
  NAND2X0_HVT U1294 ( .A1(n713), .A2(conv2_sram_rdata_weight[58]), .Y(n681) );
  NAND2X0_HVT U1295 ( .A1(n711), .A2(conv1_sram_rdata_weight[58]), .Y(n682) );
  INVX2_HVT U1296 ( .A(conv_weight_box[10]), .Y(DP_OP_424J2_126_3477_n2055) );
  NAND3X0_HVT U1297 ( .A1(n935), .A2(n936), .A3(n683), .Y(
        DP_OP_424J2_126_3477_n1180) );
  NAND2X0_HVT U1298 ( .A1(DP_OP_424J2_126_3477_n2919), .A2(
        DP_OP_424J2_126_3477_n2025), .Y(n683) );
  AND2X1_HVT U1299 ( .A1(conv_weight_box[10]), .A2(n684), .Y(
        DP_OP_424J2_126_3477_n2025) );
  INVX2_HVT U1300 ( .A(DP_OP_425J2_127_3477_n2973), .Y(n684) );
  INVX2_HVT U1301 ( .A(DP_OP_424J2_126_3477_n2927), .Y(n685) );
  AND2X2_HVT U1302 ( .A1(n1928), .A2(n688), .Y(n686) );
  INVX4_HVT U1303 ( .A(n1928), .Y(n687) );
  INVX2_HVT U1304 ( .A(conv2_sram_rdata_weight[71]), .Y(n688) );
  INVX2_HVT U1305 ( .A(conv1_sram_rdata_weight[71]), .Y(n689) );
  NBUFFX2_HVT U1306 ( .A(n34), .Y(n690) );
  NBUFFX2_HVT U1307 ( .A(n34), .Y(n691) );
  NBUFFX2_HVT U1308 ( .A(n34), .Y(n692) );
  NBUFFX2_HVT U1309 ( .A(n694), .Y(n693) );
  NAND2X0_HVT U1310 ( .A1(n843), .A2(conv1_sram_rdata_weight[0]), .Y(n696) );
  AND2X4_HVT U1311 ( .A1(n695), .A2(src_window[48]), .Y(
        DP_OP_423J2_125_3477_n3055) );
  INVX4_HVT U1312 ( .A(n34), .Y(n695) );
  INVX4_HVT U1313 ( .A(conv2_sram_rdata_weight[0]), .Y(n697) );
  NBUFFX2_HVT U1314 ( .A(n704), .Y(n698) );
  NBUFFX2_HVT U1315 ( .A(n704), .Y(n699) );
  INVX2_HVT U1316 ( .A(n7001), .Y(n1648) );
  INVX2_HVT U1317 ( .A(n701), .Y(n703) );
  INVX0_HVT U1318 ( .A(n702), .Y(n705) );
  INVX2_HVT U1319 ( .A(DP_OP_425J2_127_3477_n3024), .Y(n701) );
  NBUFFX8_HVT U1320 ( .A(DP_OP_425J2_127_3477_n3024), .Y(n704) );
  NAND2X0_HVT U1321 ( .A1(n711), .A2(conv1_sram_rdata_weight[9]), .Y(n706) );
  AND2X1_HVT U1322 ( .A1(n705), .A2(src_window[65]), .Y(n7001) );
  NBUFFX2_HVT U1323 ( .A(DP_OP_425J2_127_3477_n3024), .Y(n702) );
  OA21X2_HVT U1324 ( .A1(n711), .A2(n707), .A3(n706), .Y(
        DP_OP_425J2_127_3477_n3024) );
  INVX4_HVT U1325 ( .A(conv2_sram_rdata_weight[9]), .Y(n707) );
  OR2X1_HVT U1326 ( .A1(n708), .A2(n709), .Y(n1048) );
  NAND2X0_HVT U1327 ( .A1(n709), .A2(n708), .Y(n1047) );
  NAND2X0_HVT U1328 ( .A1(DP_OP_424J2_126_3477_n285), .A2(
        DP_OP_424J2_126_3477_n185), .Y(n708) );
  NAND2X0_HVT U1329 ( .A1(n710), .A2(DP_OP_424J2_126_3477_n190), .Y(n709) );
  NAND2X0_HVT U1330 ( .A1(n1518), .A2(DP_OP_424J2_126_3477_n187), .Y(n710) );
  NBUFFX8_HVT U1331 ( .A(n4), .Y(n711) );
  INVX2_HVT U1332 ( .A(n726), .Y(DP_OP_422J2_124_3477_n2759) );
  AND2X1_HVT U1333 ( .A1(n726), .A2(n712), .Y(DP_OP_423J2_125_3477_n2729) );
  INVX2_HVT U1334 ( .A(DP_OP_425J2_127_3477_n2401), .Y(n712) );
  INVX2_HVT U1335 ( .A(n1923), .Y(n713) );
  NBUFFX2_HVT U1336 ( .A(conv_weight_box[39]), .Y(n714) );
  AND2X1_HVT U1337 ( .A1(conv_weight_box[39]), .A2(n715), .Y(
        DP_OP_424J2_126_3477_n2737) );
  INVX2_HVT U1338 ( .A(DP_OP_422J2_124_3477_n2181), .Y(n715) );
  NAND2X0_HVT U1339 ( .A1(conv_weight_box[39]), .A2(n716), .Y(
        DP_OP_424J2_126_3477_n2734) );
  INVX2_HVT U1340 ( .A(DP_OP_422J2_124_3477_n2178), .Y(n716) );
  AND2X1_HVT U1341 ( .A1(n714), .A2(n717), .Y(DP_OP_423J2_125_3477_n2740) );
  INVX2_HVT U1342 ( .A(DP_OP_423J2_125_3477_n2756), .Y(n717) );
  AND2X1_HVT U1343 ( .A1(n714), .A2(n718), .Y(DP_OP_423J2_125_3477_n2735) );
  INVX2_HVT U1344 ( .A(DP_OP_423J2_125_3477_n2751), .Y(n718) );
  AND2X1_HVT U1345 ( .A1(n714), .A2(n719), .Y(DP_OP_423J2_125_3477_n2736) );
  INVX2_HVT U1346 ( .A(DP_OP_422J2_124_3477_n2268), .Y(n719) );
  AND2X1_HVT U1347 ( .A1(n714), .A2(n720), .Y(DP_OP_423J2_125_3477_n2737) );
  INVX2_HVT U1348 ( .A(DP_OP_425J2_127_3477_n2401), .Y(n720) );
  NAND2X0_HVT U1349 ( .A1(n714), .A2(n721), .Y(DP_OP_423J2_125_3477_n2734) );
  INVX2_HVT U1350 ( .A(DP_OP_423J2_125_3477_n2750), .Y(n721) );
  AND2X1_HVT U1351 ( .A1(n714), .A2(n722), .Y(DP_OP_424J2_126_3477_n2741) );
  INVX2_HVT U1352 ( .A(DP_OP_422J2_124_3477_n2185), .Y(n722) );
  AND2X1_HVT U1353 ( .A1(n714), .A2(n723), .Y(DP_OP_423J2_125_3477_n2739) );
  INVX2_HVT U1354 ( .A(DP_OP_424J2_126_3477_n2667), .Y(n723) );
  AND2X1_HVT U1355 ( .A1(n714), .A2(n724), .Y(DP_OP_423J2_125_3477_n2738) );
  INVX2_HVT U1356 ( .A(DP_OP_423J2_125_3477_n2754), .Y(n724) );
  AND2X4_HVT U1357 ( .A1(n714), .A2(n725), .Y(DP_OP_423J2_125_3477_n2741) );
  INVX2_HVT U1358 ( .A(DP_OP_423J2_125_3477_n2757), .Y(n725) );
  NBUFFX2_HVT U1359 ( .A(n726), .Y(n727) );
  INVX2_HVT U1360 ( .A(DP_OP_422J2_124_3477_n2185), .Y(n728) );
  AND2X1_HVT U1361 ( .A1(n726), .A2(n729), .Y(DP_OP_424J2_126_3477_n2728) );
  INVX2_HVT U1362 ( .A(DP_OP_424J2_126_3477_n2752), .Y(n729) );
  AND2X1_HVT U1363 ( .A1(n727), .A2(n730), .Y(DP_OP_423J2_125_3477_n2733) );
  INVX2_HVT U1364 ( .A(DP_OP_423J2_125_3477_n2757), .Y(n730) );
  AND2X1_HVT U1365 ( .A1(n727), .A2(n731), .Y(DP_OP_424J2_126_3477_n2731) );
  INVX2_HVT U1366 ( .A(DP_OP_422J2_124_3477_n2183), .Y(n731) );
  NAND2X0_HVT U1367 ( .A1(n727), .A2(n732), .Y(DP_OP_423J2_125_3477_n2726) );
  INVX2_HVT U1368 ( .A(DP_OP_423J2_125_3477_n2750), .Y(n732) );
  AND2X1_HVT U1369 ( .A1(n727), .A2(n733), .Y(DP_OP_425J2_127_3477_n2731) );
  INVX2_HVT U1370 ( .A(DP_OP_425J2_127_3477_n2755), .Y(n733) );
  AND2X1_HVT U1371 ( .A1(n727), .A2(n734), .Y(DP_OP_423J2_125_3477_n2727) );
  INVX2_HVT U1372 ( .A(DP_OP_423J2_125_3477_n2751), .Y(n734) );
  AND2X1_HVT U1373 ( .A1(n727), .A2(n735), .Y(DP_OP_422J2_124_3477_n2727) );
  INVX2_HVT U1374 ( .A(DP_OP_422J2_124_3477_n2751), .Y(n735) );
  AND2X4_HVT U1375 ( .A1(n727), .A2(n736), .Y(DP_OP_424J2_126_3477_n2727) );
  INVX2_HVT U1376 ( .A(DP_OP_422J2_124_3477_n2179), .Y(n736) );
  INVX0_HVT U1377 ( .A(n737), .Y(DP_OP_424J2_126_3477_n2730) );
  NBUFFX2_HVT U1378 ( .A(n726), .Y(n738) );
  INVX4_HVT U1379 ( .A(DP_OP_424J2_126_3477_n2754), .Y(n739) );
  INVX2_HVT U1380 ( .A(DP_OP_422J2_124_3477_n2753), .Y(n740) );
  AND2X1_HVT U1381 ( .A1(n738), .A2(n741), .Y(DP_OP_423J2_125_3477_n2728) );
  INVX2_HVT U1382 ( .A(DP_OP_425J2_127_3477_n2400), .Y(n741) );
  AND2X1_HVT U1383 ( .A1(n738), .A2(n742), .Y(DP_OP_425J2_127_3477_n2730) );
  INVX2_HVT U1384 ( .A(DP_OP_425J2_127_3477_n2754), .Y(n742) );
  AND2X1_HVT U1385 ( .A1(n738), .A2(n743), .Y(DP_OP_424J2_126_3477_n2729) );
  INVX2_HVT U1386 ( .A(DP_OP_422J2_124_3477_n2181), .Y(n743) );
  AND2X1_HVT U1387 ( .A1(n738), .A2(n744), .Y(DP_OP_423J2_125_3477_n2730) );
  INVX2_HVT U1388 ( .A(DP_OP_423J2_125_3477_n2754), .Y(n744) );
  AND2X1_HVT U1389 ( .A1(n738), .A2(n745), .Y(DP_OP_425J2_127_3477_n2729) );
  INVX2_HVT U1390 ( .A(DP_OP_424J2_126_3477_n2269), .Y(n745) );
  AND2X1_HVT U1391 ( .A1(n738), .A2(n746), .Y(DP_OP_424J2_126_3477_n2732) );
  INVX2_HVT U1392 ( .A(DP_OP_424J2_126_3477_n2756), .Y(n746) );
  NAND2X0_HVT U1393 ( .A1(n738), .A2(n747), .Y(DP_OP_422J2_124_3477_n2726) );
  INVX2_HVT U1394 ( .A(DP_OP_422J2_124_3477_n2750), .Y(n747) );
  NAND2X0_HVT U1395 ( .A1(n738), .A2(n748), .Y(DP_OP_424J2_126_3477_n2726) );
  INVX2_HVT U1396 ( .A(DP_OP_422J2_124_3477_n2178), .Y(n748) );
  AND2X1_HVT U1397 ( .A1(n738), .A2(n749), .Y(DP_OP_422J2_124_3477_n2731) );
  INVX2_HVT U1398 ( .A(DP_OP_424J2_126_3477_n2403), .Y(n749) );
  NAND2X0_HVT U1399 ( .A1(n738), .A2(n750), .Y(DP_OP_425J2_127_3477_n2726) );
  INVX2_HVT U1400 ( .A(DP_OP_423J2_125_3477_n2178), .Y(n750) );
  MUX21X2_HVT U1401 ( .A1(conv2_sram_rdata_weight[47]), .A2(
        conv1_sram_rdata_weight[47]), .S0(n241), .Y(conv_weight_box[32]) );
  INVX2_HVT U1402 ( .A(DP_OP_422J2_124_3477_n2448), .Y(n751) );
  INVX2_HVT U1403 ( .A(DP_OP_422J2_124_3477_n2619), .Y(n752) );
  NAND2X0_HVT U1404 ( .A1(n769), .A2(n790), .Y(n753) );
  INVX2_HVT U1405 ( .A(n791), .Y(n754) );
  INVX2_HVT U1406 ( .A(DP_OP_424J2_126_3477_n2667), .Y(n756) );
  INVX2_HVT U1407 ( .A(DP_OP_424J2_126_3477_n2669), .Y(n757) );
  NAND2X0_HVT U1408 ( .A1(n88), .A2(n758), .Y(DP_OP_424J2_126_3477_n2636) );
  INVX2_HVT U1409 ( .A(DP_OP_423J2_125_3477_n2756), .Y(n758) );
  NAND2X0_HVT U1410 ( .A1(n87), .A2(n759), .Y(DP_OP_424J2_126_3477_n2633) );
  INVX2_HVT U1411 ( .A(DP_OP_425J2_127_3477_n2401), .Y(n759) );
  NAND2X0_HVT U1412 ( .A1(n88), .A2(n760), .Y(DP_OP_424J2_126_3477_n2634) );
  INVX2_HVT U1413 ( .A(DP_OP_422J2_124_3477_n2270), .Y(n760) );
  NAND2X0_HVT U1414 ( .A1(n88), .A2(n761), .Y(DP_OP_425J2_127_3477_n2635) );
  INVX2_HVT U1415 ( .A(DP_OP_422J2_124_3477_n2799), .Y(n761) );
  NAND2X0_HVT U1416 ( .A1(n88), .A2(n762), .Y(DP_OP_424J2_126_3477_n2632) );
  INVX2_HVT U1417 ( .A(DP_OP_425J2_127_3477_n2400), .Y(n762) );
  NAND2X0_HVT U1418 ( .A1(n88), .A2(n763), .Y(DP_OP_425J2_127_3477_n2637) );
  INVX2_HVT U1419 ( .A(DP_OP_422J2_124_3477_n2801), .Y(n763) );
  NAND2X0_HVT U1420 ( .A1(n88), .A2(n764), .Y(DP_OP_425J2_127_3477_n2636) );
  INVX2_HVT U1421 ( .A(DP_OP_422J2_124_3477_n2800), .Y(n764) );
  NAND2X0_HVT U1422 ( .A1(n88), .A2(n765), .Y(DP_OP_424J2_126_3477_n2631) );
  INVX2_HVT U1423 ( .A(DP_OP_422J2_124_3477_n2267), .Y(n765) );
  NAND2X0_HVT U1424 ( .A1(n88), .A2(n766), .Y(DP_OP_425J2_127_3477_n2631) );
  INVX2_HVT U1425 ( .A(DP_OP_423J2_125_3477_n2267), .Y(n766) );
  AND2X4_HVT U1426 ( .A1(n88), .A2(n767), .Y(DP_OP_424J2_126_3477_n2630) );
  INVX2_HVT U1427 ( .A(DP_OP_423J2_125_3477_n2750), .Y(n767) );
  INVX2_HVT U1428 ( .A(n951), .Y(n952) );
  MUX21X2_HVT U1429 ( .A1(conv2_sram_rdata_weight[42]), .A2(
        conv1_sram_rdata_weight[42]), .S0(n240), .Y(conv_weight_box[28]) );
  OR2X4_HVT U1430 ( .A1(mode[0]), .A2(n951), .Y(n1923) );
  NBUFFX2_HVT U1431 ( .A(n4), .Y(n769) );
  INVX8_HVT U1432 ( .A(n1923), .Y(n1396) );
  FADDX1_HVT U1433 ( .A(DP_OP_424J2_126_3477_n1313), .B(
        DP_OP_424J2_126_3477_n1317), .CI(DP_OP_424J2_126_3477_n1474), .CO(
        DP_OP_424J2_126_3477_n1268) );
  NBUFFX2_HVT U1434 ( .A(n772), .Y(n770) );
  NBUFFX8_HVT U1435 ( .A(DP_OP_425J2_127_3477_n2539), .Y(n771) );
  NBUFFX16_HVT U1436 ( .A(DP_OP_425J2_127_3477_n2539), .Y(n772) );
  OA21X2_HVT U1437 ( .A1(n711), .A2(n774), .A3(n773), .Y(
        DP_OP_425J2_127_3477_n2539) );
  NAND2X0_HVT U1438 ( .A1(n711), .A2(conv1_sram_rdata_weight[98]), .Y(n773) );
  INVX2_HVT U1439 ( .A(conv2_sram_rdata_weight[98]), .Y(n774) );
  NBUFFX2_HVT U1440 ( .A(n30), .Y(n775) );
  NBUFFX2_HVT U1441 ( .A(n779), .Y(n776) );
  NBUFFX2_HVT U1442 ( .A(n779), .Y(n777) );
  INVX2_HVT U1443 ( .A(n779), .Y(n778) );
  NAND2X0_HVT U1444 ( .A1(n711), .A2(conv1_sram_rdata_weight[15]), .Y(n780) );
  INVX2_HVT U1445 ( .A(conv2_sram_rdata_weight[15]), .Y(n781) );
  INVX2_HVT U1446 ( .A(DP_OP_424J2_126_3477_n2752), .Y(n782) );
  INVX2_HVT U1447 ( .A(DP_OP_424J2_126_3477_n2887), .Y(n783) );
  INVX4_HVT U1448 ( .A(n844), .Y(n784) );
  INVX4_HVT U1449 ( .A(n845), .Y(n785) );
  INVX2_HVT U1450 ( .A(conv_weight_box[50]), .Y(DP_OP_425J2_127_3477_n2671) );
  AND2X1_HVT U1451 ( .A1(conv_weight_box[50]), .A2(n786), .Y(
        DP_OP_422J2_124_3477_n2645) );
  INVX2_HVT U1452 ( .A(DP_OP_422J2_124_3477_n2669), .Y(n786) );
  MUX21X1_HVT U1453 ( .A1(conv1_sram_rdata_weight[74]), .A2(
        conv2_sram_rdata_weight[74]), .S0(n1396), .Y(conv_weight_box[50]) );
  INVX4_HVT U1454 ( .A(n1923), .Y(n858) );
  INVX2_HVT U1455 ( .A(conv_weight_box[5]), .Y(DP_OP_424J2_126_3477_n3025) );
  MUX21X1_HVT U1456 ( .A1(n788), .A2(n787), .S0(n858), .Y(conv_weight_box[5])
         );
  INVX2_HVT U1457 ( .A(n847), .Y(n787) );
  INVX2_HVT U1458 ( .A(n848), .Y(n788) );
  INVX2_HVT U1459 ( .A(conv1_sram_rdata_weight[86]), .Y(n790) );
  INVX2_HVT U1460 ( .A(conv2_sram_rdata_weight[86]), .Y(n791) );
  NBUFFX2_HVT U1461 ( .A(n799), .Y(n792) );
  NBUFFX2_HVT U1462 ( .A(n799), .Y(n793) );
  NBUFFX2_HVT U1463 ( .A(n799), .Y(n794) );
  NBUFFX2_HVT U1464 ( .A(n799), .Y(n795) );
  IBUFFX32_HVT U1465 ( .A(src_window[227]), .Y(n796) );
  NBUFFX2_HVT U1466 ( .A(DP_OP_422J2_124_3477_n2407), .Y(n797) );
  NBUFFX8_HVT U1467 ( .A(DP_OP_422J2_124_3477_n2407), .Y(n798) );
  NBUFFX16_HVT U1468 ( .A(DP_OP_422J2_124_3477_n2407), .Y(n799) );
  NAND2X0_HVT U1469 ( .A1(n857), .A2(conv1_sram_rdata_weight[78]), .Y(n800) );
  NOR2X0_HVT U1470 ( .A1(n798), .A2(n796), .Y(DP_OP_423J2_125_3477_n2378) );
  OA21X2_HVT U1471 ( .A1(n857), .A2(n801), .A3(n800), .Y(
        DP_OP_422J2_124_3477_n2407) );
  INVX4_HVT U1472 ( .A(conv2_sram_rdata_weight[78]), .Y(n801) );
  AND2X1_HVT U1473 ( .A1(n1715), .A2(n1733), .Y(n805) );
  NAND3X0_HVT U1474 ( .A1(n1042), .A2(n1714), .A3(n1713), .Y(n1733) );
  OA21X1_HVT U1475 ( .A1(DP_OP_424J2_126_3477_n240), .A2(
        DP_OP_424J2_126_3477_n236), .A3(DP_OP_424J2_126_3477_n237), .Y(n1715)
         );
  AND3X1_HVT U1476 ( .A1(n804), .A2(n803), .A3(n1357), .Y(n802) );
  NAND2X0_HVT U1477 ( .A1(n807), .A2(n1067), .Y(n803) );
  NAND3X0_HVT U1478 ( .A1(n807), .A2(n1712), .A3(n1711), .Y(n804) );
  NAND3X0_HVT U1479 ( .A1(n807), .A2(n1732), .A3(n1711), .Y(n806) );
  AND2X1_HVT U1480 ( .A1(DP_OP_424J2_126_3477_n419), .A2(
        DP_OP_424J2_126_3477_n512), .Y(n1712) );
  OR2X1_HVT U1481 ( .A1(DP_OP_424J2_126_3477_n512), .A2(
        DP_OP_424J2_126_3477_n419), .Y(n1732) );
  AND2X1_HVT U1482 ( .A1(n1745), .A2(n1752), .Y(n807) );
  NAND2X0_HVT U1483 ( .A1(n1773), .A2(n1772), .Y(n808) );
  OR2X1_HVT U1484 ( .A1(DP_OP_425J2_127_3477_n822), .A2(
        DP_OP_425J2_127_3477_n649), .Y(n1773) );
  AND2X1_HVT U1485 ( .A1(n809), .A2(DP_OP_425J2_127_3477_n249), .Y(
        DP_OP_425J2_127_3477_n245) );
  NAND2X0_HVT U1486 ( .A1(DP_OP_425J2_127_3477_n250), .A2(
        DP_OP_425J2_127_3477_n295), .Y(n809) );
  INVX2_HVT U1487 ( .A(n1794), .Y(n810) );
  OR2X1_HVT U1488 ( .A1(DP_OP_425J2_127_3477_n1018), .A2(
        DP_OP_425J2_127_3477_n823), .Y(n1794) );
  AO22X1_HVT U1489 ( .A1(DP_OP_423J2_125_3477_n523), .A2(
        DP_OP_423J2_125_3477_n656), .A3(DP_OP_423J2_125_3477_n654), .A4(n811), 
        .Y(DP_OP_423J2_125_3477_n516) );
  OR2X1_HVT U1490 ( .A1(DP_OP_423J2_125_3477_n656), .A2(
        DP_OP_423J2_125_3477_n523), .Y(n811) );
  XOR3X2_HVT U1491 ( .A1(DP_OP_423J2_125_3477_n523), .A2(
        DP_OP_423J2_125_3477_n656), .A3(DP_OP_423J2_125_3477_n654), .Y(
        DP_OP_423J2_125_3477_n517) );
  INVX2_HVT U1492 ( .A(n814), .Y(DP_OP_424J2_126_3477_n259) );
  NAND2X0_HVT U1493 ( .A1(n812), .A2(DP_OP_424J2_126_3477_n260), .Y(n1736) );
  NAND2X0_HVT U1494 ( .A1(n814), .A2(n813), .Y(n812) );
  INVX2_HVT U1495 ( .A(DP_OP_424J2_126_3477_n261), .Y(n813) );
  OR2X1_HVT U1496 ( .A1(DP_OP_424J2_126_3477_n1579), .A2(
        DP_OP_424J2_126_3477_n1577), .Y(n814) );
  AND2X1_HVT U1497 ( .A1(n824), .A2(n815), .Y(DP_OP_422J2_124_3477_n2344) );
  INVX2_HVT U1498 ( .A(DP_OP_424J2_126_3477_n2580), .Y(n815) );
  AND2X1_HVT U1499 ( .A1(n824), .A2(n816), .Y(DP_OP_424J2_126_3477_n2340) );
  INVX2_HVT U1500 ( .A(DP_OP_422J2_124_3477_n2796), .Y(n816) );
  OR2X1_HVT U1501 ( .A1(DP_OP_423J2_125_3477_n2354), .A2(n825), .Y(
        DP_OP_423J2_125_3477_n2338) );
  AND2X1_HVT U1502 ( .A1(n824), .A2(n817), .Y(DP_OP_424J2_126_3477_n2345) );
  INVX2_HVT U1503 ( .A(DP_OP_423J2_125_3477_n2273), .Y(n817) );
  AND2X1_HVT U1504 ( .A1(n824), .A2(n818), .Y(DP_OP_423J2_125_3477_n2341) );
  INVX2_HVT U1505 ( .A(DP_OP_422J2_124_3477_n2709), .Y(n818) );
  AND2X1_HVT U1506 ( .A1(n824), .A2(n819), .Y(DP_OP_423J2_125_3477_n2342) );
  INVX2_HVT U1507 ( .A(DP_OP_422J2_124_3477_n2710), .Y(n819) );
  AND2X1_HVT U1508 ( .A1(n824), .A2(n820), .Y(DP_OP_425J2_127_3477_n2345) );
  INVX2_HVT U1509 ( .A(DP_OP_423J2_125_3477_n2801), .Y(n820) );
  AND2X1_HVT U1510 ( .A1(n824), .A2(n821), .Y(DP_OP_422J2_124_3477_n2345) );
  INVX2_HVT U1511 ( .A(DP_OP_423J2_125_3477_n2669), .Y(n821) );
  AND2X1_HVT U1512 ( .A1(n824), .A2(n822), .Y(DP_OP_423J2_125_3477_n2339) );
  INVX2_HVT U1513 ( .A(DP_OP_424J2_126_3477_n2443), .Y(n822) );
  AND2X1_HVT U1514 ( .A1(n824), .A2(n823), .Y(DP_OP_425J2_127_3477_n2339) );
  INVX2_HVT U1515 ( .A(DP_OP_423J2_125_3477_n2795), .Y(n823) );
  INVX2_HVT U1516 ( .A(n825), .Y(n824) );
  NBUFFX2_HVT U1517 ( .A(DP_OP_423J2_125_3477_n2364), .Y(n825) );
  FADDX1_HVT U1518 ( .A(n826), .B(DP_OP_424J2_126_3477_n2950), .CI(
        DP_OP_424J2_126_3477_n2033), .CO(DP_OP_424J2_126_3477_n1368) );
  XOR3X2_HVT U1519 ( .A1(DP_OP_424J2_126_3477_n2950), .A2(n826), .A3(
        DP_OP_424J2_126_3477_n2033), .Y(DP_OP_424J2_126_3477_n1369) );
  AND2X1_HVT U1520 ( .A1(n1387), .A2(n827), .Y(n826) );
  INVX2_HVT U1521 ( .A(DP_OP_423J2_125_3477_n2269), .Y(n827) );
  INVX2_HVT U1522 ( .A(DP_OP_423J2_125_3477_n2364), .Y(n1387) );
  FADDX1_HVT U1523 ( .A(DP_OP_424J2_126_3477_n1267), .B(
        DP_OP_424J2_126_3477_n1271), .CI(DP_OP_424J2_126_3477_n1273), .CO(
        DP_OP_424J2_126_3477_n1240) );
  INVX2_HVT U1524 ( .A(conv_weight_box[22]), .Y(DP_OP_425J2_127_3477_n2891) );
  AND2X1_HVT U1525 ( .A1(conv_weight_box[22]), .A2(n828), .Y(
        DP_OP_424J2_126_3477_n2864) );
  INVX2_HVT U1526 ( .A(DP_OP_423J2_125_3477_n2976), .Y(n828) );
  NAND2X0_HVT U1527 ( .A1(n829), .A2(n888), .Y(DP_OP_423J2_125_3477_n686) );
  NAND2X0_HVT U1528 ( .A1(n830), .A2(DP_OP_423J2_125_3477_n711), .Y(n829) );
  OR2X1_HVT U1529 ( .A1(DP_OP_423J2_125_3477_n878), .A2(
        DP_OP_423J2_125_3477_n876), .Y(n830) );
  INVX2_HVT U1530 ( .A(n832), .Y(n1231) );
  INVX2_HVT U1531 ( .A(DP_OP_423J2_125_3477_n753), .Y(n831) );
  INVX2_HVT U1532 ( .A(n1614), .Y(n833) );
  IBUFFX32_HVT U1533 ( .A(n841), .Y(n834) );
  NAND3X0_HVT U1534 ( .A1(n840), .A2(n838), .A3(n835), .Y(n_conv2_sum_b[18])
         );
  AO22X1_HVT U1535 ( .A1(n1681), .A2(n837), .A3(n836), .A4(n842), .Y(n835) );
  INVX2_HVT U1536 ( .A(n1681), .Y(n836) );
  NAND2X0_HVT U1537 ( .A1(n1674), .A2(n921), .Y(n837) );
  NAND2X0_HVT U1538 ( .A1(n1614), .A2(n839), .Y(n838) );
  AND2X1_HVT U1539 ( .A1(n1681), .A2(n921), .Y(n839) );
  NAND2X0_HVT U1540 ( .A1(n834), .A2(n833), .Y(n840) );
  OR2X1_HVT U1541 ( .A1(n842), .A2(n1674), .Y(n841) );
  INVX2_HVT U1542 ( .A(DP_OP_423J2_125_3477_n19), .Y(n842) );
  NBUFFX8_HVT U1543 ( .A(n4), .Y(n843) );
  INVX2_HVT U1544 ( .A(conv1_sram_rdata_weight[31]), .Y(n844) );
  INVX2_HVT U1545 ( .A(conv2_sram_rdata_weight[31]), .Y(n845) );
  NBUFFX8_HVT U1546 ( .A(DP_OP_424J2_126_3477_n3025), .Y(n846) );
  INVX2_HVT U1547 ( .A(conv2_sram_rdata_weight[8]), .Y(n847) );
  INVX2_HVT U1548 ( .A(conv1_sram_rdata_weight[8]), .Y(n848) );
  INVX2_HVT U1549 ( .A(DP_OP_424J2_126_3477_n3063), .Y(n849) );
  AO22X1_HVT U1550 ( .A1(DP_OP_422J2_124_3477_n1874), .A2(
        DP_OP_422J2_124_3477_n1878), .A3(DP_OP_422J2_124_3477_n1807), .A4(n850), .Y(DP_OP_422J2_124_3477_n1772) );
  NAND2X0_HVT U1551 ( .A1(n852), .A2(n851), .Y(n850) );
  INVX2_HVT U1552 ( .A(DP_OP_422J2_124_3477_n1874), .Y(n851) );
  INVX2_HVT U1553 ( .A(DP_OP_422J2_124_3477_n1878), .Y(n852) );
  XOR3X2_HVT U1554 ( .A1(DP_OP_422J2_124_3477_n1874), .A2(
        DP_OP_422J2_124_3477_n1878), .A3(DP_OP_422J2_124_3477_n1807), .Y(
        DP_OP_422J2_124_3477_n1773) );
  INVX2_HVT U1555 ( .A(conv_weight_box[22]), .Y(DP_OP_424J2_126_3477_n2891) );
  AND2X1_HVT U1556 ( .A1(conv_weight_box[22]), .A2(n853), .Y(
        DP_OP_425J2_127_3477_n2864) );
  INVX2_HVT U1557 ( .A(DP_OP_425J2_127_3477_n2888), .Y(n853) );
  MUX21X1_HVT U1558 ( .A1(n854), .A2(n1365), .S0(n1928), .Y(
        DP_OP_423J2_125_3477_n2538) );
  INVX2_HVT U1559 ( .A(conv1_sram_rdata_weight[99]), .Y(n854) );
  INVX4_HVT U1560 ( .A(conv2_sram_rdata_weight[93]), .Y(n855) );
  INVX4_HVT U1561 ( .A(conv1_sram_rdata_weight[93]), .Y(n856) );
  INVX2_HVT U1562 ( .A(DP_OP_424J2_126_3477_n2365), .Y(conv_weight_box[47]) );
  AO22X1_HVT U1563 ( .A1(n860), .A2(n859), .A3(n952), .A4(n861), .Y(
        DP_OP_424J2_126_3477_n2365) );
  INVX2_HVT U1564 ( .A(n862), .Y(n859) );
  NAND2X0_HVT U1565 ( .A1(n952), .A2(n1516), .Y(n860) );
  AND2X1_HVT U1566 ( .A1(n863), .A2(n1516), .Y(n861) );
  INVX2_HVT U1567 ( .A(n864), .Y(n862) );
  INVX2_HVT U1568 ( .A(conv2_sram_rdata_weight[68]), .Y(n863) );
  INVX2_HVT U1569 ( .A(conv1_sram_rdata_weight[68]), .Y(n864) );
  AO22X2_HVT U1570 ( .A1(n1533), .A2(n1850), .A3(n1849), .A4(n1483), .Y(n2153)
         );
  INVX2_HVT U1571 ( .A(tmp_big1[7]), .Y(n2171) );
  HADDX2_HVT U1572 ( .A0(n1267), .B0(DP_OP_424J2_126_3477_n250), .SO(
        n_conv2_sum_c[6]) );
  HADDX2_HVT U1573 ( .A0(n1222), .B0(n1737), .SO(n_conv2_sum_c[5]) );
  NOR2X2_HVT U1574 ( .A1(DP_OP_423J2_125_3477_n2801), .A2(
        DP_OP_424J2_126_3477_n2365), .Y(DP_OP_425J2_127_3477_n2353) );
  OR2X4_HVT U1575 ( .A1(DP_OP_423J2_125_3477_n2794), .A2(
        DP_OP_424J2_126_3477_n2365), .Y(DP_OP_425J2_127_3477_n2346) );
  NOR2X2_HVT U1576 ( .A1(DP_OP_423J2_125_3477_n2800), .A2(
        DP_OP_424J2_126_3477_n2365), .Y(DP_OP_425J2_127_3477_n2352) );
  NOR2X2_HVT U1577 ( .A1(DP_OP_425J2_127_3477_n2356), .A2(
        DP_OP_424J2_126_3477_n2365), .Y(DP_OP_425J2_127_3477_n2348) );
  NOR2X2_HVT U1578 ( .A1(DP_OP_425J2_127_3477_n2359), .A2(
        DP_OP_424J2_126_3477_n2365), .Y(DP_OP_425J2_127_3477_n2351) );
  OR2X4_HVT U1579 ( .A1(DP_OP_422J2_124_3477_n2354), .A2(
        DP_OP_424J2_126_3477_n2365), .Y(DP_OP_422J2_124_3477_n2346) );
  NOR2X2_HVT U1580 ( .A1(DP_OP_423J2_125_3477_n2269), .A2(
        DP_OP_424J2_126_3477_n2365), .Y(DP_OP_424J2_126_3477_n2349) );
  NOR2X2_HVT U1581 ( .A1(DP_OP_423J2_125_3477_n2267), .A2(
        DP_OP_424J2_126_3477_n2365), .Y(DP_OP_424J2_126_3477_n2347) );
  IBUFFX4_HVT U1582 ( .A(n1961), .Y(n1496) );
  OR2X2_HVT U1583 ( .A1(DP_OP_425J2_127_3477_n1968), .A2(N7), .Y(n2175) );
  OR2X1_HVT U1584 ( .A1(n1524), .A2(conv2_sum_a[11]), .Y(n2025) );
  OA22X1_HVT U1585 ( .A1(n1326), .A2(conv2_sum_a[30]), .A3(n1323), .A4(
        conv2_sum_b[31]), .Y(n865) );
  IBUFFX16_HVT U1586 ( .A(n865), .Y(n2007) );
  XOR3X2_HVT U1587 ( .A1(DP_OP_422J2_124_3477_n689), .A2(
        DP_OP_422J2_124_3477_n854), .A3(DP_OP_422J2_124_3477_n687), .Y(
        DP_OP_422J2_124_3477_n671) );
  NAND2X0_HVT U1588 ( .A1(DP_OP_422J2_124_3477_n689), .A2(
        DP_OP_422J2_124_3477_n687), .Y(n866) );
  NAND2X0_HVT U1589 ( .A1(DP_OP_422J2_124_3477_n854), .A2(
        DP_OP_422J2_124_3477_n687), .Y(n867) );
  NAND2X0_HVT U1590 ( .A1(DP_OP_422J2_124_3477_n854), .A2(
        DP_OP_422J2_124_3477_n689), .Y(n868) );
  NAND3X2_HVT U1591 ( .A1(n868), .A2(n867), .A3(n866), .Y(
        DP_OP_422J2_124_3477_n670) );
  XOR3X2_HVT U1592 ( .A1(DP_OP_422J2_124_3477_n956), .A2(
        DP_OP_422J2_124_3477_n958), .A3(DP_OP_422J2_124_3477_n962), .Y(
        DP_OP_422J2_124_3477_n753) );
  NAND2X0_HVT U1593 ( .A1(DP_OP_422J2_124_3477_n956), .A2(
        DP_OP_422J2_124_3477_n962), .Y(n869) );
  NAND2X0_HVT U1594 ( .A1(DP_OP_422J2_124_3477_n958), .A2(
        DP_OP_422J2_124_3477_n962), .Y(n870) );
  NAND2X0_HVT U1595 ( .A1(DP_OP_422J2_124_3477_n958), .A2(
        DP_OP_422J2_124_3477_n956), .Y(n871) );
  NAND3X0_HVT U1596 ( .A1(n871), .A2(n870), .A3(n869), .Y(
        DP_OP_422J2_124_3477_n752) );
  OA21X1_HVT U1597 ( .A1(n1418), .A2(n1376), .A3(n1375), .Y(n872) );
  OA21X1_HVT U1598 ( .A1(n1418), .A2(n1376), .A3(n1375), .Y(n873) );
  NBUFFX4_HVT U1599 ( .A(n872), .Y(n874) );
  NBUFFX4_HVT U1600 ( .A(n873), .Y(n875) );
  NBUFFX4_HVT U1601 ( .A(DP_OP_423J2_125_3477_n2363), .Y(n876) );
  OA21X1_HVT U1602 ( .A1(n1418), .A2(n1376), .A3(n1375), .Y(
        DP_OP_423J2_125_3477_n2363) );
  XOR3X2_HVT U1603 ( .A1(DP_OP_424J2_126_3477_n956), .A2(
        DP_OP_424J2_126_3477_n958), .A3(DP_OP_424J2_126_3477_n962), .Y(
        DP_OP_424J2_126_3477_n753) );
  NAND2X0_HVT U1604 ( .A1(DP_OP_424J2_126_3477_n956), .A2(
        DP_OP_424J2_126_3477_n962), .Y(n877) );
  NAND2X0_HVT U1605 ( .A1(DP_OP_424J2_126_3477_n958), .A2(
        DP_OP_424J2_126_3477_n962), .Y(n878) );
  NAND2X1_HVT U1606 ( .A1(DP_OP_424J2_126_3477_n958), .A2(
        DP_OP_424J2_126_3477_n956), .Y(n879) );
  NAND3X2_HVT U1607 ( .A1(n879), .A2(n878), .A3(n877), .Y(
        DP_OP_424J2_126_3477_n752) );
  XOR3X2_HVT U1608 ( .A1(DP_OP_424J2_126_3477_n686), .A2(
        DP_OP_424J2_126_3477_n684), .A3(DP_OP_424J2_126_3477_n553), .Y(
        DP_OP_424J2_126_3477_n537) );
  NAND2X0_HVT U1609 ( .A1(DP_OP_424J2_126_3477_n686), .A2(
        DP_OP_424J2_126_3477_n553), .Y(n880) );
  NAND2X0_HVT U1610 ( .A1(DP_OP_424J2_126_3477_n684), .A2(
        DP_OP_424J2_126_3477_n553), .Y(n881) );
  NAND2X0_HVT U1611 ( .A1(DP_OP_424J2_126_3477_n686), .A2(
        DP_OP_424J2_126_3477_n684), .Y(n882) );
  NAND3X0_HVT U1612 ( .A1(n882), .A2(n881), .A3(n880), .Y(
        DP_OP_424J2_126_3477_n536) );
  XOR3X2_HVT U1613 ( .A1(DP_OP_425J2_127_3477_n423), .A2(
        DP_OP_425J2_127_3477_n514), .A3(DP_OP_425J2_127_3477_n421), .Y(
        DP_OP_425J2_127_3477_n419) );
  NAND2X0_HVT U1614 ( .A1(DP_OP_425J2_127_3477_n423), .A2(
        DP_OP_425J2_127_3477_n421), .Y(n883) );
  NAND2X0_HVT U1615 ( .A1(DP_OP_425J2_127_3477_n421), .A2(
        DP_OP_425J2_127_3477_n514), .Y(n884) );
  NAND2X0_HVT U1616 ( .A1(DP_OP_425J2_127_3477_n514), .A2(
        DP_OP_425J2_127_3477_n423), .Y(n885) );
  NAND3X0_HVT U1617 ( .A1(n885), .A2(n884), .A3(n883), .Y(
        DP_OP_425J2_127_3477_n418) );
  XOR2X1_HVT U1618 ( .A1(n1580), .A2(n1259), .Y(n_conv2_sum_a[14]) );
  INVX2_HVT U1619 ( .A(n1874), .Y(n886) );
  INVX1_HVT U1620 ( .A(n1975), .Y(n887) );
  MUX21X1_HVT U1621 ( .A1(tmp_big2[14]), .A2(tmp_big1[14]), .S0(N9), .Y(
        data_out[14]) );
  XOR3X2_HVT U1622 ( .A1(DP_OP_424J2_126_3477_n1267), .A2(
        DP_OP_424J2_126_3477_n1271), .A3(DP_OP_424J2_126_3477_n1273), .Y(
        DP_OP_424J2_126_3477_n1241) );
  NAND2X0_HVT U1623 ( .A1(DP_OP_423J2_125_3477_n876), .A2(
        DP_OP_423J2_125_3477_n878), .Y(n888) );
  AND2X1_HVT U1624 ( .A1(n1633), .A2(DP_OP_423J2_125_3477_n237), .Y(n890) );
  NAND3X0_HVT U1625 ( .A1(n1448), .A2(n1447), .A3(n1446), .Y(n891) );
  XOR3X2_HVT U1626 ( .A1(DP_OP_424J2_126_3477_n1218), .A2(
        DP_OP_424J2_126_3477_n1031), .A3(DP_OP_424J2_126_3477_n1029), .Y(
        DP_OP_424J2_126_3477_n1023) );
  NAND2X0_HVT U1627 ( .A1(DP_OP_424J2_126_3477_n1218), .A2(
        DP_OP_424J2_126_3477_n1029), .Y(n893) );
  NAND2X0_HVT U1628 ( .A1(DP_OP_424J2_126_3477_n1031), .A2(
        DP_OP_424J2_126_3477_n1029), .Y(n894) );
  NAND2X0_HVT U1629 ( .A1(DP_OP_424J2_126_3477_n1218), .A2(
        DP_OP_424J2_126_3477_n1031), .Y(n895) );
  NAND3X0_HVT U1630 ( .A1(n895), .A2(n894), .A3(n893), .Y(
        DP_OP_424J2_126_3477_n1022) );
  XOR3X2_HVT U1631 ( .A1(DP_OP_424J2_126_3477_n748), .A2(
        DP_OP_424J2_126_3477_n746), .A3(DP_OP_424J2_126_3477_n752), .Y(
        DP_OP_424J2_126_3477_n579) );
  NAND2X0_HVT U1632 ( .A1(DP_OP_424J2_126_3477_n748), .A2(
        DP_OP_424J2_126_3477_n752), .Y(n896) );
  NAND2X0_HVT U1633 ( .A1(DP_OP_424J2_126_3477_n746), .A2(
        DP_OP_424J2_126_3477_n752), .Y(n897) );
  NAND2X0_HVT U1634 ( .A1(DP_OP_424J2_126_3477_n746), .A2(
        DP_OP_424J2_126_3477_n748), .Y(n898) );
  NAND3X0_HVT U1635 ( .A1(n898), .A2(n897), .A3(n896), .Y(
        DP_OP_424J2_126_3477_n578) );
  XOR3X2_HVT U1636 ( .A1(DP_OP_425J2_127_3477_n374), .A2(
        DP_OP_425J2_127_3477_n376), .A3(DP_OP_425J2_127_3477_n353), .Y(
        DP_OP_425J2_127_3477_n351) );
  NAND2X0_HVT U1637 ( .A1(DP_OP_425J2_127_3477_n353), .A2(
        DP_OP_425J2_127_3477_n374), .Y(n899) );
  NAND2X0_HVT U1638 ( .A1(DP_OP_425J2_127_3477_n376), .A2(
        DP_OP_425J2_127_3477_n353), .Y(n9001) );
  NAND2X0_HVT U1639 ( .A1(DP_OP_425J2_127_3477_n376), .A2(
        DP_OP_425J2_127_3477_n374), .Y(n901) );
  NAND3X0_HVT U1640 ( .A1(n901), .A2(n9001), .A3(n899), .Y(
        DP_OP_425J2_127_3477_n350) );
  FADDX2_HVT U1641 ( .A(DP_OP_425J2_127_3477_n428), .B(
        DP_OP_425J2_127_3477_n381), .CI(DP_OP_425J2_127_3477_n426), .CO(
        DP_OP_425J2_127_3477_n376), .S(DP_OP_425J2_127_3477_n377) );
  NOR2X0_HVT U1642 ( .A1(DP_OP_422J2_124_3477_n2796), .A2(n876), .Y(
        DP_OP_424J2_126_3477_n2332) );
  XOR3X2_HVT U1643 ( .A1(DP_OP_423J2_125_3477_n423), .A2(
        DP_OP_423J2_125_3477_n514), .A3(n942), .Y(n1476) );
  XOR3X2_HVT U1644 ( .A1(DP_OP_425J2_127_3477_n1611), .A2(
        DP_OP_425J2_127_3477_n1742), .A3(DP_OP_425J2_127_3477_n1744), .Y(
        DP_OP_425J2_127_3477_n1591) );
  NAND2X0_HVT U1645 ( .A1(DP_OP_425J2_127_3477_n1611), .A2(
        DP_OP_425J2_127_3477_n1744), .Y(n902) );
  NAND2X0_HVT U1646 ( .A1(DP_OP_425J2_127_3477_n1742), .A2(
        DP_OP_425J2_127_3477_n1744), .Y(n903) );
  NAND2X0_HVT U1647 ( .A1(DP_OP_425J2_127_3477_n1742), .A2(
        DP_OP_425J2_127_3477_n1611), .Y(n904) );
  NAND3X0_HVT U1648 ( .A1(n904), .A2(n903), .A3(n902), .Y(
        DP_OP_425J2_127_3477_n1590) );
  HADDX2_HVT U1649 ( .A0(n1519), .B0(n1223), .SO(n_conv2_sum_c[8]) );
  OA21X2_HVT U1650 ( .A1(n1519), .A2(n1268), .A3(DP_OP_424J2_126_3477_n240), 
        .Y(n1269) );
  NAND2X0_HVT U1651 ( .A1(DP_OP_423J2_125_3477_n382), .A2(
        DP_OP_423J2_125_3477_n380), .Y(n905) );
  NAND2X0_HVT U1652 ( .A1(DP_OP_423J2_125_3477_n380), .A2(
        DP_OP_423J2_125_3477_n359), .Y(n906) );
  NAND2X0_HVT U1653 ( .A1(DP_OP_423J2_125_3477_n359), .A2(
        DP_OP_423J2_125_3477_n382), .Y(n907) );
  NAND3X0_HVT U1654 ( .A1(n907), .A2(n906), .A3(n905), .Y(
        DP_OP_423J2_125_3477_n354) );
  HADDX2_HVT U1655 ( .A0(DP_OP_423J2_125_3477_n253), .B0(n1084), .SO(
        n_conv2_sum_b[5]) );
  OR2X4_HVT U1656 ( .A1(DP_OP_424J2_126_3477_n2354), .A2(n876), .Y(
        DP_OP_424J2_126_3477_n2330) );
  NOR2X2_HVT U1657 ( .A1(DP_OP_424J2_126_3477_n2712), .A2(n874), .Y(
        DP_OP_425J2_127_3477_n2336) );
  NOR2X2_HVT U1658 ( .A1(DP_OP_425J2_127_3477_n2359), .A2(n876), .Y(
        DP_OP_425J2_127_3477_n2335) );
  NOR2X2_HVT U1659 ( .A1(DP_OP_425J2_127_3477_n2356), .A2(n874), .Y(
        DP_OP_425J2_127_3477_n2332) );
  NOR2X2_HVT U1660 ( .A1(DP_OP_425J2_127_3477_n2493), .A2(n875), .Y(
        DP_OP_422J2_124_3477_n2337) );
  XOR2X2_HVT U1661 ( .A1(n1385), .A2(n908), .Y(n_conv2_sum_a[15]) );
  IBUFFX32_HVT U1662 ( .A(DP_OP_422J2_124_3477_n22), .Y(n908) );
  NBUFFX2_HVT U1663 ( .A(DP_OP_423J2_125_3477_n340), .Y(n909) );
  HADDX2_HVT U1664 ( .A0(n1202), .B0(n1666), .SO(n_conv2_sum_b[7]) );
  XOR3X2_HVT U1665 ( .A1(DP_OP_425J2_127_3477_n1020), .A2(
        DP_OP_425J2_127_3477_n827), .A3(DP_OP_425J2_127_3477_n825), .Y(
        DP_OP_425J2_127_3477_n823) );
  NAND2X0_HVT U1666 ( .A1(DP_OP_425J2_127_3477_n1020), .A2(
        DP_OP_425J2_127_3477_n825), .Y(n910) );
  NAND2X0_HVT U1667 ( .A1(DP_OP_425J2_127_3477_n825), .A2(
        DP_OP_425J2_127_3477_n827), .Y(n911) );
  NAND2X0_HVT U1668 ( .A1(DP_OP_425J2_127_3477_n827), .A2(
        DP_OP_425J2_127_3477_n1020), .Y(n912) );
  NAND3X0_HVT U1669 ( .A1(n912), .A2(n911), .A3(n910), .Y(
        DP_OP_425J2_127_3477_n822) );
  HADDX2_HVT U1670 ( .A0(n1138), .B0(DP_OP_423J2_125_3477_n250), .SO(
        n_conv2_sum_b[6]) );
  NAND2X0_HVT U1671 ( .A1(n1535), .A2(DP_OP_422J2_124_3477_n244), .Y(n913) );
  AND2X4_HVT U1672 ( .A1(n1572), .A2(n1530), .Y(n914) );
  XOR3X2_HVT U1673 ( .A1(DP_OP_425J2_127_3477_n430), .A2(
        DP_OP_425J2_127_3477_n385), .A3(DP_OP_425J2_127_3477_n383), .Y(
        DP_OP_425J2_127_3477_n379) );
  NAND2X0_HVT U1674 ( .A1(DP_OP_425J2_127_3477_n430), .A2(
        DP_OP_425J2_127_3477_n383), .Y(n915) );
  NAND2X0_HVT U1675 ( .A1(DP_OP_425J2_127_3477_n385), .A2(
        DP_OP_425J2_127_3477_n383), .Y(n916) );
  NAND2X0_HVT U1676 ( .A1(DP_OP_425J2_127_3477_n385), .A2(
        DP_OP_425J2_127_3477_n430), .Y(n917) );
  NAND3X0_HVT U1677 ( .A1(n917), .A2(n916), .A3(n915), .Y(
        DP_OP_425J2_127_3477_n378) );
  XOR3X2_HVT U1678 ( .A1(DP_OP_425J2_127_3477_n2919), .A2(
        DP_OP_425J2_127_3477_n2025), .A3(DP_OP_425J2_127_3477_n2333), .Y(
        DP_OP_425J2_127_3477_n1181) );
  NAND2X0_HVT U1679 ( .A1(DP_OP_425J2_127_3477_n2919), .A2(
        DP_OP_425J2_127_3477_n2333), .Y(n918) );
  NAND2X0_HVT U1680 ( .A1(DP_OP_425J2_127_3477_n2025), .A2(
        DP_OP_425J2_127_3477_n2333), .Y(n919) );
  NAND2X1_HVT U1681 ( .A1(DP_OP_425J2_127_3477_n2025), .A2(
        DP_OP_425J2_127_3477_n2919), .Y(n920) );
  NAND3X0_HVT U1682 ( .A1(n920), .A2(n919), .A3(n918), .Y(
        DP_OP_425J2_127_3477_n1180) );
  NOR2X2_HVT U1683 ( .A1(DP_OP_425J2_127_3477_n2357), .A2(n874), .Y(
        DP_OP_425J2_127_3477_n2333) );
  NOR2X4_HVT U1684 ( .A1(DP_OP_422J2_124_3477_n3057), .A2(n444), .Y(
        DP_OP_425J2_127_3477_n2919) );
  IBUFFX2_HVT U1685 ( .A(DP_OP_423J2_125_3477_n19), .Y(n921) );
  NAND2X2_HVT U1686 ( .A1(DP_OP_423J2_125_3477_n283), .A2(
        DP_OP_423J2_125_3477_n167), .Y(DP_OP_423J2_125_3477_n19) );
  NAND3X0_HVT U1687 ( .A1(DP_OP_422J2_124_3477_n98), .A2(
        DP_OP_422J2_124_3477_n276), .A3(n1560), .Y(n922) );
  NAND2X0_HVT U1688 ( .A1(n923), .A2(n1559), .Y(n1177) );
  INVX1_HVT U1689 ( .A(n922), .Y(n923) );
  OA21X2_HVT U1690 ( .A1(DP_OP_422J2_124_3477_n102), .A2(
        DP_OP_422J2_124_3477_n110), .A3(DP_OP_422J2_124_3477_n105), .Y(n1560)
         );
  NAND3X0_HVT U1691 ( .A1(DP_OP_422J2_124_3477_n129), .A2(
        DP_OP_422J2_124_3477_n279), .A3(n1558), .Y(n924) );
  NAND2X0_HVT U1692 ( .A1(n925), .A2(n1557), .Y(n1088) );
  INVX1_HVT U1693 ( .A(n924), .Y(n925) );
  OA21X2_HVT U1694 ( .A1(DP_OP_422J2_124_3477_n133), .A2(
        DP_OP_422J2_124_3477_n141), .A3(DP_OP_422J2_124_3477_n136), .Y(n1558)
         );
  NAND3X0_HVT U1695 ( .A1(DP_OP_422J2_124_3477_n120), .A2(n1588), .A3(n1554), 
        .Y(n926) );
  NAND2X0_HVT U1696 ( .A1(n927), .A2(n1552), .Y(n1105) );
  INVX1_HVT U1697 ( .A(n926), .Y(n927) );
  OA21X2_HVT U1698 ( .A1(DP_OP_422J2_124_3477_n124), .A2(
        DP_OP_422J2_124_3477_n141), .A3(DP_OP_422J2_124_3477_n125), .Y(n1554)
         );
  AO22X2_HVT U1699 ( .A1(DP_OP_422J2_124_3477_n274), .A2(
        DP_OP_422J2_124_3477_n78), .A3(n1561), .A4(n1562), .Y(n1260) );
  AND2X1_HVT U1700 ( .A1(DP_OP_422J2_124_3477_n272), .A2(
        DP_OP_422J2_124_3477_n52), .Y(n928) );
  XOR3X2_HVT U1701 ( .A1(DP_OP_424J2_126_3477_n666), .A2(
        DP_OP_424J2_126_3477_n668), .A3(DP_OP_424J2_126_3477_n535), .Y(
        DP_OP_424J2_126_3477_n525) );
  NAND2X0_HVT U1702 ( .A1(n3), .A2(DP_OP_424J2_126_3477_n535), .Y(n929) );
  NAND2X0_HVT U1703 ( .A1(DP_OP_424J2_126_3477_n535), .A2(
        DP_OP_424J2_126_3477_n668), .Y(n930) );
  NAND2X0_HVT U1704 ( .A1(DP_OP_424J2_126_3477_n668), .A2(n3), .Y(n931) );
  NAND3X1_HVT U1705 ( .A1(n931), .A2(n930), .A3(n929), .Y(
        DP_OP_424J2_126_3477_n524) );
  XOR3X2_HVT U1706 ( .A1(DP_OP_424J2_126_3477_n430), .A2(
        DP_OP_424J2_126_3477_n385), .A3(DP_OP_424J2_126_3477_n383), .Y(
        DP_OP_424J2_126_3477_n379) );
  NAND2X0_HVT U1707 ( .A1(DP_OP_424J2_126_3477_n430), .A2(
        DP_OP_424J2_126_3477_n383), .Y(n932) );
  NAND2X0_HVT U1708 ( .A1(DP_OP_424J2_126_3477_n385), .A2(
        DP_OP_424J2_126_3477_n383), .Y(n933) );
  NAND2X0_HVT U1709 ( .A1(DP_OP_424J2_126_3477_n385), .A2(
        DP_OP_424J2_126_3477_n430), .Y(n934) );
  NAND3X0_HVT U1710 ( .A1(n934), .A2(n933), .A3(n932), .Y(
        DP_OP_424J2_126_3477_n378) );
  XOR3X2_HVT U1711 ( .A1(DP_OP_424J2_126_3477_n2919), .A2(
        DP_OP_424J2_126_3477_n2025), .A3(DP_OP_424J2_126_3477_n2333), .Y(
        DP_OP_424J2_126_3477_n1181) );
  NAND2X0_HVT U1712 ( .A1(DP_OP_424J2_126_3477_n2919), .A2(
        DP_OP_424J2_126_3477_n2333), .Y(n935) );
  NAND2X0_HVT U1713 ( .A1(DP_OP_424J2_126_3477_n2025), .A2(
        DP_OP_424J2_126_3477_n2333), .Y(n936) );
  NOR2X2_HVT U1714 ( .A1(DP_OP_422J2_124_3477_n2797), .A2(n876), .Y(
        DP_OP_424J2_126_3477_n2333) );
  NAND3X2_HVT U1715 ( .A1(DP_OP_422J2_124_3477_n105), .A2(
        DP_OP_422J2_124_3477_n277), .A3(DP_OP_422J2_124_3477_n110), .Y(n937)
         );
  NAND2X0_HVT U1716 ( .A1(n938), .A2(n1581), .Y(n1144) );
  INVX1_HVT U1717 ( .A(n937), .Y(n938) );
  NAND2X0_HVT U1718 ( .A1(DP_OP_425J2_127_3477_n1581), .A2(
        DP_OP_425J2_127_3477_n1730), .Y(n939) );
  NAND2X0_HVT U1719 ( .A1(DP_OP_425J2_127_3477_n1583), .A2(
        DP_OP_425J2_127_3477_n1730), .Y(n940) );
  NAND2X0_HVT U1720 ( .A1(DP_OP_425J2_127_3477_n1583), .A2(
        DP_OP_425J2_127_3477_n1581), .Y(n941) );
  NAND3X0_HVT U1721 ( .A1(n941), .A2(n940), .A3(n939), .Y(
        DP_OP_425J2_127_3477_n1576) );
  OR2X2_HVT U1722 ( .A1(DP_OP_424J2_126_3477_n418), .A2(
        DP_OP_424J2_126_3477_n373), .Y(n1711) );
  NBUFFX2_HVT U1723 ( .A(DP_OP_423J2_125_3477_n421), .Y(n942) );
  INVX1_HVT U1724 ( .A(DP_OP_422J2_124_3477_n351), .Y(n1572) );
  XOR2X2_HVT U1725 ( .A1(n1569), .A2(n943), .Y(n_conv2_sum_a[31]) );
  AND2X1_HVT U1726 ( .A1(n1583), .A2(DP_OP_422J2_124_3477_n38), .Y(n943) );
  XOR2X2_HVT U1727 ( .A1(n1567), .A2(n944), .Y(n_conv2_sum_a[30]) );
  AND2X1_HVT U1728 ( .A1(n1585), .A2(DP_OP_422J2_124_3477_n47), .Y(n944) );
  AND2X1_HVT U1729 ( .A1(n1586), .A2(DP_OP_422J2_124_3477_n65), .Y(n945) );
  XOR2X2_HVT U1730 ( .A1(n1566), .A2(n946), .Y(n_conv2_sum_a[21]) );
  AND2X1_HVT U1731 ( .A1(DP_OP_422J2_124_3477_n280), .A2(
        DP_OP_422J2_124_3477_n136), .Y(n946) );
  XOR2X2_HVT U1732 ( .A1(n1521), .A2(n947), .Y(n_conv2_sum_a[20]) );
  AND2X1_HVT U1733 ( .A1(DP_OP_422J2_124_3477_n281), .A2(
        DP_OP_422J2_124_3477_n149), .Y(n947) );
  XOR2X2_HVT U1734 ( .A1(n1564), .A2(n948), .Y(n_conv2_sum_a[19]) );
  AND2X1_HVT U1735 ( .A1(DP_OP_422J2_124_3477_n282), .A2(
        DP_OP_422J2_124_3477_n156), .Y(n948) );
  XOR2X2_HVT U1736 ( .A1(n1568), .A2(n949), .Y(n_conv2_sum_a[18]) );
  AND2X1_HVT U1737 ( .A1(DP_OP_422J2_124_3477_n283), .A2(
        DP_OP_422J2_124_3477_n167), .Y(n949) );
  XOR2X2_HVT U1738 ( .A1(n1565), .A2(n950), .Y(n_conv2_sum_a[17]) );
  AND2X1_HVT U1739 ( .A1(DP_OP_422J2_124_3477_n284), .A2(
        DP_OP_422J2_124_3477_n174), .Y(n950) );
  MUX21X1_HVT U1740 ( .A1(conv2_sram_rdata_weight[22]), .A2(
        conv1_sram_rdata_weight[22]), .S0(n619), .Y(conv_weight_box[14]) );
  AOI22X2_HVT U1741 ( .A1(n619), .A2(conv1_sram_rdata_weight[55]), .A3(n1095), 
        .A4(conv2_sram_rdata_weight[55]), .Y(DP_OP_424J2_126_3477_n2274) );
  MUX21X1_HVT U1742 ( .A1(conv2_sram_rdata_weight[66]), .A2(
        conv1_sram_rdata_weight[66]), .S0(n241), .Y(conv_weight_box[45]) );
  MUX21X1_HVT U1743 ( .A1(conv2_sram_rdata_weight[85]), .A2(
        conv1_sram_rdata_weight[85]), .S0(n241), .Y(conv_weight_box[58]) );
  AND2X4_HVT U1744 ( .A1(conv_weight_box[12]), .A2(src_window[91]), .Y(
        DP_OP_422J2_124_3477_n2950) );
  AND2X4_HVT U1745 ( .A1(conv_weight_box[12]), .A2(src_window[93]), .Y(
        DP_OP_422J2_124_3477_n2948) );
  AND2X4_HVT U1746 ( .A1(conv_weight_box[12]), .A2(src_window[89]), .Y(
        DP_OP_422J2_124_3477_n2952) );
  AND2X4_HVT U1747 ( .A1(conv_weight_box[12]), .A2(src_window[92]), .Y(
        DP_OP_422J2_124_3477_n2949) );
  AND2X4_HVT U1748 ( .A1(conv_weight_box[12]), .A2(src_window[88]), .Y(
        DP_OP_422J2_124_3477_n2953) );
  AND2X4_HVT U1749 ( .A1(conv_weight_box[12]), .A2(src_window[94]), .Y(
        DP_OP_422J2_124_3477_n2947) );
  XOR2X2_HVT U1750 ( .A1(n1563), .A2(n953), .Y(n_conv2_sum_a[16]) );
  AND2X1_HVT U1751 ( .A1(DP_OP_422J2_124_3477_n285), .A2(
        DP_OP_422J2_124_3477_n185), .Y(n953) );
  NAND3X1_HVT U1752 ( .A1(n1692), .A2(n1693), .A3(n1694), .Y(
        DP_OP_423J2_125_3477_n518) );
  XOR3X2_HVT U1753 ( .A1(DP_OP_425J2_127_3477_n650), .A2(
        DP_OP_425J2_127_3477_n517), .A3(DP_OP_425J2_127_3477_n515), .Y(
        DP_OP_425J2_127_3477_n513) );
  NAND2X0_HVT U1754 ( .A1(DP_OP_425J2_127_3477_n650), .A2(
        DP_OP_425J2_127_3477_n515), .Y(n954) );
  NAND2X0_HVT U1755 ( .A1(DP_OP_425J2_127_3477_n517), .A2(
        DP_OP_425J2_127_3477_n515), .Y(n955) );
  NAND2X0_HVT U1756 ( .A1(DP_OP_425J2_127_3477_n517), .A2(
        DP_OP_425J2_127_3477_n650), .Y(n956) );
  NAND3X0_HVT U1757 ( .A1(n956), .A2(n955), .A3(n954), .Y(
        DP_OP_425J2_127_3477_n512) );
  XOR3X2_HVT U1758 ( .A1(DP_OP_425J2_127_3477_n1028), .A2(
        DP_OP_425J2_127_3477_n837), .A3(DP_OP_425J2_127_3477_n1026), .Y(
        DP_OP_425J2_127_3477_n829) );
  NAND2X0_HVT U1759 ( .A1(DP_OP_425J2_127_3477_n1028), .A2(
        DP_OP_425J2_127_3477_n1026), .Y(n957) );
  NAND2X0_HVT U1760 ( .A1(DP_OP_425J2_127_3477_n1026), .A2(
        DP_OP_425J2_127_3477_n837), .Y(n958) );
  NAND2X0_HVT U1761 ( .A1(DP_OP_425J2_127_3477_n837), .A2(
        DP_OP_425J2_127_3477_n1028), .Y(n959) );
  NAND3X0_HVT U1762 ( .A1(n959), .A2(n958), .A3(n957), .Y(
        DP_OP_425J2_127_3477_n828) );
  OR2X4_HVT U1763 ( .A1(DP_OP_425J2_127_3477_n512), .A2(
        DP_OP_425J2_127_3477_n419), .Y(n1791) );
  INVX4_HVT U1764 ( .A(n1353), .Y(n1832) );
  INVX2_HVT U1765 ( .A(n1781), .Y(n1823) );
  INVX2_HVT U1766 ( .A(n488), .Y(n2174) );
  INVX4_HVT U1767 ( .A(n1928), .Y(n1418) );
  NOR2X4_HVT U1768 ( .A1(DP_OP_422J2_124_3477_n2358), .A2(n875), .Y(
        DP_OP_422J2_124_3477_n2334) );
  NOR2X4_HVT U1769 ( .A1(DP_OP_425J2_127_3477_n2358), .A2(n874), .Y(
        DP_OP_425J2_127_3477_n2334) );
  NOR2X4_HVT U1770 ( .A1(DP_OP_422J2_124_3477_n2357), .A2(n876), .Y(
        DP_OP_422J2_124_3477_n2333) );
  NOR2X4_HVT U1771 ( .A1(DP_OP_424J2_126_3477_n2358), .A2(n874), .Y(
        DP_OP_424J2_126_3477_n2334) );
  XOR3X2_HVT U1772 ( .A1(DP_OP_422J2_124_3477_n650), .A2(
        DP_OP_422J2_124_3477_n517), .A3(DP_OP_422J2_124_3477_n515), .Y(
        DP_OP_422J2_124_3477_n513) );
  NAND2X0_HVT U1773 ( .A1(DP_OP_422J2_124_3477_n515), .A2(
        DP_OP_422J2_124_3477_n650), .Y(n960) );
  NAND2X0_HVT U1774 ( .A1(DP_OP_422J2_124_3477_n517), .A2(
        DP_OP_422J2_124_3477_n515), .Y(n961) );
  NAND2X0_HVT U1775 ( .A1(DP_OP_422J2_124_3477_n517), .A2(
        DP_OP_422J2_124_3477_n650), .Y(n962) );
  NAND3X0_HVT U1776 ( .A1(n962), .A2(n961), .A3(n960), .Y(
        DP_OP_422J2_124_3477_n512) );
  XOR3X2_HVT U1777 ( .A1(DP_OP_422J2_124_3477_n1433), .A2(
        DP_OP_422J2_124_3477_n1592), .A3(DP_OP_422J2_124_3477_n1590), .Y(
        DP_OP_422J2_124_3477_n1415) );
  NAND2X0_HVT U1778 ( .A1(DP_OP_422J2_124_3477_n1433), .A2(
        DP_OP_422J2_124_3477_n1590), .Y(n963) );
  NAND2X0_HVT U1779 ( .A1(DP_OP_422J2_124_3477_n1592), .A2(
        DP_OP_422J2_124_3477_n1590), .Y(n964) );
  NAND2X0_HVT U1780 ( .A1(DP_OP_422J2_124_3477_n1592), .A2(
        DP_OP_422J2_124_3477_n1433), .Y(n965) );
  NAND3X0_HVT U1781 ( .A1(n965), .A2(n964), .A3(n963), .Y(
        DP_OP_422J2_124_3477_n1414) );
  OR2X4_HVT U1782 ( .A1(DP_OP_423J2_125_3477_n2354), .A2(n875), .Y(
        DP_OP_423J2_125_3477_n2330) );
  OR2X4_HVT U1783 ( .A1(DP_OP_422J2_124_3477_n2222), .A2(n874), .Y(
        DP_OP_425J2_127_3477_n2330) );
  NOR2X2_HVT U1784 ( .A1(DP_OP_422J2_124_3477_n2800), .A2(n875), .Y(
        DP_OP_424J2_126_3477_n2336) );
  NOR2X2_HVT U1785 ( .A1(DP_OP_423J2_125_3477_n2668), .A2(n875), .Y(
        DP_OP_422J2_124_3477_n2336) );
  NOR2X2_HVT U1786 ( .A1(DP_OP_424J2_126_3477_n2447), .A2(n875), .Y(
        DP_OP_423J2_125_3477_n2335) );
  OR2X4_HVT U1787 ( .A1(DP_OP_422J2_124_3477_n2354), .A2(n876), .Y(
        DP_OP_422J2_124_3477_n2330) );
  NOR2X2_HVT U1788 ( .A1(DP_OP_425J2_127_3477_n2580), .A2(n875), .Y(
        DP_OP_423J2_125_3477_n2336) );
  OR2X2_HVT U1789 ( .A1(DP_OP_422J2_124_3477_n418), .A2(
        DP_OP_422J2_124_3477_n373), .Y(n1534) );
  INVX1_HVT U1790 ( .A(conv2_sram_rdata_weight[99]), .Y(n1365) );
  INVX1_HVT U1791 ( .A(conv_weight_box[35]), .Y(n1443) );
  NOR2X0_HVT U1792 ( .A1(DP_OP_423J2_125_3477_n2537), .A2(
        DP_OP_425J2_127_3477_n2539), .Y(DP_OP_423J2_125_3477_n2513) );
  NOR2X0_HVT U1793 ( .A1(DP_OP_423J2_125_3477_n2536), .A2(
        DP_OP_424J2_126_3477_n2540), .Y(DP_OP_423J2_125_3477_n2520) );
  INVX1_HVT U1794 ( .A(n1362), .Y(n1364) );
  INVX1_HVT U1795 ( .A(n1379), .Y(DP_OP_422J2_124_3477_n1929) );
  NOR2X0_HVT U1796 ( .A1(DP_OP_422J2_124_3477_n3015), .A2(n704), .Y(
        DP_OP_422J2_124_3477_n2999) );
  OR2X1_HVT U1797 ( .A1(DP_OP_425J2_127_3477_n2797), .A2(
        DP_OP_423J2_125_3477_n2802), .Y(DP_OP_425J2_127_3477_n2765) );
  OR2X1_HVT U1798 ( .A1(DP_OP_423J2_125_3477_n2090), .A2(
        DP_OP_423J2_125_3477_n2849), .Y(DP_OP_425J2_127_3477_n2830) );
  OR2X1_HVT U1799 ( .A1(DP_OP_422J2_124_3477_n2662), .A2(
        DP_OP_425J2_127_3477_n2541), .Y(DP_OP_425J2_127_3477_n2522) );
  OR2X1_HVT U1800 ( .A1(DP_OP_425J2_127_3477_n2269), .A2(
        DP_OP_424J2_126_3477_n2802), .Y(DP_OP_424J2_126_3477_n2765) );
  OR2X1_HVT U1801 ( .A1(DP_OP_424J2_126_3477_n2796), .A2(n1443), .Y(
        DP_OP_424J2_126_3477_n2764) );
  OR2X1_HVT U1802 ( .A1(DP_OP_423J2_125_3477_n2799), .A2(
        DP_OP_423J2_125_3477_n2802), .Y(DP_OP_423J2_125_3477_n2767) );
  OR2X1_HVT U1803 ( .A1(DP_OP_423J2_125_3477_n2798), .A2(
        DP_OP_424J2_126_3477_n2802), .Y(DP_OP_423J2_125_3477_n2766) );
  NOR2X0_HVT U1804 ( .A1(DP_OP_425J2_127_3477_n2312), .A2(
        DP_OP_424J2_126_3477_n2849), .Y(DP_OP_423J2_125_3477_n2832) );
  OR2X1_HVT U1805 ( .A1(DP_OP_425J2_127_3477_n2310), .A2(
        DP_OP_423J2_125_3477_n2849), .Y(DP_OP_423J2_125_3477_n2830) );
  OR2X1_HVT U1806 ( .A1(DP_OP_425J2_127_3477_n2357), .A2(n1443), .Y(
        DP_OP_423J2_125_3477_n2765) );
  AND2X1_HVT U1807 ( .A1(n1372), .A2(src_window[270]), .Y(
        DP_OP_423J2_125_3477_n2463) );
  OR2X1_HVT U1808 ( .A1(DP_OP_425J2_127_3477_n2356), .A2(
        DP_OP_424J2_126_3477_n2802), .Y(DP_OP_423J2_125_3477_n2764) );
  OR2X1_HVT U1809 ( .A1(DP_OP_422J2_124_3477_n2574), .A2(
        DP_OP_425J2_127_3477_n2495), .Y(DP_OP_423J2_125_3477_n2462) );
  OR2X1_HVT U1810 ( .A1(DP_OP_423J2_125_3477_n2795), .A2(
        DP_OP_424J2_126_3477_n2802), .Y(DP_OP_423J2_125_3477_n2763) );
  OR2X1_HVT U1811 ( .A1(DP_OP_422J2_124_3477_n2799), .A2(n1443), .Y(
        DP_OP_422J2_124_3477_n2767) );
  OR2X1_HVT U1812 ( .A1(DP_OP_422J2_124_3477_n2535), .A2(n1362), .Y(
        DP_OP_422J2_124_3477_n2503) );
  OR2X1_HVT U1813 ( .A1(DP_OP_422J2_124_3477_n2798), .A2(
        DP_OP_423J2_125_3477_n2802), .Y(DP_OP_422J2_124_3477_n2766) );
  XOR3X1_HVT U1814 ( .A1(DP_OP_422J2_124_3477_n2156), .A2(
        DP_OP_422J2_124_3477_n2163), .A3(DP_OP_422J2_124_3477_n2860), .Y(
        DP_OP_422J2_124_3477_n971) );
  NOR2X0_HVT U1815 ( .A1(DP_OP_423J2_125_3477_n2048), .A2(n704), .Y(
        DP_OP_422J2_124_3477_n3000) );
  OR2X1_HVT U1816 ( .A1(DP_OP_422J2_124_3477_n2662), .A2(
        DP_OP_424J2_126_3477_n2671), .Y(DP_OP_422J2_124_3477_n2638) );
  OR2X1_HVT U1817 ( .A1(DP_OP_425J2_127_3477_n2798), .A2(
        DP_OP_424J2_126_3477_n2802), .Y(DP_OP_425J2_127_3477_n2766) );
  NOR2X0_HVT U1818 ( .A1(DP_OP_423J2_125_3477_n2666), .A2(
        DP_OP_425J2_127_3477_n2495), .Y(DP_OP_425J2_127_3477_n2466) );
  NOR2X0_HVT U1819 ( .A1(DP_OP_423J2_125_3477_n2399), .A2(
        DP_OP_425J2_127_3477_n2541), .Y(DP_OP_425J2_127_3477_n2523) );
  NOR2X0_HVT U1820 ( .A1(DP_OP_423J2_125_3477_n2665), .A2(
        DP_OP_425J2_127_3477_n2495), .Y(DP_OP_425J2_127_3477_n2465) );
  NOR2X0_HVT U1821 ( .A1(DP_OP_422J2_124_3477_n2796), .A2(
        DP_OP_424J2_126_3477_n2671), .Y(DP_OP_425J2_127_3477_n2640) );
  NOR2X0_HVT U1822 ( .A1(DP_OP_424J2_126_3477_n2576), .A2(
        DP_OP_425J2_127_3477_n2495), .Y(DP_OP_425J2_127_3477_n2464) );
  NOR2X0_HVT U1823 ( .A1(DP_OP_424J2_126_3477_n2575), .A2(
        DP_OP_425J2_127_3477_n2495), .Y(DP_OP_425J2_127_3477_n2463) );
  OR2X1_HVT U1824 ( .A1(DP_OP_424J2_126_3477_n2354), .A2(
        DP_OP_424J2_126_3477_n2671), .Y(DP_OP_425J2_127_3477_n2638) );
  OR2X1_HVT U1825 ( .A1(DP_OP_424J2_126_3477_n2574), .A2(
        DP_OP_425J2_127_3477_n2495), .Y(DP_OP_425J2_127_3477_n2462) );
  OR2X1_HVT U1826 ( .A1(DP_OP_423J2_125_3477_n2135), .A2(
        DP_OP_423J2_125_3477_n2802), .Y(DP_OP_425J2_127_3477_n2763) );
  OR2X1_HVT U1827 ( .A1(DP_OP_424J2_126_3477_n2799), .A2(
        DP_OP_424J2_126_3477_n2802), .Y(DP_OP_424J2_126_3477_n2767) );
  OR2X1_HVT U1828 ( .A1(DP_OP_423J2_125_3477_n2886), .A2(
        DP_OP_424J2_126_3477_n2802), .Y(DP_OP_424J2_126_3477_n2766) );
  NOR2X0_HVT U1829 ( .A1(DP_OP_425J2_127_3477_n2401), .A2(
        DP_OP_424J2_126_3477_n2671), .Y(DP_OP_424J2_126_3477_n2641) );
  OR2X1_HVT U1830 ( .A1(DP_OP_424J2_126_3477_n2795), .A2(n1443), .Y(
        DP_OP_424J2_126_3477_n2763) );
  OR2X1_HVT U1831 ( .A1(DP_OP_423J2_125_3477_n2800), .A2(n1443), .Y(
        DP_OP_423J2_125_3477_n2768) );
  NOR2X0_HVT U1832 ( .A1(DP_OP_423J2_125_3477_n2794), .A2(
        DP_OP_424J2_126_3477_n2802), .Y(DP_OP_423J2_125_3477_n2762) );
  INVX1_HVT U1833 ( .A(conv_weight_box[45]), .Y(n1497) );
  INVX1_HVT U1834 ( .A(conv_weight_box[17]), .Y(DP_OP_422J2_124_3477_n2935) );
  NOR2X0_HVT U1835 ( .A1(DP_OP_422J2_124_3477_n2841), .A2(
        DP_OP_424J2_126_3477_n2849), .Y(DP_OP_422J2_124_3477_n2833) );
  NOR2X0_HVT U1836 ( .A1(DP_OP_425J2_127_3477_n2886), .A2(n704), .Y(
        DP_OP_422J2_124_3477_n3002) );
  INVX1_HVT U1837 ( .A(conv_weight_box[64]), .Y(DP_OP_422J2_124_3477_n2495) );
  OR2X1_HVT U1838 ( .A1(DP_OP_422J2_124_3477_n2537), .A2(n1336), .Y(
        DP_OP_422J2_124_3477_n2505) );
  NOR2X0_HVT U1839 ( .A1(DP_OP_422J2_124_3477_n2667), .A2(
        DP_OP_424J2_126_3477_n2671), .Y(DP_OP_422J2_124_3477_n2643) );
  NOR2X0_HVT U1840 ( .A1(DP_OP_422J2_124_3477_n2840), .A2(n1428), .Y(
        DP_OP_422J2_124_3477_n2832) );
  NOR2X0_HVT U1841 ( .A1(DP_OP_422J2_124_3477_n3017), .A2(n703), .Y(
        DP_OP_422J2_124_3477_n3001) );
  OR2X1_HVT U1842 ( .A1(DP_OP_422J2_124_3477_n3014), .A2(n704), .Y(
        DP_OP_422J2_124_3477_n2998) );
  OR2X1_HVT U1843 ( .A1(DP_OP_422J2_124_3477_n2796), .A2(n1443), .Y(
        DP_OP_422J2_124_3477_n2764) );
  NOR2X0_HVT U1844 ( .A1(DP_OP_422J2_124_3477_n2754), .A2(
        DP_OP_422J2_124_3477_n2759), .Y(DP_OP_422J2_124_3477_n2730) );
  NOR2X0_HVT U1845 ( .A1(DP_OP_424J2_126_3477_n2579), .A2(
        DP_OP_425J2_127_3477_n2495), .Y(DP_OP_425J2_127_3477_n2467) );
  OR2X1_HVT U1846 ( .A1(DP_OP_425J2_127_3477_n2800), .A2(
        DP_OP_423J2_125_3477_n2802), .Y(DP_OP_425J2_127_3477_n2768) );
  NOR2X0_HVT U1847 ( .A1(DP_OP_424J2_126_3477_n2222), .A2(n1443), .Y(
        DP_OP_425J2_127_3477_n2762) );
  AND2X1_HVT U1848 ( .A1(n1366), .A2(src_window[199]), .Y(
        DP_OP_425J2_127_3477_n2586) );
  INVX1_HVT U1849 ( .A(conv2_sram_rdata_weight[77]), .Y(n1356) );
  OR2X1_HVT U1850 ( .A1(DP_OP_422J2_124_3477_n2140), .A2(n1443), .Y(
        DP_OP_424J2_126_3477_n2768) );
  NOR2X0_HVT U1851 ( .A1(DP_OP_424J2_126_3477_n2667), .A2(
        DP_OP_424J2_126_3477_n2671), .Y(DP_OP_424J2_126_3477_n2643) );
  NOR2X0_HVT U1852 ( .A1(DP_OP_424J2_126_3477_n2794), .A2(
        DP_OP_423J2_125_3477_n2802), .Y(DP_OP_424J2_126_3477_n2762) );
  INVX1_HVT U1853 ( .A(n1720), .Y(n1373) );
  INVX1_HVT U1854 ( .A(conv_weight_box[17]), .Y(DP_OP_425J2_127_3477_n2935) );
  INVX1_HVT U1855 ( .A(conv_weight_box[20]), .Y(DP_OP_422J2_124_3477_n2143) );
  NOR2X0_HVT U1856 ( .A1(DP_OP_422J2_124_3477_n3019), .A2(n704), .Y(
        DP_OP_422J2_124_3477_n3003) );
  NOR2X0_HVT U1857 ( .A1(DP_OP_425J2_127_3477_n2493), .A2(
        DP_OP_425J2_127_3477_n2495), .Y(DP_OP_425J2_127_3477_n2469) );
  INVX1_HVT U1858 ( .A(conv_weight_box[20]), .Y(DP_OP_425J2_127_3477_n2143) );
  INVX1_HVT U1859 ( .A(conv_weight_box[50]), .Y(DP_OP_424J2_126_3477_n2671) );
  INVX1_HVT U1860 ( .A(n1779), .Y(n1377) );
  NOR2X0_HVT U1861 ( .A1(DP_OP_424J2_126_3477_n2580), .A2(
        DP_OP_425J2_127_3477_n2495), .Y(DP_OP_425J2_127_3477_n2468) );
  NOR2X0_HVT U1862 ( .A1(DP_OP_422J2_124_3477_n3019), .A2(
        DP_OP_423J2_125_3477_n2892), .Y(DP_OP_425J2_127_3477_n2871) );
  NOR2X0_HVT U1863 ( .A1(DP_OP_425J2_127_3477_n2534), .A2(
        DP_OP_425J2_127_3477_n2541), .Y(DP_OP_425J2_127_3477_n2526) );
  XOR3X1_HVT U1864 ( .A1(n1646), .A2(n1647), .A3(n1648), .Y(
        DP_OP_423J2_125_3477_n1803) );
  XOR3X1_HVT U1865 ( .A1(n1640), .A2(n1641), .A3(n1642), .Y(
        DP_OP_423J2_125_3477_n1715) );
  NOR2X0_HVT U1866 ( .A1(DP_OP_424J2_126_3477_n2184), .A2(
        DP_OP_422J2_124_3477_n2980), .Y(DP_OP_422J2_124_3477_n2960) );
  INVX4_HVT U1867 ( .A(n1531), .Y(n1532) );
  NOR2X0_HVT U1868 ( .A1(DP_OP_425J2_127_3477_n2536), .A2(
        DP_OP_425J2_127_3477_n2541), .Y(DP_OP_425J2_127_3477_n2528) );
  NOR2X0_HVT U1869 ( .A1(DP_OP_422J2_124_3477_n3021), .A2(n704), .Y(
        DP_OP_422J2_124_3477_n3005) );
  MUX21X1_HVT U1870 ( .A1(conv2_sram_rdata_weight[76]), .A2(
        conv1_sram_rdata_weight[76]), .S0(n241), .Y(conv_weight_box[51]) );
  NAND3X0_HVT U1871 ( .A1(n1468), .A2(n1469), .A3(n1470), .Y(
        DP_OP_423J2_125_3477_n1414) );
  NOR2X0_HVT U1872 ( .A1(DP_OP_423J2_125_3477_n2845), .A2(n1428), .Y(
        DP_OP_423J2_125_3477_n2837) );
  NOR2X0_HVT U1873 ( .A1(DP_OP_424J2_126_3477_n2317), .A2(
        DP_OP_424J2_126_3477_n2849), .Y(DP_OP_422J2_124_3477_n2837) );
  NOR2X0_HVT U1874 ( .A1(DP_OP_423J2_125_3477_n2097), .A2(n1428), .Y(
        DP_OP_425J2_127_3477_n2837) );
  AND2X1_HVT U1875 ( .A1(n1395), .A2(src_window[104]), .Y(
        DP_OP_425J2_127_3477_n2221) );
  INVX1_HVT U1876 ( .A(n1686), .Y(DP_OP_423J2_125_3477_n240) );
  OR2X1_HVT U1877 ( .A1(DP_OP_422J2_124_3477_n648), .A2(
        DP_OP_422J2_124_3477_n513), .Y(n1536) );
  OR2X1_HVT U1878 ( .A1(DP_OP_425J2_127_3477_n372), .A2(
        DP_OP_425J2_127_3477_n351), .Y(n1814) );
  OA21X1_HVT U1879 ( .A1(n1811), .A2(n1806), .A3(n1812), .Y(
        DP_OP_425J2_127_3477_n110) );
  OA21X1_HVT U1880 ( .A1(DP_OP_424J2_126_3477_n182), .A2(
        DP_OP_424J2_126_3477_n190), .A3(DP_OP_424J2_126_3477_n185), .Y(n1740)
         );
  OA21X1_HVT U1881 ( .A1(DP_OP_424J2_126_3477_n82), .A2(
        DP_OP_424J2_126_3477_n110), .A3(DP_OP_424J2_126_3477_n85), .Y(n1352)
         );
  AO22X1_HVT U1882 ( .A1(n1833), .A2(DP_OP_425J2_127_3477_n38), .A3(n1793), 
        .A4(n1847), .Y(n1147) );
  OA22X1_HVT U1883 ( .A1(n2067), .A2(conv2_sum_d[16]), .A3(n1906), .A4(
        conv2_sum_d[17]), .Y(n966) );
  OA222X1_HVT U1884 ( .A1(conv2_sum_d[18]), .A2(n2066), .A3(conv2_sum_d[19]), 
        .A4(n1907), .A5(n2099), .A6(n966), .Y(n967) );
  NAND2X0_HVT U1885 ( .A1(n2068), .A2(conv2_sum_c[22]), .Y(n968) );
  OA22X1_HVT U1886 ( .A1(n2062), .A2(conv2_sum_d[20]), .A3(n1908), .A4(
        conv2_sum_d[21]), .Y(n969) );
  OA222X1_HVT U1887 ( .A1(n968), .A2(conv2_sum_d[22]), .A3(conv2_sum_d[23]), 
        .A4(n1909), .A5(n2069), .A6(n969), .Y(n970) );
  OA21X1_HVT U1888 ( .A1(n2098), .A2(n967), .A3(n970), .Y(n1920) );
  NAND3X0_HVT U1889 ( .A1(tmp_big1[1]), .A2(n2176), .A3(n2175), .Y(n971) );
  NAND2X0_HVT U1890 ( .A1(n971), .A2(tmp_big2[0]), .Y(n2140) );
  INVX0_HVT U1891 ( .A(DP_OP_425J2_127_3477_n140), .Y(n972) );
  NAND2X0_HVT U1892 ( .A1(n1832), .A2(n972), .Y(n1809) );
  INVX0_HVT U1893 ( .A(tmp_big2[8]), .Y(n973) );
  INVX0_HVT U1894 ( .A(n2137), .Y(n974) );
  NAND2X0_HVT U1897 ( .A1(DP_OP_425J2_127_3477_n146), .A2(
        DP_OP_425J2_127_3477_n165), .Y(n977) );
  AO22X2_HVT U1898 ( .A1(DP_OP_425J2_127_3477_n285), .A2(
        DP_OP_425J2_127_3477_n185), .A3(n1800), .A4(DP_OP_425J2_127_3477_n190), 
        .Y(n978) );
  NAND4X0_HVT U1899 ( .A1(DP_OP_425J2_127_3477_n285), .A2(
        DP_OP_425J2_127_3477_n185), .A3(n1800), .A4(DP_OP_425J2_127_3477_n190), 
        .Y(n979) );
  NAND2X0_HVT U1900 ( .A1(n979), .A2(n978), .Y(n_conv2_sum_d[16]) );
  OA22X1_HVT U1901 ( .A1(n1985), .A2(tmp_big2[3]), .A3(tmp_big2[2]), .A4(n2139), .Y(n980) );
  AOI22X1_HVT U1902 ( .A1(n1985), .A2(tmp_big2[3]), .A3(n2167), .A4(
        tmp_big2[2]), .Y(n981) );
  OA22X1_HVT U1903 ( .A1(n1401), .A2(tmp_big1[1]), .A3(tmp_big1[0]), .A4(n2140), .Y(n982) );
  NAND2X0_HVT U1904 ( .A1(n981), .A2(n982), .Y(n983) );
  AO22X1_HVT U1905 ( .A1(n1918), .A2(tmp_big2[4]), .A3(n2170), .A4(tmp_big2[5]), .Y(n984) );
  NAND3X0_HVT U1907 ( .A1(conv2_sum_a[24]), .A2(n2044), .A3(n1296), .Y(n986)
         );
  OA21X1_HVT U1908 ( .A1(conv2_sum_b[25]), .A2(n1903), .A3(n986), .Y(n2000) );
  AO22X2_HVT U1909 ( .A1(DP_OP_425J2_127_3477_n284), .A2(
        DP_OP_425J2_127_3477_n174), .A3(n1804), .A4(n1806), .Y(n987) );
  NAND4X0_HVT U1910 ( .A1(DP_OP_425J2_127_3477_n284), .A2(
        DP_OP_425J2_127_3477_n174), .A3(n1804), .A4(n1806), .Y(n988) );
  NAND2X0_HVT U1911 ( .A1(n987), .A2(n988), .Y(n_conv2_sum_d[17]) );
  INVX0_HVT U1912 ( .A(n2060), .Y(n989) );
  INVX0_HVT U1913 ( .A(n2061), .Y(n990) );
  NAND2X0_HVT U1914 ( .A1(conv2_sum_d[24]), .A2(n1895), .Y(n991) );
  AND4X1_HVT U1915 ( .A1(n2103), .A2(n989), .A3(n990), .A4(n991), .Y(n1964) );
  OAI21X1_HVT U1916 ( .A1(conv2_sum_a[8]), .A2(n1858), .A3(n2031), .Y(n992) );
  OR3X1_HVT U1917 ( .A1(n2032), .A2(n2033), .A3(n992), .Y(n993) );
  AO22X2_HVT U1918 ( .A1(DP_OP_425J2_127_3477_n282), .A2(
        DP_OP_425J2_127_3477_n156), .A3(n1808), .A4(n1822), .Y(n994) );
  NAND4X0_HVT U1919 ( .A1(DP_OP_425J2_127_3477_n282), .A2(
        DP_OP_425J2_127_3477_n156), .A3(n1808), .A4(n1822), .Y(n995) );
  NAND2X0_HVT U1920 ( .A1(n994), .A2(n995), .Y(n_conv2_sum_d[19]) );
  NAND2X0_HVT U1921 ( .A1(n1989), .A2(n887), .Y(n996) );
  NAND2X0_HVT U1922 ( .A1(tmp_big2[7]), .A2(n2171), .Y(n997) );
  NAND2X0_HVT U1923 ( .A1(tmp_big1[6]), .A2(n997), .Y(n998) );
  OA22X1_HVT U1924 ( .A1(tmp_big2[4]), .A2(n1918), .A3(tmp_big2[5]), .A4(n2170), .Y(n999) );
  AO21X1_HVT U1925 ( .A1(n2170), .A2(tmp_big2[5]), .A3(n999), .Y(n1000) );
  OA222X1_HVT U1926 ( .A1(n998), .A2(tmp_big2[6]), .A3(tmp_big2[7]), .A4(n2171), .A5(n1000), .A6(n2141), .Y(n1933) );
  NAND3X0_HVT U1927 ( .A1(n1724), .A2(n1723), .A3(n1001), .Y(n1725) );
  AO22X2_HVT U1928 ( .A1(DP_OP_425J2_127_3477_n280), .A2(
        DP_OP_425J2_127_3477_n136), .A3(n1809), .A4(DP_OP_425J2_127_3477_n141), 
        .Y(n1002) );
  NAND4X0_HVT U1929 ( .A1(DP_OP_425J2_127_3477_n280), .A2(
        DP_OP_425J2_127_3477_n136), .A3(n1809), .A4(DP_OP_425J2_127_3477_n141), 
        .Y(n1003) );
  NAND2X0_HVT U1930 ( .A1(n1002), .A2(n1003), .Y(n_conv2_sum_d[21]) );
  NAND2X0_HVT U1931 ( .A1(n2157), .A2(tmp_big2[15]), .Y(n1004) );
  NAND2X0_HVT U1932 ( .A1(tmp_big1[14]), .A2(n1004), .Y(n1005) );
  OA22X1_HVT U1933 ( .A1(n2157), .A2(tmp_big2[15]), .A3(tmp_big2[14]), .A4(
        n1005), .Y(n1936) );
  NAND2X0_HVT U1934 ( .A1(n2103), .A2(conv2_sum_c[24]), .Y(n1006) );
  OA22X1_HVT U1935 ( .A1(conv2_sum_d[25]), .A2(n1910), .A3(conv2_sum_d[24]), 
        .A4(n1006), .Y(n2053) );
  INVX0_HVT U1936 ( .A(n2009), .Y(n1007) );
  INVX0_HVT U1937 ( .A(n2008), .Y(n1008) );
  NAND2X0_HVT U1938 ( .A1(conv2_sum_b[24]), .A2(n1888), .Y(n1009) );
  NAND4X0_HVT U1939 ( .A1(n2044), .A2(n1007), .A3(n1008), .A4(n1009), .Y(n1966) );
  NAND2X0_HVT U1941 ( .A1(DP_OP_424J2_126_3477_n146), .A2(
        DP_OP_424J2_126_3477_n165), .Y(n1011) );
  AOI22X1_HVT U1943 ( .A1(n1759), .A2(DP_OP_424J2_126_3477_n72), .A3(
        DP_OP_424J2_126_3477_n201), .A4(DP_OP_424J2_126_3477_n58), .Y(n1013)
         );
  INVX0_HVT U1944 ( .A(DP_OP_423J2_125_3477_n267), .Y(n1014) );
  AND2X1_HVT U1945 ( .A1(n1014), .A2(DP_OP_423J2_125_3477_n268), .Y(n1015) );
  HADDX1_HVT U1946 ( .A0(n1015), .B0(DP_OP_423J2_125_3477_n269), .SO(
        n_conv2_sum_b[1]) );
  AO22X2_HVT U1947 ( .A1(n1842), .A2(DP_OP_425J2_127_3477_n120), .A3(n1805), 
        .A4(n1807), .Y(n1016) );
  NAND4X0_HVT U1948 ( .A1(n1842), .A2(DP_OP_425J2_127_3477_n120), .A3(n1805), 
        .A4(n1807), .Y(n1017) );
  NAND2X0_HVT U1949 ( .A1(n1016), .A2(n1017), .Y(n_conv2_sum_d[23]) );
  NAND2X0_HVT U1950 ( .A1(n1915), .A2(conv2_sum_c[31]), .Y(n1018) );
  NAND2X0_HVT U1951 ( .A1(conv2_sum_c[30]), .A2(n1018), .Y(n2055) );
  INVX0_HVT U1952 ( .A(n2117), .Y(n1019) );
  INVX0_HVT U1953 ( .A(n2118), .Y(n1020) );
  INVX0_HVT U1954 ( .A(tmp_big1[24]), .Y(n1021) );
  NAND2X0_HVT U1955 ( .A1(tmp_big2[24]), .A2(n1021), .Y(n1022) );
  NAND4X0_HVT U1956 ( .A1(n2148), .A2(n1019), .A3(n1020), .A4(n1022), .Y(n1971) );
  NAND2X0_HVT U1958 ( .A1(DP_OP_422J2_124_3477_n146), .A2(
        DP_OP_422J2_124_3477_n165), .Y(n1024) );
  OR2X1_HVT U1959 ( .A1(DP_OP_425J2_127_3477_n115), .A2(
        DP_OP_425J2_127_3477_n145), .Y(n1025) );
  NAND2X0_HVT U1960 ( .A1(n1842), .A2(DP_OP_425J2_127_3477_n127), .Y(n1026) );
  NAND3X0_HVT U1961 ( .A1(n1025), .A2(DP_OP_425J2_127_3477_n120), .A3(n1026), 
        .Y(DP_OP_425J2_127_3477_n114) );
  OR2X1_HVT U1962 ( .A1(DP_OP_424J2_126_3477_n115), .A2(
        DP_OP_424J2_126_3477_n145), .Y(n1027) );
  NAND2X0_HVT U1963 ( .A1(n1764), .A2(DP_OP_424J2_126_3477_n127), .Y(n1028) );
  NAND3X0_HVT U1964 ( .A1(n1027), .A2(DP_OP_424J2_126_3477_n120), .A3(n1028), 
        .Y(DP_OP_424J2_126_3477_n114) );
  INVX0_HVT U1965 ( .A(n490), .Y(n1029) );
  OA221X1_HVT U1966 ( .A1(n1029), .A2(n2042), .A3(n1029), .A4(n2043), .A5(
        n2045), .Y(n1533) );
  INVX0_HVT U1967 ( .A(n1823), .Y(n1030) );
  NAND3X0_HVT U1968 ( .A1(n1783), .A2(n1782), .A3(n1030), .Y(n1784) );
  AND2X1_HVT U1969 ( .A1(DP_OP_423J2_125_3477_n265), .A2(n1676), .Y(n1031) );
  HADDX1_HVT U1970 ( .A0(n1031), .B0(DP_OP_423J2_125_3477_n266), .SO(
        n_conv2_sum_b[2]) );
  NAND2X0_HVT U1971 ( .A1(n1032), .A2(n1033), .Y(n_conv2_sum_c[17]) );
  OA22X1_HVT U1972 ( .A1(tmp_big2[26]), .A2(n2163), .A3(tmp_big2[27]), .A4(
        n2164), .Y(n1034) );
  AO21X1_HVT U1973 ( .A1(n2164), .A2(tmp_big2[27]), .A3(n1034), .Y(n1924) );
  NAND2X0_HVT U1974 ( .A1(conv2_sum_b[5]), .A2(n1852), .Y(n1035) );
  NAND2X0_HVT U1975 ( .A1(conv2_sum_a[4]), .A2(n1035), .Y(n1036) );
  OA22X1_HVT U1976 ( .A1(conv2_sum_b[5]), .A2(n1852), .A3(conv2_sum_b[4]), 
        .A4(n1036), .Y(n2038) );
  OR2X1_HVT U1977 ( .A1(DP_OP_423J2_125_3477_n115), .A2(
        DP_OP_423J2_125_3477_n145), .Y(n1037) );
  NAND2X0_HVT U1978 ( .A1(n1673), .A2(DP_OP_423J2_125_3477_n127), .Y(n1038) );
  NAND3X0_HVT U1979 ( .A1(n1037), .A2(DP_OP_423J2_125_3477_n120), .A3(n1038), 
        .Y(DP_OP_423J2_125_3477_n114) );
  NOR3X0_HVT U1980 ( .A1(n2041), .A2(n2040), .A3(n1039), .Y(n1876) );
  AOI21X1_HVT U1981 ( .A1(DP_OP_423J2_125_3477_n177), .A2(
        DP_OP_423J2_125_3477_n162), .A3(DP_OP_423J2_125_3477_n165), .Y(
        DP_OP_423J2_125_3477_n161) );
  NAND2X0_HVT U1982 ( .A1(n1588), .A2(DP_OP_422J2_124_3477_n127), .Y(n1040) );
  OR2X1_HVT U1983 ( .A1(DP_OP_422J2_124_3477_n115), .A2(
        DP_OP_422J2_124_3477_n145), .Y(n1041) );
  NAND3X0_HVT U1984 ( .A1(n1041), .A2(DP_OP_422J2_124_3477_n120), .A3(n1040), 
        .Y(DP_OP_422J2_124_3477_n114) );
  AOI22X1_HVT U1986 ( .A1(n1836), .A2(DP_OP_425J2_127_3477_n72), .A3(
        DP_OP_425J2_127_3477_n201), .A4(DP_OP_425J2_127_3477_n58), .Y(n1044)
         );
  NAND3X0_HVT U1987 ( .A1(n1832), .A2(n1835), .A3(DP_OP_425J2_127_3477_n49), 
        .Y(n1793) );
  OAI21X1_HVT U1988 ( .A1(DP_OP_424J2_126_3477_n107), .A2(
        DP_OP_424J2_126_3477_n13), .A3(DP_OP_424J2_126_3477_n110), .Y(n1750)
         );
  INVX0_HVT U1989 ( .A(DP_OP_423J2_125_3477_n259), .Y(n1045) );
  NAND2X0_HVT U1990 ( .A1(n1045), .A2(DP_OP_423J2_125_3477_n260), .Y(n1046) );
  HADDX1_HVT U1991 ( .A0(DP_OP_423J2_125_3477_n261), .B0(n1046), .SO(
        n_conv2_sum_b[3]) );
  NAND2X0_HVT U1992 ( .A1(n1047), .A2(n1048), .Y(n_conv2_sum_c[16]) );
  NAND2X0_HVT U1993 ( .A1(n1049), .A2(n1050), .Y(n_conv2_sum_c[19]) );
  NAND2X0_HVT U1994 ( .A1(n2082), .A2(conv2_sum_c[8]), .Y(n1051) );
  OA22X1_HVT U1995 ( .A1(conv2_sum_d[9]), .A2(n1993), .A3(conv2_sum_d[8]), 
        .A4(n1051), .Y(n1052) );
  NAND2X0_HVT U1996 ( .A1(n2075), .A2(n1052), .Y(n1991) );
  INVX0_HVT U1997 ( .A(n2174), .Y(n1053) );
  AO22X1_HVT U1998 ( .A1(n2174), .A2(conv2_sum_b[11]), .A3(n1053), .A4(
        conv2_sum_a[11]), .Y(tmp_big1[11]) );
  INVX0_HVT U1999 ( .A(n490), .Y(n1054) );
  OA221X2_HVT U2000 ( .A1(n1054), .A2(n2043), .A3(n1054), .A4(n2042), .A5(
        n2045), .Y(n1960) );
  NAND2X0_HVT U2001 ( .A1(n1528), .A2(DP_OP_423J2_125_3477_n286), .Y(n1055) );
  AND2X1_HVT U2002 ( .A1(n1055), .A2(DP_OP_423J2_125_3477_n198), .Y(
        DP_OP_423J2_125_3477_n190) );
  NAND2X0_HVT U2003 ( .A1(DP_OP_422J2_124_3477_n96), .A2(n1587), .Y(n1056) );
  AND2X1_HVT U2004 ( .A1(n1056), .A2(DP_OP_422J2_124_3477_n89), .Y(
        DP_OP_422J2_124_3477_n85) );
  NAND2X0_HVT U2005 ( .A1(n1525), .A2(DP_OP_422J2_124_3477_n286), .Y(n1057) );
  AND2X1_HVT U2006 ( .A1(n1057), .A2(DP_OP_422J2_124_3477_n198), .Y(
        DP_OP_422J2_124_3477_n190) );
  IBUFFX2_HVT U2007 ( .A(DP_OP_424J2_126_3477_n160), .Y(n1058) );
  AO22X1_HVT U2008 ( .A1(n1531), .A2(conv2_sum_d[0]), .A3(n1994), .A4(
        conv2_sum_c[0]), .Y(tmp_big2[0]) );
  INVX0_HVT U2009 ( .A(DP_OP_423J2_125_3477_n256), .Y(n1059) );
  NAND2X0_HVT U2010 ( .A1(n1059), .A2(DP_OP_423J2_125_3477_n257), .Y(n1060) );
  HADDX1_HVT U2011 ( .A0(n1634), .B0(n1060), .SO(n_conv2_sum_b[4]) );
  AND2X1_HVT U2012 ( .A1(DP_OP_425J2_127_3477_n257), .A2(
        DP_OP_425J2_127_3477_n297), .Y(n1061) );
  HADDX1_HVT U2013 ( .A0(n1061), .B0(n1796), .SO(n_conv2_sum_d[4]) );
  AO22X2_HVT U2014 ( .A1(n1841), .A2(DP_OP_425J2_127_3477_n89), .A3(n1810), 
        .A4(n1813), .Y(n1062) );
  NAND4X0_HVT U2015 ( .A1(n1841), .A2(DP_OP_425J2_127_3477_n89), .A3(n1810), 
        .A4(n1813), .Y(n1063) );
  NAND2X0_HVT U2016 ( .A1(n1062), .A2(n1063), .Y(n_conv2_sum_d[26]) );
  NAND2X0_HVT U2017 ( .A1(n1064), .A2(n1065), .Y(n_conv2_sum_c[21]) );
  INVX1_HVT U2018 ( .A(tmp_big1[6]), .Y(n1066) );
  AO22X1_HVT U2019 ( .A1(tmp_big2[6]), .A2(n1066), .A3(tmp_big2[7]), .A4(n2171), .Y(n2141) );
  AOI22X1_HVT U2021 ( .A1(n1671), .A2(DP_OP_423J2_125_3477_n72), .A3(n1528), 
        .A4(DP_OP_423J2_125_3477_n58), .Y(n1069) );
  NAND2X0_HVT U2023 ( .A1(DP_OP_422J2_124_3477_n75), .A2(
        DP_OP_422J2_124_3477_n114), .Y(n1071) );
  OAI21X1_HVT U2024 ( .A1(DP_OP_422J2_124_3477_n73), .A2(
        DP_OP_422J2_124_3477_n185), .A3(n1072), .Y(DP_OP_422J2_124_3477_n72)
         );
  NAND2X0_HVT U2026 ( .A1(DP_OP_424J2_126_3477_n75), .A2(
        DP_OP_424J2_126_3477_n114), .Y(n1074) );
  OAI21X1_HVT U2027 ( .A1(DP_OP_424J2_126_3477_n73), .A2(
        DP_OP_424J2_126_3477_n185), .A3(n1075), .Y(DP_OP_424J2_126_3477_n72)
         );
  NAND2X0_HVT U2028 ( .A1(n1591), .A2(DP_OP_422J2_124_3477_n266), .Y(n1076) );
  AND2X1_HVT U2029 ( .A1(n1076), .A2(DP_OP_422J2_124_3477_n265), .Y(
        DP_OP_422J2_124_3477_n261) );
  NAND3X0_HVT U2030 ( .A1(n1599), .A2(n1600), .A3(n1601), .Y(n1077) );
  NAND2X0_HVT U2031 ( .A1(n1077), .A2(DP_OP_422J2_124_3477_n351), .Y(
        DP_OP_422J2_124_3477_n217) );
  NAND3X0_HVT U2032 ( .A1(n1821), .A2(DP_OP_425J2_127_3477_n185), .A3(
        DP_OP_425J2_127_3477_n198), .Y(n1078) );
  NAND2X0_HVT U2033 ( .A1(DP_OP_425J2_127_3477_n182), .A2(
        DP_OP_425J2_127_3477_n185), .Y(n1079) );
  NAND3X0_HVT U2034 ( .A1(n1078), .A2(DP_OP_425J2_127_3477_n162), .A3(n1079), 
        .Y(n1080) );
  INVX0_HVT U2035 ( .A(DP_OP_425J2_127_3477_n165), .Y(n1081) );
  AND2X1_HVT U2036 ( .A1(n1080), .A2(n1081), .Y(n1822) );
  NAND2X0_HVT U2037 ( .A1(DP_OP_424J2_126_3477_n297), .A2(n1736), .Y(n1082) );
  NAND2X0_HVT U2038 ( .A1(DP_OP_424J2_126_3477_n257), .A2(n1082), .Y(n1737) );
  INVX0_HVT U2039 ( .A(DP_OP_424J2_126_3477_n96), .Y(n1083) );
  OA21X1_HVT U2040 ( .A1(DP_OP_424J2_126_3477_n110), .A2(
        DP_OP_424J2_126_3477_n93), .A3(n1083), .Y(n1744) );
  NAND2X0_HVT U2041 ( .A1(DP_OP_423J2_125_3477_n252), .A2(n1636), .Y(n1084) );
  INVX0_HVT U2042 ( .A(n1610), .Y(n1085) );
  AND2X1_HVT U2043 ( .A1(n1085), .A2(n1622), .Y(n1086) );
  HADDX1_HVT U2044 ( .A0(n1086), .B0(n1291), .SO(n_conv2_sum_b[10]) );
  AO22X2_HVT U2045 ( .A1(DP_OP_422J2_124_3477_n279), .A2(
        DP_OP_422J2_124_3477_n129), .A3(n1557), .A4(n1558), .Y(n1087) );
  NAND2X0_HVT U2046 ( .A1(n1087), .A2(n1088), .Y(n_conv2_sum_a[22]) );
  AND2X1_HVT U2047 ( .A1(DP_OP_425J2_127_3477_n252), .A2(n1795), .Y(n1089) );
  HADDX1_HVT U2048 ( .A0(n1089), .B0(n1797), .SO(n_conv2_sum_d[5]) );
  AO22X2_HVT U2049 ( .A1(n1836), .A2(DP_OP_425J2_127_3477_n65), .A3(n1799), 
        .A4(n1838), .Y(n1090) );
  NAND4X0_HVT U2050 ( .A1(n1836), .A2(DP_OP_425J2_127_3477_n65), .A3(n1799), 
        .A4(n1838), .Y(n1091) );
  NAND2X0_HVT U2051 ( .A1(n1090), .A2(n1091), .Y(n_conv2_sum_d[28]) );
  AND2X1_HVT U2052 ( .A1(DP_OP_424J2_126_3477_n287), .A2(
        DP_OP_424J2_126_3477_n203), .Y(n1092) );
  HADDX1_HVT U2053 ( .A0(n1092), .B0(n182), .SO(n_conv2_sum_c[14]) );
  NAND2X0_HVT U2054 ( .A1(n1093), .A2(n1094), .Y(n_conv2_sum_c[23]) );
  INVX0_HVT U2055 ( .A(n619), .Y(n1095) );
  AND4X1_HVT U2056 ( .A1(src_window[57]), .A2(conv2_sum_b[1]), .A3(
        conv_weight_box[2]), .A4(n1484), .Y(n1117) );
  AO22X1_HVT U2057 ( .A1(tmp_big2[11]), .A2(n2178), .A3(tmp_big1[11]), .A4(
        n1504), .Y(data_out[11]) );
  NAND2X0_HVT U2058 ( .A1(DP_OP_425J2_127_3477_n96), .A2(n1841), .Y(n1096) );
  AND2X1_HVT U2059 ( .A1(n1096), .A2(DP_OP_425J2_127_3477_n89), .Y(
        DP_OP_425J2_127_3477_n85) );
  AO222X1_HVT U2060 ( .A1(DP_OP_424J2_126_3477_n827), .A2(
        DP_OP_424J2_126_3477_n1020), .A3(DP_OP_424J2_126_3477_n827), .A4(
        DP_OP_424J2_126_3477_n825), .A5(DP_OP_424J2_126_3477_n1020), .A6(
        DP_OP_424J2_126_3477_n825), .Y(DP_OP_424J2_126_3477_n822) );
  AOI21X1_HVT U2061 ( .A1(DP_OP_422J2_124_3477_n177), .A2(
        DP_OP_422J2_124_3477_n111), .A3(DP_OP_422J2_124_3477_n114), .Y(
        DP_OP_422J2_124_3477_n110) );
  INVX0_HVT U2062 ( .A(DP_OP_424J2_126_3477_n214), .Y(n1097) );
  AND2X1_HVT U2063 ( .A1(DP_OP_424J2_126_3477_n219), .A2(n1097), .Y(
        DP_OP_424J2_126_3477_n212) );
  INVX0_HVT U2064 ( .A(n1773), .Y(n1098) );
  NAND2X0_HVT U2065 ( .A1(DP_OP_425J2_127_3477_n237), .A2(n1772), .Y(n1100) );
  HADDX1_HVT U2066 ( .A0(n1099), .B0(n1100), .SO(n_conv2_sum_d[9]) );
  INVX0_HVT U2067 ( .A(DP_OP_422J2_124_3477_n267), .Y(n1101) );
  AND2X1_HVT U2068 ( .A1(n1101), .A2(DP_OP_422J2_124_3477_n268), .Y(n1102) );
  HADDX1_HVT U2069 ( .A0(n1102), .B0(DP_OP_422J2_124_3477_n269), .SO(
        n_conv2_sum_a[1]) );
  AND2X1_HVT U2070 ( .A1(n1544), .A2(n1573), .Y(n1103) );
  HADDX1_HVT U2071 ( .A0(n1103), .B0(DP_OP_422J2_124_3477_n232), .SO(
        n_conv2_sum_a[10]) );
  AO22X2_HVT U2072 ( .A1(n1588), .A2(DP_OP_422J2_124_3477_n120), .A3(n1552), 
        .A4(n1554), .Y(n1104) );
  NAND2X0_HVT U2073 ( .A1(n1104), .A2(n1105), .Y(n_conv2_sum_a[23]) );
  AND2X1_HVT U2074 ( .A1(DP_OP_425J2_127_3477_n249), .A2(
        DP_OP_425J2_127_3477_n295), .Y(n1106) );
  HADDX1_HVT U2075 ( .A0(n1106), .B0(DP_OP_425J2_127_3477_n250), .SO(
        n_conv2_sum_d[6]) );
  AOI21X1_HVT U2076 ( .A1(DP_OP_425J2_127_3477_n233), .A2(
        DP_OP_425J2_127_3477_n219), .A3(DP_OP_425J2_127_3477_n220), .Y(n1107)
         );
  NAND2X0_HVT U2077 ( .A1(DP_OP_425J2_127_3477_n217), .A2(n1814), .Y(n1108) );
  HADDX1_HVT U2078 ( .A0(n1107), .B0(n1108), .SO(n_conv2_sum_d[12]) );
  AO22X2_HVT U2079 ( .A1(n1835), .A2(DP_OP_425J2_127_3477_n47), .A3(n1802), 
        .A4(n1803), .Y(n1109) );
  NAND4X0_HVT U2080 ( .A1(n1835), .A2(DP_OP_425J2_127_3477_n47), .A3(n1802), 
        .A4(n1803), .Y(n1110) );
  NAND2X0_HVT U2081 ( .A1(n1109), .A2(n1110), .Y(n_conv2_sum_d[30]) );
  NAND2X0_HVT U2082 ( .A1(n182), .A2(n1765), .Y(n1111) );
  NAND3X0_HVT U2083 ( .A1(n1755), .A2(n1111), .A3(n1112), .Y(n_conv2_sum_c[20]) );
  AO22X2_HVT U2084 ( .A1(DP_OP_424J2_126_3477_n274), .A2(
        DP_OP_424J2_126_3477_n78), .A3(n1351), .A4(n1352), .Y(n1113) );
  NAND2X0_HVT U2085 ( .A1(n1113), .A2(n1114), .Y(n_conv2_sum_c[27]) );
  FADDX1_HVT U2086 ( .A(n1115), .B(n1116), .CI(n1117), .S(
        DP_OP_423J2_125_3477_n1785) );
  INVX0_HVT U2087 ( .A(tmp_big1[25]), .Y(n1118) );
  NAND2X0_HVT U2088 ( .A1(tmp_big2[25]), .A2(n1118), .Y(n2148) );
  AOI22X1_HVT U2090 ( .A1(n1586), .A2(DP_OP_422J2_124_3477_n72), .A3(n1525), 
        .A4(DP_OP_422J2_124_3477_n58), .Y(n1120) );
  NAND2X0_HVT U2093 ( .A1(DP_OP_425J2_127_3477_n75), .A2(
        DP_OP_425J2_127_3477_n114), .Y(n1123) );
  OAI21X1_HVT U2094 ( .A1(DP_OP_425J2_127_3477_n73), .A2(
        DP_OP_425J2_127_3477_n185), .A3(n1124), .Y(DP_OP_425J2_127_3477_n72)
         );
  INVX0_HVT U2095 ( .A(n1436), .Y(n1125) );
  NAND3X0_HVT U2096 ( .A1(n1626), .A2(n1623), .A3(n1125), .Y(n1627) );
  INVX0_HVT U2097 ( .A(DP_OP_423J2_125_3477_n72), .Y(n1126) );
  OAI21X1_HVT U2098 ( .A1(DP_OP_423J2_125_3477_n190), .A2(
        DP_OP_423J2_125_3477_n69), .A3(n1126), .Y(DP_OP_423J2_125_3477_n68) );
  NAND2X0_HVT U2099 ( .A1(n1590), .A2(DP_OP_422J2_124_3477_n258), .Y(n1127) );
  AND2X1_HVT U2100 ( .A1(n1127), .A2(DP_OP_422J2_124_3477_n257), .Y(
        DP_OP_422J2_124_3477_n253) );
  NAND2X0_HVT U2101 ( .A1(n1840), .A2(DP_OP_425J2_127_3477_n266), .Y(n1128) );
  AND2X1_HVT U2102 ( .A1(n1128), .A2(DP_OP_425J2_127_3477_n265), .Y(
        DP_OP_425J2_127_3477_n261) );
  INVX0_HVT U2103 ( .A(DP_OP_425J2_127_3477_n214), .Y(n1129) );
  AND2X1_HVT U2104 ( .A1(DP_OP_425J2_127_3477_n219), .A2(n1129), .Y(
        DP_OP_425J2_127_3477_n212) );
  OAI21X1_HVT U2105 ( .A1(DP_OP_425J2_127_3477_n107), .A2(
        DP_OP_425J2_127_3477_n13), .A3(DP_OP_425J2_127_3477_n110), .Y(n1825)
         );
  INVX0_HVT U2106 ( .A(DP_OP_424J2_126_3477_n220), .Y(n1130) );
  OAI21X2_HVT U2107 ( .A1(DP_OP_424J2_126_3477_n214), .A2(n1130), .A3(
        DP_OP_424J2_126_3477_n217), .Y(DP_OP_424J2_126_3477_n213) );
  NAND3X0_HVT U2108 ( .A1(n1747), .A2(DP_OP_424J2_126_3477_n185), .A3(
        DP_OP_424J2_126_3477_n198), .Y(n1131) );
  NAND2X0_HVT U2109 ( .A1(DP_OP_424J2_126_3477_n182), .A2(
        DP_OP_424J2_126_3477_n185), .Y(n1132) );
  INVX0_HVT U2110 ( .A(DP_OP_424J2_126_3477_n165), .Y(n1133) );
  NAND3X0_HVT U2111 ( .A1(n1131), .A2(DP_OP_424J2_126_3477_n162), .A3(n1132), 
        .Y(n1134) );
  AND2X1_HVT U2112 ( .A1(n1134), .A2(n1133), .Y(n1748) );
  NAND2X0_HVT U2113 ( .A1(DP_OP_424J2_126_3477_n50), .A2(n1758), .Y(n1135) );
  AND2X1_HVT U2114 ( .A1(n1135), .A2(DP_OP_424J2_126_3477_n47), .Y(n1769) );
  INVX0_HVT U2115 ( .A(DP_OP_424J2_126_3477_n259), .Y(n1136) );
  NAND2X0_HVT U2116 ( .A1(n1136), .A2(DP_OP_424J2_126_3477_n260), .Y(n1137) );
  HADDX1_HVT U2117 ( .A0(DP_OP_424J2_126_3477_n261), .B0(n1137), .SO(
        n_conv2_sum_c[3]) );
  AND2X1_HVT U2118 ( .A1(DP_OP_423J2_125_3477_n249), .A2(
        DP_OP_423J2_125_3477_n295), .Y(n1138) );
  NAND2X0_HVT U2119 ( .A1(n1612), .A2(DP_OP_423J2_125_3477_n240), .Y(n1139) );
  HADDX1_HVT U2120 ( .A0(n71), .B0(n1139), .SO(n_conv2_sum_b[8]) );
  AND2X1_HVT U2121 ( .A1(DP_OP_422J2_124_3477_n265), .A2(n1591), .Y(n1140) );
  HADDX1_HVT U2122 ( .A0(n1140), .B0(DP_OP_422J2_124_3477_n266), .SO(
        n_conv2_sum_a[2]) );
  AOI21X1_HVT U2123 ( .A1(DP_OP_422J2_124_3477_n232), .A2(n1544), .A3(n6), .Y(
        n1141) );
  NAND2X0_HVT U2124 ( .A1(DP_OP_422J2_124_3477_n226), .A2(n1534), .Y(n1142) );
  HADDX1_HVT U2125 ( .A0(n1141), .B0(n1142), .SO(n_conv2_sum_a[11]) );
  AO22X2_HVT U2126 ( .A1(DP_OP_422J2_124_3477_n277), .A2(
        DP_OP_422J2_124_3477_n105), .A3(n1581), .A4(DP_OP_422J2_124_3477_n110), 
        .Y(n1143) );
  NAND2X0_HVT U2127 ( .A1(n1143), .A2(n1144), .Y(n_conv2_sum_a[24]) );
  NAND2X0_HVT U2128 ( .A1(DP_OP_425J2_127_3477_n244), .A2(n1794), .Y(n1145) );
  HADDX1_HVT U2129 ( .A0(DP_OP_425J2_127_3477_n245), .B0(n1145), .SO(
        n_conv2_sum_d[7]) );
  AND2X1_HVT U2130 ( .A1(DP_OP_425J2_127_3477_n287), .A2(
        DP_OP_425J2_127_3477_n203), .Y(n1146) );
  HADDX1_HVT U2131 ( .A0(n1146), .B0(n1823), .SO(n_conv2_sum_d[14]) );
  NAND4X0_HVT U2132 ( .A1(n1833), .A2(DP_OP_425J2_127_3477_n38), .A3(n1793), 
        .A4(n1847), .Y(n1148) );
  NAND2X0_HVT U2133 ( .A1(n1147), .A2(n1148), .Y(n_conv2_sum_d[31]) );
  INVX0_HVT U2134 ( .A(n1712), .Y(n1149) );
  AND2X1_HVT U2135 ( .A1(n1149), .A2(n1732), .Y(n1150) );
  HADDX1_HVT U2136 ( .A0(n1150), .B0(DP_OP_424J2_126_3477_n233), .SO(
        n_conv2_sum_c[10]) );
  AND2X1_HVT U2137 ( .A1(DP_OP_424J2_126_3477_n110), .A2(n1749), .Y(n1151) );
  NAND2X0_HVT U2138 ( .A1(n1152), .A2(n1153), .Y(n_conv2_sum_c[28]) );
  INVX0_HVT U2139 ( .A(n843), .Y(n1154) );
  INVX0_HVT U2140 ( .A(tmp_big1[22]), .Y(n1155) );
  AO22X1_HVT U2141 ( .A1(tmp_big2[23]), .A2(n2162), .A3(tmp_big2[22]), .A4(
        n1155), .Y(n2126) );
  NAND2X0_HVT U2142 ( .A1(n2039), .A2(conv2_sum_a[16]), .Y(n1156) );
  OA22X1_HVT U2143 ( .A1(conv2_sum_b[17]), .A2(n1899), .A3(conv2_sum_b[16]), 
        .A4(n1156), .Y(n2015) );
  NAND2X0_HVT U2144 ( .A1(DP_OP_423J2_125_3477_n75), .A2(
        DP_OP_423J2_125_3477_n114), .Y(n1157) );
  OAI21X1_HVT U2146 ( .A1(DP_OP_423J2_125_3477_n73), .A2(
        DP_OP_423J2_125_3477_n185), .A3(n1159), .Y(DP_OP_423J2_125_3477_n72)
         );
  NAND2X0_HVT U2147 ( .A1(DP_OP_424J2_126_3477_n96), .A2(n1763), .Y(n1160) );
  AND2X1_HVT U2148 ( .A1(n1160), .A2(DP_OP_424J2_126_3477_n89), .Y(
        DP_OP_424J2_126_3477_n85) );
  NAND2X0_HVT U2149 ( .A1(n1762), .A2(DP_OP_424J2_126_3477_n266), .Y(n1161) );
  AND2X1_HVT U2150 ( .A1(n1161), .A2(DP_OP_424J2_126_3477_n265), .Y(
        DP_OP_424J2_126_3477_n261) );
  INVX0_HVT U2151 ( .A(DP_OP_425J2_127_3477_n127), .Y(n1162) );
  OA21X1_HVT U2152 ( .A1(DP_OP_425J2_127_3477_n141), .A2(
        DP_OP_425J2_127_3477_n124), .A3(n1162), .Y(n1807) );
  AO22X1_HVT U2153 ( .A1(conv2_sum_a[4]), .A2(n1437), .A3(conv2_sum_b[4]), 
        .A4(n1533), .Y(tmp_big1[4]) );
  INVX0_HVT U2154 ( .A(n1612), .Y(n1163) );
  OA21X1_HVT U2155 ( .A1(n71), .A2(n1163), .A3(DP_OP_423J2_125_3477_n240), .Y(
        n1164) );
  NAND2X0_HVT U2156 ( .A1(DP_OP_423J2_125_3477_n237), .A2(n1611), .Y(n1165) );
  HADDX1_HVT U2157 ( .A0(n1164), .B0(n1165), .SO(n_conv2_sum_b[9]) );
  AOI21X1_HVT U2158 ( .A1(n1291), .A2(n1622), .A3(n1610), .Y(n1166) );
  NAND2X0_HVT U2159 ( .A1(DP_OP_423J2_125_3477_n226), .A2(n1609), .Y(n1167) );
  HADDX1_HVT U2160 ( .A0(n1166), .B0(n1167), .SO(n_conv2_sum_b[11]) );
  INVX0_HVT U2161 ( .A(n1528), .Y(n1168) );
  AND2X1_HVT U2162 ( .A1(n1168), .A2(n1677), .Y(n1169) );
  HADDX1_HVT U2163 ( .A0(n1169), .B0(n1436), .SO(n_conv2_sum_b[14]) );
  INVX0_HVT U2164 ( .A(DP_OP_422J2_124_3477_n259), .Y(n1170) );
  NAND2X0_HVT U2165 ( .A1(n1170), .A2(DP_OP_422J2_124_3477_n260), .Y(n1171) );
  HADDX1_HVT U2166 ( .A0(DP_OP_422J2_124_3477_n261), .B0(n1171), .SO(
        n_conv2_sum_a[3]) );
  NAND2X0_HVT U2167 ( .A1(DP_OP_422J2_124_3477_n244), .A2(n1579), .Y(n1172) );
  HADDX1_HVT U2168 ( .A0(DP_OP_422J2_124_3477_n245), .B0(n1172), .SO(
        n_conv2_sum_a[7]) );
  AOI21X1_HVT U2169 ( .A1(DP_OP_422J2_124_3477_n232), .A2(
        DP_OP_422J2_124_3477_n219), .A3(DP_OP_422J2_124_3477_n220), .Y(n1173)
         );
  INVX0_HVT U2170 ( .A(n914), .Y(n1174) );
  NAND2X0_HVT U2171 ( .A1(n1174), .A2(DP_OP_422J2_124_3477_n217), .Y(n1175) );
  HADDX1_HVT U2172 ( .A0(n1173), .B0(n1175), .SO(n_conv2_sum_a[12]) );
  AO22X2_HVT U2173 ( .A1(DP_OP_422J2_124_3477_n276), .A2(
        DP_OP_422J2_124_3477_n98), .A3(n1559), .A4(n1560), .Y(n1176) );
  NAND2X0_HVT U2174 ( .A1(n1176), .A2(n1177), .Y(n_conv2_sum_a[25]) );
  AND2X1_HVT U2175 ( .A1(DP_OP_425J2_127_3477_n265), .A2(n1840), .Y(n1178) );
  HADDX1_HVT U2176 ( .A0(n1178), .B0(DP_OP_425J2_127_3477_n266), .SO(
        n_conv2_sum_d[2]) );
  NAND2X0_HVT U2177 ( .A1(n1773), .A2(DP_OP_425J2_127_3477_n240), .Y(n1179) );
  AOI21X1_HVT U2178 ( .A1(DP_OP_425J2_127_3477_n233), .A2(
        DP_OP_425J2_127_3477_n212), .A3(DP_OP_425J2_127_3477_n213), .Y(n1180)
         );
  NAND2X0_HVT U2179 ( .A1(DP_OP_425J2_127_3477_n210), .A2(n1827), .Y(n1181) );
  HADDX1_HVT U2180 ( .A0(n1180), .B0(n1181), .SO(n_conv2_sum_d[13]) );
  NAND2X0_HVT U2181 ( .A1(n1823), .A2(n1843), .Y(n1182) );
  OR2X2_HVT U2182 ( .A1(n1823), .A2(n1829), .Y(n1183) );
  NAND3X0_HVT U2183 ( .A1(n1830), .A2(n1182), .A3(n1183), .Y(n_conv2_sum_d[20]) );
  AO22X1_HVT U2184 ( .A1(DP_OP_425J2_127_3477_n274), .A2(
        DP_OP_425J2_127_3477_n78), .A3(n1367), .A4(n1368), .Y(n1184) );
  NAND4X0_HVT U2185 ( .A1(DP_OP_425J2_127_3477_n274), .A2(
        DP_OP_425J2_127_3477_n78), .A3(n1367), .A4(n1368), .Y(n1185) );
  NAND2X0_HVT U2186 ( .A1(n1184), .A2(n1185), .Y(n_conv2_sum_d[27]) );
  NAND2X0_HVT U2187 ( .A1(DP_OP_424J2_126_3477_n244), .A2(n1734), .Y(n1186) );
  HADDX1_HVT U2188 ( .A0(DP_OP_424J2_126_3477_n245), .B0(n1186), .SO(
        n_conv2_sum_c[7]) );
  AOI21X1_HVT U2189 ( .A1(DP_OP_424J2_126_3477_n233), .A2(n1732), .A3(n1712), 
        .Y(n1187) );
  NAND2X0_HVT U2190 ( .A1(DP_OP_424J2_126_3477_n226), .A2(n1711), .Y(n1188) );
  HADDX1_HVT U2191 ( .A0(n1187), .B0(n1188), .SO(n_conv2_sum_c[11]) );
  NAND2X0_HVT U2192 ( .A1(n1189), .A2(n1190), .Y(n_conv2_sum_c[29]) );
  FADDX1_HVT U2193 ( .A(DP_OP_423J2_125_3477_n968), .B(
        DP_OP_423J2_125_3477_n970), .CI(n1191), .S(DP_OP_423J2_125_3477_n749)
         );
  INVX0_HVT U2194 ( .A(n92), .Y(n1192) );
  AOI22X2_HVT U2195 ( .A1(n92), .A2(conv1_sram_rdata_weight[37]), .A3(n1192), 
        .A4(conv2_sram_rdata_weight[37]), .Y(DP_OP_425J2_127_3477_n2188) );
  NAND2X0_HVT U2196 ( .A1(n2159), .A2(tmp_big2[19]), .Y(n1193) );
  NAND2X0_HVT U2197 ( .A1(tmp_big1[18]), .A2(n1193), .Y(n1194) );
  OA22X1_HVT U2198 ( .A1(n2159), .A2(tmp_big2[19]), .A3(tmp_big2[18]), .A4(
        n1194), .Y(n1943) );
  INVX1_HVT U2199 ( .A(tmp_big2[24]), .Y(n1195) );
  AND2X1_HVT U2200 ( .A1(tmp_big1[24]), .A2(n1195), .Y(n1925) );
  NAND2X0_HVT U2201 ( .A1(DP_OP_423J2_125_3477_n146), .A2(
        DP_OP_423J2_125_3477_n165), .Y(n1196) );
  AOI22X1_HVT U2203 ( .A1(n488), .A2(conv2_sum_a[3]), .A3(n2174), .A4(
        conv2_sum_b[3]), .Y(n1985) );
  INVX1_HVT U2204 ( .A(n1436), .Y(n1198) );
  NAND3X0_HVT U2205 ( .A1(n1616), .A2(n1615), .A3(n1198), .Y(n1617) );
  INVX0_HVT U2206 ( .A(DP_OP_422J2_124_3477_n72), .Y(n1199) );
  OAI21X1_HVT U2207 ( .A1(DP_OP_422J2_124_3477_n190), .A2(
        DP_OP_422J2_124_3477_n69), .A3(n1199), .Y(DP_OP_422J2_124_3477_n68) );
  INVX0_HVT U2208 ( .A(DP_OP_425J2_127_3477_n220), .Y(n1200) );
  OAI21X2_HVT U2209 ( .A1(DP_OP_425J2_127_3477_n214), .A2(n1200), .A3(
        DP_OP_425J2_127_3477_n217), .Y(DP_OP_425J2_127_3477_n213) );
  INVX0_HVT U2210 ( .A(DP_OP_425J2_127_3477_n96), .Y(n1201) );
  OA21X1_HVT U2211 ( .A1(DP_OP_425J2_127_3477_n110), .A2(
        DP_OP_425J2_127_3477_n93), .A3(n1201), .Y(n1813) );
  AND2X1_HVT U2212 ( .A1(n1665), .A2(DP_OP_423J2_125_3477_n244), .Y(n1202) );
  INVX0_HVT U2213 ( .A(n1522), .Y(n1203) );
  NAND2X0_HVT U2214 ( .A1(DP_OP_423J2_125_3477_n217), .A2(n1655), .Y(n1205) );
  HADDX1_HVT U2215 ( .A0(n1204), .B0(n1205), .SO(n_conv2_sum_b[12]) );
  INVX0_HVT U2216 ( .A(DP_OP_422J2_124_3477_n251), .Y(n1206) );
  NAND2X0_HVT U2217 ( .A1(n1206), .A2(DP_OP_422J2_124_3477_n252), .Y(n1207) );
  HADDX1_HVT U2218 ( .A0(DP_OP_422J2_124_3477_n253), .B0(n1207), .SO(
        n_conv2_sum_a[5]) );
  NAND2X0_HVT U2219 ( .A1(n1537), .A2(DP_OP_422J2_124_3477_n240), .Y(n1208) );
  HADDX1_HVT U2220 ( .A0(DP_OP_422J2_124_3477_n241), .B0(n1208), .SO(
        n_conv2_sum_a[8]) );
  AOI21X1_HVT U2221 ( .A1(DP_OP_422J2_124_3477_n232), .A2(
        DP_OP_422J2_124_3477_n212), .A3(DP_OP_422J2_124_3477_n213), .Y(n1209)
         );
  INVX0_HVT U2222 ( .A(DP_OP_422J2_124_3477_n209), .Y(n1210) );
  NAND2X0_HVT U2223 ( .A1(n1210), .A2(DP_OP_422J2_124_3477_n210), .Y(n1211) );
  HADDX1_HVT U2224 ( .A0(n1209), .B0(n1211), .SO(n_conv2_sum_a[13]) );
  AO22X2_HVT U2225 ( .A1(n1587), .A2(DP_OP_422J2_124_3477_n89), .A3(n1555), 
        .A4(n1556), .Y(n1212) );
  NAND4X0_HVT U2226 ( .A1(n1555), .A2(DP_OP_422J2_124_3477_n89), .A3(n1587), 
        .A4(n1556), .Y(n1213) );
  NAND2X0_HVT U2227 ( .A1(n1212), .A2(n1213), .Y(n_conv2_sum_a[26]) );
  INVX0_HVT U2228 ( .A(DP_OP_425J2_127_3477_n259), .Y(n1214) );
  NAND2X0_HVT U2229 ( .A1(n1214), .A2(DP_OP_425J2_127_3477_n260), .Y(n1215) );
  HADDX1_HVT U2230 ( .A0(DP_OP_425J2_127_3477_n261), .B0(n1215), .SO(
        n_conv2_sum_d[3]) );
  INVX0_HVT U2231 ( .A(n1771), .Y(n1216) );
  AND2X1_HVT U2232 ( .A1(n1216), .A2(n1791), .Y(n1217) );
  HADDX1_HVT U2233 ( .A0(n1217), .B0(DP_OP_425J2_127_3477_n233), .SO(
        n_conv2_sum_d[10]) );
  AO22X2_HVT U2234 ( .A1(DP_OP_425J2_127_3477_n272), .A2(
        DP_OP_425J2_127_3477_n52), .A3(n1801), .A4(DP_OP_425J2_127_3477_n57), 
        .Y(n1218) );
  NAND4X0_HVT U2235 ( .A1(DP_OP_425J2_127_3477_n272), .A2(
        DP_OP_425J2_127_3477_n52), .A3(n1801), .A4(DP_OP_425J2_127_3477_n57), 
        .Y(n1219) );
  NAND2X0_HVT U2236 ( .A1(n1218), .A2(n1219), .Y(n_conv2_sum_d[29]) );
  INVX0_HVT U2237 ( .A(DP_OP_424J2_126_3477_n267), .Y(n1220) );
  AND2X1_HVT U2238 ( .A1(n1220), .A2(DP_OP_424J2_126_3477_n268), .Y(n1221) );
  HADDX1_HVT U2239 ( .A0(n1221), .B0(DP_OP_424J2_126_3477_n269), .SO(
        n_conv2_sum_c[1]) );
  AND2X1_HVT U2240 ( .A1(DP_OP_424J2_126_3477_n252), .A2(n1735), .Y(n1222) );
  NAND2X0_HVT U2241 ( .A1(n1714), .A2(DP_OP_424J2_126_3477_n240), .Y(n1223) );
  AOI21X1_HVT U2242 ( .A1(DP_OP_424J2_126_3477_n233), .A2(
        DP_OP_424J2_126_3477_n219), .A3(DP_OP_424J2_126_3477_n220), .Y(n1224)
         );
  NAND2X0_HVT U2243 ( .A1(DP_OP_424J2_126_3477_n217), .A2(n1745), .Y(n1225) );
  HADDX1_HVT U2244 ( .A0(n1224), .B0(n1225), .SO(n_conv2_sum_c[12]) );
  AO22X2_HVT U2245 ( .A1(DP_OP_424J2_126_3477_n276), .A2(
        DP_OP_424J2_126_3477_n98), .A3(n1349), .A4(n1348), .Y(n1226) );
  NAND2X0_HVT U2246 ( .A1(n1226), .A2(n1227), .Y(n_conv2_sum_c[25]) );
  NAND2X0_HVT U2247 ( .A1(n1228), .A2(n1229), .Y(n_conv2_sum_c[30]) );
  INVX1_HVT U2248 ( .A(n1514), .Y(n1512) );
  NAND2X0_HVT U2249 ( .A1(DP_OP_423J2_125_3477_n969), .A2(
        DP_OP_423J2_125_3477_n953), .Y(n1230) );
  AO222X1_HVT U2250 ( .A1(DP_OP_423J2_125_3477_n749), .A2(
        DP_OP_423J2_125_3477_n753), .A3(DP_OP_423J2_125_3477_n749), .A4(n1231), 
        .A5(DP_OP_423J2_125_3477_n753), .A6(n1231), .Y(
        DP_OP_423J2_125_3477_n710) );
  FADDX1_HVT U2251 ( .A(DP_OP_422J2_124_3477_n1498), .B(
        DP_OP_422J2_124_3477_n1486), .CI(DP_OP_422J2_124_3477_n1488), .S(n1232) );
  FADDX1_HVT U2252 ( .A(DP_OP_422J2_124_3477_n1281), .B(
        DP_OP_422J2_124_3477_n1448), .CI(n1232), .S(DP_OP_422J2_124_3477_n1249) );
  FADDX1_HVT U2253 ( .A(DP_OP_425J2_127_3477_n1675), .B(
        DP_OP_425J2_127_3477_n1727), .CI(n1233), .S(DP_OP_425J2_127_3477_n1637) );
  NAND2X0_HVT U2254 ( .A1(DP_OP_423J2_125_3477_n96), .A2(n1672), .Y(n1234) );
  AND2X1_HVT U2255 ( .A1(n1234), .A2(DP_OP_423J2_125_3477_n89), .Y(
        DP_OP_423J2_125_3477_n85) );
  INVX0_HVT U2256 ( .A(n2170), .Y(n1235) );
  AO22X1_HVT U2257 ( .A1(N9), .A2(n1235), .A3(tmp_big2[5]), .A4(n2178), .Y(
        data_out[5]) );
  NAND2X0_HVT U2258 ( .A1(n1676), .A2(DP_OP_423J2_125_3477_n266), .Y(n1236) );
  AND2X1_HVT U2259 ( .A1(n1236), .A2(DP_OP_423J2_125_3477_n265), .Y(
        DP_OP_423J2_125_3477_n261) );
  INVX0_HVT U2260 ( .A(DP_OP_423J2_125_3477_n17), .Y(n1237) );
  AND2X1_HVT U2261 ( .A1(n1638), .A2(n1237), .Y(n1424) );
  NAND2X0_HVT U2262 ( .A1(DP_OP_423J2_125_3477_n50), .A2(n1670), .Y(n1238) );
  AND2X1_HVT U2263 ( .A1(n1238), .A2(DP_OP_423J2_125_3477_n47), .Y(n1680) );
  INVX0_HVT U2264 ( .A(n914), .Y(n1239) );
  AND2X1_HVT U2265 ( .A1(DP_OP_422J2_124_3477_n219), .A2(n1239), .Y(
        DP_OP_422J2_124_3477_n212) );
  INVX0_HVT U2266 ( .A(DP_OP_422J2_124_3477_n171), .Y(n1240) );
  AND2X1_HVT U2267 ( .A1(DP_OP_422J2_124_3477_n176), .A2(n1240), .Y(
        DP_OP_422J2_124_3477_n169) );
  NAND2X0_HVT U2268 ( .A1(n1585), .A2(DP_OP_422J2_124_3477_n50), .Y(n1241) );
  NAND2X0_HVT U2269 ( .A1(DP_OP_422J2_124_3477_n47), .A2(n1241), .Y(n1594) );
  INVX0_HVT U2270 ( .A(DP_OP_425J2_127_3477_n72), .Y(n1242) );
  OA21X1_HVT U2271 ( .A1(DP_OP_425J2_127_3477_n190), .A2(
        DP_OP_425J2_127_3477_n69), .A3(n1242), .Y(n1838) );
  NAND2X0_HVT U2272 ( .A1(DP_OP_425J2_127_3477_n50), .A2(n1835), .Y(n1243) );
  AND2X1_HVT U2273 ( .A1(n1243), .A2(DP_OP_425J2_127_3477_n47), .Y(n1847) );
  INVX0_HVT U2274 ( .A(DP_OP_424J2_126_3477_n127), .Y(n1244) );
  OA21X1_HVT U2275 ( .A1(DP_OP_424J2_126_3477_n141), .A2(
        DP_OP_424J2_126_3477_n124), .A3(n1244), .Y(n1741) );
  INVX0_HVT U2276 ( .A(DP_OP_424J2_126_3477_n72), .Y(n1245) );
  OA21X1_HVT U2277 ( .A1(DP_OP_424J2_126_3477_n190), .A2(
        DP_OP_424J2_126_3477_n69), .A3(n1245), .Y(n1761) );
  INVX0_HVT U2278 ( .A(DP_OP_425J2_127_3477_n267), .Y(n1246) );
  AND2X1_HVT U2279 ( .A1(n1246), .A2(DP_OP_425J2_127_3477_n268), .Y(n1247) );
  HADDX1_HVT U2280 ( .A0(n1247), .B0(DP_OP_425J2_127_3477_n269), .SO(
        n_conv2_sum_d[1]) );
  AOI21X1_HVT U2281 ( .A1(n1291), .A2(DP_OP_423J2_125_3477_n212), .A3(
        DP_OP_423J2_125_3477_n213), .Y(n1248) );
  NAND2X0_HVT U2282 ( .A1(DP_OP_423J2_125_3477_n210), .A2(n1656), .Y(n1249) );
  HADDX1_HVT U2283 ( .A0(n1248), .B0(n1249), .SO(n_conv2_sum_b[13]) );
  AO22X1_HVT U2284 ( .A1(DP_OP_423J2_125_3477_n279), .A2(
        DP_OP_423J2_125_3477_n129), .A3(n1657), .A4(n1658), .Y(n1250) );
  NAND2X0_HVT U2285 ( .A1(n1251), .A2(n1250), .Y(n_conv2_sum_b[22]) );
  AND2X1_HVT U2286 ( .A1(DP_OP_422J2_124_3477_n257), .A2(n1590), .Y(n1252) );
  HADDX1_HVT U2287 ( .A0(n1252), .B0(DP_OP_422J2_124_3477_n258), .SO(
        n_conv2_sum_a[4]) );
  INVX0_HVT U2288 ( .A(DP_OP_422J2_124_3477_n248), .Y(n1253) );
  NAND2X0_HVT U2289 ( .A1(n1253), .A2(DP_OP_422J2_124_3477_n249), .Y(n1254) );
  HADDX1_HVT U2290 ( .A0(n1577), .B0(n1254), .SO(n_conv2_sum_a[6]) );
  INVX0_HVT U2291 ( .A(n1537), .Y(n1255) );
  NAND2X0_HVT U2292 ( .A1(DP_OP_422J2_124_3477_n237), .A2(n1536), .Y(n1257) );
  HADDX1_HVT U2293 ( .A0(n1256), .B0(n1257), .SO(n_conv2_sum_a[9]) );
  INVX0_HVT U2294 ( .A(n1525), .Y(n1258) );
  NAND2X0_HVT U2295 ( .A1(n1258), .A2(n1592), .Y(n1259) );
  NAND4X0_HVT U2296 ( .A1(n1561), .A2(DP_OP_422J2_124_3477_n78), .A3(
        DP_OP_422J2_124_3477_n274), .A4(n1562), .Y(n1261) );
  NAND2X0_HVT U2297 ( .A1(n1260), .A2(n1261), .Y(n_conv2_sum_a[27]) );
  AOI21X1_HVT U2298 ( .A1(DP_OP_425J2_127_3477_n233), .A2(n1791), .A3(n1771), 
        .Y(n1262) );
  NAND2X0_HVT U2299 ( .A1(DP_OP_425J2_127_3477_n226), .A2(n1770), .Y(n1263) );
  HADDX1_HVT U2300 ( .A0(n1262), .B0(n1263), .SO(n_conv2_sum_d[11]) );
  AND2X1_HVT U2301 ( .A1(DP_OP_425J2_127_3477_n110), .A2(n1824), .Y(n1264) );
  AO222X1_HVT U2302 ( .A1(n1781), .A2(n1264), .A3(n1823), .A4(n1844), .A5(
        n1826), .A6(n1825), .Y(n_conv2_sum_d[24]) );
  AND2X1_HVT U2303 ( .A1(DP_OP_424J2_126_3477_n265), .A2(n1762), .Y(n1265) );
  HADDX1_HVT U2304 ( .A0(n1265), .B0(DP_OP_424J2_126_3477_n266), .SO(
        n_conv2_sum_c[2]) );
  AND2X1_HVT U2305 ( .A1(DP_OP_424J2_126_3477_n257), .A2(
        DP_OP_424J2_126_3477_n297), .Y(n1266) );
  HADDX1_HVT U2306 ( .A0(n1266), .B0(n1736), .SO(n_conv2_sum_c[4]) );
  AND2X1_HVT U2307 ( .A1(DP_OP_424J2_126_3477_n249), .A2(
        DP_OP_424J2_126_3477_n295), .Y(n1267) );
  INVX0_HVT U2308 ( .A(n1714), .Y(n1268) );
  NAND2X0_HVT U2309 ( .A1(DP_OP_424J2_126_3477_n237), .A2(n1713), .Y(n1270) );
  HADDX1_HVT U2310 ( .A0(n1269), .B0(n1270), .SO(n_conv2_sum_c[9]) );
  AOI21X1_HVT U2311 ( .A1(DP_OP_424J2_126_3477_n233), .A2(
        DP_OP_424J2_126_3477_n212), .A3(DP_OP_424J2_126_3477_n213), .Y(n1271)
         );
  NAND2X0_HVT U2312 ( .A1(DP_OP_424J2_126_3477_n210), .A2(n1752), .Y(n1272) );
  HADDX1_HVT U2313 ( .A0(n1271), .B0(n1272), .SO(n_conv2_sum_c[13]) );
  AO22X1_HVT U2314 ( .A1(n1763), .A2(DP_OP_424J2_126_3477_n89), .A3(n1374), 
        .A4(n1744), .Y(n1273) );
  NAND2X0_HVT U2315 ( .A1(n1273), .A2(n1274), .Y(n_conv2_sum_c[26]) );
  NAND2X0_HVT U2316 ( .A1(n1275), .A2(n1276), .Y(n_conv2_sum_c[31]) );
  MUX21X1_HVT U2317 ( .A1(conv2_sram_rdata_weight[48]), .A2(
        conv1_sram_rdata_weight[48]), .S0(n345), .Y(conv_weight_box[33]) );
  INVX1_HVT U2318 ( .A(conv_weight_box[34]), .Y(DP_OP_423J2_125_3477_n2803) );
  INVX1_HVT U2319 ( .A(conv_weight_box[34]), .Y(n1444) );
  INVX2_HVT U2320 ( .A(conv_weight_box[31]), .Y(DP_OP_424J2_126_3477_n2231) );
  INVX2_HVT U2321 ( .A(conv_weight_box[31]), .Y(DP_OP_425J2_127_3477_n2231) );
  INVX2_HVT U2322 ( .A(DP_OP_424J2_126_3477_n2274), .Y(n1371) );
  NBUFFX4_HVT U2323 ( .A(DP_OP_424J2_126_3477_n2274), .Y(n1370) );
  INVX4_HVT U2324 ( .A(n1371), .Y(n1338) );
  MUX21X1_HVT U2325 ( .A1(conv2_sram_rdata_weight[54]), .A2(
        conv1_sram_rdata_weight[54]), .S0(n1418), .Y(conv_weight_box[38]) );
  INVX1_HVT U2326 ( .A(conv_weight_box[38]), .Y(n1427) );
  INVX2_HVT U2327 ( .A(conv_weight_box[37]), .Y(DP_OP_422J2_124_3477_n2276) );
  INVX2_HVT U2328 ( .A(conv_weight_box[37]), .Y(DP_OP_424J2_126_3477_n2276) );
  MUX21X1_HVT U2329 ( .A1(conv2_sram_rdata_weight[13]), .A2(
        conv1_sram_rdata_weight[13]), .S0(n241), .Y(conv_weight_box[9]) );
  MUX21X1_HVT U2330 ( .A1(conv1_sram_rdata_weight[44]), .A2(
        conv2_sram_rdata_weight[44]), .S0(n1396), .Y(conv_weight_box[30]) );
  INVX1_HVT U2331 ( .A(conv_weight_box[30]), .Y(DP_OP_423J2_125_3477_n2233) );
  INVX4_HVT U2332 ( .A(n1384), .Y(n1425) );
  MUX21X1_HVT U2333 ( .A1(conv2_sram_rdata_weight[36]), .A2(
        conv1_sram_rdata_weight[36]), .S0(n1418), .Y(conv_weight_box[24]) );
  MUX21X1_HVT U2334 ( .A1(conv2_sram_rdata_weight[39]), .A2(
        conv1_sram_rdata_weight[39]), .S0(n619), .Y(conv_weight_box[25]) );
  INVX2_HVT U2335 ( .A(conv_weight_box[58]), .Y(DP_OP_423J2_125_3477_n2452) );
  INVX2_HVT U2336 ( .A(conv_weight_box[58]), .Y(n1488) );
  INVX2_HVT U2337 ( .A(conv_weight_box[4]), .Y(DP_OP_423J2_125_3477_n2010) );
  INVX2_HVT U2338 ( .A(conv_weight_box[4]), .Y(DP_OP_424J2_126_3477_n2010) );
  INVX2_HVT U2339 ( .A(conv_weight_box[2]), .Y(DP_OP_422J2_124_3477_n2013) );
  INVX2_HVT U2340 ( .A(conv_weight_box[57]), .Y(DP_OP_425J2_127_3477_n2453) );
  INVX4_HVT U2341 ( .A(conv_weight_box[56]), .Y(n1331) );
  MUX21X1_HVT U2342 ( .A1(conv2_sram_rdata_weight[67]), .A2(
        conv1_sram_rdata_weight[67]), .S0(n92), .Y(conv_weight_box[46]) );
  MUX21X1_HVT U2343 ( .A1(conv2_sram_rdata_weight[61]), .A2(
        conv1_sram_rdata_weight[61]), .S0(n1418), .Y(conv_weight_box[42]) );
  INVX1_HVT U2344 ( .A(conv_weight_box[50]), .Y(n1400) );
  INVX2_HVT U2345 ( .A(DP_OP_425J2_127_3477_n2188), .Y(n1388) );
  AND3X1_HVT U2346 ( .A1(n1816), .A2(n1818), .A3(n1839), .Y(n1277) );
  INVX1_HVT U2347 ( .A(conv_weight_box[64]), .Y(DP_OP_425J2_127_3477_n2495) );
  AND2X1_HVT U2348 ( .A1(n2050), .A2(n2049), .Y(n1290) );
  INVX1_HVT U2349 ( .A(n1380), .Y(DP_OP_424J2_126_3477_n320) );
  NOR2X4_HVT U2350 ( .A1(n1279), .A2(DP_OP_422J2_124_3477_n2), .Y(n1295) );
  INVX1_HVT U2351 ( .A(n1381), .Y(DP_OP_425J2_127_3477_n330) );
  INVX1_HVT U2352 ( .A(n1382), .Y(DP_OP_423J2_125_3477_n312) );
  INVX1_HVT U2353 ( .A(n1383), .Y(DP_OP_422J2_124_3477_n306) );
  INVX1_HVT U2354 ( .A(n1331), .Y(n1332) );
  OA21X2_HVT U2355 ( .A1(n4), .A2(n1356), .A3(n1355), .Y(n1333) );
  INVX2_HVT U2356 ( .A(DP_OP_423J2_125_3477_n2538), .Y(n1363) );
  INVX0_HVT U2357 ( .A(n1363), .Y(n1334) );
  INVX0_HVT U2358 ( .A(n1363), .Y(n1335) );
  INVX1_HVT U2359 ( .A(n1363), .Y(n1336) );
  INVX1_HVT U2360 ( .A(n1378), .Y(n1340) );
  INVX2_HVT U2361 ( .A(n1378), .Y(n1341) );
  INVX2_HVT U2362 ( .A(n1378), .Y(n1342) );
  INVX1_HVT U2363 ( .A(n1388), .Y(n1343) );
  INVX2_HVT U2364 ( .A(n1388), .Y(n1344) );
  INVX2_HVT U2365 ( .A(n1388), .Y(n1345) );
  MUX21X1_HVT U2366 ( .A1(conv1_sram_rdata_weight[51]), .A2(
        conv2_sram_rdata_weight[51]), .S0(n1396), .Y(conv_weight_box[35]) );
  MUX21X1_HVT U2367 ( .A1(conv1_sram_rdata_weight[96]), .A2(
        conv2_sram_rdata_weight[96]), .S0(n1396), .Y(conv_weight_box[66]) );
  XNOR2X2_HVT U2368 ( .A1(n1520), .A2(DP_OP_425J2_127_3477_n12), .Y(
        n_conv2_sum_d[25]) );
  INVX1_HVT U2369 ( .A(tmp_big1[4]), .Y(n1918) );
  NOR2X2_HVT U2370 ( .A1(DP_OP_425J2_127_3477_n2357), .A2(n1386), .Y(
        DP_OP_425J2_127_3477_n2341) );
  OR2X2_HVT U2371 ( .A1(DP_OP_424J2_126_3477_n3019), .A2(n30), .Y(
        DP_OP_425J2_127_3477_n2019) );
  NOR2X4_HVT U2372 ( .A1(DP_OP_422J2_124_3477_n2356), .A2(
        DP_OP_423J2_125_3477_n2364), .Y(DP_OP_422J2_124_3477_n2340) );
  NOR2X4_HVT U2373 ( .A1(DP_OP_422J2_124_3477_n2357), .A2(
        DP_OP_423J2_125_3477_n2364), .Y(DP_OP_422J2_124_3477_n2341) );
  NOR2X0_HVT U2374 ( .A1(DP_OP_424J2_126_3477_n2136), .A2(
        DP_OP_423J2_125_3477_n2891), .Y(DP_OP_425J2_127_3477_n2860) );
  NBUFFX4_HVT U2375 ( .A(DP_OP_423J2_125_3477_n2364), .Y(n1386) );
  MUX21X2_HVT U2376 ( .A1(tmp_big2[15]), .A2(tmp_big1[15]), .S0(N9), .Y(
        data_out[15]) );
  OA21X2_HVT U2377 ( .A1(n4), .A2(n1356), .A3(n1355), .Y(n1346) );
  INVX2_HVT U2378 ( .A(n585), .Y(DP_OP_422J2_124_3477_n2142) );
  MUX21X1_HVT U2379 ( .A1(conv2_sram_rdata_weight[92]), .A2(
        conv1_sram_rdata_weight[92]), .S0(n241), .Y(conv_weight_box[62]) );
  MUX21X2_HVT U2380 ( .A1(conv2_sram_rdata_weight[95]), .A2(
        conv1_sram_rdata_weight[95]), .S0(n843), .Y(conv_weight_box[65]) );
  OA22X1_HVT U2381 ( .A1(n1929), .A2(n1485), .A3(n1931), .A4(n1930), .Y(
        DP_OP_423J2_125_3477_n2364) );
  OR2X1_HVT U2382 ( .A1(DP_OP_424J2_126_3477_n648), .A2(
        DP_OP_424J2_126_3477_n513), .Y(n1713) );
  AND2X4_HVT U2383 ( .A1(conv_weight_box[12]), .A2(src_window[90]), .Y(
        DP_OP_422J2_124_3477_n2951) );
  NAND2X0_HVT U2384 ( .A1(conv_weight_box[12]), .A2(src_window[95]), .Y(
        DP_OP_422J2_124_3477_n2946) );
  AO22X1_HVT U2385 ( .A1(DP_OP_422J2_124_3477_n547), .A2(
        DP_OP_422J2_124_3477_n680), .A3(n1347), .A4(DP_OP_422J2_124_3477_n678), 
        .Y(DP_OP_422J2_124_3477_n532) );
  OR2X1_HVT U2386 ( .A1(DP_OP_422J2_124_3477_n680), .A2(
        DP_OP_422J2_124_3477_n547), .Y(n1347) );
  XOR3X2_HVT U2387 ( .A1(DP_OP_422J2_124_3477_n547), .A2(
        DP_OP_422J2_124_3477_n680), .A3(DP_OP_422J2_124_3477_n678), .Y(
        DP_OP_422J2_124_3477_n533) );
  OA21X1_HVT U2388 ( .A1(DP_OP_424J2_126_3477_n102), .A2(
        DP_OP_424J2_126_3477_n110), .A3(DP_OP_424J2_126_3477_n105), .Y(n1348)
         );
  OA21X2_HVT U2389 ( .A1(n1742), .A2(n1740), .A3(n1743), .Y(
        DP_OP_424J2_126_3477_n110) );
  NBUFFX2_HVT U2390 ( .A(conv_weight_box[16]), .Y(n1350) );
  AND2X1_HVT U2391 ( .A1(conv_weight_box[16]), .A2(src_window[116]), .Y(
        DP_OP_422J2_124_3477_n2913) );
  NAND2X0_HVT U2392 ( .A1(n1350), .A2(src_window[119]), .Y(
        DP_OP_422J2_124_3477_n2910) );
  AND2X1_HVT U2393 ( .A1(n1350), .A2(src_window[117]), .Y(
        DP_OP_422J2_124_3477_n2912) );
  AND2X1_HVT U2394 ( .A1(n1350), .A2(src_window[113]), .Y(
        DP_OP_422J2_124_3477_n2916) );
  AND2X1_HVT U2395 ( .A1(n1350), .A2(src_window[112]), .Y(
        DP_OP_422J2_124_3477_n2917) );
  AND2X1_HVT U2396 ( .A1(n1350), .A2(src_window[118]), .Y(
        DP_OP_422J2_124_3477_n2911) );
  AND2X1_HVT U2397 ( .A1(n1350), .A2(src_window[114]), .Y(
        DP_OP_422J2_124_3477_n2915) );
  AND2X4_HVT U2398 ( .A1(n1350), .A2(src_window[115]), .Y(
        DP_OP_422J2_124_3477_n2914) );
  MUX21X1_HVT U2399 ( .A1(conv2_sum_d[5]), .A2(conv2_sum_c[5]), .S0(N7), .Y(
        tmp_big2[5]) );
  AO22X1_HVT U2400 ( .A1(n1851), .A2(n1533), .A3(n1437), .A4(n1852), .Y(n2170)
         );
  AND2X1_HVT U2401 ( .A1(n1354), .A2(n1277), .Y(n1353) );
  NAND2X0_HVT U2402 ( .A1(n1819), .A2(n1820), .Y(n1354) );
  NAND2X0_HVT U2403 ( .A1(n1832), .A2(DP_OP_425J2_127_3477_n158), .Y(n1808) );
  OA21X2_HVT U2404 ( .A1(n1923), .A2(n1356), .A3(n1355), .Y(
        DP_OP_424J2_126_3477_n2408) );
  NAND2X0_HVT U2405 ( .A1(n857), .A2(conv1_sram_rdata_weight[77]), .Y(n1355)
         );
  OA21X1_HVT U2406 ( .A1(DP_OP_424J2_126_3477_n209), .A2(
        DP_OP_424J2_126_3477_n217), .A3(DP_OP_424J2_126_3477_n210), .Y(n1357)
         );
  NAND2X0_HVT U2407 ( .A1(DP_OP_424J2_126_3477_n351), .A2(
        DP_OP_424J2_126_3477_n372), .Y(DP_OP_424J2_126_3477_n217) );
  AND2X1_HVT U2408 ( .A1(conv_weight_box[64]), .A2(src_window[275]), .Y(
        DP_OP_422J2_124_3477_n2466) );
  MUX21X1_HVT U2409 ( .A1(conv1_sram_rdata_weight[94]), .A2(
        conv2_sram_rdata_weight[94]), .S0(n1515), .Y(conv_weight_box[64]) );
  AO22X1_HVT U2410 ( .A1(DP_OP_425J2_127_3477_n523), .A2(
        DP_OP_425J2_127_3477_n656), .A3(n1358), .A4(DP_OP_425J2_127_3477_n654), 
        .Y(DP_OP_425J2_127_3477_n516) );
  OR2X1_HVT U2411 ( .A1(DP_OP_425J2_127_3477_n523), .A2(
        DP_OP_425J2_127_3477_n656), .Y(n1358) );
  XOR3X2_HVT U2412 ( .A1(DP_OP_425J2_127_3477_n523), .A2(
        DP_OP_425J2_127_3477_n656), .A3(DP_OP_425J2_127_3477_n654), .Y(
        DP_OP_425J2_127_3477_n517) );
  AO22X1_HVT U2413 ( .A1(DP_OP_422J2_124_3477_n518), .A2(
        DP_OP_422J2_124_3477_n425), .A3(n1359), .A4(n1360), .Y(
        DP_OP_422J2_124_3477_n420) );
  OR2X1_HVT U2414 ( .A1(DP_OP_422J2_124_3477_n518), .A2(
        DP_OP_422J2_124_3477_n425), .Y(n1359) );
  XOR3X2_HVT U2415 ( .A1(DP_OP_422J2_124_3477_n425), .A2(
        DP_OP_422J2_124_3477_n518), .A3(n1360), .Y(DP_OP_422J2_124_3477_n421)
         );
  NAND3X0_HVT U2416 ( .A1(n1510), .A2(n1511), .A3(n1509), .Y(n1360) );
  INVX2_HVT U2417 ( .A(n1361), .Y(DP_OP_425J2_127_3477_n2458) );
  NAND2X0_HVT U2418 ( .A1(conv_weight_box[65]), .A2(src_window[218]), .Y(
        DP_OP_425J2_127_3477_n2459) );
  AND2X1_HVT U2419 ( .A1(conv_weight_box[65]), .A2(src_window[219]), .Y(n1361)
         );
  NAND2X0_HVT U2420 ( .A1(conv_weight_box[65]), .A2(src_window[220]), .Y(
        DP_OP_425J2_127_3477_n2457) );
  NAND2X0_HVT U2421 ( .A1(n464), .A2(src_window[216]), .Y(
        DP_OP_425J2_127_3477_n2461) );
  NAND2X0_HVT U2422 ( .A1(n464), .A2(src_window[217]), .Y(
        DP_OP_425J2_127_3477_n2460) );
  NAND2X0_HVT U2423 ( .A1(n464), .A2(src_window[221]), .Y(
        DP_OP_425J2_127_3477_n2456) );
  NAND2X0_HVT U2424 ( .A1(n464), .A2(src_window[222]), .Y(
        DP_OP_425J2_127_3477_n2455) );
  AND2X4_HVT U2425 ( .A1(conv_weight_box[65]), .A2(src_window[223]), .Y(
        DP_OP_425J2_127_3477_n2454) );
  AND2X1_HVT U2426 ( .A1(n1350), .A2(src_window[61]), .Y(
        DP_OP_425J2_127_3477_n2912) );
  AND2X1_HVT U2427 ( .A1(conv_weight_box[16]), .A2(src_window[62]), .Y(
        DP_OP_425J2_127_3477_n2911) );
  NAND2X0_HVT U2428 ( .A1(n1350), .A2(src_window[63]), .Y(
        DP_OP_425J2_127_3477_n2910) );
  AND2X1_HVT U2429 ( .A1(n1350), .A2(src_window[57]), .Y(
        DP_OP_425J2_127_3477_n2916) );
  AND2X1_HVT U2430 ( .A1(n1350), .A2(src_window[60]), .Y(
        DP_OP_425J2_127_3477_n2913) );
  AND2X1_HVT U2431 ( .A1(n1350), .A2(src_window[56]), .Y(
        DP_OP_425J2_127_3477_n2917) );
  AND2X1_HVT U2432 ( .A1(n1350), .A2(src_window[58]), .Y(
        DP_OP_425J2_127_3477_n2915) );
  AND2X4_HVT U2433 ( .A1(n1350), .A2(src_window[59]), .Y(
        DP_OP_425J2_127_3477_n2914) );
  NBUFFX2_HVT U2434 ( .A(DP_OP_423J2_125_3477_n2538), .Y(n1362) );
  NAND2X0_HVT U2435 ( .A1(n1364), .A2(src_window[275]), .Y(
        DP_OP_423J2_125_3477_n2502) );
  NAND2X0_HVT U2436 ( .A1(conv_weight_box[56]), .A2(src_window[194]), .Y(
        DP_OP_425J2_127_3477_n2591) );
  NAND2X0_HVT U2437 ( .A1(n1332), .A2(src_window[192]), .Y(
        DP_OP_425J2_127_3477_n2593) );
  NAND2X0_HVT U2438 ( .A1(n1332), .A2(src_window[197]), .Y(
        DP_OP_425J2_127_3477_n2588) );
  NAND2X0_HVT U2439 ( .A1(n1366), .A2(src_window[196]), .Y(
        DP_OP_425J2_127_3477_n2589) );
  NAND2X0_HVT U2440 ( .A1(n1366), .A2(src_window[193]), .Y(
        DP_OP_425J2_127_3477_n2592) );
  NAND2X0_HVT U2441 ( .A1(n1366), .A2(src_window[195]), .Y(
        DP_OP_425J2_127_3477_n2590) );
  NAND2X0_HVT U2442 ( .A1(n1366), .A2(src_window[198]), .Y(
        DP_OP_425J2_127_3477_n2587) );
  NAND2X0_HVT U2443 ( .A1(n1832), .A2(DP_OP_425J2_127_3477_n80), .Y(n1367) );
  OA21X2_HVT U2444 ( .A1(DP_OP_425J2_127_3477_n82), .A2(
        DP_OP_425J2_127_3477_n110), .A3(DP_OP_425J2_127_3477_n85), .Y(n1368)
         );
  AO22X1_HVT U2445 ( .A1(DP_OP_422J2_124_3477_n1291), .A2(
        DP_OP_422J2_124_3477_n1289), .A3(n1369), .A4(
        DP_OP_422J2_124_3477_n1458), .Y(DP_OP_422J2_124_3477_n1256) );
  OR2X1_HVT U2446 ( .A1(DP_OP_422J2_124_3477_n1291), .A2(
        DP_OP_422J2_124_3477_n1289), .Y(n1369) );
  XOR3X2_HVT U2447 ( .A1(DP_OP_422J2_124_3477_n1289), .A2(
        DP_OP_422J2_124_3477_n1291), .A3(DP_OP_422J2_124_3477_n1458), .Y(
        DP_OP_422J2_124_3477_n1257) );
  NAND2X0_HVT U2448 ( .A1(conv2_sum_b[25]), .A2(n1903), .Y(n2044) );
  NBUFFX2_HVT U2449 ( .A(conv_weight_box[64]), .Y(n1372) );
  AND2X1_HVT U2450 ( .A1(conv_weight_box[64]), .A2(src_window[227]), .Y(
        DP_OP_424J2_126_3477_n2466) );
  AND2X1_HVT U2451 ( .A1(n1372), .A2(src_window[230]), .Y(
        DP_OP_424J2_126_3477_n2463) );
  AND2X1_HVT U2452 ( .A1(n1372), .A2(src_window[226]), .Y(
        DP_OP_424J2_126_3477_n2467) );
  AND2X1_HVT U2453 ( .A1(n1372), .A2(src_window[225]), .Y(
        DP_OP_424J2_126_3477_n2468) );
  AND2X1_HVT U2454 ( .A1(n1372), .A2(src_window[224]), .Y(
        DP_OP_424J2_126_3477_n2469) );
  AND2X1_HVT U2455 ( .A1(n1372), .A2(src_window[269]), .Y(
        DP_OP_423J2_125_3477_n2464) );
  AND2X1_HVT U2456 ( .A1(n1372), .A2(src_window[229]), .Y(
        DP_OP_424J2_126_3477_n2464) );
  NAND2X0_HVT U2457 ( .A1(n1372), .A2(src_window[231]), .Y(
        DP_OP_424J2_126_3477_n2462) );
  AND2X1_HVT U2458 ( .A1(n1372), .A2(src_window[228]), .Y(
        DP_OP_424J2_126_3477_n2465) );
  AO22X1_HVT U2459 ( .A1(n1373), .A2(n1718), .A3(n1719), .A4(
        DP_OP_424J2_126_3477_n2922), .Y(DP_OP_424J2_126_3477_n1682) );
  XOR3X2_HVT U2460 ( .A1(n1716), .A2(n1373), .A3(n1717), .Y(
        DP_OP_424J2_126_3477_n1683) );
  OR2X1_HVT U2461 ( .A1(DP_OP_424J2_126_3477_n2976), .A2(
        DP_OP_424J2_126_3477_n2979), .Y(n1720) );
  NAND2X0_HVT U2462 ( .A1(n1418), .A2(conv1_sram_rdata_weight[70]), .Y(n1375)
         );
  INVX2_HVT U2463 ( .A(conv2_sram_rdata_weight[70]), .Y(n1376) );
  AO22X1_HVT U2464 ( .A1(n1377), .A2(n1777), .A3(n1778), .A4(
        DP_OP_425J2_127_3477_n2922), .Y(DP_OP_425J2_127_3477_n1682) );
  XOR3X2_HVT U2465 ( .A1(n1775), .A2(n1377), .A3(n1776), .Y(
        DP_OP_425J2_127_3477_n1683) );
  OR2X2_HVT U2466 ( .A1(n857), .A2(n1871), .Y(n1384) );
  OR2X1_HVT U2467 ( .A1(n1853), .A2(DP_OP_422J2_124_3477_n2), .Y(n1379) );
  AND2X1_HVT U2468 ( .A1(conv_weight_box[43]), .A2(src_window[204]), .Y(
        DP_OP_422J2_124_3477_n2289) );
  AND2X1_HVT U2469 ( .A1(conv_weight_box[43]), .A2(src_window[205]), .Y(
        DP_OP_422J2_124_3477_n2288) );
  NAND2X0_HVT U2470 ( .A1(conv_weight_box[43]), .A2(src_window[207]), .Y(
        DP_OP_422J2_124_3477_n2286) );
  AND2X1_HVT U2471 ( .A1(conv_weight_box[43]), .A2(src_window[206]), .Y(
        DP_OP_422J2_124_3477_n2287) );
  AND2X1_HVT U2472 ( .A1(conv_weight_box[43]), .A2(src_window[203]), .Y(
        DP_OP_422J2_124_3477_n2290) );
  AND2X1_HVT U2473 ( .A1(conv_weight_box[43]), .A2(src_window[202]), .Y(
        DP_OP_422J2_124_3477_n2291) );
  AND2X1_HVT U2474 ( .A1(conv_weight_box[43]), .A2(src_window[201]), .Y(
        DP_OP_422J2_124_3477_n2292) );
  AND2X4_HVT U2475 ( .A1(conv_weight_box[43]), .A2(src_window[200]), .Y(
        DP_OP_422J2_124_3477_n2293) );
  AO21X1_HVT U2476 ( .A1(DP_OP_422J2_124_3477_n4), .A2(n1592), .A3(n1525), .Y(
        n1385) );
  AND2X1_HVT U2477 ( .A1(conv_weight_box[30]), .A2(src_window[114]), .Y(
        DP_OP_424J2_126_3477_n2219) );
  NAND2X0_HVT U2478 ( .A1(n1390), .A2(n1389), .Y(n1393) );
  AND3X1_HVT U2479 ( .A1(n1394), .A2(n1609), .A3(n1622), .Y(n1389) );
  AND2X1_HVT U2480 ( .A1(n1656), .A2(n1655), .Y(n1394) );
  NAND2X0_HVT U2481 ( .A1(n1633), .A2(DP_OP_423J2_125_3477_n237), .Y(n1391) );
  NBUFFX2_HVT U2482 ( .A(conv_weight_box[30]), .Y(n1395) );
  NAND2X0_HVT U2483 ( .A1(conv_weight_box[30]), .A2(src_window[111]), .Y(
        DP_OP_425J2_127_3477_n2214) );
  AND2X1_HVT U2484 ( .A1(n1395), .A2(src_window[106]), .Y(
        DP_OP_425J2_127_3477_n2219) );
  AND2X1_HVT U2485 ( .A1(n1395), .A2(src_window[110]), .Y(
        DP_OP_425J2_127_3477_n2215) );
  AND2X1_HVT U2486 ( .A1(n1395), .A2(src_window[109]), .Y(
        DP_OP_425J2_127_3477_n2216) );
  AND2X1_HVT U2487 ( .A1(n1395), .A2(src_window[105]), .Y(
        DP_OP_425J2_127_3477_n2220) );
  AND2X1_HVT U2488 ( .A1(n1395), .A2(src_window[108]), .Y(
        DP_OP_425J2_127_3477_n2217) );
  AND2X1_HVT U2489 ( .A1(n1395), .A2(src_window[107]), .Y(
        DP_OP_425J2_127_3477_n2218) );
  INVX2_HVT U2490 ( .A(n1960), .Y(n1483) );
  MUX21X2_HVT U2491 ( .A1(conv2_sum_b[17]), .A2(conv2_sum_a[17]), .S0(n1483), 
        .Y(tmp_big1[17]) );
  INVX4_HVT U2492 ( .A(conv_weight_box[51]), .Y(DP_OP_423J2_125_3477_n2409) );
  MUX21X2_HVT U2493 ( .A1(conv2_sram_rdata_weight[43]), .A2(
        conv1_sram_rdata_weight[43]), .S0(n619), .Y(conv_weight_box[29]) );
  MUX21X2_HVT U2494 ( .A1(conv2_sram_rdata_weight[32]), .A2(
        conv1_sram_rdata_weight[32]), .S0(n619), .Y(conv_weight_box[21]) );
  NAND2X0_HVT U2495 ( .A1(n1290), .A2(n2107), .Y(n2060) );
  XOR3X2_HVT U2496 ( .A1(DP_OP_423J2_125_3477_n1047), .A2(
        DP_OP_423J2_125_3477_n1232), .A3(DP_OP_423J2_125_3477_n1230), .Y(
        DP_OP_423J2_125_3477_n1033) );
  NAND2X0_HVT U2497 ( .A1(DP_OP_423J2_125_3477_n1047), .A2(
        DP_OP_423J2_125_3477_n1230), .Y(n1397) );
  NAND2X0_HVT U2498 ( .A1(DP_OP_423J2_125_3477_n1232), .A2(
        DP_OP_423J2_125_3477_n1230), .Y(n1398) );
  NAND2X0_HVT U2499 ( .A1(DP_OP_423J2_125_3477_n1232), .A2(
        DP_OP_423J2_125_3477_n1047), .Y(n1399) );
  NAND3X0_HVT U2500 ( .A1(n1399), .A2(n1398), .A3(n1397), .Y(
        DP_OP_423J2_125_3477_n1032) );
  OR2X4_HVT U2501 ( .A1(DP_OP_423J2_125_3477_n335), .A2(n909), .Y(n1677) );
  MUX21X2_HVT U2502 ( .A1(conv2_sum_b[7]), .A2(conv2_sum_a[7]), .S0(n1974), 
        .Y(tmp_big1[7]) );
  INVX1_HVT U2503 ( .A(n1534), .Y(n1575) );
  XNOR2X2_HVT U2504 ( .A1(n1831), .A2(DP_OP_425J2_127_3477_n15), .Y(
        n_conv2_sum_d[22]) );
  INVX1_HVT U2505 ( .A(n2177), .Y(n1401) );
  OR2X2_HVT U2506 ( .A1(DP_OP_424J2_126_3477_n2933), .A2(n1432), .Y(n1514) );
  MUX21X2_HVT U2507 ( .A1(conv2_sum_b[6]), .A2(conv2_sum_a[6]), .S0(n1502), 
        .Y(tmp_big1[6]) );
  XOR3X2_HVT U2508 ( .A1(DP_OP_422J2_124_3477_n1258), .A2(
        DP_OP_422J2_124_3477_n1077), .A3(DP_OP_422J2_124_3477_n1254), .Y(
        DP_OP_422J2_124_3477_n1051) );
  NAND2X0_HVT U2509 ( .A1(DP_OP_422J2_124_3477_n1258), .A2(
        DP_OP_422J2_124_3477_n1254), .Y(n1402) );
  NAND2X0_HVT U2510 ( .A1(DP_OP_422J2_124_3477_n1077), .A2(
        DP_OP_422J2_124_3477_n1254), .Y(n1403) );
  NAND2X0_HVT U2511 ( .A1(DP_OP_422J2_124_3477_n1077), .A2(
        DP_OP_422J2_124_3477_n1258), .Y(n1404) );
  NAND3X0_HVT U2512 ( .A1(n1404), .A2(n1403), .A3(n1402), .Y(
        DP_OP_422J2_124_3477_n1050) );
  XOR3X2_HVT U2513 ( .A1(DP_OP_422J2_124_3477_n1656), .A2(
        DP_OP_422J2_124_3477_n1654), .A3(DP_OP_422J2_124_3477_n1652), .Y(
        DP_OP_422J2_124_3477_n1461) );
  NAND2X0_HVT U2514 ( .A1(DP_OP_422J2_124_3477_n1656), .A2(
        DP_OP_422J2_124_3477_n1654), .Y(n1405) );
  NAND2X0_HVT U2515 ( .A1(DP_OP_422J2_124_3477_n1652), .A2(
        DP_OP_422J2_124_3477_n1654), .Y(n1406) );
  NAND2X0_HVT U2516 ( .A1(DP_OP_422J2_124_3477_n1652), .A2(
        DP_OP_422J2_124_3477_n1656), .Y(n1407) );
  NAND3X0_HVT U2517 ( .A1(n1407), .A2(n1406), .A3(n1405), .Y(
        DP_OP_422J2_124_3477_n1460) );
  MUX21X1_HVT U2518 ( .A1(conv2_sum_a[8]), .A2(conv2_sum_b[8]), .S0(n1960), 
        .Y(tmp_big1[8]) );
  NOR2X0_HVT U2519 ( .A1(DP_OP_423J2_125_3477_n2669), .A2(n1400), .Y(
        DP_OP_423J2_125_3477_n2645) );
  NOR2X0_HVT U2520 ( .A1(DP_OP_423J2_125_3477_n2668), .A2(n1400), .Y(
        DP_OP_423J2_125_3477_n2644) );
  NOR2X0_HVT U2521 ( .A1(DP_OP_423J2_125_3477_n2269), .A2(
        DP_OP_424J2_126_3477_n2671), .Y(DP_OP_425J2_127_3477_n2641) );
  NOR2X2_HVT U2522 ( .A1(DP_OP_424J2_126_3477_n2576), .A2(n1400), .Y(
        DP_OP_423J2_125_3477_n2640) );
  OR2X1_HVT U2523 ( .A1(DP_OP_425J2_127_3477_n2801), .A2(n1443), .Y(
        DP_OP_425J2_127_3477_n2769) );
  NOR2X0_HVT U2524 ( .A1(DP_OP_422J2_124_3477_n2794), .A2(n1443), .Y(
        DP_OP_422J2_124_3477_n2762) );
  OR2X1_HVT U2525 ( .A1(DP_OP_422J2_124_3477_n2797), .A2(n1443), .Y(
        DP_OP_422J2_124_3477_n2765) );
  OR2X1_HVT U2526 ( .A1(DP_OP_425J2_127_3477_n2799), .A2(n1443), .Y(
        DP_OP_425J2_127_3477_n2767) );
  MUX21X2_HVT U2527 ( .A1(conv2_sram_rdata_weight[41]), .A2(
        conv1_sram_rdata_weight[41]), .S0(n843), .Y(conv_weight_box[27]) );
  OR2X4_HVT U2528 ( .A1(DP_OP_422J2_124_3477_n2354), .A2(n1400), .Y(
        DP_OP_423J2_125_3477_n2638) );
  OR2X4_HVT U2529 ( .A1(DP_OP_423J2_125_3477_n2750), .A2(
        DP_OP_425J2_127_3477_n2671), .Y(DP_OP_424J2_126_3477_n2638) );
  NOR2X4_HVT U2530 ( .A1(DP_OP_423J2_125_3477_n2667), .A2(n1400), .Y(
        DP_OP_423J2_125_3477_n2643) );
  NOR2X2_HVT U2531 ( .A1(DP_OP_422J2_124_3477_n2800), .A2(n1400), .Y(
        DP_OP_425J2_127_3477_n2644) );
  NOR2X4_HVT U2532 ( .A1(DP_OP_424J2_126_3477_n2575), .A2(
        DP_OP_425J2_127_3477_n2671), .Y(DP_OP_423J2_125_3477_n2639) );
  NOR2X2_HVT U2533 ( .A1(DP_OP_422J2_124_3477_n2795), .A2(
        DP_OP_425J2_127_3477_n2671), .Y(DP_OP_425J2_127_3477_n2639) );
  NOR2X4_HVT U2534 ( .A1(DP_OP_425J2_127_3477_n2404), .A2(n1400), .Y(
        DP_OP_424J2_126_3477_n2644) );
  INVX4_HVT U2535 ( .A(n1960), .Y(n1502) );
  NOR2X2_HVT U2536 ( .A1(DP_OP_423J2_125_3477_n2887), .A2(
        DP_OP_423J2_125_3477_n2892), .Y(DP_OP_423J2_125_3477_n2871) );
  OR2X2_HVT U2537 ( .A1(DP_OP_423J2_125_3477_n2053), .A2(n30), .Y(
        DP_OP_423J2_125_3477_n2021) );
  OR2X2_HVT U2538 ( .A1(DP_OP_425J2_127_3477_n2796), .A2(
        DP_OP_424J2_126_3477_n2802), .Y(DP_OP_425J2_127_3477_n2764) );
  XOR3X2_HVT U2539 ( .A1(DP_OP_423J2_125_3477_n1248), .A2(
        DP_OP_423J2_125_3477_n1246), .A3(DP_OP_423J2_125_3477_n1250), .Y(
        DP_OP_423J2_125_3477_n1045) );
  NAND2X0_HVT U2540 ( .A1(DP_OP_423J2_125_3477_n1248), .A2(
        DP_OP_423J2_125_3477_n1250), .Y(n1408) );
  NAND2X0_HVT U2541 ( .A1(DP_OP_423J2_125_3477_n1246), .A2(
        DP_OP_423J2_125_3477_n1250), .Y(n1409) );
  NAND2X0_HVT U2542 ( .A1(DP_OP_423J2_125_3477_n1246), .A2(
        DP_OP_423J2_125_3477_n1248), .Y(n1410) );
  NAND3X0_HVT U2543 ( .A1(n1410), .A2(n1409), .A3(n1408), .Y(
        DP_OP_423J2_125_3477_n1044) );
  MUX21X2_HVT U2544 ( .A1(conv2_sram_rdata_weight[10]), .A2(
        conv1_sram_rdata_weight[10]), .S0(n241), .Y(conv_weight_box[6]) );
  MUX21X2_HVT U2545 ( .A1(conv2_sram_rdata_weight[97]), .A2(
        conv1_sram_rdata_weight[97]), .S0(n241), .Y(conv_weight_box[67]) );
  MUX21X2_HVT U2546 ( .A1(conv2_sram_rdata_weight[79]), .A2(
        conv1_sram_rdata_weight[79]), .S0(n241), .Y(conv_weight_box[52]) );
  MUX21X2_HVT U2547 ( .A1(conv2_sram_rdata_weight[46]), .A2(
        conv1_sram_rdata_weight[46]), .S0(n241), .Y(conv_weight_box[31]) );
  NOR2X0_HVT U2548 ( .A1(DP_OP_423J2_125_3477_n2317), .A2(
        DP_OP_425J2_127_3477_n2320), .Y(DP_OP_423J2_125_3477_n2301) );
  NAND2X0_HVT U2549 ( .A1(DP_OP_422J2_124_3477_n2156), .A2(
        DP_OP_422J2_124_3477_n2860), .Y(n1411) );
  NAND2X0_HVT U2550 ( .A1(DP_OP_422J2_124_3477_n2163), .A2(
        DP_OP_422J2_124_3477_n2860), .Y(n1412) );
  NAND2X0_HVT U2551 ( .A1(DP_OP_422J2_124_3477_n2163), .A2(
        DP_OP_422J2_124_3477_n2156), .Y(n1413) );
  NAND3X0_HVT U2552 ( .A1(n1413), .A2(n1412), .A3(n1411), .Y(
        DP_OP_422J2_124_3477_n970) );
  NBUFFX2_HVT U2553 ( .A(DP_OP_422J2_124_3477_n654), .Y(n1414) );
  NOR2X2_HVT U2554 ( .A1(DP_OP_422J2_124_3477_n2884), .A2(
        DP_OP_424J2_126_3477_n2891), .Y(DP_OP_422J2_124_3477_n2860) );
  NOR2X2_HVT U2555 ( .A1(DP_OP_422J2_124_3477_n2179), .A2(
        DP_OP_425J2_127_3477_n2188), .Y(DP_OP_422J2_124_3477_n2163) );
  NAND2X0_HVT U2556 ( .A1(DP_OP_425J2_127_3477_n2864), .A2(
        DP_OP_425J2_127_3477_n2871), .Y(n1415) );
  NAND2X0_HVT U2557 ( .A1(DP_OP_425J2_127_3477_n2350), .A2(
        DP_OP_425J2_127_3477_n2871), .Y(n1416) );
  NAND2X0_HVT U2558 ( .A1(DP_OP_425J2_127_3477_n2350), .A2(
        DP_OP_425J2_127_3477_n2864), .Y(n1417) );
  NAND3X0_HVT U2559 ( .A1(n1417), .A2(n1416), .A3(n1415), .Y(
        DP_OP_425J2_127_3477_n1676) );
  OR2X2_HVT U2560 ( .A1(DP_OP_425J2_127_3477_n2882), .A2(
        DP_OP_423J2_125_3477_n2892), .Y(DP_OP_425J2_127_3477_n2866) );
  MUX21X2_HVT U2561 ( .A1(conv2_sram_rdata_weight[53]), .A2(
        conv1_sram_rdata_weight[53]), .S0(n843), .Y(conv_weight_box[37]) );
  MUX21X2_HVT U2562 ( .A1(conv2_sram_rdata_weight[84]), .A2(
        conv1_sram_rdata_weight[84]), .S0(n843), .Y(conv_weight_box[57]) );
  OR2X2_HVT U2563 ( .A1(DP_OP_425J2_127_3477_n418), .A2(
        DP_OP_425J2_127_3477_n373), .Y(n1770) );
  XOR3X2_HVT U2564 ( .A1(DP_OP_425J2_127_3477_n424), .A2(
        DP_OP_425J2_127_3477_n379), .A3(DP_OP_425J2_127_3477_n422), .Y(
        DP_OP_425J2_127_3477_n375) );
  INVX4_HVT U2565 ( .A(n1503), .Y(n1481) );
  INVX2_HVT U2566 ( .A(n1505), .Y(n1503) );
  INVX2_HVT U2567 ( .A(conv_weight_box[27]), .Y(DP_OP_425J2_127_3477_n2848) );
  MUX21X2_HVT U2568 ( .A1(conv2_sum_b[15]), .A2(conv2_sum_a[15]), .S0(n1429), 
        .Y(tmp_big1[15]) );
  MUX21X2_HVT U2569 ( .A1(conv2_sum_b[24]), .A2(conv2_sum_a[24]), .S0(n1974), 
        .Y(tmp_big1[24]) );
  XOR3X2_HVT U2570 ( .A1(DP_OP_424J2_126_3477_n379), .A2(
        DP_OP_424J2_126_3477_n424), .A3(DP_OP_424J2_126_3477_n422), .Y(
        DP_OP_424J2_126_3477_n375) );
  INVX1_HVT U2571 ( .A(n1713), .Y(DP_OP_424J2_126_3477_n236) );
  NOR2X2_HVT U2572 ( .A1(DP_OP_425J2_127_3477_n2756), .A2(
        DP_OP_422J2_124_3477_n2759), .Y(DP_OP_425J2_127_3477_n2732) );
  NOR2X2_HVT U2573 ( .A1(DP_OP_423J2_125_3477_n2756), .A2(
        DP_OP_422J2_124_3477_n2759), .Y(DP_OP_423J2_125_3477_n2732) );
  NAND2X0_HVT U2574 ( .A1(n1639), .A2(DP_OP_423J2_125_3477_n17), .Y(n1419) );
  NAND2X0_HVT U2575 ( .A1(n1424), .A2(n1637), .Y(n1420) );
  NAND2X0_HVT U2576 ( .A1(n1419), .A2(n1420), .Y(n_conv2_sum_b[20]) );
  XOR3X2_HVT U2577 ( .A1(DP_OP_423J2_125_3477_n2520), .A2(
        DP_OP_423J2_125_3477_n2513), .A3(DP_OP_423J2_125_3477_n2733), .Y(
        DP_OP_423J2_125_3477_n1805) );
  NAND2X0_HVT U2578 ( .A1(DP_OP_423J2_125_3477_n2520), .A2(
        DP_OP_423J2_125_3477_n2733), .Y(n1421) );
  NAND2X0_HVT U2579 ( .A1(DP_OP_423J2_125_3477_n2513), .A2(
        DP_OP_423J2_125_3477_n2733), .Y(n1422) );
  NAND2X0_HVT U2580 ( .A1(DP_OP_423J2_125_3477_n2513), .A2(
        DP_OP_423J2_125_3477_n2520), .Y(n1423) );
  NAND3X0_HVT U2581 ( .A1(n1423), .A2(n1422), .A3(n1421), .Y(
        DP_OP_423J2_125_3477_n1804) );
  MUX21X2_HVT U2582 ( .A1(tmp_big2[21]), .A2(tmp_big1[21]), .S0(n1504), .Y(
        data_out[21]) );
  NBUFFX4_HVT U2583 ( .A(n1505), .Y(n1504) );
  MUX21X2_HVT U2584 ( .A1(tmp_big2[28]), .A2(tmp_big1[28]), .S0(n1967), .Y(
        data_out[28]) );
  INVX2_HVT U2585 ( .A(conv_weight_box[20]), .Y(DP_OP_424J2_126_3477_n2143) );
  NOR2X4_HVT U2586 ( .A1(DP_OP_423J2_125_3477_n2006), .A2(
        DP_OP_422J2_124_3477_n2935), .Y(DP_OP_425J2_127_3477_n2906) );
  NOR2X4_HVT U2587 ( .A1(DP_OP_424J2_126_3477_n2092), .A2(
        DP_OP_422J2_124_3477_n2935), .Y(DP_OP_425J2_127_3477_n2904) );
  OR2X2_HVT U2588 ( .A1(DP_OP_422J2_124_3477_n2533), .A2(n1334), .Y(
        DP_OP_422J2_124_3477_n2501) );
  NOR2X2_HVT U2589 ( .A1(DP_OP_422J2_124_3477_n2530), .A2(n1362), .Y(
        DP_OP_422J2_124_3477_n2498) );
  OR2X2_HVT U2590 ( .A1(DP_OP_422J2_124_3477_n2536), .A2(n1335), .Y(
        DP_OP_422J2_124_3477_n2504) );
  INVX8_HVT U2591 ( .A(n1425), .Y(DP_OP_422J2_124_3477_n2) );
  MUX21X2_HVT U2592 ( .A1(conv2_sram_rdata_weight[7]), .A2(
        conv1_sram_rdata_weight[7]), .S0(n241), .Y(conv_weight_box[4]) );
  AND2X1_HVT U2593 ( .A1(conv_weight_box[15]), .A2(src_window[96]), .Y(n1640)
         );
  AND2X1_HVT U2594 ( .A1(conv_weight_box[15]), .A2(src_window[104]), .Y(n1547)
         );
  MUX21X2_HVT U2595 ( .A1(conv2_sram_rdata_weight[23]), .A2(
        conv1_sram_rdata_weight[23]), .S0(n241), .Y(conv_weight_box[15]) );
  OR2X2_HVT U2596 ( .A1(DP_OP_425J2_127_3477_n2933), .A2(
        DP_OP_423J2_125_3477_n2010), .Y(DP_OP_423J2_125_3477_n1977) );
  OR2X4_HVT U2597 ( .A1(DP_OP_423J2_125_3477_n2005), .A2(
        DP_OP_423J2_125_3477_n2010), .Y(DP_OP_423J2_125_3477_n1973) );
  OR2X4_HVT U2598 ( .A1(DP_OP_423J2_125_3477_n2006), .A2(
        DP_OP_423J2_125_3477_n2010), .Y(DP_OP_423J2_125_3477_n1974) );
  OR2X4_HVT U2599 ( .A1(DP_OP_423J2_125_3477_n2003), .A2(
        DP_OP_423J2_125_3477_n2010), .Y(DP_OP_423J2_125_3477_n1971) );
  INVX1_HVT U2600 ( .A(n2059), .Y(n2107) );
  INVX2_HVT U2601 ( .A(conv_weight_box[45]), .Y(DP_OP_422J2_124_3477_n2715) );
  NOR2X2_HVT U2602 ( .A1(DP_OP_422J2_124_3477_n2490), .A2(n772), .Y(
        DP_OP_423J2_125_3477_n2510) );
  NOR2X2_HVT U2603 ( .A1(DP_OP_422J2_124_3477_n2488), .A2(n772), .Y(
        DP_OP_423J2_125_3477_n2508) );
  NOR2X2_HVT U2604 ( .A1(DP_OP_422J2_124_3477_n2489), .A2(n772), .Y(
        DP_OP_423J2_125_3477_n2509) );
  NOR2X2_HVT U2605 ( .A1(DP_OP_422J2_124_3477_n2491), .A2(n772), .Y(
        DP_OP_423J2_125_3477_n2511) );
  MUX21X2_HVT U2606 ( .A1(conv2_sum_b[2]), .A2(conv2_sum_a[2]), .S0(n1502), 
        .Y(tmp_big1[2]) );
  INVX1_HVT U2607 ( .A(conv_weight_box[52]), .Y(n1426) );
  INVX2_HVT U2608 ( .A(conv_weight_box[52]), .Y(n1433) );
  INVX2_HVT U2609 ( .A(conv_weight_box[16]), .Y(DP_OP_423J2_125_3477_n2936) );
  OR2X4_HVT U2610 ( .A1(DP_OP_422J2_124_3477_n2006), .A2(
        DP_OP_424J2_126_3477_n2010), .Y(DP_OP_422J2_124_3477_n1974) );
  NOR2X4_HVT U2611 ( .A1(DP_OP_424J2_126_3477_n2185), .A2(
        DP_OP_425J2_127_3477_n2980), .Y(DP_OP_422J2_124_3477_n2961) );
  NOR2X2_HVT U2612 ( .A1(DP_OP_424J2_126_3477_n2005), .A2(n1431), .Y(
        DP_OP_424J2_126_3477_n1997) );
  NOR2X4_HVT U2613 ( .A1(DP_OP_423J2_125_3477_n2005), .A2(
        DP_OP_422J2_124_3477_n2013), .Y(DP_OP_423J2_125_3477_n1997) );
  NOR2X2_HVT U2614 ( .A1(DP_OP_424J2_126_3477_n3057), .A2(
        DP_OP_422J2_124_3477_n2013), .Y(DP_OP_425J2_127_3477_n1995) );
  OR2X4_HVT U2615 ( .A1(DP_OP_424J2_126_3477_n2002), .A2(
        DP_OP_422J2_124_3477_n2013), .Y(DP_OP_424J2_126_3477_n1994) );
  OR2X4_HVT U2616 ( .A1(DP_OP_424J2_126_3477_n2090), .A2(
        DP_OP_422J2_124_3477_n2935), .Y(DP_OP_425J2_127_3477_n2902) );
  OR2X4_HVT U2617 ( .A1(DP_OP_422J2_124_3477_n2926), .A2(
        DP_OP_422J2_124_3477_n2935), .Y(DP_OP_422J2_124_3477_n2902) );
  NOR2X4_HVT U2618 ( .A1(DP_OP_423J2_125_3477_n2003), .A2(
        DP_OP_422J2_124_3477_n2935), .Y(DP_OP_425J2_127_3477_n2903) );
  NOR2X2_HVT U2619 ( .A1(DP_OP_424J2_126_3477_n2929), .A2(
        DP_OP_422J2_124_3477_n2935), .Y(DP_OP_424J2_126_3477_n2905) );
  OR2X4_HVT U2620 ( .A1(DP_OP_422J2_124_3477_n2795), .A2(
        DP_OP_423J2_125_3477_n2802), .Y(DP_OP_422J2_124_3477_n2763) );
  OR2X4_HVT U2621 ( .A1(DP_OP_422J2_124_3477_n2970), .A2(
        DP_OP_424J2_126_3477_n2980), .Y(DP_OP_422J2_124_3477_n2954) );
  NOR2X2_HVT U2622 ( .A1(DP_OP_422J2_124_3477_n2975), .A2(
        DP_OP_425J2_127_3477_n2980), .Y(DP_OP_422J2_124_3477_n2959) );
  NOR2X2_HVT U2623 ( .A1(DP_OP_422J2_124_3477_n2973), .A2(
        DP_OP_425J2_127_3477_n2980), .Y(DP_OP_422J2_124_3477_n2957) );
  NOR2X2_HVT U2624 ( .A1(DP_OP_422J2_124_3477_n2971), .A2(
        DP_OP_424J2_126_3477_n2980), .Y(DP_OP_422J2_124_3477_n2955) );
  OR2X2_HVT U2625 ( .A1(DP_OP_425J2_127_3477_n2002), .A2(
        DP_OP_422J2_124_3477_n2013), .Y(DP_OP_425J2_127_3477_n1994) );
  INVX2_HVT U2626 ( .A(N7), .Y(n1531) );
  INVX4_HVT U2627 ( .A(conv_weight_box[2]), .Y(DP_OP_423J2_125_3477_n2013) );
  AND2X4_HVT U2628 ( .A1(conv_weight_box[2]), .A2(src_window[65]), .Y(
        DP_OP_422J2_124_3477_n2000) );
  MUX21X2_HVT U2629 ( .A1(conv2_sram_rdata_weight[83]), .A2(
        conv1_sram_rdata_weight[83]), .S0(n240), .Y(conv_weight_box[56]) );
  INVX1_HVT U2630 ( .A(conv_weight_box[35]), .Y(DP_OP_424J2_126_3477_n2802) );
  INVX1_HVT U2631 ( .A(conv_weight_box[26]), .Y(n1428) );
  INVX2_HVT U2632 ( .A(conv_weight_box[17]), .Y(n1432) );
  INVX2_HVT U2633 ( .A(conv_weight_box[56]), .Y(DP_OP_422J2_124_3477_n2626) );
  INVX2_HVT U2634 ( .A(n1960), .Y(n1429) );
  INVX2_HVT U2635 ( .A(n1960), .Y(n1430) );
  INVX8_HVT U2636 ( .A(DP_OP_422J2_124_3477_n2), .Y(n1484) );
  XOR3X2_HVT U2637 ( .A1(DP_OP_424J2_126_3477_n1455), .A2(
        DP_OP_424J2_126_3477_n1453), .A3(DP_OP_424J2_126_3477_n1449), .Y(
        DP_OP_424J2_126_3477_n1425) );
  XOR3X2_HVT U2638 ( .A1(DP_OP_422J2_124_3477_n656), .A2(
        DP_OP_422J2_124_3477_n523), .A3(n1414), .Y(DP_OP_422J2_124_3477_n517)
         );
  XOR3X2_HVT U2639 ( .A1(DP_OP_425J2_127_3477_n1455), .A2(
        DP_OP_425J2_127_3477_n1453), .A3(DP_OP_425J2_127_3477_n1449), .Y(
        DP_OP_425J2_127_3477_n1425) );
  AND2X4_HVT U2640 ( .A1(conv_weight_box[17]), .A2(src_window[110]), .Y(
        DP_OP_423J2_125_3477_n2903) );
  AND2X4_HVT U2641 ( .A1(conv_weight_box[17]), .A2(src_window[106]), .Y(
        DP_OP_423J2_125_3477_n2907) );
  AND2X4_HVT U2642 ( .A1(conv_weight_box[17]), .A2(src_window[107]), .Y(
        DP_OP_423J2_125_3477_n2906) );
  AND2X4_HVT U2643 ( .A1(conv_weight_box[17]), .A2(src_window[108]), .Y(
        DP_OP_423J2_125_3477_n2905) );
  AND2X4_HVT U2644 ( .A1(conv_weight_box[17]), .A2(src_window[109]), .Y(
        DP_OP_423J2_125_3477_n2904) );
  AND2X4_HVT U2645 ( .A1(conv_weight_box[17]), .A2(src_window[105]), .Y(
        DP_OP_423J2_125_3477_n2908) );
  AND2X4_HVT U2646 ( .A1(conv_weight_box[17]), .A2(src_window[104]), .Y(
        DP_OP_423J2_125_3477_n2909) );
  INVX1_HVT U2647 ( .A(conv_weight_box[2]), .Y(n1431) );
  NOR2X2_HVT U2648 ( .A1(DP_OP_424J2_126_3477_n2667), .A2(
        DP_OP_422J2_124_3477_n2759), .Y(DP_OP_423J2_125_3477_n2731) );
  NAND2X0_HVT U2649 ( .A1(n1792), .A2(n1774), .Y(DP_OP_425J2_127_3477_n233) );
  INVX0_HVT U2650 ( .A(DP_OP_423J2_125_3477_n71), .Y(DP_OP_423J2_125_3477_n69)
         );
  OAI21X1_HVT U2651 ( .A1(DP_OP_425J2_127_3477_n261), .A2(
        DP_OP_425J2_127_3477_n259), .A3(DP_OP_425J2_127_3477_n260), .Y(n1796)
         );
  INVX1_HVT U2652 ( .A(n1533), .Y(n1437) );
  INVX2_HVT U2653 ( .A(n1960), .Y(n1974) );
  MUX21X1_HVT U2654 ( .A1(conv2_sum_b[1]), .A2(conv2_sum_a[1]), .S0(n488), .Y(
        tmp_big1[1]) );
  OR2X1_HVT U2655 ( .A1(DP_OP_422J2_124_3477_n3015), .A2(n1507), .Y(
        DP_OP_422J2_124_3477_n2983) );
  OR2X1_HVT U2656 ( .A1(DP_OP_422J2_124_3477_n2838), .A2(
        DP_OP_422J2_124_3477_n2847), .Y(DP_OP_422J2_124_3477_n2814) );
  OR2X1_HVT U2657 ( .A1(DP_OP_422J2_124_3477_n2179), .A2(
        DP_OP_424J2_126_3477_n2758), .Y(DP_OP_424J2_126_3477_n2719) );
  OR2X1_HVT U2658 ( .A1(DP_OP_424J2_126_3477_n2574), .A2(n671), .Y(
        DP_OP_424J2_126_3477_n2550) );
  OR2X1_HVT U2659 ( .A1(DP_OP_423J2_125_3477_n2090), .A2(n621), .Y(
        DP_OP_423J2_125_3477_n2082) );
  OR2X1_HVT U2660 ( .A1(DP_OP_423J2_125_3477_n3056), .A2(n621), .Y(
        DP_OP_425J2_127_3477_n2082) );
  OR2X2_HVT U2661 ( .A1(DP_OP_422J2_124_3477_n2091), .A2(n1439), .Y(
        DP_OP_422J2_124_3477_n2059) );
  OR2X1_HVT U2662 ( .A1(DP_OP_423J2_125_3477_n2227), .A2(
        DP_OP_425J2_127_3477_n2230), .Y(DP_OP_423J2_125_3477_n2195) );
  OR2X1_HVT U2663 ( .A1(DP_OP_422J2_124_3477_n2223), .A2(
        DP_OP_422J2_124_3477_n2230), .Y(DP_OP_422J2_124_3477_n2191) );
  NOR2X0_HVT U2664 ( .A1(DP_OP_423J2_125_3477_n3057), .A2(n621), .Y(
        DP_OP_425J2_127_3477_n2083) );
  NOR2X1_HVT U2665 ( .A1(DP_OP_424J2_126_3477_n3020), .A2(
        DP_OP_425J2_127_3477_n3023), .Y(DP_OP_424J2_126_3477_n2996) );
  OR2X1_HVT U2666 ( .A1(DP_OP_425J2_127_3477_n2843), .A2(n1439), .Y(
        DP_OP_423J2_125_3477_n2063) );
  OR2X1_HVT U2667 ( .A1(DP_OP_423J2_125_3477_n3059), .A2(n1439), .Y(
        DP_OP_425J2_127_3477_n2061) );
  OR2X1_HVT U2668 ( .A1(DP_OP_424J2_126_3477_n2005), .A2(n1507), .Y(
        DP_OP_425J2_127_3477_n2985) );
  OR2X1_HVT U2669 ( .A1(DP_OP_423J2_125_3477_n2750), .A2(
        DP_OP_422J2_124_3477_n2409), .Y(DP_OP_425J2_127_3477_n2390) );
  OR2X1_HVT U2670 ( .A1(DP_OP_424J2_126_3477_n2269), .A2(
        DP_OP_422J2_124_3477_n2758), .Y(DP_OP_425J2_127_3477_n2721) );
  OR2X1_HVT U2671 ( .A1(DP_OP_425J2_127_3477_n2048), .A2(n1507), .Y(
        DP_OP_424J2_126_3477_n2984) );
  OR2X1_HVT U2672 ( .A1(DP_OP_425J2_127_3477_n2046), .A2(n1475), .Y(
        DP_OP_425J2_127_3477_n2038) );
  NOR2X1_HVT U2673 ( .A1(DP_OP_425J2_127_3477_n2053), .A2(n1475), .Y(
        DP_OP_425J2_127_3477_n2045) );
  OR2X1_HVT U2674 ( .A1(DP_OP_425J2_127_3477_n2933), .A2(n1439), .Y(
        DP_OP_424J2_126_3477_n2065) );
  NOR2X1_HVT U2675 ( .A1(DP_OP_425J2_127_3477_n2712), .A2(n1440), .Y(
        DP_OP_425J2_127_3477_n2688) );
  OR2X1_HVT U2676 ( .A1(DP_OP_423J2_125_3477_n2008), .A2(
        DP_OP_423J2_125_3477_n2010), .Y(DP_OP_423J2_125_3477_n1976) );
  NOR2X1_HVT U2677 ( .A1(DP_OP_424J2_126_3477_n2927), .A2(
        DP_OP_425J2_127_3477_n2935), .Y(DP_OP_424J2_126_3477_n2903) );
  OR2X1_HVT U2678 ( .A1(DP_OP_424J2_126_3477_n2003), .A2(
        DP_OP_424J2_126_3477_n2010), .Y(DP_OP_424J2_126_3477_n1971) );
  NOR2X1_HVT U2679 ( .A1(DP_OP_423J2_125_3477_n2447), .A2(n789), .Y(
        DP_OP_423J2_125_3477_n2423) );
  OR2X1_HVT U2680 ( .A1(DP_OP_423J2_125_3477_n2708), .A2(
        DP_OP_422J2_124_3477_n2626), .Y(DP_OP_424J2_126_3477_n2588) );
  NOR2X1_HVT U2681 ( .A1(DP_OP_423J2_125_3477_n2053), .A2(
        DP_OP_425J2_127_3477_n2057), .Y(DP_OP_423J2_125_3477_n2045) );
  OR2X1_HVT U2682 ( .A1(DP_OP_423J2_125_3477_n3063), .A2(n1439), .Y(
        DP_OP_425J2_127_3477_n2065) );
  OR2X1_HVT U2683 ( .A1(DP_OP_422J2_124_3477_n2751), .A2(n1433), .Y(
        DP_OP_424J2_126_3477_n2367) );
  OR2X1_HVT U2684 ( .A1(DP_OP_423J2_125_3477_n2003), .A2(
        DP_OP_425J2_127_3477_n2098), .Y(DP_OP_424J2_126_3477_n2059) );
  OR2X1_HVT U2685 ( .A1(DP_OP_422J2_124_3477_n2090), .A2(n1438), .Y(
        DP_OP_424J2_126_3477_n2814) );
  OR2X1_HVT U2686 ( .A1(DP_OP_424J2_126_3477_n2619), .A2(n1331), .Y(
        DP_OP_424J2_126_3477_n2587) );
  OR2X1_HVT U2687 ( .A1(DP_OP_422J2_124_3477_n2002), .A2(n1432), .Y(
        DP_OP_424J2_126_3477_n2902) );
  OR2X1_HVT U2688 ( .A1(DP_OP_425J2_127_3477_n2574), .A2(n671), .Y(
        DP_OP_425J2_127_3477_n2550) );
  OR2X1_HVT U2689 ( .A1(DP_OP_424J2_126_3477_n2928), .A2(n1507), .Y(
        DP_OP_423J2_125_3477_n2984) );
  OR2X1_HVT U2690 ( .A1(DP_OP_425J2_127_3477_n2448), .A2(
        DP_OP_422J2_124_3477_n2626), .Y(DP_OP_424J2_126_3477_n2592) );
  OR2X1_HVT U2691 ( .A1(DP_OP_424J2_126_3477_n2090), .A2(n621), .Y(
        DP_OP_424J2_126_3477_n2082) );
  OR2X1_HVT U2692 ( .A1(DP_OP_422J2_124_3477_n2618), .A2(
        DP_OP_423J2_125_3477_n2452), .Y(DP_OP_423J2_125_3477_n2426) );
  OR2X1_HVT U2693 ( .A1(DP_OP_424J2_126_3477_n2267), .A2(
        DP_OP_423J2_125_3477_n2758), .Y(DP_OP_425J2_127_3477_n2719) );
  OR2X1_HVT U2694 ( .A1(DP_OP_422J2_124_3477_n2442), .A2(n671), .Y(
        DP_OP_423J2_125_3477_n2550) );
  OR2X1_HVT U2695 ( .A1(DP_OP_425J2_127_3477_n2138), .A2(n1507), .Y(
        DP_OP_423J2_125_3477_n2986) );
  OR2X2_HVT U2696 ( .A1(DP_OP_423J2_125_3477_n3060), .A2(n1439), .Y(
        DP_OP_425J2_127_3477_n2062) );
  OR2X1_HVT U2697 ( .A1(DP_OP_422J2_124_3477_n3058), .A2(
        DP_OP_423J2_125_3477_n2010), .Y(DP_OP_423J2_125_3477_n1972) );
  OR2X1_HVT U2698 ( .A1(DP_OP_424J2_126_3477_n3060), .A2(
        DP_OP_425J2_127_3477_n2010), .Y(DP_OP_425J2_127_3477_n1974) );
  OR2X1_HVT U2699 ( .A1(DP_OP_422J2_124_3477_n2270), .A2(n1433), .Y(
        DP_OP_425J2_127_3477_n2370) );
  OR2X2_HVT U2700 ( .A1(DP_OP_423J2_125_3477_n3057), .A2(n1439), .Y(
        DP_OP_425J2_127_3477_n2059) );
  OR2X1_HVT U2701 ( .A1(DP_OP_422J2_124_3477_n2093), .A2(n1439), .Y(
        DP_OP_422J2_124_3477_n2061) );
  OR2X1_HVT U2702 ( .A1(DP_OP_423J2_125_3477_n2931), .A2(n1439), .Y(
        DP_OP_422J2_124_3477_n2063) );
  OR2X1_HVT U2703 ( .A1(DP_OP_424J2_126_3477_n2095), .A2(n1439), .Y(
        DP_OP_424J2_126_3477_n2063) );
  NOR2X0_HVT U2704 ( .A1(DP_OP_422J2_124_3477_n2839), .A2(n1440), .Y(
        DP_OP_425J2_127_3477_n2683) );
  OR2X2_HVT U2705 ( .A1(DP_OP_425J2_127_3477_n2839), .A2(n1439), .Y(
        DP_OP_423J2_125_3477_n2059) );
  OR2X1_HVT U2706 ( .A1(DP_OP_423J2_125_3477_n2706), .A2(n1497), .Y(
        DP_OP_423J2_125_3477_n2682) );
  NOR2X1_HVT U2707 ( .A1(DP_OP_425J2_127_3477_n2359), .A2(n1440), .Y(
        DP_OP_424J2_126_3477_n2687) );
  OR2X1_HVT U2708 ( .A1(DP_OP_424J2_126_3477_n2574), .A2(
        DP_OP_422J2_124_3477_n2585), .Y(DP_OP_424J2_126_3477_n2566) );
  OR2X1_HVT U2709 ( .A1(DP_OP_423J2_125_3477_n2222), .A2(n1497), .Y(
        DP_OP_425J2_127_3477_n2682) );
  OR2X1_HVT U2710 ( .A1(DP_OP_424J2_126_3477_n3057), .A2(
        DP_OP_425J2_127_3477_n2010), .Y(DP_OP_425J2_127_3477_n1971) );
  OR2X1_HVT U2711 ( .A1(DP_OP_424J2_126_3477_n2004), .A2(n1507), .Y(
        DP_OP_425J2_127_3477_n2984) );
  NOR2X0_HVT U2712 ( .A1(DP_OP_422J2_124_3477_n2839), .A2(
        DP_OP_425J2_127_3477_n2231), .Y(DP_OP_423J2_125_3477_n2199) );
  NOR2X1_HVT U2713 ( .A1(DP_OP_424J2_126_3477_n2927), .A2(
        DP_OP_424J2_126_3477_n3023), .Y(DP_OP_423J2_125_3477_n2991) );
  OR2X1_HVT U2714 ( .A1(DP_OP_425J2_127_3477_n2092), .A2(n1439), .Y(
        DP_OP_425J2_127_3477_n2060) );
  NOR2X0_HVT U2715 ( .A1(DP_OP_422J2_124_3477_n2840), .A2(n1438), .Y(
        DP_OP_422J2_124_3477_n2816) );
  NOR2X0_HVT U2716 ( .A1(DP_OP_422J2_124_3477_n2622), .A2(n789), .Y(
        DP_OP_423J2_125_3477_n2422) );
  OR2X1_HVT U2717 ( .A1(DP_OP_422J2_124_3477_n2751), .A2(
        DP_OP_422J2_124_3477_n2758), .Y(DP_OP_422J2_124_3477_n2719) );
  OR2X1_HVT U2718 ( .A1(DP_OP_424J2_126_3477_n2622), .A2(
        DP_OP_422J2_124_3477_n2626), .Y(DP_OP_424J2_126_3477_n2590) );
  NOR2X0_HVT U2719 ( .A1(DP_OP_424J2_126_3477_n2003), .A2(
        DP_OP_423J2_125_3477_n2013), .Y(DP_OP_424J2_126_3477_n1995) );
  OR2X1_HVT U2720 ( .A1(DP_OP_422J2_124_3477_n2181), .A2(
        DP_OP_424J2_126_3477_n2758), .Y(DP_OP_424J2_126_3477_n2721) );
  OR2X1_HVT U2721 ( .A1(DP_OP_422J2_124_3477_n2574), .A2(n671), .Y(
        DP_OP_422J2_124_3477_n2550) );
  OR2X1_HVT U2722 ( .A1(DP_OP_422J2_124_3477_n3060), .A2(
        DP_OP_425J2_127_3477_n2098), .Y(DP_OP_424J2_126_3477_n2062) );
  OR2X1_HVT U2723 ( .A1(DP_OP_422J2_124_3477_n2882), .A2(
        DP_OP_423J2_125_3477_n2892), .Y(DP_OP_422J2_124_3477_n2866) );
  OR2X1_HVT U2724 ( .A1(DP_OP_425J2_127_3477_n2050), .A2(n1507), .Y(
        DP_OP_424J2_126_3477_n2986) );
  OR2X1_HVT U2725 ( .A1(DP_OP_422J2_124_3477_n3021), .A2(n1507), .Y(
        DP_OP_422J2_124_3477_n2989) );
  OR2X1_HVT U2726 ( .A1(DP_OP_422J2_124_3477_n2092), .A2(n1439), .Y(
        DP_OP_422J2_124_3477_n2060) );
  OR2X1_HVT U2727 ( .A1(DP_OP_422J2_124_3477_n2754), .A2(n1433), .Y(
        DP_OP_424J2_126_3477_n2370) );
  OR2X1_HVT U2728 ( .A1(DP_OP_424J2_126_3477_n2006), .A2(
        DP_OP_424J2_126_3477_n2010), .Y(DP_OP_424J2_126_3477_n1974) );
  OR2X1_HVT U2729 ( .A1(DP_OP_424J2_126_3477_n2136), .A2(n1507), .Y(
        DP_OP_422J2_124_3477_n2984) );
  OR2X1_HVT U2730 ( .A1(DP_OP_422J2_124_3477_n2313), .A2(
        DP_OP_422J2_124_3477_n2626), .Y(DP_OP_424J2_126_3477_n2589) );
  NOR2X1_HVT U2731 ( .A1(DP_OP_423J2_125_3477_n2798), .A2(n1440), .Y(
        DP_OP_424J2_126_3477_n2686) );
  NOR2X0_HVT U2732 ( .A1(DP_OP_422J2_124_3477_n2223), .A2(n597), .Y(
        DP_OP_424J2_126_3477_n2699) );
  OR2X1_HVT U2733 ( .A1(DP_OP_423J2_125_3477_n2794), .A2(n597), .Y(
        DP_OP_424J2_126_3477_n2698) );
  NOR2X0_HVT U2734 ( .A1(DP_OP_422J2_124_3477_n2619), .A2(
        DP_OP_422J2_124_3477_n2629), .Y(DP_OP_422J2_124_3477_n2611) );
  OR2X1_HVT U2735 ( .A1(DP_OP_422J2_124_3477_n2618), .A2(
        DP_OP_422J2_124_3477_n2629), .Y(DP_OP_422J2_124_3477_n2610) );
  INVX1_HVT U2736 ( .A(conv_weight_box[18]), .Y(n1442) );
  NOR2X1_HVT U2737 ( .A1(DP_OP_423J2_125_3477_n2795), .A2(
        DP_OP_422J2_124_3477_n2803), .Y(DP_OP_423J2_125_3477_n2771) );
  NOR2X0_HVT U2738 ( .A1(DP_OP_423J2_125_3477_n2619), .A2(
        DP_OP_423J2_125_3477_n2629), .Y(DP_OP_423J2_125_3477_n2611) );
  INVX2_HVT U2739 ( .A(conv_weight_box[28]), .Y(n1438) );
  INVX1_HVT U2740 ( .A(conv_weight_box[54]), .Y(n1441) );
  OR2X1_HVT U2741 ( .A1(DP_OP_423J2_125_3477_n2310), .A2(
        DP_OP_423J2_125_3477_n2321), .Y(DP_OP_423J2_125_3477_n2302) );
  NOR2X0_HVT U2742 ( .A1(DP_OP_422J2_124_3477_n2795), .A2(n1444), .Y(
        DP_OP_422J2_124_3477_n2771) );
  OR2X2_HVT U2743 ( .A1(DP_OP_422J2_124_3477_n2794), .A2(
        DP_OP_422J2_124_3477_n2803), .Y(DP_OP_422J2_124_3477_n2770) );
  OR2X1_HVT U2744 ( .A1(DP_OP_423J2_125_3477_n2618), .A2(
        DP_OP_423J2_125_3477_n2629), .Y(DP_OP_423J2_125_3477_n2610) );
  INVX1_HVT U2745 ( .A(conv_weight_box[33]), .Y(DP_OP_422J2_124_3477_n2805) );
  INVX1_HVT U2746 ( .A(conv_weight_box[33]), .Y(DP_OP_423J2_125_3477_n2805) );
  MUX21X1_HVT U2747 ( .A1(conv2_sram_rdata_weight[81]), .A2(
        conv1_sram_rdata_weight[81]), .S0(n241), .Y(conv_weight_box[54]) );
  INVX1_HVT U2748 ( .A(srstn), .Y(n1434) );
  INVX0_HVT U2749 ( .A(src_window[168]), .Y(DP_OP_422J2_124_3477_n2801) );
  INVX2_HVT U2750 ( .A(n1614), .Y(n1436) );
  INVX0_HVT U2751 ( .A(DP_OP_423J2_125_3477_n222), .Y(n1523) );
  INVX0_HVT U2752 ( .A(n1623), .Y(n1630) );
  INVX0_HVT U2753 ( .A(DP_OP_423J2_125_3477_n220), .Y(
        DP_OP_423J2_125_3477_n222) );
  NAND2X0_HVT U2754 ( .A1(n1733), .A2(n1715), .Y(DP_OP_424J2_126_3477_n233) );
  INVX0_HVT U2755 ( .A(DP_OP_422J2_124_3477_n141), .Y(
        DP_OP_422J2_124_3477_n139) );
  MUX21X1_HVT U2756 ( .A1(tmp_big2[23]), .A2(tmp_big1[23]), .S0(n1482), .Y(
        data_out[23]) );
  MUX21X1_HVT U2757 ( .A1(tmp_big2[27]), .A2(tmp_big1[27]), .S0(n1967), .Y(
        data_out[27]) );
  INVX0_HVT U2758 ( .A(DP_OP_424J2_126_3477_n109), .Y(
        DP_OP_424J2_126_3477_n107) );
  INVX0_HVT U2759 ( .A(DP_OP_425J2_127_3477_n109), .Y(
        DP_OP_425J2_127_3477_n107) );
  INVX0_HVT U2760 ( .A(n1625), .Y(DP_OP_423J2_125_3477_n141) );
  INVX0_HVT U2761 ( .A(DP_OP_423J2_125_3477_n122), .Y(n1628) );
  INVX0_HVT U2762 ( .A(DP_OP_425J2_127_3477_n160), .Y(
        DP_OP_425J2_127_3477_n158) );
  INVX0_HVT U2763 ( .A(n913), .Y(DP_OP_422J2_124_3477_n241) );
  INVX0_HVT U2764 ( .A(DP_OP_422J2_124_3477_n160), .Y(
        DP_OP_422J2_124_3477_n158) );
  INVX0_HVT U2765 ( .A(DP_OP_422J2_124_3477_n161), .Y(
        DP_OP_422J2_124_3477_n159) );
  INVX0_HVT U2766 ( .A(DP_OP_423J2_125_3477_n161), .Y(
        DP_OP_423J2_125_3477_n159) );
  INVX0_HVT U2767 ( .A(DP_OP_424J2_126_3477_n140), .Y(
        DP_OP_424J2_126_3477_n138) );
  INVX0_HVT U2768 ( .A(DP_OP_422J2_124_3477_n140), .Y(
        DP_OP_422J2_124_3477_n138) );
  INVX0_HVT U2769 ( .A(DP_OP_422J2_124_3477_n109), .Y(
        DP_OP_422J2_124_3477_n107) );
  INVX0_HVT U2770 ( .A(DP_OP_422J2_124_3477_n177), .Y(
        DP_OP_422J2_124_3477_n179) );
  MUX21X1_HVT U2771 ( .A1(tmp_big2[8]), .A2(tmp_big1[8]), .S0(n1482), .Y(
        data_out[8]) );
  INVX0_HVT U2772 ( .A(DP_OP_423J2_125_3477_n140), .Y(
        DP_OP_423J2_125_3477_n138) );
  INVX0_HVT U2773 ( .A(DP_OP_423J2_125_3477_n160), .Y(
        DP_OP_423J2_125_3477_n158) );
  INVX0_HVT U2774 ( .A(DP_OP_423J2_125_3477_n109), .Y(
        DP_OP_423J2_125_3477_n107) );
  INVX0_HVT U2775 ( .A(DP_OP_423J2_125_3477_n110), .Y(
        DP_OP_423J2_125_3477_n108) );
  INVX0_HVT U2776 ( .A(DP_OP_425J2_127_3477_n50), .Y(n1803) );
  NBUFFX2_HVT U2777 ( .A(n1481), .Y(n1967) );
  INVX0_HVT U2778 ( .A(DP_OP_425J2_127_3477_n176), .Y(
        DP_OP_425J2_127_3477_n178) );
  INVX0_HVT U2779 ( .A(DP_OP_424J2_126_3477_n176), .Y(
        DP_OP_424J2_126_3477_n178) );
  INVX0_HVT U2780 ( .A(DP_OP_424J2_126_3477_n50), .Y(n1739) );
  INVX0_HVT U2781 ( .A(DP_OP_422J2_124_3477_n190), .Y(
        DP_OP_422J2_124_3477_n188) );
  INVX0_HVT U2782 ( .A(n1655), .Y(DP_OP_423J2_125_3477_n214) );
  INVX0_HVT U2783 ( .A(DP_OP_425J2_127_3477_n56), .Y(DP_OP_425J2_127_3477_n54)
         );
  INVX0_HVT U2784 ( .A(DP_OP_422J2_124_3477_n189), .Y(
        DP_OP_422J2_124_3477_n187) );
  INVX0_HVT U2785 ( .A(DP_OP_422J2_124_3477_n57), .Y(DP_OP_422J2_124_3477_n55)
         );
  INVX0_HVT U2786 ( .A(DP_OP_422J2_124_3477_n56), .Y(DP_OP_422J2_124_3477_n54)
         );
  INVX0_HVT U2787 ( .A(DP_OP_424J2_126_3477_n189), .Y(
        DP_OP_424J2_126_3477_n187) );
  INVX0_HVT U2788 ( .A(DP_OP_425J2_127_3477_n189), .Y(
        DP_OP_425J2_127_3477_n187) );
  INVX2_HVT U2789 ( .A(n1503), .Y(n1482) );
  INVX0_HVT U2790 ( .A(DP_OP_423J2_125_3477_n177), .Y(
        DP_OP_423J2_125_3477_n179) );
  INVX1_HVT U2791 ( .A(N9), .Y(n2178) );
  INVX0_HVT U2792 ( .A(DP_OP_423J2_125_3477_n176), .Y(
        DP_OP_423J2_125_3477_n178) );
  INVX0_HVT U2793 ( .A(DP_OP_424J2_126_3477_n56), .Y(DP_OP_424J2_126_3477_n54)
         );
  INVX0_HVT U2794 ( .A(DP_OP_423J2_125_3477_n67), .Y(n1619) );
  AND2X1_HVT U2795 ( .A1(DP_OP_424J2_126_3477_n287), .A2(
        DP_OP_424J2_126_3477_n22), .Y(n1726) );
  INVX0_HVT U2796 ( .A(n1745), .Y(DP_OP_424J2_126_3477_n214) );
  INVX0_HVT U2797 ( .A(DP_OP_425J2_127_3477_n226), .Y(n1817) );
  INVX0_HVT U2798 ( .A(DP_OP_424J2_126_3477_n22), .Y(n1724) );
  INVX0_HVT U2799 ( .A(DP_OP_423J2_125_3477_n190), .Y(
        DP_OP_423J2_125_3477_n188) );
  INVX0_HVT U2800 ( .A(DP_OP_424J2_126_3477_n201), .Y(n1723) );
  INVX0_HVT U2801 ( .A(n1814), .Y(DP_OP_425J2_127_3477_n214) );
  AND2X1_HVT U2802 ( .A1(DP_OP_425J2_127_3477_n287), .A2(
        DP_OP_425J2_127_3477_n22), .Y(n1785) );
  INVX0_HVT U2803 ( .A(DP_OP_425J2_127_3477_n201), .Y(n1782) );
  INVX0_HVT U2804 ( .A(n1772), .Y(DP_OP_425J2_127_3477_n236) );
  INVX0_HVT U2805 ( .A(DP_OP_423J2_125_3477_n57), .Y(DP_OP_423J2_125_3477_n55)
         );
  INVX0_HVT U2806 ( .A(DP_OP_423J2_125_3477_n56), .Y(DP_OP_423J2_125_3477_n54)
         );
  INVX0_HVT U2807 ( .A(DP_OP_423J2_125_3477_n189), .Y(
        DP_OP_423J2_125_3477_n187) );
  INVX0_HVT U2808 ( .A(DP_OP_422J2_124_3477_n245), .Y(n1578) );
  INVX1_HVT U2809 ( .A(DP_OP_424J2_126_3477_n202), .Y(
        DP_OP_424J2_126_3477_n287) );
  INVX0_HVT U2810 ( .A(DP_OP_425J2_127_3477_n22), .Y(n1783) );
  INVX1_HVT U2811 ( .A(DP_OP_425J2_127_3477_n202), .Y(
        DP_OP_425J2_127_3477_n287) );
  OR2X1_HVT U2812 ( .A1(DP_OP_422J2_124_3477_n335), .A2(
        DP_OP_422J2_124_3477_n340), .Y(n1592) );
  XOR3X1_HVT U2813 ( .A1(DP_OP_424J2_126_3477_n423), .A2(
        DP_OP_424J2_126_3477_n514), .A3(DP_OP_424J2_126_3477_n421), .Y(
        DP_OP_424J2_126_3477_n419) );
  INVX0_HVT U2814 ( .A(n1971), .Y(n1968) );
  INVX0_HVT U2815 ( .A(DP_OP_425J2_127_3477_n252), .Y(n1798) );
  INVX0_HVT U2816 ( .A(DP_OP_424J2_126_3477_n252), .Y(n1738) );
  INVX0_HVT U2817 ( .A(DP_OP_423J2_125_3477_n182), .Y(
        DP_OP_423J2_125_3477_n285) );
  INVX0_HVT U2818 ( .A(DP_OP_425J2_127_3477_n182), .Y(
        DP_OP_425J2_127_3477_n285) );
  INVX0_HVT U2819 ( .A(DP_OP_425J2_127_3477_n257), .Y(
        DP_OP_425J2_127_3477_n255) );
  INVX0_HVT U2820 ( .A(DP_OP_422J2_124_3477_n182), .Y(
        DP_OP_422J2_124_3477_n285) );
  INVX0_HVT U2821 ( .A(DP_OP_424J2_126_3477_n182), .Y(
        DP_OP_424J2_126_3477_n285) );
  FADDX1_HVT U2822 ( .A(DP_OP_422J2_124_3477_n667), .B(
        DP_OP_422J2_124_3477_n834), .CI(DP_OP_422J2_124_3477_n665), .CO(
        DP_OP_422J2_124_3477_n656), .S(DP_OP_422J2_124_3477_n657) );
  INVX0_HVT U2823 ( .A(n2144), .Y(n1941) );
  INVX0_HVT U2824 ( .A(n2116), .Y(n2169) );
  INVX0_HVT U2825 ( .A(n2145), .Y(n1945) );
  FADDX1_HVT U2826 ( .A(DP_OP_423J2_125_3477_n536), .B(
        DP_OP_423J2_125_3477_n443), .CI(DP_OP_423J2_125_3477_n534), .CO(
        DP_OP_423J2_125_3477_n432), .S(DP_OP_423J2_125_3477_n433) );
  INVX0_HVT U2827 ( .A(DP_OP_424J2_126_3477_n111), .Y(n1742) );
  INVX0_HVT U2828 ( .A(DP_OP_422J2_124_3477_n144), .Y(
        DP_OP_422J2_124_3477_n142) );
  INVX0_HVT U2829 ( .A(DP_OP_422J2_124_3477_n96), .Y(DP_OP_422J2_124_3477_n94)
         );
  INVX0_HVT U2830 ( .A(DP_OP_422J2_124_3477_n127), .Y(
        DP_OP_422J2_124_3477_n125) );
  INVX0_HVT U2831 ( .A(DP_OP_422J2_124_3477_n126), .Y(
        DP_OP_422J2_124_3477_n124) );
  INVX0_HVT U2832 ( .A(DP_OP_424J2_126_3477_n144), .Y(
        DP_OP_424J2_126_3477_n142) );
  INVX0_HVT U2833 ( .A(tmp_big1[18]), .Y(n2158) );
  INVX0_HVT U2834 ( .A(n2156), .Y(tmp_big1[13]) );
  AOI22X1_HVT U2835 ( .A1(tmp_big2[14]), .A2(n1976), .A3(tmp_big2[15]), .A4(
        n2157), .Y(n2135) );
  INVX0_HVT U2836 ( .A(tmp_big1[28]), .Y(n2165) );
  INVX0_HVT U2837 ( .A(tmp_big2[25]), .Y(n1926) );
  INVX0_HVT U2838 ( .A(tmp_big1[30]), .Y(n2168) );
  INVX0_HVT U2839 ( .A(n2164), .Y(tmp_big1[27]) );
  INVX0_HVT U2840 ( .A(tmp_big1[12]), .Y(n2155) );
  INVX0_HVT U2841 ( .A(tmp_big1[20]), .Y(n2160) );
  INVX0_HVT U2842 ( .A(DP_OP_422J2_124_3477_n269), .Y(DP_OP_422J2_124_3477_n5)
         );
  INVX0_HVT U2843 ( .A(DP_OP_425J2_127_3477_n111), .Y(n1811) );
  INVX0_HVT U2844 ( .A(DP_OP_422J2_124_3477_n51), .Y(DP_OP_422J2_124_3477_n272) );
  INVX0_HVT U2845 ( .A(DP_OP_423J2_125_3477_n269), .Y(DP_OP_423J2_125_3477_n5)
         );
  INVX0_HVT U2846 ( .A(DP_OP_422J2_124_3477_n133), .Y(
        DP_OP_422J2_124_3477_n280) );
  INVX0_HVT U2847 ( .A(DP_OP_422J2_124_3477_n153), .Y(
        DP_OP_422J2_124_3477_n282) );
  INVX0_HVT U2848 ( .A(DP_OP_422J2_124_3477_n166), .Y(
        DP_OP_422J2_124_3477_n283) );
  INVX0_HVT U2849 ( .A(DP_OP_422J2_124_3477_n102), .Y(
        DP_OP_422J2_124_3477_n277) );
  INVX0_HVT U2850 ( .A(DP_OP_425J2_127_3477_n269), .Y(DP_OP_425J2_127_3477_n5)
         );
  INVX0_HVT U2851 ( .A(DP_OP_422J2_124_3477_n171), .Y(
        DP_OP_422J2_124_3477_n284) );
  INVX0_HVT U2852 ( .A(DP_OP_422J2_124_3477_n97), .Y(DP_OP_422J2_124_3477_n276) );
  INVX0_HVT U2853 ( .A(DP_OP_422J2_124_3477_n128), .Y(
        DP_OP_422J2_124_3477_n279) );
  INVX0_HVT U2854 ( .A(DP_OP_422J2_124_3477_n148), .Y(
        DP_OP_422J2_124_3477_n281) );
  INVX0_HVT U2855 ( .A(DP_OP_424J2_126_3477_n19), .Y(n1477) );
  INVX0_HVT U2856 ( .A(DP_OP_422J2_124_3477_n77), .Y(DP_OP_422J2_124_3477_n274) );
  INVX0_HVT U2857 ( .A(DP_OP_425J2_127_3477_n13), .Y(n1824) );
  INVX0_HVT U2858 ( .A(DP_OP_425J2_127_3477_n144), .Y(
        DP_OP_425J2_127_3477_n142) );
  INVX0_HVT U2859 ( .A(DP_OP_425J2_127_3477_n77), .Y(DP_OP_425J2_127_3477_n274) );
  INVX0_HVT U2860 ( .A(DP_OP_424J2_126_3477_n269), .Y(DP_OP_424J2_126_3477_n5)
         );
  INVX0_HVT U2861 ( .A(DP_OP_424J2_126_3477_n13), .Y(n1749) );
  INVX0_HVT U2862 ( .A(DP_OP_424J2_126_3477_n17), .Y(n1753) );
  INVX0_HVT U2863 ( .A(DP_OP_424J2_126_3477_n171), .Y(
        DP_OP_424J2_126_3477_n284) );
  NAND2X0_HVT U2864 ( .A1(DP_OP_424J2_126_3477_n283), .A2(
        DP_OP_424J2_126_3477_n167), .Y(DP_OP_424J2_126_3477_n19) );
  INVX0_HVT U2865 ( .A(DP_OP_424J2_126_3477_n51), .Y(DP_OP_424J2_126_3477_n272) );
  INVX0_HVT U2866 ( .A(DP_OP_424J2_126_3477_n77), .Y(DP_OP_424J2_126_3477_n274) );
  INVX0_HVT U2867 ( .A(tmp_big1[9]), .Y(n1979) );
  INVX0_HVT U2868 ( .A(DP_OP_423J2_125_3477_n144), .Y(
        DP_OP_423J2_125_3477_n142) );
  INVX0_HVT U2869 ( .A(DP_OP_423J2_125_3477_n77), .Y(DP_OP_423J2_125_3477_n274) );
  INVX0_HVT U2870 ( .A(DP_OP_423J2_125_3477_n51), .Y(DP_OP_423J2_125_3477_n272) );
  INVX0_HVT U2871 ( .A(tmp_big2[16]), .Y(n2151) );
  INVX0_HVT U2872 ( .A(DP_OP_425J2_127_3477_n17), .Y(n1828) );
  INVX0_HVT U2873 ( .A(DP_OP_425J2_127_3477_n19), .Y(n1453) );
  INVX0_HVT U2874 ( .A(DP_OP_425J2_127_3477_n126), .Y(
        DP_OP_425J2_127_3477_n124) );
  INVX0_HVT U2875 ( .A(DP_OP_423J2_125_3477_n126), .Y(
        DP_OP_423J2_125_3477_n124) );
  INVX0_HVT U2876 ( .A(DP_OP_423J2_125_3477_n127), .Y(
        DP_OP_423J2_125_3477_n125) );
  INVX0_HVT U2877 ( .A(DP_OP_424J2_126_3477_n126), .Y(
        DP_OP_424J2_126_3477_n124) );
  INVX0_HVT U2878 ( .A(DP_OP_423J2_125_3477_n96), .Y(DP_OP_423J2_125_3477_n94)
         );
  INVX0_HVT U2879 ( .A(DP_OP_424J2_126_3477_n166), .Y(
        DP_OP_424J2_126_3477_n283) );
  INVX0_HVT U2880 ( .A(DP_OP_425J2_127_3477_n51), .Y(DP_OP_425J2_127_3477_n272) );
  XOR3X1_HVT U2881 ( .A1(DP_OP_423J2_125_3477_n953), .A2(
        DP_OP_423J2_125_3477_n969), .A3(DP_OP_423J2_125_3477_n977), .Y(
        DP_OP_423J2_125_3477_n913) );
  XOR3X1_HVT U2882 ( .A1(DP_OP_422J2_124_3477_n1696), .A2(
        DP_OP_422J2_124_3477_n1662), .A3(DP_OP_422J2_124_3477_n1672), .Y(
        DP_OP_422J2_124_3477_n1495) );
  INVX0_HVT U2883 ( .A(DP_OP_423J2_125_3477_n97), .Y(DP_OP_423J2_125_3477_n276) );
  INVX0_HVT U2884 ( .A(DP_OP_423J2_125_3477_n102), .Y(
        DP_OP_423J2_125_3477_n277) );
  INVX1_HVT U2885 ( .A(n1961), .Y(n1994) );
  INVX0_HVT U2886 ( .A(DP_OP_423J2_125_3477_n128), .Y(
        DP_OP_423J2_125_3477_n279) );
  INVX0_HVT U2887 ( .A(DP_OP_423J2_125_3477_n133), .Y(
        DP_OP_423J2_125_3477_n280) );
  INVX0_HVT U2888 ( .A(DP_OP_425J2_127_3477_n166), .Y(
        DP_OP_425J2_127_3477_n283) );
  INVX0_HVT U2889 ( .A(DP_OP_423J2_125_3477_n148), .Y(
        DP_OP_423J2_125_3477_n281) );
  INVX0_HVT U2890 ( .A(DP_OP_425J2_127_3477_n97), .Y(DP_OP_425J2_127_3477_n276) );
  INVX0_HVT U2891 ( .A(DP_OP_425J2_127_3477_n102), .Y(
        DP_OP_425J2_127_3477_n277) );
  INVX0_HVT U2892 ( .A(DP_OP_424J2_126_3477_n97), .Y(DP_OP_424J2_126_3477_n276) );
  INVX0_HVT U2893 ( .A(DP_OP_424J2_126_3477_n102), .Y(
        DP_OP_424J2_126_3477_n277) );
  INVX0_HVT U2894 ( .A(DP_OP_424J2_126_3477_n128), .Y(
        DP_OP_424J2_126_3477_n279) );
  INVX0_HVT U2895 ( .A(DP_OP_425J2_127_3477_n128), .Y(
        DP_OP_425J2_127_3477_n279) );
  INVX0_HVT U2896 ( .A(DP_OP_424J2_126_3477_n133), .Y(
        DP_OP_424J2_126_3477_n280) );
  INVX0_HVT U2897 ( .A(DP_OP_424J2_126_3477_n148), .Y(
        DP_OP_424J2_126_3477_n281) );
  INVX0_HVT U2898 ( .A(DP_OP_425J2_127_3477_n133), .Y(
        DP_OP_425J2_127_3477_n280) );
  INVX0_HVT U2899 ( .A(DP_OP_424J2_126_3477_n153), .Y(
        DP_OP_424J2_126_3477_n282) );
  INVX0_HVT U2900 ( .A(DP_OP_425J2_127_3477_n148), .Y(
        DP_OP_425J2_127_3477_n281) );
  INVX0_HVT U2901 ( .A(DP_OP_423J2_125_3477_n153), .Y(
        DP_OP_423J2_125_3477_n282) );
  XOR3X1_HVT U2902 ( .A1(DP_OP_423J2_125_3477_n1668), .A2(
        DP_OP_423J2_125_3477_n1692), .A3(DP_OP_423J2_125_3477_n1694), .Y(
        DP_OP_423J2_125_3477_n1493) );
  INVX0_HVT U2903 ( .A(DP_OP_423J2_125_3477_n166), .Y(
        DP_OP_423J2_125_3477_n283) );
  INVX0_HVT U2904 ( .A(DP_OP_423J2_125_3477_n171), .Y(
        DP_OP_423J2_125_3477_n284) );
  INVX0_HVT U2905 ( .A(DP_OP_425J2_127_3477_n153), .Y(
        DP_OP_425J2_127_3477_n282) );
  INVX0_HVT U2906 ( .A(DP_OP_425J2_127_3477_n171), .Y(
        DP_OP_425J2_127_3477_n284) );
  INVX0_HVT U2907 ( .A(n1775), .Y(n1777) );
  INVX0_HVT U2908 ( .A(n1538), .Y(n1540) );
  XOR3X1_HVT U2909 ( .A1(DP_OP_422J2_124_3477_n2952), .A2(n1538), .A3(n1539), 
        .Y(DP_OP_422J2_124_3477_n1683) );
  INVX0_HVT U2910 ( .A(n1716), .Y(n1718) );
  XOR3X1_HVT U2911 ( .A1(DP_OP_422J2_124_3477_n2695), .A2(
        DP_OP_422J2_124_3477_n2688), .A3(DP_OP_422J2_124_3477_n1834), .Y(
        DP_OP_422J2_124_3477_n1661) );
  FADDX1_HVT U2912 ( .A(DP_OP_423J2_125_3477_n2087), .B(
        DP_OP_423J2_125_3477_n2080), .CI(DP_OP_423J2_125_3477_n2117), .CO(
        DP_OP_423J2_125_3477_n1828), .S(DP_OP_423J2_125_3477_n1829) );
  OR2X1_HVT U2913 ( .A1(DP_OP_425J2_127_3477_n2002), .A2(
        DP_OP_425J2_127_3477_n3066), .Y(DP_OP_424J2_126_3477_n3040) );
  NOR2X1_HVT U2914 ( .A1(DP_OP_424J2_126_3477_n2405), .A2(
        DP_OP_425J2_127_3477_n2409), .Y(DP_OP_424J2_126_3477_n2397) );
  OR2X1_HVT U2915 ( .A1(DP_OP_423J2_125_3477_n3061), .A2(
        DP_OP_423J2_125_3477_n2098), .Y(DP_OP_425J2_127_3477_n2063) );
  NOR2X0_HVT U2916 ( .A1(DP_OP_422J2_124_3477_n2715), .A2(
        DP_OP_424J2_126_3477_n2712), .Y(DP_OP_424J2_126_3477_n2688) );
  OR2X1_HVT U2917 ( .A1(DP_OP_424J2_126_3477_n2752), .A2(
        DP_OP_424J2_126_3477_n2758), .Y(DP_OP_424J2_126_3477_n2720) );
  OR2X1_HVT U2918 ( .A1(DP_OP_422J2_124_3477_n2838), .A2(
        DP_OP_422J2_124_3477_n2320), .Y(DP_OP_424J2_126_3477_n2294) );
  OR2X1_HVT U2919 ( .A1(DP_OP_425J2_127_3477_n2755), .A2(
        DP_OP_423J2_125_3477_n2758), .Y(DP_OP_425J2_127_3477_n2723) );
  OR2X1_HVT U2920 ( .A1(DP_OP_422J2_124_3477_n2398), .A2(n1487), .Y(
        DP_OP_424J2_126_3477_n2514) );
  OR2X1_HVT U2921 ( .A1(DP_OP_422J2_124_3477_n2618), .A2(n1499), .Y(
        DP_OP_422J2_124_3477_n2602) );
  NOR2X1_HVT U2922 ( .A1(DP_OP_423J2_125_3477_n2053), .A2(n1501), .Y(
        DP_OP_424J2_126_3477_n2133) );
  NOR2X1_HVT U2923 ( .A1(DP_OP_425J2_127_3477_n2933), .A2(n621), .Y(
        DP_OP_424J2_126_3477_n2089) );
  OR2X1_HVT U2924 ( .A1(DP_OP_422J2_124_3477_n2530), .A2(n1486), .Y(
        DP_OP_422J2_124_3477_n2514) );
  OR2X1_HVT U2925 ( .A1(DP_OP_424J2_126_3477_n2400), .A2(
        DP_OP_422J2_124_3477_n2758), .Y(DP_OP_422J2_124_3477_n2720) );
  OR2X1_HVT U2926 ( .A1(DP_OP_422J2_124_3477_n3056), .A2(
        DP_OP_423J2_125_3477_n3066), .Y(DP_OP_422J2_124_3477_n3040) );
  OR2X1_HVT U2927 ( .A1(DP_OP_422J2_124_3477_n2310), .A2(
        DP_OP_425J2_127_3477_n2320), .Y(DP_OP_422J2_124_3477_n2294) );
  OR2X1_HVT U2928 ( .A1(DP_OP_424J2_126_3477_n2794), .A2(
        DP_OP_423J2_125_3477_n2804), .Y(DP_OP_424J2_126_3477_n2778) );
  NOR2X0_HVT U2929 ( .A1(DP_OP_422J2_124_3477_n3014), .A2(n1507), .Y(
        DP_OP_422J2_124_3477_n2982) );
  OR2X1_HVT U2930 ( .A1(DP_OP_424J2_126_3477_n2092), .A2(
        DP_OP_425J2_127_3477_n2098), .Y(DP_OP_424J2_126_3477_n2060) );
  NOR2X0_HVT U2931 ( .A1(DP_OP_422J2_124_3477_n2090), .A2(
        DP_OP_425J2_127_3477_n2098), .Y(DP_OP_422J2_124_3477_n2058) );
  NOR2X1_HVT U2932 ( .A1(DP_OP_423J2_125_3477_n2625), .A2(n1499), .Y(
        DP_OP_423J2_125_3477_n2609) );
  NOR2X1_HVT U2933 ( .A1(DP_OP_423J2_125_3477_n3063), .A2(
        DP_OP_423J2_125_3477_n3066), .Y(DP_OP_423J2_125_3477_n3047) );
  NOR2X1_HVT U2934 ( .A1(DP_OP_424J2_126_3477_n2623), .A2(n1499), .Y(
        DP_OP_424J2_126_3477_n2607) );
  OR2X1_HVT U2935 ( .A1(DP_OP_423J2_125_3477_n2090), .A2(
        DP_OP_425J2_127_3477_n2847), .Y(DP_OP_425J2_127_3477_n2814) );
  OR2X1_HVT U2936 ( .A1(DP_OP_424J2_126_3477_n2002), .A2(
        DP_OP_422J2_124_3477_n3023), .Y(DP_OP_425J2_127_3477_n2990) );
  OR2X1_HVT U2937 ( .A1(DP_OP_422J2_124_3477_n2090), .A2(
        DP_OP_424J2_126_3477_n2231), .Y(DP_OP_425J2_127_3477_n2198) );
  OR2X1_HVT U2938 ( .A1(DP_OP_422J2_124_3477_n2222), .A2(
        DP_OP_425J2_127_3477_n2231), .Y(DP_OP_422J2_124_3477_n2198) );
  NOR2X0_HVT U2939 ( .A1(DP_OP_424J2_126_3477_n2002), .A2(
        DP_OP_424J2_126_3477_n2010), .Y(DP_OP_424J2_126_3477_n1970) );
  OR2X1_HVT U2940 ( .A1(DP_OP_422J2_124_3477_n3014), .A2(
        DP_OP_422J2_124_3477_n3023), .Y(DP_OP_422J2_124_3477_n2990) );
  NOR2X0_HVT U2941 ( .A1(DP_OP_422J2_124_3477_n2178), .A2(
        DP_OP_424J2_126_3477_n2758), .Y(DP_OP_424J2_126_3477_n2718) );
  NOR2X0_HVT U2942 ( .A1(DP_OP_424J2_126_3477_n2090), .A2(
        DP_OP_423J2_125_3477_n2098), .Y(DP_OP_424J2_126_3477_n2058) );
  NOR2X0_HVT U2943 ( .A1(DP_OP_425J2_127_3477_n2046), .A2(n1506), .Y(
        DP_OP_424J2_126_3477_n2982) );
  OR2X1_HVT U2944 ( .A1(DP_OP_424J2_126_3477_n2004), .A2(
        DP_OP_424J2_126_3477_n2010), .Y(DP_OP_424J2_126_3477_n1972) );
  NOR2X1_HVT U2945 ( .A1(DP_OP_422J2_124_3477_n2092), .A2(
        DP_OP_422J2_124_3477_n2231), .Y(DP_OP_425J2_127_3477_n2200) );
  OR2X1_HVT U2946 ( .A1(DP_OP_423J2_125_3477_n2794), .A2(
        DP_OP_422J2_124_3477_n2715), .Y(DP_OP_424J2_126_3477_n2682) );
  NOR2X1_HVT U2947 ( .A1(DP_OP_423J2_125_3477_n2399), .A2(n1487), .Y(
        DP_OP_425J2_127_3477_n2515) );
  OR2X1_HVT U2948 ( .A1(DP_OP_425J2_127_3477_n2046), .A2(
        DP_OP_425J2_127_3477_n3023), .Y(DP_OP_424J2_126_3477_n2990) );
  OR2X1_HVT U2949 ( .A1(DP_OP_423J2_125_3477_n2666), .A2(
        DP_OP_422J2_124_3477_n2585), .Y(n1716) );
  OR2X1_HVT U2950 ( .A1(DP_OP_424J2_126_3477_n2222), .A2(
        DP_OP_422J2_124_3477_n2231), .Y(DP_OP_424J2_126_3477_n2198) );
  OR2X1_HVT U2951 ( .A1(DP_OP_423J2_125_3477_n3021), .A2(
        DP_OP_423J2_125_3477_n3022), .Y(DP_OP_423J2_125_3477_n2989) );
  NOR2X1_HVT U2952 ( .A1(DP_OP_422J2_124_3477_n2224), .A2(
        DP_OP_425J2_127_3477_n2231), .Y(DP_OP_422J2_124_3477_n2200) );
  OR2X1_HVT U2953 ( .A1(DP_OP_423J2_125_3477_n2706), .A2(n1498), .Y(
        DP_OP_424J2_126_3477_n2602) );
  OR2X1_HVT U2954 ( .A1(DP_OP_424J2_126_3477_n2400), .A2(n1433), .Y(
        DP_OP_424J2_126_3477_n2368) );
  NOR2X1_HVT U2955 ( .A1(DP_OP_424J2_126_3477_n2004), .A2(
        DP_OP_425J2_127_3477_n3023), .Y(DP_OP_425J2_127_3477_n2992) );
  NOR2X1_HVT U2956 ( .A1(DP_OP_423J2_125_3477_n2311), .A2(n1498), .Y(
        DP_OP_425J2_127_3477_n2603) );
  NOR2X1_HVT U2957 ( .A1(DP_OP_424J2_126_3477_n3015), .A2(
        DP_OP_422J2_124_3477_n3023), .Y(DP_OP_424J2_126_3477_n2991) );
  NOR2X1_HVT U2958 ( .A1(DP_OP_422J2_124_3477_n2927), .A2(
        DP_OP_425J2_127_3477_n2231), .Y(DP_OP_424J2_126_3477_n2199) );
  OR2X1_HVT U2959 ( .A1(DP_OP_423J2_125_3477_n2798), .A2(
        DP_OP_423J2_125_3477_n2230), .Y(DP_OP_422J2_124_3477_n2194) );
  NOR2X1_HVT U2960 ( .A1(DP_OP_425J2_127_3477_n2576), .A2(n671), .Y(
        DP_OP_425J2_127_3477_n2552) );
  NOR2X0_HVT U2961 ( .A1(DP_OP_422J2_124_3477_n2750), .A2(n1433), .Y(
        DP_OP_424J2_126_3477_n2366) );
  NOR2X1_HVT U2962 ( .A1(DP_OP_422J2_124_3477_n2578), .A2(n671), .Y(
        DP_OP_422J2_124_3477_n2554) );
  NOR2X1_HVT U2963 ( .A1(DP_OP_422J2_124_3477_n3059), .A2(
        DP_OP_425J2_127_3477_n3066), .Y(DP_OP_422J2_124_3477_n3043) );
  OR2X1_HVT U2964 ( .A1(DP_OP_425J2_127_3477_n2801), .A2(
        DP_OP_422J2_124_3477_n2230), .Y(DP_OP_424J2_126_3477_n2197) );
  NOR2X1_HVT U2965 ( .A1(DP_OP_425J2_127_3477_n2049), .A2(
        DP_OP_425J2_127_3477_n3023), .Y(DP_OP_424J2_126_3477_n2993) );
  NOR2X1_HVT U2966 ( .A1(DP_OP_423J2_125_3477_n3061), .A2(n621), .Y(
        DP_OP_425J2_127_3477_n2087) );
  NOR2X1_HVT U2967 ( .A1(DP_OP_424J2_126_3477_n3019), .A2(n1475), .Y(
        DP_OP_425J2_127_3477_n2043) );
  OR2X1_HVT U2968 ( .A1(DP_OP_424J2_126_3477_n2005), .A2(
        DP_OP_424J2_126_3477_n2010), .Y(DP_OP_424J2_126_3477_n1973) );
  NOR2X1_HVT U2969 ( .A1(DP_OP_423J2_125_3477_n2316), .A2(n1499), .Y(
        DP_OP_425J2_127_3477_n2608) );
  NOR2X0_HVT U2970 ( .A1(DP_OP_425J2_127_3477_n2002), .A2(
        DP_OP_425J2_127_3477_n2010), .Y(DP_OP_425J2_127_3477_n1970) );
  OR2X1_HVT U2971 ( .A1(DP_OP_423J2_125_3477_n2005), .A2(
        DP_OP_423J2_125_3477_n2098), .Y(DP_OP_424J2_126_3477_n2061) );
  NOR2X1_HVT U2972 ( .A1(DP_OP_425J2_127_3477_n2048), .A2(
        DP_OP_424J2_126_3477_n2057), .Y(DP_OP_425J2_127_3477_n2040) );
  OR2X1_HVT U2973 ( .A1(DP_OP_422J2_124_3477_n2750), .A2(
        DP_OP_424J2_126_3477_n2409), .Y(DP_OP_424J2_126_3477_n2390) );
  NOR2X1_HVT U2974 ( .A1(DP_OP_424J2_126_3477_n2845), .A2(
        DP_OP_424J2_126_3477_n2231), .Y(DP_OP_425J2_127_3477_n2205) );
  NOR2X0_HVT U2975 ( .A1(DP_OP_422J2_124_3477_n2882), .A2(
        DP_OP_424J2_126_3477_n2758), .Y(DP_OP_425J2_127_3477_n2718) );
  OR2X1_HVT U2976 ( .A1(DP_OP_422J2_124_3477_n2753), .A2(
        DP_OP_422J2_124_3477_n2406), .Y(DP_OP_424J2_126_3477_n2369) );
  NOR2X0_HVT U2977 ( .A1(DP_OP_423J2_125_3477_n3056), .A2(
        DP_OP_425J2_127_3477_n2098), .Y(DP_OP_425J2_127_3477_n2058) );
  NOR2X0_HVT U2978 ( .A1(DP_OP_424J2_126_3477_n2002), .A2(n1507), .Y(
        DP_OP_425J2_127_3477_n2982) );
  NOR2X1_HVT U2979 ( .A1(DP_OP_425J2_127_3477_n2577), .A2(n671), .Y(
        DP_OP_425J2_127_3477_n2553) );
  NOR2X1_HVT U2980 ( .A1(DP_OP_425J2_127_3477_n2580), .A2(
        DP_OP_424J2_126_3477_n2585), .Y(DP_OP_425J2_127_3477_n2572) );
  OR2X1_HVT U2981 ( .A1(DP_OP_424J2_126_3477_n3058), .A2(
        DP_OP_425J2_127_3477_n2010), .Y(DP_OP_425J2_127_3477_n1972) );
  OR2X1_HVT U2982 ( .A1(DP_OP_422J2_124_3477_n2183), .A2(
        DP_OP_424J2_126_3477_n2758), .Y(DP_OP_424J2_126_3477_n2723) );
  OR2X1_HVT U2983 ( .A1(DP_OP_424J2_126_3477_n3019), .A2(
        DP_OP_423J2_125_3477_n3022), .Y(DP_OP_424J2_126_3477_n2987) );
  NOR2X1_HVT U2984 ( .A1(DP_OP_425J2_127_3477_n2977), .A2(
        DP_OP_424J2_126_3477_n2057), .Y(DP_OP_424J2_126_3477_n2045) );
  NOR2X1_HVT U2985 ( .A1(DP_OP_425J2_127_3477_n3063), .A2(
        DP_OP_423J2_125_3477_n3066), .Y(DP_OP_425J2_127_3477_n3047) );
  NOR2X1_HVT U2986 ( .A1(DP_OP_423J2_125_3477_n2317), .A2(n1499), .Y(
        DP_OP_425J2_127_3477_n2609) );
  OR2X1_HVT U2987 ( .A1(DP_OP_425J2_127_3477_n3056), .A2(
        DP_OP_424J2_126_3477_n3066), .Y(DP_OP_425J2_127_3477_n3040) );
  NOR2X1_HVT U2988 ( .A1(DP_OP_423J2_125_3477_n3062), .A2(n621), .Y(
        DP_OP_425J2_127_3477_n2088) );
  NOR2X1_HVT U2989 ( .A1(DP_OP_425J2_127_3477_n2448), .A2(n1499), .Y(
        DP_OP_424J2_126_3477_n2608) );
  NOR2X1_HVT U2990 ( .A1(DP_OP_422J2_124_3477_n2669), .A2(n1487), .Y(
        DP_OP_425J2_127_3477_n2521) );
  NOR2X1_HVT U2991 ( .A1(DP_OP_424J2_126_3477_n3020), .A2(
        DP_OP_425J2_127_3477_n2057), .Y(DP_OP_425J2_127_3477_n2044) );
  NOR2X1_HVT U2992 ( .A1(DP_OP_425J2_127_3477_n2048), .A2(
        DP_OP_422J2_124_3477_n3023), .Y(DP_OP_424J2_126_3477_n2992) );
  NOR2X1_HVT U2993 ( .A1(DP_OP_423J2_125_3477_n2005), .A2(n621), .Y(
        DP_OP_424J2_126_3477_n2085) );
  NOR2X1_HVT U2994 ( .A1(DP_OP_424J2_126_3477_n2622), .A2(n1498), .Y(
        DP_OP_424J2_126_3477_n2606) );
  NOR2X1_HVT U2995 ( .A1(DP_OP_424J2_126_3477_n2006), .A2(
        DP_OP_424J2_126_3477_n3023), .Y(DP_OP_425J2_127_3477_n2994) );
  NOR2X1_HVT U2996 ( .A1(DP_OP_425J2_127_3477_n2577), .A2(
        DP_OP_422J2_124_3477_n2585), .Y(DP_OP_425J2_127_3477_n2569) );
  NOR2X1_HVT U2997 ( .A1(DP_OP_424J2_126_3477_n2315), .A2(
        DP_OP_422J2_124_3477_n2715), .Y(DP_OP_425J2_127_3477_n2687) );
  NOR2X1_HVT U2998 ( .A1(DP_OP_425J2_127_3477_n2049), .A2(
        DP_OP_424J2_126_3477_n2057), .Y(DP_OP_425J2_127_3477_n2041) );
  NOR2X1_HVT U2999 ( .A1(DP_OP_425J2_127_3477_n2973), .A2(
        DP_OP_425J2_127_3477_n2057), .Y(DP_OP_424J2_126_3477_n2041) );
  NOR2X1_HVT U3000 ( .A1(DP_OP_425J2_127_3477_n3060), .A2(
        DP_OP_425J2_127_3477_n3066), .Y(DP_OP_425J2_127_3477_n3044) );
  NOR2X1_HVT U3001 ( .A1(DP_OP_424J2_126_3477_n2051), .A2(
        DP_OP_425J2_127_3477_n2057), .Y(DP_OP_424J2_126_3477_n2043) );
  NOR2X1_HVT U3002 ( .A1(DP_OP_425J2_127_3477_n2622), .A2(n1498), .Y(
        DP_OP_425J2_127_3477_n2606) );
  NOR2X1_HVT U3003 ( .A1(DP_OP_423J2_125_3477_n3059), .A2(n621), .Y(
        DP_OP_425J2_127_3477_n2085) );
  NOR2X1_HVT U3004 ( .A1(DP_OP_423J2_125_3477_n2665), .A2(
        DP_OP_424J2_126_3477_n2585), .Y(DP_OP_424J2_126_3477_n2569) );
  NOR2X1_HVT U3005 ( .A1(DP_OP_425J2_127_3477_n2401), .A2(
        DP_OP_422J2_124_3477_n2409), .Y(DP_OP_425J2_127_3477_n2393) );
  NOR2X1_HVT U3006 ( .A1(DP_OP_425J2_127_3477_n3019), .A2(
        DP_OP_422J2_124_3477_n3023), .Y(DP_OP_425J2_127_3477_n2995) );
  OR2X1_HVT U3007 ( .A1(DP_OP_425J2_127_3477_n3020), .A2(n1507), .Y(
        DP_OP_425J2_127_3477_n2988) );
  OR2X1_HVT U3008 ( .A1(DP_OP_423J2_125_3477_n3062), .A2(
        DP_OP_423J2_125_3477_n2098), .Y(DP_OP_425J2_127_3477_n2064) );
  OR2X1_HVT U3009 ( .A1(DP_OP_425J2_127_3477_n2404), .A2(
        DP_OP_422J2_124_3477_n2406), .Y(DP_OP_425J2_127_3477_n2372) );
  OR2X1_HVT U3010 ( .A1(DP_OP_423J2_125_3477_n2932), .A2(
        DP_OP_425J2_127_3477_n2230), .Y(DP_OP_425J2_127_3477_n2196) );
  NOR2X1_HVT U3011 ( .A1(DP_OP_424J2_126_3477_n3019), .A2(
        DP_OP_425J2_127_3477_n3023), .Y(DP_OP_424J2_126_3477_n2995) );
  NOR2X1_HVT U3012 ( .A1(DP_OP_424J2_126_3477_n2532), .A2(n1486), .Y(
        DP_OP_424J2_126_3477_n2516) );
  NOR2X1_HVT U3013 ( .A1(DP_OP_423J2_125_3477_n2708), .A2(n1499), .Y(
        DP_OP_424J2_126_3477_n2604) );
  OR2X1_HVT U3014 ( .A1(DP_OP_423J2_125_3477_n2008), .A2(
        DP_OP_425J2_127_3477_n2098), .Y(DP_OP_424J2_126_3477_n2064) );
  NOR2X1_HVT U3015 ( .A1(DP_OP_422J2_124_3477_n2664), .A2(n1486), .Y(
        DP_OP_425J2_127_3477_n2516) );
  NOR2X1_HVT U3016 ( .A1(DP_OP_423J2_125_3477_n2665), .A2(n671), .Y(
        DP_OP_424J2_126_3477_n2553) );
  OR2X1_HVT U3017 ( .A1(DP_OP_422J2_124_3477_n2756), .A2(n1426), .Y(
        DP_OP_424J2_126_3477_n2372) );
  NOR2X0_HVT U3018 ( .A1(DP_OP_422J2_124_3477_n3057), .A2(n621), .Y(
        DP_OP_424J2_126_3477_n2083) );
  NOR2X1_HVT U3019 ( .A1(DP_OP_422J2_124_3477_n2093), .A2(
        DP_OP_422J2_124_3477_n2847), .Y(DP_OP_424J2_126_3477_n2817) );
  NOR2X1_HVT U3020 ( .A1(DP_OP_424J2_126_3477_n2003), .A2(
        DP_OP_422J2_124_3477_n3023), .Y(DP_OP_425J2_127_3477_n2991) );
  NOR2X1_HVT U3021 ( .A1(DP_OP_425J2_127_3477_n2710), .A2(n1497), .Y(
        DP_OP_425J2_127_3477_n2686) );
  NOR2X1_HVT U3022 ( .A1(DP_OP_422J2_124_3477_n2091), .A2(
        DP_OP_422J2_124_3477_n2231), .Y(DP_OP_425J2_127_3477_n2199) );
  NOR2X1_HVT U3023 ( .A1(DP_OP_424J2_126_3477_n3063), .A2(
        DP_OP_424J2_126_3477_n3066), .Y(DP_OP_424J2_126_3477_n3047) );
  NOR2X1_HVT U3024 ( .A1(DP_OP_425J2_127_3477_n2449), .A2(n1498), .Y(
        DP_OP_424J2_126_3477_n2609) );
  NOR2X1_HVT U3025 ( .A1(DP_OP_422J2_124_3477_n2405), .A2(n1486), .Y(
        DP_OP_424J2_126_3477_n2521) );
  NOR2X1_HVT U3026 ( .A1(DP_OP_424J2_126_3477_n3059), .A2(
        DP_OP_423J2_125_3477_n3066), .Y(DP_OP_424J2_126_3477_n3043) );
  NOR2X1_HVT U3027 ( .A1(DP_OP_425J2_127_3477_n2972), .A2(
        DP_OP_424J2_126_3477_n2057), .Y(DP_OP_424J2_126_3477_n2040) );
  NOR2X1_HVT U3028 ( .A1(DP_OP_423J2_125_3477_n2097), .A2(n621), .Y(
        DP_OP_423J2_125_3477_n2089) );
  NOR2X1_HVT U3029 ( .A1(DP_OP_425J2_127_3477_n2976), .A2(
        DP_OP_424J2_126_3477_n2057), .Y(DP_OP_424J2_126_3477_n2044) );
  NOR2X1_HVT U3030 ( .A1(DP_OP_425J2_127_3477_n2801), .A2(n1500), .Y(
        DP_OP_423J2_125_3477_n2133) );
  NOR2X1_HVT U3031 ( .A1(DP_OP_425J2_127_3477_n2050), .A2(
        DP_OP_424J2_126_3477_n3023), .Y(DP_OP_424J2_126_3477_n2994) );
  NOR2X0_HVT U3032 ( .A1(DP_OP_423J2_125_3477_n2750), .A2(n1433), .Y(
        DP_OP_425J2_127_3477_n2366) );
  NOR2X1_HVT U3033 ( .A1(DP_OP_424J2_126_3477_n2619), .A2(n1499), .Y(
        DP_OP_424J2_126_3477_n2603) );
  OR2X1_HVT U3034 ( .A1(DP_OP_424J2_126_3477_n2268), .A2(
        DP_OP_424J2_126_3477_n2758), .Y(DP_OP_425J2_127_3477_n2720) );
  NOR2X1_HVT U3035 ( .A1(DP_OP_424J2_126_3477_n2576), .A2(n671), .Y(
        DP_OP_424J2_126_3477_n2552) );
  OR2X1_HVT U3036 ( .A1(DP_OP_424J2_126_3477_n2486), .A2(n1487), .Y(
        DP_OP_425J2_127_3477_n2514) );
  NOR2X1_HVT U3037 ( .A1(DP_OP_424J2_126_3477_n2580), .A2(
        DP_OP_424J2_126_3477_n2585), .Y(DP_OP_424J2_126_3477_n2572) );
  NOR2X1_HVT U3038 ( .A1(DP_OP_423J2_125_3477_n2315), .A2(n1498), .Y(
        DP_OP_425J2_127_3477_n2607) );
  NOR2X1_HVT U3039 ( .A1(DP_OP_425J2_127_3477_n2841), .A2(
        DP_OP_422J2_124_3477_n2847), .Y(DP_OP_425J2_127_3477_n2817) );
  NOR2X1_HVT U3040 ( .A1(DP_OP_422J2_124_3477_n2093), .A2(
        DP_OP_425J2_127_3477_n2231), .Y(DP_OP_425J2_127_3477_n2201) );
  NOR2X1_HVT U3041 ( .A1(DP_OP_424J2_126_3477_n2005), .A2(
        DP_OP_424J2_126_3477_n3023), .Y(DP_OP_425J2_127_3477_n2993) );
  OR2X1_HVT U3042 ( .A1(DP_OP_425J2_127_3477_n2578), .A2(
        DP_OP_422J2_124_3477_n2585), .Y(n1775) );
  OR2X1_HVT U3043 ( .A1(DP_OP_424J2_126_3477_n2222), .A2(
        DP_OP_423J2_125_3477_n2804), .Y(DP_OP_425J2_127_3477_n2778) );
  NOR2X1_HVT U3044 ( .A1(DP_OP_424J2_126_3477_n2669), .A2(
        DP_OP_425J2_127_3477_n2409), .Y(DP_OP_425J2_127_3477_n2397) );
  NOR2X1_HVT U3045 ( .A1(DP_OP_423J2_125_3477_n3063), .A2(n621), .Y(
        DP_OP_425J2_127_3477_n2089) );
  OR2X1_HVT U3046 ( .A1(DP_OP_423J2_125_3477_n2310), .A2(n1498), .Y(
        DP_OP_425J2_127_3477_n2602) );
  OR2X1_HVT U3047 ( .A1(DP_OP_424J2_126_3477_n2403), .A2(n1433), .Y(
        DP_OP_424J2_126_3477_n2371) );
  NOR2X1_HVT U3048 ( .A1(DP_OP_424J2_126_3477_n2136), .A2(n1500), .Y(
        DP_OP_424J2_126_3477_n2128) );
  OR2X1_HVT U3049 ( .A1(DP_OP_424J2_126_3477_n3059), .A2(
        DP_OP_425J2_127_3477_n2010), .Y(DP_OP_425J2_127_3477_n1973) );
  OR2X1_HVT U3050 ( .A1(DP_OP_423J2_125_3477_n2401), .A2(n1433), .Y(
        DP_OP_423J2_125_3477_n2369) );
  NOR2X0_HVT U3051 ( .A1(DP_OP_424J2_126_3477_n2090), .A2(
        DP_OP_423J2_125_3477_n2010), .Y(DP_OP_423J2_125_3477_n1970) );
  OR2X1_HVT U3052 ( .A1(DP_OP_423J2_125_3477_n2400), .A2(n1433), .Y(
        DP_OP_423J2_125_3477_n2368) );
  OR2X1_HVT U3053 ( .A1(DP_OP_423J2_125_3477_n2618), .A2(n1499), .Y(
        DP_OP_423J2_125_3477_n2602) );
  NOR2X1_HVT U3054 ( .A1(DP_OP_425J2_127_3477_n2796), .A2(n1501), .Y(
        DP_OP_423J2_125_3477_n2128) );
  NOR2X1_HVT U3055 ( .A1(DP_OP_422J2_124_3477_n2405), .A2(
        DP_OP_422J2_124_3477_n2409), .Y(DP_OP_422J2_124_3477_n2397) );
  XOR3X1_HVT U3056 ( .A1(n1546), .A2(n1547), .A3(n1548), .Y(
        DP_OP_422J2_124_3477_n1715) );
  NOR2X1_HVT U3057 ( .A1(DP_OP_423J2_125_3477_n3019), .A2(
        DP_OP_422J2_124_3477_n3023), .Y(DP_OP_423J2_125_3477_n2995) );
  NOR2X1_HVT U3058 ( .A1(DP_OP_423J2_125_3477_n3060), .A2(
        DP_OP_425J2_127_3477_n3066), .Y(DP_OP_423J2_125_3477_n3044) );
  NOR2X1_HVT U3059 ( .A1(DP_OP_422J2_124_3477_n3063), .A2(
        DP_OP_424J2_126_3477_n3066), .Y(DP_OP_422J2_124_3477_n3047) );
  NOR2X1_HVT U3060 ( .A1(DP_OP_422J2_124_3477_n2625), .A2(n1498), .Y(
        DP_OP_422J2_124_3477_n2609) );
  NOR2X1_HVT U3061 ( .A1(DP_OP_422J2_124_3477_n2444), .A2(n671), .Y(
        DP_OP_423J2_125_3477_n2552) );
  NOR2X1_HVT U3062 ( .A1(DP_OP_422J2_124_3477_n2622), .A2(n1499), .Y(
        DP_OP_422J2_124_3477_n2606) );
  NOR2X0_HVT U3063 ( .A1(DP_OP_423J2_125_3477_n2401), .A2(
        DP_OP_423J2_125_3477_n2409), .Y(DP_OP_423J2_125_3477_n2393) );
  OR2X1_HVT U3064 ( .A1(DP_OP_425J2_127_3477_n2840), .A2(
        DP_OP_423J2_125_3477_n2098), .Y(DP_OP_423J2_125_3477_n2060) );
  NOR2X1_HVT U3065 ( .A1(DP_OP_422J2_124_3477_n2049), .A2(n1475), .Y(
        DP_OP_422J2_124_3477_n2041) );
  NOR2X0_HVT U3066 ( .A1(DP_OP_423J2_125_3477_n3014), .A2(n1506), .Y(
        DP_OP_423J2_125_3477_n2982) );
  NOR2X0_HVT U3067 ( .A1(DP_OP_423J2_125_3477_n2090), .A2(
        DP_OP_423J2_125_3477_n2098), .Y(DP_OP_423J2_125_3477_n2058) );
  OR2X1_HVT U3068 ( .A1(DP_OP_423J2_125_3477_n2799), .A2(
        DP_OP_425J2_127_3477_n2230), .Y(DP_OP_422J2_124_3477_n2195) );
  NOR2X1_HVT U3069 ( .A1(DP_OP_422J2_124_3477_n2577), .A2(n670), .Y(
        DP_OP_422J2_124_3477_n2553) );
  OR2X1_HVT U3070 ( .A1(DP_OP_422J2_124_3477_n2756), .A2(
        DP_OP_422J2_124_3477_n2758), .Y(DP_OP_422J2_124_3477_n2724) );
  OR2X1_HVT U3071 ( .A1(DP_OP_425J2_127_3477_n2310), .A2(
        DP_OP_422J2_124_3477_n2847), .Y(DP_OP_423J2_125_3477_n2814) );
  OR2X1_HVT U3072 ( .A1(DP_OP_423J2_125_3477_n3019), .A2(
        DP_OP_423J2_125_3477_n3022), .Y(DP_OP_423J2_125_3477_n2987) );
  OR2X1_HVT U3073 ( .A1(DP_OP_422J2_124_3477_n3019), .A2(
        DP_OP_423J2_125_3477_n3022), .Y(DP_OP_422J2_124_3477_n2987) );
  NOR2X1_HVT U3074 ( .A1(DP_OP_423J2_125_3477_n2843), .A2(
        DP_OP_425J2_127_3477_n2847), .Y(DP_OP_423J2_125_3477_n2819) );
  OR2X1_HVT U3075 ( .A1(DP_OP_423J2_125_3477_n3056), .A2(
        DP_OP_423J2_125_3477_n3066), .Y(DP_OP_423J2_125_3477_n3040) );
  OR2X1_HVT U3076 ( .A1(DP_OP_424J2_126_3477_n2403), .A2(
        DP_OP_422J2_124_3477_n2758), .Y(DP_OP_422J2_124_3477_n2723) );
  NOR2X0_HVT U3077 ( .A1(DP_OP_425J2_127_3477_n2311), .A2(
        DP_OP_422J2_124_3477_n2847), .Y(DP_OP_423J2_125_3477_n2815) );
  OR2X1_HVT U3078 ( .A1(DP_OP_423J2_125_3477_n2399), .A2(
        DP_OP_422J2_124_3477_n2406), .Y(DP_OP_423J2_125_3477_n2367) );
  NOR2X1_HVT U3079 ( .A1(DP_OP_423J2_125_3477_n2841), .A2(
        DP_OP_422J2_124_3477_n2847), .Y(DP_OP_423J2_125_3477_n2817) );
  NOR2X1_HVT U3080 ( .A1(DP_OP_422J2_124_3477_n3060), .A2(
        DP_OP_423J2_125_3477_n3066), .Y(DP_OP_422J2_124_3477_n3044) );
  NOR2X1_HVT U3081 ( .A1(DP_OP_423J2_125_3477_n2620), .A2(n1499), .Y(
        DP_OP_423J2_125_3477_n2604) );
  NOR2X1_HVT U3082 ( .A1(DP_OP_422J2_124_3477_n2620), .A2(n1498), .Y(
        DP_OP_422J2_124_3477_n2604) );
  NOR2X1_HVT U3083 ( .A1(DP_OP_424J2_126_3477_n2845), .A2(n621), .Y(
        DP_OP_422J2_124_3477_n2089) );
  NOR2X1_HVT U3084 ( .A1(DP_OP_422J2_124_3477_n2404), .A2(
        DP_OP_425J2_127_3477_n2409), .Y(DP_OP_422J2_124_3477_n2396) );
  OR2X1_HVT U3085 ( .A1(DP_OP_423J2_125_3477_n2404), .A2(n1433), .Y(
        DP_OP_423J2_125_3477_n2372) );
  NOR2X1_HVT U3086 ( .A1(DP_OP_423J2_125_3477_n2795), .A2(
        DP_OP_423J2_125_3477_n2804), .Y(DP_OP_423J2_125_3477_n2779) );
  OR2X1_HVT U3087 ( .A1(DP_OP_422J2_124_3477_n2486), .A2(n1487), .Y(
        DP_OP_423J2_125_3477_n2514) );
  OR2X1_HVT U3088 ( .A1(DP_OP_422J2_124_3477_n2574), .A2(n1491), .Y(
        DP_OP_423J2_125_3477_n2470) );
  NOR2X1_HVT U3089 ( .A1(DP_OP_423J2_125_3477_n2619), .A2(n1498), .Y(
        DP_OP_423J2_125_3477_n2603) );
  NOR2X1_HVT U3090 ( .A1(DP_OP_423J2_125_3477_n2800), .A2(
        DP_OP_425J2_127_3477_n2231), .Y(DP_OP_422J2_124_3477_n2204) );
  NOR2X1_HVT U3091 ( .A1(DP_OP_422J2_124_3477_n2669), .A2(n279), .Y(
        DP_OP_422J2_124_3477_n2653) );
  NOR2X1_HVT U3092 ( .A1(DP_OP_423J2_125_3477_n2447), .A2(n1498), .Y(
        DP_OP_422J2_124_3477_n2607) );
  OR2X1_HVT U3093 ( .A1(DP_OP_424J2_126_3477_n2712), .A2(
        DP_OP_423J2_125_3477_n2230), .Y(DP_OP_422J2_124_3477_n2196) );
  OR2X1_HVT U3094 ( .A1(DP_OP_423J2_125_3477_n2094), .A2(
        DP_OP_423J2_125_3477_n2098), .Y(DP_OP_423J2_125_3477_n2062) );
  NOR2X1_HVT U3095 ( .A1(DP_OP_422J2_124_3477_n2537), .A2(n1486), .Y(
        DP_OP_422J2_124_3477_n2521) );
  OR2X1_HVT U3096 ( .A1(DP_OP_424J2_126_3477_n2932), .A2(
        DP_OP_423J2_125_3477_n3022), .Y(DP_OP_423J2_125_3477_n2988) );
  NOR2X1_HVT U3097 ( .A1(DP_OP_423J2_125_3477_n2886), .A2(
        DP_OP_425J2_127_3477_n2891), .Y(DP_OP_423J2_125_3477_n2862) );
  NOR2X1_HVT U3098 ( .A1(DP_OP_425J2_127_3477_n3021), .A2(
        DP_OP_423J2_125_3477_n2013), .Y(DP_OP_424J2_126_3477_n2001) );
  NOR2X0_HVT U3099 ( .A1(DP_OP_422J2_124_3477_n2620), .A2(n789), .Y(
        DP_OP_423J2_125_3477_n2420) );
  NOR2X1_HVT U3100 ( .A1(DP_OP_425J2_127_3477_n2268), .A2(
        DP_OP_425J2_127_3477_n2891), .Y(DP_OP_423J2_125_3477_n2860) );
  NOR2X1_HVT U3101 ( .A1(DP_OP_424J2_126_3477_n3060), .A2(
        DP_OP_423J2_125_3477_n2013), .Y(DP_OP_425J2_127_3477_n1998) );
  NOR2X0_HVT U3102 ( .A1(DP_OP_422J2_124_3477_n2621), .A2(n789), .Y(
        DP_OP_423J2_125_3477_n2421) );
  OR2X1_HVT U3103 ( .A1(DP_OP_423J2_125_3477_n2623), .A2(
        DP_OP_422J2_124_3477_n2626), .Y(DP_OP_423J2_125_3477_n2591) );
  AND2X1_HVT U3104 ( .A1(conv_weight_box[28]), .A2(src_window[149]), .Y(
        DP_OP_423J2_125_3477_n2816) );
  NOR2X1_HVT U3105 ( .A1(DP_OP_424J2_126_3477_n3058), .A2(
        DP_OP_422J2_124_3477_n2013), .Y(DP_OP_425J2_127_3477_n1996) );
  NOR2X1_HVT U3106 ( .A1(DP_OP_424J2_126_3477_n3059), .A2(n1431), .Y(
        DP_OP_425J2_127_3477_n1997) );
  NOR2X1_HVT U3107 ( .A1(DP_OP_423J2_125_3477_n2182), .A2(
        DP_OP_423J2_125_3477_n2892), .Y(DP_OP_422J2_124_3477_n2870) );
  OR2X1_HVT U3108 ( .A1(DP_OP_424J2_126_3477_n2794), .A2(
        DP_OP_424J2_126_3477_n2891), .Y(DP_OP_423J2_125_3477_n2858) );
  NOR2X1_HVT U3109 ( .A1(DP_OP_422J2_124_3477_n2625), .A2(n789), .Y(
        DP_OP_423J2_125_3477_n2425) );
  NOR2X1_HVT U3110 ( .A1(DP_OP_423J2_125_3477_n2887), .A2(
        DP_OP_423J2_125_3477_n2891), .Y(DP_OP_423J2_125_3477_n2863) );
  INVX1_HVT U3111 ( .A(conv_weight_box[18]), .Y(n1501) );
  NOR2X1_HVT U3112 ( .A1(DP_OP_422J2_124_3477_n2665), .A2(
        DP_OP_424J2_126_3477_n2671), .Y(DP_OP_422J2_124_3477_n2641) );
  INVX1_HVT U3113 ( .A(conv_weight_box[7]), .Y(n1507) );
  NOR2X1_HVT U3114 ( .A1(DP_OP_422J2_124_3477_n2888), .A2(
        DP_OP_423J2_125_3477_n2892), .Y(DP_OP_422J2_124_3477_n2872) );
  NOR2X0_HVT U3115 ( .A1(DP_OP_422J2_124_3477_n2310), .A2(
        DP_OP_422J2_124_3477_n2626), .Y(DP_OP_424J2_126_3477_n2586) );
  NOR2X1_HVT U3116 ( .A1(DP_OP_422J2_124_3477_n2137), .A2(
        DP_OP_424J2_126_3477_n2891), .Y(DP_OP_423J2_125_3477_n2861) );
  INVX1_HVT U3117 ( .A(conv_weight_box[18]), .Y(n1500) );
  OR2X1_HVT U3118 ( .A1(DP_OP_424J2_126_3477_n2623), .A2(n1331), .Y(
        DP_OP_424J2_126_3477_n2591) );
  INVX1_HVT U3119 ( .A(conv_weight_box[40]), .Y(DP_OP_423J2_125_3477_n2758) );
  NOR2X1_HVT U3120 ( .A1(DP_OP_422J2_124_3477_n2889), .A2(
        DP_OP_423J2_125_3477_n2892), .Y(DP_OP_422J2_124_3477_n2873) );
  NOR2X1_HVT U3121 ( .A1(DP_OP_424J2_126_3477_n2928), .A2(n1432), .Y(
        DP_OP_424J2_126_3477_n2904) );
  NOR2X1_HVT U3122 ( .A1(DP_OP_425J2_127_3477_n2138), .A2(
        DP_OP_425J2_127_3477_n2935), .Y(DP_OP_424J2_126_3477_n2906) );
  NOR2X1_HVT U3123 ( .A1(DP_OP_423J2_125_3477_n3019), .A2(n1432), .Y(
        DP_OP_424J2_126_3477_n2907) );
  NOR2X1_HVT U3124 ( .A1(DP_OP_424J2_126_3477_n2004), .A2(n1431), .Y(
        DP_OP_424J2_126_3477_n1996) );
  NOR2X1_HVT U3125 ( .A1(DP_OP_425J2_127_3477_n2272), .A2(
        DP_OP_425J2_127_3477_n2891), .Y(DP_OP_423J2_125_3477_n2864) );
  INVX1_HVT U3126 ( .A(conv_weight_box[7]), .Y(n1506) );
  NOR2X1_HVT U3127 ( .A1(DP_OP_424J2_126_3477_n2006), .A2(
        DP_OP_422J2_124_3477_n2013), .Y(DP_OP_424J2_126_3477_n1998) );
  OR2X1_HVT U3128 ( .A1(DP_OP_423J2_125_3477_n2447), .A2(
        DP_OP_422J2_124_3477_n2626), .Y(DP_OP_422J2_124_3477_n2591) );
  NOR2X1_HVT U3129 ( .A1(DP_OP_422J2_124_3477_n2885), .A2(
        DP_OP_423J2_125_3477_n2892), .Y(DP_OP_422J2_124_3477_n2869) );
  NOR2X1_HVT U3130 ( .A1(DP_OP_423J2_125_3477_n2404), .A2(n1400), .Y(
        DP_OP_422J2_124_3477_n2644) );
  NOR2X0_HVT U3131 ( .A1(DP_OP_425J2_127_3477_n2534), .A2(
        DP_OP_425J2_127_3477_n2671), .Y(DP_OP_422J2_124_3477_n2642) );
  INVX1_HVT U3132 ( .A(conv_weight_box[52]), .Y(DP_OP_422J2_124_3477_n2406) );
  NOR2X0_HVT U3133 ( .A1(DP_OP_422J2_124_3477_n2883), .A2(
        DP_OP_423J2_125_3477_n2892), .Y(DP_OP_422J2_124_3477_n2867) );
  INVX0_HVT U3134 ( .A(n1648), .Y(n1652) );
  INVX0_HVT U3135 ( .A(n1647), .Y(n1650) );
  NOR2X1_HVT U3136 ( .A1(DP_OP_424J2_126_3477_n3063), .A2(
        DP_OP_423J2_125_3477_n2013), .Y(DP_OP_425J2_127_3477_n2001) );
  INVX1_HVT U3137 ( .A(DP_OP_424J2_126_3477_n2791), .Y(n1513) );
  NOR2X1_HVT U3138 ( .A1(DP_OP_422J2_124_3477_n2313), .A2(n597), .Y(
        DP_OP_423J2_125_3477_n2701) );
  NOR2X1_HVT U3139 ( .A1(DP_OP_423J2_125_3477_n2624), .A2(
        DP_OP_423J2_125_3477_n2629), .Y(DP_OP_423J2_125_3477_n2616) );
  NOR2X1_HVT U3140 ( .A1(DP_OP_423J2_125_3477_n2316), .A2(
        DP_OP_423J2_125_3477_n2321), .Y(DP_OP_423J2_125_3477_n2308) );
  NOR2X1_HVT U3141 ( .A1(DP_OP_423J2_125_3477_n2621), .A2(
        DP_OP_423J2_125_3477_n2629), .Y(DP_OP_423J2_125_3477_n2613) );
  NOR2X1_HVT U3142 ( .A1(DP_OP_422J2_124_3477_n2621), .A2(
        DP_OP_422J2_124_3477_n2629), .Y(DP_OP_422J2_124_3477_n2613) );
  NOR2X1_HVT U3143 ( .A1(DP_OP_422J2_124_3477_n2751), .A2(n1333), .Y(
        DP_OP_424J2_126_3477_n2383) );
  NOR2X1_HVT U3144 ( .A1(DP_OP_424J2_126_3477_n2669), .A2(n1346), .Y(
        DP_OP_425J2_127_3477_n2389) );
  INVX2_HVT U3145 ( .A(conv_weight_box[15]), .Y(n1439) );
  INVX2_HVT U3146 ( .A(conv_weight_box[45]), .Y(n1440) );
  NOR2X1_HVT U3147 ( .A1(DP_OP_425J2_127_3477_n2622), .A2(
        DP_OP_423J2_125_3477_n2321), .Y(DP_OP_423J2_125_3477_n2306) );
  NOR2X1_HVT U3148 ( .A1(DP_OP_423J2_125_3477_n2620), .A2(
        DP_OP_423J2_125_3477_n2629), .Y(DP_OP_423J2_125_3477_n2612) );
  INVX0_HVT U3149 ( .A(DP_OP_422J2_124_3477_n2952), .Y(n1542) );
  NOR2X1_HVT U3150 ( .A1(DP_OP_423J2_125_3477_n2801), .A2(n597), .Y(
        DP_OP_424J2_126_3477_n2705) );
  NOR2X1_HVT U3151 ( .A1(DP_OP_425J2_127_3477_n2621), .A2(
        DP_OP_423J2_125_3477_n2321), .Y(DP_OP_423J2_125_3477_n2305) );
  INVX1_HVT U3152 ( .A(n1425), .Y(n1508) );
  NOR2X1_HVT U3153 ( .A1(DP_OP_425J2_127_3477_n2620), .A2(
        DP_OP_423J2_125_3477_n2321), .Y(DP_OP_423J2_125_3477_n2304) );
  NOR2X1_HVT U3154 ( .A1(DP_OP_424J2_126_3477_n2405), .A2(n1346), .Y(
        DP_OP_424J2_126_3477_n2389) );
  NOR2X1_HVT U3155 ( .A1(DP_OP_424J2_126_3477_n2712), .A2(n597), .Y(
        DP_OP_424J2_126_3477_n2704) );
  NOR2X1_HVT U3156 ( .A1(DP_OP_423J2_125_3477_n2448), .A2(
        DP_OP_422J2_124_3477_n2629), .Y(DP_OP_422J2_124_3477_n2616) );
  NOR2X1_HVT U3157 ( .A1(DP_OP_422J2_124_3477_n2754), .A2(
        DP_OP_424J2_126_3477_n2408), .Y(DP_OP_424J2_126_3477_n2386) );
  NOR2X1_HVT U3158 ( .A1(DP_OP_423J2_125_3477_n2625), .A2(
        DP_OP_423J2_125_3477_n2629), .Y(DP_OP_423J2_125_3477_n2617) );
  NOR2X1_HVT U3159 ( .A1(DP_OP_422J2_124_3477_n2797), .A2(n1444), .Y(
        DP_OP_422J2_124_3477_n2773) );
  NOR2X1_HVT U3160 ( .A1(DP_OP_423J2_125_3477_n2447), .A2(
        DP_OP_422J2_124_3477_n2629), .Y(DP_OP_422J2_124_3477_n2615) );
  AND2X1_HVT U3161 ( .A1(conv_weight_box[47]), .A2(src_window[208]), .Y(
        DP_OP_423J2_125_3477_n2353) );
  NOR2X1_HVT U3162 ( .A1(DP_OP_422J2_124_3477_n2225), .A2(n597), .Y(
        DP_OP_424J2_126_3477_n2701) );
  NOR2X1_HVT U3163 ( .A1(DP_OP_423J2_125_3477_n2317), .A2(
        DP_OP_423J2_125_3477_n2321), .Y(DP_OP_423J2_125_3477_n2309) );
  NOR2X1_HVT U3164 ( .A1(DP_OP_425J2_127_3477_n2799), .A2(
        DP_OP_423J2_125_3477_n2803), .Y(DP_OP_425J2_127_3477_n2775) );
  NOR2X1_HVT U3165 ( .A1(DP_OP_422J2_124_3477_n2625), .A2(
        DP_OP_422J2_124_3477_n2629), .Y(DP_OP_422J2_124_3477_n2617) );
  NOR2X1_HVT U3166 ( .A1(DP_OP_422J2_124_3477_n2620), .A2(
        DP_OP_422J2_124_3477_n2629), .Y(DP_OP_422J2_124_3477_n2612) );
  OR2X1_HVT U3167 ( .A1(DP_OP_424J2_126_3477_n2794), .A2(
        DP_OP_422J2_124_3477_n2803), .Y(DP_OP_424J2_126_3477_n2770) );
  NOR2X0_HVT U3168 ( .A1(DP_OP_423J2_125_3477_n2751), .A2(n1333), .Y(
        DP_OP_425J2_127_3477_n2383) );
  NOR2X1_HVT U3169 ( .A1(DP_OP_423J2_125_3477_n2315), .A2(
        DP_OP_423J2_125_3477_n2321), .Y(DP_OP_423J2_125_3477_n2307) );
  INVX1_HVT U3170 ( .A(conv_weight_box[9]), .Y(DP_OP_422J2_124_3477_n2056) );
  MUX21X1_HVT U3171 ( .A1(conv2_sram_rdata_weight[88]), .A2(
        conv1_sram_rdata_weight[88]), .S0(n1485), .Y(conv_weight_box[60]) );
  INVX1_HVT U3172 ( .A(conv_weight_box[9]), .Y(DP_OP_425J2_127_3477_n2056) );
  OR2X1_HVT U3173 ( .A1(DP_OP_422J2_124_3477_n2926), .A2(
        DP_OP_422J2_124_3477_n2803), .Y(DP_OP_425J2_127_3477_n2770) );
  MUX21X1_HVT U3174 ( .A1(conv2_sram_rdata_weight[11]), .A2(
        conv1_sram_rdata_weight[11]), .S0(n241), .Y(conv_weight_box[7]) );
  NOR2X1_HVT U3175 ( .A1(DP_OP_423J2_125_3477_n2623), .A2(
        DP_OP_423J2_125_3477_n2629), .Y(DP_OP_423J2_125_3477_n2615) );
  NOR2X1_HVT U3176 ( .A1(DP_OP_423J2_125_3477_n2754), .A2(n1333), .Y(
        DP_OP_425J2_127_3477_n2386) );
  NOR2X1_HVT U3177 ( .A1(DP_OP_425J2_127_3477_n2796), .A2(
        DP_OP_423J2_125_3477_n2803), .Y(DP_OP_425J2_127_3477_n2772) );
  NOR2X1_HVT U3178 ( .A1(DP_OP_423J2_125_3477_n2135), .A2(
        DP_OP_422J2_124_3477_n2803), .Y(DP_OP_425J2_127_3477_n2771) );
  MUX21X1_HVT U3179 ( .A1(conv2_sram_rdata_weight[21]), .A2(
        conv1_sram_rdata_weight[21]), .S0(n241), .Y(conv_weight_box[13]) );
  INVX0_HVT U3180 ( .A(n1646), .Y(n1649) );
  NOR2X1_HVT U3181 ( .A1(DP_OP_423J2_125_3477_n2800), .A2(
        DP_OP_423J2_125_3477_n2803), .Y(DP_OP_423J2_125_3477_n2776) );
  OR2X1_HVT U3182 ( .A1(DP_OP_422J2_124_3477_n2051), .A2(
        DP_OP_425J2_127_3477_n2186), .Y(DP_OP_425J2_127_3477_n2151) );
  INVX1_HVT U3183 ( .A(conv_weight_box[41]), .Y(DP_OP_422J2_124_3477_n2321) );
  INVX1_HVT U3184 ( .A(conv_weight_box[29]), .Y(DP_OP_425J2_127_3477_n2846) );
  INVX1_HVT U3185 ( .A(conv_weight_box[25]), .Y(DP_OP_422J2_124_3477_n2186) );
  INVX1_HVT U3186 ( .A(conv_weight_box[53]), .Y(DP_OP_423J2_125_3477_n2629) );
  INVX1_HVT U3187 ( .A(conv_weight_box[29]), .Y(DP_OP_424J2_126_3477_n2846) );
  INVX1_HVT U3188 ( .A(conv_weight_box[53]), .Y(DP_OP_422J2_124_3477_n2629) );
  MUX21X1_HVT U3189 ( .A1(conv2_sram_rdata_weight[63]), .A2(
        conv1_sram_rdata_weight[63]), .S0(n92), .Y(conv_weight_box[44]) );
  MUX21X1_HVT U3190 ( .A1(conv2_sram_rdata_weight[57]), .A2(
        conv1_sram_rdata_weight[57]), .S0(n345), .Y(conv_weight_box[39]) );
  INVX1_HVT U3191 ( .A(srstn), .Y(n1445) );
  INVX0_HVT U3192 ( .A(n2081), .Y(n2105) );
  INVX0_HVT U3193 ( .A(n2069), .Y(n2106) );
  INVX0_HVT U3194 ( .A(n2022), .Y(n2047) );
  INVX0_HVT U3195 ( .A(n2030), .Y(n2046) );
  AO22X1_HVT U3196 ( .A1(conv2_sum_b[10]), .A2(n1849), .A3(conv2_sum_b[11]), 
        .A4(n1973), .Y(n2033) );
  XOR3X2_HVT U3197 ( .A1(DP_OP_423J2_125_3477_n824), .A2(
        DP_OP_423J2_125_3477_n653), .A3(DP_OP_423J2_125_3477_n651), .Y(
        DP_OP_423J2_125_3477_n649) );
  NAND2X0_HVT U3198 ( .A1(DP_OP_423J2_125_3477_n824), .A2(
        DP_OP_423J2_125_3477_n651), .Y(n1446) );
  NAND2X0_HVT U3199 ( .A1(DP_OP_423J2_125_3477_n653), .A2(
        DP_OP_423J2_125_3477_n651), .Y(n1447) );
  NAND2X0_HVT U3200 ( .A1(DP_OP_423J2_125_3477_n653), .A2(
        DP_OP_423J2_125_3477_n824), .Y(n1448) );
  NAND3X0_HVT U3201 ( .A1(n1448), .A2(n1447), .A3(n1446), .Y(
        DP_OP_423J2_125_3477_n648) );
  OR2X1_HVT U3202 ( .A1(DP_OP_422J2_124_3477_n3029), .A2(
        DP_OP_422J2_124_3477_n2502), .Y(DP_OP_422J2_124_3477_n1210) );
  NAND2X0_HVT U3203 ( .A1(DP_OP_424J2_126_3477_n514), .A2(
        DP_OP_424J2_126_3477_n423), .Y(n1449) );
  XOR3X2_HVT U3204 ( .A1(DP_OP_425J2_127_3477_n831), .A2(
        DP_OP_425J2_127_3477_n1022), .A3(DP_OP_425J2_127_3477_n829), .Y(
        DP_OP_425J2_127_3477_n825) );
  NAND2X0_HVT U3205 ( .A1(DP_OP_425J2_127_3477_n831), .A2(
        DP_OP_425J2_127_3477_n829), .Y(n1450) );
  NAND2X0_HVT U3206 ( .A1(DP_OP_425J2_127_3477_n1022), .A2(
        DP_OP_425J2_127_3477_n829), .Y(n1451) );
  NAND2X0_HVT U3207 ( .A1(DP_OP_425J2_127_3477_n1022), .A2(
        DP_OP_425J2_127_3477_n831), .Y(n1452) );
  NAND2X0_HVT U3208 ( .A1(DP_OP_425J2_127_3477_n168), .A2(n1453), .Y(n1454) );
  NAND2X0_HVT U3209 ( .A1(n1454), .A2(n1455), .Y(n_conv2_sum_d[18]) );
  XOR3X2_HVT U3210 ( .A1(DP_OP_422J2_124_3477_n1120), .A2(
        DP_OP_422J2_124_3477_n1132), .A3(DP_OP_422J2_124_3477_n1134), .Y(
        DP_OP_422J2_124_3477_n901) );
  NAND2X0_HVT U3211 ( .A1(DP_OP_422J2_124_3477_n1120), .A2(
        DP_OP_422J2_124_3477_n1134), .Y(n1456) );
  NAND2X0_HVT U3212 ( .A1(DP_OP_422J2_124_3477_n1132), .A2(
        DP_OP_422J2_124_3477_n1134), .Y(n1457) );
  NAND2X0_HVT U3213 ( .A1(DP_OP_422J2_124_3477_n1132), .A2(
        DP_OP_422J2_124_3477_n1120), .Y(n1458) );
  NAND3X0_HVT U3214 ( .A1(n1458), .A2(n1457), .A3(n1456), .Y(
        DP_OP_422J2_124_3477_n900) );
  XOR3X2_HVT U3215 ( .A1(DP_OP_422J2_124_3477_n2649), .A2(
        DP_OP_422J2_124_3477_n2612), .A3(DP_OP_422J2_124_3477_n2605), .Y(
        DP_OP_422J2_124_3477_n1333) );
  NAND2X0_HVT U3216 ( .A1(DP_OP_422J2_124_3477_n2649), .A2(
        DP_OP_422J2_124_3477_n2605), .Y(n1459) );
  NAND2X0_HVT U3217 ( .A1(DP_OP_422J2_124_3477_n2612), .A2(
        DP_OP_422J2_124_3477_n2605), .Y(n1460) );
  NAND2X0_HVT U3218 ( .A1(DP_OP_422J2_124_3477_n2612), .A2(
        DP_OP_422J2_124_3477_n2649), .Y(n1461) );
  NAND3X0_HVT U3219 ( .A1(n1461), .A2(n1460), .A3(n1459), .Y(
        DP_OP_422J2_124_3477_n1332) );
  XOR3X2_HVT U3220 ( .A1(DP_OP_422J2_124_3477_n359), .A2(
        DP_OP_422J2_124_3477_n382), .A3(DP_OP_422J2_124_3477_n380), .Y(
        DP_OP_422J2_124_3477_n355) );
  NAND2X0_HVT U3221 ( .A1(DP_OP_422J2_124_3477_n359), .A2(
        DP_OP_422J2_124_3477_n380), .Y(n1462) );
  NAND2X0_HVT U3222 ( .A1(DP_OP_422J2_124_3477_n382), .A2(
        DP_OP_422J2_124_3477_n380), .Y(n1463) );
  NAND2X0_HVT U3223 ( .A1(DP_OP_422J2_124_3477_n382), .A2(
        DP_OP_422J2_124_3477_n359), .Y(n1464) );
  NAND3X0_HVT U3224 ( .A1(n1464), .A2(n1463), .A3(n1462), .Y(
        DP_OP_422J2_124_3477_n354) );
  XOR3X2_HVT U3225 ( .A1(DP_OP_423J2_125_3477_n650), .A2(
        DP_OP_423J2_125_3477_n517), .A3(DP_OP_423J2_125_3477_n515), .Y(
        DP_OP_423J2_125_3477_n513) );
  NAND2X0_HVT U3226 ( .A1(DP_OP_423J2_125_3477_n650), .A2(
        DP_OP_423J2_125_3477_n515), .Y(n1465) );
  NAND2X0_HVT U3227 ( .A1(DP_OP_423J2_125_3477_n517), .A2(
        DP_OP_423J2_125_3477_n515), .Y(n1466) );
  NAND2X0_HVT U3228 ( .A1(DP_OP_423J2_125_3477_n517), .A2(
        DP_OP_423J2_125_3477_n650), .Y(n1467) );
  XOR3X2_HVT U3229 ( .A1(DP_OP_423J2_125_3477_n1433), .A2(
        DP_OP_423J2_125_3477_n1592), .A3(DP_OP_423J2_125_3477_n1590), .Y(
        DP_OP_423J2_125_3477_n1415) );
  NAND2X0_HVT U3230 ( .A1(DP_OP_423J2_125_3477_n1433), .A2(
        DP_OP_423J2_125_3477_n1592), .Y(n1468) );
  NAND2X0_HVT U3231 ( .A1(DP_OP_423J2_125_3477_n1433), .A2(
        DP_OP_423J2_125_3477_n1590), .Y(n1469) );
  NAND2X0_HVT U3232 ( .A1(DP_OP_423J2_125_3477_n1590), .A2(
        DP_OP_423J2_125_3477_n1592), .Y(n1470) );
  XOR2X1_HVT U3233 ( .A1(DP_OP_423J2_125_3477_n1235), .A2(
        DP_OP_423J2_125_3477_n1412), .Y(n1471) );
  XOR2X1_HVT U3234 ( .A1(n1471), .A2(DP_OP_423J2_125_3477_n1414), .Y(
        DP_OP_423J2_125_3477_n1223) );
  NAND2X0_HVT U3235 ( .A1(DP_OP_423J2_125_3477_n1235), .A2(
        DP_OP_423J2_125_3477_n1412), .Y(n1472) );
  NAND2X0_HVT U3236 ( .A1(DP_OP_423J2_125_3477_n1235), .A2(
        DP_OP_423J2_125_3477_n1414), .Y(n1473) );
  NAND2X0_HVT U3237 ( .A1(DP_OP_423J2_125_3477_n1412), .A2(
        DP_OP_423J2_125_3477_n1414), .Y(n1474) );
  NAND3X0_HVT U3238 ( .A1(n1473), .A2(n1472), .A3(n1474), .Y(
        DP_OP_423J2_125_3477_n1222) );
  INVX1_HVT U3239 ( .A(conv_weight_box[8]), .Y(n1475) );
  MUX21X1_HVT U3240 ( .A1(conv2_sram_rdata_weight[12]), .A2(
        conv1_sram_rdata_weight[12]), .S0(n240), .Y(conv_weight_box[8]) );
  MUX21X1_HVT U3241 ( .A1(conv2_sram_rdata_weight[28]), .A2(
        conv1_sram_rdata_weight[28]), .S0(n241), .Y(conv_weight_box[18]) );
  INVX1_HVT U3242 ( .A(conv_weight_box[32]), .Y(DP_OP_423J2_125_3477_n2230) );
  NOR2X0_HVT U3243 ( .A1(DP_OP_424J2_126_3477_n2795), .A2(
        DP_OP_425J2_127_3477_n2891), .Y(DP_OP_423J2_125_3477_n2859) );
  OR2X1_HVT U3244 ( .A1(DP_OP_425J2_127_3477_n2970), .A2(
        DP_OP_424J2_126_3477_n2057), .Y(DP_OP_424J2_126_3477_n2038) );
  OR2X1_HVT U3245 ( .A1(DP_OP_422J2_124_3477_n512), .A2(
        DP_OP_422J2_124_3477_n419), .Y(n1544) );
  NAND2X0_HVT U3246 ( .A1(DP_OP_423J2_125_3477_n1020), .A2(
        DP_OP_423J2_125_3477_n825), .Y(n1478) );
  NAND2X0_HVT U3247 ( .A1(DP_OP_423J2_125_3477_n827), .A2(
        DP_OP_423J2_125_3477_n825), .Y(n1479) );
  NAND2X0_HVT U3248 ( .A1(DP_OP_423J2_125_3477_n827), .A2(
        DP_OP_423J2_125_3477_n1020), .Y(n1480) );
  NAND3X0_HVT U3249 ( .A1(n1480), .A2(n1479), .A3(n1478), .Y(
        DP_OP_423J2_125_3477_n822) );
  OR2X1_HVT U3250 ( .A1(DP_OP_423J2_125_3477_n2052), .A2(n1506), .Y(
        DP_OP_422J2_124_3477_n2988) );
  NOR2X4_HVT U3251 ( .A1(DP_OP_422J2_124_3477_n2663), .A2(n1400), .Y(
        DP_OP_422J2_124_3477_n2639) );
  INVX2_HVT U3252 ( .A(srstn), .Y(n1494) );
  INVX1_HVT U3253 ( .A(srstn), .Y(n1495) );
  INVX2_HVT U3254 ( .A(srstn), .Y(n1493) );
  INVX2_HVT U3255 ( .A(srstn), .Y(n1492) );
  INVX1_HVT U3256 ( .A(conv_weight_box[34]), .Y(DP_OP_422J2_124_3477_n2803) );
  MUX21X1_HVT U3257 ( .A1(conv2_sram_rdata_weight[59]), .A2(
        conv1_sram_rdata_weight[59]), .S0(n1418), .Y(conv_weight_box[40]) );
  MUX21X1_HVT U3258 ( .A1(conv2_sram_rdata_weight[30]), .A2(
        conv1_sram_rdata_weight[30]), .S0(n1418), .Y(conv_weight_box[20]) );
  INVX1_HVT U3259 ( .A(conv_weight_box[67]), .Y(n1486) );
  INVX1_HVT U3260 ( .A(conv_weight_box[67]), .Y(n1487) );
  INVX1_HVT U3261 ( .A(conv_weight_box[67]), .Y(DP_OP_424J2_126_3477_n2540) );
  INVX1_HVT U3262 ( .A(conv_weight_box[58]), .Y(n1489) );
  INVX1_HVT U3263 ( .A(conv_weight_box[63]), .Y(DP_OP_423J2_125_3477_n2496) );
  INVX1_HVT U3264 ( .A(conv_weight_box[42]), .Y(DP_OP_423J2_125_3477_n2320) );
  NOR2X0_HVT U3265 ( .A1(DP_OP_422J2_124_3477_n2224), .A2(
        DP_OP_422J2_124_3477_n2717), .Y(DP_OP_424J2_126_3477_n2700) );
  OR2X1_HVT U3266 ( .A1(DP_OP_424J2_126_3477_n2311), .A2(
        DP_OP_425J2_127_3477_n2230), .Y(DP_OP_423J2_125_3477_n2191) );
  NOR2X0_HVT U3267 ( .A1(DP_OP_423J2_125_3477_n2222), .A2(
        DP_OP_423J2_125_3477_n2230), .Y(DP_OP_423J2_125_3477_n2190) );
  NOR2X0_HVT U3268 ( .A1(DP_OP_422J2_124_3477_n2222), .A2(
        DP_OP_422J2_124_3477_n2230), .Y(DP_OP_422J2_124_3477_n2190) );
  OR2X1_HVT U3269 ( .A1(DP_OP_425J2_127_3477_n2708), .A2(
        DP_OP_425J2_127_3477_n2230), .Y(DP_OP_423J2_125_3477_n2192) );
  OR2X1_HVT U3270 ( .A1(DP_OP_422J2_124_3477_n2224), .A2(
        DP_OP_423J2_125_3477_n2230), .Y(DP_OP_422J2_124_3477_n2192) );
  OR2X1_HVT U3271 ( .A1(DP_OP_425J2_127_3477_n2710), .A2(
        DP_OP_423J2_125_3477_n2230), .Y(DP_OP_423J2_125_3477_n2194) );
  OR2X1_HVT U3272 ( .A1(DP_OP_423J2_125_3477_n2228), .A2(
        DP_OP_422J2_124_3477_n2230), .Y(DP_OP_423J2_125_3477_n2196) );
  MUX21X1_HVT U3273 ( .A1(conv2_sum_d[22]), .A2(conv2_sum_c[22]), .S0(n1496), 
        .Y(tmp_big2[22]) );
  MUX21X1_HVT U3274 ( .A1(conv2_sum_d[8]), .A2(conv2_sum_c[8]), .S0(n1994), 
        .Y(tmp_big2[8]) );
  OR2X1_HVT U3275 ( .A1(DP_OP_425J2_127_3477_n2574), .A2(n1497), .Y(
        DP_OP_422J2_124_3477_n2682) );
  NOR2X0_HVT U3276 ( .A1(DP_OP_422J2_124_3477_n2223), .A2(n1440), .Y(
        DP_OP_424J2_126_3477_n2683) );
  OR2X1_HVT U3277 ( .A1(DP_OP_422J2_124_3477_n2750), .A2(n1346), .Y(
        DP_OP_424J2_126_3477_n2382) );
  OR2X1_HVT U3278 ( .A1(DP_OP_423J2_125_3477_n2750), .A2(
        DP_OP_424J2_126_3477_n2408), .Y(DP_OP_425J2_127_3477_n2382) );
  OR2X1_HVT U3279 ( .A1(DP_OP_425J2_127_3477_n2574), .A2(
        DP_OP_422J2_124_3477_n2585), .Y(DP_OP_425J2_127_3477_n2566) );
  INVX1_HVT U3280 ( .A(conv_weight_box[60]), .Y(DP_OP_423J2_125_3477_n2585) );
  INVX1_HVT U3281 ( .A(conv_weight_box[54]), .Y(n1498) );
  INVX1_HVT U3282 ( .A(conv_weight_box[54]), .Y(n1499) );
  OR2X1_HVT U3283 ( .A1(DP_OP_425J2_127_3477_n2882), .A2(n1442), .Y(
        DP_OP_424J2_126_3477_n2126) );
  OR2X1_HVT U3284 ( .A1(DP_OP_423J2_125_3477_n3014), .A2(n1501), .Y(
        DP_OP_425J2_127_3477_n2126) );
  NOR2X0_HVT U3285 ( .A1(DP_OP_425J2_127_3477_n2883), .A2(n1442), .Y(
        DP_OP_424J2_126_3477_n2127) );
  OR2X1_HVT U3286 ( .A1(DP_OP_424J2_126_3477_n2222), .A2(n1501), .Y(
        DP_OP_423J2_125_3477_n2126) );
  INVX1_HVT U3287 ( .A(conv_weight_box[13]), .Y(DP_OP_423J2_125_3477_n2100) );
  AND2X1_HVT U3288 ( .A1(n1972), .A2(n1970), .Y(n1505) );
  INVX1_HVT U3289 ( .A(conv_weight_box[7]), .Y(DP_OP_423J2_125_3477_n3022) );
  NAND2X0_HVT U3290 ( .A1(DP_OP_422J2_124_3477_n523), .A2(
        DP_OP_422J2_124_3477_n656), .Y(n1509) );
  NAND2X0_HVT U3291 ( .A1(DP_OP_422J2_124_3477_n654), .A2(
        DP_OP_422J2_124_3477_n523), .Y(n1510) );
  NAND2X0_HVT U3292 ( .A1(DP_OP_422J2_124_3477_n654), .A2(
        DP_OP_422J2_124_3477_n656), .Y(n1511) );
  FADDX1_HVT U3293 ( .A(n1512), .B(DP_OP_424J2_126_3477_n2821), .CI(
        DP_OP_424J2_126_3477_n2791), .CO(DP_OP_424J2_126_3477_n1788) );
  XOR3X2_HVT U3294 ( .A1(DP_OP_424J2_126_3477_n2821), .A2(n1514), .A3(n1513), 
        .Y(DP_OP_424J2_126_3477_n1789) );
  NAND2X0_HVT U3295 ( .A1(conv_weight_box[47]), .A2(src_window[215]), .Y(
        DP_OP_423J2_125_3477_n2346) );
  AND2X1_HVT U3296 ( .A1(conv_weight_box[47]), .A2(src_window[213]), .Y(
        DP_OP_423J2_125_3477_n2348) );
  AND2X1_HVT U3297 ( .A1(conv_weight_box[47]), .A2(src_window[210]), .Y(
        DP_OP_423J2_125_3477_n2351) );
  AND2X1_HVT U3298 ( .A1(conv_weight_box[47]), .A2(src_window[211]), .Y(
        DP_OP_423J2_125_3477_n2350) );
  AND2X1_HVT U3299 ( .A1(conv_weight_box[47]), .A2(src_window[212]), .Y(
        DP_OP_423J2_125_3477_n2349) );
  AND2X1_HVT U3300 ( .A1(conv_weight_box[47]), .A2(src_window[214]), .Y(
        DP_OP_423J2_125_3477_n2347) );
  AND2X1_HVT U3301 ( .A1(conv_weight_box[47]), .A2(src_window[209]), .Y(
        DP_OP_423J2_125_3477_n2352) );
  NAND2X0_HVT U3302 ( .A1(conv_weight_box[17]), .A2(src_window[111]), .Y(
        DP_OP_423J2_125_3477_n2902) );
  AO21X1_HVT U3303 ( .A1(n1832), .A2(DP_OP_425J2_127_3477_n100), .A3(
        DP_OP_425J2_127_3477_n101), .Y(n1520) );
  XOR2X2_HVT U3304 ( .A1(n1664), .A2(DP_OP_423J2_125_3477_n7), .Y(
        n_conv2_sum_b[30]) );
  XOR2X2_HVT U3305 ( .A1(n1667), .A2(DP_OP_423J2_125_3477_n8), .Y(
        n_conv2_sum_b[29]) );
  XOR2X2_HVT U3306 ( .A1(n1662), .A2(DP_OP_423J2_125_3477_n16), .Y(
        n_conv2_sum_b[21]) );
  XOR2X2_HVT U3307 ( .A1(n1663), .A2(DP_OP_423J2_125_3477_n18), .Y(
        n_conv2_sum_b[19]) );
  XOR2X2_HVT U3308 ( .A1(n1661), .A2(DP_OP_423J2_125_3477_n20), .Y(
        n_conv2_sum_b[17]) );
  XOR2X2_HVT U3309 ( .A1(n1659), .A2(DP_OP_423J2_125_3477_n21), .Y(
        n_conv2_sum_b[16]) );
  XOR2X2_HVT U3310 ( .A1(n1608), .A2(DP_OP_423J2_125_3477_n22), .Y(
        n_conv2_sum_b[15]) );
  XOR2X2_HVT U3311 ( .A1(n1660), .A2(DP_OP_423J2_125_3477_n13), .Y(
        n_conv2_sum_b[24]) );
  AND2X1_HVT U3312 ( .A1(src_window[144]), .A2(conv_weight_box[28]), .Y(
        DP_OP_423J2_125_3477_n2821) );
  AO21X1_HVT U3313 ( .A1(n1517), .A2(DP_OP_422J2_124_3477_n151), .A3(
        DP_OP_422J2_124_3477_n152), .Y(n1521) );
  NAND2X0_HVT U3314 ( .A1(n1622), .A2(n1609), .Y(n1522) );
  OR2X4_HVT U3315 ( .A1(DP_OP_422J2_124_3477_n2267), .A2(n1426), .Y(
        DP_OP_425J2_127_3477_n2367) );
  OR2X2_HVT U3316 ( .A1(DP_OP_425J2_127_3477_n2401), .A2(
        DP_OP_422J2_124_3477_n2406), .Y(DP_OP_425J2_127_3477_n2369) );
  OR2X2_HVT U3317 ( .A1(DP_OP_425J2_127_3477_n2400), .A2(
        DP_OP_422J2_124_3477_n2406), .Y(DP_OP_425J2_127_3477_n2368) );
  OR2X2_HVT U3318 ( .A1(DP_OP_422J2_124_3477_n2401), .A2(n1426), .Y(
        DP_OP_422J2_124_3477_n2369) );
  INVX2_HVT U3319 ( .A(DP_OP_423J2_125_3477_n4), .Y(n1614) );
  AND2X1_HVT U3320 ( .A1(DP_OP_422J2_124_3477_n340), .A2(
        DP_OP_422J2_124_3477_n335), .Y(n1525) );
  XOR2X2_HVT U3321 ( .A1(n1526), .A2(n1527), .Y(n_conv2_sum_b[27]) );
  AO21X1_HVT U3322 ( .A1(DP_OP_423J2_125_3477_n4), .A2(
        DP_OP_423J2_125_3477_n80), .A3(DP_OP_423J2_125_3477_n81), .Y(n1526) );
  AND2X1_HVT U3323 ( .A1(DP_OP_423J2_125_3477_n274), .A2(
        DP_OP_423J2_125_3477_n78), .Y(n1527) );
  AND2X1_HVT U3324 ( .A1(DP_OP_423J2_125_3477_n340), .A2(
        DP_OP_423J2_125_3477_n335), .Y(n1528) );
  MUX21X1_HVT U3325 ( .A1(tmp_big2[19]), .A2(tmp_big1[19]), .S0(n1481), .Y(
        data_out[19]) );
  NAND2X0_HVT U3326 ( .A1(tmp_big2[13]), .A2(n2156), .Y(n1529) );
  OR2X2_HVT U3327 ( .A1(DP_OP_425J2_127_3477_n2534), .A2(
        DP_OP_422J2_124_3477_n2406), .Y(DP_OP_423J2_125_3477_n2370) );
  AND3X1_HVT U3328 ( .A1(n1601), .A2(n1600), .A3(n1599), .Y(n1530) );
  NOR2X0_HVT U3329 ( .A1(DP_OP_423J2_125_3477_n2842), .A2(n1438), .Y(
        DP_OP_423J2_125_3477_n2818) );
  INVX1_HVT U3330 ( .A(DP_OP_422J2_124_3477_n1728), .Y(
        DP_OP_422J2_124_3477_n1729) );
  INVX1_HVT U3331 ( .A(src_window[71]), .Y(DP_OP_422J2_124_3477_n2002) );
  INVX1_HVT U3332 ( .A(src_window[70]), .Y(DP_OP_422J2_124_3477_n2003) );
  INVX1_HVT U3333 ( .A(src_window[69]), .Y(DP_OP_422J2_124_3477_n2004) );
  INVX1_HVT U3334 ( .A(src_window[68]), .Y(DP_OP_422J2_124_3477_n2005) );
  INVX1_HVT U3335 ( .A(src_window[67]), .Y(DP_OP_422J2_124_3477_n2006) );
  INVX1_HVT U3336 ( .A(src_window[66]), .Y(DP_OP_422J2_124_3477_n2007) );
  INVX1_HVT U3337 ( .A(src_window[87]), .Y(DP_OP_422J2_124_3477_n2046) );
  INVX1_HVT U3338 ( .A(src_window[86]), .Y(DP_OP_422J2_124_3477_n2047) );
  INVX1_HVT U3339 ( .A(src_window[85]), .Y(DP_OP_422J2_124_3477_n2048) );
  INVX1_HVT U3340 ( .A(src_window[84]), .Y(DP_OP_422J2_124_3477_n2049) );
  INVX1_HVT U3341 ( .A(src_window[82]), .Y(DP_OP_422J2_124_3477_n2051) );
  INVX1_HVT U3342 ( .A(src_window[111]), .Y(DP_OP_422J2_124_3477_n2090) );
  INVX1_HVT U3343 ( .A(src_window[110]), .Y(DP_OP_422J2_124_3477_n2091) );
  INVX1_HVT U3344 ( .A(src_window[109]), .Y(DP_OP_422J2_124_3477_n2092) );
  INVX1_HVT U3345 ( .A(src_window[108]), .Y(DP_OP_422J2_124_3477_n2093) );
  INVX1_HVT U3346 ( .A(src_window[127]), .Y(DP_OP_422J2_124_3477_n2134) );
  INVX1_HVT U3347 ( .A(src_window[126]), .Y(DP_OP_422J2_124_3477_n2135) );
  INVX1_HVT U3348 ( .A(src_window[124]), .Y(DP_OP_422J2_124_3477_n2137) );
  INVX1_HVT U3349 ( .A(src_window[123]), .Y(DP_OP_422J2_124_3477_n2138) );
  INVX1_HVT U3350 ( .A(src_window[121]), .Y(DP_OP_422J2_124_3477_n2140) );
  INVX1_HVT U3351 ( .A(src_window[143]), .Y(DP_OP_422J2_124_3477_n2178) );
  INVX1_HVT U3352 ( .A(src_window[142]), .Y(DP_OP_422J2_124_3477_n2179) );
  INVX1_HVT U3353 ( .A(src_window[140]), .Y(DP_OP_422J2_124_3477_n2181) );
  INVX1_HVT U3354 ( .A(src_window[138]), .Y(DP_OP_422J2_124_3477_n2183) );
  INVX1_HVT U3355 ( .A(src_window[136]), .Y(DP_OP_422J2_124_3477_n2185) );
  INVX1_HVT U3356 ( .A(src_window[167]), .Y(DP_OP_422J2_124_3477_n2222) );
  INVX1_HVT U3357 ( .A(src_window[166]), .Y(DP_OP_422J2_124_3477_n2223) );
  INVX1_HVT U3358 ( .A(src_window[165]), .Y(DP_OP_422J2_124_3477_n2224) );
  INVX1_HVT U3359 ( .A(src_window[164]), .Y(DP_OP_422J2_124_3477_n2225) );
  INVX1_HVT U3360 ( .A(src_window[183]), .Y(DP_OP_422J2_124_3477_n2266) );
  INVX1_HVT U3361 ( .A(src_window[182]), .Y(DP_OP_422J2_124_3477_n2267) );
  INVX1_HVT U3362 ( .A(src_window[181]), .Y(DP_OP_422J2_124_3477_n2268) );
  INVX1_HVT U3363 ( .A(src_window[180]), .Y(DP_OP_422J2_124_3477_n2269) );
  INVX1_HVT U3364 ( .A(src_window[179]), .Y(DP_OP_422J2_124_3477_n2270) );
  INVX1_HVT U3365 ( .A(src_window[207]), .Y(DP_OP_422J2_124_3477_n2310) );
  INVX1_HVT U3366 ( .A(src_window[206]), .Y(DP_OP_422J2_124_3477_n2311) );
  INVX1_HVT U3367 ( .A(src_window[205]), .Y(DP_OP_422J2_124_3477_n2312) );
  INVX1_HVT U3368 ( .A(src_window[204]), .Y(DP_OP_422J2_124_3477_n2313) );
  INVX1_HVT U3369 ( .A(src_window[203]), .Y(DP_OP_422J2_124_3477_n2314) );
  INVX1_HVT U3370 ( .A(src_window[223]), .Y(DP_OP_422J2_124_3477_n2354) );
  INVX1_HVT U3371 ( .A(src_window[222]), .Y(DP_OP_422J2_124_3477_n2355) );
  INVX1_HVT U3372 ( .A(src_window[221]), .Y(DP_OP_422J2_124_3477_n2356) );
  INVX1_HVT U3373 ( .A(src_window[220]), .Y(DP_OP_422J2_124_3477_n2357) );
  INVX1_HVT U3374 ( .A(src_window[219]), .Y(DP_OP_422J2_124_3477_n2358) );
  INVX1_HVT U3375 ( .A(src_window[239]), .Y(DP_OP_422J2_124_3477_n2398) );
  INVX1_HVT U3376 ( .A(src_window[238]), .Y(DP_OP_422J2_124_3477_n2399) );
  INVX1_HVT U3377 ( .A(src_window[236]), .Y(DP_OP_422J2_124_3477_n2401) );
  INVX1_HVT U3378 ( .A(src_window[233]), .Y(DP_OP_422J2_124_3477_n2404) );
  INVX1_HVT U3379 ( .A(src_window[232]), .Y(DP_OP_422J2_124_3477_n2405) );
  INVX1_HVT U3380 ( .A(src_window[263]), .Y(DP_OP_422J2_124_3477_n2442) );
  INVX1_HVT U3381 ( .A(src_window[262]), .Y(DP_OP_422J2_124_3477_n2443) );
  INVX1_HVT U3382 ( .A(src_window[261]), .Y(DP_OP_422J2_124_3477_n2444) );
  INVX1_HVT U3383 ( .A(src_window[260]), .Y(DP_OP_422J2_124_3477_n2445) );
  INVX1_HVT U3384 ( .A(src_window[259]), .Y(DP_OP_422J2_124_3477_n2446) );
  INVX1_HVT U3385 ( .A(src_window[257]), .Y(DP_OP_422J2_124_3477_n2448) );
  INVX1_HVT U3386 ( .A(src_window[279]), .Y(DP_OP_422J2_124_3477_n2486) );
  INVX1_HVT U3387 ( .A(src_window[277]), .Y(DP_OP_422J2_124_3477_n2488) );
  INVX1_HVT U3388 ( .A(src_window[276]), .Y(DP_OP_422J2_124_3477_n2489) );
  INVX1_HVT U3389 ( .A(src_window[275]), .Y(DP_OP_422J2_124_3477_n2490) );
  INVX1_HVT U3390 ( .A(src_window[274]), .Y(DP_OP_422J2_124_3477_n2491) );
  INVX1_HVT U3391 ( .A(src_window[287]), .Y(DP_OP_422J2_124_3477_n2530) );
  INVX1_HVT U3392 ( .A(src_window[286]), .Y(DP_OP_422J2_124_3477_n2531) );
  INVX1_HVT U3393 ( .A(src_window[285]), .Y(DP_OP_422J2_124_3477_n2532) );
  INVX1_HVT U3394 ( .A(src_window[284]), .Y(DP_OP_422J2_124_3477_n2533) );
  INVX1_HVT U3395 ( .A(src_window[283]), .Y(DP_OP_422J2_124_3477_n2534) );
  INVX1_HVT U3396 ( .A(src_window[282]), .Y(DP_OP_422J2_124_3477_n2535) );
  INVX1_HVT U3397 ( .A(src_window[281]), .Y(DP_OP_422J2_124_3477_n2536) );
  INVX1_HVT U3398 ( .A(src_window[280]), .Y(DP_OP_422J2_124_3477_n2537) );
  INVX1_HVT U3399 ( .A(src_window[271]), .Y(DP_OP_422J2_124_3477_n2574) );
  INVX1_HVT U3400 ( .A(src_window[270]), .Y(DP_OP_422J2_124_3477_n2575) );
  INVX1_HVT U3401 ( .A(src_window[269]), .Y(DP_OP_422J2_124_3477_n2576) );
  INVX1_HVT U3402 ( .A(src_window[268]), .Y(DP_OP_422J2_124_3477_n2577) );
  INVX1_HVT U3403 ( .A(src_window[267]), .Y(DP_OP_422J2_124_3477_n2578) );
  INVX1_HVT U3404 ( .A(src_window[266]), .Y(DP_OP_422J2_124_3477_n2579) );
  INVX1_HVT U3405 ( .A(src_window[265]), .Y(DP_OP_422J2_124_3477_n2580) );
  INVX1_HVT U3406 ( .A(src_window[255]), .Y(DP_OP_422J2_124_3477_n2618) );
  INVX1_HVT U3407 ( .A(src_window[254]), .Y(DP_OP_422J2_124_3477_n2619) );
  INVX1_HVT U3408 ( .A(src_window[253]), .Y(DP_OP_422J2_124_3477_n2620) );
  INVX1_HVT U3409 ( .A(src_window[252]), .Y(DP_OP_422J2_124_3477_n2621) );
  INVX1_HVT U3410 ( .A(src_window[251]), .Y(DP_OP_422J2_124_3477_n2622) );
  INVX1_HVT U3411 ( .A(src_window[248]), .Y(DP_OP_422J2_124_3477_n2625) );
  INVX1_HVT U3412 ( .A(src_window[231]), .Y(DP_OP_422J2_124_3477_n2662) );
  INVX1_HVT U3413 ( .A(src_window[230]), .Y(DP_OP_422J2_124_3477_n2663) );
  INVX1_HVT U3414 ( .A(src_window[229]), .Y(DP_OP_422J2_124_3477_n2664) );
  INVX1_HVT U3415 ( .A(src_window[228]), .Y(DP_OP_422J2_124_3477_n2665) );
  INVX1_HVT U3416 ( .A(src_window[226]), .Y(DP_OP_422J2_124_3477_n2667) );
  INVX1_HVT U3417 ( .A(src_window[224]), .Y(DP_OP_422J2_124_3477_n2669) );
  INVX1_HVT U3418 ( .A(conv_weight_box[49]), .Y(DP_OP_422J2_124_3477_n2673) );
  INVX1_HVT U3419 ( .A(src_window[214]), .Y(DP_OP_422J2_124_3477_n2707) );
  INVX1_HVT U3420 ( .A(src_window[213]), .Y(DP_OP_422J2_124_3477_n2708) );
  INVX1_HVT U3421 ( .A(src_window[212]), .Y(DP_OP_422J2_124_3477_n2709) );
  INVX1_HVT U3422 ( .A(src_window[211]), .Y(DP_OP_422J2_124_3477_n2710) );
  INVX1_HVT U3423 ( .A(src_window[209]), .Y(DP_OP_422J2_124_3477_n2712) );
  INVX1_HVT U3424 ( .A(src_window[191]), .Y(DP_OP_422J2_124_3477_n2750) );
  INVX1_HVT U3425 ( .A(src_window[190]), .Y(DP_OP_422J2_124_3477_n2751) );
  INVX1_HVT U3426 ( .A(src_window[188]), .Y(DP_OP_422J2_124_3477_n2753) );
  INVX1_HVT U3427 ( .A(src_window[187]), .Y(DP_OP_422J2_124_3477_n2754) );
  INVX1_HVT U3428 ( .A(src_window[185]), .Y(DP_OP_422J2_124_3477_n2756) );
  INVX1_HVT U3429 ( .A(src_window[175]), .Y(DP_OP_422J2_124_3477_n2794) );
  INVX1_HVT U3430 ( .A(src_window[174]), .Y(DP_OP_422J2_124_3477_n2795) );
  INVX1_HVT U3431 ( .A(src_window[173]), .Y(DP_OP_422J2_124_3477_n2796) );
  INVX1_HVT U3432 ( .A(src_window[172]), .Y(DP_OP_422J2_124_3477_n2797) );
  INVX1_HVT U3433 ( .A(src_window[171]), .Y(DP_OP_422J2_124_3477_n2798) );
  INVX1_HVT U3434 ( .A(src_window[170]), .Y(DP_OP_422J2_124_3477_n2799) );
  INVX1_HVT U3435 ( .A(src_window[169]), .Y(DP_OP_422J2_124_3477_n2800) );
  INVX1_HVT U3436 ( .A(src_window[159]), .Y(DP_OP_422J2_124_3477_n2838) );
  INVX1_HVT U3437 ( .A(src_window[158]), .Y(DP_OP_422J2_124_3477_n2839) );
  INVX1_HVT U3438 ( .A(src_window[157]), .Y(DP_OP_422J2_124_3477_n2840) );
  INVX1_HVT U3439 ( .A(src_window[156]), .Y(DP_OP_422J2_124_3477_n2841) );
  INVX1_HVT U3440 ( .A(src_window[155]), .Y(DP_OP_422J2_124_3477_n2842) );
  INVX1_HVT U3441 ( .A(src_window[135]), .Y(DP_OP_422J2_124_3477_n2882) );
  INVX1_HVT U3442 ( .A(src_window[134]), .Y(DP_OP_422J2_124_3477_n2883) );
  INVX1_HVT U3443 ( .A(src_window[133]), .Y(DP_OP_422J2_124_3477_n2884) );
  INVX1_HVT U3444 ( .A(src_window[132]), .Y(DP_OP_422J2_124_3477_n2885) );
  INVX1_HVT U3445 ( .A(src_window[130]), .Y(DP_OP_422J2_124_3477_n2887) );
  INVX1_HVT U3446 ( .A(src_window[129]), .Y(DP_OP_422J2_124_3477_n2888) );
  INVX1_HVT U3447 ( .A(src_window[128]), .Y(DP_OP_422J2_124_3477_n2889) );
  INVX1_HVT U3448 ( .A(src_window[119]), .Y(DP_OP_422J2_124_3477_n2926) );
  INVX1_HVT U3449 ( .A(src_window[118]), .Y(DP_OP_422J2_124_3477_n2927) );
  INVX1_HVT U3450 ( .A(src_window[117]), .Y(DP_OP_422J2_124_3477_n2928) );
  INVX1_HVT U3451 ( .A(src_window[116]), .Y(DP_OP_422J2_124_3477_n2929) );
  INVX1_HVT U3452 ( .A(src_window[115]), .Y(DP_OP_422J2_124_3477_n2930) );
  INVX1_HVT U3453 ( .A(src_window[95]), .Y(DP_OP_422J2_124_3477_n2970) );
  INVX1_HVT U3454 ( .A(src_window[94]), .Y(DP_OP_422J2_124_3477_n2971) );
  INVX1_HVT U3455 ( .A(src_window[93]), .Y(DP_OP_422J2_124_3477_n2972) );
  INVX1_HVT U3456 ( .A(src_window[92]), .Y(DP_OP_422J2_124_3477_n2973) );
  INVX1_HVT U3457 ( .A(src_window[91]), .Y(DP_OP_422J2_124_3477_n2974) );
  INVX1_HVT U3458 ( .A(src_window[90]), .Y(DP_OP_422J2_124_3477_n2975) );
  INVX1_HVT U3459 ( .A(src_window[79]), .Y(DP_OP_422J2_124_3477_n3014) );
  INVX1_HVT U3460 ( .A(src_window[78]), .Y(DP_OP_422J2_124_3477_n3015) );
  INVX1_HVT U3461 ( .A(src_window[76]), .Y(DP_OP_422J2_124_3477_n3017) );
  INVX1_HVT U3462 ( .A(src_window[74]), .Y(DP_OP_422J2_124_3477_n3019) );
  INVX1_HVT U3463 ( .A(src_window[72]), .Y(DP_OP_422J2_124_3477_n3021) );
  INVX1_HVT U3464 ( .A(DP_OP_422J2_124_3477_n302), .Y(
        DP_OP_422J2_124_3477_n303) );
  INVX1_HVT U3465 ( .A(DP_OP_422J2_124_3477_n304), .Y(
        DP_OP_422J2_124_3477_n305) );
  INVX1_HVT U3466 ( .A(src_window[63]), .Y(DP_OP_422J2_124_3477_n3056) );
  INVX1_HVT U3467 ( .A(src_window[62]), .Y(DP_OP_422J2_124_3477_n3057) );
  INVX1_HVT U3468 ( .A(src_window[61]), .Y(DP_OP_422J2_124_3477_n3058) );
  INVX1_HVT U3469 ( .A(src_window[60]), .Y(DP_OP_422J2_124_3477_n3059) );
  INVX1_HVT U3470 ( .A(src_window[59]), .Y(DP_OP_422J2_124_3477_n3060) );
  INVX1_HVT U3471 ( .A(src_window[56]), .Y(DP_OP_422J2_124_3477_n3063) );
  INVX1_HVT U3472 ( .A(DP_OP_422J2_124_3477_n308), .Y(
        DP_OP_422J2_124_3477_n309) );
  INVX1_HVT U3473 ( .A(DP_OP_422J2_124_3477_n310), .Y(
        DP_OP_422J2_124_3477_n311) );
  INVX1_HVT U3474 ( .A(DP_OP_422J2_124_3477_n312), .Y(
        DP_OP_422J2_124_3477_n313) );
  INVX1_HVT U3475 ( .A(DP_OP_422J2_124_3477_n314), .Y(
        DP_OP_422J2_124_3477_n315) );
  INVX1_HVT U3476 ( .A(DP_OP_422J2_124_3477_n316), .Y(
        DP_OP_422J2_124_3477_n317) );
  INVX1_HVT U3477 ( .A(DP_OP_422J2_124_3477_n318), .Y(
        DP_OP_422J2_124_3477_n319) );
  INVX1_HVT U3478 ( .A(DP_OP_422J2_124_3477_n320), .Y(
        DP_OP_422J2_124_3477_n321) );
  INVX1_HVT U3479 ( .A(DP_OP_422J2_124_3477_n322), .Y(
        DP_OP_422J2_124_3477_n323) );
  INVX1_HVT U3480 ( .A(DP_OP_422J2_124_3477_n324), .Y(
        DP_OP_422J2_124_3477_n325) );
  INVX1_HVT U3481 ( .A(DP_OP_422J2_124_3477_n326), .Y(
        DP_OP_422J2_124_3477_n327) );
  INVX1_HVT U3482 ( .A(DP_OP_422J2_124_3477_n328), .Y(
        DP_OP_422J2_124_3477_n329) );
  INVX1_HVT U3483 ( .A(DP_OP_422J2_124_3477_n330), .Y(
        DP_OP_422J2_124_3477_n331) );
  INVX1_HVT U3484 ( .A(DP_OP_422J2_124_3477_n510), .Y(
        DP_OP_422J2_124_3477_n511) );
  INVX1_HVT U3485 ( .A(DP_OP_422J2_124_3477_n71), .Y(DP_OP_422J2_124_3477_n69)
         );
  INVX1_HVT U3486 ( .A(DP_OP_422J2_124_3477_n820), .Y(
        DP_OP_422J2_124_3477_n821) );
  INVX1_HVT U3487 ( .A(DP_OP_422J2_124_3477_n95), .Y(DP_OP_422J2_124_3477_n93)
         );
  NAND2X0_HVT U3488 ( .A1(DP_OP_422J2_124_3477_n649), .A2(
        DP_OP_422J2_124_3477_n822), .Y(DP_OP_422J2_124_3477_n240) );
  NAND2X0_HVT U3489 ( .A1(n1538), .A2(n1542), .Y(n1541) );
  AO22X1_HVT U3490 ( .A1(DP_OP_422J2_124_3477_n2952), .A2(n1540), .A3(
        DP_OP_422J2_124_3477_n2922), .A4(n1541), .Y(DP_OP_422J2_124_3477_n1682) );
  XOR3X2_HVT U3491 ( .A1(DP_OP_422J2_124_3477_n379), .A2(
        DP_OP_422J2_124_3477_n424), .A3(DP_OP_422J2_124_3477_n422), .Y(
        DP_OP_422J2_124_3477_n375) );
  OR2X1_HVT U3492 ( .A1(DP_OP_422J2_124_3477_n424), .A2(
        DP_OP_422J2_124_3477_n379), .Y(n1543) );
  AO22X1_HVT U3493 ( .A1(DP_OP_422J2_124_3477_n379), .A2(
        DP_OP_422J2_124_3477_n424), .A3(DP_OP_422J2_124_3477_n422), .A4(n1543), 
        .Y(DP_OP_422J2_124_3477_n374) );
  NAND2X0_HVT U3494 ( .A1(n1535), .A2(DP_OP_422J2_124_3477_n244), .Y(
        DP_OP_422J2_124_3477_n242) );
  NAND2X0_HVT U3495 ( .A1(conv_weight_box[35]), .A2(src_window[168]), .Y(n1548) );
  NAND2X0_HVT U3496 ( .A1(n1546), .A2(n1547), .Y(n1549) );
  NAND2X0_HVT U3497 ( .A1(n1549), .A2(n1548), .Y(n1550) );
  OR2X1_HVT U3498 ( .A1(n1547), .A2(n1546), .Y(n1551) );
  NAND2X0_HVT U3499 ( .A1(n1550), .A2(n1551), .Y(DP_OP_422J2_124_3477_n1714)
         );
  NAND2X0_HVT U3500 ( .A1(DP_OP_422J2_124_3477_n4), .A2(
        DP_OP_422J2_124_3477_n122), .Y(n1552) );
  NAND2X0_HVT U3501 ( .A1(DP_OP_422J2_124_3477_n4), .A2(
        DP_OP_422J2_124_3477_n91), .Y(n1555) );
  NAND2X0_HVT U3502 ( .A1(DP_OP_422J2_124_3477_n4), .A2(
        DP_OP_422J2_124_3477_n131), .Y(n1557) );
  NAND2X0_HVT U3503 ( .A1(DP_OP_422J2_124_3477_n4), .A2(
        DP_OP_422J2_124_3477_n100), .Y(n1559) );
  NAND2X0_HVT U3504 ( .A1(DP_OP_422J2_124_3477_n4), .A2(
        DP_OP_422J2_124_3477_n80), .Y(n1561) );
  AO21X1_HVT U3505 ( .A1(n1517), .A2(DP_OP_422J2_124_3477_n187), .A3(
        DP_OP_422J2_124_3477_n188), .Y(n1563) );
  AO21X1_HVT U3506 ( .A1(n1517), .A2(DP_OP_422J2_124_3477_n158), .A3(
        DP_OP_422J2_124_3477_n159), .Y(n1564) );
  AO21X1_HVT U3507 ( .A1(DP_OP_422J2_124_3477_n4), .A2(
        DP_OP_422J2_124_3477_n176), .A3(DP_OP_422J2_124_3477_n177), .Y(n1565)
         );
  AO21X1_HVT U3508 ( .A1(DP_OP_422J2_124_3477_n4), .A2(
        DP_OP_422J2_124_3477_n138), .A3(DP_OP_422J2_124_3477_n139), .Y(n1566)
         );
  AO21X1_HVT U3509 ( .A1(n1517), .A2(DP_OP_422J2_124_3477_n49), .A3(
        DP_OP_422J2_124_3477_n50), .Y(n1567) );
  AO21X1_HVT U3510 ( .A1(n1517), .A2(DP_OP_422J2_124_3477_n169), .A3(
        DP_OP_422J2_124_3477_n170), .Y(n1568) );
  AO21X1_HVT U3511 ( .A1(n1517), .A2(n1595), .A3(n1594), .Y(n1569) );
  NAND2X0_HVT U3512 ( .A1(conv_weight_box[29]), .A2(src_window[152]), .Y(
        DP_OP_422J2_124_3477_n2813) );
  NAND2X0_HVT U3513 ( .A1(conv_weight_box[32]), .A2(src_window[160]), .Y(
        DP_OP_422J2_124_3477_n2197) );
  AND2X1_HVT U3514 ( .A1(conv_weight_box[37]), .A2(src_window[182]), .Y(
        DP_OP_422J2_124_3477_n2251) );
  OR2X1_HVT U3515 ( .A1(DP_OP_422J2_124_3477_n2688), .A2(
        DP_OP_422J2_124_3477_n2695), .Y(n1571) );
  AO22X1_HVT U3516 ( .A1(DP_OP_422J2_124_3477_n2688), .A2(
        DP_OP_422J2_124_3477_n2695), .A3(DP_OP_422J2_124_3477_n1834), .A4(
        n1571), .Y(DP_OP_422J2_124_3477_n1660) );
  AND2X1_HVT U3517 ( .A1(n1572), .A2(n1530), .Y(DP_OP_422J2_124_3477_n214) );
  NAND2X0_HVT U3518 ( .A1(n1573), .A2(DP_OP_422J2_124_3477_n226), .Y(n1574) );
  NAND2X0_HVT U3519 ( .A1(n1575), .A2(DP_OP_422J2_124_3477_n226), .Y(n1576) );
  OA21X1_HVT U3520 ( .A1(n1577), .A2(DP_OP_422J2_124_3477_n248), .A3(
        DP_OP_422J2_124_3477_n249), .Y(DP_OP_422J2_124_3477_n245) );
  OR2X1_HVT U3521 ( .A1(DP_OP_422J2_124_3477_n1018), .A2(
        DP_OP_422J2_124_3477_n823), .Y(n1579) );
  NAND2X0_HVT U3522 ( .A1(n1578), .A2(n1579), .Y(n1535) );
  NAND2X0_HVT U3523 ( .A1(DP_OP_422J2_124_3477_n419), .A2(
        DP_OP_422J2_124_3477_n512), .Y(n1573) );
  NAND2X0_HVT U3524 ( .A1(DP_OP_422J2_124_3477_n4), .A2(
        DP_OP_422J2_124_3477_n107), .Y(n1581) );
  XOR3X2_HVT U3525 ( .A1(DP_OP_422J2_124_3477_n943), .A2(
        DP_OP_422J2_124_3477_n1108), .A3(DP_OP_422J2_124_3477_n1098), .Y(
        DP_OP_422J2_124_3477_n891) );
  OR2X1_HVT U3526 ( .A1(DP_OP_422J2_124_3477_n943), .A2(
        DP_OP_422J2_124_3477_n1108), .Y(n1582) );
  AO22X1_HVT U3527 ( .A1(DP_OP_422J2_124_3477_n1108), .A2(
        DP_OP_422J2_124_3477_n943), .A3(n1582), .A4(DP_OP_422J2_124_3477_n1098), .Y(DP_OP_422J2_124_3477_n890) );
  OR2X1_HVT U3528 ( .A1(DP_OP_422J2_124_3477_n302), .A2(n1584), .Y(n1583) );
  OR2X1_HVT U3529 ( .A1(DP_OP_422J2_124_3477_n304), .A2(
        DP_OP_422J2_124_3477_n303), .Y(n1585) );
  OR2X1_HVT U3530 ( .A1(DP_OP_422J2_124_3477_n308), .A2(n1383), .Y(n1586) );
  OR2X1_HVT U3531 ( .A1(DP_OP_422J2_124_3477_n312), .A2(
        DP_OP_422J2_124_3477_n311), .Y(n1587) );
  OR2X1_HVT U3532 ( .A1(DP_OP_422J2_124_3477_n318), .A2(
        DP_OP_422J2_124_3477_n317), .Y(n1588) );
  INVX1_HVT U3533 ( .A(n1536), .Y(DP_OP_422J2_124_3477_n236) );
  OR2X1_HVT U3534 ( .A1(DP_OP_422J2_124_3477_n1403), .A2(
        DP_OP_422J2_124_3477_n1401), .Y(n1590) );
  OR2X1_HVT U3535 ( .A1(DP_OP_422J2_124_3477_n1733), .A2(
        DP_OP_422J2_124_3477_n1731), .Y(n1591) );
  AND2X1_HVT U3536 ( .A1(n1536), .A2(n1537), .Y(n1593) );
  AND2X1_HVT U3537 ( .A1(DP_OP_422J2_124_3477_n49), .A2(n1585), .Y(n1595) );
  INVX1_HVT U3538 ( .A(conv_weight_box[29]), .Y(DP_OP_422J2_124_3477_n2846) );
  INVX1_HVT U3539 ( .A(conv_weight_box[32]), .Y(DP_OP_422J2_124_3477_n2230) );
  OR2X1_HVT U3540 ( .A1(DP_OP_422J2_124_3477_n2578), .A2(
        DP_OP_422J2_124_3477_n2585), .Y(n1538) );
  INVX1_HVT U3541 ( .A(DP_OP_422J2_124_3477_n2922), .Y(n1539) );
  OA21X1_HVT U3542 ( .A1(DP_OP_422J2_124_3477_n209), .A2(
        DP_OP_422J2_124_3477_n217), .A3(DP_OP_422J2_124_3477_n210), .Y(n1589)
         );
  OA21X1_HVT U3543 ( .A1(DP_OP_422J2_124_3477_n93), .A2(
        DP_OP_422J2_124_3477_n110), .A3(DP_OP_422J2_124_3477_n94), .Y(n1556)
         );
  NAND2X0_HVT U3544 ( .A1(DP_OP_422J2_124_3477_n177), .A2(
        DP_OP_422J2_124_3477_n142), .Y(n1553) );
  AND2X1_HVT U3545 ( .A1(n1553), .A2(DP_OP_422J2_124_3477_n145), .Y(
        DP_OP_422J2_124_3477_n141) );
  OA21X1_HVT U3546 ( .A1(DP_OP_422J2_124_3477_n82), .A2(
        DP_OP_422J2_124_3477_n110), .A3(DP_OP_422J2_124_3477_n85), .Y(n1562)
         );
  INVX1_HVT U3547 ( .A(conv_weight_box[11]), .Y(DP_OP_422J2_124_3477_n2980) );
  INVX1_HVT U3548 ( .A(DP_OP_422J2_124_3477_n233), .Y(
        DP_OP_422J2_124_3477_n232) );
  INVX1_HVT U3549 ( .A(conv_weight_box[36]), .Y(DP_OP_422J2_124_3477_n2277) );
  INVX1_HVT U3550 ( .A(conv_weight_box[42]), .Y(DP_OP_422J2_124_3477_n2320) );
  INVX1_HVT U3551 ( .A(conv_weight_box[21]), .Y(DP_OP_422J2_124_3477_n2893) );
  INVX1_HVT U3552 ( .A(conv_weight_box[62]), .Y(DP_OP_422J2_124_3477_n2497) );
  OR2X1_HVT U3553 ( .A1(DP_OP_422J2_124_3477_n822), .A2(
        DP_OP_422J2_124_3477_n649), .Y(n1537) );
  INVX1_HVT U3554 ( .A(conv_weight_box[38]), .Y(DP_OP_422J2_124_3477_n2275) );
  INVX1_HVT U3555 ( .A(conv_weight_box[66]), .Y(DP_OP_422J2_124_3477_n2541) );
  INVX1_HVT U3556 ( .A(conv_weight_box[51]), .Y(DP_OP_422J2_124_3477_n2409) );
  INVX1_HVT U3557 ( .A(conv_weight_box[19]), .Y(DP_OP_422J2_124_3477_n2144) );
  INVX1_HVT U3558 ( .A(conv_weight_box[24]), .Y(DP_OP_422J2_124_3477_n2189) );
  INVX1_HVT U3559 ( .A(conv_weight_box[13]), .Y(DP_OP_422J2_124_3477_n2100) );
  INVX1_HVT U3560 ( .A(conv_weight_box[60]), .Y(DP_OP_422J2_124_3477_n2585) );
  INVX1_HVT U3561 ( .A(conv_weight_box[31]), .Y(DP_OP_422J2_124_3477_n2231) );
  INVX1_HVT U3562 ( .A(DP_OP_422J2_124_3477_n338), .Y(
        DP_OP_422J2_124_3477_n339) );
  INVX1_HVT U3563 ( .A(conv_weight_box[6]), .Y(DP_OP_422J2_124_3477_n3023) );
  INVX1_HVT U3564 ( .A(conv_weight_box[10]), .Y(DP_OP_422J2_124_3477_n2055) );
  INVX1_HVT U3565 ( .A(conv_weight_box[3]), .Y(DP_OP_422J2_124_3477_n2011) );
  INVX1_HVT U3566 ( .A(conv_weight_box[40]), .Y(DP_OP_422J2_124_3477_n2758) );
  INVX1_HVT U3567 ( .A(conv_weight_box[55]), .Y(DP_OP_422J2_124_3477_n2627) );
  INVX1_HVT U3568 ( .A(conv_weight_box[61]), .Y(DP_OP_422J2_124_3477_n2582) );
  INVX1_HVT U3569 ( .A(conv_weight_box[48]), .Y(DP_OP_422J2_124_3477_n2362) );
  INVX1_HVT U3570 ( .A(conv_weight_box[46]), .Y(DP_OP_422J2_124_3477_n2714) );
  INVX1_HVT U3571 ( .A(conv_weight_box[44]), .Y(DP_OP_422J2_124_3477_n2318) );
  INVX1_HVT U3572 ( .A(DP_OP_422J2_124_3477_n197), .Y(
        DP_OP_422J2_124_3477_n286) );
  INVX2_HVT U3573 ( .A(conv_weight_box[28]), .Y(DP_OP_422J2_124_3477_n2847) );
  NAND3X0_HVT U3574 ( .A1(n1596), .A2(n1597), .A3(n1598), .Y(
        DP_OP_422J2_124_3477_n1044) );
  NAND2X0_HVT U3575 ( .A1(DP_OP_422J2_124_3477_n1246), .A2(
        DP_OP_422J2_124_3477_n1248), .Y(n1596) );
  NAND2X0_HVT U3576 ( .A1(DP_OP_422J2_124_3477_n1246), .A2(
        DP_OP_422J2_124_3477_n1250), .Y(n1597) );
  NAND2X0_HVT U3577 ( .A1(DP_OP_422J2_124_3477_n1248), .A2(
        DP_OP_422J2_124_3477_n1250), .Y(n1598) );
  NAND2X0_HVT U3578 ( .A1(DP_OP_422J2_124_3477_n377), .A2(
        DP_OP_422J2_124_3477_n420), .Y(n1599) );
  NAND2X0_HVT U3579 ( .A1(DP_OP_422J2_124_3477_n375), .A2(
        DP_OP_422J2_124_3477_n377), .Y(n1600) );
  NAND2X0_HVT U3580 ( .A1(DP_OP_422J2_124_3477_n375), .A2(
        DP_OP_422J2_124_3477_n420), .Y(n1601) );
  XOR3X2_HVT U3581 ( .A1(DP_OP_422J2_124_3477_n420), .A2(
        DP_OP_422J2_124_3477_n377), .A3(DP_OP_422J2_124_3477_n375), .Y(
        DP_OP_422J2_124_3477_n373) );
  NAND3X0_HVT U3582 ( .A1(n1602), .A2(n1603), .A3(n1604), .Y(
        DP_OP_422J2_124_3477_n1494) );
  NAND2X0_HVT U3583 ( .A1(DP_OP_422J2_124_3477_n1662), .A2(
        DP_OP_422J2_124_3477_n1696), .Y(n1602) );
  NAND2X0_HVT U3584 ( .A1(DP_OP_422J2_124_3477_n1662), .A2(
        DP_OP_422J2_124_3477_n1672), .Y(n1603) );
  NAND2X0_HVT U3585 ( .A1(DP_OP_422J2_124_3477_n1696), .A2(
        DP_OP_422J2_124_3477_n1672), .Y(n1604) );
  NAND3X0_HVT U3586 ( .A1(n1605), .A2(n1606), .A3(n1607), .Y(
        DP_OP_422J2_124_3477_n1282) );
  NAND2X0_HVT U3587 ( .A1(DP_OP_422J2_124_3477_n1486), .A2(
        DP_OP_422J2_124_3477_n1488), .Y(n1605) );
  NAND2X0_HVT U3588 ( .A1(DP_OP_422J2_124_3477_n1486), .A2(
        DP_OP_422J2_124_3477_n1498), .Y(n1606) );
  NAND2X0_HVT U3589 ( .A1(DP_OP_422J2_124_3477_n1488), .A2(
        DP_OP_422J2_124_3477_n1498), .Y(n1607) );
  NOR2X0_HVT U3590 ( .A1(DP_OP_422J2_124_3477_n2795), .A2(
        DP_OP_423J2_125_3477_n2804), .Y(DP_OP_422J2_124_3477_n2779) );
  INVX1_HVT U3591 ( .A(DP_OP_423J2_125_3477_n1728), .Y(
        DP_OP_423J2_125_3477_n1729) );
  INVX1_HVT U3592 ( .A(DP_OP_423J2_125_3477_n197), .Y(
        DP_OP_423J2_125_3477_n286) );
  INVX1_HVT U3593 ( .A(src_window[62]), .Y(DP_OP_423J2_125_3477_n2003) );
  INVX1_HVT U3594 ( .A(src_window[60]), .Y(DP_OP_423J2_125_3477_n2005) );
  INVX1_HVT U3595 ( .A(src_window[59]), .Y(DP_OP_423J2_125_3477_n2006) );
  INVX1_HVT U3596 ( .A(src_window[58]), .Y(DP_OP_423J2_125_3477_n2007) );
  INVX1_HVT U3597 ( .A(src_window[57]), .Y(DP_OP_423J2_125_3477_n2008) );
  INVX1_HVT U3598 ( .A(src_window[77]), .Y(DP_OP_423J2_125_3477_n2048) );
  INVX1_HVT U3599 ( .A(src_window[74]), .Y(DP_OP_423J2_125_3477_n2051) );
  INVX1_HVT U3600 ( .A(src_window[73]), .Y(DP_OP_423J2_125_3477_n2052) );
  INVX1_HVT U3601 ( .A(src_window[72]), .Y(DP_OP_423J2_125_3477_n2053) );
  INVX1_HVT U3602 ( .A(src_window[103]), .Y(DP_OP_423J2_125_3477_n2090) );
  INVX1_HVT U3603 ( .A(src_window[99]), .Y(DP_OP_423J2_125_3477_n2094) );
  INVX1_HVT U3604 ( .A(src_window[97]), .Y(DP_OP_423J2_125_3477_n2096) );
  INVX1_HVT U3605 ( .A(src_window[96]), .Y(DP_OP_423J2_125_3477_n2097) );
  INVX1_HVT U3606 ( .A(src_window[118]), .Y(DP_OP_423J2_125_3477_n2135) );
  INVX1_HVT U3607 ( .A(src_window[113]), .Y(DP_OP_423J2_125_3477_n2140) );
  INVX1_HVT U3608 ( .A(src_window[135]), .Y(DP_OP_423J2_125_3477_n2178) );
  INVX1_HVT U3609 ( .A(src_window[131]), .Y(DP_OP_423J2_125_3477_n2182) );
  INVX1_HVT U3610 ( .A(src_window[128]), .Y(DP_OP_423J2_125_3477_n2185) );
  INVX1_HVT U3611 ( .A(src_window[159]), .Y(DP_OP_423J2_125_3477_n2222) );
  INVX1_HVT U3612 ( .A(src_window[156]), .Y(DP_OP_423J2_125_3477_n2225) );
  INVX1_HVT U3613 ( .A(src_window[154]), .Y(DP_OP_423J2_125_3477_n2227) );
  INVX1_HVT U3614 ( .A(src_window[153]), .Y(DP_OP_423J2_125_3477_n2228) );
  INVX1_HVT U3615 ( .A(src_window[152]), .Y(DP_OP_423J2_125_3477_n2229) );
  INVX1_HVT U3616 ( .A(src_window[174]), .Y(DP_OP_423J2_125_3477_n2267) );
  INVX1_HVT U3617 ( .A(src_window[173]), .Y(DP_OP_423J2_125_3477_n2268) );
  INVX1_HVT U3618 ( .A(src_window[172]), .Y(DP_OP_423J2_125_3477_n2269) );
  INVX1_HVT U3619 ( .A(src_window[170]), .Y(DP_OP_423J2_125_3477_n2271) );
  INVX1_HVT U3620 ( .A(src_window[169]), .Y(DP_OP_423J2_125_3477_n2272) );
  INVX1_HVT U3621 ( .A(src_window[168]), .Y(DP_OP_423J2_125_3477_n2273) );
  INVX1_HVT U3622 ( .A(conv_weight_box[36]), .Y(DP_OP_423J2_125_3477_n2277) );
  INVX1_HVT U3623 ( .A(src_window[199]), .Y(DP_OP_423J2_125_3477_n2310) );
  INVX1_HVT U3624 ( .A(src_window[198]), .Y(DP_OP_423J2_125_3477_n2311) );
  INVX1_HVT U3625 ( .A(src_window[194]), .Y(DP_OP_423J2_125_3477_n2315) );
  INVX1_HVT U3626 ( .A(src_window[193]), .Y(DP_OP_423J2_125_3477_n2316) );
  INVX1_HVT U3627 ( .A(src_window[192]), .Y(DP_OP_423J2_125_3477_n2317) );
  INVX1_HVT U3628 ( .A(src_window[215]), .Y(DP_OP_423J2_125_3477_n2354) );
  INVX1_HVT U3629 ( .A(src_window[208]), .Y(DP_OP_423J2_125_3477_n2361) );
  INVX1_HVT U3630 ( .A(src_window[230]), .Y(DP_OP_423J2_125_3477_n2399) );
  INVX1_HVT U3631 ( .A(src_window[229]), .Y(DP_OP_423J2_125_3477_n2400) );
  INVX1_HVT U3632 ( .A(src_window[228]), .Y(DP_OP_423J2_125_3477_n2401) );
  INVX1_HVT U3633 ( .A(src_window[225]), .Y(DP_OP_423J2_125_3477_n2404) );
  INVX1_HVT U3634 ( .A(src_window[224]), .Y(DP_OP_423J2_125_3477_n2405) );
  INVX1_HVT U3635 ( .A(src_window[250]), .Y(DP_OP_423J2_125_3477_n2447) );
  INVX1_HVT U3636 ( .A(src_window[249]), .Y(DP_OP_423J2_125_3477_n2448) );
  INVX1_HVT U3637 ( .A(src_window[264]), .Y(DP_OP_423J2_125_3477_n2493) );
  INVX1_HVT U3638 ( .A(src_window[278]), .Y(DP_OP_423J2_125_3477_n2531) );
  INVX1_HVT U3639 ( .A(src_window[273]), .Y(DP_OP_423J2_125_3477_n2536) );
  INVX1_HVT U3640 ( .A(src_window[272]), .Y(DP_OP_423J2_125_3477_n2537) );
  INVX1_HVT U3641 ( .A(src_window[258]), .Y(DP_OP_423J2_125_3477_n2579) );
  INVX1_HVT U3642 ( .A(src_window[256]), .Y(DP_OP_423J2_125_3477_n2581) );
  INVX1_HVT U3643 ( .A(src_window[247]), .Y(DP_OP_423J2_125_3477_n2618) );
  INVX1_HVT U3644 ( .A(src_window[246]), .Y(DP_OP_423J2_125_3477_n2619) );
  INVX1_HVT U3645 ( .A(src_window[245]), .Y(DP_OP_423J2_125_3477_n2620) );
  INVX1_HVT U3646 ( .A(src_window[244]), .Y(DP_OP_423J2_125_3477_n2621) );
  INVX1_HVT U3647 ( .A(src_window[243]), .Y(DP_OP_423J2_125_3477_n2622) );
  INVX1_HVT U3648 ( .A(src_window[242]), .Y(DP_OP_423J2_125_3477_n2623) );
  INVX1_HVT U3649 ( .A(src_window[241]), .Y(DP_OP_423J2_125_3477_n2624) );
  INVX1_HVT U3650 ( .A(src_window[240]), .Y(DP_OP_423J2_125_3477_n2625) );
  INVX1_HVT U3651 ( .A(src_window[220]), .Y(DP_OP_423J2_125_3477_n2665) );
  INVX1_HVT U3652 ( .A(src_window[219]), .Y(DP_OP_423J2_125_3477_n2666) );
  INVX1_HVT U3653 ( .A(src_window[218]), .Y(DP_OP_423J2_125_3477_n2667) );
  INVX1_HVT U3654 ( .A(src_window[217]), .Y(DP_OP_423J2_125_3477_n2668) );
  INVX1_HVT U3655 ( .A(src_window[216]), .Y(DP_OP_423J2_125_3477_n2669) );
  INVX1_HVT U3656 ( .A(src_window[207]), .Y(DP_OP_423J2_125_3477_n2706) );
  INVX1_HVT U3657 ( .A(src_window[205]), .Y(DP_OP_423J2_125_3477_n2708) );
  INVX1_HVT U3658 ( .A(src_window[201]), .Y(DP_OP_423J2_125_3477_n2712) );
  INVX1_HVT U3659 ( .A(src_window[200]), .Y(DP_OP_423J2_125_3477_n2713) );
  INVX1_HVT U3660 ( .A(src_window[183]), .Y(DP_OP_423J2_125_3477_n2750) );
  INVX1_HVT U3661 ( .A(src_window[182]), .Y(DP_OP_423J2_125_3477_n2751) );
  INVX1_HVT U3662 ( .A(src_window[179]), .Y(DP_OP_423J2_125_3477_n2754) );
  INVX1_HVT U3663 ( .A(src_window[177]), .Y(DP_OP_423J2_125_3477_n2756) );
  INVX1_HVT U3664 ( .A(src_window[176]), .Y(DP_OP_423J2_125_3477_n2757) );
  INVX1_HVT U3665 ( .A(src_window[167]), .Y(DP_OP_423J2_125_3477_n2794) );
  INVX1_HVT U3666 ( .A(src_window[166]), .Y(DP_OP_423J2_125_3477_n2795) );
  INVX1_HVT U3667 ( .A(src_window[163]), .Y(DP_OP_423J2_125_3477_n2798) );
  INVX1_HVT U3668 ( .A(src_window[162]), .Y(DP_OP_423J2_125_3477_n2799) );
  INVX1_HVT U3669 ( .A(src_window[161]), .Y(DP_OP_423J2_125_3477_n2800) );
  INVX1_HVT U3670 ( .A(src_window[160]), .Y(DP_OP_423J2_125_3477_n2801) );
  INVX1_HVT U3671 ( .A(src_window[148]), .Y(DP_OP_423J2_125_3477_n2841) );
  INVX1_HVT U3672 ( .A(src_window[147]), .Y(DP_OP_423J2_125_3477_n2842) );
  INVX1_HVT U3673 ( .A(src_window[146]), .Y(DP_OP_423J2_125_3477_n2843) );
  INVX1_HVT U3674 ( .A(src_window[145]), .Y(DP_OP_423J2_125_3477_n2844) );
  INVX1_HVT U3675 ( .A(src_window[144]), .Y(DP_OP_423J2_125_3477_n2845) );
  INVX1_HVT U3676 ( .A(conv_weight_box[26]), .Y(DP_OP_423J2_125_3477_n2849) );
  INVX1_HVT U3677 ( .A(src_window[123]), .Y(DP_OP_423J2_125_3477_n2886) );
  INVX1_HVT U3678 ( .A(src_window[122]), .Y(DP_OP_423J2_125_3477_n2887) );
  INVX1_HVT U3679 ( .A(src_window[120]), .Y(DP_OP_423J2_125_3477_n2889) );
  INVX1_HVT U3680 ( .A(src_window[106]), .Y(DP_OP_423J2_125_3477_n2931) );
  INVX1_HVT U3681 ( .A(src_window[105]), .Y(DP_OP_423J2_125_3477_n2932) );
  INVX1_HVT U3682 ( .A(src_window[84]), .Y(DP_OP_423J2_125_3477_n2973) );
  INVX1_HVT U3683 ( .A(src_window[81]), .Y(DP_OP_423J2_125_3477_n2976) );
  INVX1_HVT U3684 ( .A(src_window[71]), .Y(DP_OP_423J2_125_3477_n3014) );
  INVX1_HVT U3685 ( .A(src_window[66]), .Y(DP_OP_423J2_125_3477_n3019) );
  INVX1_HVT U3686 ( .A(src_window[64]), .Y(DP_OP_423J2_125_3477_n3021) );
  INVX1_HVT U3687 ( .A(DP_OP_423J2_125_3477_n302), .Y(
        DP_OP_423J2_125_3477_n303) );
  INVX1_HVT U3688 ( .A(DP_OP_423J2_125_3477_n304), .Y(
        DP_OP_423J2_125_3477_n305) );
  INVX1_HVT U3689 ( .A(src_window[55]), .Y(DP_OP_423J2_125_3477_n3056) );
  INVX1_HVT U3690 ( .A(src_window[54]), .Y(DP_OP_423J2_125_3477_n3057) );
  INVX1_HVT U3691 ( .A(src_window[52]), .Y(DP_OP_423J2_125_3477_n3059) );
  INVX1_HVT U3692 ( .A(src_window[51]), .Y(DP_OP_423J2_125_3477_n3060) );
  INVX1_HVT U3693 ( .A(src_window[50]), .Y(DP_OP_423J2_125_3477_n3061) );
  INVX1_HVT U3694 ( .A(src_window[49]), .Y(DP_OP_423J2_125_3477_n3062) );
  INVX1_HVT U3695 ( .A(src_window[48]), .Y(DP_OP_423J2_125_3477_n3063) );
  INVX1_HVT U3696 ( .A(conv_weight_box[0]), .Y(DP_OP_423J2_125_3477_n3066) );
  INVX1_HVT U3697 ( .A(DP_OP_423J2_125_3477_n306), .Y(
        DP_OP_423J2_125_3477_n307) );
  INVX1_HVT U3698 ( .A(DP_OP_423J2_125_3477_n308), .Y(
        DP_OP_423J2_125_3477_n309) );
  INVX1_HVT U3699 ( .A(DP_OP_423J2_125_3477_n310), .Y(
        DP_OP_423J2_125_3477_n311) );
  INVX1_HVT U3700 ( .A(DP_OP_423J2_125_3477_n314), .Y(
        DP_OP_423J2_125_3477_n315) );
  INVX1_HVT U3701 ( .A(DP_OP_423J2_125_3477_n316), .Y(
        DP_OP_423J2_125_3477_n317) );
  INVX1_HVT U3702 ( .A(DP_OP_423J2_125_3477_n318), .Y(
        DP_OP_423J2_125_3477_n319) );
  INVX1_HVT U3703 ( .A(DP_OP_423J2_125_3477_n320), .Y(
        DP_OP_423J2_125_3477_n321) );
  INVX1_HVT U3704 ( .A(DP_OP_423J2_125_3477_n322), .Y(
        DP_OP_423J2_125_3477_n323) );
  INVX1_HVT U3705 ( .A(DP_OP_423J2_125_3477_n324), .Y(
        DP_OP_423J2_125_3477_n325) );
  INVX1_HVT U3706 ( .A(DP_OP_423J2_125_3477_n326), .Y(
        DP_OP_423J2_125_3477_n327) );
  INVX1_HVT U3707 ( .A(DP_OP_423J2_125_3477_n328), .Y(
        DP_OP_423J2_125_3477_n329) );
  INVX1_HVT U3708 ( .A(DP_OP_423J2_125_3477_n330), .Y(
        DP_OP_423J2_125_3477_n331) );
  INVX1_HVT U3709 ( .A(DP_OP_423J2_125_3477_n510), .Y(
        DP_OP_423J2_125_3477_n511) );
  INVX1_HVT U3710 ( .A(DP_OP_423J2_125_3477_n820), .Y(
        DP_OP_423J2_125_3477_n821) );
  INVX1_HVT U3711 ( .A(DP_OP_423J2_125_3477_n95), .Y(DP_OP_423J2_125_3477_n93)
         );
  AO21X1_HVT U3712 ( .A1(DP_OP_423J2_125_3477_n4), .A2(n1677), .A3(n1528), .Y(
        n1608) );
  XOR3X2_HVT U3713 ( .A1(DP_OP_423J2_125_3477_n379), .A2(
        DP_OP_423J2_125_3477_n424), .A3(DP_OP_423J2_125_3477_n422), .Y(
        DP_OP_423J2_125_3477_n375) );
  OR2X1_HVT U3714 ( .A1(DP_OP_423J2_125_3477_n424), .A2(
        DP_OP_423J2_125_3477_n379), .Y(n1613) );
  AO22X1_HVT U3715 ( .A1(DP_OP_423J2_125_3477_n379), .A2(
        DP_OP_423J2_125_3477_n424), .A3(DP_OP_423J2_125_3477_n422), .A4(n1613), 
        .Y(DP_OP_423J2_125_3477_n374) );
  NAND2X0_HVT U3716 ( .A1(n1436), .A2(n1678), .Y(n1618) );
  NAND2X0_HVT U3717 ( .A1(n1619), .A2(n1616), .Y(n1620) );
  AO22X1_HVT U3718 ( .A1(n1615), .A2(n1620), .A3(DP_OP_423J2_125_3477_n68), 
        .A4(n1616), .Y(n1621) );
  NAND3X0_HVT U3719 ( .A1(n1617), .A2(n1618), .A3(n1621), .Y(n_conv2_sum_b[28]) );
  NAND2X0_HVT U3720 ( .A1(DP_OP_423J2_125_3477_n177), .A2(
        DP_OP_423J2_125_3477_n142), .Y(n1624) );
  NAND2X0_HVT U3721 ( .A1(n1624), .A2(DP_OP_423J2_125_3477_n145), .Y(n1625) );
  NAND2X0_HVT U3722 ( .A1(n1628), .A2(n1626), .Y(n1629) );
  AO22X1_HVT U3723 ( .A1(n1623), .A2(n1629), .A3(n1630), .A4(n1626), .Y(n1631)
         );
  NAND2X0_HVT U3724 ( .A1(n1436), .A2(n1679), .Y(n1632) );
  NAND3X0_HVT U3725 ( .A1(n1627), .A2(n1631), .A3(n1632), .Y(n_conv2_sum_b[23]) );
  NAND2X0_HVT U3726 ( .A1(n1611), .A2(n1686), .Y(n1633) );
  XOR3X2_HVT U3727 ( .A1(DP_OP_423J2_125_3477_n1830), .A2(
        DP_OP_423J2_125_3477_n1828), .A3(DP_OP_423J2_125_3477_n1808), .Y(
        DP_OP_423J2_125_3477_n1657) );
  FADDX1_HVT U3728 ( .A(DP_OP_423J2_125_3477_n1828), .B(
        DP_OP_423J2_125_3477_n1830), .CI(DP_OP_423J2_125_3477_n1808), .CO(
        DP_OP_423J2_125_3477_n1656) );
  OA21X1_HVT U3729 ( .A1(DP_OP_423J2_125_3477_n261), .A2(
        DP_OP_423J2_125_3477_n259), .A3(DP_OP_423J2_125_3477_n260), .Y(n1634)
         );
  OA21X1_HVT U3730 ( .A1(n1634), .A2(DP_OP_423J2_125_3477_n256), .A3(
        DP_OP_423J2_125_3477_n257), .Y(DP_OP_423J2_125_3477_n253) );
  OR2X1_HVT U3731 ( .A1(DP_OP_423J2_125_3477_n1215), .A2(
        DP_OP_423J2_125_3477_n1213), .Y(n1636) );
  NAND2X0_HVT U3732 ( .A1(DP_OP_423J2_125_3477_n151), .A2(
        DP_OP_423J2_125_3477_n4), .Y(n1637) );
  NAND2X0_HVT U3733 ( .A1(n1637), .A2(n1638), .Y(n1639) );
  NAND2X0_HVT U3734 ( .A1(conv_weight_box[35]), .A2(src_window[160]), .Y(n1642) );
  NAND2X0_HVT U3735 ( .A1(n1640), .A2(n1641), .Y(n1643) );
  NAND2X0_HVT U3736 ( .A1(n1643), .A2(n1642), .Y(n1644) );
  OR2X1_HVT U3737 ( .A1(n1641), .A2(n1640), .Y(n1645) );
  NAND2X0_HVT U3738 ( .A1(n1644), .A2(n1645), .Y(DP_OP_423J2_125_3477_n1714)
         );
  AND2X1_HVT U3739 ( .A1(conv_weight_box[66]), .A2(src_window[274]), .Y(n1647)
         );
  NAND2X0_HVT U3740 ( .A1(n1650), .A2(n1646), .Y(n1651) );
  AO22X1_HVT U3741 ( .A1(n1649), .A2(n1647), .A3(n1651), .A4(n1652), .Y(
        DP_OP_423J2_125_3477_n1802) );
  NAND2X0_HVT U3742 ( .A1(n1425), .A2(conv2_sum_b[1]), .Y(n1653) );
  AND2X1_HVT U3743 ( .A1(conv_weight_box[2]), .A2(src_window[57]), .Y(n1654)
         );
  AO21X1_HVT U3744 ( .A1(DP_OP_423J2_125_3477_n4), .A2(
        DP_OP_423J2_125_3477_n187), .A3(DP_OP_423J2_125_3477_n188), .Y(n1659)
         );
  AO21X1_HVT U3745 ( .A1(DP_OP_423J2_125_3477_n4), .A2(
        DP_OP_423J2_125_3477_n107), .A3(DP_OP_423J2_125_3477_n108), .Y(n1660)
         );
  AO21X1_HVT U3746 ( .A1(DP_OP_423J2_125_3477_n4), .A2(
        DP_OP_423J2_125_3477_n176), .A3(DP_OP_423J2_125_3477_n177), .Y(n1661)
         );
  AO21X1_HVT U3747 ( .A1(DP_OP_423J2_125_3477_n4), .A2(
        DP_OP_423J2_125_3477_n138), .A3(n1625), .Y(n1662) );
  AO21X1_HVT U3748 ( .A1(DP_OP_423J2_125_3477_n4), .A2(
        DP_OP_423J2_125_3477_n158), .A3(DP_OP_423J2_125_3477_n159), .Y(n1663)
         );
  AO21X1_HVT U3749 ( .A1(DP_OP_423J2_125_3477_n4), .A2(
        DP_OP_423J2_125_3477_n49), .A3(DP_OP_423J2_125_3477_n50), .Y(n1664) );
  AND2X1_HVT U3750 ( .A1(conv_weight_box[64]), .A2(src_window[265]), .Y(
        DP_OP_423J2_125_3477_n2468) );
  OR2X1_HVT U3751 ( .A1(DP_OP_423J2_125_3477_n3029), .A2(
        DP_OP_423J2_125_3477_n2502), .Y(DP_OP_423J2_125_3477_n1210) );
  OR2X1_HVT U3752 ( .A1(DP_OP_423J2_125_3477_n648), .A2(
        DP_OP_423J2_125_3477_n513), .Y(n1611) );
  AO21X1_HVT U3753 ( .A1(DP_OP_423J2_125_3477_n4), .A2(
        DP_OP_423J2_125_3477_n54), .A3(DP_OP_423J2_125_3477_n55), .Y(n1667) );
  OR2X1_HVT U3754 ( .A1(DP_OP_423J2_125_3477_n512), .A2(n1476), .Y(n1622) );
  OR2X1_HVT U3755 ( .A1(DP_OP_423J2_125_3477_n302), .A2(n1669), .Y(n1668) );
  OR2X1_HVT U3756 ( .A1(DP_OP_423J2_125_3477_n304), .A2(
        DP_OP_423J2_125_3477_n303), .Y(n1670) );
  OR2X1_HVT U3757 ( .A1(DP_OP_423J2_125_3477_n308), .A2(
        DP_OP_423J2_125_3477_n307), .Y(n1671) );
  OR2X1_HVT U3758 ( .A1(DP_OP_423J2_125_3477_n312), .A2(
        DP_OP_423J2_125_3477_n311), .Y(n1672) );
  OR2X1_HVT U3759 ( .A1(DP_OP_423J2_125_3477_n318), .A2(
        DP_OP_423J2_125_3477_n317), .Y(n1673) );
  INVX1_HVT U3760 ( .A(DP_OP_423J2_125_3477_n68), .Y(n1615) );
  OR2X1_HVT U3761 ( .A1(DP_OP_423J2_125_3477_n171), .A2(
        DP_OP_423J2_125_3477_n178), .Y(n1674) );
  INVX1_HVT U3762 ( .A(DP_OP_423J2_125_3477_n209), .Y(n1656) );
  OR2X1_HVT U3763 ( .A1(DP_OP_423J2_125_3477_n1733), .A2(
        DP_OP_423J2_125_3477_n1731), .Y(n1676) );
  AND2X1_HVT U3764 ( .A1(DP_OP_423J2_125_3477_n67), .A2(
        DP_OP_423J2_125_3477_n9), .Y(n1678) );
  OA21X1_HVT U3765 ( .A1(DP_OP_423J2_125_3477_n171), .A2(
        DP_OP_423J2_125_3477_n179), .A3(DP_OP_423J2_125_3477_n174), .Y(n1681)
         );
  AND2X1_HVT U3766 ( .A1(DP_OP_423J2_125_3477_n49), .A2(n1670), .Y(n1682) );
  INVX1_HVT U3767 ( .A(conv_weight_box[35]), .Y(DP_OP_423J2_125_3477_n2802) );
  INVX1_HVT U3768 ( .A(conv_weight_box[15]), .Y(DP_OP_423J2_125_3477_n2098) );
  INVX1_HVT U3769 ( .A(DP_OP_423J2_125_3477_n253), .Y(n1635) );
  OA21X1_HVT U3770 ( .A1(DP_OP_423J2_125_3477_n153), .A2(
        DP_OP_423J2_125_3477_n161), .A3(DP_OP_423J2_125_3477_n156), .Y(n1638)
         );
  OA21X1_HVT U3771 ( .A1(DP_OP_423J2_125_3477_n133), .A2(
        DP_OP_423J2_125_3477_n141), .A3(DP_OP_423J2_125_3477_n136), .Y(n1658)
         );
  OA21X1_HVT U3772 ( .A1(DP_OP_423J2_125_3477_n124), .A2(
        DP_OP_423J2_125_3477_n141), .A3(DP_OP_423J2_125_3477_n125), .Y(n1623)
         );
  INVX1_HVT U3773 ( .A(DP_OP_423J2_125_3477_n14), .Y(n1626) );
  AND2X1_HVT U3774 ( .A1(DP_OP_423J2_125_3477_n122), .A2(
        DP_OP_423J2_125_3477_n14), .Y(n1679) );
  INVX1_HVT U3775 ( .A(DP_OP_423J2_125_3477_n9), .Y(n1616) );
  OA21X1_HVT U3776 ( .A1(DP_OP_423J2_125_3477_n209), .A2(
        DP_OP_423J2_125_3477_n217), .A3(DP_OP_423J2_125_3477_n210), .Y(n1675)
         );
  INVX1_HVT U3777 ( .A(conv_weight_box[5]), .Y(DP_OP_423J2_125_3477_n3025) );
  INVX1_HVT U3778 ( .A(conv_weight_box[41]), .Y(DP_OP_423J2_125_3477_n2321) );
  XNOR2X1_HVT U3779 ( .A1(n1653), .A2(n1654), .Y(DP_OP_423J2_125_3477_n1897)
         );
  OR2X1_HVT U3780 ( .A1(DP_OP_423J2_125_3477_n372), .A2(
        DP_OP_423J2_125_3477_n351), .Y(n1655) );
  INVX1_HVT U3781 ( .A(DP_OP_423J2_125_3477_n338), .Y(
        DP_OP_423J2_125_3477_n339) );
  INVX1_HVT U3782 ( .A(conv_weight_box[55]), .Y(DP_OP_423J2_125_3477_n2627) );
  INVX1_HVT U3783 ( .A(conv_weight_box[1]), .Y(DP_OP_423J2_125_3477_n3065) );
  INVX1_HVT U3784 ( .A(conv_weight_box[14]), .Y(DP_OP_423J2_125_3477_n2099) );
  INVX1_HVT U3785 ( .A(conv_weight_box[48]), .Y(DP_OP_423J2_125_3477_n2362) );
  INVX1_HVT U3786 ( .A(conv_weight_box[44]), .Y(DP_OP_423J2_125_3477_n2318) );
  INVX1_HVT U3787 ( .A(conv_weight_box[23]), .Y(DP_OP_423J2_125_3477_n2890) );
  NAND3X0_HVT U3788 ( .A1(n1683), .A2(n1684), .A3(n1685), .Y(
        DP_OP_423J2_125_3477_n1282) );
  NAND2X0_HVT U3789 ( .A1(DP_OP_423J2_125_3477_n1488), .A2(
        DP_OP_423J2_125_3477_n1486), .Y(n1683) );
  NAND2X0_HVT U3790 ( .A1(DP_OP_423J2_125_3477_n1488), .A2(
        DP_OP_423J2_125_3477_n1498), .Y(n1684) );
  NAND2X0_HVT U3791 ( .A1(DP_OP_423J2_125_3477_n1486), .A2(
        DP_OP_423J2_125_3477_n1498), .Y(n1685) );
  XOR3X2_HVT U3792 ( .A1(DP_OP_423J2_125_3477_n1486), .A2(
        DP_OP_423J2_125_3477_n1498), .A3(DP_OP_423J2_125_3477_n1488), .Y(
        DP_OP_423J2_125_3477_n1283) );
  AND2X1_HVT U3793 ( .A1(DP_OP_423J2_125_3477_n649), .A2(
        DP_OP_423J2_125_3477_n822), .Y(n1686) );
  AND2X1_HVT U3794 ( .A1(n1672), .A2(DP_OP_423J2_125_3477_n89), .Y(n1687) );
  AO21X1_HVT U3795 ( .A1(DP_OP_423J2_125_3477_n4), .A2(
        DP_OP_423J2_125_3477_n91), .A3(DP_OP_423J2_125_3477_n92), .Y(n1688) );
  XOR2X2_HVT U3796 ( .A1(n1688), .A2(n1687), .Y(n_conv2_sum_b[26]) );
  OR2X1_HVT U3797 ( .A1(DP_OP_423J2_125_3477_n822), .A2(
        DP_OP_423J2_125_3477_n649), .Y(n1612) );
  XOR3X2_HVT U3798 ( .A1(DP_OP_423J2_125_3477_n2251), .A2(
        DP_OP_423J2_125_3477_n2816), .A3(DP_OP_423J2_125_3477_n2244), .Y(
        DP_OP_423J2_125_3477_n967) );
  NAND3X0_HVT U3799 ( .A1(n1689), .A2(n1690), .A3(n1691), .Y(
        DP_OP_423J2_125_3477_n1492) );
  NAND2X0_HVT U3800 ( .A1(DP_OP_423J2_125_3477_n1692), .A2(
        DP_OP_423J2_125_3477_n1668), .Y(n1689) );
  NAND2X0_HVT U3801 ( .A1(DP_OP_423J2_125_3477_n1692), .A2(
        DP_OP_423J2_125_3477_n1694), .Y(n1690) );
  NAND2X0_HVT U3802 ( .A1(DP_OP_423J2_125_3477_n1668), .A2(
        DP_OP_423J2_125_3477_n1694), .Y(n1691) );
  NAND2X0_HVT U3803 ( .A1(DP_OP_423J2_125_3477_n527), .A2(
        DP_OP_423J2_125_3477_n658), .Y(n1692) );
  NAND2X0_HVT U3804 ( .A1(DP_OP_423J2_125_3477_n527), .A2(
        DP_OP_423J2_125_3477_n525), .Y(n1693) );
  NAND2X0_HVT U3805 ( .A1(DP_OP_423J2_125_3477_n658), .A2(
        DP_OP_423J2_125_3477_n525), .Y(n1694) );
  XOR3X2_HVT U3806 ( .A1(DP_OP_423J2_125_3477_n658), .A2(
        DP_OP_423J2_125_3477_n527), .A3(DP_OP_423J2_125_3477_n525), .Y(
        DP_OP_423J2_125_3477_n519) );
  NAND3X0_HVT U3807 ( .A1(n1695), .A2(n1696), .A3(n1697), .Y(
        DP_OP_423J2_125_3477_n1256) );
  NAND2X0_HVT U3808 ( .A1(DP_OP_423J2_125_3477_n1289), .A2(
        DP_OP_423J2_125_3477_n1291), .Y(n1695) );
  NAND2X0_HVT U3809 ( .A1(DP_OP_423J2_125_3477_n1289), .A2(
        DP_OP_423J2_125_3477_n1458), .Y(n1696) );
  NAND2X0_HVT U3810 ( .A1(DP_OP_423J2_125_3477_n1291), .A2(
        DP_OP_423J2_125_3477_n1458), .Y(n1697) );
  XOR3X2_HVT U3811 ( .A1(DP_OP_423J2_125_3477_n1289), .A2(
        DP_OP_423J2_125_3477_n1291), .A3(DP_OP_423J2_125_3477_n1458), .Y(
        DP_OP_423J2_125_3477_n1257) );
  NAND3X0_HVT U3812 ( .A1(n1698), .A2(n1699), .A3(n1700), .Y(
        DP_OP_423J2_125_3477_n442) );
  NAND2X0_HVT U3813 ( .A1(DP_OP_423J2_125_3477_n552), .A2(
        DP_OP_423J2_125_3477_n457), .Y(n1698) );
  NAND2X0_HVT U3814 ( .A1(DP_OP_423J2_125_3477_n552), .A2(
        DP_OP_423J2_125_3477_n550), .Y(n1699) );
  NAND2X0_HVT U3815 ( .A1(DP_OP_423J2_125_3477_n457), .A2(
        DP_OP_423J2_125_3477_n550), .Y(n1700) );
  XOR3X2_HVT U3816 ( .A1(DP_OP_423J2_125_3477_n457), .A2(
        DP_OP_423J2_125_3477_n552), .A3(DP_OP_423J2_125_3477_n550), .Y(
        DP_OP_423J2_125_3477_n443) );
  NAND3X0_HVT U3817 ( .A1(n1701), .A2(n1702), .A3(n1703), .Y(
        DP_OP_423J2_125_3477_n834) );
  NAND2X0_HVT U3818 ( .A1(DP_OP_423J2_125_3477_n847), .A2(
        DP_OP_423J2_125_3477_n1034), .Y(n1701) );
  NAND2X0_HVT U3819 ( .A1(DP_OP_423J2_125_3477_n847), .A2(
        DP_OP_423J2_125_3477_n1036), .Y(n1702) );
  NAND2X0_HVT U3820 ( .A1(DP_OP_423J2_125_3477_n1034), .A2(
        DP_OP_423J2_125_3477_n1036), .Y(n1703) );
  XOR3X2_HVT U3821 ( .A1(DP_OP_423J2_125_3477_n1034), .A2(
        DP_OP_423J2_125_3477_n847), .A3(DP_OP_423J2_125_3477_n1036), .Y(
        DP_OP_423J2_125_3477_n835) );
  NAND3X0_HVT U3822 ( .A1(n1704), .A2(n1705), .A3(n1706), .Y(
        DP_OP_423J2_125_3477_n906) );
  NAND2X0_HVT U3823 ( .A1(DP_OP_423J2_125_3477_n981), .A2(
        DP_OP_423J2_125_3477_n983), .Y(n1704) );
  NAND2X0_HVT U3824 ( .A1(DP_OP_423J2_125_3477_n981), .A2(
        DP_OP_423J2_125_3477_n979), .Y(n1705) );
  NAND2X0_HVT U3825 ( .A1(DP_OP_423J2_125_3477_n983), .A2(
        DP_OP_423J2_125_3477_n979), .Y(n1706) );
  XOR3X2_HVT U3826 ( .A1(DP_OP_423J2_125_3477_n983), .A2(
        DP_OP_423J2_125_3477_n981), .A3(DP_OP_423J2_125_3477_n979), .Y(
        DP_OP_423J2_125_3477_n907) );
  NAND2X0_HVT U3827 ( .A1(DP_OP_423J2_125_3477_n969), .A2(
        DP_OP_423J2_125_3477_n977), .Y(n1707) );
  NAND2X0_HVT U3828 ( .A1(DP_OP_423J2_125_3477_n953), .A2(
        DP_OP_423J2_125_3477_n977), .Y(n1708) );
  AND2X1_HVT U3829 ( .A1(DP_OP_423J2_125_3477_n276), .A2(
        DP_OP_423J2_125_3477_n98), .Y(n1709) );
  AO21X1_HVT U3830 ( .A1(DP_OP_423J2_125_3477_n4), .A2(
        DP_OP_423J2_125_3477_n100), .A3(DP_OP_423J2_125_3477_n101), .Y(n1710)
         );
  XOR2X2_HVT U3831 ( .A1(n1710), .A2(n1709), .Y(n_conv2_sum_b[25]) );
  INVX1_HVT U3832 ( .A(DP_OP_424J2_126_3477_n1728), .Y(
        DP_OP_424J2_126_3477_n1729) );
  INVX1_HVT U3833 ( .A(DP_OP_424J2_126_3477_n197), .Y(
        DP_OP_424J2_126_3477_n286) );
  INVX1_HVT U3834 ( .A(src_window[23]), .Y(DP_OP_424J2_126_3477_n2002) );
  INVX1_HVT U3835 ( .A(src_window[22]), .Y(DP_OP_424J2_126_3477_n2003) );
  INVX1_HVT U3836 ( .A(src_window[21]), .Y(DP_OP_424J2_126_3477_n2004) );
  INVX1_HVT U3837 ( .A(src_window[20]), .Y(DP_OP_424J2_126_3477_n2005) );
  INVX1_HVT U3838 ( .A(src_window[19]), .Y(DP_OP_424J2_126_3477_n2006) );
  INVX1_HVT U3839 ( .A(DP_OP_424J2_126_3477_n203), .Y(
        DP_OP_424J2_126_3477_n201) );
  INVX1_HVT U3840 ( .A(conv_weight_box[3]), .Y(DP_OP_424J2_126_3477_n2011) );
  INVX1_HVT U3841 ( .A(src_window[34]), .Y(DP_OP_424J2_126_3477_n2051) );
  INVX1_HVT U3842 ( .A(conv_weight_box[9]), .Y(DP_OP_424J2_126_3477_n2056) );
  INVX1_HVT U3843 ( .A(src_window[63]), .Y(DP_OP_424J2_126_3477_n2090) );
  INVX1_HVT U3844 ( .A(src_window[61]), .Y(DP_OP_424J2_126_3477_n2092) );
  INVX1_HVT U3845 ( .A(src_window[58]), .Y(DP_OP_424J2_126_3477_n2095) );
  INVX1_HVT U3846 ( .A(conv_weight_box[14]), .Y(DP_OP_424J2_126_3477_n2099) );
  INVX1_HVT U3847 ( .A(conv_weight_box[13]), .Y(DP_OP_424J2_126_3477_n2100) );
  INVX1_HVT U3848 ( .A(src_window[77]), .Y(DP_OP_424J2_126_3477_n2136) );
  INVX1_HVT U3849 ( .A(src_window[75]), .Y(DP_OP_424J2_126_3477_n2138) );
  INVX1_HVT U3850 ( .A(conv_weight_box[19]), .Y(DP_OP_424J2_126_3477_n2144) );
  INVX1_HVT U3851 ( .A(src_window[89]), .Y(DP_OP_424J2_126_3477_n2184) );
  INVX1_HVT U3852 ( .A(src_window[88]), .Y(DP_OP_424J2_126_3477_n2185) );
  INVX1_HVT U3853 ( .A(conv_weight_box[25]), .Y(DP_OP_424J2_126_3477_n2186) );
  INVX1_HVT U3854 ( .A(conv_weight_box[24]), .Y(DP_OP_424J2_126_3477_n2189) );
  INVX1_HVT U3855 ( .A(src_window[119]), .Y(DP_OP_424J2_126_3477_n2222) );
  INVX1_HVT U3856 ( .A(src_window[134]), .Y(DP_OP_424J2_126_3477_n2267) );
  INVX1_HVT U3857 ( .A(src_window[133]), .Y(DP_OP_424J2_126_3477_n2268) );
  INVX1_HVT U3858 ( .A(src_window[132]), .Y(DP_OP_424J2_126_3477_n2269) );
  INVX1_HVT U3859 ( .A(conv_weight_box[38]), .Y(DP_OP_424J2_126_3477_n2275) );
  INVX1_HVT U3860 ( .A(src_window[158]), .Y(DP_OP_424J2_126_3477_n2311) );
  INVX1_HVT U3861 ( .A(src_window[154]), .Y(DP_OP_424J2_126_3477_n2315) );
  INVX1_HVT U3862 ( .A(src_window[152]), .Y(DP_OP_424J2_126_3477_n2317) );
  INVX1_HVT U3863 ( .A(conv_weight_box[44]), .Y(DP_OP_424J2_126_3477_n2318) );
  INVX1_HVT U3864 ( .A(src_window[175]), .Y(DP_OP_424J2_126_3477_n2354) );
  INVX1_HVT U3865 ( .A(src_window[171]), .Y(DP_OP_424J2_126_3477_n2358) );
  INVX1_HVT U3866 ( .A(src_window[189]), .Y(DP_OP_424J2_126_3477_n2400) );
  INVX1_HVT U3867 ( .A(src_window[186]), .Y(DP_OP_424J2_126_3477_n2403) );
  INVX1_HVT U3868 ( .A(src_window[184]), .Y(DP_OP_424J2_126_3477_n2405) );
  INVX1_HVT U3869 ( .A(src_window[214]), .Y(DP_OP_424J2_126_3477_n2443) );
  INVX1_HVT U3870 ( .A(src_window[210]), .Y(DP_OP_424J2_126_3477_n2447) );
  INVX1_HVT U3871 ( .A(src_window[231]), .Y(DP_OP_424J2_126_3477_n2486) );
  INVX1_HVT U3872 ( .A(src_window[226]), .Y(DP_OP_424J2_126_3477_n2491) );
  INVX1_HVT U3873 ( .A(conv_weight_box[62]), .Y(DP_OP_424J2_126_3477_n2497) );
  INVX1_HVT U3874 ( .A(src_window[237]), .Y(DP_OP_424J2_126_3477_n2532) );
  INVX1_HVT U3875 ( .A(src_window[235]), .Y(DP_OP_424J2_126_3477_n2534) );
  INVX1_HVT U3876 ( .A(src_window[234]), .Y(DP_OP_424J2_126_3477_n2535) );
  INVX1_HVT U3877 ( .A(src_window[223]), .Y(DP_OP_424J2_126_3477_n2574) );
  INVX1_HVT U3878 ( .A(src_window[222]), .Y(DP_OP_424J2_126_3477_n2575) );
  INVX1_HVT U3879 ( .A(src_window[221]), .Y(DP_OP_424J2_126_3477_n2576) );
  INVX1_HVT U3880 ( .A(src_window[218]), .Y(DP_OP_424J2_126_3477_n2579) );
  INVX1_HVT U3881 ( .A(src_window[217]), .Y(DP_OP_424J2_126_3477_n2580) );
  INVX1_HVT U3882 ( .A(src_window[206]), .Y(DP_OP_424J2_126_3477_n2619) );
  INVX1_HVT U3883 ( .A(src_window[203]), .Y(DP_OP_424J2_126_3477_n2622) );
  INVX1_HVT U3884 ( .A(src_window[202]), .Y(DP_OP_424J2_126_3477_n2623) );
  INVX1_HVT U3885 ( .A(conv_weight_box[55]), .Y(DP_OP_424J2_126_3477_n2627) );
  INVX1_HVT U3886 ( .A(conv_weight_box[53]), .Y(DP_OP_424J2_126_3477_n2629) );
  INVX1_HVT U3887 ( .A(src_window[178]), .Y(DP_OP_424J2_126_3477_n2667) );
  INVX1_HVT U3888 ( .A(src_window[176]), .Y(DP_OP_424J2_126_3477_n2669) );
  INVX1_HVT U3889 ( .A(conv_weight_box[49]), .Y(DP_OP_424J2_126_3477_n2673) );
  INVX1_HVT U3890 ( .A(src_window[161]), .Y(DP_OP_424J2_126_3477_n2712) );
  INVX1_HVT U3891 ( .A(src_window[141]), .Y(DP_OP_424J2_126_3477_n2752) );
  INVX1_HVT U3892 ( .A(src_window[139]), .Y(DP_OP_424J2_126_3477_n2754) );
  INVX1_HVT U3893 ( .A(src_window[137]), .Y(DP_OP_424J2_126_3477_n2756) );
  INVX1_HVT U3894 ( .A(conv_weight_box[40]), .Y(DP_OP_424J2_126_3477_n2758) );
  INVX1_HVT U3895 ( .A(src_window[127]), .Y(DP_OP_424J2_126_3477_n2794) );
  INVX1_HVT U3896 ( .A(src_window[126]), .Y(DP_OP_424J2_126_3477_n2795) );
  INVX1_HVT U3897 ( .A(src_window[125]), .Y(DP_OP_424J2_126_3477_n2796) );
  INVX1_HVT U3898 ( .A(src_window[122]), .Y(DP_OP_424J2_126_3477_n2799) );
  INVX1_HVT U3899 ( .A(src_window[120]), .Y(DP_OP_424J2_126_3477_n2801) );
  INVX1_HVT U3900 ( .A(conv_weight_box[33]), .Y(DP_OP_424J2_126_3477_n2805) );
  INVX1_HVT U3901 ( .A(src_window[104]), .Y(DP_OP_424J2_126_3477_n2845) );
  INVX1_HVT U3902 ( .A(conv_weight_box[26]), .Y(DP_OP_424J2_126_3477_n2849) );
  INVX1_HVT U3903 ( .A(src_window[87]), .Y(DP_OP_424J2_126_3477_n2882) );
  INVX1_HVT U3904 ( .A(src_window[86]), .Y(DP_OP_424J2_126_3477_n2883) );
  INVX1_HVT U3905 ( .A(src_window[83]), .Y(DP_OP_424J2_126_3477_n2886) );
  INVX1_HVT U3906 ( .A(src_window[82]), .Y(DP_OP_424J2_126_3477_n2887) );
  INVX1_HVT U3907 ( .A(src_window[80]), .Y(DP_OP_424J2_126_3477_n2889) );
  INVX1_HVT U3908 ( .A(conv_weight_box[23]), .Y(DP_OP_424J2_126_3477_n2890) );
  INVX1_HVT U3909 ( .A(conv_weight_box[21]), .Y(DP_OP_424J2_126_3477_n2893) );
  INVX1_HVT U3910 ( .A(src_window[70]), .Y(DP_OP_424J2_126_3477_n2927) );
  INVX1_HVT U3911 ( .A(src_window[69]), .Y(DP_OP_424J2_126_3477_n2928) );
  INVX1_HVT U3912 ( .A(src_window[68]), .Y(DP_OP_424J2_126_3477_n2929) );
  INVX1_HVT U3913 ( .A(src_window[65]), .Y(DP_OP_424J2_126_3477_n2932) );
  INVX1_HVT U3914 ( .A(src_window[64]), .Y(DP_OP_424J2_126_3477_n2933) );
  INVX1_HVT U3915 ( .A(conv_weight_box[16]), .Y(DP_OP_424J2_126_3477_n2936) );
  INVX1_HVT U3916 ( .A(src_window[47]), .Y(DP_OP_424J2_126_3477_n2970) );
  INVX1_HVT U3917 ( .A(src_window[46]), .Y(DP_OP_424J2_126_3477_n2971) );
  INVX1_HVT U3918 ( .A(src_window[45]), .Y(DP_OP_424J2_126_3477_n2972) );
  INVX1_HVT U3919 ( .A(src_window[44]), .Y(DP_OP_424J2_126_3477_n2973) );
  INVX1_HVT U3920 ( .A(src_window[43]), .Y(DP_OP_424J2_126_3477_n2974) );
  INVX1_HVT U3921 ( .A(src_window[42]), .Y(DP_OP_424J2_126_3477_n2975) );
  INVX1_HVT U3922 ( .A(src_window[41]), .Y(DP_OP_424J2_126_3477_n2976) );
  INVX1_HVT U3923 ( .A(src_window[40]), .Y(DP_OP_424J2_126_3477_n2977) );
  INVX1_HVT U3924 ( .A(conv_weight_box[11]), .Y(DP_OP_424J2_126_3477_n2980) );
  INVX1_HVT U3925 ( .A(src_window[30]), .Y(DP_OP_424J2_126_3477_n3015) );
  INVX1_HVT U3926 ( .A(src_window[26]), .Y(DP_OP_424J2_126_3477_n3019) );
  INVX1_HVT U3927 ( .A(src_window[25]), .Y(DP_OP_424J2_126_3477_n3020) );
  INVX1_HVT U3928 ( .A(conv_weight_box[6]), .Y(DP_OP_424J2_126_3477_n3023) );
  INVX1_HVT U3929 ( .A(DP_OP_424J2_126_3477_n302), .Y(
        DP_OP_424J2_126_3477_n303) );
  INVX1_HVT U3930 ( .A(DP_OP_424J2_126_3477_n304), .Y(
        DP_OP_424J2_126_3477_n305) );
  INVX1_HVT U3931 ( .A(src_window[14]), .Y(DP_OP_424J2_126_3477_n3057) );
  INVX1_HVT U3932 ( .A(src_window[13]), .Y(DP_OP_424J2_126_3477_n3058) );
  INVX1_HVT U3933 ( .A(src_window[12]), .Y(DP_OP_424J2_126_3477_n3059) );
  INVX1_HVT U3934 ( .A(src_window[11]), .Y(DP_OP_424J2_126_3477_n3060) );
  INVX1_HVT U3935 ( .A(src_window[8]), .Y(DP_OP_424J2_126_3477_n3063) );
  INVX1_HVT U3936 ( .A(conv_weight_box[1]), .Y(DP_OP_424J2_126_3477_n3065) );
  INVX1_HVT U3937 ( .A(conv_weight_box[0]), .Y(DP_OP_424J2_126_3477_n3066) );
  INVX1_HVT U3938 ( .A(DP_OP_424J2_126_3477_n306), .Y(
        DP_OP_424J2_126_3477_n307) );
  INVX1_HVT U3939 ( .A(DP_OP_424J2_126_3477_n308), .Y(
        DP_OP_424J2_126_3477_n309) );
  INVX1_HVT U3940 ( .A(DP_OP_424J2_126_3477_n310), .Y(
        DP_OP_424J2_126_3477_n311) );
  INVX1_HVT U3941 ( .A(DP_OP_424J2_126_3477_n312), .Y(
        DP_OP_424J2_126_3477_n313) );
  INVX1_HVT U3942 ( .A(DP_OP_424J2_126_3477_n314), .Y(
        DP_OP_424J2_126_3477_n315) );
  INVX1_HVT U3943 ( .A(DP_OP_424J2_126_3477_n316), .Y(
        DP_OP_424J2_126_3477_n317) );
  INVX1_HVT U3944 ( .A(DP_OP_424J2_126_3477_n318), .Y(
        DP_OP_424J2_126_3477_n319) );
  INVX1_HVT U3945 ( .A(DP_OP_424J2_126_3477_n322), .Y(
        DP_OP_424J2_126_3477_n323) );
  INVX1_HVT U3946 ( .A(DP_OP_424J2_126_3477_n324), .Y(
        DP_OP_424J2_126_3477_n325) );
  INVX1_HVT U3947 ( .A(DP_OP_424J2_126_3477_n326), .Y(
        DP_OP_424J2_126_3477_n327) );
  INVX1_HVT U3948 ( .A(DP_OP_424J2_126_3477_n328), .Y(
        DP_OP_424J2_126_3477_n329) );
  INVX1_HVT U3949 ( .A(DP_OP_424J2_126_3477_n330), .Y(
        DP_OP_424J2_126_3477_n331) );
  INVX1_HVT U3950 ( .A(DP_OP_424J2_126_3477_n71), .Y(DP_OP_424J2_126_3477_n69)
         );
  INVX1_HVT U3951 ( .A(DP_OP_424J2_126_3477_n820), .Y(
        DP_OP_424J2_126_3477_n821) );
  INVX1_HVT U3952 ( .A(DP_OP_424J2_126_3477_n95), .Y(DP_OP_424J2_126_3477_n93)
         );
  NAND2X0_HVT U3953 ( .A1(DP_OP_424J2_126_3477_n649), .A2(
        DP_OP_424J2_126_3477_n822), .Y(DP_OP_424J2_126_3477_n240) );
  NAND2X0_HVT U3954 ( .A1(n1716), .A2(n1720), .Y(n1719) );
  OR2X1_HVT U3955 ( .A1(DP_OP_424J2_126_3477_n424), .A2(
        DP_OP_424J2_126_3477_n379), .Y(n1721) );
  AO22X1_HVT U3956 ( .A1(DP_OP_424J2_126_3477_n379), .A2(
        DP_OP_424J2_126_3477_n424), .A3(DP_OP_424J2_126_3477_n422), .A4(n1721), 
        .Y(DP_OP_424J2_126_3477_n374) );
  NAND2X0_HVT U3957 ( .A1(n182), .A2(n1726), .Y(n1727) );
  OR2X1_HVT U3958 ( .A1(DP_OP_424J2_126_3477_n22), .A2(n1723), .Y(n1728) );
  NAND2X0_HVT U3959 ( .A1(DP_OP_424J2_126_3477_n202), .A2(n1724), .Y(n1729) );
  NAND2X0_HVT U3960 ( .A1(n1729), .A2(n1723), .Y(n1730) );
  NAND2X0_HVT U3961 ( .A1(n1728), .A2(n1730), .Y(n1731) );
  NAND3X0_HVT U3962 ( .A1(n1725), .A2(n1727), .A3(n1731), .Y(n_conv2_sum_c[15]) );
  OR2X1_HVT U3963 ( .A1(DP_OP_424J2_126_3477_n822), .A2(
        DP_OP_424J2_126_3477_n649), .Y(n1714) );
  OR2X1_HVT U3964 ( .A1(DP_OP_424J2_126_3477_n1021), .A2(
        DP_OP_424J2_126_3477_n1019), .Y(DP_OP_424J2_126_3477_n295) );
  OR2X1_HVT U3965 ( .A1(DP_OP_424J2_126_3477_n1215), .A2(
        DP_OP_424J2_126_3477_n1213), .Y(n1735) );
  OR2X1_HVT U3966 ( .A1(DP_OP_424J2_126_3477_n1403), .A2(
        DP_OP_424J2_126_3477_n1401), .Y(DP_OP_424J2_126_3477_n297) );
  AO21X1_HVT U3967 ( .A1(n1735), .A2(n1737), .A3(n1738), .Y(
        DP_OP_424J2_126_3477_n250) );
  FADDX1_HVT U3968 ( .A(DP_OP_424J2_126_3477_n1455), .B(
        DP_OP_424J2_126_3477_n1449), .CI(DP_OP_424J2_126_3477_n1453), .CO(
        DP_OP_424J2_126_3477_n1424) );
  NAND2X0_HVT U3969 ( .A1(n1712), .A2(n1711), .Y(n1746) );
  NAND2X0_HVT U3970 ( .A1(n1746), .A2(DP_OP_424J2_126_3477_n226), .Y(
        DP_OP_424J2_126_3477_n220) );
  AND2X1_HVT U3971 ( .A1(n1732), .A2(n1711), .Y(DP_OP_424J2_126_3477_n219) );
  NAND2X0_HVT U3972 ( .A1(DP_OP_424J2_126_3477_n201), .A2(
        DP_OP_424J2_126_3477_n286), .Y(n1747) );
  AND2X1_HVT U3973 ( .A1(n1747), .A2(DP_OP_424J2_126_3477_n198), .Y(
        DP_OP_424J2_126_3477_n190) );
  OR2X1_HVT U3974 ( .A1(DP_OP_424J2_126_3477_n13), .A2(
        DP_OP_424J2_126_3477_n110), .Y(n1751) );
  NAND2X0_HVT U3975 ( .A1(n1768), .A2(n1753), .Y(n1754) );
  OA22X1_HVT U3976 ( .A1(n1768), .A2(n1753), .A3(n1754), .A4(
        DP_OP_424J2_126_3477_n151), .Y(n1755) );
  OR2X1_HVT U3977 ( .A1(DP_OP_424J2_126_3477_n302), .A2(n1757), .Y(n1756) );
  OR2X1_HVT U3978 ( .A1(DP_OP_424J2_126_3477_n304), .A2(
        DP_OP_424J2_126_3477_n303), .Y(n1758) );
  OR2X1_HVT U3979 ( .A1(DP_OP_424J2_126_3477_n308), .A2(
        DP_OP_424J2_126_3477_n307), .Y(n1759) );
  OR2X1_HVT U3980 ( .A1(DP_OP_424J2_126_3477_n171), .A2(
        DP_OP_424J2_126_3477_n178), .Y(n1760) );
  INVX1_HVT U3981 ( .A(DP_OP_424J2_126_3477_n209), .Y(n1752) );
  OR2X1_HVT U3982 ( .A1(DP_OP_424J2_126_3477_n1733), .A2(
        DP_OP_424J2_126_3477_n1731), .Y(n1762) );
  OR2X1_HVT U3983 ( .A1(DP_OP_424J2_126_3477_n312), .A2(
        DP_OP_424J2_126_3477_n311), .Y(n1763) );
  OR2X1_HVT U3984 ( .A1(DP_OP_424J2_126_3477_n318), .A2(
        DP_OP_424J2_126_3477_n317), .Y(n1764) );
  AND2X1_HVT U3985 ( .A1(DP_OP_424J2_126_3477_n151), .A2(
        DP_OP_424J2_126_3477_n17), .Y(n1765) );
  AND2X1_HVT U3986 ( .A1(DP_OP_424J2_126_3477_n107), .A2(
        DP_OP_424J2_126_3477_n13), .Y(n1766) );
  OA21X1_HVT U3987 ( .A1(DP_OP_424J2_126_3477_n153), .A2(n1748), .A3(
        DP_OP_424J2_126_3477_n156), .Y(n1768) );
  INVX1_HVT U3988 ( .A(DP_OP_424J2_126_3477_n2922), .Y(n1717) );
  OA21X1_HVT U3989 ( .A1(DP_OP_424J2_126_3477_n171), .A2(n1740), .A3(
        DP_OP_424J2_126_3477_n174), .Y(n1767) );
  INVX1_HVT U3990 ( .A(DP_OP_424J2_126_3477_n114), .Y(n1743) );
  OA21X1_HVT U3991 ( .A1(DP_OP_424J2_126_3477_n144), .A2(n1740), .A3(
        DP_OP_424J2_126_3477_n145), .Y(DP_OP_424J2_126_3477_n141) );
  INVX1_HVT U3992 ( .A(conv_weight_box[66]), .Y(DP_OP_424J2_126_3477_n2541) );
  INVX1_HVT U3993 ( .A(conv_weight_box[60]), .Y(DP_OP_424J2_126_3477_n2585) );
  INVX1_HVT U3994 ( .A(conv_weight_box[8]), .Y(DP_OP_424J2_126_3477_n2057) );
  INVX1_HVT U3995 ( .A(conv_weight_box[51]), .Y(DP_OP_424J2_126_3477_n2409) );
  OR2X1_HVT U3996 ( .A1(DP_OP_424J2_126_3477_n372), .A2(
        DP_OP_424J2_126_3477_n351), .Y(n1745) );
  INVX1_HVT U3997 ( .A(n1518), .Y(n1722) );
  INVX1_HVT U3998 ( .A(DP_OP_424J2_126_3477_n338), .Y(
        DP_OP_424J2_126_3477_n339) );
  INVX1_HVT U3999 ( .A(DP_OP_425J2_127_3477_n1728), .Y(
        DP_OP_425J2_127_3477_n1729) );
  INVX1_HVT U4000 ( .A(DP_OP_425J2_127_3477_n197), .Y(
        DP_OP_425J2_127_3477_n286) );
  INVX1_HVT U4001 ( .A(src_window[15]), .Y(DP_OP_425J2_127_3477_n2002) );
  INVX1_HVT U4002 ( .A(src_window[10]), .Y(DP_OP_425J2_127_3477_n2007) );
  INVX1_HVT U4003 ( .A(src_window[9]), .Y(DP_OP_425J2_127_3477_n2008) );
  INVX1_HVT U4004 ( .A(DP_OP_425J2_127_3477_n203), .Y(
        DP_OP_425J2_127_3477_n201) );
  INVX1_HVT U4005 ( .A(conv_weight_box[3]), .Y(DP_OP_425J2_127_3477_n2011) );
  INVX1_HVT U4006 ( .A(src_window[31]), .Y(DP_OP_425J2_127_3477_n2046) );
  INVX1_HVT U4007 ( .A(src_window[29]), .Y(DP_OP_425J2_127_3477_n2048) );
  INVX1_HVT U4008 ( .A(src_window[28]), .Y(DP_OP_425J2_127_3477_n2049) );
  INVX1_HVT U4009 ( .A(src_window[27]), .Y(DP_OP_425J2_127_3477_n2050) );
  INVX1_HVT U4010 ( .A(src_window[24]), .Y(DP_OP_425J2_127_3477_n2053) );
  INVX1_HVT U4011 ( .A(conv_weight_box[10]), .Y(DP_OP_425J2_127_3477_n2055) );
  INVX1_HVT U4012 ( .A(src_window[53]), .Y(DP_OP_425J2_127_3477_n2092) );
  INVX1_HVT U4013 ( .A(conv_weight_box[15]), .Y(DP_OP_425J2_127_3477_n2098) );
  INVX1_HVT U4014 ( .A(conv_weight_box[14]), .Y(DP_OP_425J2_127_3477_n2099) );
  INVX1_HVT U4015 ( .A(src_window[67]), .Y(DP_OP_425J2_127_3477_n2138) );
  INVX1_HVT U4016 ( .A(conv_weight_box[19]), .Y(DP_OP_425J2_127_3477_n2144) );
  INVX1_HVT U4017 ( .A(src_window[85]), .Y(DP_OP_425J2_127_3477_n2180) );
  INVX1_HVT U4018 ( .A(src_window[83]), .Y(DP_OP_425J2_127_3477_n2182) );
  INVX1_HVT U4019 ( .A(src_window[81]), .Y(DP_OP_425J2_127_3477_n2184) );
  INVX1_HVT U4020 ( .A(src_window[80]), .Y(DP_OP_425J2_127_3477_n2185) );
  INVX1_HVT U4021 ( .A(conv_weight_box[25]), .Y(DP_OP_425J2_127_3477_n2186) );
  INVX1_HVT U4022 ( .A(conv_weight_box[24]), .Y(DP_OP_425J2_127_3477_n2189) );
  INVX1_HVT U4023 ( .A(src_window[107]), .Y(DP_OP_425J2_127_3477_n2226) );
  INVX1_HVT U4024 ( .A(conv_weight_box[32]), .Y(DP_OP_425J2_127_3477_n2230) );
  INVX1_HVT U4025 ( .A(src_window[125]), .Y(DP_OP_425J2_127_3477_n2268) );
  INVX1_HVT U4026 ( .A(src_window[124]), .Y(DP_OP_425J2_127_3477_n2269) );
  INVX1_HVT U4027 ( .A(src_window[121]), .Y(DP_OP_425J2_127_3477_n2272) );
  INVX1_HVT U4028 ( .A(src_window[151]), .Y(DP_OP_425J2_127_3477_n2310) );
  INVX1_HVT U4029 ( .A(src_window[150]), .Y(DP_OP_425J2_127_3477_n2311) );
  INVX1_HVT U4030 ( .A(src_window[149]), .Y(DP_OP_425J2_127_3477_n2312) );
  INVX1_HVT U4031 ( .A(conv_weight_box[42]), .Y(DP_OP_425J2_127_3477_n2320) );
  INVX1_HVT U4032 ( .A(conv_weight_box[41]), .Y(DP_OP_425J2_127_3477_n2321) );
  INVX1_HVT U4033 ( .A(src_window[165]), .Y(DP_OP_425J2_127_3477_n2356) );
  INVX1_HVT U4034 ( .A(src_window[164]), .Y(DP_OP_425J2_127_3477_n2357) );
  INVX1_HVT U4035 ( .A(src_window[163]), .Y(DP_OP_425J2_127_3477_n2358) );
  INVX1_HVT U4036 ( .A(src_window[162]), .Y(DP_OP_425J2_127_3477_n2359) );
  INVX1_HVT U4037 ( .A(src_window[181]), .Y(DP_OP_425J2_127_3477_n2400) );
  INVX1_HVT U4038 ( .A(src_window[180]), .Y(DP_OP_425J2_127_3477_n2401) );
  INVX1_HVT U4039 ( .A(src_window[178]), .Y(DP_OP_425J2_127_3477_n2403) );
  INVX1_HVT U4040 ( .A(src_window[177]), .Y(DP_OP_425J2_127_3477_n2404) );
  INVX1_HVT U4041 ( .A(src_window[204]), .Y(DP_OP_425J2_127_3477_n2445) );
  INVX1_HVT U4042 ( .A(src_window[202]), .Y(DP_OP_425J2_127_3477_n2447) );
  INVX1_HVT U4043 ( .A(src_window[201]), .Y(DP_OP_425J2_127_3477_n2448) );
  INVX1_HVT U4044 ( .A(src_window[200]), .Y(DP_OP_425J2_127_3477_n2449) );
  INVX1_HVT U4045 ( .A(src_window[216]), .Y(DP_OP_425J2_127_3477_n2493) );
  INVX1_HVT U4046 ( .A(conv_weight_box[62]), .Y(DP_OP_425J2_127_3477_n2497) );
  INVX1_HVT U4047 ( .A(src_window[227]), .Y(DP_OP_425J2_127_3477_n2534) );
  INVX1_HVT U4048 ( .A(src_window[225]), .Y(DP_OP_425J2_127_3477_n2536) );
  INVX1_HVT U4049 ( .A(src_window[215]), .Y(DP_OP_425J2_127_3477_n2574) );
  INVX1_HVT U4050 ( .A(src_window[213]), .Y(DP_OP_425J2_127_3477_n2576) );
  INVX1_HVT U4051 ( .A(src_window[212]), .Y(DP_OP_425J2_127_3477_n2577) );
  INVX1_HVT U4052 ( .A(src_window[211]), .Y(DP_OP_425J2_127_3477_n2578) );
  INVX1_HVT U4053 ( .A(src_window[210]), .Y(DP_OP_425J2_127_3477_n2579) );
  INVX1_HVT U4054 ( .A(src_window[209]), .Y(DP_OP_425J2_127_3477_n2580) );
  INVX1_HVT U4055 ( .A(src_window[208]), .Y(DP_OP_425J2_127_3477_n2581) );
  INVX1_HVT U4056 ( .A(conv_weight_box[61]), .Y(DP_OP_425J2_127_3477_n2582) );
  INVX1_HVT U4057 ( .A(src_window[197]), .Y(DP_OP_425J2_127_3477_n2620) );
  INVX1_HVT U4058 ( .A(src_window[196]), .Y(DP_OP_425J2_127_3477_n2621) );
  INVX1_HVT U4059 ( .A(src_window[195]), .Y(DP_OP_425J2_127_3477_n2622) );
  INVX1_HVT U4060 ( .A(conv_weight_box[49]), .Y(DP_OP_425J2_127_3477_n2673) );
  INVX1_HVT U4061 ( .A(src_window[157]), .Y(DP_OP_425J2_127_3477_n2708) );
  INVX1_HVT U4062 ( .A(src_window[155]), .Y(DP_OP_425J2_127_3477_n2710) );
  INVX1_HVT U4063 ( .A(src_window[153]), .Y(DP_OP_425J2_127_3477_n2712) );
  INVX1_HVT U4064 ( .A(src_window[131]), .Y(DP_OP_425J2_127_3477_n2754) );
  INVX1_HVT U4065 ( .A(src_window[130]), .Y(DP_OP_425J2_127_3477_n2755) );
  INVX1_HVT U4066 ( .A(src_window[129]), .Y(DP_OP_425J2_127_3477_n2756) );
  INVX1_HVT U4067 ( .A(conv_weight_box[39]), .Y(DP_OP_425J2_127_3477_n2760) );
  INVX1_HVT U4068 ( .A(src_window[117]), .Y(DP_OP_425J2_127_3477_n2796) );
  INVX1_HVT U4069 ( .A(src_window[116]), .Y(DP_OP_425J2_127_3477_n2797) );
  INVX1_HVT U4070 ( .A(src_window[115]), .Y(DP_OP_425J2_127_3477_n2798) );
  INVX1_HVT U4071 ( .A(src_window[114]), .Y(DP_OP_425J2_127_3477_n2799) );
  INVX1_HVT U4072 ( .A(src_window[113]), .Y(DP_OP_425J2_127_3477_n2800) );
  INVX1_HVT U4073 ( .A(src_window[112]), .Y(DP_OP_425J2_127_3477_n2801) );
  INVX1_HVT U4074 ( .A(src_window[102]), .Y(DP_OP_425J2_127_3477_n2839) );
  INVX1_HVT U4075 ( .A(src_window[101]), .Y(DP_OP_425J2_127_3477_n2840) );
  INVX1_HVT U4076 ( .A(src_window[100]), .Y(DP_OP_425J2_127_3477_n2841) );
  INVX1_HVT U4077 ( .A(src_window[98]), .Y(DP_OP_425J2_127_3477_n2843) );
  INVX1_HVT U4078 ( .A(conv_weight_box[28]), .Y(DP_OP_425J2_127_3477_n2847) );
  INVX1_HVT U4079 ( .A(src_window[79]), .Y(DP_OP_425J2_127_3477_n2882) );
  INVX1_HVT U4080 ( .A(src_window[78]), .Y(DP_OP_425J2_127_3477_n2883) );
  INVX1_HVT U4081 ( .A(src_window[76]), .Y(DP_OP_425J2_127_3477_n2885) );
  INVX1_HVT U4082 ( .A(src_window[75]), .Y(DP_OP_425J2_127_3477_n2886) );
  INVX1_HVT U4083 ( .A(src_window[73]), .Y(DP_OP_425J2_127_3477_n2888) );
  INVX1_HVT U4084 ( .A(conv_weight_box[21]), .Y(DP_OP_425J2_127_3477_n2893) );
  INVX1_HVT U4085 ( .A(src_window[56]), .Y(DP_OP_425J2_127_3477_n2933) );
  INVX1_HVT U4086 ( .A(src_window[39]), .Y(DP_OP_425J2_127_3477_n2970) );
  INVX1_HVT U4087 ( .A(src_window[38]), .Y(DP_OP_425J2_127_3477_n2971) );
  INVX1_HVT U4088 ( .A(src_window[37]), .Y(DP_OP_425J2_127_3477_n2972) );
  INVX1_HVT U4089 ( .A(src_window[36]), .Y(DP_OP_425J2_127_3477_n2973) );
  INVX1_HVT U4090 ( .A(src_window[35]), .Y(DP_OP_425J2_127_3477_n2974) );
  INVX1_HVT U4091 ( .A(src_window[33]), .Y(DP_OP_425J2_127_3477_n2976) );
  INVX1_HVT U4092 ( .A(src_window[32]), .Y(DP_OP_425J2_127_3477_n2977) );
  INVX1_HVT U4093 ( .A(conv_weight_box[11]), .Y(DP_OP_425J2_127_3477_n2980) );
  INVX1_HVT U4094 ( .A(src_window[18]), .Y(DP_OP_425J2_127_3477_n3019) );
  INVX1_HVT U4095 ( .A(src_window[17]), .Y(DP_OP_425J2_127_3477_n3020) );
  INVX1_HVT U4096 ( .A(src_window[16]), .Y(DP_OP_425J2_127_3477_n3021) );
  INVX1_HVT U4097 ( .A(conv_weight_box[6]), .Y(DP_OP_425J2_127_3477_n3023) );
  INVX1_HVT U4098 ( .A(DP_OP_425J2_127_3477_n302), .Y(
        DP_OP_425J2_127_3477_n303) );
  INVX1_HVT U4099 ( .A(DP_OP_425J2_127_3477_n304), .Y(
        DP_OP_425J2_127_3477_n305) );
  INVX1_HVT U4100 ( .A(src_window[7]), .Y(DP_OP_425J2_127_3477_n3056) );
  INVX1_HVT U4101 ( .A(src_window[6]), .Y(DP_OP_425J2_127_3477_n3057) );
  INVX1_HVT U4102 ( .A(src_window[5]), .Y(DP_OP_425J2_127_3477_n3058) );
  INVX1_HVT U4103 ( .A(src_window[4]), .Y(DP_OP_425J2_127_3477_n3059) );
  INVX1_HVT U4104 ( .A(src_window[3]), .Y(DP_OP_425J2_127_3477_n3060) );
  INVX1_HVT U4105 ( .A(src_window[2]), .Y(DP_OP_425J2_127_3477_n3061) );
  INVX1_HVT U4106 ( .A(src_window[1]), .Y(DP_OP_425J2_127_3477_n3062) );
  INVX1_HVT U4107 ( .A(src_window[0]), .Y(DP_OP_425J2_127_3477_n3063) );
  INVX1_HVT U4108 ( .A(conv_weight_box[1]), .Y(DP_OP_425J2_127_3477_n3065) );
  INVX1_HVT U4109 ( .A(conv_weight_box[0]), .Y(DP_OP_425J2_127_3477_n3066) );
  INVX1_HVT U4110 ( .A(DP_OP_425J2_127_3477_n306), .Y(
        DP_OP_425J2_127_3477_n307) );
  INVX1_HVT U4111 ( .A(DP_OP_425J2_127_3477_n308), .Y(
        DP_OP_425J2_127_3477_n309) );
  INVX1_HVT U4112 ( .A(DP_OP_425J2_127_3477_n310), .Y(
        DP_OP_425J2_127_3477_n311) );
  INVX1_HVT U4113 ( .A(DP_OP_425J2_127_3477_n312), .Y(
        DP_OP_425J2_127_3477_n313) );
  INVX1_HVT U4114 ( .A(DP_OP_425J2_127_3477_n314), .Y(
        DP_OP_425J2_127_3477_n315) );
  INVX1_HVT U4115 ( .A(DP_OP_425J2_127_3477_n316), .Y(
        DP_OP_425J2_127_3477_n317) );
  INVX1_HVT U4116 ( .A(DP_OP_425J2_127_3477_n318), .Y(
        DP_OP_425J2_127_3477_n319) );
  INVX1_HVT U4117 ( .A(DP_OP_425J2_127_3477_n320), .Y(
        DP_OP_425J2_127_3477_n321) );
  INVX1_HVT U4118 ( .A(DP_OP_425J2_127_3477_n322), .Y(
        DP_OP_425J2_127_3477_n323) );
  INVX1_HVT U4119 ( .A(DP_OP_425J2_127_3477_n324), .Y(
        DP_OP_425J2_127_3477_n325) );
  INVX1_HVT U4120 ( .A(DP_OP_425J2_127_3477_n326), .Y(
        DP_OP_425J2_127_3477_n327) );
  INVX1_HVT U4121 ( .A(DP_OP_425J2_127_3477_n328), .Y(
        DP_OP_425J2_127_3477_n329) );
  INVX1_HVT U4122 ( .A(DP_OP_425J2_127_3477_n510), .Y(
        DP_OP_425J2_127_3477_n511) );
  INVX1_HVT U4123 ( .A(DP_OP_425J2_127_3477_n71), .Y(DP_OP_425J2_127_3477_n69)
         );
  INVX1_HVT U4124 ( .A(DP_OP_425J2_127_3477_n820), .Y(
        DP_OP_425J2_127_3477_n821) );
  INVX1_HVT U4125 ( .A(DP_OP_425J2_127_3477_n95), .Y(DP_OP_425J2_127_3477_n93)
         );
  NAND2X0_HVT U4126 ( .A1(DP_OP_425J2_127_3477_n649), .A2(
        DP_OP_425J2_127_3477_n822), .Y(DP_OP_425J2_127_3477_n240) );
  NAND2X0_HVT U4127 ( .A1(n1775), .A2(n1779), .Y(n1778) );
  OR2X1_HVT U4128 ( .A1(DP_OP_425J2_127_3477_n424), .A2(
        DP_OP_425J2_127_3477_n379), .Y(n1780) );
  AO22X1_HVT U4129 ( .A1(DP_OP_425J2_127_3477_n379), .A2(
        DP_OP_425J2_127_3477_n424), .A3(DP_OP_425J2_127_3477_n422), .A4(n1780), 
        .Y(DP_OP_425J2_127_3477_n374) );
  NAND2X0_HVT U4130 ( .A1(n1823), .A2(n1785), .Y(n1786) );
  OR2X1_HVT U4131 ( .A1(DP_OP_425J2_127_3477_n22), .A2(n1782), .Y(n1787) );
  NAND2X0_HVT U4132 ( .A1(DP_OP_425J2_127_3477_n202), .A2(n1783), .Y(n1788) );
  NAND2X0_HVT U4133 ( .A1(n1788), .A2(n1782), .Y(n1789) );
  NAND2X0_HVT U4134 ( .A1(n1787), .A2(n1789), .Y(n1790) );
  NAND3X0_HVT U4135 ( .A1(n1784), .A2(n1786), .A3(n1790), .Y(n_conv2_sum_d[15]) );
  OR2X1_HVT U4136 ( .A1(DP_OP_425J2_127_3477_n1021), .A2(
        DP_OP_425J2_127_3477_n1019), .Y(DP_OP_425J2_127_3477_n295) );
  OR2X1_HVT U4137 ( .A1(DP_OP_425J2_127_3477_n1215), .A2(
        DP_OP_425J2_127_3477_n1213), .Y(n1795) );
  OR2X1_HVT U4138 ( .A1(DP_OP_425J2_127_3477_n1403), .A2(
        DP_OP_425J2_127_3477_n1401), .Y(DP_OP_425J2_127_3477_n297) );
  AO21X1_HVT U4139 ( .A1(DP_OP_425J2_127_3477_n297), .A2(n1796), .A3(
        DP_OP_425J2_127_3477_n255), .Y(n1797) );
  AO21X1_HVT U4140 ( .A1(n1795), .A2(n1797), .A3(n1798), .Y(
        DP_OP_425J2_127_3477_n250) );
  FADDX1_HVT U4141 ( .A(DP_OP_425J2_127_3477_n1453), .B(
        DP_OP_425J2_127_3477_n1449), .CI(DP_OP_425J2_127_3477_n1455), .CO(
        DP_OP_425J2_127_3477_n1424) );
  NAND2X0_HVT U4142 ( .A1(n1832), .A2(DP_OP_425J2_127_3477_n67), .Y(n1799) );
  NAND2X0_HVT U4143 ( .A1(n1832), .A2(DP_OP_425J2_127_3477_n187), .Y(n1800) );
  NAND2X0_HVT U4144 ( .A1(n1832), .A2(DP_OP_425J2_127_3477_n54), .Y(n1801) );
  NAND2X0_HVT U4145 ( .A1(n1832), .A2(DP_OP_425J2_127_3477_n49), .Y(n1802) );
  NAND2X0_HVT U4146 ( .A1(n1832), .A2(DP_OP_425J2_127_3477_n176), .Y(n1804) );
  NAND2X0_HVT U4147 ( .A1(n1832), .A2(DP_OP_425J2_127_3477_n122), .Y(n1805) );
  NAND2X0_HVT U4148 ( .A1(n1832), .A2(DP_OP_425J2_127_3477_n91), .Y(n1810) );
  NAND2X0_HVT U4149 ( .A1(n1771), .A2(n1770), .Y(n1815) );
  NAND2X0_HVT U4150 ( .A1(n1815), .A2(DP_OP_425J2_127_3477_n226), .Y(
        DP_OP_425J2_127_3477_n220) );
  NAND2X0_HVT U4151 ( .A1(DP_OP_425J2_127_3477_n207), .A2(n1817), .Y(n1818) );
  OA21X1_HVT U4152 ( .A1(DP_OP_425J2_127_3477_n240), .A2(
        DP_OP_425J2_127_3477_n236), .A3(DP_OP_425J2_127_3477_n237), .Y(n1774)
         );
  NAND2X0_HVT U4153 ( .A1(n1792), .A2(n1774), .Y(n1819) );
  AND3X1_HVT U4154 ( .A1(n1791), .A2(n1770), .A3(DP_OP_425J2_127_3477_n207), 
        .Y(n1820) );
  AND2X1_HVT U4155 ( .A1(n1791), .A2(n1770), .Y(DP_OP_425J2_127_3477_n219) );
  NAND2X0_HVT U4156 ( .A1(DP_OP_425J2_127_3477_n201), .A2(
        DP_OP_425J2_127_3477_n286), .Y(n1821) );
  OA21X1_HVT U4157 ( .A1(DP_OP_425J2_127_3477_n182), .A2(
        DP_OP_425J2_127_3477_n190), .A3(DP_OP_425J2_127_3477_n185), .Y(n1806)
         );
  AND2X1_HVT U4158 ( .A1(n1821), .A2(DP_OP_425J2_127_3477_n198), .Y(
        DP_OP_425J2_127_3477_n190) );
  OR2X1_HVT U4159 ( .A1(DP_OP_425J2_127_3477_n13), .A2(
        DP_OP_425J2_127_3477_n110), .Y(n1826) );
  AND2X1_HVT U4160 ( .A1(n1814), .A2(n1827), .Y(DP_OP_425J2_127_3477_n207) );
  AND2X1_HVT U4161 ( .A1(DP_OP_425J2_127_3477_n419), .A2(
        DP_OP_425J2_127_3477_n512), .Y(n1771) );
  NAND3X0_HVT U4162 ( .A1(DP_OP_425J2_127_3477_n207), .A2(n1771), .A3(n1770), 
        .Y(n1816) );
  NAND2X0_HVT U4163 ( .A1(n1846), .A2(n1828), .Y(n1829) );
  OA22X1_HVT U4164 ( .A1(n1846), .A2(n1828), .A3(n1829), .A4(
        DP_OP_425J2_127_3477_n151), .Y(n1830) );
  AO21X1_HVT U4165 ( .A1(DP_OP_425J2_127_3477_n131), .A2(n1832), .A3(
        DP_OP_425J2_127_3477_n132), .Y(n1831) );
  OR2X1_HVT U4166 ( .A1(DP_OP_425J2_127_3477_n302), .A2(n1834), .Y(n1833) );
  OR2X1_HVT U4167 ( .A1(DP_OP_425J2_127_3477_n304), .A2(
        DP_OP_425J2_127_3477_n303), .Y(n1835) );
  OR2X1_HVT U4168 ( .A1(DP_OP_425J2_127_3477_n308), .A2(
        DP_OP_425J2_127_3477_n307), .Y(n1836) );
  OR2X1_HVT U4169 ( .A1(DP_OP_425J2_127_3477_n171), .A2(
        DP_OP_425J2_127_3477_n178), .Y(n1837) );
  INVX1_HVT U4170 ( .A(DP_OP_425J2_127_3477_n209), .Y(n1827) );
  OR2X1_HVT U4171 ( .A1(DP_OP_425J2_127_3477_n1733), .A2(
        DP_OP_425J2_127_3477_n1731), .Y(n1840) );
  OR2X1_HVT U4172 ( .A1(DP_OP_425J2_127_3477_n312), .A2(
        DP_OP_425J2_127_3477_n311), .Y(n1841) );
  OR2X1_HVT U4173 ( .A1(DP_OP_425J2_127_3477_n318), .A2(
        DP_OP_425J2_127_3477_n317), .Y(n1842) );
  AND2X1_HVT U4174 ( .A1(DP_OP_425J2_127_3477_n151), .A2(
        DP_OP_425J2_127_3477_n17), .Y(n1843) );
  AND2X1_HVT U4175 ( .A1(DP_OP_425J2_127_3477_n107), .A2(
        DP_OP_425J2_127_3477_n13), .Y(n1844) );
  OA21X1_HVT U4176 ( .A1(DP_OP_425J2_127_3477_n153), .A2(n1822), .A3(
        DP_OP_425J2_127_3477_n156), .Y(n1846) );
  INVX1_HVT U4177 ( .A(conv2_sum_d[1]), .Y(DP_OP_425J2_127_3477_n1968) );
  INVX1_HVT U4178 ( .A(DP_OP_425J2_127_3477_n2922), .Y(n1776) );
  OA21X1_HVT U4179 ( .A1(DP_OP_425J2_127_3477_n209), .A2(
        DP_OP_425J2_127_3477_n217), .A3(DP_OP_425J2_127_3477_n210), .Y(n1839)
         );
  OA21X1_HVT U4180 ( .A1(DP_OP_425J2_127_3477_n171), .A2(n1806), .A3(
        DP_OP_425J2_127_3477_n174), .Y(n1845) );
  INVX1_HVT U4181 ( .A(DP_OP_425J2_127_3477_n114), .Y(n1812) );
  OA21X1_HVT U4182 ( .A1(DP_OP_425J2_127_3477_n144), .A2(n1806), .A3(
        DP_OP_425J2_127_3477_n145), .Y(DP_OP_425J2_127_3477_n141) );
  INVX1_HVT U4183 ( .A(conv_weight_box[51]), .Y(DP_OP_425J2_127_3477_n2409) );
  INVX1_HVT U4184 ( .A(conv_weight_box[66]), .Y(DP_OP_425J2_127_3477_n2541) );
  INVX1_HVT U4185 ( .A(conv_weight_box[5]), .Y(DP_OP_425J2_127_3477_n3025) );
  INVX1_HVT U4186 ( .A(DP_OP_425J2_127_3477_n338), .Y(
        DP_OP_425J2_127_3477_n339) );
  INVX1_HVT U4187 ( .A(conv_weight_box[4]), .Y(DP_OP_425J2_127_3477_n2010) );
  OR2X1_HVT U4188 ( .A1(DP_OP_425J2_127_3477_n648), .A2(
        DP_OP_425J2_127_3477_n513), .Y(n1772) );
  MUX21X2_HVT U4189 ( .A1(conv2_sram_rdata_weight[26]), .A2(
        conv1_sram_rdata_weight[26]), .S0(n345), .Y(conv_weight_box[17]) );
  NAND2X4_HVT U4190 ( .A1(n2149), .A2(n2150), .Y(N9) );
  MUX21X1_HVT U4191 ( .A1(conv2_sram_rdata_weight[2]), .A2(
        conv1_sram_rdata_weight[2]), .S0(n92), .Y(conv_weight_box[1]) );
  MUX21X1_HVT U4192 ( .A1(conv2_sram_rdata_weight[82]), .A2(
        conv1_sram_rdata_weight[82]), .S0(n619), .Y(conv_weight_box[55]) );
  MUX21X1_HVT U4193 ( .A1(tmp_big2[9]), .A2(tmp_big1[9]), .S0(N9), .Y(
        data_out[9]) );
  MUX21X1_HVT U4194 ( .A1(tmp_big2[10]), .A2(tmp_big1[10]), .S0(N9), .Y(
        data_out[10]) );
  MUX21X1_HVT U4195 ( .A1(conv2_sram_rdata_weight[6]), .A2(
        conv1_sram_rdata_weight[6]), .S0(n92), .Y(conv_weight_box[3]) );
  MUX21X1_HVT U4196 ( .A1(conv2_sram_rdata_weight[14]), .A2(
        conv1_sram_rdata_weight[14]), .S0(n92), .Y(conv_weight_box[10]) );
  MUX21X1_HVT U4197 ( .A1(tmp_big2[31]), .A2(tmp_big1[31]), .S0(n1504), .Y(
        data_out[31]) );
  MUX21X1_HVT U4198 ( .A1(tmp_big2[30]), .A2(tmp_big1[30]), .S0(n1504), .Y(
        data_out[30]) );
  MUX21X1_HVT U4199 ( .A1(conv2_sram_rdata_weight[25]), .A2(
        conv1_sram_rdata_weight[25]), .S0(n619), .Y(conv_weight_box[16]) );
  MUX21X1_HVT U4200 ( .A1(conv2_sram_rdata_weight[29]), .A2(
        conv1_sram_rdata_weight[29]), .S0(n619), .Y(conv_weight_box[19]) );
  MUX21X1_HVT U4201 ( .A1(conv2_sram_rdata_weight[17]), .A2(
        conv1_sram_rdata_weight[17]), .S0(n345), .Y(conv_weight_box[11]) );
  MUX21X1_HVT U4202 ( .A1(tmp_big2[29]), .A2(tmp_big1[29]), .S0(n1504), .Y(
        data_out[29]) );
  MUX21X1_HVT U4203 ( .A1(tmp_big2[26]), .A2(tmp_big1[26]), .S0(n1504), .Y(
        data_out[26]) );
  MUX21X1_HVT U4204 ( .A1(tmp_big2[6]), .A2(tmp_big1[6]), .S0(N9), .Y(
        data_out[6]) );
  MUX21X1_HVT U4205 ( .A1(tmp_big2[25]), .A2(tmp_big1[25]), .S0(n1504), .Y(
        data_out[25]) );
  MUX21X1_HVT U4206 ( .A1(tmp_big2[24]), .A2(tmp_big1[24]), .S0(n1504), .Y(
        data_out[24]) );
  MUX21X1_HVT U4207 ( .A1(tmp_big2[22]), .A2(tmp_big1[22]), .S0(n1481), .Y(
        data_out[22]) );
  MUX21X1_HVT U4208 ( .A1(conv2_sum_b[31]), .A2(conv2_sum_a[31]), .S0(n1437), 
        .Y(tmp_big1[31]) );
  MUX21X1_HVT U4209 ( .A1(conv2_sram_rdata_weight[1]), .A2(
        conv1_sram_rdata_weight[1]), .S0(n1418), .Y(conv_weight_box[0]) );
  MUX21X1_HVT U4210 ( .A1(conv2_sum_d[31]), .A2(conv2_sum_c[31]), .S0(n1532), 
        .Y(tmp_big2[31]) );
  MUX21X1_HVT U4211 ( .A1(conv2_sum_d[30]), .A2(conv2_sum_c[30]), .S0(n1496), 
        .Y(tmp_big2[30]) );
  MUX21X1_HVT U4212 ( .A1(n1881), .A2(n1882), .S0(n1430), .Y(n2164) );
  MUX21X1_HVT U4213 ( .A1(conv2_sum_b[0]), .A2(conv2_sum_a[0]), .S0(n1974), 
        .Y(tmp_big1[0]) );
  MUX21X1_HVT U4214 ( .A1(conv2_sum_d[3]), .A2(conv2_sum_c[3]), .S0(N7), .Y(
        tmp_big2[3]) );
  MUX21X1_HVT U4215 ( .A1(conv2_sum_d[2]), .A2(conv2_sum_c[2]), .S0(n1994), 
        .Y(tmp_big2[2]) );
  MUX21X1_HVT U4216 ( .A1(conv2_sum_d[4]), .A2(conv2_sum_c[4]), .S0(n1994), 
        .Y(tmp_big2[4]) );
  MUX21X2_HVT U4217 ( .A1(conv2_sram_rdata_weight[4]), .A2(
        conv1_sram_rdata_weight[4]), .S0(n345), .Y(conv_weight_box[2]) );
  INVX1_HVT U4218 ( .A(tmp_big1[29]), .Y(n2166) );
  INVX1_HVT U4219 ( .A(tmp_big2[31]), .Y(n2152) );
  INVX1_HVT U4220 ( .A(tmp_big1[23]), .Y(n2162) );
  INVX1_HVT U4221 ( .A(tmp_big1[21]), .Y(n2161) );
  INVX1_HVT U4222 ( .A(tmp_big1[19]), .Y(n2159) );
  INVX1_HVT U4223 ( .A(n2153), .Y(tmp_big1[10]) );
  AO21X1_HVT U4224 ( .A1(n2174), .A2(conv2_sum_b[9]), .A3(n2173), .Y(
        tmp_big1[9]) );
  AO22X1_HVT U4225 ( .A1(tmp_big2[10]), .A2(n2153), .A3(tmp_big2[11]), .A4(
        n2154), .Y(n2137) );
  INVX1_HVT U4226 ( .A(tmp_big1[11]), .Y(n2154) );
  INVX1_HVT U4227 ( .A(tmp_big1[15]), .Y(n2157) );
  INVX1_HVT U4228 ( .A(n1964), .Y(n1962) );
  AO22X1_HVT U4229 ( .A1(conv2_sum_d[10]), .A2(n1860), .A3(conv2_sum_d[11]), 
        .A4(n1982), .Y(n2085) );
  INVX1_HVT U4230 ( .A(conv2_sram_rdata_weight[69]), .Y(n1929) );
  INVX1_HVT U4231 ( .A(n1485), .Y(n1930) );
  INVX1_HVT U4232 ( .A(conv1_sram_rdata_weight[69]), .Y(n1931) );
  AOI22X1_HVT U4233 ( .A1(tmp_big1[25]), .A2(n1926), .A3(n1925), .A4(n2148), 
        .Y(n1848) );
  INVX1_HVT U4234 ( .A(tmp_big1[26]), .Y(n2163) );
  AOI22X1_HVT U4235 ( .A1(conv2_sum_a[13]), .A2(n1880), .A3(n1919), .A4(n2023), 
        .Y(n1870) );
  NOR3X0_HVT U4236 ( .A1(channel[2]), .A2(channel[3]), .A3(n2172), .Y(n1871)
         );
  AOI22X1_HVT U4237 ( .A1(conv2_sum_b[6]), .A2(n1861), .A3(conv2_sum_b[7]), 
        .A4(n1853), .Y(n1873) );
  NOR3X0_HVT U4238 ( .A1(n2099), .A2(n2098), .A3(n2097), .Y(n1875) );
  NOR3X0_HVT U4239 ( .A1(n2145), .A2(n2144), .A3(n2143), .Y(n1877) );
  NAND2X0_HVT U4240 ( .A1(n1952), .A2(n1951), .Y(n1878) );
  MUX21X1_HVT U4241 ( .A1(conv2_sum_b[22]), .A2(conv2_sum_a[22]), .S0(n1974), 
        .Y(tmp_big1[22]) );
  MUX21X1_HVT U4242 ( .A1(conv1_sram_rdata_weight[18]), .A2(
        conv2_sram_rdata_weight[18]), .S0(n1515), .Y(conv_weight_box[12]) );
  NAND2X0_HVT U4243 ( .A1(n1879), .A2(conv2_sum_b[13]), .Y(n2023) );
  AND2X1_HVT U4244 ( .A1(n1857), .A2(conv2_sum_a[12]), .Y(n1919) );
  NAND2X0_HVT U4245 ( .A1(n2100), .A2(n2102), .Y(n1921) );
  AND2X1_HVT U4246 ( .A1(n1964), .A2(n1875), .Y(n1922) );
  OA21X1_HVT U4247 ( .A1(n1848), .A2(n2118), .A3(n1924), .Y(n2114) );
  MUX21X1_HVT U4248 ( .A1(conv2_sum_b[26]), .A2(conv2_sum_a[26]), .S0(n1483), 
        .Y(tmp_big1[26]) );
  NAND2X0_HVT U4249 ( .A1(n2156), .A2(tmp_big2[13]), .Y(n2128) );
  MUX21X1_HVT U4250 ( .A1(n1879), .A2(n1880), .S0(n1533), .Y(n2156) );
  OR2X1_HVT U4251 ( .A1(n1927), .A2(n2126), .Y(n2144) );
  NAND2X0_HVT U4252 ( .A1(n2121), .A2(n2120), .Y(n1927) );
  AO22X1_HVT U4253 ( .A1(n619), .A2(conv1_sram_rdata_weight[72]), .A3(n1930), 
        .A4(conv2_sram_rdata_weight[72]), .Y(conv_weight_box[49]) );
  NAND4X0_HVT U4254 ( .A1(n1948), .A2(n1950), .A3(n1933), .A4(n1932), .Y(n1939) );
  AND2X1_HVT U4255 ( .A1(n1936), .A2(n1934), .Y(n1950) );
  NAND2X0_HVT U4256 ( .A1(n1935), .A2(n2135), .Y(n1934) );
  OAI22X1_HVT U4257 ( .A1(tmp_big2[13]), .A2(n2156), .A3(tmp_big2[12]), .A4(
        n2127), .Y(n1935) );
  NAND2X0_HVT U4258 ( .A1(n1937), .A2(n1952), .Y(n1948) );
  NAND2X0_HVT U4259 ( .A1(n1949), .A2(n2134), .Y(n1937) );
  NAND3X0_HVT U4260 ( .A1(n1939), .A2(n1938), .A3(n1877), .Y(n2146) );
  NAND3X0_HVT U4261 ( .A1(n1948), .A2(n1878), .A3(n1950), .Y(n1938) );
  NAND2X0_HVT U4262 ( .A1(n2146), .A2(n2147), .Y(n1969) );
  AND2X1_HVT U4263 ( .A1(n1947), .A2(n1940), .Y(n2147) );
  NAND2X0_HVT U4264 ( .A1(n1942), .A2(n1941), .Y(n1940) );
  NAND2X0_HVT U4265 ( .A1(n1944), .A2(n1943), .Y(n1942) );
  NAND2X0_HVT U4266 ( .A1(n1946), .A2(n1945), .Y(n1944) );
  OA21X1_HVT U4267 ( .A1(n2126), .A2(n2125), .A3(n2124), .Y(n1947) );
  OR2X1_HVT U4268 ( .A1(n2137), .A2(n2133), .Y(n1949) );
  AND2X1_HVT U4269 ( .A1(n2135), .A2(n1953), .Y(n1952) );
  AND2X1_HVT U4270 ( .A1(n2129), .A2(n1529), .Y(n1953) );
  NAND3X0_HVT U4271 ( .A1(n1955), .A2(n1876), .A3(n1954), .Y(n2042) );
  NAND2X0_HVT U4272 ( .A1(n1957), .A2(n1873), .Y(n1956) );
  OA21X1_HVT U4273 ( .A1(n2032), .A2(n2029), .A3(n1959), .Y(n1958) );
  OA21X1_HVT U4274 ( .A1(n2030), .A2(n1870), .A3(n2028), .Y(n1959) );
  NAND2X0_HVT U4275 ( .A1(n2102), .A2(n2101), .Y(n1963) );
  NAND2X0_HVT U4276 ( .A1(n1969), .A2(n1968), .Y(n2149) );
  NAND2X0_HVT U4277 ( .A1(n2150), .A2(n1971), .Y(n1970) );
  NAND3X0_HVT U4278 ( .A1(n2146), .A2(n2150), .A3(n2147), .Y(n1972) );
  INVX1_HVT U4279 ( .A(n1976), .Y(tmp_big1[14]) );
  MUX21X1_HVT U4280 ( .A1(n1977), .A2(n1978), .S0(n1430), .Y(n1976) );
  INVX1_HVT U4281 ( .A(n1985), .Y(tmp_big1[3]) );
  INVX1_HVT U4282 ( .A(tmp_big1[2]), .Y(n2167) );
  OR2X1_HVT U4283 ( .A1(n1984), .A2(n886), .Y(n2031) );
  OR2X1_HVT U4284 ( .A1(n1986), .A2(conv2_sum_c[11]), .Y(n2073) );
  AOI21X1_HVT U4285 ( .A1(n2174), .A2(conv2_sum_b[9]), .A3(n2173), .Y(n1990)
         );
  NAND2X0_HVT U4286 ( .A1(n2075), .A2(n2085), .Y(n1992) );
  NAND2X0_HVT U4287 ( .A1(n1991), .A2(n1992), .Y(n2079) );
  NAND2X0_HVT U4288 ( .A1(conv2_sum_b[29]), .A2(n1916), .Y(n1996) );
  NAND2X0_HVT U4289 ( .A1(conv2_sum_a[28]), .A2(n1996), .Y(n1995) );
  OA22X1_HVT U4290 ( .A1(n1916), .A2(conv2_sum_b[29]), .A3(n1995), .A4(
        conv2_sum_b[28]), .Y(n2006) );
  NAND2X0_HVT U4291 ( .A1(conv2_sum_b[28]), .A2(n1890), .Y(n1997) );
  NAND3X0_HVT U4292 ( .A1(n1997), .A2(n865), .A3(n1996), .Y(n2008) );
  NAND2X0_HVT U4293 ( .A1(conv2_sum_b[27]), .A2(n1882), .Y(n1998) );
  NAND2X0_HVT U4294 ( .A1(conv2_sum_a[26]), .A2(n1998), .Y(n1999) );
  OA22X1_HVT U4295 ( .A1(conv2_sum_b[27]), .A2(n1882), .A3(conv2_sum_b[26]), 
        .A4(n1999), .Y(n2001) );
  AO22X1_HVT U4296 ( .A1(conv2_sum_b[26]), .A2(n1889), .A3(conv2_sum_b[27]), 
        .A4(n1882), .Y(n2009) );
  AO22X1_HVT U4297 ( .A1(n2001), .A2(n2000), .A3(n2001), .A4(n2009), .Y(n2005)
         );
  NAND2X0_HVT U4298 ( .A1(conv2_sum_a[31]), .A2(n1914), .Y(n2002) );
  NAND2X0_HVT U4299 ( .A1(conv2_sum_a[30]), .A2(n2002), .Y(n2003) );
  OA22X1_HVT U4300 ( .A1(n1914), .A2(conv2_sum_a[31]), .A3(n2003), .A4(
        conv2_sum_b[30]), .Y(n2004) );
  AO22X1_HVT U4301 ( .A1(conv2_sum_b[22]), .A2(n1887), .A3(conv2_sum_b[23]), 
        .A4(n1902), .Y(n2022) );
  NAND2X0_HVT U4302 ( .A1(conv2_sum_b[21]), .A2(n1901), .Y(n2011) );
  NAND2X0_HVT U4303 ( .A1(conv2_sum_a[20]), .A2(n2011), .Y(n2010) );
  OA22X1_HVT U4304 ( .A1(n1901), .A2(conv2_sum_b[21]), .A3(n2010), .A4(
        conv2_sum_b[20]), .Y(n2021) );
  NAND2X0_HVT U4305 ( .A1(conv2_sum_b[20]), .A2(n1886), .Y(n2012) );
  NAND3X0_HVT U4306 ( .A1(n2012), .A2(n2047), .A3(n2011), .Y(n2040) );
  NAND2X0_HVT U4307 ( .A1(conv2_sum_b[19]), .A2(n1900), .Y(n2013) );
  NAND2X0_HVT U4308 ( .A1(conv2_sum_a[18]), .A2(n2013), .Y(n2014) );
  OA22X1_HVT U4309 ( .A1(conv2_sum_b[19]), .A2(n1900), .A3(conv2_sum_b[18]), 
        .A4(n2014), .Y(n2016) );
  NAND2X0_HVT U4310 ( .A1(conv2_sum_b[17]), .A2(n1899), .Y(n2039) );
  AO22X1_HVT U4311 ( .A1(conv2_sum_b[18]), .A2(n1885), .A3(conv2_sum_b[19]), 
        .A4(n1900), .Y(n2041) );
  AO22X1_HVT U4312 ( .A1(n2016), .A2(n2015), .A3(n2016), .A4(n2041), .Y(n2020)
         );
  NAND2X0_HVT U4313 ( .A1(conv2_sum_b[23]), .A2(n1902), .Y(n2017) );
  NAND2X0_HVT U4314 ( .A1(conv2_sum_a[22]), .A2(n2017), .Y(n2018) );
  OA22X1_HVT U4315 ( .A1(n1902), .A2(conv2_sum_b[23]), .A3(n2018), .A4(
        conv2_sum_b[22]), .Y(n2019) );
  AO22X1_HVT U4316 ( .A1(conv2_sum_b[14]), .A2(n1978), .A3(conv2_sum_b[15]), 
        .A4(n1898), .Y(n2030) );
  NAND2X0_HVT U4317 ( .A1(conv2_sum_b[12]), .A2(n1864), .Y(n2024) );
  NAND3X0_HVT U4318 ( .A1(n2024), .A2(n2046), .A3(n2023), .Y(n2032) );
  NAND2X0_HVT U4319 ( .A1(conv2_sum_b[15]), .A2(n1898), .Y(n2026) );
  NAND2X0_HVT U4320 ( .A1(conv2_sum_a[14]), .A2(n2026), .Y(n2027) );
  OA22X1_HVT U4321 ( .A1(n1898), .A2(conv2_sum_b[15]), .A3(n2027), .A4(
        conv2_sum_b[14]), .Y(n2028) );
  AO22X1_HVT U4322 ( .A1(conv2_sum_b[5]), .A2(n1852), .A3(conv2_sum_b[4]), 
        .A4(n1863), .Y(n2034) );
  NAND2X0_HVT U4323 ( .A1(conv2_sum_b[7]), .A2(n1853), .Y(n2035) );
  NAND2X0_HVT U4324 ( .A1(conv2_sum_a[6]), .A2(n2035), .Y(n2036) );
  OA22X1_HVT U4325 ( .A1(n1853), .A2(conv2_sum_b[7]), .A3(n2036), .A4(
        conv2_sum_b[6]), .Y(n2037) );
  OA221X1_HVT U4326 ( .A1(n2005), .A2(n2008), .A3(n2006), .A4(n2007), .A5(
        n2004), .Y(n2045) );
  AO22X1_HVT U4327 ( .A1(conv2_sum_d[30]), .A2(n1913), .A3(conv2_sum_c[31]), 
        .A4(n1915), .Y(n2059) );
  NAND2X0_HVT U4328 ( .A1(conv2_sum_d[29]), .A2(n1917), .Y(n2049) );
  NAND2X0_HVT U4329 ( .A1(conv2_sum_c[28]), .A2(n2049), .Y(n2048) );
  OA22X1_HVT U4330 ( .A1(n1917), .A2(conv2_sum_d[29]), .A3(n2048), .A4(
        conv2_sum_d[28]), .Y(n2058) );
  NAND2X0_HVT U4331 ( .A1(conv2_sum_d[28]), .A2(n1897), .Y(n2050) );
  NAND2X0_HVT U4332 ( .A1(conv2_sum_d[27]), .A2(n1911), .Y(n2051) );
  NAND2X0_HVT U4333 ( .A1(conv2_sum_c[26]), .A2(n2051), .Y(n2052) );
  OA22X1_HVT U4334 ( .A1(conv2_sum_d[27]), .A2(n1911), .A3(conv2_sum_d[26]), 
        .A4(n2052), .Y(n2054) );
  NAND2X0_HVT U4335 ( .A1(conv2_sum_d[25]), .A2(n1910), .Y(n2103) );
  AO22X1_HVT U4336 ( .A1(conv2_sum_d[26]), .A2(n1896), .A3(conv2_sum_d[27]), 
        .A4(n1911), .Y(n2061) );
  AO22X1_HVT U4337 ( .A1(n2054), .A2(n2053), .A3(n2054), .A4(n2061), .Y(n2057)
         );
  OA22X1_HVT U4338 ( .A1(n1915), .A2(conv2_sum_c[31]), .A3(n2055), .A4(
        conv2_sum_d[30]), .Y(n2056) );
  AO22X1_HVT U4339 ( .A1(conv2_sum_d[22]), .A2(n1894), .A3(conv2_sum_d[23]), 
        .A4(n1909), .Y(n2069) );
  NAND2X0_HVT U4340 ( .A1(conv2_sum_d[21]), .A2(n1908), .Y(n2063) );
  NAND2X0_HVT U4341 ( .A1(conv2_sum_c[20]), .A2(n2063), .Y(n2062) );
  NAND2X0_HVT U4342 ( .A1(conv2_sum_d[20]), .A2(n1893), .Y(n2064) );
  NAND3X0_HVT U4343 ( .A1(n2064), .A2(n2106), .A3(n2063), .Y(n2098) );
  NAND2X0_HVT U4344 ( .A1(conv2_sum_d[19]), .A2(n1907), .Y(n2065) );
  NAND2X0_HVT U4345 ( .A1(conv2_sum_c[18]), .A2(n2065), .Y(n2066) );
  NAND2X0_HVT U4346 ( .A1(conv2_sum_d[17]), .A2(n1906), .Y(n2096) );
  NAND2X0_HVT U4347 ( .A1(conv2_sum_c[16]), .A2(n2096), .Y(n2067) );
  AO22X1_HVT U4348 ( .A1(conv2_sum_d[18]), .A2(n1892), .A3(conv2_sum_d[19]), 
        .A4(n1907), .Y(n2099) );
  NAND2X0_HVT U4349 ( .A1(conv2_sum_d[23]), .A2(n1909), .Y(n2068) );
  AO22X1_HVT U4350 ( .A1(conv2_sum_d[14]), .A2(n1891), .A3(conv2_sum_d[15]), 
        .A4(n1905), .Y(n2081) );
  NAND2X0_HVT U4351 ( .A1(conv2_sum_d[13]), .A2(n1904), .Y(n2071) );
  NAND2X0_HVT U4352 ( .A1(conv2_sum_c[12]), .A2(n2071), .Y(n2070) );
  OA22X1_HVT U4353 ( .A1(n1904), .A2(conv2_sum_d[13]), .A3(n2070), .A4(
        conv2_sum_d[12]), .Y(n2080) );
  NAND2X0_HVT U4354 ( .A1(conv2_sum_d[12]), .A2(n1868), .Y(n2072) );
  NAND3X0_HVT U4355 ( .A1(n2072), .A2(n2105), .A3(n2071), .Y(n2084) );
  NAND2X0_HVT U4356 ( .A1(conv2_sum_c[10]), .A2(n2073), .Y(n2074) );
  OA22X1_HVT U4357 ( .A1(conv2_sum_d[11]), .A2(n1982), .A3(conv2_sum_d[10]), 
        .A4(n2074), .Y(n2075) );
  NAND2X0_HVT U4358 ( .A1(conv2_sum_d[9]), .A2(n1993), .Y(n2082) );
  NAND2X0_HVT U4359 ( .A1(conv2_sum_d[15]), .A2(n1905), .Y(n2076) );
  NAND2X0_HVT U4360 ( .A1(conv2_sum_c[14]), .A2(n2076), .Y(n2077) );
  OA22X1_HVT U4361 ( .A1(n1905), .A2(conv2_sum_d[15]), .A3(n2077), .A4(
        conv2_sum_d[14]), .Y(n2078) );
  OAI21X1_HVT U4362 ( .A1(conv2_sum_c[8]), .A2(n1856), .A3(n2082), .Y(n2083)
         );
  OR3X1_HVT U4363 ( .A1(n2085), .A2(n2084), .A3(n2083), .Y(n2101) );
  AO22X1_HVT U4364 ( .A1(conv2_sum_d[2]), .A2(n1865), .A3(conv2_sum_d[3]), 
        .A4(n1988), .Y(n2087) );
  AO22X1_HVT U4365 ( .A1(conv2_sum_d[5]), .A2(n1854), .A3(conv2_sum_d[4]), 
        .A4(n1859), .Y(n2086) );
  AO22X1_HVT U4366 ( .A1(conv2_sum_d[6]), .A2(n1862), .A3(conv2_sum_d[7]), 
        .A4(n1855), .Y(n2094) );
  NAND2X0_HVT U4367 ( .A1(conv2_sum_d[5]), .A2(n1854), .Y(n2088) );
  NAND2X0_HVT U4368 ( .A1(conv2_sum_c[4]), .A2(n2088), .Y(n2089) );
  OA22X1_HVT U4369 ( .A1(n2089), .A2(conv2_sum_d[4]), .A3(n1854), .A4(
        conv2_sum_d[5]), .Y(n2093) );
  NAND2X0_HVT U4370 ( .A1(conv2_sum_d[7]), .A2(n1855), .Y(n2090) );
  NAND2X0_HVT U4371 ( .A1(conv2_sum_c[6]), .A2(n2090), .Y(n2091) );
  OA22X1_HVT U4372 ( .A1(n1855), .A2(conv2_sum_d[7]), .A3(n2091), .A4(
        conv2_sum_d[6]), .Y(n2092) );
  OA221X1_HVT U4373 ( .A1(n2094), .A2(n2095), .A3(n2093), .A4(n2094), .A5(
        n2092), .Y(n2100) );
  OAI21X1_HVT U4374 ( .A1(conv2_sum_c[16]), .A2(n1884), .A3(n2096), .Y(n2097)
         );
  OA221X1_HVT U4375 ( .A1(n2057), .A2(n2060), .A3(n2058), .A4(n2059), .A5(
        n2056), .Y(n2104) );
  OA221X1_HVT U4376 ( .A1(n2084), .A2(n2079), .A3(n2080), .A4(n2081), .A5(
        n2078), .Y(n2102) );
  AO22X1_HVT U4377 ( .A1(tmp_big2[30]), .A2(n2168), .A3(tmp_big1[31]), .A4(
        n2152), .Y(n2116) );
  NAND2X0_HVT U4378 ( .A1(tmp_big2[29]), .A2(n2166), .Y(n2109) );
  NAND2X0_HVT U4379 ( .A1(tmp_big1[28]), .A2(n2109), .Y(n2108) );
  OA22X1_HVT U4380 ( .A1(n2166), .A2(tmp_big2[29]), .A3(n2108), .A4(
        tmp_big2[28]), .Y(n2115) );
  NAND2X0_HVT U4381 ( .A1(tmp_big2[28]), .A2(n2165), .Y(n2110) );
  NAND3X0_HVT U4382 ( .A1(n2110), .A2(n2169), .A3(n2109), .Y(n2117) );
  AO22X1_HVT U4383 ( .A1(tmp_big2[26]), .A2(n2163), .A3(tmp_big2[27]), .A4(
        n2164), .Y(n2118) );
  NAND2X0_HVT U4384 ( .A1(tmp_big1[31]), .A2(n2152), .Y(n2111) );
  NAND2X0_HVT U4385 ( .A1(tmp_big1[30]), .A2(n2111), .Y(n2112) );
  OA22X1_HVT U4386 ( .A1(n2152), .A2(tmp_big1[31]), .A3(n2112), .A4(
        tmp_big2[30]), .Y(n2113) );
  NAND2X0_HVT U4387 ( .A1(tmp_big2[21]), .A2(n2161), .Y(n2120) );
  NAND2X0_HVT U4388 ( .A1(tmp_big1[20]), .A2(n2120), .Y(n2119) );
  OA22X1_HVT U4389 ( .A1(n2161), .A2(tmp_big2[21]), .A3(n2119), .A4(
        tmp_big2[20]), .Y(n2125) );
  NAND2X0_HVT U4390 ( .A1(tmp_big2[20]), .A2(n2160), .Y(n2121) );
  AO22X1_HVT U4391 ( .A1(tmp_big2[18]), .A2(n2158), .A3(tmp_big2[19]), .A4(
        n2159), .Y(n2145) );
  NAND2X0_HVT U4392 ( .A1(tmp_big2[23]), .A2(n2162), .Y(n2122) );
  NAND2X0_HVT U4393 ( .A1(tmp_big1[22]), .A2(n2122), .Y(n2123) );
  OA22X1_HVT U4394 ( .A1(n2162), .A2(tmp_big2[23]), .A3(n2123), .A4(
        tmp_big2[22]), .Y(n2124) );
  NAND2X0_HVT U4395 ( .A1(tmp_big1[12]), .A2(n2128), .Y(n2127) );
  NAND2X0_HVT U4396 ( .A1(tmp_big2[12]), .A2(n2155), .Y(n2129) );
  NAND2X0_HVT U4397 ( .A1(tmp_big2[11]), .A2(n2154), .Y(n2130) );
  NAND2X0_HVT U4398 ( .A1(tmp_big1[10]), .A2(n2130), .Y(n2131) );
  OA22X1_HVT U4399 ( .A1(tmp_big2[11]), .A2(n2154), .A3(tmp_big2[10]), .A4(
        n2131), .Y(n2134) );
  NAND2X0_HVT U4400 ( .A1(tmp_big2[9]), .A2(n1990), .Y(n2136) );
  NAND2X0_HVT U4401 ( .A1(tmp_big1[8]), .A2(n2136), .Y(n2132) );
  OA22X1_HVT U4402 ( .A1(n1979), .A2(tmp_big2[9]), .A3(n2132), .A4(tmp_big2[8]), .Y(n2133) );
  NAND2X0_HVT U4403 ( .A1(tmp_big2[3]), .A2(n1985), .Y(n2138) );
  NAND2X0_HVT U4404 ( .A1(n2138), .A2(tmp_big1[2]), .Y(n2139) );
  OAI21X1_HVT U4405 ( .A1(tmp_big1[16]), .A2(n2151), .A3(n2142), .Y(n2143) );
  OA221X1_HVT U4406 ( .A1(n2114), .A2(n2117), .A3(n2115), .A4(n2116), .A5(
        n2113), .Y(n2150) );
  OR3X1_HVT U4407 ( .A1(channel[4]), .A2(channel[0]), .A3(channel[1]), .Y(
        n2172) );
  MUX21X1_HVT U4408 ( .A1(conv2_sum_b[30]), .A2(conv2_sum_a[30]), .S0(n1430), 
        .Y(tmp_big1[30]) );
  MUX21X1_HVT U4409 ( .A1(conv2_sum_b[29]), .A2(conv2_sum_a[29]), .S0(n1483), 
        .Y(tmp_big1[29]) );
  MUX21X1_HVT U4410 ( .A1(conv2_sum_b[28]), .A2(conv2_sum_a[28]), .S0(n1437), 
        .Y(tmp_big1[28]) );
  MUX21X1_HVT U4411 ( .A1(conv2_sum_b[25]), .A2(conv2_sum_a[25]), .S0(n1502), 
        .Y(tmp_big1[25]) );
  MUX21X1_HVT U4412 ( .A1(conv2_sum_b[23]), .A2(conv2_sum_a[23]), .S0(n1483), 
        .Y(tmp_big1[23]) );
  MUX21X1_HVT U4413 ( .A1(conv2_sum_b[21]), .A2(conv2_sum_a[21]), .S0(n1430), 
        .Y(tmp_big1[21]) );
  MUX21X1_HVT U4414 ( .A1(conv2_sum_b[20]), .A2(conv2_sum_a[20]), .S0(n1429), 
        .Y(tmp_big1[20]) );
  MUX21X1_HVT U4415 ( .A1(conv2_sum_b[19]), .A2(conv2_sum_a[19]), .S0(n1429), 
        .Y(tmp_big1[19]) );
  MUX21X1_HVT U4416 ( .A1(conv2_sum_b[18]), .A2(conv2_sum_a[18]), .S0(n1437), 
        .Y(tmp_big1[18]) );
  MUX21X1_HVT U4417 ( .A1(conv2_sum_b[16]), .A2(conv2_sum_a[16]), .S0(n1437), 
        .Y(tmp_big1[16]) );
  MUX21X1_HVT U4418 ( .A1(conv2_sum_b[12]), .A2(conv2_sum_a[12]), .S0(n1429), 
        .Y(tmp_big1[12]) );
  MUX21X1_HVT U4419 ( .A1(conv2_sum_d[29]), .A2(conv2_sum_c[29]), .S0(n1532), 
        .Y(tmp_big2[29]) );
  MUX21X1_HVT U4420 ( .A1(conv2_sum_d[28]), .A2(conv2_sum_c[28]), .S0(n1496), 
        .Y(tmp_big2[28]) );
  MUX21X1_HVT U4421 ( .A1(conv2_sum_d[27]), .A2(conv2_sum_c[27]), .S0(n1532), 
        .Y(tmp_big2[27]) );
  MUX21X1_HVT U4422 ( .A1(conv2_sum_d[26]), .A2(conv2_sum_c[26]), .S0(n1994), 
        .Y(tmp_big2[26]) );
  MUX21X1_HVT U4423 ( .A1(conv2_sum_d[25]), .A2(conv2_sum_c[25]), .S0(n1532), 
        .Y(tmp_big2[25]) );
  MUX21X1_HVT U4424 ( .A1(conv2_sum_d[24]), .A2(conv2_sum_c[24]), .S0(n1496), 
        .Y(tmp_big2[24]) );
  MUX21X1_HVT U4425 ( .A1(conv2_sum_d[23]), .A2(conv2_sum_c[23]), .S0(n1532), 
        .Y(tmp_big2[23]) );
  MUX21X1_HVT U4426 ( .A1(conv2_sum_d[21]), .A2(conv2_sum_c[21]), .S0(n1532), 
        .Y(tmp_big2[21]) );
  MUX21X1_HVT U4427 ( .A1(conv2_sum_d[20]), .A2(conv2_sum_c[20]), .S0(n1496), 
        .Y(tmp_big2[20]) );
  MUX21X1_HVT U4428 ( .A1(conv2_sum_d[19]), .A2(conv2_sum_c[19]), .S0(n1532), 
        .Y(tmp_big2[19]) );
  MUX21X1_HVT U4429 ( .A1(conv2_sum_d[18]), .A2(conv2_sum_c[18]), .S0(n1994), 
        .Y(tmp_big2[18]) );
  MUX21X1_HVT U4430 ( .A1(conv2_sum_d[16]), .A2(conv2_sum_c[16]), .S0(n1994), 
        .Y(tmp_big2[16]) );
  MUX21X1_HVT U4431 ( .A1(conv2_sum_d[15]), .A2(conv2_sum_c[15]), .S0(n1532), 
        .Y(tmp_big2[15]) );
  MUX21X1_HVT U4432 ( .A1(conv2_sum_d[14]), .A2(conv2_sum_c[14]), .S0(n1496), 
        .Y(tmp_big2[14]) );
  MUX21X1_HVT U4433 ( .A1(conv2_sum_d[13]), .A2(conv2_sum_c[13]), .S0(N7), .Y(
        tmp_big2[13]) );
  MUX21X1_HVT U4434 ( .A1(conv2_sum_d[12]), .A2(conv2_sum_c[12]), .S0(n1496), 
        .Y(tmp_big2[12]) );
  MUX21X1_HVT U4435 ( .A1(conv2_sum_d[11]), .A2(conv2_sum_c[11]), .S0(n1532), 
        .Y(tmp_big2[11]) );
  MUX21X1_HVT U4436 ( .A1(conv2_sum_d[10]), .A2(conv2_sum_c[10]), .S0(n1496), 
        .Y(tmp_big2[10]) );
  MUX21X1_HVT U4437 ( .A1(conv2_sum_d[7]), .A2(conv2_sum_c[7]), .S0(N7), .Y(
        tmp_big2[7]) );
  MUX21X1_HVT U4438 ( .A1(conv2_sum_d[6]), .A2(conv2_sum_c[6]), .S0(n1994), 
        .Y(tmp_big2[6]) );
  NAND2X0_HVT U4439 ( .A1(N7), .A2(conv2_sum_c[1]), .Y(n2176) );
  MUX21X1_HVT U4440 ( .A1(tmp_big2[0]), .A2(tmp_big1[0]), .S0(n1967), .Y(
        data_out[0]) );
  NAND2X0_HVT U4441 ( .A1(n2176), .A2(n2175), .Y(n2177) );
  MUX21X1_HVT U4442 ( .A1(n2177), .A2(tmp_big1[1]), .S0(n1967), .Y(data_out[1]) );
  MUX21X1_HVT U4443 ( .A1(tmp_big2[2]), .A2(tmp_big1[2]), .S0(n1967), .Y(
        data_out[2]) );
  MUX21X1_HVT U4444 ( .A1(tmp_big2[3]), .A2(tmp_big1[3]), .S0(n1967), .Y(
        data_out[3]) );
  MUX21X1_HVT U4445 ( .A1(tmp_big2[4]), .A2(tmp_big1[4]), .S0(n1967), .Y(
        data_out[4]) );
  MUX21X1_HVT U4446 ( .A1(tmp_big2[7]), .A2(tmp_big1[7]), .S0(n1504), .Y(
        data_out[7]) );
  MUX21X1_HVT U4447 ( .A1(tmp_big2[12]), .A2(tmp_big1[12]), .S0(n1504), .Y(
        data_out[12]) );
  MUX21X1_HVT U4448 ( .A1(tmp_big2[13]), .A2(tmp_big1[13]), .S0(n1481), .Y(
        data_out[13]) );
  MUX21X1_HVT U4449 ( .A1(tmp_big2[16]), .A2(tmp_big1[16]), .S0(n1482), .Y(
        data_out[16]) );
  MUX21X1_HVT U4450 ( .A1(tmp_big2[17]), .A2(tmp_big1[17]), .S0(n1482), .Y(
        data_out[17]) );
  MUX21X1_HVT U4451 ( .A1(tmp_big2[18]), .A2(tmp_big1[18]), .S0(n1482), .Y(
        data_out[18]) );
  MUX21X1_HVT U4452 ( .A1(tmp_big2[20]), .A2(tmp_big1[20]), .S0(n1504), .Y(
        data_out[20]) );
endmodule


module quantize ( clk, srstn, bias_data, mode, quantized_data, ori_data_31_, 
        ori_data_30_, ori_data_29_, ori_data_28_, ori_data_27_, ori_data_26_, 
        ori_data_25_, ori_data_24_, ori_data_23_, ori_data_22_, ori_data_21_, 
        ori_data_20_, ori_data_19_, ori_data_18_, ori_data_17_, ori_data_16_, 
        ori_data_15_, ori_data_14_, ori_data_13_, ori_data_12_, ori_data_11_, 
        ori_data_10_, ori_data_9_, ori_data_8_, ori_data_7_, ori_data_6_, 
        ori_data_5_ );
  input [3:0] bias_data;
  input [1:0] mode;
  output [7:0] quantized_data;
  input clk, srstn, ori_data_31_, ori_data_30_, ori_data_29_, ori_data_28_,
         ori_data_27_, ori_data_26_, ori_data_25_, ori_data_24_, ori_data_23_,
         ori_data_22_, ori_data_21_, ori_data_20_, ori_data_19_, ori_data_18_,
         ori_data_17_, ori_data_16_, ori_data_15_, ori_data_14_, ori_data_13_,
         ori_data_12_, ori_data_11_, ori_data_10_, ori_data_9_, ori_data_8_,
         ori_data_7_, ori_data_6_, ori_data_5_;
  wire   N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N59, N60, N61, N113, N114, N115, N116, N117, N118, N119,
         N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130,
         N131, n13, DP_OP_26J6_124_4249_n594, DP_OP_26J6_124_4249_n593,
         DP_OP_26J6_124_4249_n592, DP_OP_26J6_124_4249_n590,
         DP_OP_26J6_124_4249_n588, DP_OP_26J6_124_4249_n586,
         DP_OP_26J6_124_4249_n584, DP_OP_26J6_124_4249_n582,
         DP_OP_26J6_124_4249_n580, DP_OP_26J6_124_4249_n578,
         DP_OP_26J6_124_4249_n576, DP_OP_26J6_124_4249_n571,
         DP_OP_26J6_124_4249_n570, DP_OP_26J6_124_4249_n568,
         DP_OP_26J6_124_4249_n567, DP_OP_26J6_124_4249_n566,
         DP_OP_26J6_124_4249_n560, DP_OP_26J6_124_4249_n559,
         DP_OP_26J6_124_4249_n558, DP_OP_26J6_124_4249_n553,
         DP_OP_26J6_124_4249_n552, DP_OP_26J6_124_4249_n545,
         DP_OP_26J6_124_4249_n544, DP_OP_26J6_124_4249_n543,
         DP_OP_26J6_124_4249_n538, DP_OP_26J6_124_4249_n537,
         DP_OP_26J6_124_4249_n536, DP_OP_26J6_124_4249_n535,
         DP_OP_26J6_124_4249_n530, DP_OP_26J6_124_4249_n527,
         DP_OP_26J6_124_4249_n526, DP_OP_26J6_124_4249_n525,
         DP_OP_26J6_124_4249_n524, DP_OP_26J6_124_4249_n523,
         DP_OP_26J6_124_4249_n520, DP_OP_26J6_124_4249_n519,
         DP_OP_26J6_124_4249_n518, DP_OP_26J6_124_4249_n517,
         DP_OP_26J6_124_4249_n508, DP_OP_26J6_124_4249_n507,
         DP_OP_26J6_124_4249_n506, DP_OP_26J6_124_4249_n501,
         DP_OP_26J6_124_4249_n500, DP_OP_26J6_124_4249_n498,
         DP_OP_26J6_124_4249_n497, DP_OP_26J6_124_4249_n496,
         DP_OP_26J6_124_4249_n495, DP_OP_26J6_124_4249_n490,
         DP_OP_26J6_124_4249_n488, DP_OP_26J6_124_4249_n487,
         DP_OP_26J6_124_4249_n485, DP_OP_26J6_124_4249_n484,
         DP_OP_26J6_124_4249_n479, DP_OP_26J6_124_4249_n478,
         DP_OP_26J6_124_4249_n477, DP_OP_26J6_124_4249_n476,
         DP_OP_26J6_124_4249_n475, DP_OP_26J6_124_4249_n474,
         DP_OP_26J6_124_4249_n473, DP_OP_26J6_124_4249_n468,
         DP_OP_26J6_124_4249_n466, DP_OP_26J6_124_4249_n465,
         DP_OP_26J6_124_4249_n464, DP_OP_26J6_124_4249_n463,
         DP_OP_26J6_124_4249_n462, DP_OP_26J6_124_4249_n458,
         DP_OP_26J6_124_4249_n457, DP_OP_26J6_124_4249_n456,
         DP_OP_26J6_124_4249_n455, DP_OP_26J6_124_4249_n454,
         DP_OP_26J6_124_4249_n452, DP_OP_26J6_124_4249_n447,
         DP_OP_26J6_124_4249_n446, DP_OP_26J6_124_4249_n445,
         DP_OP_26J6_124_4249_n442, DP_OP_26J6_124_4249_n441,
         DP_OP_26J6_124_4249_n440, DP_OP_26J6_124_4249_n436,
         DP_OP_26J6_124_4249_n435, DP_OP_26J6_124_4249_n434,
         DP_OP_26J6_124_4249_n432, DP_OP_26J6_124_4249_n431,
         DP_OP_26J6_124_4249_n421, DP_OP_26J6_124_4249_n420,
         DP_OP_26J6_124_4249_n415, DP_OP_26J6_124_4249_n414,
         DP_OP_26J6_124_4249_n413, DP_OP_26J6_124_4249_n412,
         DP_OP_26J6_124_4249_n411, DP_OP_26J6_124_4249_n410,
         DP_OP_26J6_124_4249_n409, DP_OP_26J6_124_4249_n404,
         DP_OP_26J6_124_4249_n402, DP_OP_26J6_124_4249_n401,
         DP_OP_26J6_124_4249_n399, DP_OP_26J6_124_4249_n398,
         DP_OP_26J6_124_4249_n397, DP_OP_26J6_124_4249_n396,
         DP_OP_26J6_124_4249_n393, DP_OP_26J6_124_4249_n392,
         DP_OP_26J6_124_4249_n391, DP_OP_26J6_124_4249_n390,
         DP_OP_26J6_124_4249_n389, DP_OP_26J6_124_4249_n388,
         DP_OP_26J6_124_4249_n387, DP_OP_26J6_124_4249_n382,
         DP_OP_26J6_124_4249_n380, DP_OP_26J6_124_4249_n379,
         DP_OP_26J6_124_4249_n377, DP_OP_26J6_124_4249_n376,
         DP_OP_26J6_124_4249_n373, DP_OP_26J6_124_4249_n372,
         DP_OP_26J6_124_4249_n371, DP_OP_26J6_124_4249_n370,
         DP_OP_26J6_124_4249_n369, DP_OP_26J6_124_4249_n368,
         DP_OP_26J6_124_4249_n367, DP_OP_26J6_124_4249_n366,
         DP_OP_26J6_124_4249_n361, DP_OP_26J6_124_4249_n360,
         DP_OP_26J6_124_4249_n359, DP_OP_26J6_124_4249_n358,
         DP_OP_26J6_124_4249_n357, DP_OP_26J6_124_4249_n356,
         DP_OP_26J6_124_4249_n355, DP_OP_26J6_124_4249_n354,
         DP_OP_26J6_124_4249_n352, DP_OP_26J6_124_4249_n350,
         DP_OP_26J6_124_4249_n349, DP_OP_26J6_124_4249_n348,
         DP_OP_26J6_124_4249_n347, DP_OP_26J6_124_4249_n346,
         DP_OP_26J6_124_4249_n345, DP_OP_26J6_124_4249_n344,
         DP_OP_26J6_124_4249_n342, DP_OP_26J6_124_4249_n336,
         DP_OP_26J6_124_4249_n335, DP_OP_26J6_124_4249_n333,
         DP_OP_26J6_124_4249_n331, DP_OP_26J6_124_4249_n325,
         DP_OP_26J6_124_4249_n324, DP_OP_26J6_124_4249_n323,
         DP_OP_26J6_124_4249_n322, DP_OP_26J6_124_4249_n320,
         DP_OP_26J6_124_4249_n319, DP_OP_26J6_124_4249_n318,
         DP_OP_26J6_124_4249_n317, DP_OP_26J6_124_4249_n316,
         DP_OP_26J6_124_4249_n315, DP_OP_26J6_124_4249_n314,
         DP_OP_26J6_124_4249_n313, DP_OP_26J6_124_4249_n312,
         DP_OP_26J6_124_4249_n311, DP_OP_26J6_124_4249_n310,
         DP_OP_26J6_124_4249_n309, DP_OP_26J6_124_4249_n308,
         DP_OP_26J6_124_4249_n307, DP_OP_26J6_124_4249_n306,
         DP_OP_26J6_124_4249_n304, DP_OP_26J6_124_4249_n303,
         DP_OP_26J6_124_4249_n302, DP_OP_26J6_124_4249_n301,
         DP_OP_26J6_124_4249_n300, DP_OP_26J6_124_4249_n299,
         DP_OP_26J6_124_4249_n298, DP_OP_26J6_124_4249_n297,
         DP_OP_26J6_124_4249_n296, DP_OP_26J6_124_4249_n295,
         DP_OP_26J6_124_4249_n291, DP_OP_26J6_124_4249_n290,
         DP_OP_26J6_124_4249_n289, DP_OP_26J6_124_4249_n287,
         DP_OP_26J6_124_4249_n285, DP_OP_26J6_124_4249_n283,
         DP_OP_26J6_124_4249_n281, DP_OP_26J6_124_4249_n279,
         DP_OP_26J6_124_4249_n277, DP_OP_26J6_124_4249_n271,
         DP_OP_26J6_124_4249_n265, DP_OP_26J6_124_4249_n263,
         DP_OP_26J6_124_4249_n262, DP_OP_26J6_124_4249_n261,
         DP_OP_26J6_124_4249_n260, DP_OP_26J6_124_4249_n259,
         DP_OP_26J6_124_4249_n258, DP_OP_26J6_124_4249_n253,
         DP_OP_26J6_124_4249_n252, DP_OP_26J6_124_4249_n251,
         DP_OP_26J6_124_4249_n250, DP_OP_26J6_124_4249_n249,
         DP_OP_26J6_124_4249_n248, DP_OP_26J6_124_4249_n247,
         DP_OP_26J6_124_4249_n246, DP_OP_26J6_124_4249_n245,
         DP_OP_26J6_124_4249_n238, DP_OP_26J6_124_4249_n237,
         DP_OP_26J6_124_4249_n236, DP_OP_26J6_124_4249_n233,
         DP_OP_26J6_124_4249_n232, DP_OP_26J6_124_4249_n231,
         DP_OP_26J6_124_4249_n230, DP_OP_26J6_124_4249_n229,
         DP_OP_26J6_124_4249_n228, DP_OP_26J6_124_4249_n223,
         DP_OP_26J6_124_4249_n222, DP_OP_26J6_124_4249_n221,
         DP_OP_26J6_124_4249_n220, DP_OP_26J6_124_4249_n219,
         DP_OP_26J6_124_4249_n218, DP_OP_26J6_124_4249_n217,
         DP_OP_26J6_124_4249_n216, DP_OP_26J6_124_4249_n215,
         DP_OP_26J6_124_4249_n214, DP_OP_26J6_124_4249_n213,
         DP_OP_26J6_124_4249_n211, DP_OP_26J6_124_4249_n210,
         DP_OP_26J6_124_4249_n201, DP_OP_26J6_124_4249_n200,
         DP_OP_26J6_124_4249_n199, DP_OP_26J6_124_4249_n194,
         DP_OP_26J6_124_4249_n193, DP_OP_26J6_124_4249_n192,
         DP_OP_26J6_124_4249_n191, DP_OP_26J6_124_4249_n190,
         DP_OP_26J6_124_4249_n189, DP_OP_26J6_124_4249_n188,
         DP_OP_26J6_124_4249_n183, DP_OP_26J6_124_4249_n181,
         DP_OP_26J6_124_4249_n180, DP_OP_26J6_124_4249_n179,
         DP_OP_26J6_124_4249_n178, DP_OP_26J6_124_4249_n177,
         DP_OP_26J6_124_4249_n175, DP_OP_26J6_124_4249_n172,
         DP_OP_26J6_124_4249_n171, DP_OP_26J6_124_4249_n170,
         DP_OP_26J6_124_4249_n169, DP_OP_26J6_124_4249_n168,
         DP_OP_26J6_124_4249_n167, DP_OP_26J6_124_4249_n166,
         DP_OP_26J6_124_4249_n161, DP_OP_26J6_124_4249_n159,
         DP_OP_26J6_124_4249_n158, DP_OP_26J6_124_4249_n157,
         DP_OP_26J6_124_4249_n156, DP_OP_26J6_124_4249_n155,
         DP_OP_26J6_124_4249_n152, DP_OP_26J6_124_4249_n151,
         DP_OP_26J6_124_4249_n150, DP_OP_26J6_124_4249_n149,
         DP_OP_26J6_124_4249_n148, DP_OP_26J6_124_4249_n147,
         DP_OP_26J6_124_4249_n146, DP_OP_26J6_124_4249_n145,
         DP_OP_26J6_124_4249_n140, DP_OP_26J6_124_4249_n139,
         DP_OP_26J6_124_4249_n138, DP_OP_26J6_124_4249_n137,
         DP_OP_26J6_124_4249_n136, DP_OP_26J6_124_4249_n135,
         DP_OP_26J6_124_4249_n134, DP_OP_26J6_124_4249_n133,
         DP_OP_26J6_124_4249_n132, DP_OP_26J6_124_4249_n131,
         DP_OP_26J6_124_4249_n130, DP_OP_26J6_124_4249_n129,
         DP_OP_26J6_124_4249_n128, DP_OP_26J6_124_4249_n127,
         DP_OP_26J6_124_4249_n125, DP_OP_26J6_124_4249_n124,
         DP_OP_26J6_124_4249_n114, DP_OP_26J6_124_4249_n113,
         DP_OP_26J6_124_4249_n108, DP_OP_26J6_124_4249_n107,
         DP_OP_26J6_124_4249_n106, DP_OP_26J6_124_4249_n103,
         DP_OP_26J6_124_4249_n102, DP_OP_26J6_124_4249_n97,
         DP_OP_26J6_124_4249_n96, DP_OP_26J6_124_4249_n95,
         DP_OP_26J6_124_4249_n94, DP_OP_26J6_124_4249_n93,
         DP_OP_26J6_124_4249_n92, DP_OP_26J6_124_4249_n91,
         DP_OP_26J6_124_4249_n90, DP_OP_26J6_124_4249_n89,
         DP_OP_26J6_124_4249_n86, DP_OP_26J6_124_4249_n85,
         DP_OP_26J6_124_4249_n84, DP_OP_26J6_124_4249_n83,
         DP_OP_26J6_124_4249_n82, DP_OP_26J6_124_4249_n81,
         DP_OP_26J6_124_4249_n80, DP_OP_26J6_124_4249_n75,
         DP_OP_26J6_124_4249_n74, DP_OP_26J6_124_4249_n73,
         DP_OP_26J6_124_4249_n72, DP_OP_26J6_124_4249_n71,
         DP_OP_26J6_124_4249_n70, DP_OP_26J6_124_4249_n69,
         DP_OP_26J6_124_4249_n66, DP_OP_26J6_124_4249_n65,
         DP_OP_26J6_124_4249_n64, DP_OP_26J6_124_4249_n63,
         DP_OP_26J6_124_4249_n59, DP_OP_26J6_124_4249_n54,
         DP_OP_26J6_124_4249_n53, DP_OP_26J6_124_4249_n52,
         DP_OP_26J6_124_4249_n51, DP_OP_26J6_124_4249_n50,
         DP_OP_26J6_124_4249_n49, DP_OP_26J6_124_4249_n48,
         DP_OP_26J6_124_4249_n47, DP_OP_26J6_124_4249_n46,
         DP_OP_26J6_124_4249_n45, DP_OP_26J6_124_4249_n44,
         DP_OP_26J6_124_4249_n43, DP_OP_26J6_124_4249_n42,
         DP_OP_26J6_124_4249_n41, DP_OP_26J6_124_4249_n33,
         DP_OP_26J6_124_4249_n32, DP_OP_26J6_124_4249_n31,
         DP_OP_26J6_124_4249_n30, DP_OP_26J6_124_4249_n25,
         DP_OP_26J6_124_4249_n24, DP_OP_26J6_124_4249_n23,
         DP_OP_26J6_124_4249_n22, DP_OP_26J6_124_4249_n21,
         DP_OP_26J6_124_4249_n20, DP_OP_26J6_124_4249_n19,
         DP_OP_26J6_124_4249_n18, DP_OP_26J6_124_4249_n17,
         DP_OP_26J6_124_4249_n16, DP_OP_26J6_124_4249_n15,
         DP_OP_26J6_124_4249_n14, DP_OP_26J6_124_4249_n13,
         DP_OP_26J6_124_4249_n12, DP_OP_26J6_124_4249_n11,
         DP_OP_26J6_124_4249_n10, DP_OP_26J6_124_4249_n9,
         DP_OP_26J6_124_4249_n8, DP_OP_26J6_124_4249_n7,
         DP_OP_26J6_124_4249_n6, DP_OP_26J6_124_4249_n4,
         DP_OP_26J6_124_4249_n2, DP_OP_26J6_124_4249_n1, n1, n2, n3, n4, n5,
         n6, n7, n9, n10, n11, n12, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n430, n440, n450, n460, n470, n480,
         n490, n510, n520, n530, n540, n550, n560, n570, n580, n590, n600,
         n610, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n92, n93, n94, n95, n96, n97, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n1130, n1140,
         n1150, n1160, n1170, n1180, n1190, n1200, n1210, n1220, n1230, n1240,
         n1250, n1260, n1270, n1280, n1290, n1300, n1310, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188;
  wire   [7:0] n_quantized_data;

  DFFSSRX1_HVT quantized_data_reg_7_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[7]), .CLK(clk), .Q(quantized_data[7]) );
  DFFSSRX1_HVT quantized_data_reg_6_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[6]), .CLK(clk), .Q(quantized_data[6]) );
  DFFSSRX1_HVT quantized_data_reg_5_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[5]), .CLK(clk), .Q(quantized_data[5]) );
  DFFSSRX1_HVT quantized_data_reg_4_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[4]), .CLK(clk), .Q(quantized_data[4]) );
  DFFSSRX1_HVT quantized_data_reg_3_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[3]), .CLK(clk), .Q(quantized_data[3]) );
  DFFSSRX1_HVT quantized_data_reg_2_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[2]), .CLK(clk), .Q(quantized_data[2]) );
  DFFSSRX1_HVT quantized_data_reg_1_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[1]), .CLK(clk), .Q(quantized_data[1]) );
  DFFSSRX1_HVT quantized_data_reg_0_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[0]), .CLK(clk), .Q(quantized_data[0]) );
  XNOR2X2_HVT DP_OP_26J6_124_4249_U2 ( .A1(DP_OP_26J6_124_4249_n31), .A2(
        DP_OP_26J6_124_4249_n2), .Y(N131) );
  XNOR2X2_HVT DP_OP_26J6_124_4249_U322 ( .A1(DP_OP_26J6_124_4249_n323), .A2(
        DP_OP_26J6_124_4249_n295), .Y(N61) );
  XNOR2X2_HVT DP_OP_26J6_124_4249_U17 ( .A1(DP_OP_26J6_124_4249_n49), .A2(
        DP_OP_26J6_124_4249_n4), .Y(N129) );
  XNOR2X2_HVT DP_OP_26J6_124_4249_U425 ( .A1(DP_OP_26J6_124_4249_n411), .A2(
        DP_OP_26J6_124_4249_n303), .Y(N53) );
  XNOR2X2_HVT DP_OP_26J6_124_4249_U341 ( .A1(DP_OP_26J6_124_4249_n345), .A2(
        DP_OP_26J6_124_4249_n297), .Y(N59) );
  XNOR2X2_HVT DP_OP_26J6_124_4249_U397 ( .A1(DP_OP_26J6_124_4249_n389), .A2(
        DP_OP_26J6_124_4249_n301), .Y(N55) );
  XNOR2X2_HVT DP_OP_26J6_124_4249_U369 ( .A1(DP_OP_26J6_124_4249_n367), .A2(
        DP_OP_26J6_124_4249_n299), .Y(N57) );
  XNOR2X2_HVT DP_OP_26J6_124_4249_U355 ( .A1(DP_OP_26J6_124_4249_n356), .A2(
        DP_OP_26J6_124_4249_n298), .Y(N58) );
  XNOR2X2_HVT DP_OP_26J6_124_4249_U535 ( .A1(DP_OP_26J6_124_4249_n497), .A2(
        DP_OP_26J6_124_4249_n311), .Y(N45) );
  XNOR2X2_HVT DP_OP_26J6_124_4249_U549 ( .A1(DP_OP_26J6_124_4249_n508), .A2(
        DP_OP_26J6_124_4249_n312), .Y(N44) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U296 ( .A1(DP_OP_26J6_124_4249_n258), .A2(
        DP_OP_26J6_124_4249_n260), .A3(DP_OP_26J6_124_4249_n259), .Y(
        DP_OP_26J6_124_4249_n253) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U36 ( .A1(DP_OP_26J6_124_4249_n54), .A2(
        DP_OP_26J6_124_4249_n66), .A3(DP_OP_26J6_124_4249_n59), .Y(
        DP_OP_26J6_124_4249_n53) );
  XOR2X1_HVT DP_OP_26J6_124_4249_U239 ( .A1(DP_OP_26J6_124_4249_n220), .A2(
        DP_OP_26J6_124_4249_n20), .Y(N113) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U253 ( .A1(DP_OP_26J6_124_4249_n223), .A2(
        DP_OP_26J6_124_4249_n233), .A3(DP_OP_26J6_124_4249_n228), .Y(
        DP_OP_26J6_124_4249_n222) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U146 ( .A1(DP_OP_26J6_124_4249_n140), .A2(
        DP_OP_26J6_124_4249_n152), .A3(DP_OP_26J6_124_4249_n145), .Y(
        DP_OP_26J6_124_4249_n139) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U26 ( .A1(DP_OP_26J6_124_4249_n59), .A2(
        DP_OP_26J6_124_4249_n47), .A3(DP_OP_26J6_124_4249_n48), .Y(
        DP_OP_26J6_124_4249_n46) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U54 ( .A1(DP_OP_26J6_124_4249_n81), .A2(
        DP_OP_26J6_124_4249_n69), .A3(DP_OP_26J6_124_4249_n70), .Y(
        DP_OP_26J6_124_4249_n64) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U82 ( .A1(DP_OP_26J6_124_4249_n103), .A2(
        DP_OP_26J6_124_4249_n91), .A3(DP_OP_26J6_124_4249_n92), .Y(
        DP_OP_26J6_124_4249_n90) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U136 ( .A1(DP_OP_26J6_124_4249_n145), .A2(
        DP_OP_26J6_124_4249_n133), .A3(DP_OP_26J6_124_4249_n134), .Y(
        DP_OP_26J6_124_4249_n132) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U245 ( .A1(DP_OP_26J6_124_4249_n228), .A2(
        DP_OP_26J6_124_4249_n218), .A3(DP_OP_26J6_124_4249_n219), .Y(
        DP_OP_26J6_124_4249_n217) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U374 ( .A1(DP_OP_26J6_124_4249_n361), .A2(
        DP_OP_26J6_124_4249_n373), .A3(DP_OP_26J6_124_4249_n366), .Y(
        DP_OP_26J6_124_4249_n360) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U392 ( .A1(DP_OP_26J6_124_4249_n388), .A2(
        DP_OP_26J6_124_4249_n376), .A3(DP_OP_26J6_124_4249_n377), .Y(
        DP_OP_26J6_124_4249_n371) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U484 ( .A1(DP_OP_26J6_124_4249_n447), .A2(
        n103), .A3(DP_OP_26J6_124_4249_n452), .Y(DP_OP_26J6_124_4249_n446) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U583 ( .A1(DP_OP_26J6_124_4249_n535), .A2(
        DP_OP_26J6_124_4249_n525), .A3(DP_OP_26J6_124_4249_n526), .Y(
        DP_OP_26J6_124_4249_n524) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U649 ( .A1(ori_data_6_), .A2(bias_data[1]), 
        .Y(DP_OP_26J6_124_4249_n570) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U646 ( .A1(n1200), .A2(
        DP_OP_26J6_124_4249_n570), .Y(DP_OP_26J6_124_4249_n320) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U639 ( .A1(n1180), .A2(
        DP_OP_26J6_124_4249_n566), .Y(DP_OP_26J6_124_4249_n319) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U632 ( .A1(ori_data_8_), .A2(n1260), .Y(
        DP_OP_26J6_124_4249_n559) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U629 ( .A1(n1170), .A2(
        DP_OP_26J6_124_4249_n559), .Y(DP_OP_26J6_124_4249_n318) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U623 ( .A1(ori_data_9_), .A2(n1270), .Y(
        DP_OP_26J6_124_4249_n553) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U620 ( .A1(DP_OP_26J6_124_4249_n594), .A2(
        DP_OP_26J6_124_4249_n553), .Y(DP_OP_26J6_124_4249_n317) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U611 ( .A1(ori_data_10_), .A2(n1280), .Y(
        DP_OP_26J6_124_4249_n544) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U610 ( .A1(n1260), .A2(ori_data_10_), .Y(
        DP_OP_26J6_124_4249_n543) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U608 ( .A1(DP_OP_26J6_124_4249_n593), .A2(
        DP_OP_26J6_124_4249_n544), .Y(DP_OP_26J6_124_4249_n316) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U606 ( .A1(DP_OP_26J6_124_4249_n543), .A2(
        DP_OP_26J6_124_4249_n552), .Y(DP_OP_26J6_124_4249_n537) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U599 ( .A1(ori_data_11_), .A2(n1270), .Y(
        DP_OP_26J6_124_4249_n535) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U596 ( .A1(DP_OP_26J6_124_4249_n592), .A2(
        DP_OP_26J6_124_4249_n535), .Y(DP_OP_26J6_124_4249_n315) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U587 ( .A1(ori_data_12_), .A2(n1250), .Y(
        DP_OP_26J6_124_4249_n526) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U586 ( .A1(n1260), .A2(ori_data_12_), .Y(
        DP_OP_26J6_124_4249_n525) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U584 ( .A1(DP_OP_26J6_124_4249_n287), .A2(
        DP_OP_26J6_124_4249_n526), .Y(DP_OP_26J6_124_4249_n314) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U582 ( .A1(DP_OP_26J6_124_4249_n530), .A2(
        DP_OP_26J6_124_4249_n525), .Y(DP_OP_26J6_124_4249_n523) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U576 ( .A1(ori_data_13_), .A2(n1270), .Y(
        DP_OP_26J6_124_4249_n518) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U575 ( .A1(n1280), .A2(ori_data_13_), .Y(
        DP_OP_26J6_124_4249_n517) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U573 ( .A1(DP_OP_26J6_124_4249_n590), .A2(
        DP_OP_26J6_124_4249_n518), .Y(DP_OP_26J6_124_4249_n313) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U562 ( .A1(ori_data_14_), .A2(n1250), .Y(
        DP_OP_26J6_124_4249_n507) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U561 ( .A1(bias_data[3]), .A2(ori_data_14_), 
        .Y(DP_OP_26J6_124_4249_n506) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U559 ( .A1(DP_OP_26J6_124_4249_n285), .A2(
        DP_OP_26J6_124_4249_n507), .Y(DP_OP_26J6_124_4249_n312) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U557 ( .A1(DP_OP_26J6_124_4249_n506), .A2(
        DP_OP_26J6_124_4249_n517), .Y(DP_OP_26J6_124_4249_n500) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U548 ( .A1(n1240), .A2(ori_data_15_), .Y(
        DP_OP_26J6_124_4249_n496) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U545 ( .A1(DP_OP_26J6_124_4249_n588), .A2(
        DP_OP_26J6_124_4249_n496), .Y(DP_OP_26J6_124_4249_n311) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U538 ( .A1(DP_OP_26J6_124_4249_n501), .A2(
        DP_OP_26J6_124_4249_n588), .A3(DP_OP_26J6_124_4249_n490), .Y(
        DP_OP_26J6_124_4249_n488) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U537 ( .A1(DP_OP_26J6_124_4249_n500), .A2(
        DP_OP_26J6_124_4249_n588), .Y(DP_OP_26J6_124_4249_n487) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U534 ( .A1(ori_data_16_), .A2(n1270), .Y(
        DP_OP_26J6_124_4249_n485) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U533 ( .A1(n1280), .A2(ori_data_16_), .Y(
        DP_OP_26J6_124_4249_n484) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U531 ( .A1(DP_OP_26J6_124_4249_n283), .A2(
        DP_OP_26J6_124_4249_n485), .Y(DP_OP_26J6_124_4249_n310) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U520 ( .A1(ori_data_17_), .A2(n1260), .Y(
        DP_OP_26J6_124_4249_n474) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U517 ( .A1(DP_OP_26J6_124_4249_n586), .A2(
        DP_OP_26J6_124_4249_n474), .Y(DP_OP_26J6_124_4249_n309) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U509 ( .A1(DP_OP_26J6_124_4249_n478), .A2(
        DP_OP_26J6_124_4249_n586), .Y(DP_OP_26J6_124_4249_n465) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U506 ( .A1(ori_data_18_), .A2(n1270), .Y(
        DP_OP_26J6_124_4249_n463) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U505 ( .A1(n1260), .A2(ori_data_18_), .Y(
        DP_OP_26J6_124_4249_n462) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U503 ( .A1(DP_OP_26J6_124_4249_n281), .A2(
        DP_OP_26J6_124_4249_n463), .Y(DP_OP_26J6_124_4249_n308) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U501 ( .A1(DP_OP_26J6_124_4249_n462), .A2(
        DP_OP_26J6_124_4249_n473), .Y(DP_OP_26J6_124_4249_n456) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U496 ( .A1(DP_OP_26J6_124_4249_n479), .A2(
        DP_OP_26J6_124_4249_n456), .A3(DP_OP_26J6_124_4249_n457), .Y(
        DP_OP_26J6_124_4249_n455) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U495 ( .A1(DP_OP_26J6_124_4249_n478), .A2(
        DP_OP_26J6_124_4249_n456), .Y(DP_OP_26J6_124_4249_n454) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U492 ( .A1(n1240), .A2(ori_data_19_), .Y(
        DP_OP_26J6_124_4249_n452) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U489 ( .A1(DP_OP_26J6_124_4249_n584), .A2(
        DP_OP_26J6_124_4249_n452), .Y(DP_OP_26J6_124_4249_n307) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U483 ( .A1(DP_OP_26J6_124_4249_n447), .A2(
        DP_OP_26J6_124_4249_n458), .Y(DP_OP_26J6_124_4249_n445) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U478 ( .A1(ori_data_20_), .A2(n1260), .Y(
        DP_OP_26J6_124_4249_n441) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U475 ( .A1(DP_OP_26J6_124_4249_n279), .A2(
        DP_OP_26J6_124_4249_n441), .Y(DP_OP_26J6_124_4249_n306) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U469 ( .A1(DP_OP_26J6_124_4249_n436), .A2(
        DP_OP_26J6_124_4249_n476), .Y(DP_OP_26J6_124_4249_n434) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U466 ( .A1(ori_data_21_), .A2(n1260), .Y(
        DP_OP_26J6_124_4249_n432) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U452 ( .A1(ori_data_22_), .A2(n1270), .Y(
        DP_OP_26J6_124_4249_n421) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U451 ( .A1(n1280), .A2(ori_data_22_), .Y(
        DP_OP_26J6_124_4249_n420) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U449 ( .A1(DP_OP_26J6_124_4249_n277), .A2(
        DP_OP_26J6_124_4249_n421), .Y(DP_OP_26J6_124_4249_n304) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U447 ( .A1(DP_OP_26J6_124_4249_n420), .A2(
        DP_OP_26J6_124_4249_n431), .Y(DP_OP_26J6_124_4249_n414) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U438 ( .A1(ori_data_23_), .A2(bias_data[3]), 
        .Y(DP_OP_26J6_124_4249_n410) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U437 ( .A1(n1260), .A2(ori_data_23_), .Y(
        DP_OP_26J6_124_4249_n409) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U435 ( .A1(DP_OP_26J6_124_4249_n580), .A2(
        DP_OP_26J6_124_4249_n410), .Y(DP_OP_26J6_124_4249_n303) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U428 ( .A1(DP_OP_26J6_124_4249_n415), .A2(
        DP_OP_26J6_124_4249_n580), .A3(DP_OP_26J6_124_4249_n404), .Y(
        DP_OP_26J6_124_4249_n402) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U427 ( .A1(DP_OP_26J6_124_4249_n414), .A2(
        DP_OP_26J6_124_4249_n580), .Y(DP_OP_26J6_124_4249_n401) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U424 ( .A1(ori_data_24_), .A2(n1250), .Y(
        DP_OP_26J6_124_4249_n399) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U421 ( .A1(DP_OP_26J6_124_4249_n96), .A2(
        DP_OP_26J6_124_4249_n399), .Y(DP_OP_26J6_124_4249_n302) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U419 ( .A1(DP_OP_26J6_124_4249_n398), .A2(
        DP_OP_26J6_124_4249_n409), .Y(DP_OP_26J6_124_4249_n396) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U418 ( .A1(DP_OP_26J6_124_4249_n415), .A2(
        DP_OP_26J6_124_4249_n396), .A3(DP_OP_26J6_124_4249_n397), .Y(
        DP_OP_26J6_124_4249_n391) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U417 ( .A1(DP_OP_26J6_124_4249_n414), .A2(
        DP_OP_26J6_124_4249_n396), .Y(DP_OP_26J6_124_4249_n390) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U410 ( .A1(ori_data_25_), .A2(n1280), .Y(
        DP_OP_26J6_124_4249_n388) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U407 ( .A1(DP_OP_26J6_124_4249_n578), .A2(
        DP_OP_26J6_124_4249_n388), .Y(DP_OP_26J6_124_4249_n301) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U400 ( .A1(DP_OP_26J6_124_4249_n393), .A2(
        DP_OP_26J6_124_4249_n578), .A3(DP_OP_26J6_124_4249_n382), .Y(
        DP_OP_26J6_124_4249_n380) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U399 ( .A1(DP_OP_26J6_124_4249_n392), .A2(
        DP_OP_26J6_124_4249_n578), .Y(DP_OP_26J6_124_4249_n379) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U396 ( .A1(ori_data_26_), .A2(n1270), .Y(
        DP_OP_26J6_124_4249_n377) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U393 ( .A1(DP_OP_26J6_124_4249_n74), .A2(
        DP_OP_26J6_124_4249_n377), .Y(DP_OP_26J6_124_4249_n300) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U391 ( .A1(DP_OP_26J6_124_4249_n376), .A2(
        DP_OP_26J6_124_4249_n387), .Y(DP_OP_26J6_124_4249_n370) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U386 ( .A1(DP_OP_26J6_124_4249_n393), .A2(
        DP_OP_26J6_124_4249_n370), .A3(DP_OP_26J6_124_4249_n371), .Y(
        DP_OP_26J6_124_4249_n369) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U385 ( .A1(DP_OP_26J6_124_4249_n392), .A2(
        DP_OP_26J6_124_4249_n370), .Y(DP_OP_26J6_124_4249_n368) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U382 ( .A1(ori_data_27_), .A2(n1260), .Y(
        DP_OP_26J6_124_4249_n366) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U381 ( .A1(n1280), .A2(ori_data_27_), .Y(
        DP_OP_26J6_124_4249_n361) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U379 ( .A1(DP_OP_26J6_124_4249_n576), .A2(
        DP_OP_26J6_124_4249_n366), .Y(DP_OP_26J6_124_4249_n299) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U373 ( .A1(DP_OP_26J6_124_4249_n361), .A2(
        DP_OP_26J6_124_4249_n372), .Y(DP_OP_26J6_124_4249_n359) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U372 ( .A1(DP_OP_26J6_124_4249_n393), .A2(
        DP_OP_26J6_124_4249_n359), .A3(DP_OP_26J6_124_4249_n360), .Y(
        DP_OP_26J6_124_4249_n358) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U371 ( .A1(DP_OP_26J6_124_4249_n359), .A2(
        DP_OP_26J6_124_4249_n392), .Y(DP_OP_26J6_124_4249_n357) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U368 ( .A1(ori_data_28_), .A2(n1280), .Y(
        DP_OP_26J6_124_4249_n355) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U367 ( .A1(n1280), .A2(ori_data_28_), .Y(
        DP_OP_26J6_124_4249_n354) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U365 ( .A1(DP_OP_26J6_124_4249_n271), .A2(
        DP_OP_26J6_124_4249_n355), .Y(DP_OP_26J6_124_4249_n298) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U363 ( .A1(DP_OP_26J6_124_4249_n354), .A2(
        DP_OP_26J6_124_4249_n361), .Y(DP_OP_26J6_124_4249_n352) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U361 ( .A1(DP_OP_26J6_124_4249_n370), .A2(
        DP_OP_26J6_124_4249_n352), .Y(DP_OP_26J6_124_4249_n350) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U359 ( .A1(DP_OP_26J6_124_4249_n350), .A2(
        DP_OP_26J6_124_4249_n390), .Y(DP_OP_26J6_124_4249_n348) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U354 ( .A1(ori_data_29_), .A2(n1270), .Y(
        DP_OP_26J6_124_4249_n344) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U351 ( .A1(n148), .A2(
        DP_OP_26J6_124_4249_n344), .Y(DP_OP_26J6_124_4249_n297) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U344 ( .A1(DP_OP_26J6_124_4249_n349), .A2(
        n148), .A3(DP_OP_26J6_124_4249_n342), .Y(DP_OP_26J6_124_4249_n336) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U343 ( .A1(DP_OP_26J6_124_4249_n348), .A2(
        n148), .Y(DP_OP_26J6_124_4249_n335) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U340 ( .A1(ori_data_30_), .A2(n1260), .Y(
        DP_OP_26J6_124_4249_n333) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U337 ( .A1(n146), .A2(
        DP_OP_26J6_124_4249_n333), .Y(DP_OP_26J6_124_4249_n296) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U330 ( .A1(DP_OP_26J6_124_4249_n349), .A2(
        n147), .A3(n143), .Y(DP_OP_26J6_124_4249_n325) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U329 ( .A1(DP_OP_26J6_124_4249_n348), .A2(
        n147), .Y(DP_OP_26J6_124_4249_n324) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U326 ( .A1(ori_data_31_), .A2(n1280), .Y(
        DP_OP_26J6_124_4249_n322) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U323 ( .A1(n142), .A2(
        DP_OP_26J6_124_4249_n322), .Y(DP_OP_26J6_124_4249_n295) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U312 ( .A1(ori_data_6_), .A2(ori_data_5_), 
        .Y(DP_OP_26J6_124_4249_n263) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U307 ( .A1(DP_OP_26J6_124_4249_n262), .A2(
        DP_OP_26J6_124_4249_n263), .Y(DP_OP_26J6_124_4249_n261) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U304 ( .A1(ori_data_8_), .A2(bias_data[0]), 
        .Y(DP_OP_26J6_124_4249_n259) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U301 ( .A1(DP_OP_26J6_124_4249_n291), .A2(
        DP_OP_26J6_124_4249_n259), .Y(DP_OP_26J6_124_4249_n25) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U294 ( .A1(ori_data_9_), .A2(bias_data[1]), 
        .Y(DP_OP_26J6_124_4249_n252) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U291 ( .A1(DP_OP_26J6_124_4249_n290), .A2(
        DP_OP_26J6_124_4249_n252), .Y(DP_OP_26J6_124_4249_n24) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U289 ( .A1(DP_OP_26J6_124_4249_n251), .A2(
        DP_OP_26J6_124_4249_n258), .Y(DP_OP_26J6_124_4249_n249) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U288 ( .A1(DP_OP_26J6_124_4249_n249), .A2(
        DP_OP_26J6_124_4249_n261), .A3(DP_OP_26J6_124_4249_n250), .Y(
        DP_OP_26J6_124_4249_n248) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U285 ( .A1(ori_data_10_), .A2(bias_data[2]), 
        .Y(DP_OP_26J6_124_4249_n246) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U282 ( .A1(DP_OP_26J6_124_4249_n289), .A2(
        DP_OP_26J6_124_4249_n246), .Y(DP_OP_26J6_124_4249_n23) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U273 ( .A1(ori_data_11_), .A2(bias_data[3]), 
        .Y(DP_OP_26J6_124_4249_n237) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U272 ( .A1(n1230), .A2(ori_data_11_), .Y(
        DP_OP_26J6_124_4249_n236) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U270 ( .A1(DP_OP_26J6_124_4249_n592), .A2(
        DP_OP_26J6_124_4249_n237), .Y(DP_OP_26J6_124_4249_n22) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U268 ( .A1(DP_OP_26J6_124_4249_n236), .A2(
        DP_OP_26J6_124_4249_n245), .Y(DP_OP_26J6_124_4249_n230) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U261 ( .A1(ori_data_12_), .A2(n1250), .Y(
        DP_OP_26J6_124_4249_n228) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U258 ( .A1(DP_OP_26J6_124_4249_n287), .A2(
        DP_OP_26J6_124_4249_n228), .Y(DP_OP_26J6_124_4249_n21) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U252 ( .A1(DP_OP_26J6_124_4249_n223), .A2(
        DP_OP_26J6_124_4249_n232), .Y(DP_OP_26J6_124_4249_n221) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U251 ( .A1(DP_OP_26J6_124_4249_n247), .A2(
        DP_OP_26J6_124_4249_n221), .A3(DP_OP_26J6_124_4249_n222), .Y(
        DP_OP_26J6_124_4249_n220) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U249 ( .A1(ori_data_13_), .A2(bias_data[3]), 
        .Y(DP_OP_26J6_124_4249_n219) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U248 ( .A1(bias_data[3]), .A2(ori_data_13_), 
        .Y(DP_OP_26J6_124_4249_n218) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U246 ( .A1(DP_OP_26J6_124_4249_n590), .A2(
        DP_OP_26J6_124_4249_n219), .Y(DP_OP_26J6_124_4249_n20) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U244 ( .A1(DP_OP_26J6_124_4249_n218), .A2(
        DP_OP_26J6_124_4249_n223), .Y(DP_OP_26J6_124_4249_n216) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U242 ( .A1(DP_OP_26J6_124_4249_n216), .A2(
        DP_OP_26J6_124_4249_n230), .Y(DP_OP_26J6_124_4249_n214) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U238 ( .A1(ori_data_14_), .A2(n1240), .Y(
        DP_OP_26J6_124_4249_n211) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U235 ( .A1(DP_OP_26J6_124_4249_n285), .A2(
        DP_OP_26J6_124_4249_n211), .Y(DP_OP_26J6_124_4249_n19) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U224 ( .A1(n1240), .A2(ori_data_15_), .Y(
        DP_OP_26J6_124_4249_n200) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U223 ( .A1(n1230), .A2(ori_data_15_), .Y(
        DP_OP_26J6_124_4249_n199) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U221 ( .A1(DP_OP_26J6_124_4249_n588), .A2(
        DP_OP_26J6_124_4249_n200), .Y(DP_OP_26J6_124_4249_n18) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U219 ( .A1(DP_OP_26J6_124_4249_n199), .A2(
        DP_OP_26J6_124_4249_n210), .Y(DP_OP_26J6_124_4249_n193) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U210 ( .A1(ori_data_16_), .A2(n1250), .Y(
        DP_OP_26J6_124_4249_n189) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U209 ( .A1(n1280), .A2(ori_data_16_), .Y(
        DP_OP_26J6_124_4249_n188) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U207 ( .A1(DP_OP_26J6_124_4249_n283), .A2(
        DP_OP_26J6_124_4249_n189), .Y(DP_OP_26J6_124_4249_n17) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U199 ( .A1(DP_OP_26J6_124_4249_n193), .A2(
        DP_OP_26J6_124_4249_n283), .Y(DP_OP_26J6_124_4249_n180) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U196 ( .A1(ori_data_17_), .A2(n1240), .Y(
        DP_OP_26J6_124_4249_n178) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U195 ( .A1(n1280), .A2(ori_data_17_), .Y(
        DP_OP_26J6_124_4249_n177) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U193 ( .A1(DP_OP_26J6_124_4249_n586), .A2(
        DP_OP_26J6_124_4249_n178), .Y(DP_OP_26J6_124_4249_n16) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U191 ( .A1(DP_OP_26J6_124_4249_n177), .A2(
        DP_OP_26J6_124_4249_n188), .Y(DP_OP_26J6_124_4249_n175) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U189 ( .A1(DP_OP_26J6_124_4249_n193), .A2(
        DP_OP_26J6_124_4249_n175), .Y(DP_OP_26J6_124_4249_n169) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U182 ( .A1(ori_data_18_), .A2(n1240), .Y(
        DP_OP_26J6_124_4249_n167) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U181 ( .A1(bias_data[3]), .A2(ori_data_18_), 
        .Y(DP_OP_26J6_124_4249_n166) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U179 ( .A1(DP_OP_26J6_124_4249_n281), .A2(
        DP_OP_26J6_124_4249_n167), .Y(DP_OP_26J6_124_4249_n15) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U172 ( .A1(DP_OP_26J6_124_4249_n172), .A2(
        DP_OP_26J6_124_4249_n281), .A3(DP_OP_26J6_124_4249_n161), .Y(
        DP_OP_26J6_124_4249_n159) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U171 ( .A1(DP_OP_26J6_124_4249_n171), .A2(
        DP_OP_26J6_124_4249_n281), .Y(DP_OP_26J6_124_4249_n158) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U168 ( .A1(ori_data_19_), .A2(n1230), .Y(
        DP_OP_26J6_124_4249_n156) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U167 ( .A1(n1250), .A2(ori_data_19_), .Y(
        DP_OP_26J6_124_4249_n155) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U165 ( .A1(DP_OP_26J6_124_4249_n584), .A2(
        DP_OP_26J6_124_4249_n156), .Y(DP_OP_26J6_124_4249_n14) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U157 ( .A1(DP_OP_26J6_124_4249_n171), .A2(
        DP_OP_26J6_124_4249_n149), .Y(DP_OP_26J6_124_4249_n147) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U154 ( .A1(ori_data_20_), .A2(n1240), .Y(
        DP_OP_26J6_124_4249_n145) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U153 ( .A1(n1250), .A2(ori_data_20_), .Y(
        DP_OP_26J6_124_4249_n140) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U151 ( .A1(DP_OP_26J6_124_4249_n279), .A2(
        DP_OP_26J6_124_4249_n145), .Y(DP_OP_26J6_124_4249_n13) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U145 ( .A1(DP_OP_26J6_124_4249_n140), .A2(
        DP_OP_26J6_124_4249_n151), .Y(DP_OP_26J6_124_4249_n138) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U144 ( .A1(DP_OP_26J6_124_4249_n172), .A2(
        DP_OP_26J6_124_4249_n138), .A3(DP_OP_26J6_124_4249_n139), .Y(
        DP_OP_26J6_124_4249_n137) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U143 ( .A1(DP_OP_26J6_124_4249_n138), .A2(
        DP_OP_26J6_124_4249_n171), .Y(DP_OP_26J6_124_4249_n136) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U140 ( .A1(ori_data_21_), .A2(n1240), .Y(
        DP_OP_26J6_124_4249_n134) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U137 ( .A1(DP_OP_26J6_124_4249_n582), .A2(
        DP_OP_26J6_124_4249_n134), .Y(DP_OP_26J6_124_4249_n12) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U135 ( .A1(DP_OP_26J6_124_4249_n133), .A2(
        DP_OP_26J6_124_4249_n140), .Y(DP_OP_26J6_124_4249_n131) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U134 ( .A1(DP_OP_26J6_124_4249_n150), .A2(
        DP_OP_26J6_124_4249_n131), .A3(DP_OP_26J6_124_4249_n132), .Y(
        DP_OP_26J6_124_4249_n130) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U133 ( .A1(DP_OP_26J6_124_4249_n149), .A2(
        DP_OP_26J6_124_4249_n131), .Y(DP_OP_26J6_124_4249_n129) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U131 ( .A1(DP_OP_26J6_124_4249_n129), .A2(
        DP_OP_26J6_124_4249_n169), .Y(DP_OP_26J6_124_4249_n127) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U128 ( .A1(ori_data_22_), .A2(n1230), .Y(
        DP_OP_26J6_124_4249_n125) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U125 ( .A1(DP_OP_26J6_124_4249_n277), .A2(
        DP_OP_26J6_124_4249_n125), .Y(DP_OP_26J6_124_4249_n11) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U114 ( .A1(ori_data_23_), .A2(n1250), .Y(
        DP_OP_26J6_124_4249_n114) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U113 ( .A1(n1230), .A2(ori_data_23_), .Y(
        DP_OP_26J6_124_4249_n113) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U111 ( .A1(DP_OP_26J6_124_4249_n580), .A2(
        DP_OP_26J6_124_4249_n114), .Y(DP_OP_26J6_124_4249_n10) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U109 ( .A1(DP_OP_26J6_124_4249_n113), .A2(
        DP_OP_26J6_124_4249_n124), .Y(DP_OP_26J6_124_4249_n107) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U100 ( .A1(ori_data_24_), .A2(n1250), .Y(
        DP_OP_26J6_124_4249_n103) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U99 ( .A1(n1230), .A2(ori_data_24_), .Y(
        DP_OP_26J6_124_4249_n102) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U97 ( .A1(DP_OP_26J6_124_4249_n96), .A2(
        DP_OP_26J6_124_4249_n103), .Y(DP_OP_26J6_124_4249_n9) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U90 ( .A1(DP_OP_26J6_124_4249_n108), .A2(
        DP_OP_26J6_124_4249_n96), .A3(DP_OP_26J6_124_4249_n97), .Y(
        DP_OP_26J6_124_4249_n95) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U89 ( .A1(DP_OP_26J6_124_4249_n107), .A2(
        DP_OP_26J6_124_4249_n96), .Y(DP_OP_26J6_124_4249_n94) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U86 ( .A1(ori_data_25_), .A2(n1250), .Y(
        DP_OP_26J6_124_4249_n92) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U83 ( .A1(DP_OP_26J6_124_4249_n578), .A2(
        DP_OP_26J6_124_4249_n92), .Y(DP_OP_26J6_124_4249_n8) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U81 ( .A1(DP_OP_26J6_124_4249_n91), .A2(
        DP_OP_26J6_124_4249_n102), .Y(DP_OP_26J6_124_4249_n89) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U80 ( .A1(DP_OP_26J6_124_4249_n108), .A2(
        DP_OP_26J6_124_4249_n89), .A3(DP_OP_26J6_124_4249_n90), .Y(
        DP_OP_26J6_124_4249_n84) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U79 ( .A1(DP_OP_26J6_124_4249_n107), .A2(
        DP_OP_26J6_124_4249_n89), .Y(DP_OP_26J6_124_4249_n83) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U72 ( .A1(ori_data_26_), .A2(n1250), .Y(
        DP_OP_26J6_124_4249_n81) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U71 ( .A1(bias_data[3]), .A2(ori_data_26_), 
        .Y(DP_OP_26J6_124_4249_n80) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U69 ( .A1(DP_OP_26J6_124_4249_n74), .A2(
        DP_OP_26J6_124_4249_n81), .Y(DP_OP_26J6_124_4249_n7) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U62 ( .A1(DP_OP_26J6_124_4249_n86), .A2(
        DP_OP_26J6_124_4249_n74), .A3(DP_OP_26J6_124_4249_n75), .Y(
        DP_OP_26J6_124_4249_n73) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U61 ( .A1(DP_OP_26J6_124_4249_n85), .A2(
        DP_OP_26J6_124_4249_n74), .Y(DP_OP_26J6_124_4249_n72) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U58 ( .A1(ori_data_27_), .A2(bias_data[3]), 
        .Y(DP_OP_26J6_124_4249_n70) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U57 ( .A1(bias_data[3]), .A2(ori_data_27_), 
        .Y(DP_OP_26J6_124_4249_n69) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U55 ( .A1(DP_OP_26J6_124_4249_n576), .A2(
        DP_OP_26J6_124_4249_n70), .Y(DP_OP_26J6_124_4249_n6) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U53 ( .A1(DP_OP_26J6_124_4249_n69), .A2(
        DP_OP_26J6_124_4249_n80), .Y(DP_OP_26J6_124_4249_n63) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U44 ( .A1(ori_data_28_), .A2(n1240), .Y(
        DP_OP_26J6_124_4249_n59) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U43 ( .A1(n1230), .A2(ori_data_28_), .Y(
        DP_OP_26J6_124_4249_n54) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U35 ( .A1(DP_OP_26J6_124_4249_n54), .A2(
        DP_OP_26J6_124_4249_n65), .Y(DP_OP_26J6_124_4249_n52) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U34 ( .A1(DP_OP_26J6_124_4249_n86), .A2(
        DP_OP_26J6_124_4249_n52), .A3(DP_OP_26J6_124_4249_n53), .Y(
        DP_OP_26J6_124_4249_n51) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U33 ( .A1(DP_OP_26J6_124_4249_n52), .A2(
        DP_OP_26J6_124_4249_n85), .Y(DP_OP_26J6_124_4249_n50) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U30 ( .A1(ori_data_29_), .A2(n1230), .Y(
        DP_OP_26J6_124_4249_n48) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U27 ( .A1(n148), .A2(DP_OP_26J6_124_4249_n48), .Y(DP_OP_26J6_124_4249_n4) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U25 ( .A1(DP_OP_26J6_124_4249_n47), .A2(
        DP_OP_26J6_124_4249_n54), .Y(DP_OP_26J6_124_4249_n45) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U24 ( .A1(DP_OP_26J6_124_4249_n64), .A2(
        DP_OP_26J6_124_4249_n45), .A3(DP_OP_26J6_124_4249_n46), .Y(
        DP_OP_26J6_124_4249_n44) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U23 ( .A1(DP_OP_26J6_124_4249_n63), .A2(
        DP_OP_26J6_124_4249_n45), .Y(DP_OP_26J6_124_4249_n43) );
  AOI21X1_HVT DP_OP_26J6_124_4249_U10 ( .A1(DP_OP_26J6_124_4249_n42), .A2(n144), .A3(DP_OP_26J6_124_4249_n331), .Y(DP_OP_26J6_124_4249_n33) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U9 ( .A1(DP_OP_26J6_124_4249_n41), .A2(n144), 
        .Y(DP_OP_26J6_124_4249_n32) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U6 ( .A1(ori_data_31_), .A2(n1240), .Y(
        DP_OP_26J6_124_4249_n30) );
  NAND2X0_HVT DP_OP_26J6_124_4249_U3 ( .A1(n141), .A2(DP_OP_26J6_124_4249_n30), 
        .Y(DP_OP_26J6_124_4249_n2) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U423 ( .A1(n1280), .A2(ori_data_24_), .Y(
        DP_OP_26J6_124_4249_n398) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U85 ( .A1(n1230), .A2(ori_data_25_), .Y(
        DP_OP_26J6_124_4249_n91) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U260 ( .A1(n1250), .A2(ori_data_12_), .Y(
        DP_OP_26J6_124_4249_n223) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U29 ( .A1(n1240), .A2(ori_data_29_), .Y(
        DP_OP_26J6_124_4249_n47) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U284 ( .A1(bias_data[2]), .A2(ori_data_10_), 
        .Y(DP_OP_26J6_124_4249_n245) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U395 ( .A1(n1270), .A2(ori_data_26_), .Y(
        DP_OP_26J6_124_4249_n376) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U607 ( .A1(DP_OP_26J6_124_4249_n553), .A2(
        DP_OP_26J6_124_4249_n543), .A3(DP_OP_26J6_124_4249_n544), .Y(
        DP_OP_26J6_124_4249_n538) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U303 ( .A1(bias_data[0]), .A2(ori_data_8_), 
        .Y(DP_OP_26J6_124_4249_n258) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U127 ( .A1(n1240), .A2(ori_data_22_), .Y(
        DP_OP_26J6_124_4249_n124) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U448 ( .A1(DP_OP_26J6_124_4249_n432), .A2(
        DP_OP_26J6_124_4249_n420), .A3(DP_OP_26J6_124_4249_n421), .Y(
        DP_OP_26J6_124_4249_n415) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U269 ( .A1(DP_OP_26J6_124_4249_n246), .A2(
        DP_OP_26J6_124_4249_n236), .A3(DP_OP_26J6_124_4249_n237), .Y(
        DP_OP_26J6_124_4249_n231) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U110 ( .A1(DP_OP_26J6_124_4249_n125), .A2(
        DP_OP_26J6_124_4249_n113), .A3(DP_OP_26J6_124_4249_n114), .Y(
        DP_OP_26J6_124_4249_n108) );
  OAI21X1_HVT DP_OP_26J6_124_4249_U22 ( .A1(DP_OP_26J6_124_4249_n43), .A2(
        DP_OP_26J6_124_4249_n84), .A3(DP_OP_26J6_124_4249_n44), .Y(
        DP_OP_26J6_124_4249_n42) );
  XNOR2X1_HVT DP_OP_26J6_124_4249_U155 ( .A1(DP_OP_26J6_124_4249_n157), .A2(
        DP_OP_26J6_124_4249_n14), .Y(N119) );
  XNOR2X1_HVT DP_OP_26J6_124_4249_U59 ( .A1(DP_OP_26J6_124_4249_n82), .A2(
        DP_OP_26J6_124_4249_n7), .Y(N126) );
  XNOR2X1_HVT DP_OP_26J6_124_4249_U169 ( .A1(DP_OP_26J6_124_4249_n168), .A2(
        DP_OP_26J6_124_4249_n15), .Y(N118) );
  XNOR2X1_HVT DP_OP_26J6_124_4249_U73 ( .A1(DP_OP_26J6_124_4249_n93), .A2(
        DP_OP_26J6_124_4249_n8), .Y(N125) );
  XNOR2X1_HVT DP_OP_26J6_124_4249_U129 ( .A1(DP_OP_26J6_124_4249_n135), .A2(
        DP_OP_26J6_124_4249_n12), .Y(N121) );
  XNOR2X1_HVT DP_OP_26J6_124_4249_U183 ( .A1(DP_OP_26J6_124_4249_n179), .A2(
        DP_OP_26J6_124_4249_n16), .Y(N117) );
  XNOR2X1_HVT DP_OP_26J6_124_4249_U45 ( .A1(DP_OP_26J6_124_4249_n71), .A2(
        DP_OP_26J6_124_4249_n6), .Y(N127) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U477 ( .A1(n1260), .A2(ori_data_20_), .Y(
        DP_OP_26J6_124_4249_n440) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U622 ( .A1(n1260), .A2(ori_data_9_), .Y(
        DP_OP_26J6_124_4249_n552) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U293 ( .A1(bias_data[1]), .A2(ori_data_9_), 
        .Y(DP_OP_26J6_124_4249_n251) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U139 ( .A1(n1230), .A2(ori_data_21_), .Y(
        DP_OP_26J6_124_4249_n133) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U465 ( .A1(n1260), .A2(ori_data_21_), .Y(
        DP_OP_26J6_124_4249_n431) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U237 ( .A1(n1240), .A2(ori_data_14_), .Y(
        DP_OP_26J6_124_4249_n210) );
  NOR2X1_HVT DP_OP_26J6_124_4249_U409 ( .A1(n1270), .A2(ori_data_25_), .Y(
        DP_OP_26J6_124_4249_n387) );
  NOR2X0_HVT DP_OP_26J6_124_4249_U21 ( .A1(DP_OP_26J6_124_4249_n43), .A2(
        DP_OP_26J6_124_4249_n83), .Y(DP_OP_26J6_124_4249_n41) );
  AOI22X1_HVT U3 ( .A1(DP_OP_26J6_124_4249_n64), .A2(1'b1), .A3(
        DP_OP_26J6_124_4249_n86), .A4(DP_OP_26J6_124_4249_n63), .Y(n29) );
  OA221X1_HVT U4 ( .A1(1'b0), .A2(DP_OP_26J6_124_4249_n535), .A3(
        DP_OP_26J6_124_4249_n530), .A4(n95), .A5(n97), .Y(
        DP_OP_26J6_124_4249_n527) );
  OA221X1_HVT U5 ( .A1(1'b0), .A2(DP_OP_26J6_124_4249_n355), .A3(
        DP_OP_26J6_124_4249_n366), .A4(DP_OP_26J6_124_4249_n354), .A5(n510), 
        .Y(n520) );
  AOI21X1_HVT U6 ( .A1(n139), .A2(DP_OP_26J6_124_4249_n537), .A3(
        DP_OP_26J6_124_4249_n538), .Y(DP_OP_26J6_124_4249_n536) );
  NAND2X1_HVT U7 ( .A1(n110), .A2(n109), .Y(n139) );
  NAND3X2_HVT U8 ( .A1(n430), .A2(n440), .A3(n450), .Y(n188) );
  NBUFFX2_HVT U9 ( .A(DP_OP_26J6_124_4249_n213), .Y(n1) );
  NAND2X0_HVT U10 ( .A1(n2), .A2(DP_OP_26J6_124_4249_n192), .Y(
        DP_OP_26J6_124_4249_n190) );
  NAND2X0_HVT U11 ( .A1(DP_OP_26J6_124_4249_n213), .A2(n3), .Y(n2) );
  INVX2_HVT U12 ( .A(DP_OP_26J6_124_4249_n191), .Y(n3) );
  NAND2X0_HVT U13 ( .A1(n4), .A2(DP_OP_26J6_124_4249_n211), .Y(
        DP_OP_26J6_124_4249_n201) );
  NAND2X0_HVT U14 ( .A1(n1), .A2(n5), .Y(n4) );
  INVX2_HVT U15 ( .A(DP_OP_26J6_124_4249_n210), .Y(n5) );
  NAND2X0_HVT U16 ( .A1(n6), .A2(DP_OP_26J6_124_4249_n181), .Y(
        DP_OP_26J6_124_4249_n179) );
  NAND2X0_HVT U17 ( .A1(n1), .A2(n7), .Y(n6) );
  INVX2_HVT U18 ( .A(DP_OP_26J6_124_4249_n180), .Y(n7) );
  NAND2X0_HVT U19 ( .A1(n9), .A2(DP_OP_26J6_124_4249_n170), .Y(
        DP_OP_26J6_124_4249_n168) );
  NAND2X0_HVT U20 ( .A1(n1), .A2(n10), .Y(n9) );
  INVX2_HVT U21 ( .A(DP_OP_26J6_124_4249_n169), .Y(n10) );
  XNOR2X2_HVT U22 ( .A1(n1), .A2(DP_OP_26J6_124_4249_n19), .Y(N114) );
  NAND2X0_HVT U23 ( .A1(DP_OP_26J6_124_4249_n148), .A2(n11), .Y(
        DP_OP_26J6_124_4249_n146) );
  NAND2X0_HVT U24 ( .A1(n1), .A2(n12), .Y(n11) );
  INVX2_HVT U25 ( .A(DP_OP_26J6_124_4249_n147), .Y(n12) );
  NAND2X0_HVT U26 ( .A1(DP_OP_26J6_124_4249_n159), .A2(n14), .Y(
        DP_OP_26J6_124_4249_n157) );
  NAND2X0_HVT U27 ( .A1(n1), .A2(n15), .Y(n14) );
  INVX2_HVT U28 ( .A(DP_OP_26J6_124_4249_n158), .Y(n15) );
  NAND2X0_HVT U29 ( .A1(DP_OP_26J6_124_4249_n137), .A2(n16), .Y(
        DP_OP_26J6_124_4249_n135) );
  NAND2X0_HVT U30 ( .A1(n1), .A2(n17), .Y(n16) );
  INVX2_HVT U31 ( .A(DP_OP_26J6_124_4249_n136), .Y(n17) );
  OR3X1_HVT U32 ( .A1(n26), .A2(n24), .A3(n18), .Y(n41) );
  NAND3X0_HVT U33 ( .A1(n22), .A2(n20), .A3(n19), .Y(n18) );
  INVX2_HVT U34 ( .A(N51), .Y(n19) );
  NOR2X0_HVT U35 ( .A1(N49), .A2(N50), .Y(n20) );
  XNOR2X2_HVT U36 ( .A1(DP_OP_26J6_124_4249_n442), .A2(
        DP_OP_26J6_124_4249_n306), .Y(N50) );
  XOR2X2_HVT U37 ( .A1(n21), .A2(DP_OP_26J6_124_4249_n307), .Y(N49) );
  OA21X1_HVT U38 ( .A1(DP_OP_26J6_124_4249_n454), .A2(DP_OP_26J6_124_4249_n519), .A3(DP_OP_26J6_124_4249_n455), .Y(n21) );
  INVX2_HVT U39 ( .A(N56), .Y(n22) );
  XOR2X2_HVT U40 ( .A1(n23), .A2(DP_OP_26J6_124_4249_n300), .Y(N56) );
  OA21X1_HVT U41 ( .A1(DP_OP_26J6_124_4249_n379), .A2(n134), .A3(
        DP_OP_26J6_124_4249_n380), .Y(n23) );
  AND2X1_HVT U42 ( .A1(n108), .A2(n100), .Y(n134) );
  OR3X1_HVT U43 ( .A1(N46), .A2(N47), .A3(n25), .Y(n24) );
  OR3X1_HVT U44 ( .A1(N43), .A2(n185), .A3(N48), .Y(n25) );
  XNOR2X2_HVT U45 ( .A1(DP_OP_26J6_124_4249_n464), .A2(
        DP_OP_26J6_124_4249_n308), .Y(N48) );
  XNOR2X2_HVT U46 ( .A1(DP_OP_26J6_124_4249_n475), .A2(
        DP_OP_26J6_124_4249_n309), .Y(N47) );
  XOR2X2_HVT U47 ( .A1(n137), .A2(DP_OP_26J6_124_4249_n310), .Y(N46) );
  OR2X1_HVT U48 ( .A1(N44), .A2(N45), .Y(n26) );
  INVX2_HVT U49 ( .A(DP_OP_26J6_124_4249_n520), .Y(DP_OP_26J6_124_4249_n519)
         );
  NAND2X0_HVT U50 ( .A1(n27), .A2(DP_OP_26J6_124_4249_n466), .Y(
        DP_OP_26J6_124_4249_n464) );
  NAND2X0_HVT U51 ( .A1(n28), .A2(DP_OP_26J6_124_4249_n520), .Y(n27) );
  AO21X1_HVT U52 ( .A1(n1310), .A2(n139), .A3(n132), .Y(
        DP_OP_26J6_124_4249_n520) );
  INVX2_HVT U53 ( .A(DP_OP_26J6_124_4249_n465), .Y(n28) );
  INVX2_HVT U54 ( .A(n1150), .Y(DP_OP_26J6_124_4249_n1) );
  NAND2X0_HVT U55 ( .A1(n30), .A2(n29), .Y(n92) );
  NAND2X0_HVT U56 ( .A1(n1150), .A2(n31), .Y(n30) );
  INVX2_HVT U57 ( .A(n32), .Y(n31) );
  NAND2X0_HVT U58 ( .A1(DP_OP_26J6_124_4249_n85), .A2(DP_OP_26J6_124_4249_n63), 
        .Y(n32) );
  OR2X2_HVT U59 ( .A1(DP_OP_26J6_124_4249_n129), .A2(DP_OP_26J6_124_4249_n170), 
        .Y(n33) );
  NAND2X0_HVT U60 ( .A1(n33), .A2(DP_OP_26J6_124_4249_n130), .Y(
        DP_OP_26J6_124_4249_n128) );
  OAI21X2_HVT U61 ( .A1(DP_OP_26J6_124_4249_n167), .A2(
        DP_OP_26J6_124_4249_n155), .A3(DP_OP_26J6_124_4249_n156), .Y(
        DP_OP_26J6_124_4249_n150) );
  OR2X1_HVT U62 ( .A1(n34), .A2(n92), .Y(n36) );
  IBUFFX32_HVT U63 ( .A(n93), .Y(n34) );
  NAND2X0_HVT U64 ( .A1(n35), .A2(n92), .Y(n37) );
  NAND2X0_HVT U65 ( .A1(n36), .A2(n37), .Y(N128) );
  INVX1_HVT U66 ( .A(n93), .Y(n35) );
  OR2X4_HVT U67 ( .A1(DP_OP_26J6_124_4249_n177), .A2(DP_OP_26J6_124_4249_n189), 
        .Y(n38) );
  AND3X1_HVT U68 ( .A1(DP_OP_26J6_124_4249_n178), .A2(n38), .A3(n82), .Y(
        DP_OP_26J6_124_4249_n170) );
  AOI21X2_HVT U69 ( .A1(DP_OP_26J6_124_4249_n194), .A2(
        DP_OP_26J6_124_4249_n283), .A3(DP_OP_26J6_124_4249_n183), .Y(
        DP_OP_26J6_124_4249_n181) );
  INVX1_HVT U70 ( .A(n187), .Y(n39) );
  INVX2_HVT U71 ( .A(n39), .Y(n40) );
  INVX1_HVT U72 ( .A(n100), .Y(DP_OP_26J6_124_4249_n435) );
  INVX1_HVT U73 ( .A(n1210), .Y(DP_OP_26J6_124_4249_n571) );
  OR3X1_HVT U74 ( .A1(n149), .A2(n155), .A3(n41), .Y(n42) );
  OR3X1_HVT U75 ( .A1(n150), .A2(n154), .A3(n42), .Y(n430) );
  INVX0_HVT U76 ( .A(n_quantized_data[7]), .Y(n440) );
  OR3X1_HVT U77 ( .A1(n165), .A2(n164), .A3(n163), .Y(n450) );
  NAND2X0_HVT U78 ( .A1(bias_data[3]), .A2(ori_data_30_), .Y(n460) );
  AND2X1_HVT U79 ( .A1(n460), .A2(n144), .Y(n470) );
  INVX0_HVT U80 ( .A(DP_OP_26J6_124_4249_n1), .Y(n480) );
  AO21X1_HVT U81 ( .A1(DP_OP_26J6_124_4249_n41), .A2(n480), .A3(
        DP_OP_26J6_124_4249_n42), .Y(n490) );
  HADDX1_HVT U82 ( .A0(n470), .B0(n490), .SO(N130) );
  NAND2X0_HVT U84 ( .A1(DP_OP_26J6_124_4249_n352), .A2(
        DP_OP_26J6_124_4249_n371), .Y(n510) );
  OAI21X2_HVT U85 ( .A1(DP_OP_26J6_124_4249_n350), .A2(
        DP_OP_26J6_124_4249_n391), .A3(n520), .Y(DP_OP_26J6_124_4249_n349) );
  INVX0_HVT U86 ( .A(mode[0]), .Y(n530) );
  AND2X1_HVT U87 ( .A1(mode[1]), .A2(n530), .Y(n184) );
  HADDX1_HVT U88 ( .A0(DP_OP_26J6_124_4249_n320), .B0(DP_OP_26J6_124_4249_n571), .SO(n540) );
  NAND4X0_HVT U89 ( .A1(n184), .A2(n99), .A3(n153), .A4(n540), .Y(n550) );
  INVX0_HVT U90 ( .A(DP_OP_26J6_124_4249_n265), .Y(n560) );
  HADDX1_HVT U91 ( .A0(ori_data_5_), .B0(n560), .SO(n570) );
  NAND4X0_HVT U92 ( .A1(n1300), .A2(n40), .A3(n185), .A4(n570), .Y(n580) );
  NAND3X0_HVT U93 ( .A1(n188), .A2(n550), .A3(n580), .Y(n_quantized_data[0])
         );
  HADDX1_HVT U94 ( .A0(DP_OP_26J6_124_4249_n567), .B0(DP_OP_26J6_124_4249_n319), .SO(n590) );
  NAND4X0_HVT U95 ( .A1(n184), .A2(n99), .A3(n153), .A4(n590), .Y(n600) );
  HADDX1_HVT U96 ( .A0(DP_OP_26J6_124_4249_n263), .B0(DP_OP_26J6_124_4249_n262), .SO(n610) );
  NAND4X0_HVT U97 ( .A1(n40), .A2(n1300), .A3(n185), .A4(n610), .Y(n62) );
  NAND3X0_HVT U98 ( .A1(n188), .A2(n600), .A3(n62), .Y(n_quantized_data[1]) );
  XNOR2X1_HVT U99 ( .A1(DP_OP_26J6_124_4249_n560), .A2(
        DP_OP_26J6_124_4249_n318), .Y(n63) );
  NAND4X0_HVT U100 ( .A1(n99), .A2(n184), .A3(n153), .A4(n63), .Y(n64) );
  HADDX1_HVT U101 ( .A0(DP_OP_26J6_124_4249_n260), .B0(DP_OP_26J6_124_4249_n25), .SO(n65) );
  NAND4X0_HVT U102 ( .A1(n40), .A2(n186), .A3(n185), .A4(n65), .Y(n66) );
  NAND3X0_HVT U103 ( .A1(n188), .A2(n64), .A3(n66), .Y(n_quantized_data[2]) );
  INVX0_HVT U104 ( .A(n139), .Y(n67) );
  HADDX1_HVT U105 ( .A0(DP_OP_26J6_124_4249_n317), .B0(n67), .SO(n68) );
  NAND4X0_HVT U106 ( .A1(n99), .A2(n184), .A3(n153), .A4(n68), .Y(n69) );
  XNOR2X1_HVT U107 ( .A1(DP_OP_26J6_124_4249_n253), .A2(
        DP_OP_26J6_124_4249_n24), .Y(n70) );
  NAND4X0_HVT U108 ( .A1(n1300), .A2(n40), .A3(n185), .A4(n70), .Y(n71) );
  NAND3X0_HVT U109 ( .A1(n188), .A2(n69), .A3(n71), .Y(n_quantized_data[3]) );
  HADDX1_HVT U110 ( .A0(DP_OP_26J6_124_4249_n545), .B0(
        DP_OP_26J6_124_4249_n316), .SO(n72) );
  NAND4X0_HVT U111 ( .A1(n184), .A2(n99), .A3(n153), .A4(n72), .Y(n73) );
  INVX0_HVT U112 ( .A(DP_OP_26J6_124_4249_n247), .Y(n74) );
  HADDX1_HVT U113 ( .A0(DP_OP_26J6_124_4249_n23), .B0(n74), .SO(n75) );
  NAND4X0_HVT U114 ( .A1(n186), .A2(n40), .A3(n185), .A4(n75), .Y(n76) );
  NAND3X0_HVT U115 ( .A1(n188), .A2(n73), .A3(n76), .Y(n_quantized_data[4]) );
  INVX0_HVT U116 ( .A(n104), .Y(n77) );
  NAND2X0_HVT U117 ( .A1(DP_OP_26J6_124_4249_n456), .A2(n77), .Y(
        DP_OP_26J6_124_4249_n436) );
  HADDX1_HVT U118 ( .A0(DP_OP_26J6_124_4249_n536), .B0(
        DP_OP_26J6_124_4249_n315), .SO(n78) );
  NAND4X0_HVT U119 ( .A1(n184), .A2(n99), .A3(n153), .A4(n78), .Y(n79) );
  HADDX1_HVT U120 ( .A0(DP_OP_26J6_124_4249_n238), .B0(DP_OP_26J6_124_4249_n22), .SO(n80) );
  NAND4X0_HVT U121 ( .A1(n40), .A2(n1300), .A3(n185), .A4(n80), .Y(n81) );
  NAND3X0_HVT U122 ( .A1(n188), .A2(n79), .A3(n81), .Y(n_quantized_data[5]) );
  NAND2X0_HVT U123 ( .A1(DP_OP_26J6_124_4249_n175), .A2(
        DP_OP_26J6_124_4249_n194), .Y(n82) );
  INVX0_HVT U124 ( .A(n106), .Y(n83) );
  NAND2X0_HVT U125 ( .A1(DP_OP_26J6_124_4249_n500), .A2(n83), .Y(
        DP_OP_26J6_124_4249_n476) );
  INVX0_HVT U126 ( .A(n1180), .Y(n84) );
  OAI21X1_HVT U127 ( .A1(DP_OP_26J6_124_4249_n567), .A2(n84), .A3(
        DP_OP_26J6_124_4249_n566), .Y(DP_OP_26J6_124_4249_n560) );
  NAND2X0_HVT U128 ( .A1(n139), .A2(DP_OP_26J6_124_4249_n594), .Y(n85) );
  AND2X1_HVT U129 ( .A1(n85), .A2(DP_OP_26J6_124_4249_n553), .Y(
        DP_OP_26J6_124_4249_n545) );
  HADDX1_HVT U130 ( .A0(DP_OP_26J6_124_4249_n527), .B0(
        DP_OP_26J6_124_4249_n314), .SO(n86) );
  NAND4X0_HVT U131 ( .A1(n184), .A2(n99), .A3(n153), .A4(n86), .Y(n87) );
  HADDX1_HVT U132 ( .A0(DP_OP_26J6_124_4249_n229), .B0(DP_OP_26J6_124_4249_n21), .SO(n88) );
  NAND4X0_HVT U133 ( .A1(n40), .A2(n186), .A3(n185), .A4(n88), .Y(n89) );
  NAND3X0_HVT U134 ( .A1(n188), .A2(n87), .A3(n89), .Y(n_quantized_data[6]) );
  NAND2X0_HVT U135 ( .A1(DP_OP_26J6_124_4249_n582), .A2(
        DP_OP_26J6_124_4249_n432), .Y(n90) );
  HADDX1_HVT U136 ( .A0(n135), .B0(n90), .SO(N51) );
  AND2X1_HVT U138 ( .A1(DP_OP_26J6_124_4249_n271), .A2(DP_OP_26J6_124_4249_n59), .Y(n93) );
  NAND2X0_HVT U139 ( .A1(DP_OP_26J6_124_4249_n247), .A2(
        DP_OP_26J6_124_4249_n289), .Y(n94) );
  AND2X1_HVT U140 ( .A1(n94), .A2(DP_OP_26J6_124_4249_n246), .Y(
        DP_OP_26J6_124_4249_n238) );
  INVX0_HVT U141 ( .A(DP_OP_26J6_124_4249_n538), .Y(n95) );
  INVX0_HVT U142 ( .A(DP_OP_26J6_124_4249_n530), .Y(n96) );
  NAND3X0_HVT U143 ( .A1(n139), .A2(DP_OP_26J6_124_4249_n537), .A3(n96), .Y(
        n97) );
  AO22X1_HVT U145 ( .A1(n184), .A2(N61), .A3(n185), .A4(N131), .Y(
        n_quantized_data[7]) );
  NAND2X0_HVT U146 ( .A1(n171), .A2(N61), .Y(n99) );
  OAI21X2_HVT U147 ( .A1(DP_OP_26J6_124_4249_n211), .A2(
        DP_OP_26J6_124_4249_n199), .A3(DP_OP_26J6_124_4249_n200), .Y(
        DP_OP_26J6_124_4249_n194) );
  INVX1_HVT U148 ( .A(n103), .Y(DP_OP_26J6_124_4249_n457) );
  INVX1_HVT U149 ( .A(n107), .Y(DP_OP_26J6_124_4249_n501) );
  INVX1_HVT U150 ( .A(n1170), .Y(DP_OP_26J6_124_4249_n558) );
  NOR2X4_HVT U151 ( .A1(n1230), .A2(ori_data_15_), .Y(DP_OP_26J6_124_4249_n495) );
  OA21X1_HVT U152 ( .A1(DP_OP_26J6_124_4249_n436), .A2(
        DP_OP_26J6_124_4249_n477), .A3(n101), .Y(n100) );
  OA21X1_HVT U153 ( .A1(n104), .A2(n103), .A3(n102), .Y(n101) );
  OA21X1_HVT U154 ( .A1(DP_OP_26J6_124_4249_n452), .A2(
        DP_OP_26J6_124_4249_n440), .A3(DP_OP_26J6_124_4249_n441), .Y(n102) );
  OA21X1_HVT U155 ( .A1(DP_OP_26J6_124_4249_n474), .A2(
        DP_OP_26J6_124_4249_n462), .A3(DP_OP_26J6_124_4249_n463), .Y(n103) );
  OR2X1_HVT U156 ( .A1(DP_OP_26J6_124_4249_n447), .A2(DP_OP_26J6_124_4249_n440), .Y(n104) );
  OA21X1_HVT U157 ( .A1(n107), .A2(n106), .A3(n105), .Y(
        DP_OP_26J6_124_4249_n477) );
  OA21X1_HVT U158 ( .A1(DP_OP_26J6_124_4249_n496), .A2(
        DP_OP_26J6_124_4249_n484), .A3(DP_OP_26J6_124_4249_n485), .Y(n105) );
  OR2X1_HVT U159 ( .A1(DP_OP_26J6_124_4249_n495), .A2(DP_OP_26J6_124_4249_n484), .Y(n106) );
  OA21X1_HVT U160 ( .A1(DP_OP_26J6_124_4249_n518), .A2(
        DP_OP_26J6_124_4249_n506), .A3(DP_OP_26J6_124_4249_n507), .Y(n107) );
  NAND2X0_HVT U161 ( .A1(DP_OP_26J6_124_4249_n520), .A2(
        DP_OP_26J6_124_4249_n434), .Y(n108) );
  OA21X1_HVT U162 ( .A1(DP_OP_26J6_124_4249_n566), .A2(
        DP_OP_26J6_124_4249_n558), .A3(DP_OP_26J6_124_4249_n559), .Y(n109) );
  NAND2X0_HVT U163 ( .A1(n1160), .A2(DP_OP_26J6_124_4249_n568), .Y(n110) );
  OR2X1_HVT U164 ( .A1(N124), .A2(N123), .Y(n156) );
  XNOR2X2_HVT U165 ( .A1(n111), .A2(DP_OP_26J6_124_4249_n10), .Y(N123) );
  NAND2X0_HVT U166 ( .A1(n112), .A2(DP_OP_26J6_124_4249_n125), .Y(n111) );
  NAND2X0_HVT U167 ( .A1(n1150), .A2(DP_OP_26J6_124_4249_n277), .Y(n112) );
  XNOR2X2_HVT U168 ( .A1(n1130), .A2(DP_OP_26J6_124_4249_n9), .Y(N124) );
  NAND2X0_HVT U169 ( .A1(n1140), .A2(DP_OP_26J6_124_4249_n106), .Y(n1130) );
  NAND2X0_HVT U170 ( .A1(n1150), .A2(DP_OP_26J6_124_4249_n107), .Y(n1140) );
  AO21X1_HVT U171 ( .A1(DP_OP_26J6_124_4249_n213), .A2(
        DP_OP_26J6_124_4249_n127), .A3(DP_OP_26J6_124_4249_n128), .Y(n1150) );
  NAND2X0_HVT U172 ( .A1(ori_data_7_), .A2(bias_data[2]), .Y(
        DP_OP_26J6_124_4249_n566) );
  AND2X1_HVT U173 ( .A1(n1180), .A2(n1170), .Y(n1160) );
  OR2X1_HVT U174 ( .A1(n1270), .A2(ori_data_8_), .Y(n1170) );
  OR2X1_HVT U175 ( .A1(bias_data[2]), .A2(ori_data_7_), .Y(n1180) );
  NAND2X0_HVT U176 ( .A1(n1190), .A2(DP_OP_26J6_124_4249_n570), .Y(
        DP_OP_26J6_124_4249_n568) );
  NAND2X0_HVT U177 ( .A1(n1210), .A2(n1200), .Y(n1190) );
  OR2X1_HVT U178 ( .A1(bias_data[1]), .A2(ori_data_6_), .Y(n1200) );
  OR2X1_HVT U179 ( .A1(bias_data[0]), .A2(ori_data_5_), .Y(n1210) );
  XNOR2X2_HVT U180 ( .A1(DP_OP_26J6_124_4249_n201), .A2(
        DP_OP_26J6_124_4249_n18), .Y(N115) );
  XNOR2X2_HVT U181 ( .A1(DP_OP_26J6_124_4249_n146), .A2(
        DP_OP_26J6_124_4249_n13), .Y(N120) );
  OAI21X2_HVT U182 ( .A1(DP_OP_26J6_124_4249_n259), .A2(
        DP_OP_26J6_124_4249_n251), .A3(DP_OP_26J6_124_4249_n252), .Y(
        DP_OP_26J6_124_4249_n250) );
  XOR2X2_HVT U183 ( .A1(n1220), .A2(DP_OP_26J6_124_4249_n302), .Y(N54) );
  OA21X2_HVT U184 ( .A1(DP_OP_26J6_124_4249_n401), .A2(n134), .A3(
        DP_OP_26J6_124_4249_n402), .Y(n1220) );
  XOR2X2_HVT U185 ( .A1(n1290), .A2(DP_OP_26J6_124_4249_n296), .Y(N60) );
  IBUFFX2_HVT U186 ( .A(DP_OP_26J6_124_4249_n568), .Y(DP_OP_26J6_124_4249_n567) );
  AOI21X2_HVT U187 ( .A1(DP_OP_26J6_124_4249_n520), .A2(
        DP_OP_26J6_124_4249_n434), .A3(DP_OP_26J6_124_4249_n435), .Y(n135) );
  OA21X2_HVT U188 ( .A1(DP_OP_26J6_124_4249_n487), .A2(
        DP_OP_26J6_124_4249_n519), .A3(DP_OP_26J6_124_4249_n488), .Y(n137) );
  OAI21X2_HVT U189 ( .A1(DP_OP_26J6_124_4249_n357), .A2(n134), .A3(
        DP_OP_26J6_124_4249_n358), .Y(DP_OP_26J6_124_4249_n356) );
  OAI21X2_HVT U190 ( .A1(DP_OP_26J6_124_4249_n368), .A2(n134), .A3(
        DP_OP_26J6_124_4249_n369), .Y(DP_OP_26J6_124_4249_n367) );
  OAI21X2_HVT U191 ( .A1(DP_OP_26J6_124_4249_n346), .A2(n134), .A3(
        DP_OP_26J6_124_4249_n347), .Y(DP_OP_26J6_124_4249_n345) );
  OAI21X2_HVT U192 ( .A1(DP_OP_26J6_124_4249_n390), .A2(n134), .A3(
        DP_OP_26J6_124_4249_n391), .Y(DP_OP_26J6_124_4249_n389) );
  OAI21X2_HVT U193 ( .A1(DP_OP_26J6_124_4249_n498), .A2(
        DP_OP_26J6_124_4249_n519), .A3(n107), .Y(DP_OP_26J6_124_4249_n497) );
  OAI21X2_HVT U194 ( .A1(DP_OP_26J6_124_4249_n517), .A2(
        DP_OP_26J6_124_4249_n519), .A3(DP_OP_26J6_124_4249_n518), .Y(
        DP_OP_26J6_124_4249_n508) );
  INVX0_HVT U195 ( .A(DP_OP_26J6_124_4249_n166), .Y(DP_OP_26J6_124_4249_n281)
         );
  NOR2X0_HVT U196 ( .A1(bias_data[3]), .A2(ori_data_19_), .Y(
        DP_OP_26J6_124_4249_n447) );
  OR2X1_HVT U197 ( .A1(n152), .A2(n151), .Y(n153) );
  INVX0_HVT U198 ( .A(N61), .Y(n151) );
  XOR2X1_HVT U199 ( .A1(n140), .A2(DP_OP_26J6_124_4249_n304), .Y(N52) );
  INVX0_HVT U200 ( .A(DP_OP_26J6_124_4249_n349), .Y(DP_OP_26J6_124_4249_n347)
         );
  OAI21X1_HVT U201 ( .A1(DP_OP_26J6_124_4249_n412), .A2(n135), .A3(
        DP_OP_26J6_124_4249_n413), .Y(DP_OP_26J6_124_4249_n411) );
  INVX0_HVT U202 ( .A(DP_OP_26J6_124_4249_n348), .Y(DP_OP_26J6_124_4249_n346)
         );
  INVX0_HVT U203 ( .A(DP_OP_26J6_124_4249_n83), .Y(DP_OP_26J6_124_4249_n85) );
  INVX0_HVT U204 ( .A(DP_OP_26J6_124_4249_n108), .Y(DP_OP_26J6_124_4249_n106)
         );
  AOI21X1_HVT U205 ( .A1(DP_OP_26J6_124_4249_n172), .A2(
        DP_OP_26J6_124_4249_n149), .A3(DP_OP_26J6_124_4249_n150), .Y(
        DP_OP_26J6_124_4249_n148) );
  INVX0_HVT U206 ( .A(DP_OP_26J6_124_4249_n390), .Y(DP_OP_26J6_124_4249_n392)
         );
  INVX0_HVT U207 ( .A(DP_OP_26J6_124_4249_n63), .Y(DP_OP_26J6_124_4249_n65) );
  INVX0_HVT U208 ( .A(DP_OP_26J6_124_4249_n476), .Y(DP_OP_26J6_124_4249_n478)
         );
  INVX0_HVT U209 ( .A(DP_OP_26J6_124_4249_n64), .Y(DP_OP_26J6_124_4249_n66) );
  INVX0_HVT U210 ( .A(DP_OP_26J6_124_4249_n477), .Y(DP_OP_26J6_124_4249_n479)
         );
  INVX0_HVT U211 ( .A(DP_OP_26J6_124_4249_n169), .Y(DP_OP_26J6_124_4249_n171)
         );
  INVX0_HVT U212 ( .A(DP_OP_26J6_124_4249_n170), .Y(DP_OP_26J6_124_4249_n172)
         );
  INVX0_HVT U213 ( .A(DP_OP_26J6_124_4249_n410), .Y(DP_OP_26J6_124_4249_n404)
         );
  INVX0_HVT U214 ( .A(DP_OP_26J6_124_4249_n500), .Y(DP_OP_26J6_124_4249_n498)
         );
  INVX0_HVT U215 ( .A(DP_OP_26J6_124_4249_n361), .Y(DP_OP_26J6_124_4249_n576)
         );
  OAI21X1_HVT U216 ( .A1(DP_OP_26J6_124_4249_n410), .A2(
        DP_OP_26J6_124_4249_n398), .A3(DP_OP_26J6_124_4249_n399), .Y(
        DP_OP_26J6_124_4249_n397) );
  INVX0_HVT U217 ( .A(DP_OP_26J6_124_4249_n54), .Y(DP_OP_26J6_124_4249_n271)
         );
  INVX0_HVT U218 ( .A(DP_OP_26J6_124_4249_n149), .Y(DP_OP_26J6_124_4249_n151)
         );
  INVX0_HVT U219 ( .A(DP_OP_26J6_124_4249_n456), .Y(DP_OP_26J6_124_4249_n458)
         );
  INVX0_HVT U220 ( .A(DP_OP_26J6_124_4249_n415), .Y(DP_OP_26J6_124_4249_n413)
         );
  INVX0_HVT U221 ( .A(DP_OP_26J6_124_4249_n231), .Y(DP_OP_26J6_124_4249_n233)
         );
  INVX0_HVT U222 ( .A(DP_OP_26J6_124_4249_n150), .Y(DP_OP_26J6_124_4249_n152)
         );
  INVX0_HVT U223 ( .A(DP_OP_26J6_124_4249_n414), .Y(DP_OP_26J6_124_4249_n412)
         );
  INVX0_HVT U224 ( .A(DP_OP_26J6_124_4249_n230), .Y(DP_OP_26J6_124_4249_n232)
         );
  INVX0_HVT U225 ( .A(DP_OP_26J6_124_4249_n447), .Y(DP_OP_26J6_124_4249_n584)
         );
  INVX0_HVT U226 ( .A(DP_OP_26J6_124_4249_n124), .Y(DP_OP_26J6_124_4249_n277)
         );
  INVX0_HVT U227 ( .A(DP_OP_26J6_124_4249_n370), .Y(DP_OP_26J6_124_4249_n372)
         );
  INVX0_HVT U228 ( .A(DP_OP_26J6_124_4249_n371), .Y(DP_OP_26J6_124_4249_n373)
         );
  INVX0_HVT U229 ( .A(DP_OP_26J6_124_4249_n258), .Y(DP_OP_26J6_124_4249_n291)
         );
  INVX0_HVT U230 ( .A(DP_OP_26J6_124_4249_n194), .Y(DP_OP_26J6_124_4249_n192)
         );
  INVX0_HVT U231 ( .A(DP_OP_26J6_124_4249_n188), .Y(DP_OP_26J6_124_4249_n283)
         );
  INVX0_HVT U232 ( .A(DP_OP_26J6_124_4249_n167), .Y(DP_OP_26J6_124_4249_n161)
         );
  INVX0_HVT U233 ( .A(DP_OP_26J6_124_4249_n189), .Y(DP_OP_26J6_124_4249_n183)
         );
  INVX0_HVT U234 ( .A(DP_OP_26J6_124_4249_n474), .Y(DP_OP_26J6_124_4249_n468)
         );
  INVX0_HVT U235 ( .A(DP_OP_26J6_124_4249_n473), .Y(DP_OP_26J6_124_4249_n586)
         );
  INVX0_HVT U236 ( .A(DP_OP_26J6_124_4249_n530), .Y(DP_OP_26J6_124_4249_n592)
         );
  INVX0_HVT U237 ( .A(DP_OP_26J6_124_4249_n193), .Y(DP_OP_26J6_124_4249_n191)
         );
  INVX0_HVT U238 ( .A(DP_OP_26J6_124_4249_n517), .Y(DP_OP_26J6_124_4249_n590)
         );
  INVX0_HVT U239 ( .A(DP_OP_26J6_124_4249_n543), .Y(DP_OP_26J6_124_4249_n593)
         );
  INVX0_HVT U240 ( .A(DP_OP_26J6_124_4249_n431), .Y(DP_OP_26J6_124_4249_n582)
         );
  INVX0_HVT U241 ( .A(DP_OP_26J6_124_4249_n388), .Y(DP_OP_26J6_124_4249_n382)
         );
  INVX0_HVT U242 ( .A(DP_OP_26J6_124_4249_n251), .Y(DP_OP_26J6_124_4249_n290)
         );
  INVX0_HVT U243 ( .A(DP_OP_26J6_124_4249_n495), .Y(DP_OP_26J6_124_4249_n588)
         );
  INVX0_HVT U244 ( .A(DP_OP_26J6_124_4249_n496), .Y(DP_OP_26J6_124_4249_n490)
         );
  INVX0_HVT U245 ( .A(DP_OP_26J6_124_4249_n140), .Y(DP_OP_26J6_124_4249_n279)
         );
  NOR2X0_HVT U246 ( .A1(n1270), .A2(ori_data_17_), .Y(DP_OP_26J6_124_4249_n473) );
  INVX0_HVT U247 ( .A(DP_OP_26J6_124_4249_n210), .Y(DP_OP_26J6_124_4249_n285)
         );
  INVX0_HVT U248 ( .A(DP_OP_26J6_124_4249_n223), .Y(DP_OP_26J6_124_4249_n287)
         );
  INVX0_HVT U249 ( .A(DP_OP_26J6_124_4249_n103), .Y(DP_OP_26J6_124_4249_n97)
         );
  INVX0_HVT U250 ( .A(DP_OP_26J6_124_4249_n344), .Y(DP_OP_26J6_124_4249_n342)
         );
  INVX0_HVT U251 ( .A(DP_OP_26J6_124_4249_n333), .Y(DP_OP_26J6_124_4249_n331)
         );
  INVX0_HVT U252 ( .A(DP_OP_26J6_124_4249_n81), .Y(DP_OP_26J6_124_4249_n75) );
  INVX0_HVT U253 ( .A(ori_data_6_), .Y(DP_OP_26J6_124_4249_n265) );
  INVX1_HVT U254 ( .A(n133), .Y(n1260) );
  INVX1_HVT U255 ( .A(n133), .Y(n1270) );
  INVX1_HVT U256 ( .A(n133), .Y(n1280) );
  INVX1_HVT U257 ( .A(n133), .Y(n1250) );
  INVX1_HVT U258 ( .A(n133), .Y(n1230) );
  INVX1_HVT U259 ( .A(n133), .Y(n1240) );
  INVX1_HVT U260 ( .A(bias_data[3]), .Y(n133) );
  INVX0_HVT U261 ( .A(srstn), .Y(n13) );
  OAI21X2_HVT U262 ( .A1(DP_OP_26J6_124_4249_n1), .A2(DP_OP_26J6_124_4249_n32), 
        .A3(DP_OP_26J6_124_4249_n33), .Y(DP_OP_26J6_124_4249_n31) );
  OA21X1_HVT U263 ( .A1(DP_OP_26J6_124_4249_n335), .A2(n135), .A3(
        DP_OP_26J6_124_4249_n336), .Y(n1290) );
  NAND2X0_HVT U264 ( .A1(n183), .A2(N131), .Y(n1300) );
  AND2X1_HVT U265 ( .A1(DP_OP_26J6_124_4249_n537), .A2(
        DP_OP_26J6_124_4249_n523), .Y(n1310) );
  AO21X1_HVT U266 ( .A1(DP_OP_26J6_124_4249_n538), .A2(
        DP_OP_26J6_124_4249_n523), .A3(DP_OP_26J6_124_4249_n524), .Y(n132) );
  INVX1_HVT U267 ( .A(DP_OP_26J6_124_4249_n245), .Y(DP_OP_26J6_124_4249_n289)
         );
  INVX1_HVT U268 ( .A(DP_OP_26J6_124_4249_n248), .Y(DP_OP_26J6_124_4249_n247)
         );
  INVX1_HVT U269 ( .A(DP_OP_26J6_124_4249_n261), .Y(DP_OP_26J6_124_4249_n260)
         );
  INVX1_HVT U270 ( .A(ori_data_7_), .Y(DP_OP_26J6_124_4249_n262) );
  INVX1_HVT U271 ( .A(DP_OP_26J6_124_4249_n80), .Y(DP_OP_26J6_124_4249_n74) );
  INVX1_HVT U272 ( .A(DP_OP_26J6_124_4249_n102), .Y(DP_OP_26J6_124_4249_n96)
         );
  INVX1_HVT U273 ( .A(DP_OP_26J6_124_4249_n387), .Y(DP_OP_26J6_124_4249_n578)
         );
  INVX1_HVT U274 ( .A(DP_OP_26J6_124_4249_n391), .Y(DP_OP_26J6_124_4249_n393)
         );
  INVX1_HVT U275 ( .A(DP_OP_26J6_124_4249_n409), .Y(DP_OP_26J6_124_4249_n580)
         );
  INVX1_HVT U276 ( .A(DP_OP_26J6_124_4249_n552), .Y(DP_OP_26J6_124_4249_n594)
         );
  INVX1_HVT U277 ( .A(DP_OP_26J6_124_4249_n84), .Y(DP_OP_26J6_124_4249_n86) );
  XOR2X1_HVT U278 ( .A1(DP_OP_26J6_124_4249_n1), .A2(DP_OP_26J6_124_4249_n11), 
        .Y(N122) );
  NAND2X0_HVT U279 ( .A1(n136), .A2(DP_OP_26J6_124_4249_n215), .Y(
        DP_OP_26J6_124_4249_n213) );
  OR2X1_HVT U280 ( .A1(DP_OP_26J6_124_4249_n214), .A2(DP_OP_26J6_124_4249_n248), .Y(n136) );
  AO21X1_HVT U281 ( .A1(n145), .A2(DP_OP_26J6_124_4249_n520), .A3(n138), .Y(
        DP_OP_26J6_124_4249_n442) );
  OR2X1_HVT U282 ( .A1(n1230), .A2(ori_data_31_), .Y(n141) );
  OR2X1_HVT U283 ( .A1(n1270), .A2(ori_data_31_), .Y(n142) );
  AO21X1_HVT U284 ( .A1(n146), .A2(DP_OP_26J6_124_4249_n342), .A3(
        DP_OP_26J6_124_4249_n331), .Y(n143) );
  OR2X1_HVT U285 ( .A1(n1250), .A2(ori_data_30_), .Y(n144) );
  AND2X1_HVT U286 ( .A1(DP_OP_26J6_124_4249_n445), .A2(
        DP_OP_26J6_124_4249_n478), .Y(n145) );
  OR2X1_HVT U287 ( .A1(n1280), .A2(ori_data_30_), .Y(n146) );
  AND2X1_HVT U288 ( .A1(n148), .A2(n146), .Y(n147) );
  OR2X1_HVT U289 ( .A1(n1260), .A2(ori_data_29_), .Y(n148) );
  NOR2X0_HVT U290 ( .A1(n1280), .A2(ori_data_11_), .Y(DP_OP_26J6_124_4249_n530) );
  AOI21X1_HVT U291 ( .A1(DP_OP_26J6_124_4249_n479), .A2(
        DP_OP_26J6_124_4249_n586), .A3(DP_OP_26J6_124_4249_n468), .Y(
        DP_OP_26J6_124_4249_n466) );
  AO21X1_HVT U292 ( .A1(DP_OP_26J6_124_4249_n479), .A2(
        DP_OP_26J6_124_4249_n445), .A3(DP_OP_26J6_124_4249_n446), .Y(n138) );
  OA21X1_HVT U293 ( .A1(DP_OP_26J6_124_4249_n431), .A2(n134), .A3(
        DP_OP_26J6_124_4249_n432), .Y(n140) );
  AOI21X1_HVT U294 ( .A1(DP_OP_26J6_124_4249_n231), .A2(
        DP_OP_26J6_124_4249_n216), .A3(DP_OP_26J6_124_4249_n217), .Y(
        DP_OP_26J6_124_4249_n215) );
  NOR2X0_HVT U295 ( .A1(DP_OP_26J6_124_4249_n155), .A2(
        DP_OP_26J6_124_4249_n166), .Y(DP_OP_26J6_124_4249_n149) );
  AOI21X1_HVT U296 ( .A1(DP_OP_26J6_124_4249_n247), .A2(
        DP_OP_26J6_124_4249_n230), .A3(DP_OP_26J6_124_4249_n231), .Y(
        DP_OP_26J6_124_4249_n229) );
  XOR2X1_HVT U297 ( .A1(DP_OP_26J6_124_4249_n519), .A2(
        DP_OP_26J6_124_4249_n313), .Y(N43) );
  OAI21X1_HVT U298 ( .A1(DP_OP_26J6_124_4249_n50), .A2(DP_OP_26J6_124_4249_n1), 
        .A3(DP_OP_26J6_124_4249_n51), .Y(DP_OP_26J6_124_4249_n49) );
  XNOR2X2_HVT U299 ( .A1(DP_OP_26J6_124_4249_n190), .A2(
        DP_OP_26J6_124_4249_n17), .Y(N116) );
  OAI21X1_HVT U300 ( .A1(DP_OP_26J6_124_4249_n72), .A2(DP_OP_26J6_124_4249_n1), 
        .A3(DP_OP_26J6_124_4249_n73), .Y(DP_OP_26J6_124_4249_n71) );
  OAI21X1_HVT U301 ( .A1(DP_OP_26J6_124_4249_n94), .A2(DP_OP_26J6_124_4249_n1), 
        .A3(DP_OP_26J6_124_4249_n95), .Y(DP_OP_26J6_124_4249_n93) );
  OAI21X1_HVT U302 ( .A1(DP_OP_26J6_124_4249_n83), .A2(DP_OP_26J6_124_4249_n1), 
        .A3(DP_OP_26J6_124_4249_n84), .Y(DP_OP_26J6_124_4249_n82) );
  OAI21X1_HVT U303 ( .A1(DP_OP_26J6_124_4249_n324), .A2(n135), .A3(
        DP_OP_26J6_124_4249_n325), .Y(DP_OP_26J6_124_4249_n323) );
  OAI21X2_HVT U304 ( .A1(DP_OP_26J6_124_4249_n476), .A2(
        DP_OP_26J6_124_4249_n519), .A3(DP_OP_26J6_124_4249_n477), .Y(
        DP_OP_26J6_124_4249_n475) );
  INVX1_HVT U305 ( .A(n184), .Y(n185) );
  OR2X1_HVT U306 ( .A1(N59), .A2(N53), .Y(n149) );
  OR2X1_HVT U307 ( .A1(N60), .A2(N52), .Y(n150) );
  AND3X1_HVT U308 ( .A1(n175), .A2(n174), .A3(N55), .Y(n152) );
  OR2X1_HVT U309 ( .A1(N54), .A2(N58), .Y(n154) );
  OR2X1_HVT U310 ( .A1(N57), .A2(N55), .Y(n155) );
  OR2X1_HVT U311 ( .A1(N130), .A2(N125), .Y(n165) );
  OR3X1_HVT U312 ( .A1(N127), .A2(N126), .A3(n156), .Y(n164) );
  OR2X1_HVT U313 ( .A1(N115), .A2(N120), .Y(n157) );
  OR3X1_HVT U314 ( .A1(N119), .A2(N117), .A3(n157), .Y(n162) );
  OR3X1_HVT U315 ( .A1(n184), .A2(N113), .A3(N114), .Y(n158) );
  OR3X1_HVT U316 ( .A1(N122), .A2(n158), .A3(N116), .Y(n159) );
  OR3X1_HVT U317 ( .A1(N121), .A2(N118), .A3(n159), .Y(n161) );
  OR2X1_HVT U318 ( .A1(N128), .A2(N129), .Y(n160) );
  OR3X1_HVT U319 ( .A1(n162), .A2(n161), .A3(n160), .Y(n163) );
  NAND2X0_HVT U320 ( .A1(N56), .A2(N60), .Y(n170) );
  NAND2X0_HVT U321 ( .A1(N54), .A2(N52), .Y(n169) );
  AND2X1_HVT U322 ( .A1(N47), .A2(N45), .Y(n166) );
  AND3X1_HVT U323 ( .A1(n166), .A2(N49), .A3(N50), .Y(n167) );
  NAND2X0_HVT U324 ( .A1(n167), .A2(N58), .Y(n168) );
  OR3X1_HVT U325 ( .A1(n170), .A2(n169), .A3(n168), .Y(n171) );
  AND2X1_HVT U326 ( .A1(N48), .A2(N46), .Y(n173) );
  AND3X1_HVT U327 ( .A1(N44), .A2(N43), .A3(N51), .Y(n172) );
  AND3X1_HVT U328 ( .A1(N53), .A2(n173), .A3(n172), .Y(n175) );
  AND2X1_HVT U329 ( .A1(N59), .A2(N57), .Y(n174) );
  NAND2X0_HVT U330 ( .A1(N123), .A2(N130), .Y(n178) );
  NAND2X0_HVT U331 ( .A1(N128), .A2(N129), .Y(n177) );
  NAND2X0_HVT U332 ( .A1(N127), .A2(N124), .Y(n176) );
  OR3X1_HVT U333 ( .A1(n178), .A2(n177), .A3(n176), .Y(n179) );
  NAND2X0_HVT U334 ( .A1(n179), .A2(N131), .Y(n187) );
  AND3X1_HVT U335 ( .A1(N122), .A2(N114), .A3(N113), .Y(n180) );
  AND4X1_HVT U336 ( .A1(n180), .A2(N121), .A3(N118), .A4(N116), .Y(n182) );
  AND4X1_HVT U337 ( .A1(N119), .A2(N117), .A3(N115), .A4(N120), .Y(n181) );
  NAND4X0_HVT U338 ( .A1(n182), .A2(n181), .A3(N126), .A4(N125), .Y(n183) );
  NAND2X0_HVT U339 ( .A1(n183), .A2(N131), .Y(n186) );
endmodule


module conv_top ( clk, srstn, conv_start, fc_done, sram_rdata_a0, 
        sram_rdata_a1, sram_rdata_a2, sram_rdata_a3, sram_rdata_a4, 
        sram_rdata_a5, sram_rdata_a6, sram_rdata_a7, sram_rdata_a8, 
        sram_rdata_b0, sram_rdata_b1, sram_rdata_b2, sram_rdata_b3, 
        sram_rdata_b4, sram_rdata_b5, sram_rdata_b6, sram_rdata_b7, 
        sram_rdata_b8, sram_rdata_weight, sram_raddr_weight, sram_raddr_a0, 
        sram_raddr_a1, sram_raddr_a2, sram_raddr_a3, sram_raddr_a4, 
        sram_raddr_a5, sram_raddr_a6, sram_raddr_a7, sram_raddr_a8, 
        sram_write_enable_b0, sram_write_enable_b1, sram_write_enable_b2, 
        sram_write_enable_b3, sram_write_enable_b4, sram_write_enable_b5, 
        sram_write_enable_b6, sram_write_enable_b7, sram_write_enable_b8, 
        sram_bytemask_b, sram_waddr_b, sram_wdata_b, sram_raddr_b0, 
        sram_raddr_b1, sram_raddr_b2, sram_raddr_b3, sram_raddr_b4, 
        sram_raddr_b5, sram_raddr_b6, sram_raddr_b7, sram_raddr_b8, 
        sram_write_enable_c0, sram_write_enable_c1, sram_write_enable_c2, 
        sram_write_enable_c3, sram_write_enable_c4, sram_bytemask_c, 
        sram_waddr_c, sram_wdata_c, sram_write_enable_d0, sram_write_enable_d1, 
        sram_write_enable_d2, sram_write_enable_d3, sram_write_enable_d4, 
        sram_bytemask_d, sram_waddr_d, sram_wdata_d, conv1_done, conv_done, 
        mem_sel );
  input [31:0] sram_rdata_a0;
  input [31:0] sram_rdata_a1;
  input [31:0] sram_rdata_a2;
  input [31:0] sram_rdata_a3;
  input [31:0] sram_rdata_a4;
  input [31:0] sram_rdata_a5;
  input [31:0] sram_rdata_a6;
  input [31:0] sram_rdata_a7;
  input [31:0] sram_rdata_a8;
  input [31:0] sram_rdata_b0;
  input [31:0] sram_rdata_b1;
  input [31:0] sram_rdata_b2;
  input [31:0] sram_rdata_b3;
  input [31:0] sram_rdata_b4;
  input [31:0] sram_rdata_b5;
  input [31:0] sram_rdata_b6;
  input [31:0] sram_rdata_b7;
  input [31:0] sram_rdata_b8;
  input [99:0] sram_rdata_weight;
  output [16:0] sram_raddr_weight;
  output [9:0] sram_raddr_a0;
  output [9:0] sram_raddr_a1;
  output [9:0] sram_raddr_a2;
  output [9:0] sram_raddr_a3;
  output [9:0] sram_raddr_a4;
  output [9:0] sram_raddr_a5;
  output [9:0] sram_raddr_a6;
  output [9:0] sram_raddr_a7;
  output [9:0] sram_raddr_a8;
  output [3:0] sram_bytemask_b;
  output [9:0] sram_waddr_b;
  output [7:0] sram_wdata_b;
  output [9:0] sram_raddr_b0;
  output [9:0] sram_raddr_b1;
  output [9:0] sram_raddr_b2;
  output [9:0] sram_raddr_b3;
  output [9:0] sram_raddr_b4;
  output [9:0] sram_raddr_b5;
  output [9:0] sram_raddr_b6;
  output [9:0] sram_raddr_b7;
  output [9:0] sram_raddr_b8;
  output [3:0] sram_bytemask_c;
  output [9:0] sram_waddr_c;
  output [7:0] sram_wdata_c;
  output [3:0] sram_bytemask_d;
  output [9:0] sram_waddr_d;
  output [7:0] sram_wdata_d;
  input clk, srstn, conv_start, fc_done;
  output sram_write_enable_b0, sram_write_enable_b1, sram_write_enable_b2,
         sram_write_enable_b3, sram_write_enable_b4, sram_write_enable_b5,
         sram_write_enable_b6, sram_write_enable_b7, sram_write_enable_b8,
         sram_write_enable_c0, sram_write_enable_c1, sram_write_enable_c2,
         sram_write_enable_c3, sram_write_enable_c4, sram_write_enable_d0,
         sram_write_enable_d1, sram_write_enable_d2, sram_write_enable_d3,
         sram_write_enable_d4, conv1_done, conv_done, mem_sel;
  wire   load_conv1_bias_enable, conv1_bias_set_16_, conv1_bias_set_15_,
         conv1_bias_set_14_, conv1_bias_set_13_, conv1_bias_set_12_,
         conv1_bias_set_11_, conv1_bias_set_10_, conv1_bias_set_9_,
         conv1_bias_set_8_, conv1_bias_set_7_, conv1_bias_set_6_,
         conv1_bias_set_5_, conv1_bias_set_4_, conv1_bias_set_3_,
         conv1_bias_set_2_, conv1_bias_set_1_, conv1_bias_set_0_, set_7_,
         set_6_, set_5_, set_4_, set_3_, set_2_, set_1_, set_0_,
         load_conv2_bias0_enable, load_conv2_bias1_enable, data_out_31_,
         data_out_30_, data_out_29_, data_out_28_, data_out_27_, data_out_26_,
         data_out_25_, data_out_24_, data_out_23_, data_out_22_, data_out_21_,
         data_out_20_, data_out_19_, data_out_18_, data_out_17_, data_out_16_,
         data_out_15_, data_out_14_, data_out_13_, data_out_12_, data_out_11_,
         data_out_10_, data_out_9_, data_out_8_, data_out_7_, data_out_6_,
         data_out_5_, data_out_4_, data_out_3_, data_out_2_, data_out_1_,
         data_out_0_, n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [1:0] mode;
  wire   [3:0] box_sel;
  wire   [4:0] channel;
  wire   [99:0] conv1_weight;
  wire   [99:0] weight;
  wire   [287:0] src_window;
  wire   [3:0] bias_data;

  fsm fsm ( .clk(clk), .srstn(n5), .conv_start(conv_start), .conv1_done(
        conv1_done), .conv_done(conv_done), .fc_done(fc_done), .mode(mode), 
        .mem_sel(mem_sel) );
  conv_control conv_control ( .clk(clk), .srstn(n5), .mode({n7, n1}), 
        .mem_sel(mem_sel), .conv1_done(conv1_done), .sram_raddr_weight(
        sram_raddr_weight), .box_sel(box_sel), .load_conv1_bias_enable(
        load_conv1_bias_enable), .conv1_bias_set({conv1_bias_set_16_, 
        conv1_bias_set_15_, conv1_bias_set_14_, conv1_bias_set_13_, 
        conv1_bias_set_12_, conv1_bias_set_11_, conv1_bias_set_10_, 
        conv1_bias_set_9_, conv1_bias_set_8_, conv1_bias_set_7_, 
        conv1_bias_set_6_, conv1_bias_set_5_, conv1_bias_set_4_, 
        conv1_bias_set_3_, conv1_bias_set_2_, conv1_bias_set_1_, 
        conv1_bias_set_0_}), .sram_raddr_a0(sram_raddr_a0), .sram_raddr_a1(
        sram_raddr_a1), .sram_raddr_a2(sram_raddr_a2), .sram_raddr_a3(
        sram_raddr_a3), .sram_raddr_a4(sram_raddr_a4), .sram_raddr_a5(
        sram_raddr_a5), .sram_raddr_a6(sram_raddr_a6), .sram_raddr_a7(
        sram_raddr_a7), .sram_raddr_a8(sram_raddr_a8), .sram_write_enable_b0(
        sram_write_enable_b0), .sram_write_enable_b1(sram_write_enable_b1), 
        .sram_write_enable_b2(sram_write_enable_b2), .sram_write_enable_b3(
        sram_write_enable_b3), .sram_write_enable_b4(sram_write_enable_b4), 
        .sram_write_enable_b5(sram_write_enable_b5), .sram_write_enable_b6(
        sram_write_enable_b6), .sram_write_enable_b7(sram_write_enable_b7), 
        .sram_write_enable_b8(sram_write_enable_b8), .sram_bytemask_b(
        sram_bytemask_b), .sram_waddr_b(sram_waddr_b), .conv_done(conv_done), 
        .channel(channel), .set({set_7_, set_6_, set_5_, set_4_, set_3_, 
        set_2_, set_1_, set_0_}), .load_conv2_bias0_enable(
        load_conv2_bias0_enable), .load_conv2_bias1_enable(
        load_conv2_bias1_enable), .sram_raddr_b0(sram_raddr_b0), 
        .sram_raddr_b1(sram_raddr_b1), .sram_raddr_b2(sram_raddr_b2), 
        .sram_raddr_b3(sram_raddr_b3), .sram_raddr_b4(sram_raddr_b4), 
        .sram_raddr_b5(sram_raddr_b5), .sram_raddr_b6(sram_raddr_b6), 
        .sram_raddr_b7(sram_raddr_b7), .sram_raddr_b8(sram_raddr_b8), 
        .sram_write_enable_c0(sram_write_enable_c0), .sram_write_enable_c1(
        sram_write_enable_c1), .sram_write_enable_c2(sram_write_enable_c2), 
        .sram_write_enable_c3(sram_write_enable_c3), .sram_write_enable_c4(
        sram_write_enable_c4), .sram_bytemask_c(sram_bytemask_c), 
        .sram_waddr_c(sram_waddr_c), .sram_write_enable_d0(
        sram_write_enable_d0), .sram_write_enable_d1(sram_write_enable_d1), 
        .sram_write_enable_d2(sram_write_enable_d2), .sram_write_enable_d3(
        sram_write_enable_d3), .sram_write_enable_d4(sram_write_enable_d4), 
        .sram_bytemask_d(sram_bytemask_d), .sram_waddr_d(sram_waddr_d) );
  data_reg data_reg ( .clk(clk), .srstn(n4), .mode({n7, n1}), .box_sel(box_sel), .sram_rdata_a0(sram_rdata_a0), .sram_rdata_a1(sram_rdata_a1), 
        .sram_rdata_a2(sram_rdata_a2), .sram_rdata_a3(sram_rdata_a3), 
        .sram_rdata_a4(sram_rdata_a4), .sram_rdata_a5(sram_rdata_a5), 
        .sram_rdata_a6(sram_rdata_a6), .sram_rdata_a7(sram_rdata_a7), 
        .sram_rdata_a8(sram_rdata_a8), .sram_rdata_b0(sram_rdata_b0), 
        .sram_rdata_b1(sram_rdata_b1), .sram_rdata_b2(sram_rdata_b2), 
        .sram_rdata_b3(sram_rdata_b3), .sram_rdata_b4(sram_rdata_b4), 
        .sram_rdata_b5(sram_rdata_b5), .sram_rdata_b6(sram_rdata_b6), 
        .sram_rdata_b7(sram_rdata_b7), .sram_rdata_b8(sram_rdata_b8), 
        .sram_rdata_weight(sram_rdata_weight), .conv1_weight(conv1_weight), 
        .weight(weight), .src_window(src_window) );
  bias_sel bias_sel ( .clk(clk), .srstn(n3), .mode({n7, n1}), 
        .load_conv1_bias_enable(load_conv1_bias_enable), 
        .load_conv2_bias0_enable(load_conv2_bias0_enable), 
        .load_conv2_bias1_enable(load_conv2_bias1_enable), .sram_rdata_weight(
        sram_rdata_weight), .bias_data(bias_data), .conv1_bias_set_5_(
        conv1_bias_set_5_), .conv1_bias_set_4_(conv1_bias_set_4_), 
        .conv1_bias_set_3_(conv1_bias_set_3_), .conv1_bias_set_2_(
        conv1_bias_set_2_), .conv1_bias_set_1_(conv1_bias_set_1_), 
        .conv1_bias_set_0_(conv1_bias_set_0_), .set_5_(set_5_), .set_4_(set_4_), .set_3_(set_3_), .set_2_(set_2_), .set_1_(set_1_), .set_0_(set_0_) );
  multiply_compare multiply_compare ( .clk(clk), .srstn(n6), .mode(mode), 
        .channel(channel), .conv1_sram_rdata_weight(conv1_weight), 
        .conv2_sram_rdata_weight(weight), .src_window(src_window), .data_out({
        data_out_31_, data_out_30_, data_out_29_, data_out_28_, data_out_27_, 
        data_out_26_, data_out_25_, data_out_24_, data_out_23_, data_out_22_, 
        data_out_21_, data_out_20_, data_out_19_, data_out_18_, data_out_17_, 
        data_out_16_, data_out_15_, data_out_14_, data_out_13_, data_out_12_, 
        data_out_11_, data_out_10_, data_out_9_, data_out_8_, data_out_7_, 
        data_out_6_, data_out_5_, data_out_4_, data_out_3_, data_out_2_, 
        data_out_1_, data_out_0_}) );
  quantize quantize ( .clk(clk), .srstn(n4), .bias_data(bias_data), .mode({n7, 
        n1}), .quantized_data(sram_wdata_c), .ori_data_31_(data_out_31_), 
        .ori_data_30_(data_out_30_), .ori_data_29_(data_out_29_), 
        .ori_data_28_(data_out_28_), .ori_data_27_(data_out_27_), 
        .ori_data_26_(data_out_26_), .ori_data_25_(data_out_25_), 
        .ori_data_24_(data_out_24_), .ori_data_23_(data_out_23_), 
        .ori_data_22_(data_out_22_), .ori_data_21_(data_out_21_), 
        .ori_data_20_(data_out_20_), .ori_data_19_(data_out_19_), 
        .ori_data_18_(data_out_18_), .ori_data_17_(data_out_17_), 
        .ori_data_16_(data_out_16_), .ori_data_15_(data_out_15_), 
        .ori_data_14_(data_out_14_), .ori_data_13_(data_out_13_), 
        .ori_data_12_(data_out_12_), .ori_data_11_(data_out_11_), 
        .ori_data_10_(data_out_10_), .ori_data_9_(data_out_9_), .ori_data_8_(
        data_out_8_), .ori_data_7_(data_out_7_), .ori_data_6_(data_out_6_), 
        .ori_data_5_(data_out_5_) );
  NBUFFX4_HVT U1 ( .A(mode[0]), .Y(n1) );
  INVX1_HVT U2 ( .A(n2), .Y(n6) );
  INVX2_HVT U3 ( .A(n2), .Y(n3) );
  INVX8_HVT U4 ( .A(n2), .Y(n5) );
  INVX8_HVT U5 ( .A(srstn), .Y(n2) );
  INVX1_HVT U6 ( .A(n2), .Y(n4) );
  DELLN1X2_HVT U7 ( .A(sram_wdata_c[0]), .Y(sram_wdata_d[0]) );
  DELLN1X2_HVT U8 ( .A(sram_wdata_c[1]), .Y(sram_wdata_b[1]) );
  DELLN1X2_HVT U9 ( .A(sram_wdata_c[2]), .Y(sram_wdata_b[2]) );
  DELLN1X2_HVT U10 ( .A(sram_wdata_c[3]), .Y(sram_wdata_d[3]) );
  DELLN1X2_HVT U11 ( .A(sram_wdata_c[4]), .Y(sram_wdata_d[4]) );
  DELLN1X2_HVT U12 ( .A(sram_wdata_c[5]), .Y(sram_wdata_b[5]) );
  DELLN1X2_HVT U13 ( .A(sram_wdata_c[6]), .Y(sram_wdata_d[6]) );
  DELLN1X2_HVT U14 ( .A(sram_wdata_c[7]), .Y(sram_wdata_d[7]) );
  IBUFFX2_HVT U15 ( .A(mode[1]), .Y(n8) );
  INVX1_HVT U16 ( .A(n8), .Y(n7) );
  NBUFFX2_HVT U17 ( .A(sram_wdata_c[2]), .Y(sram_wdata_d[2]) );
  NBUFFX2_HVT U18 ( .A(sram_wdata_c[5]), .Y(sram_wdata_d[5]) );
  NBUFFX2_HVT U19 ( .A(sram_wdata_c[6]), .Y(sram_wdata_b[6]) );
  NBUFFX2_HVT U20 ( .A(sram_wdata_c[1]), .Y(sram_wdata_d[1]) );
  NBUFFX2_HVT U21 ( .A(sram_wdata_c[3]), .Y(sram_wdata_b[3]) );
  NBUFFX2_HVT U22 ( .A(sram_wdata_c[7]), .Y(sram_wdata_b[7]) );
  NBUFFX2_HVT U23 ( .A(sram_wdata_c[4]), .Y(sram_wdata_b[4]) );
  NBUFFX2_HVT U24 ( .A(sram_wdata_c[0]), .Y(sram_wdata_b[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fc_controller_mydesign_0 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net21976, n1;

  AND2X1_HVT main_gate ( .A1(net21976), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n1), .D(EN), .Q(net21976) );
  INVX0_HVT U1 ( .A(CLK), .Y(n1) );
endmodule


module SNPS_CLOCK_GATE_HIGH_fc_controller_mydesign_1 ( CLK, EN, ENCLK );
  input CLK, EN;
  output ENCLK;
  wire   net21976, n2;

  AND2X1_HVT main_gate ( .A1(net21976), .A2(CLK), .Y(ENCLK) );
  LATCHX1_HVT latch ( .CLK(n2), .D(EN), .Q(net21976) );
  INVX0_HVT U1 ( .A(CLK), .Y(n2) );
endmodule


module fc_controller ( clk, srstn, conv_done, mem_sel, accumulate_reset, 
        fc_state, sram_sel, sram_raddr_c0, sram_raddr_c1, sram_raddr_c2, 
        sram_raddr_c3, sram_raddr_c4, sram_raddr_d0, sram_raddr_d1, 
        sram_raddr_d2, sram_raddr_d3, sram_raddr_d4, sram_raddr_e0, 
        sram_raddr_e1, sram_raddr_e2, sram_raddr_e3, sram_raddr_e4, 
        sram_write_enable_e0, sram_write_enable_e1, sram_write_enable_e2, 
        sram_write_enable_e3, sram_write_enable_e4, sram_write_enable_f, 
        sram_waddr, sram_bytemask, sram_raddr_weight, fc1_done, fc2_done );
  output [1:0] sram_sel;
  output [5:0] sram_raddr_c0;
  output [5:0] sram_raddr_c1;
  output [5:0] sram_raddr_c2;
  output [5:0] sram_raddr_c3;
  output [5:0] sram_raddr_c4;
  output [5:0] sram_raddr_d0;
  output [5:0] sram_raddr_d1;
  output [5:0] sram_raddr_d2;
  output [5:0] sram_raddr_d3;
  output [5:0] sram_raddr_d4;
  output [4:0] sram_raddr_e0;
  output [4:0] sram_raddr_e1;
  output [4:0] sram_raddr_e2;
  output [4:0] sram_raddr_e3;
  output [4:0] sram_raddr_e4;
  output [5:0] sram_waddr;
  output [3:0] sram_bytemask;
  output [14:0] sram_raddr_weight;
  input clk, srstn, conv_done, mem_sel;
  output accumulate_reset, fc_state, sram_write_enable_e0,
         sram_write_enable_e1, sram_write_enable_e2, sram_write_enable_e3,
         sram_write_enable_e4, sram_write_enable_f, fc1_done, fc2_done;
  wire   n_sram_sel_0_, n_write_enable, write_enable, write_e_sram_cnt_2_,
         n_write_enable_delay3, n_write_enable_delay1, n_write_enable_delay2,
         fetch_done, n_data_addr_complete, data_addr_complete, busy,
         n_conv_done_record, conv_done_record, N414, net21993, net21999,
         net22004, net22007, net22010, net22013, net22016, net22019, net22024,
         net22026, net22027, net22028, net22031, n17, n54, n55, n58, n60, n69,
         n99, n127, n128, n129, n1, n2, n5, n6, n7, n8, n10, n11, n12, n13,
         n18, n19, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n42, n43, n44, n45, n46, n48,
         n49, n50, n51, n52, n53, n56, n57, n59, n61, n62, n63, n64, n65, n66,
         n67, n68, n70, n71, n72, n73, n74, n149, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261;
  wire   [2:0] n_state;
  wire   [1:0] state;
  wire   [1:0] bytemask_sel;
  wire   [13:0] n_weight_cnt;
  wire   [5:1] n_row_cnt;

  SNPS_CLOCK_GATE_HIGH_fc_controller_mydesign_0 clk_gate_sram_waddr_reg ( 
        .CLK(clk), .EN(net21993), .ENCLK(net22019) );
  SNPS_CLOCK_GATE_HIGH_fc_controller_mydesign_1 clk_gate_write_e_sram_cnt_reg ( 
        .CLK(clk), .EN(net22024), .ENCLK(net22031) );
  DFFSSRX1_HVT state_reg_0_ ( .D(1'b0), .SETB(n36), .RSTB(n_state[0]), .CLK(
        clk), .Q(state[0]), .QN(n53) );
  DFFSSRX1_HVT n_write_enable_delay2_reg ( .D(1'b0), .SETB(n37), .RSTB(
        n_write_enable_delay3), .CLK(clk), .Q(n_write_enable_delay2) );
  DFFSSRX1_HVT n_write_enable_delay1_reg ( .D(1'b0), .SETB(n36), .RSTB(
        n_write_enable_delay2), .CLK(clk), .Q(n_write_enable_delay1) );
  DFFSSRX1_HVT n_write_enable_reg ( .D(1'b0), .SETB(n36), .RSTB(
        n_write_enable_delay1), .CLK(clk), .Q(n_write_enable), .QN(n44) );
  DFFSSRX1_HVT write_enable_reg ( .D(1'b0), .SETB(n37), .RSTB(n_write_enable), 
        .CLK(clk), .Q(write_enable), .QN(n59) );
  DFFSSRX1_HVT state_reg_2_ ( .D(1'b0), .SETB(n36), .RSTB(n_state[2]), .CLK(
        clk), .Q(n57), .QN(n69) );
  DFFSSRX1_HVT state_reg_1_ ( .D(1'b0), .SETB(n36), .RSTB(n_state[1]), .CLK(
        clk), .Q(state[1]) );
  DFFSSRX1_HVT data_addr_complete_reg ( .D(1'b0), .SETB(n36), .RSTB(
        n_data_addr_complete), .CLK(clk), .Q(data_addr_complete), .QN(n74) );
  DFFSSRX1_HVT row_cnt_reg_5_ ( .D(1'b0), .SETB(n36), .RSTB(n_row_cnt[5]), 
        .CLK(clk), .Q(sram_raddr_d3[5]), .QN(n52) );
  DFFSSRX1_HVT row_cnt_reg_4_ ( .D(1'b0), .SETB(n36), .RSTB(n_row_cnt[4]), 
        .CLK(clk), .Q(sram_raddr_e3[4]), .QN(n50) );
  DFFSSRX1_HVT row_cnt_reg_3_ ( .D(1'b0), .SETB(n37), .RSTB(n_row_cnt[3]), 
        .CLK(clk), .Q(sram_raddr_e3[3]), .QN(n45) );
  DFFSSRX1_HVT row_cnt_reg_2_ ( .D(1'b0), .SETB(n36), .RSTB(n_row_cnt[2]), 
        .CLK(clk), .Q(sram_raddr_e3[2]), .QN(n46) );
  DFFSSRX1_HVT row_cnt_reg_1_ ( .D(1'b0), .SETB(n36), .RSTB(n_row_cnt[1]), 
        .CLK(clk), .Q(sram_raddr_e3[1]), .QN(n56) );
  DFFSSRX1_HVT row_cnt_reg_0_ ( .D(1'b0), .SETB(n37), .RSTB(n210), .CLK(clk), 
        .Q(sram_raddr_e3[0]), .QN(n51) );
  DFFSSRX1_HVT weight_cnt_reg_12_ ( .D(1'b0), .SETB(n36), .RSTB(n60), .CLK(clk), .Q(sram_raddr_weight[12]) );
  DFFSSRX1_HVT weight_cnt_reg_0_ ( .D(1'b0), .SETB(n36), .RSTB(n_weight_cnt[0]), .CLK(clk), .Q(sram_raddr_weight[0]), .QN(n61) );
  DFFSSRX1_HVT weight_cnt_reg_10_ ( .D(1'b0), .SETB(n37), .RSTB(n200), .CLK(
        clk), .Q(sram_raddr_weight[10]), .QN(n67) );
  DFFSSRX1_HVT weight_cnt_reg_11_ ( .D(1'b0), .SETB(n36), .RSTB(n201), .CLK(
        clk), .Q(sram_raddr_weight[11]), .QN(n68) );
  DFFSSRX1_HVT weight_cnt_reg_3_ ( .D(1'b0), .SETB(n36), .RSTB(n202), .CLK(clk), .Q(sram_raddr_weight[3]), .QN(n71) );
  DFFSSRX1_HVT weight_cnt_reg_4_ ( .D(1'b0), .SETB(n36), .RSTB(n205), .CLK(clk), .Q(sram_raddr_weight[4]), .QN(n62) );
  DFFSSRX1_HVT weight_cnt_reg_6_ ( .D(1'b0), .SETB(n37), .RSTB(n206), .CLK(clk), .Q(sram_raddr_weight[6]), .QN(n72) );
  DFFSSRX1_HVT weight_cnt_reg_5_ ( .D(1'b0), .SETB(n37), .RSTB(n_weight_cnt[5]), .CLK(clk), .Q(sram_raddr_weight[5]) );
  DFFSSRX1_HVT weight_cnt_reg_8_ ( .D(1'b0), .SETB(n37), .RSTB(n203), .CLK(clk), .Q(sram_raddr_weight[8]) );
  DFFSSRX1_HVT weight_cnt_reg_9_ ( .D(1'b0), .SETB(n36), .RSTB(n199), .CLK(clk), .Q(sram_raddr_weight[9]), .QN(n66) );
  DFFSSRX1_HVT weight_cnt_reg_7_ ( .D(1'b0), .SETB(n36), .RSTB(n207), .CLK(clk), .Q(sram_raddr_weight[7]), .QN(n64) );
  DFFSSRX1_HVT weight_cnt_reg_14_ ( .D(1'b0), .SETB(n37), .RSTB(n209), .CLK(
        clk), .Q(sram_raddr_weight[14]), .QN(n63) );
  DFFSSRX1_HVT weight_cnt_reg_13_ ( .D(1'b0), .SETB(n36), .RSTB(
        n_weight_cnt[13]), .CLK(clk), .Q(sram_raddr_weight[13]) );
  DFFSSRX1_HVT weight_cnt_reg_1_ ( .D(1'b0), .SETB(n37), .RSTB(n_weight_cnt[1]), .CLK(clk), .Q(sram_raddr_weight[1]) );
  DFFSSRX1_HVT weight_cnt_reg_2_ ( .D(1'b0), .SETB(n36), .RSTB(n204), .CLK(clk), .Q(sram_raddr_weight[2]), .QN(n65) );
  DFFSSRX1_HVT sram_sel_reg_0_ ( .D(1'b0), .SETB(n37), .RSTB(n_sram_sel_0_), 
        .CLK(clk), .Q(sram_sel[0]) );
  DFFSSRX1_HVT sram_sel_reg_1_ ( .D(n17), .SETB(n99), .RSTB(srstn), .CLK(clk), 
        .Q(sram_sel[1]) );
  DFFSSRX1_HVT fetch_done_reg ( .D(1'b0), .SETB(n37), .RSTB(n129), .CLK(clk), 
        .Q(fetch_done), .QN(n73) );
  DFFSSRX1_HVT fc2_done_reg ( .D(1'b0), .SETB(n37), .RSTB(n208), .CLK(clk), 
        .Q(fc2_done), .QN(n58) );
  DFFSSRX1_HVT fc1_done_reg ( .D(1'b0), .SETB(n37), .RSTB(n211), .CLK(clk), 
        .Q(fc1_done) );
  DFFSSRX1_HVT bytemask_sel_reg_0_ ( .D(1'b0), .SETB(n36), .RSTB(n128), .CLK(
        clk), .Q(bytemask_sel[0]), .QN(n49) );
  DFFSSRX1_HVT bytemask_sel_reg_1_ ( .D(1'b0), .SETB(n37), .RSTB(n127), .CLK(
        clk), .Q(bytemask_sel[1]), .QN(n43) );
  DFFSSRX1_HVT write_e_sram_cnt_reg_0_ ( .D(1'b0), .SETB(n36), .RSTB(net22028), 
        .CLK(net22031), .Q(n42), .QN(n55) );
  DFFSSRX1_HVT write_e_sram_cnt_reg_1_ ( .D(1'b0), .SETB(n37), .RSTB(net22027), 
        .CLK(net22031), .Q(n48), .QN(n54) );
  DFFSSRX1_HVT write_e_sram_cnt_reg_2_ ( .D(1'b0), .SETB(n37), .RSTB(net22026), 
        .CLK(net22031), .Q(write_e_sram_cnt_2_) );
  DFFSSRX1_HVT sram_waddr_reg_0_ ( .D(1'b0), .SETB(n37), .RSTB(net22016), 
        .CLK(net22019), .Q(sram_waddr[0]) );
  DFFSSRX1_HVT sram_waddr_reg_1_ ( .D(1'b0), .SETB(n37), .RSTB(net22013), 
        .CLK(net22019), .Q(sram_waddr[1]) );
  DFFSSRX1_HVT sram_waddr_reg_2_ ( .D(1'b0), .SETB(n37), .RSTB(net22010), 
        .CLK(net22019), .Q(sram_waddr[2]) );
  DFFSSRX1_HVT sram_waddr_reg_3_ ( .D(1'b0), .SETB(n36), .RSTB(net22007), 
        .CLK(net22019), .Q(sram_waddr[3]) );
  DFFSSRX1_HVT sram_waddr_reg_4_ ( .D(1'b0), .SETB(n36), .RSTB(net22004), 
        .CLK(net22019), .Q(sram_waddr[4]) );
  DFFSSRX1_HVT sram_waddr_reg_5_ ( .D(1'b0), .SETB(n37), .RSTB(net21999), 
        .CLK(net22019), .Q(sram_waddr[5]), .QN(n70) );
  DFFSSRX1_HVT busy_reg ( .D(1'b0), .SETB(n37), .RSTB(N414), .CLK(clk), .Q(
        busy) );
  DFFSSRX1_HVT conv_done_record_reg ( .D(1'b0), .SETB(n36), .RSTB(
        n_conv_done_record), .CLK(clk), .Q(conv_done_record) );
  OA221X1_HVT U3 ( .A1(1'b0), .A2(n175), .A3(n172), .A4(sram_raddr_e3[2]), 
        .A5(n19), .Y(n_row_cnt[2]) );
  OA221X1_HVT U4 ( .A1(1'b0), .A2(n249), .A3(sram_waddr[3]), .A4(n18), .A5(
        n252), .Y(net22007) );
  OA221X1_HVT U5 ( .A1(1'b0), .A2(n238), .A3(sram_raddr_weight[12]), .A4(n239), 
        .A5(n196), .Y(n60) );
  OA221X1_HVT U6 ( .A1(1'b0), .A2(n248), .A3(sram_waddr[4]), .A4(n247), .A5(
        n252), .Y(net22004) );
  OA221X1_HVT U7 ( .A1(1'b0), .A2(n196), .A3(sram_raddr_weight[8]), .A4(n225), 
        .A5(n224), .Y(n203) );
  OA221X1_HVT U8 ( .A1(1'b0), .A2(n237), .A3(sram_raddr_weight[13]), .A4(n220), 
        .A5(n196), .Y(n_weight_cnt[13]) );
  OA221X1_HVT U9 ( .A1(1'b0), .A2(n196), .A3(sram_raddr_weight[1]), .A4(
        sram_raddr_weight[0]), .A5(n219), .Y(n_weight_cnt[1]) );
  INVX0_HVT U10 ( .A(state[1]), .Y(n1) );
  NAND2X0_HVT U11 ( .A1(n162), .A2(n1), .Y(n169) );
  NOR4X1_HVT U12 ( .A1(state[0]), .A2(state[1]), .A3(n57), .A4(busy), .Y(n2)
         );
  AO222X1_HVT U13 ( .A1(n194), .A2(n73), .A3(n211), .A4(n198), .A5(n218), .A6(
        n2), .Y(n163) );
  INVX0_HVT U16 ( .A(n63), .Y(n5) );
  INVX0_HVT U17 ( .A(n237), .Y(n6) );
  OA221X1_HVT U18 ( .A1(n63), .A2(n237), .A3(n5), .A4(n6), .A5(n196), .Y(n209)
         );
  INVX0_HVT U19 ( .A(n64), .Y(n7) );
  INVX0_HVT U20 ( .A(n228), .Y(n8) );
  OA221X1_HVT U21 ( .A1(n64), .A2(n228), .A3(n7), .A4(n8), .A5(n196), .Y(n207)
         );
  NAND3X0_HVT U23 ( .A1(sram_waddr[3]), .A2(sram_waddr[4]), .A3(n251), .Y(n10)
         );
  OR3X1_HVT U24 ( .A1(sram_waddr[0]), .A2(sram_waddr[5]), .A3(n10), .Y(n11) );
  AO221X1_HVT U25 ( .A1(n198), .A2(sram_waddr[2]), .A3(n198), .A4(n11), .A5(
        n189), .Y(n252) );
  INVX0_HVT U26 ( .A(n232), .Y(n12) );
  INVX0_HVT U27 ( .A(n62), .Y(n13) );
  OA221X1_HVT U28 ( .A1(n232), .A2(n62), .A3(n12), .A4(n13), .A5(n196), .Y(
        n205) );
  INVX0_HVT U32 ( .A(n250), .Y(n18) );
  INVX0_HVT U33 ( .A(n173), .Y(n19) );
  NAND3X0_HVT U35 ( .A1(srstn), .A2(n197), .A3(n198), .Y(net22024) );
  AO21X1_HVT U36 ( .A1(sram_waddr[1]), .A2(sram_waddr[0]), .A3(sram_waddr[2]), 
        .Y(n21) );
  AND3X1_HVT U37 ( .A1(n250), .A2(n252), .A3(n21), .Y(net22010) );
  INVX0_HVT U38 ( .A(n173), .Y(n22) );
  INVX0_HVT U39 ( .A(sram_raddr_e3[3]), .Y(n23) );
  OA221X1_HVT U40 ( .A1(n173), .A2(sram_raddr_e3[3]), .A3(n22), .A4(n23), .A5(
        n175), .Y(n_row_cnt[3]) );
  AO21X1_HVT U41 ( .A1(n59), .A2(bytemask_sel[1]), .A3(sram_bytemask[1]), .Y(
        n24) );
  OA221X1_HVT U42 ( .A1(n24), .A2(sram_bytemask[2]), .A3(n24), .A4(
        write_enable), .A5(n58), .Y(n127) );
  INVX0_HVT U43 ( .A(n174), .Y(n25) );
  INVX0_HVT U44 ( .A(sram_raddr_e3[4]), .Y(n26) );
  OA221X1_HVT U45 ( .A1(n174), .A2(sram_raddr_e3[4]), .A3(n25), .A4(n26), .A5(
        n175), .Y(n_row_cnt[4]) );
  NOR4X0_HVT U46 ( .A1(sram_raddr_weight[0]), .A2(sram_raddr_weight[1]), .A3(
        n240), .A4(n204), .Y(n27) );
  NAND4X0_HVT U47 ( .A1(n203), .A2(n202), .A3(n205), .A4(n27), .Y(n28) );
  OR3X1_HVT U48 ( .A1(n206), .A2(n207), .A3(n28), .Y(n29) );
  NAND3X0_HVT U49 ( .A1(n200), .A2(n199), .A3(n201), .Y(n30) );
  NOR4X0_HVT U50 ( .A1(n60), .A2(n_weight_cnt[13]), .A3(n29), .A4(n30), .Y(n31) );
  OA221X1_HVT U51 ( .A1(data_addr_complete), .A2(n209), .A3(data_addr_complete), .A4(n31), .A5(n189), .Y(n_data_addr_complete) );
  INVX0_HVT U52 ( .A(bytemask_sel[0]), .Y(n32) );
  INVX0_HVT U53 ( .A(write_enable), .Y(n33) );
  OA221X1_HVT U54 ( .A1(bytemask_sel[0]), .A2(write_enable), .A3(n32), .A4(n33), .A5(n58), .Y(n128) );
  NAND2X0_HVT U55 ( .A1(n174), .A2(sram_raddr_e3[4]), .Y(n34) );
  HADDX1_HVT U56 ( .A0(n52), .B0(n34), .SO(n35) );
  AND2X1_HVT U57 ( .A1(n175), .A2(n35), .Y(n_row_cnt[5]) );
  INVX1_HVT U58 ( .A(n233), .Y(n239) );
  INVX2_HVT U59 ( .A(srstn), .Y(n36) );
  INVX0_HVT U60 ( .A(n238), .Y(n220) );
  INVX0_HVT U61 ( .A(n235), .Y(n234) );
  INVX0_HVT U62 ( .A(n222), .Y(n236) );
  INVX0_HVT U63 ( .A(n224), .Y(n223) );
  INVX0_HVT U64 ( .A(n228), .Y(n221) );
  INVX0_HVT U65 ( .A(n226), .Y(n229) );
  INVX0_HVT U66 ( .A(n248), .Y(n246) );
  INVX0_HVT U67 ( .A(n39), .Y(sram_raddr_e2[0]) );
  INVX0_HVT U68 ( .A(n39), .Y(sram_raddr_e4[0]) );
  INVX0_HVT U69 ( .A(n38), .Y(sram_raddr_e4[1]) );
  INVX0_HVT U70 ( .A(n50), .Y(sram_raddr_e1[4]) );
  INVX0_HVT U71 ( .A(n56), .Y(sram_raddr_e1[1]) );
  INVX0_HVT U72 ( .A(n50), .Y(sram_raddr_e4[4]) );
  INVX0_HVT U73 ( .A(n39), .Y(sram_raddr_c1[0]) );
  INVX0_HVT U74 ( .A(n39), .Y(sram_raddr_d4[0]) );
  INVX0_HVT U75 ( .A(n56), .Y(sram_raddr_d4[1]) );
  INVX0_HVT U76 ( .A(n40), .Y(sram_raddr_c2[4]) );
  INVX0_HVT U77 ( .A(n40), .Y(sram_raddr_d4[4]) );
  INVX0_HVT U78 ( .A(n38), .Y(sram_raddr_c2[1]) );
  INVX0_HVT U79 ( .A(n51), .Y(sram_raddr_c2[0]) );
  INVX0_HVT U80 ( .A(n40), .Y(sram_raddr_c3[4]) );
  INVX0_HVT U81 ( .A(n38), .Y(sram_raddr_c3[1]) );
  INVX0_HVT U82 ( .A(n51), .Y(sram_raddr_c3[0]) );
  INVX0_HVT U83 ( .A(n51), .Y(sram_raddr_d3[0]) );
  INVX0_HVT U84 ( .A(n50), .Y(sram_raddr_c4[4]) );
  INVX0_HVT U85 ( .A(n38), .Y(sram_raddr_c4[1]) );
  INVX0_HVT U86 ( .A(n39), .Y(sram_raddr_c4[0]) );
  INVX0_HVT U87 ( .A(n56), .Y(sram_raddr_d3[1]) );
  INVX0_HVT U88 ( .A(n40), .Y(sram_raddr_d0[4]) );
  INVX0_HVT U89 ( .A(n40), .Y(sram_raddr_d3[4]) );
  INVX0_HVT U90 ( .A(n38), .Y(sram_raddr_d0[1]) );
  INVX0_HVT U91 ( .A(n39), .Y(sram_raddr_d2[0]) );
  INVX0_HVT U92 ( .A(n39), .Y(sram_raddr_d0[0]) );
  INVX0_HVT U93 ( .A(n40), .Y(sram_raddr_e2[4]) );
  INVX0_HVT U94 ( .A(n39), .Y(sram_raddr_e1[0]) );
  INVX0_HVT U95 ( .A(n56), .Y(sram_raddr_d2[1]) );
  INVX0_HVT U96 ( .A(n40), .Y(sram_raddr_d1[4]) );
  INVX0_HVT U97 ( .A(n56), .Y(sram_raddr_d1[1]) );
  INVX0_HVT U98 ( .A(n40), .Y(sram_raddr_d2[4]) );
  INVX0_HVT U99 ( .A(n39), .Y(sram_raddr_d1[0]) );
  INVX0_HVT U100 ( .A(n56), .Y(sram_raddr_e2[1]) );
  INVX0_HVT U101 ( .A(n40), .Y(sram_raddr_c0[4]) );
  INVX0_HVT U102 ( .A(n38), .Y(sram_raddr_c0[1]) );
  INVX0_HVT U103 ( .A(n39), .Y(sram_raddr_e0[0]) );
  INVX0_HVT U104 ( .A(n39), .Y(sram_raddr_c0[0]) );
  INVX0_HVT U105 ( .A(n40), .Y(sram_raddr_c1[4]) );
  INVX0_HVT U106 ( .A(n56), .Y(sram_raddr_e0[1]) );
  INVX0_HVT U107 ( .A(n40), .Y(sram_raddr_e0[4]) );
  INVX0_HVT U108 ( .A(n38), .Y(sram_raddr_c1[1]) );
  INVX0_HVT U109 ( .A(n164), .Y(n166) );
  INVX0_HVT U110 ( .A(n215), .Y(n216) );
  INVX0_HVT U111 ( .A(n189), .Y(n185) );
  INVX0_HVT U112 ( .A(sram_waddr[1]), .Y(n251) );
  INVX0_HVT U113 ( .A(sram_waddr[0]), .Y(n253) );
  INVX0_HVT U114 ( .A(n191), .Y(sram_raddr_e4[2]) );
  INVX0_HVT U115 ( .A(n167), .Y(sram_raddr_e4[3]) );
  INVX0_HVT U116 ( .A(n149), .Y(sram_raddr_d4[5]) );
  INVX0_HVT U117 ( .A(n232), .Y(n230) );
  INVX0_HVT U118 ( .A(n149), .Y(sram_raddr_d2[5]) );
  INVX0_HVT U119 ( .A(n149), .Y(sram_raddr_d1[5]) );
  INVX0_HVT U120 ( .A(n149), .Y(sram_raddr_d0[5]) );
  INVX0_HVT U121 ( .A(n149), .Y(sram_raddr_c4[5]) );
  INVX0_HVT U122 ( .A(n149), .Y(sram_raddr_c3[5]) );
  INVX0_HVT U123 ( .A(n149), .Y(sram_raddr_c2[5]) );
  INVX0_HVT U124 ( .A(n191), .Y(sram_raddr_c1[2]) );
  INVX0_HVT U125 ( .A(n167), .Y(sram_raddr_c1[3]) );
  INVX0_HVT U126 ( .A(n149), .Y(sram_raddr_c1[5]) );
  INVX0_HVT U127 ( .A(n191), .Y(sram_raddr_c0[2]) );
  INVX0_HVT U128 ( .A(n167), .Y(sram_raddr_c0[3]) );
  INVX0_HVT U129 ( .A(n149), .Y(sram_raddr_c0[5]) );
  INVX0_HVT U130 ( .A(n46), .Y(sram_raddr_e2[2]) );
  INVX0_HVT U131 ( .A(n45), .Y(sram_raddr_e2[3]) );
  INVX0_HVT U132 ( .A(n46), .Y(sram_raddr_e1[2]) );
  INVX0_HVT U133 ( .A(n45), .Y(sram_raddr_e1[3]) );
  INVX0_HVT U134 ( .A(n46), .Y(sram_raddr_e0[2]) );
  INVX0_HVT U135 ( .A(n45), .Y(sram_raddr_e0[3]) );
  INVX0_HVT U136 ( .A(n46), .Y(sram_raddr_d4[2]) );
  INVX0_HVT U137 ( .A(n45), .Y(sram_raddr_d4[3]) );
  INVX0_HVT U138 ( .A(n46), .Y(sram_raddr_d3[2]) );
  INVX0_HVT U139 ( .A(n45), .Y(sram_raddr_d3[3]) );
  INVX0_HVT U140 ( .A(n46), .Y(sram_raddr_d2[2]) );
  INVX0_HVT U141 ( .A(n45), .Y(sram_raddr_d2[3]) );
  INVX0_HVT U142 ( .A(n46), .Y(sram_raddr_d1[2]) );
  INVX0_HVT U143 ( .A(n45), .Y(sram_raddr_d1[3]) );
  INVX0_HVT U144 ( .A(n46), .Y(sram_raddr_d0[2]) );
  INVX0_HVT U145 ( .A(n45), .Y(sram_raddr_d0[3]) );
  INVX0_HVT U146 ( .A(n46), .Y(sram_raddr_c4[2]) );
  INVX0_HVT U147 ( .A(n45), .Y(sram_raddr_c4[3]) );
  INVX0_HVT U148 ( .A(n46), .Y(sram_raddr_c3[2]) );
  INVX0_HVT U149 ( .A(n45), .Y(sram_raddr_c3[3]) );
  INVX0_HVT U150 ( .A(n46), .Y(sram_raddr_c2[2]) );
  INVX0_HVT U151 ( .A(n45), .Y(sram_raddr_c2[3]) );
  INVX2_HVT U152 ( .A(srstn), .Y(n37) );
  INVX1_HVT U153 ( .A(sram_raddr_e3[1]), .Y(n38) );
  INVX1_HVT U154 ( .A(sram_raddr_e3[0]), .Y(n39) );
  INVX1_HVT U155 ( .A(sram_raddr_e3[4]), .Y(n40) );
  INVX1_HVT U156 ( .A(n169), .Y(n194) );
  NAND3X0_HVT U157 ( .A1(n164), .A2(n187), .A3(n169), .Y(n196) );
  INVX1_HVT U158 ( .A(n198), .Y(n187) );
  AND2X1_HVT U159 ( .A1(n159), .A2(n53), .Y(n198) );
  INVX1_HVT U160 ( .A(sram_raddr_d3[5]), .Y(n149) );
  INVX1_HVT U161 ( .A(sram_raddr_e3[2]), .Y(n191) );
  INVX1_HVT U162 ( .A(sram_raddr_e3[3]), .Y(n167) );
  AO21X1_HVT U163 ( .A1(n189), .A2(n178), .A3(n163), .Y(n_state[0]) );
  AND2X1_HVT U164 ( .A1(n49), .A2(n43), .Y(sram_bytemask[3]) );
  AND2X1_HVT U165 ( .A1(bytemask_sel[0]), .A2(n43), .Y(sram_bytemask[2]) );
  NAND2X0_HVT U166 ( .A1(n195), .A2(n44), .Y(accumulate_reset) );
  NAND3X0_HVT U167 ( .A1(n194), .A2(n193), .A3(n192), .Y(n195) );
  AND2X1_HVT U168 ( .A1(bytemask_sel[0]), .A2(bytemask_sel[1]), .Y(
        sram_bytemask[0]) );
  INVX1_HVT U169 ( .A(n249), .Y(n247) );
  INVX1_HVT U170 ( .A(n178), .Y(n208) );
  NOR4X1_HVT U171 ( .A1(sram_raddr_weight[11]), .A2(sram_raddr_weight[10]), 
        .A3(sram_raddr_weight[9]), .A4(n214), .Y(n259) );
  OR2X1_HVT U172 ( .A1(n59), .A2(n244), .Y(n178) );
  AND2X1_HVT U173 ( .A1(state[1]), .A2(n69), .Y(n159) );
  NAND2X0_HVT U174 ( .A1(n178), .A2(n159), .Y(n161) );
  AND2X1_HVT U175 ( .A1(state[0]), .A2(n69), .Y(n162) );
  NAND2X0_HVT U176 ( .A1(n194), .A2(fetch_done), .Y(n160) );
  NAND3X0_HVT U177 ( .A1(n161), .A2(n187), .A3(n160), .Y(n_state[1]) );
  AND2X1_HVT U178 ( .A1(n162), .A2(state[1]), .Y(n189) );
  AND4X1_HVT U179 ( .A1(n258), .A2(write_enable), .A3(n241), .A4(
        sram_raddr_weight[0]), .Y(n211) );
  OR3X1_HVT U180 ( .A1(n189), .A2(n163), .A3(n_state[1]), .Y(N414) );
  NAND2X0_HVT U181 ( .A1(n189), .A2(n74), .Y(n164) );
  AND2X1_HVT U182 ( .A1(n196), .A2(n61), .Y(n_weight_cnt[0]) );
  AND4X1_HVT U183 ( .A1(n56), .A2(n52), .A3(n51), .A4(sram_raddr_e3[4]), .Y(
        n165) );
  NAND3X0_HVT U184 ( .A1(n165), .A2(sram_raddr_e3[3]), .A3(n191), .Y(n176) );
  NAND2X0_HVT U185 ( .A1(n166), .A2(n176), .Y(n170) );
  AND2X1_HVT U186 ( .A1(sram_raddr_e3[1]), .A2(sram_raddr_e3[0]), .Y(n172) );
  AND2X1_HVT U187 ( .A1(n172), .A2(sram_raddr_e3[2]), .Y(n173) );
  AND2X1_HVT U188 ( .A1(n167), .A2(n50), .Y(n193) );
  NAND3X0_HVT U189 ( .A1(n173), .A2(sram_raddr_d3[5]), .A3(n193), .Y(n177) );
  NAND2X0_HVT U190 ( .A1(n177), .A2(n198), .Y(n168) );
  NAND3X0_HVT U191 ( .A1(n170), .A2(n169), .A3(n168), .Y(n175) );
  AND2X1_HVT U192 ( .A1(n175), .A2(n51), .Y(n210) );
  AND2X1_HVT U193 ( .A1(n56), .A2(sram_raddr_e3[0]), .Y(n171) );
  AO22X1_HVT U194 ( .A1(n171), .A2(n175), .A3(n210), .A4(sram_raddr_e3[1]), 
        .Y(n_row_cnt[1]) );
  AND2X1_HVT U195 ( .A1(n173), .A2(sram_raddr_e3[3]), .Y(n174) );
  OAI22X1_HVT U196 ( .A1(n187), .A2(n177), .A3(n185), .A4(n176), .Y(
        n_write_enable_delay3) );
  AND2X1_HVT U197 ( .A1(n208), .A2(n189), .Y(n_state[2]) );
  NAND2X0_HVT U198 ( .A1(n226), .A2(n72), .Y(n179) );
  AND3X1_HVT U199 ( .A1(n179), .A2(n228), .A3(n196), .Y(n206) );
  NAND2X0_HVT U200 ( .A1(n219), .A2(n65), .Y(n180) );
  AND3X1_HVT U201 ( .A1(n196), .A2(n231), .A3(n180), .Y(n204) );
  NAND2X0_HVT U202 ( .A1(n231), .A2(n71), .Y(n181) );
  AND3X1_HVT U203 ( .A1(n196), .A2(n232), .A3(n181), .Y(n202) );
  NAND2X0_HVT U204 ( .A1(n68), .A2(n235), .Y(n182) );
  AND3X1_HVT U205 ( .A1(n196), .A2(n233), .A3(n182), .Y(n201) );
  NAND2X0_HVT U206 ( .A1(n67), .A2(n222), .Y(n183) );
  AND3X1_HVT U207 ( .A1(n196), .A2(n235), .A3(n183), .Y(n200) );
  NAND2X0_HVT U208 ( .A1(n66), .A2(n224), .Y(n184) );
  AND3X1_HVT U209 ( .A1(n196), .A2(n222), .A3(n184), .Y(n199) );
  AND3X1_HVT U210 ( .A1(n198), .A2(n261), .A3(n55), .Y(net22028) );
  NAND2X0_HVT U211 ( .A1(n187), .A2(n185), .Y(n186) );
  NAND2X0_HVT U212 ( .A1(write_enable), .A2(sram_bytemask[0]), .Y(n197) );
  AND2X1_HVT U213 ( .A1(n198), .A2(n261), .Y(n188) );
  AO21X1_HVT U214 ( .A1(n186), .A2(n197), .A3(n188), .Y(n245) );
  OR3X1_HVT U215 ( .A1(write_e_sram_cnt_2_), .A2(n256), .A3(n187), .Y(n255) );
  NAND3X0_HVT U216 ( .A1(n188), .A2(write_e_sram_cnt_2_), .A3(n256), .Y(n254)
         );
  NAND2X0_HVT U217 ( .A1(n198), .A2(write_enable), .Y(n190) );
  NOR2X0_HVT U218 ( .A1(write_e_sram_cnt_2_), .A2(n190), .Y(n260) );
  NAND2X0_HVT U219 ( .A1(n189), .A2(write_enable), .Y(sram_write_enable_f) );
  OR2X1_HVT U220 ( .A1(n261), .A2(n190), .Y(sram_write_enable_e4) );
  AND4X1_HVT U221 ( .A1(n191), .A2(n52), .A3(n51), .A4(sram_raddr_e3[1]), .Y(
        n192) );
  AND3X1_HVT U222 ( .A1(n198), .A2(n256), .A3(n257), .Y(net22027) );
  AND2X1_HVT U223 ( .A1(n240), .A2(n196), .Y(n_weight_cnt[5]) );
  OR4X1_HVT U224 ( .A1(sram_raddr_weight[7]), .A2(sram_raddr_weight[6]), .A3(
        sram_raddr_weight[4]), .A4(sram_raddr_weight[2]), .Y(n212) );
  OR3X1_HVT U225 ( .A1(sram_raddr_weight[8]), .A2(sram_raddr_weight[3]), .A3(
        n212), .Y(n213) );
  OR3X1_HVT U226 ( .A1(sram_raddr_weight[13]), .A2(sram_raddr_weight[12]), 
        .A3(n213), .Y(n215) );
  NOR3X0_HVT U227 ( .A1(sram_raddr_weight[0]), .A2(sram_raddr_weight[1]), .A3(
        n215), .Y(n242) );
  OR2X1_HVT U228 ( .A1(sram_raddr_weight[14]), .A2(sram_raddr_weight[5]), .Y(
        n214) );
  NAND2X0_HVT U229 ( .A1(n242), .A2(n259), .Y(n244) );
  AND2X1_HVT U230 ( .A1(sram_raddr_weight[1]), .A2(n216), .Y(n258) );
  AND3X1_HVT U231 ( .A1(sram_raddr_weight[14]), .A2(sram_raddr_weight[11]), 
        .A3(sram_raddr_weight[5]), .Y(n217) );
  AND3X1_HVT U232 ( .A1(sram_raddr_weight[10]), .A2(sram_raddr_weight[9]), 
        .A3(n217), .Y(n241) );
  OR2X1_HVT U233 ( .A1(conv_done_record), .A2(conv_done), .Y(n218) );
  AND2X1_HVT U234 ( .A1(n_state[1]), .A2(n_state[0]), .Y(fc_state) );
  AND2X1_HVT U235 ( .A1(busy), .A2(n218), .Y(n_conv_done_record) );
  NAND2X0_HVT U237 ( .A1(sram_raddr_weight[0]), .A2(sram_raddr_weight[1]), .Y(
        n219) );
  NAND3X0_HVT U238 ( .A1(sram_raddr_weight[2]), .A2(sram_raddr_weight[0]), 
        .A3(sram_raddr_weight[1]), .Y(n231) );
  NAND4X0_HVT U239 ( .A1(sram_raddr_weight[3]), .A2(sram_raddr_weight[2]), 
        .A3(sram_raddr_weight[0]), .A4(sram_raddr_weight[1]), .Y(n232) );
  AND2X1_HVT U240 ( .A1(sram_raddr_weight[4]), .A2(n230), .Y(n227) );
  NAND2X0_HVT U241 ( .A1(sram_raddr_weight[5]), .A2(n227), .Y(n226) );
  NAND2X0_HVT U242 ( .A1(sram_raddr_weight[6]), .A2(n229), .Y(n228) );
  AND2X1_HVT U243 ( .A1(sram_raddr_weight[7]), .A2(n221), .Y(n225) );
  NAND2X0_HVT U244 ( .A1(sram_raddr_weight[8]), .A2(n225), .Y(n224) );
  NAND2X0_HVT U245 ( .A1(sram_raddr_weight[9]), .A2(n223), .Y(n222) );
  NAND2X0_HVT U246 ( .A1(sram_raddr_weight[10]), .A2(n236), .Y(n235) );
  NAND2X0_HVT U247 ( .A1(sram_raddr_weight[11]), .A2(n234), .Y(n233) );
  NAND2X0_HVT U248 ( .A1(sram_raddr_weight[12]), .A2(n239), .Y(n238) );
  NAND2X0_HVT U249 ( .A1(sram_raddr_weight[13]), .A2(n220), .Y(n237) );
  OA21X1_HVT U250 ( .A1(sram_raddr_weight[5]), .A2(n227), .A3(n226), .Y(n240)
         );
  AND2X1_HVT U251 ( .A1(n242), .A2(n241), .Y(n17) );
  NAND2X0_HVT U252 ( .A1(sram_sel[0]), .A2(n244), .Y(n243) );
  OAI22X1_HVT U253 ( .A1(n17), .A2(n243), .A3(mem_sel), .A4(n244), .Y(
        n_sram_sel_0_) );
  NAND2X0_HVT U254 ( .A1(sram_sel[1]), .A2(n244), .Y(n99) );
  NAND3X0_HVT U255 ( .A1(n55), .A2(n54), .A3(write_e_sram_cnt_2_), .Y(n261) );
  NAND2X0_HVT U256 ( .A1(srstn), .A2(n245), .Y(net21993) );
  NAND4X0_HVT U257 ( .A1(sram_waddr[2]), .A2(sram_waddr[0]), .A3(sram_waddr[1]), .A4(sram_waddr[3]), .Y(n249) );
  NAND2X0_HVT U258 ( .A1(sram_waddr[4]), .A2(n247), .Y(n248) );
  OA221X1_HVT U259 ( .A1(sram_waddr[5]), .A2(n246), .A3(n70), .A4(n248), .A5(
        n252), .Y(net21999) );
  NAND3X0_HVT U260 ( .A1(sram_waddr[2]), .A2(sram_waddr[0]), .A3(sram_waddr[1]), .Y(n250) );
  OA221X1_HVT U261 ( .A1(sram_waddr[1]), .A2(sram_waddr[0]), .A3(n251), .A4(
        n253), .A5(n252), .Y(net22013) );
  AND2X1_HVT U262 ( .A1(n253), .A2(n252), .Y(net22016) );
  NAND2X0_HVT U263 ( .A1(n42), .A2(n48), .Y(n256) );
  NAND2X0_HVT U264 ( .A1(n255), .A2(n254), .Y(net22026) );
  NAND2X0_HVT U265 ( .A1(n55), .A2(n54), .Y(n257) );
  AND3X1_HVT U266 ( .A1(n259), .A2(n258), .A3(n61), .Y(n129) );
  AND2X1_HVT U267 ( .A1(bytemask_sel[1]), .A2(n49), .Y(sram_bytemask[1]) );
  NAND3X0_HVT U268 ( .A1(n55), .A2(n54), .A3(n260), .Y(sram_write_enable_e0)
         );
  NAND3X0_HVT U269 ( .A1(n54), .A2(n260), .A3(n42), .Y(sram_write_enable_e1)
         );
  NAND3X0_HVT U270 ( .A1(n55), .A2(n260), .A3(n48), .Y(sram_write_enable_e2)
         );
  NAND3X0_HVT U271 ( .A1(n260), .A2(n42), .A3(n48), .Y(sram_write_enable_e3)
         );
endmodule


module fc_data_reg ( clk, srstn, sram_rdata_c0, sram_rdata_c1, sram_rdata_c2, 
        sram_rdata_c3, sram_rdata_c4, sram_rdata_d0, sram_rdata_d1, 
        sram_rdata_d2, sram_rdata_d3, sram_rdata_d4, sram_rdata_e0, 
        sram_rdata_e1, sram_rdata_e2, sram_rdata_e3, sram_rdata_e4, sram_sel, 
        src_window );
  input [31:0] sram_rdata_c0;
  input [31:0] sram_rdata_c1;
  input [31:0] sram_rdata_c2;
  input [31:0] sram_rdata_c3;
  input [31:0] sram_rdata_c4;
  input [31:0] sram_rdata_d0;
  input [31:0] sram_rdata_d1;
  input [31:0] sram_rdata_d2;
  input [31:0] sram_rdata_d3;
  input [31:0] sram_rdata_d4;
  input [31:0] sram_rdata_e0;
  input [31:0] sram_rdata_e1;
  input [31:0] sram_rdata_e2;
  input [31:0] sram_rdata_e3;
  input [31:0] sram_rdata_e4;
  input [1:0] sram_sel;
  output [159:0] src_window;
  input clk, srstn;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44;
  wire   [159:0] n_src_box;

  DFFSSRX1_HVT src_box_reg_159_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[159]), 
        .CLK(clk), .Q(src_window[159]) );
  DFFSSRX1_HVT src_box_reg_158_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[158]), 
        .CLK(clk), .Q(src_window[158]) );
  DFFSSRX1_HVT src_box_reg_157_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[157]), 
        .CLK(clk), .Q(src_window[157]) );
  DFFSSRX1_HVT src_box_reg_156_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[156]), 
        .CLK(clk), .Q(src_window[156]) );
  DFFSSRX1_HVT src_box_reg_155_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[155]), 
        .CLK(clk), .Q(src_window[155]) );
  DFFSSRX1_HVT src_box_reg_154_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[154]), 
        .CLK(clk), .Q(src_window[154]) );
  DFFSSRX1_HVT src_box_reg_153_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[153]), 
        .CLK(clk), .Q(src_window[153]) );
  DFFSSRX1_HVT src_box_reg_152_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[152]), 
        .CLK(clk), .Q(src_window[152]) );
  DFFSSRX1_HVT src_box_reg_151_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[151]), 
        .CLK(clk), .Q(src_window[151]) );
  DFFSSRX1_HVT src_box_reg_150_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[150]), 
        .CLK(clk), .Q(src_window[150]) );
  DFFSSRX1_HVT src_box_reg_149_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[149]), 
        .CLK(clk), .Q(src_window[149]) );
  DFFSSRX1_HVT src_box_reg_148_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[148]), 
        .CLK(clk), .Q(src_window[148]) );
  DFFSSRX1_HVT src_box_reg_147_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[147]), 
        .CLK(clk), .Q(src_window[147]) );
  DFFSSRX1_HVT src_box_reg_146_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[146]), 
        .CLK(clk), .Q(src_window[146]) );
  DFFSSRX1_HVT src_box_reg_145_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[145]), 
        .CLK(clk), .Q(src_window[145]) );
  DFFSSRX1_HVT src_box_reg_144_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[144]), 
        .CLK(clk), .Q(src_window[144]) );
  DFFSSRX1_HVT src_box_reg_143_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[143]), 
        .CLK(clk), .Q(src_window[143]) );
  DFFSSRX1_HVT src_box_reg_142_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[142]), 
        .CLK(clk), .Q(src_window[142]) );
  DFFSSRX1_HVT src_box_reg_141_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[141]), 
        .CLK(clk), .Q(src_window[141]) );
  DFFSSRX1_HVT src_box_reg_140_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[140]), 
        .CLK(clk), .Q(src_window[140]) );
  DFFSSRX1_HVT src_box_reg_139_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[139]), 
        .CLK(clk), .Q(src_window[139]) );
  DFFSSRX1_HVT src_box_reg_138_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[138]), 
        .CLK(clk), .Q(src_window[138]) );
  DFFSSRX1_HVT src_box_reg_137_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[137]), 
        .CLK(clk), .Q(src_window[137]) );
  DFFSSRX1_HVT src_box_reg_136_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[136]), 
        .CLK(clk), .Q(src_window[136]) );
  DFFSSRX1_HVT src_box_reg_135_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[135]), 
        .CLK(clk), .Q(src_window[135]) );
  DFFSSRX1_HVT src_box_reg_134_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[134]), 
        .CLK(clk), .Q(src_window[134]) );
  DFFSSRX1_HVT src_box_reg_133_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[133]), 
        .CLK(clk), .Q(src_window[133]) );
  DFFSSRX1_HVT src_box_reg_132_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[132]), 
        .CLK(clk), .Q(src_window[132]) );
  DFFSSRX1_HVT src_box_reg_131_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[131]), 
        .CLK(clk), .Q(src_window[131]) );
  DFFSSRX1_HVT src_box_reg_130_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[130]), 
        .CLK(clk), .Q(src_window[130]) );
  DFFSSRX1_HVT src_box_reg_129_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[129]), 
        .CLK(clk), .Q(src_window[129]) );
  DFFSSRX1_HVT src_box_reg_128_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[128]), 
        .CLK(clk), .Q(src_window[128]) );
  DFFSSRX1_HVT src_box_reg_127_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[127]), 
        .CLK(clk), .Q(src_window[127]) );
  DFFSSRX1_HVT src_box_reg_126_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[126]), 
        .CLK(clk), .Q(src_window[126]) );
  DFFSSRX1_HVT src_box_reg_125_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[125]), 
        .CLK(clk), .Q(src_window[125]) );
  DFFSSRX1_HVT src_box_reg_124_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[124]), 
        .CLK(clk), .Q(src_window[124]) );
  DFFSSRX1_HVT src_box_reg_123_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[123]), 
        .CLK(clk), .Q(src_window[123]) );
  DFFSSRX1_HVT src_box_reg_122_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[122]), 
        .CLK(clk), .Q(src_window[122]) );
  DFFSSRX1_HVT src_box_reg_121_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[121]), 
        .CLK(clk), .Q(src_window[121]) );
  DFFSSRX1_HVT src_box_reg_120_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[120]), 
        .CLK(clk), .Q(src_window[120]) );
  DFFSSRX1_HVT src_box_reg_119_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[119]), 
        .CLK(clk), .Q(src_window[119]) );
  DFFSSRX1_HVT src_box_reg_118_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[118]), 
        .CLK(clk), .Q(src_window[118]) );
  DFFSSRX1_HVT src_box_reg_117_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[117]), 
        .CLK(clk), .Q(src_window[117]) );
  DFFSSRX1_HVT src_box_reg_116_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[116]), 
        .CLK(clk), .Q(src_window[116]) );
  DFFSSRX1_HVT src_box_reg_115_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[115]), 
        .CLK(clk), .Q(src_window[115]) );
  DFFSSRX1_HVT src_box_reg_114_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[114]), 
        .CLK(clk), .Q(src_window[114]) );
  DFFSSRX1_HVT src_box_reg_113_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[113]), 
        .CLK(clk), .Q(src_window[113]) );
  DFFSSRX1_HVT src_box_reg_112_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[112]), 
        .CLK(clk), .Q(src_window[112]) );
  DFFSSRX1_HVT src_box_reg_111_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[111]), 
        .CLK(clk), .Q(src_window[111]) );
  DFFSSRX1_HVT src_box_reg_110_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[110]), 
        .CLK(clk), .Q(src_window[110]) );
  DFFSSRX1_HVT src_box_reg_109_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[109]), 
        .CLK(clk), .Q(src_window[109]) );
  DFFSSRX1_HVT src_box_reg_108_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[108]), 
        .CLK(clk), .Q(src_window[108]) );
  DFFSSRX1_HVT src_box_reg_107_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[107]), 
        .CLK(clk), .Q(src_window[107]) );
  DFFSSRX1_HVT src_box_reg_106_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[106]), 
        .CLK(clk), .Q(src_window[106]) );
  DFFSSRX1_HVT src_box_reg_105_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[105]), 
        .CLK(clk), .Q(src_window[105]) );
  DFFSSRX1_HVT src_box_reg_104_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[104]), 
        .CLK(clk), .Q(src_window[104]) );
  DFFSSRX1_HVT src_box_reg_103_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[103]), 
        .CLK(clk), .Q(src_window[103]) );
  DFFSSRX1_HVT src_box_reg_102_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[102]), 
        .CLK(clk), .Q(src_window[102]) );
  DFFSSRX1_HVT src_box_reg_101_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[101]), 
        .CLK(clk), .Q(src_window[101]) );
  DFFSSRX1_HVT src_box_reg_100_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[100]), 
        .CLK(clk), .Q(src_window[100]) );
  DFFSSRX1_HVT src_box_reg_99_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[99]), 
        .CLK(clk), .Q(src_window[99]) );
  DFFSSRX1_HVT src_box_reg_98_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[98]), 
        .CLK(clk), .Q(src_window[98]) );
  DFFSSRX1_HVT src_box_reg_97_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[97]), 
        .CLK(clk), .Q(src_window[97]) );
  DFFSSRX1_HVT src_box_reg_96_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[96]), 
        .CLK(clk), .Q(src_window[96]) );
  DFFSSRX1_HVT src_box_reg_95_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[95]), 
        .CLK(clk), .Q(src_window[95]) );
  DFFSSRX1_HVT src_box_reg_94_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[94]), 
        .CLK(clk), .Q(src_window[94]) );
  DFFSSRX1_HVT src_box_reg_93_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[93]), 
        .CLK(clk), .Q(src_window[93]) );
  DFFSSRX1_HVT src_box_reg_92_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[92]), 
        .CLK(clk), .Q(src_window[92]) );
  DFFSSRX1_HVT src_box_reg_91_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[91]), 
        .CLK(clk), .Q(src_window[91]) );
  DFFSSRX1_HVT src_box_reg_90_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[90]), 
        .CLK(clk), .Q(src_window[90]) );
  DFFSSRX1_HVT src_box_reg_89_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[89]), 
        .CLK(clk), .Q(src_window[89]) );
  DFFSSRX1_HVT src_box_reg_88_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[88]), 
        .CLK(clk), .Q(src_window[88]) );
  DFFSSRX1_HVT src_box_reg_87_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[87]), 
        .CLK(clk), .Q(src_window[87]) );
  DFFSSRX1_HVT src_box_reg_86_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[86]), 
        .CLK(clk), .Q(src_window[86]) );
  DFFSSRX1_HVT src_box_reg_85_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[85]), 
        .CLK(clk), .Q(src_window[85]) );
  DFFSSRX1_HVT src_box_reg_84_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[84]), 
        .CLK(clk), .Q(src_window[84]) );
  DFFSSRX1_HVT src_box_reg_83_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[83]), 
        .CLK(clk), .Q(src_window[83]) );
  DFFSSRX1_HVT src_box_reg_82_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[82]), 
        .CLK(clk), .Q(src_window[82]) );
  DFFSSRX1_HVT src_box_reg_81_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[81]), 
        .CLK(clk), .Q(src_window[81]) );
  DFFSSRX1_HVT src_box_reg_80_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[80]), 
        .CLK(clk), .Q(src_window[80]) );
  DFFSSRX1_HVT src_box_reg_79_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[79]), 
        .CLK(clk), .Q(src_window[79]) );
  DFFSSRX1_HVT src_box_reg_78_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[78]), 
        .CLK(clk), .Q(src_window[78]) );
  DFFSSRX1_HVT src_box_reg_77_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[77]), 
        .CLK(clk), .Q(src_window[77]) );
  DFFSSRX1_HVT src_box_reg_76_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[76]), 
        .CLK(clk), .Q(src_window[76]) );
  DFFSSRX1_HVT src_box_reg_75_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[75]), 
        .CLK(clk), .Q(src_window[75]) );
  DFFSSRX1_HVT src_box_reg_74_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[74]), 
        .CLK(clk), .Q(src_window[74]) );
  DFFSSRX1_HVT src_box_reg_73_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[73]), 
        .CLK(clk), .Q(src_window[73]) );
  DFFSSRX1_HVT src_box_reg_72_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[72]), 
        .CLK(clk), .Q(src_window[72]) );
  DFFSSRX1_HVT src_box_reg_71_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[71]), 
        .CLK(clk), .Q(src_window[71]) );
  DFFSSRX1_HVT src_box_reg_70_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[70]), 
        .CLK(clk), .Q(src_window[70]) );
  DFFSSRX1_HVT src_box_reg_69_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[69]), 
        .CLK(clk), .Q(src_window[69]) );
  DFFSSRX1_HVT src_box_reg_68_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[68]), 
        .CLK(clk), .Q(src_window[68]) );
  DFFSSRX1_HVT src_box_reg_67_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[67]), 
        .CLK(clk), .Q(src_window[67]) );
  DFFSSRX1_HVT src_box_reg_66_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[66]), 
        .CLK(clk), .Q(src_window[66]) );
  DFFSSRX1_HVT src_box_reg_65_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[65]), 
        .CLK(clk), .Q(src_window[65]) );
  DFFSSRX1_HVT src_box_reg_64_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[64]), 
        .CLK(clk), .Q(src_window[64]) );
  DFFSSRX1_HVT src_box_reg_63_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[63]), 
        .CLK(clk), .Q(src_window[63]) );
  DFFSSRX1_HVT src_box_reg_62_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[62]), 
        .CLK(clk), .Q(src_window[62]) );
  DFFSSRX1_HVT src_box_reg_61_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[61]), 
        .CLK(clk), .Q(src_window[61]) );
  DFFSSRX1_HVT src_box_reg_60_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[60]), 
        .CLK(clk), .Q(src_window[60]) );
  DFFSSRX1_HVT src_box_reg_59_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[59]), 
        .CLK(clk), .Q(src_window[59]) );
  DFFSSRX1_HVT src_box_reg_58_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[58]), 
        .CLK(clk), .Q(src_window[58]) );
  DFFSSRX1_HVT src_box_reg_57_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[57]), 
        .CLK(clk), .Q(src_window[57]) );
  DFFSSRX1_HVT src_box_reg_56_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[56]), 
        .CLK(clk), .Q(src_window[56]) );
  DFFSSRX1_HVT src_box_reg_55_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[55]), 
        .CLK(clk), .Q(src_window[55]) );
  DFFSSRX1_HVT src_box_reg_54_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[54]), 
        .CLK(clk), .Q(src_window[54]) );
  DFFSSRX1_HVT src_box_reg_53_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[53]), 
        .CLK(clk), .Q(src_window[53]) );
  DFFSSRX1_HVT src_box_reg_52_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[52]), 
        .CLK(clk), .Q(src_window[52]) );
  DFFSSRX1_HVT src_box_reg_51_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[51]), 
        .CLK(clk), .Q(src_window[51]) );
  DFFSSRX1_HVT src_box_reg_50_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[50]), 
        .CLK(clk), .Q(src_window[50]) );
  DFFSSRX1_HVT src_box_reg_49_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[49]), 
        .CLK(clk), .Q(src_window[49]) );
  DFFSSRX1_HVT src_box_reg_48_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[48]), 
        .CLK(clk), .Q(src_window[48]) );
  DFFSSRX1_HVT src_box_reg_47_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[47]), 
        .CLK(clk), .Q(src_window[47]) );
  DFFSSRX1_HVT src_box_reg_46_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[46]), 
        .CLK(clk), .Q(src_window[46]) );
  DFFSSRX1_HVT src_box_reg_45_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[45]), 
        .CLK(clk), .Q(src_window[45]) );
  DFFSSRX1_HVT src_box_reg_44_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[44]), 
        .CLK(clk), .Q(src_window[44]) );
  DFFSSRX1_HVT src_box_reg_43_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[43]), 
        .CLK(clk), .Q(src_window[43]) );
  DFFSSRX1_HVT src_box_reg_42_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[42]), 
        .CLK(clk), .Q(src_window[42]) );
  DFFSSRX1_HVT src_box_reg_41_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[41]), 
        .CLK(clk), .Q(src_window[41]) );
  DFFSSRX1_HVT src_box_reg_40_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[40]), 
        .CLK(clk), .Q(src_window[40]) );
  DFFSSRX1_HVT src_box_reg_39_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[39]), 
        .CLK(clk), .Q(src_window[39]) );
  DFFSSRX1_HVT src_box_reg_38_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[38]), 
        .CLK(clk), .Q(src_window[38]) );
  DFFSSRX1_HVT src_box_reg_37_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[37]), 
        .CLK(clk), .Q(src_window[37]) );
  DFFSSRX1_HVT src_box_reg_36_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[36]), 
        .CLK(clk), .Q(src_window[36]) );
  DFFSSRX1_HVT src_box_reg_35_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[35]), 
        .CLK(clk), .Q(src_window[35]) );
  DFFSSRX1_HVT src_box_reg_34_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[34]), 
        .CLK(clk), .Q(src_window[34]) );
  DFFSSRX1_HVT src_box_reg_33_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[33]), 
        .CLK(clk), .Q(src_window[33]) );
  DFFSSRX1_HVT src_box_reg_32_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[32]), 
        .CLK(clk), .Q(src_window[32]) );
  DFFSSRX1_HVT src_box_reg_31_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[31]), 
        .CLK(clk), .Q(src_window[31]) );
  DFFSSRX1_HVT src_box_reg_30_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[30]), 
        .CLK(clk), .Q(src_window[30]) );
  DFFSSRX1_HVT src_box_reg_29_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[29]), 
        .CLK(clk), .Q(src_window[29]) );
  DFFSSRX1_HVT src_box_reg_28_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[28]), 
        .CLK(clk), .Q(src_window[28]) );
  DFFSSRX1_HVT src_box_reg_27_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[27]), 
        .CLK(clk), .Q(src_window[27]) );
  DFFSSRX1_HVT src_box_reg_26_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[26]), 
        .CLK(clk), .Q(src_window[26]) );
  DFFSSRX1_HVT src_box_reg_25_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[25]), 
        .CLK(clk), .Q(src_window[25]) );
  DFFSSRX1_HVT src_box_reg_24_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[24]), 
        .CLK(clk), .Q(src_window[24]) );
  DFFSSRX1_HVT src_box_reg_23_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[23]), 
        .CLK(clk), .Q(src_window[23]) );
  DFFSSRX1_HVT src_box_reg_22_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[22]), 
        .CLK(clk), .Q(src_window[22]) );
  DFFSSRX1_HVT src_box_reg_21_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[21]), 
        .CLK(clk), .Q(src_window[21]) );
  DFFSSRX1_HVT src_box_reg_20_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[20]), 
        .CLK(clk), .Q(src_window[20]) );
  DFFSSRX1_HVT src_box_reg_19_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[19]), 
        .CLK(clk), .Q(src_window[19]) );
  DFFSSRX1_HVT src_box_reg_18_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[18]), 
        .CLK(clk), .Q(src_window[18]) );
  DFFSSRX1_HVT src_box_reg_17_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[17]), 
        .CLK(clk), .Q(src_window[17]) );
  DFFSSRX1_HVT src_box_reg_16_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[16]), 
        .CLK(clk), .Q(src_window[16]) );
  DFFSSRX1_HVT src_box_reg_15_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[15]), 
        .CLK(clk), .Q(src_window[15]) );
  DFFSSRX1_HVT src_box_reg_14_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[14]), 
        .CLK(clk), .Q(src_window[14]) );
  DFFSSRX1_HVT src_box_reg_13_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[13]), 
        .CLK(clk), .Q(src_window[13]) );
  DFFSSRX1_HVT src_box_reg_12_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[12]), 
        .CLK(clk), .Q(src_window[12]) );
  DFFSSRX1_HVT src_box_reg_11_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[11]), 
        .CLK(clk), .Q(src_window[11]) );
  DFFSSRX1_HVT src_box_reg_10_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[10]), 
        .CLK(clk), .Q(src_window[10]) );
  DFFSSRX1_HVT src_box_reg_9_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[9]), 
        .CLK(clk), .Q(src_window[9]) );
  DFFSSRX1_HVT src_box_reg_8_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[8]), 
        .CLK(clk), .Q(src_window[8]) );
  DFFSSRX1_HVT src_box_reg_7_ ( .D(1'b0), .SETB(n27), .RSTB(n_src_box[7]), 
        .CLK(clk), .Q(src_window[7]) );
  DFFSSRX1_HVT src_box_reg_6_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[6]), 
        .CLK(clk), .Q(src_window[6]) );
  DFFSSRX1_HVT src_box_reg_5_ ( .D(1'b0), .SETB(n1), .RSTB(n_src_box[5]), 
        .CLK(clk), .Q(src_window[5]) );
  DFFSSRX1_HVT src_box_reg_4_ ( .D(1'b0), .SETB(n30), .RSTB(n_src_box[4]), 
        .CLK(clk), .Q(src_window[4]) );
  DFFSSRX1_HVT src_box_reg_3_ ( .D(1'b0), .SETB(n29), .RSTB(n_src_box[3]), 
        .CLK(clk), .Q(src_window[3]) );
  DFFSSRX1_HVT src_box_reg_2_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[2]), 
        .CLK(clk), .Q(src_window[2]) );
  DFFSSRX1_HVT src_box_reg_1_ ( .D(1'b0), .SETB(n44), .RSTB(n_src_box[1]), 
        .CLK(clk), .Q(src_window[1]) );
  DFFSSRX1_HVT src_box_reg_0_ ( .D(1'b0), .SETB(n28), .RSTB(n_src_box[0]), 
        .CLK(clk), .Q(src_window[0]) );
  NAND2X0_HVT U3 ( .A1(n39), .A2(sram_sel[0]), .Y(n43) );
  NAND2X0_HVT U4 ( .A1(n40), .A2(sram_sel[1]), .Y(n42) );
  OR2X1_HVT U5 ( .A1(sram_sel[1]), .A2(sram_sel[0]), .Y(n41) );
  INVX0_HVT U6 ( .A(n43), .Y(n7) );
  INVX0_HVT U7 ( .A(n43), .Y(n6) );
  INVX1_HVT U8 ( .A(n43), .Y(n34) );
  INVX1_HVT U9 ( .A(n42), .Y(n31) );
  INVX2_HVT U10 ( .A(n26), .Y(n1) );
  INVX2_HVT U11 ( .A(srstn), .Y(n44) );
  INVX1_HVT U12 ( .A(n42), .Y(n22) );
  INVX1_HVT U13 ( .A(n42), .Y(n18) );
  INVX1_HVT U14 ( .A(n43), .Y(n9) );
  INVX1_HVT U15 ( .A(n42), .Y(n19) );
  INVX1_HVT U16 ( .A(n42), .Y(n25) );
  INVX1_HVT U17 ( .A(n43), .Y(n10) );
  INVX1_HVT U18 ( .A(n43), .Y(n8) );
  INVX1_HVT U19 ( .A(n43), .Y(n11) );
  INVX1_HVT U20 ( .A(n43), .Y(n4) );
  INVX1_HVT U21 ( .A(n42), .Y(n24) );
  INVX1_HVT U22 ( .A(n42), .Y(n20) );
  INVX1_HVT U23 ( .A(n43), .Y(n5) );
  INVX1_HVT U24 ( .A(n42), .Y(n21) );
  INVX1_HVT U25 ( .A(n42), .Y(n23) );
  INVX1_HVT U26 ( .A(n41), .Y(n17) );
  INVX1_HVT U27 ( .A(n12), .Y(n13) );
  INVX1_HVT U28 ( .A(n41), .Y(n14) );
  INVX1_HVT U29 ( .A(n41), .Y(n15) );
  INVX1_HVT U30 ( .A(n41), .Y(n2) );
  INVX1_HVT U31 ( .A(n41), .Y(n16) );
  INVX1_HVT U32 ( .A(n41), .Y(n3) );
  INVX1_HVT U33 ( .A(n38), .Y(n12) );
  INVX2_HVT U34 ( .A(n26), .Y(n29) );
  INVX2_HVT U35 ( .A(n26), .Y(n27) );
  INVX0_HVT U36 ( .A(sram_sel[0]), .Y(n40) );
  INVX0_HVT U37 ( .A(sram_sel[1]), .Y(n39) );
  INVX2_HVT U38 ( .A(n26), .Y(n30) );
  INVX2_HVT U39 ( .A(n26), .Y(n28) );
  INVX1_HVT U40 ( .A(n43), .Y(n35) );
  INVX2_HVT U41 ( .A(n41), .Y(n37) );
  INVX2_HVT U42 ( .A(n41), .Y(n38) );
  INVX2_HVT U43 ( .A(n41), .Y(n36) );
  INVX1_HVT U44 ( .A(n42), .Y(n33) );
  INVX1_HVT U45 ( .A(n42), .Y(n32) );
  INVX1_HVT U46 ( .A(n44), .Y(n26) );
  AO222X1_HVT U47 ( .A1(n4), .A2(sram_rdata_d4[0]), .A3(n2), .A4(
        sram_rdata_c4[0]), .A5(n31), .A6(sram_rdata_e4[0]), .Y(n_src_box[0])
         );
  AO222X1_HVT U48 ( .A1(n10), .A2(sram_rdata_d4[1]), .A3(n31), .A4(
        sram_rdata_e4[1]), .A5(sram_rdata_c4[1]), .A6(n13), .Y(n_src_box[1])
         );
  AO222X1_HVT U49 ( .A1(n6), .A2(sram_rdata_d4[2]), .A3(n21), .A4(
        sram_rdata_e4[2]), .A5(sram_rdata_c4[2]), .A6(n2), .Y(n_src_box[2]) );
  AO222X1_HVT U50 ( .A1(n8), .A2(sram_rdata_d4[3]), .A3(n31), .A4(
        sram_rdata_e4[3]), .A5(sram_rdata_c4[3]), .A6(n36), .Y(n_src_box[3])
         );
  AO222X1_HVT U51 ( .A1(n8), .A2(sram_rdata_d4[4]), .A3(n32), .A4(
        sram_rdata_e4[4]), .A5(sram_rdata_c4[4]), .A6(n17), .Y(n_src_box[4])
         );
  AO222X1_HVT U52 ( .A1(n34), .A2(sram_rdata_d4[5]), .A3(n21), .A4(
        sram_rdata_e4[5]), .A5(sram_rdata_c4[5]), .A6(n38), .Y(n_src_box[5])
         );
  AO222X1_HVT U53 ( .A1(n9), .A2(sram_rdata_d4[6]), .A3(n24), .A4(
        sram_rdata_e4[6]), .A5(sram_rdata_c4[6]), .A6(n37), .Y(n_src_box[6])
         );
  AO222X1_HVT U54 ( .A1(n6), .A2(sram_rdata_d4[7]), .A3(n23), .A4(
        sram_rdata_e4[7]), .A5(sram_rdata_c4[7]), .A6(n14), .Y(n_src_box[7])
         );
  AO222X1_HVT U55 ( .A1(n11), .A2(sram_rdata_d4[8]), .A3(n22), .A4(
        sram_rdata_e4[8]), .A5(sram_rdata_c4[8]), .A6(n15), .Y(n_src_box[8])
         );
  AO222X1_HVT U56 ( .A1(n35), .A2(sram_rdata_d4[9]), .A3(n18), .A4(
        sram_rdata_e4[9]), .A5(sram_rdata_c4[9]), .A6(n13), .Y(n_src_box[9])
         );
  AO222X1_HVT U57 ( .A1(n4), .A2(sram_rdata_d4[10]), .A3(n20), .A4(
        sram_rdata_e4[10]), .A5(sram_rdata_c4[10]), .A6(n17), .Y(n_src_box[10]) );
  AO222X1_HVT U58 ( .A1(n7), .A2(sram_rdata_d4[11]), .A3(n25), .A4(
        sram_rdata_e4[11]), .A5(sram_rdata_c4[11]), .A6(n16), .Y(n_src_box[11]) );
  AO222X1_HVT U59 ( .A1(n7), .A2(sram_rdata_d4[12]), .A3(n20), .A4(
        sram_rdata_e4[12]), .A5(sram_rdata_c4[12]), .A6(n16), .Y(n_src_box[12]) );
  AO222X1_HVT U60 ( .A1(n7), .A2(sram_rdata_d4[13]), .A3(n33), .A4(
        sram_rdata_e4[13]), .A5(sram_rdata_c4[13]), .A6(n36), .Y(n_src_box[13]) );
  AO222X1_HVT U61 ( .A1(n5), .A2(sram_rdata_d4[14]), .A3(n25), .A4(
        sram_rdata_e4[14]), .A5(sram_rdata_c4[14]), .A6(n3), .Y(n_src_box[14])
         );
  AO222X1_HVT U62 ( .A1(n9), .A2(sram_rdata_d4[15]), .A3(n24), .A4(
        sram_rdata_e4[15]), .A5(sram_rdata_c4[15]), .A6(n16), .Y(n_src_box[15]) );
  AO222X1_HVT U63 ( .A1(n35), .A2(sram_rdata_d4[16]), .A3(n32), .A4(
        sram_rdata_e4[16]), .A5(sram_rdata_c4[16]), .A6(n2), .Y(n_src_box[16])
         );
  AO222X1_HVT U64 ( .A1(n34), .A2(sram_rdata_d4[17]), .A3(n31), .A4(
        sram_rdata_e4[17]), .A5(sram_rdata_c4[17]), .A6(n37), .Y(n_src_box[17]) );
  AO222X1_HVT U65 ( .A1(n5), .A2(sram_rdata_d4[18]), .A3(n33), .A4(
        sram_rdata_e4[18]), .A5(sram_rdata_c4[18]), .A6(n17), .Y(n_src_box[18]) );
  AO222X1_HVT U66 ( .A1(n10), .A2(sram_rdata_d4[19]), .A3(n21), .A4(
        sram_rdata_e4[19]), .A5(sram_rdata_c4[19]), .A6(n37), .Y(n_src_box[19]) );
  AO222X1_HVT U67 ( .A1(n8), .A2(sram_rdata_d4[20]), .A3(n18), .A4(
        sram_rdata_e4[20]), .A5(sram_rdata_c4[20]), .A6(n14), .Y(n_src_box[20]) );
  AO222X1_HVT U68 ( .A1(n6), .A2(sram_rdata_d4[21]), .A3(n33), .A4(
        sram_rdata_e4[21]), .A5(sram_rdata_c4[21]), .A6(n36), .Y(n_src_box[21]) );
  AO222X1_HVT U69 ( .A1(n34), .A2(sram_rdata_d4[22]), .A3(n24), .A4(
        sram_rdata_e4[22]), .A5(sram_rdata_c4[22]), .A6(n38), .Y(n_src_box[22]) );
  AO222X1_HVT U70 ( .A1(n10), .A2(sram_rdata_d4[23]), .A3(n22), .A4(
        sram_rdata_e4[23]), .A5(sram_rdata_c4[23]), .A6(n17), .Y(n_src_box[23]) );
  AO222X1_HVT U71 ( .A1(n5), .A2(sram_rdata_d4[24]), .A3(n20), .A4(
        sram_rdata_e4[24]), .A5(sram_rdata_c4[24]), .A6(n38), .Y(n_src_box[24]) );
  AO222X1_HVT U72 ( .A1(n5), .A2(sram_rdata_d4[25]), .A3(n25), .A4(
        sram_rdata_e4[25]), .A5(sram_rdata_c4[25]), .A6(n17), .Y(n_src_box[25]) );
  AO222X1_HVT U73 ( .A1(n7), .A2(sram_rdata_d4[26]), .A3(n24), .A4(
        sram_rdata_e4[26]), .A5(sram_rdata_c4[26]), .A6(n3), .Y(n_src_box[26])
         );
  AO222X1_HVT U74 ( .A1(n10), .A2(sram_rdata_d4[27]), .A3(n21), .A4(
        sram_rdata_e4[27]), .A5(sram_rdata_c4[27]), .A6(n15), .Y(n_src_box[27]) );
  AO222X1_HVT U75 ( .A1(n9), .A2(sram_rdata_d4[28]), .A3(n21), .A4(
        sram_rdata_e4[28]), .A5(sram_rdata_c4[28]), .A6(n13), .Y(n_src_box[28]) );
  AO222X1_HVT U76 ( .A1(n34), .A2(sram_rdata_d4[29]), .A3(n18), .A4(
        sram_rdata_e4[29]), .A5(sram_rdata_c4[29]), .A6(n38), .Y(n_src_box[29]) );
  AO222X1_HVT U77 ( .A1(n5), .A2(sram_rdata_d4[30]), .A3(n25), .A4(
        sram_rdata_e4[30]), .A5(sram_rdata_c4[30]), .A6(n2), .Y(n_src_box[30])
         );
  AO222X1_HVT U78 ( .A1(n35), .A2(sram_rdata_d4[31]), .A3(n23), .A4(
        sram_rdata_e4[31]), .A5(sram_rdata_c4[31]), .A6(n15), .Y(n_src_box[31]) );
  AO222X1_HVT U79 ( .A1(n9), .A2(sram_rdata_d3[0]), .A3(n22), .A4(
        sram_rdata_e3[0]), .A5(sram_rdata_c3[0]), .A6(n13), .Y(n_src_box[32])
         );
  AO222X1_HVT U80 ( .A1(n35), .A2(sram_rdata_d3[1]), .A3(n21), .A4(
        sram_rdata_e3[1]), .A5(sram_rdata_c3[1]), .A6(n14), .Y(n_src_box[33])
         );
  AO222X1_HVT U81 ( .A1(n11), .A2(sram_rdata_d3[2]), .A3(n33), .A4(
        sram_rdata_e3[2]), .A5(sram_rdata_c3[2]), .A6(n14), .Y(n_src_box[34])
         );
  AO222X1_HVT U82 ( .A1(n4), .A2(sram_rdata_d3[3]), .A3(n22), .A4(
        sram_rdata_e3[3]), .A5(sram_rdata_c3[3]), .A6(n14), .Y(n_src_box[35])
         );
  AO222X1_HVT U83 ( .A1(n6), .A2(sram_rdata_d3[4]), .A3(n32), .A4(
        sram_rdata_e3[4]), .A5(sram_rdata_c3[4]), .A6(n14), .Y(n_src_box[36])
         );
  AO222X1_HVT U84 ( .A1(n6), .A2(sram_rdata_d3[5]), .A3(n31), .A4(
        sram_rdata_e3[5]), .A5(sram_rdata_c3[5]), .A6(n36), .Y(n_src_box[37])
         );
  AO222X1_HVT U85 ( .A1(n4), .A2(sram_rdata_d3[6]), .A3(n32), .A4(
        sram_rdata_e3[6]), .A5(sram_rdata_c3[6]), .A6(n2), .Y(n_src_box[38])
         );
  AO222X1_HVT U86 ( .A1(n11), .A2(sram_rdata_d3[7]), .A3(n25), .A4(
        sram_rdata_e3[7]), .A5(sram_rdata_c3[7]), .A6(n37), .Y(n_src_box[39])
         );
  AO222X1_HVT U87 ( .A1(n4), .A2(sram_rdata_d3[8]), .A3(n18), .A4(
        sram_rdata_e3[8]), .A5(sram_rdata_c3[8]), .A6(n3), .Y(n_src_box[40])
         );
  AO222X1_HVT U88 ( .A1(n34), .A2(sram_rdata_d3[9]), .A3(n31), .A4(
        sram_rdata_e3[9]), .A5(sram_rdata_c3[9]), .A6(n37), .Y(n_src_box[41])
         );
  AO222X1_HVT U89 ( .A1(n9), .A2(sram_rdata_d3[10]), .A3(n18), .A4(
        sram_rdata_e3[10]), .A5(sram_rdata_c3[10]), .A6(n37), .Y(n_src_box[42]) );
  AO222X1_HVT U90 ( .A1(n11), .A2(sram_rdata_d3[11]), .A3(n32), .A4(
        sram_rdata_e3[11]), .A5(sram_rdata_c3[11]), .A6(n38), .Y(n_src_box[43]) );
  AO222X1_HVT U91 ( .A1(n10), .A2(sram_rdata_d3[12]), .A3(n31), .A4(
        sram_rdata_e3[12]), .A5(sram_rdata_c3[12]), .A6(n14), .Y(n_src_box[44]) );
  AO222X1_HVT U92 ( .A1(n7), .A2(sram_rdata_d3[13]), .A3(n25), .A4(
        sram_rdata_e3[13]), .A5(sram_rdata_c3[13]), .A6(n15), .Y(n_src_box[45]) );
  AO222X1_HVT U93 ( .A1(n34), .A2(sram_rdata_d3[14]), .A3(n21), .A4(
        sram_rdata_e3[14]), .A5(sram_rdata_c3[14]), .A6(n37), .Y(n_src_box[46]) );
  AO222X1_HVT U94 ( .A1(n8), .A2(sram_rdata_d3[15]), .A3(n23), .A4(
        sram_rdata_e3[15]), .A5(sram_rdata_c3[15]), .A6(n15), .Y(n_src_box[47]) );
  AO222X1_HVT U95 ( .A1(n5), .A2(sram_rdata_d3[16]), .A3(n22), .A4(
        sram_rdata_e3[16]), .A5(sram_rdata_c3[16]), .A6(n17), .Y(n_src_box[48]) );
  AO222X1_HVT U96 ( .A1(n6), .A2(sram_rdata_d3[17]), .A3(n18), .A4(
        sram_rdata_e3[17]), .A5(sram_rdata_c3[17]), .A6(n2), .Y(n_src_box[49])
         );
  AO222X1_HVT U97 ( .A1(n7), .A2(sram_rdata_d3[18]), .A3(n18), .A4(
        sram_rdata_e3[18]), .A5(sram_rdata_c3[18]), .A6(n2), .Y(n_src_box[50])
         );
  AO222X1_HVT U98 ( .A1(n8), .A2(sram_rdata_d3[19]), .A3(n33), .A4(
        sram_rdata_e3[19]), .A5(sram_rdata_c3[19]), .A6(n17), .Y(n_src_box[51]) );
  AO222X1_HVT U99 ( .A1(n10), .A2(sram_rdata_d3[20]), .A3(n25), .A4(
        sram_rdata_e3[20]), .A5(sram_rdata_c3[20]), .A6(n16), .Y(n_src_box[52]) );
  AO222X1_HVT U100 ( .A1(n34), .A2(sram_rdata_d3[21]), .A3(n19), .A4(
        sram_rdata_e3[21]), .A5(sram_rdata_c3[21]), .A6(n38), .Y(n_src_box[53]) );
  AO222X1_HVT U101 ( .A1(n10), .A2(sram_rdata_d3[22]), .A3(n25), .A4(
        sram_rdata_e3[22]), .A5(sram_rdata_c3[22]), .A6(n15), .Y(n_src_box[54]) );
  AO222X1_HVT U102 ( .A1(n7), .A2(sram_rdata_d3[23]), .A3(n32), .A4(
        sram_rdata_e3[23]), .A5(sram_rdata_c3[23]), .A6(n16), .Y(n_src_box[55]) );
  AO222X1_HVT U103 ( .A1(n11), .A2(sram_rdata_d3[24]), .A3(n18), .A4(
        sram_rdata_e3[24]), .A5(sram_rdata_c3[24]), .A6(n16), .Y(n_src_box[56]) );
  AO222X1_HVT U104 ( .A1(n35), .A2(sram_rdata_d3[25]), .A3(n19), .A4(
        sram_rdata_e3[25]), .A5(sram_rdata_c3[25]), .A6(n36), .Y(n_src_box[57]) );
  AO222X1_HVT U105 ( .A1(n9), .A2(sram_rdata_d3[26]), .A3(n19), .A4(
        sram_rdata_e3[26]), .A5(sram_rdata_c3[26]), .A6(n15), .Y(n_src_box[58]) );
  AO222X1_HVT U106 ( .A1(n6), .A2(sram_rdata_d3[27]), .A3(n23), .A4(
        sram_rdata_e3[27]), .A5(sram_rdata_c3[27]), .A6(n16), .Y(n_src_box[59]) );
  AO222X1_HVT U107 ( .A1(n4), .A2(sram_rdata_d3[28]), .A3(n19), .A4(
        sram_rdata_e3[28]), .A5(sram_rdata_c3[28]), .A6(n36), .Y(n_src_box[60]) );
  AO222X1_HVT U108 ( .A1(n34), .A2(sram_rdata_d3[29]), .A3(n22), .A4(
        sram_rdata_e3[29]), .A5(sram_rdata_c3[29]), .A6(n36), .Y(n_src_box[61]) );
  AO222X1_HVT U109 ( .A1(n6), .A2(sram_rdata_d3[30]), .A3(n22), .A4(
        sram_rdata_e3[30]), .A5(sram_rdata_c3[30]), .A6(n3), .Y(n_src_box[62])
         );
  AO222X1_HVT U110 ( .A1(n9), .A2(sram_rdata_d3[31]), .A3(n23), .A4(
        sram_rdata_e3[31]), .A5(sram_rdata_c3[31]), .A6(n3), .Y(n_src_box[63])
         );
  AO222X1_HVT U111 ( .A1(n5), .A2(sram_rdata_d2[0]), .A3(n22), .A4(
        sram_rdata_e2[0]), .A5(sram_rdata_c2[0]), .A6(n2), .Y(n_src_box[64])
         );
  AO222X1_HVT U112 ( .A1(n35), .A2(sram_rdata_d2[1]), .A3(n31), .A4(
        sram_rdata_e2[1]), .A5(sram_rdata_c2[1]), .A6(n37), .Y(n_src_box[65])
         );
  AO222X1_HVT U113 ( .A1(n4), .A2(sram_rdata_d2[2]), .A3(n32), .A4(
        sram_rdata_e2[2]), .A5(sram_rdata_c2[2]), .A6(n38), .Y(n_src_box[66])
         );
  AO222X1_HVT U114 ( .A1(n8), .A2(sram_rdata_d2[3]), .A3(n31), .A4(
        sram_rdata_e2[3]), .A5(sram_rdata_c2[3]), .A6(n37), .Y(n_src_box[67])
         );
  AO222X1_HVT U115 ( .A1(n8), .A2(sram_rdata_d2[4]), .A3(n19), .A4(
        sram_rdata_e2[4]), .A5(sram_rdata_c2[4]), .A6(n15), .Y(n_src_box[68])
         );
  AO222X1_HVT U116 ( .A1(n6), .A2(sram_rdata_d2[5]), .A3(n32), .A4(
        sram_rdata_e2[5]), .A5(sram_rdata_c2[5]), .A6(n15), .Y(n_src_box[69])
         );
  AO222X1_HVT U117 ( .A1(n34), .A2(sram_rdata_d2[6]), .A3(n32), .A4(
        sram_rdata_e2[6]), .A5(sram_rdata_c2[6]), .A6(n38), .Y(n_src_box[70])
         );
  AO222X1_HVT U118 ( .A1(n8), .A2(sram_rdata_d2[7]), .A3(n20), .A4(
        sram_rdata_e2[7]), .A5(sram_rdata_c2[7]), .A6(n17), .Y(n_src_box[71])
         );
  AO222X1_HVT U119 ( .A1(n7), .A2(sram_rdata_d2[8]), .A3(n22), .A4(
        sram_rdata_e2[8]), .A5(sram_rdata_c2[8]), .A6(n13), .Y(n_src_box[72])
         );
  AO222X1_HVT U120 ( .A1(n5), .A2(sram_rdata_d2[9]), .A3(n33), .A4(
        sram_rdata_e2[9]), .A5(sram_rdata_c2[9]), .A6(n14), .Y(n_src_box[73])
         );
  AO222X1_HVT U121 ( .A1(n6), .A2(sram_rdata_d2[10]), .A3(n25), .A4(
        sram_rdata_e2[10]), .A5(sram_rdata_c2[10]), .A6(n2), .Y(n_src_box[74])
         );
  AO222X1_HVT U122 ( .A1(n10), .A2(sram_rdata_d2[11]), .A3(n20), .A4(
        sram_rdata_e2[11]), .A5(sram_rdata_c2[11]), .A6(n38), .Y(n_src_box[75]) );
  AO222X1_HVT U123 ( .A1(n11), .A2(sram_rdata_d2[12]), .A3(n18), .A4(
        sram_rdata_e2[12]), .A5(sram_rdata_c2[12]), .A6(n14), .Y(n_src_box[76]) );
  AO222X1_HVT U124 ( .A1(n6), .A2(sram_rdata_d2[13]), .A3(n20), .A4(
        sram_rdata_e2[13]), .A5(sram_rdata_c2[13]), .A6(n38), .Y(n_src_box[77]) );
  AO222X1_HVT U125 ( .A1(n4), .A2(sram_rdata_d2[14]), .A3(n24), .A4(
        sram_rdata_e2[14]), .A5(sram_rdata_c2[14]), .A6(n16), .Y(n_src_box[78]) );
  AO222X1_HVT U126 ( .A1(n35), .A2(sram_rdata_d2[15]), .A3(n20), .A4(
        sram_rdata_e2[15]), .A5(sram_rdata_c2[15]), .A6(n17), .Y(n_src_box[79]) );
  AO222X1_HVT U127 ( .A1(n9), .A2(sram_rdata_d2[16]), .A3(n23), .A4(
        sram_rdata_e2[16]), .A5(sram_rdata_c2[16]), .A6(n13), .Y(n_src_box[80]) );
  AO222X1_HVT U128 ( .A1(n35), .A2(sram_rdata_d2[17]), .A3(n18), .A4(
        sram_rdata_e2[17]), .A5(sram_rdata_c2[17]), .A6(n3), .Y(n_src_box[81])
         );
  AO222X1_HVT U129 ( .A1(n8), .A2(sram_rdata_d2[18]), .A3(n22), .A4(
        sram_rdata_e2[18]), .A5(sram_rdata_c2[18]), .A6(n16), .Y(n_src_box[82]) );
  AO222X1_HVT U130 ( .A1(n9), .A2(sram_rdata_d2[19]), .A3(n24), .A4(
        sram_rdata_e2[19]), .A5(sram_rdata_c2[19]), .A6(n14), .Y(n_src_box[83]) );
  AO222X1_HVT U131 ( .A1(n6), .A2(sram_rdata_d2[20]), .A3(n33), .A4(
        sram_rdata_e2[20]), .A5(sram_rdata_c2[20]), .A6(n36), .Y(n_src_box[84]) );
  AO222X1_HVT U132 ( .A1(n34), .A2(sram_rdata_d2[21]), .A3(n19), .A4(
        sram_rdata_e2[21]), .A5(sram_rdata_c2[21]), .A6(n36), .Y(n_src_box[85]) );
  AO222X1_HVT U133 ( .A1(n5), .A2(sram_rdata_d2[22]), .A3(n33), .A4(
        sram_rdata_e2[22]), .A5(sram_rdata_c2[22]), .A6(n3), .Y(n_src_box[86])
         );
  AO222X1_HVT U134 ( .A1(n11), .A2(sram_rdata_d2[23]), .A3(n25), .A4(
        sram_rdata_e2[23]), .A5(sram_rdata_c2[23]), .A6(n14), .Y(n_src_box[87]) );
  AO222X1_HVT U135 ( .A1(n4), .A2(sram_rdata_d2[24]), .A3(n20), .A4(
        sram_rdata_e2[24]), .A5(sram_rdata_c2[24]), .A6(n3), .Y(n_src_box[88])
         );
  AO222X1_HVT U136 ( .A1(n35), .A2(sram_rdata_d2[25]), .A3(n31), .A4(
        sram_rdata_e2[25]), .A5(sram_rdata_c2[25]), .A6(n37), .Y(n_src_box[89]) );
  AO222X1_HVT U137 ( .A1(n10), .A2(sram_rdata_d2[26]), .A3(n21), .A4(
        sram_rdata_e2[26]), .A5(sram_rdata_c2[26]), .A6(n37), .Y(n_src_box[90]) );
  AO222X1_HVT U138 ( .A1(n9), .A2(sram_rdata_d2[27]), .A3(n23), .A4(
        sram_rdata_e2[27]), .A5(sram_rdata_c2[27]), .A6(n38), .Y(n_src_box[91]) );
  AO222X1_HVT U139 ( .A1(n10), .A2(sram_rdata_d2[28]), .A3(n31), .A4(
        sram_rdata_e2[28]), .A5(sram_rdata_c2[28]), .A6(n3), .Y(n_src_box[92])
         );
  AO222X1_HVT U140 ( .A1(n7), .A2(sram_rdata_d2[29]), .A3(n22), .A4(
        sram_rdata_e2[29]), .A5(sram_rdata_c2[29]), .A6(n36), .Y(n_src_box[93]) );
  AO222X1_HVT U141 ( .A1(n34), .A2(sram_rdata_d2[30]), .A3(n24), .A4(
        sram_rdata_e2[30]), .A5(sram_rdata_c2[30]), .A6(n37), .Y(n_src_box[94]) );
  AO222X1_HVT U142 ( .A1(n11), .A2(sram_rdata_d2[31]), .A3(n24), .A4(
        sram_rdata_e2[31]), .A5(sram_rdata_c2[31]), .A6(n15), .Y(n_src_box[95]) );
  AO222X1_HVT U143 ( .A1(n5), .A2(sram_rdata_d1[0]), .A3(n25), .A4(
        sram_rdata_e1[0]), .A5(sram_rdata_c1[0]), .A6(n16), .Y(n_src_box[96])
         );
  AO222X1_HVT U144 ( .A1(n8), .A2(sram_rdata_d1[1]), .A3(n31), .A4(
        sram_rdata_e1[1]), .A5(sram_rdata_c1[1]), .A6(n13), .Y(n_src_box[97])
         );
  AO222X1_HVT U145 ( .A1(n4), .A2(sram_rdata_d1[2]), .A3(n19), .A4(
        sram_rdata_e1[2]), .A5(sram_rdata_c1[2]), .A6(n2), .Y(n_src_box[98])
         );
  AO222X1_HVT U146 ( .A1(n8), .A2(sram_rdata_d1[3]), .A3(n32), .A4(
        sram_rdata_e1[3]), .A5(sram_rdata_c1[3]), .A6(n17), .Y(n_src_box[99])
         );
  AO222X1_HVT U147 ( .A1(n8), .A2(sram_rdata_d1[4]), .A3(n33), .A4(
        sram_rdata_e1[4]), .A5(sram_rdata_c1[4]), .A6(n3), .Y(n_src_box[100])
         );
  AO222X1_HVT U148 ( .A1(n7), .A2(sram_rdata_d1[5]), .A3(n21), .A4(
        sram_rdata_e1[5]), .A5(sram_rdata_c1[5]), .A6(n38), .Y(n_src_box[101])
         );
  AO222X1_HVT U149 ( .A1(n8), .A2(sram_rdata_d1[6]), .A3(n21), .A4(
        sram_rdata_e1[6]), .A5(sram_rdata_c1[6]), .A6(n17), .Y(n_src_box[102])
         );
  AO222X1_HVT U150 ( .A1(n35), .A2(sram_rdata_d1[7]), .A3(n24), .A4(
        sram_rdata_e1[7]), .A5(sram_rdata_c1[7]), .A6(n14), .Y(n_src_box[103])
         );
  AO222X1_HVT U151 ( .A1(n11), .A2(sram_rdata_d1[8]), .A3(n21), .A4(
        sram_rdata_e1[8]), .A5(sram_rdata_c1[8]), .A6(n2), .Y(n_src_box[104])
         );
  AO222X1_HVT U152 ( .A1(n35), .A2(sram_rdata_d1[9]), .A3(n23), .A4(
        sram_rdata_e1[9]), .A5(sram_rdata_c1[9]), .A6(n16), .Y(n_src_box[105])
         );
  AO222X1_HVT U153 ( .A1(n9), .A2(sram_rdata_d1[10]), .A3(n19), .A4(
        sram_rdata_e1[10]), .A5(sram_rdata_c1[10]), .A6(n17), .Y(
        n_src_box[106]) );
  AO222X1_HVT U154 ( .A1(n11), .A2(sram_rdata_d1[11]), .A3(n25), .A4(
        sram_rdata_e1[11]), .A5(sram_rdata_c1[11]), .A6(n16), .Y(
        n_src_box[107]) );
  AO222X1_HVT U155 ( .A1(n4), .A2(sram_rdata_d1[12]), .A3(n18), .A4(
        sram_rdata_e1[12]), .A5(sram_rdata_c1[12]), .A6(n38), .Y(
        n_src_box[108]) );
  AO222X1_HVT U156 ( .A1(n34), .A2(sram_rdata_d1[13]), .A3(n32), .A4(
        sram_rdata_e1[13]), .A5(sram_rdata_c1[13]), .A6(n36), .Y(
        n_src_box[109]) );
  AO222X1_HVT U157 ( .A1(n7), .A2(sram_rdata_d1[14]), .A3(n23), .A4(
        sram_rdata_e1[14]), .A5(sram_rdata_c1[14]), .A6(n3), .Y(n_src_box[110]) );
  AO222X1_HVT U158 ( .A1(n9), .A2(sram_rdata_d1[15]), .A3(n22), .A4(
        sram_rdata_e1[15]), .A5(sram_rdata_c1[15]), .A6(n37), .Y(
        n_src_box[111]) );
  AO222X1_HVT U159 ( .A1(n4), .A2(sram_rdata_d1[16]), .A3(n33), .A4(
        sram_rdata_e1[16]), .A5(sram_rdata_c1[16]), .A6(n2), .Y(n_src_box[112]) );
  AO222X1_HVT U160 ( .A1(n35), .A2(sram_rdata_d1[17]), .A3(n31), .A4(
        sram_rdata_e1[17]), .A5(sram_rdata_c1[17]), .A6(n2), .Y(n_src_box[113]) );
  AO222X1_HVT U161 ( .A1(n9), .A2(sram_rdata_d1[18]), .A3(n33), .A4(
        sram_rdata_e1[18]), .A5(sram_rdata_c1[18]), .A6(n2), .Y(n_src_box[114]) );
  AO222X1_HVT U162 ( .A1(n10), .A2(sram_rdata_d1[19]), .A3(n20), .A4(
        sram_rdata_e1[19]), .A5(sram_rdata_c1[19]), .A6(n37), .Y(
        n_src_box[115]) );
  AO222X1_HVT U163 ( .A1(n8), .A2(sram_rdata_d1[20]), .A3(n20), .A4(
        sram_rdata_e1[20]), .A5(sram_rdata_c1[20]), .A6(n16), .Y(
        n_src_box[116]) );
  AO222X1_HVT U164 ( .A1(n6), .A2(sram_rdata_d1[21]), .A3(n33), .A4(
        sram_rdata_e1[21]), .A5(sram_rdata_c1[21]), .A6(n37), .Y(
        n_src_box[117]) );
  AO222X1_HVT U165 ( .A1(n34), .A2(sram_rdata_d1[22]), .A3(n23), .A4(
        sram_rdata_e1[22]), .A5(sram_rdata_c1[22]), .A6(n38), .Y(
        n_src_box[118]) );
  AO222X1_HVT U166 ( .A1(n11), .A2(sram_rdata_d1[23]), .A3(n21), .A4(
        sram_rdata_e1[23]), .A5(sram_rdata_c1[23]), .A6(n17), .Y(
        n_src_box[119]) );
  AO222X1_HVT U167 ( .A1(n7), .A2(sram_rdata_d1[24]), .A3(n22), .A4(
        sram_rdata_e1[24]), .A5(sram_rdata_c1[24]), .A6(n14), .Y(
        n_src_box[120]) );
  AO222X1_HVT U168 ( .A1(n4), .A2(sram_rdata_d1[25]), .A3(n24), .A4(
        sram_rdata_e1[25]), .A5(sram_rdata_c1[25]), .A6(n14), .Y(
        n_src_box[121]) );
  AO222X1_HVT U169 ( .A1(n5), .A2(sram_rdata_d1[26]), .A3(n19), .A4(
        sram_rdata_e1[26]), .A5(sram_rdata_c1[26]), .A6(n36), .Y(
        n_src_box[122]) );
  AO222X1_HVT U170 ( .A1(n10), .A2(sram_rdata_d1[27]), .A3(n19), .A4(
        sram_rdata_e1[27]), .A5(sram_rdata_c1[27]), .A6(n15), .Y(
        n_src_box[123]) );
  AO222X1_HVT U171 ( .A1(n9), .A2(sram_rdata_d1[28]), .A3(n19), .A4(
        sram_rdata_e1[28]), .A5(sram_rdata_c1[28]), .A6(n13), .Y(
        n_src_box[124]) );
  AO222X1_HVT U172 ( .A1(n6), .A2(sram_rdata_d1[29]), .A3(n18), .A4(
        sram_rdata_e1[29]), .A5(sram_rdata_c1[29]), .A6(n3), .Y(n_src_box[125]) );
  AO222X1_HVT U173 ( .A1(n4), .A2(sram_rdata_d1[30]), .A3(n23), .A4(
        sram_rdata_e1[30]), .A5(sram_rdata_c1[30]), .A6(n36), .Y(
        n_src_box[126]) );
  AO222X1_HVT U174 ( .A1(n35), .A2(sram_rdata_d1[31]), .A3(n23), .A4(
        sram_rdata_e1[31]), .A5(sram_rdata_c1[31]), .A6(n15), .Y(
        n_src_box[127]) );
  AO222X1_HVT U175 ( .A1(n9), .A2(sram_rdata_d0[0]), .A3(n24), .A4(
        sram_rdata_e0[0]), .A5(sram_rdata_c0[0]), .A6(n13), .Y(n_src_box[128])
         );
  AO222X1_HVT U176 ( .A1(n35), .A2(sram_rdata_d0[1]), .A3(n19), .A4(
        sram_rdata_e0[1]), .A5(sram_rdata_c0[1]), .A6(n36), .Y(n_src_box[129])
         );
  AO222X1_HVT U177 ( .A1(n5), .A2(sram_rdata_d0[2]), .A3(n32), .A4(
        sram_rdata_e0[2]), .A5(sram_rdata_c0[2]), .A6(n14), .Y(n_src_box[130])
         );
  AO222X1_HVT U178 ( .A1(n10), .A2(sram_rdata_d0[3]), .A3(n22), .A4(
        sram_rdata_e0[3]), .A5(sram_rdata_c0[3]), .A6(n14), .Y(n_src_box[131])
         );
  AO222X1_HVT U179 ( .A1(n6), .A2(sram_rdata_d0[4]), .A3(n32), .A4(
        sram_rdata_e0[4]), .A5(sram_rdata_c0[4]), .A6(n37), .Y(n_src_box[132])
         );
  AO222X1_HVT U180 ( .A1(n34), .A2(sram_rdata_d0[5]), .A3(n31), .A4(
        sram_rdata_e0[5]), .A5(sram_rdata_c0[5]), .A6(n38), .Y(n_src_box[133])
         );
  AO222X1_HVT U181 ( .A1(n6), .A2(sram_rdata_d0[6]), .A3(n32), .A4(
        sram_rdata_e0[6]), .A5(sram_rdata_c0[6]), .A6(n36), .Y(n_src_box[134])
         );
  AO222X1_HVT U182 ( .A1(n11), .A2(sram_rdata_d0[7]), .A3(n20), .A4(
        sram_rdata_e0[7]), .A5(sram_rdata_c0[7]), .A6(n13), .Y(n_src_box[135])
         );
  AO222X1_HVT U183 ( .A1(n7), .A2(sram_rdata_d0[8]), .A3(n19), .A4(
        sram_rdata_e0[8]), .A5(sram_rdata_c0[8]), .A6(n3), .Y(n_src_box[136])
         );
  AO222X1_HVT U184 ( .A1(n35), .A2(sram_rdata_d0[9]), .A3(n31), .A4(
        sram_rdata_e0[9]), .A5(sram_rdata_c0[9]), .A6(n2), .Y(n_src_box[137])
         );
  AO222X1_HVT U185 ( .A1(n7), .A2(sram_rdata_d0[10]), .A3(n20), .A4(
        sram_rdata_e0[10]), .A5(sram_rdata_c0[10]), .A6(n3), .Y(n_src_box[138]) );
  AO222X1_HVT U186 ( .A1(n11), .A2(sram_rdata_d0[11]), .A3(n18), .A4(
        sram_rdata_e0[11]), .A5(sram_rdata_c0[11]), .A6(n17), .Y(
        n_src_box[139]) );
  AO222X1_HVT U187 ( .A1(n10), .A2(sram_rdata_d0[12]), .A3(n31), .A4(
        sram_rdata_e0[12]), .A5(sram_rdata_c0[12]), .A6(n15), .Y(
        n_src_box[140]) );
  AO222X1_HVT U188 ( .A1(n7), .A2(sram_rdata_d0[13]), .A3(n23), .A4(
        sram_rdata_e0[13]), .A5(sram_rdata_c0[13]), .A6(n17), .Y(
        n_src_box[141]) );
  AO222X1_HVT U189 ( .A1(n34), .A2(sram_rdata_d0[14]), .A3(n20), .A4(
        sram_rdata_e0[14]), .A5(sram_rdata_c0[14]), .A6(n37), .Y(
        n_src_box[142]) );
  AO222X1_HVT U190 ( .A1(n5), .A2(sram_rdata_d0[15]), .A3(n24), .A4(
        sram_rdata_e0[15]), .A5(sram_rdata_c0[15]), .A6(n15), .Y(
        n_src_box[143]) );
  AO222X1_HVT U191 ( .A1(n5), .A2(sram_rdata_d0[16]), .A3(n24), .A4(
        sram_rdata_e0[16]), .A5(sram_rdata_c0[16]), .A6(n15), .Y(
        n_src_box[144]) );
  AO222X1_HVT U192 ( .A1(n11), .A2(sram_rdata_d0[17]), .A3(n21), .A4(
        sram_rdata_e0[17]), .A5(sram_rdata_c0[17]), .A6(n16), .Y(
        n_src_box[145]) );
  AO222X1_HVT U193 ( .A1(n5), .A2(sram_rdata_d0[18]), .A3(n20), .A4(
        sram_rdata_e0[18]), .A5(sram_rdata_c0[18]), .A6(n36), .Y(
        n_src_box[146]) );
  AO222X1_HVT U194 ( .A1(n8), .A2(sram_rdata_d0[19]), .A3(n33), .A4(
        sram_rdata_e0[19]), .A5(sram_rdata_c0[19]), .A6(n38), .Y(
        n_src_box[147]) );
  AO222X1_HVT U195 ( .A1(n10), .A2(sram_rdata_d0[20]), .A3(n24), .A4(
        sram_rdata_e0[20]), .A5(sram_rdata_c0[20]), .A6(n17), .Y(
        n_src_box[148]) );
  AO222X1_HVT U196 ( .A1(n7), .A2(sram_rdata_d0[21]), .A3(n19), .A4(
        sram_rdata_e0[21]), .A5(sram_rdata_c0[21]), .A6(n3), .Y(n_src_box[149]) );
  AO222X1_HVT U197 ( .A1(n11), .A2(sram_rdata_d0[22]), .A3(n25), .A4(
        sram_rdata_e0[22]), .A5(sram_rdata_c0[22]), .A6(n36), .Y(
        n_src_box[150]) );
  AO222X1_HVT U198 ( .A1(n5), .A2(sram_rdata_d0[23]), .A3(n33), .A4(
        sram_rdata_e0[23]), .A5(sram_rdata_c0[23]), .A6(n3), .Y(n_src_box[151]) );
  AO222X1_HVT U199 ( .A1(n11), .A2(sram_rdata_d0[24]), .A3(n23), .A4(
        sram_rdata_e0[24]), .A5(sram_rdata_c0[24]), .A6(n2), .Y(n_src_box[152]) );
  AO222X1_HVT U200 ( .A1(n35), .A2(sram_rdata_d0[25]), .A3(n18), .A4(
        sram_rdata_e0[25]), .A5(sram_rdata_c0[25]), .A6(n13), .Y(
        n_src_box[153]) );
  AO222X1_HVT U201 ( .A1(n10), .A2(sram_rdata_d0[26]), .A3(n22), .A4(
        sram_rdata_e0[26]), .A5(sram_rdata_c0[26]), .A6(n15), .Y(
        n_src_box[154]) );
  AO222X1_HVT U202 ( .A1(n8), .A2(sram_rdata_d0[27]), .A3(n23), .A4(
        sram_rdata_e0[27]), .A5(sram_rdata_c0[27]), .A6(n16), .Y(
        n_src_box[155]) );
  AO222X1_HVT U203 ( .A1(n4), .A2(sram_rdata_d0[28]), .A3(n21), .A4(
        sram_rdata_e0[28]), .A5(sram_rdata_c0[28]), .A6(n38), .Y(
        n_src_box[156]) );
  AO222X1_HVT U204 ( .A1(n34), .A2(sram_rdata_d0[29]), .A3(n25), .A4(
        sram_rdata_e0[29]), .A5(sram_rdata_c0[29]), .A6(n37), .Y(
        n_src_box[157]) );
  AO222X1_HVT U205 ( .A1(n4), .A2(sram_rdata_d0[30]), .A3(n24), .A4(
        sram_rdata_e0[30]), .A5(sram_rdata_c0[30]), .A6(n36), .Y(
        n_src_box[158]) );
  AO222X1_HVT U206 ( .A1(n9), .A2(sram_rdata_d0[31]), .A3(n25), .A4(
        sram_rdata_e0[31]), .A5(sram_rdata_c0[31]), .A6(n16), .Y(
        n_src_box[159]) );
endmodule


module fc_multiplier_accumulator ( clk, srstn, src_window, sram_rdata_weight, 
        accumulate_reset, data_out );
  input [159:0] src_window;
  input [79:0] sram_rdata_weight;
  output [22:0] data_out;
  input clk, srstn, accumulate_reset;
  wire   DP_OP_102J5_124_3590_n2411, DP_OP_102J5_124_3590_n2379,
         DP_OP_102J5_124_3590_n2378, DP_OP_102J5_124_3590_n2377,
         DP_OP_102J5_124_3590_n2376, DP_OP_102J5_124_3590_n2375,
         DP_OP_102J5_124_3590_n2374, DP_OP_102J5_124_3590_n2373,
         DP_OP_102J5_124_3590_n2372, DP_OP_102J5_124_3590_n2371,
         DP_OP_102J5_124_3590_n2370, DP_OP_102J5_124_3590_n2369,
         DP_OP_102J5_124_3590_n2368, DP_OP_102J5_124_3590_n2367,
         DP_OP_102J5_124_3590_n2366, DP_OP_102J5_124_3590_n2365,
         DP_OP_102J5_124_3590_n2364, DP_OP_102J5_124_3590_n2363,
         DP_OP_102J5_124_3590_n2362, DP_OP_102J5_124_3590_n2361,
         DP_OP_102J5_124_3590_n2360, DP_OP_102J5_124_3590_n2359,
         DP_OP_102J5_124_3590_n2358, DP_OP_102J5_124_3590_n2357,
         DP_OP_102J5_124_3590_n2356, DP_OP_102J5_124_3590_n2355,
         DP_OP_102J5_124_3590_n2354, DP_OP_102J5_124_3590_n2353,
         DP_OP_102J5_124_3590_n2352, DP_OP_102J5_124_3590_n2351,
         DP_OP_102J5_124_3590_n2350, DP_OP_102J5_124_3590_n2349,
         DP_OP_102J5_124_3590_n2348, DP_OP_102J5_124_3590_n2347,
         DP_OP_102J5_124_3590_n2346, DP_OP_102J5_124_3590_n2345,
         DP_OP_102J5_124_3590_n2344, DP_OP_102J5_124_3590_n2343,
         DP_OP_102J5_124_3590_n2342, DP_OP_102J5_124_3590_n2341,
         DP_OP_102J5_124_3590_n2336, DP_OP_102J5_124_3590_n2335,
         DP_OP_102J5_124_3590_n2334, DP_OP_102J5_124_3590_n2333,
         DP_OP_102J5_124_3590_n2332, DP_OP_102J5_124_3590_n2331,
         DP_OP_102J5_124_3590_n2330, DP_OP_102J5_124_3590_n2329,
         DP_OP_102J5_124_3590_n2328, DP_OP_102J5_124_3590_n2327,
         DP_OP_102J5_124_3590_n2326, DP_OP_102J5_124_3590_n2325,
         DP_OP_102J5_124_3590_n2324, DP_OP_102J5_124_3590_n2323,
         DP_OP_102J5_124_3590_n2322, DP_OP_102J5_124_3590_n2321,
         DP_OP_102J5_124_3590_n2320, DP_OP_102J5_124_3590_n2319,
         DP_OP_102J5_124_3590_n2318, DP_OP_102J5_124_3590_n2317,
         DP_OP_102J5_124_3590_n2316, DP_OP_102J5_124_3590_n2315,
         DP_OP_102J5_124_3590_n2314, DP_OP_102J5_124_3590_n2313,
         DP_OP_102J5_124_3590_n2312, DP_OP_102J5_124_3590_n2311,
         DP_OP_102J5_124_3590_n2310, DP_OP_102J5_124_3590_n2309,
         DP_OP_102J5_124_3590_n2308, DP_OP_102J5_124_3590_n2307,
         DP_OP_102J5_124_3590_n2306, DP_OP_102J5_124_3590_n2305,
         DP_OP_102J5_124_3590_n2304, DP_OP_102J5_124_3590_n2303,
         DP_OP_102J5_124_3590_n2302, DP_OP_102J5_124_3590_n2301,
         DP_OP_102J5_124_3590_n2300, DP_OP_102J5_124_3590_n2299,
         DP_OP_102J5_124_3590_n2298, DP_OP_102J5_124_3590_n2297,
         DP_OP_102J5_124_3590_n2292, DP_OP_102J5_124_3590_n2291,
         DP_OP_102J5_124_3590_n2290, DP_OP_102J5_124_3590_n2289,
         DP_OP_102J5_124_3590_n2288, DP_OP_102J5_124_3590_n2287,
         DP_OP_102J5_124_3590_n2286, DP_OP_102J5_124_3590_n2285,
         DP_OP_102J5_124_3590_n2284, DP_OP_102J5_124_3590_n2283,
         DP_OP_102J5_124_3590_n2282, DP_OP_102J5_124_3590_n2281,
         DP_OP_102J5_124_3590_n2280, DP_OP_102J5_124_3590_n2279,
         DP_OP_102J5_124_3590_n2278, DP_OP_102J5_124_3590_n2277,
         DP_OP_102J5_124_3590_n2276, DP_OP_102J5_124_3590_n2275,
         DP_OP_102J5_124_3590_n2274, DP_OP_102J5_124_3590_n2273,
         DP_OP_102J5_124_3590_n2272, DP_OP_102J5_124_3590_n2271,
         DP_OP_102J5_124_3590_n2270, DP_OP_102J5_124_3590_n2269,
         DP_OP_102J5_124_3590_n2268, DP_OP_102J5_124_3590_n2267,
         DP_OP_102J5_124_3590_n2266, DP_OP_102J5_124_3590_n2265,
         DP_OP_102J5_124_3590_n2264, DP_OP_102J5_124_3590_n2263,
         DP_OP_102J5_124_3590_n2262, DP_OP_102J5_124_3590_n2261,
         DP_OP_102J5_124_3590_n2260, DP_OP_102J5_124_3590_n2259,
         DP_OP_102J5_124_3590_n2258, DP_OP_102J5_124_3590_n2257,
         DP_OP_102J5_124_3590_n2256, DP_OP_102J5_124_3590_n2255,
         DP_OP_102J5_124_3590_n2254, DP_OP_102J5_124_3590_n2253,
         DP_OP_102J5_124_3590_n2248, DP_OP_102J5_124_3590_n2247,
         DP_OP_102J5_124_3590_n2246, DP_OP_102J5_124_3590_n2245,
         DP_OP_102J5_124_3590_n2244, DP_OP_102J5_124_3590_n2243,
         DP_OP_102J5_124_3590_n2242, DP_OP_102J5_124_3590_n2241,
         DP_OP_102J5_124_3590_n2240, DP_OP_102J5_124_3590_n2239,
         DP_OP_102J5_124_3590_n2238, DP_OP_102J5_124_3590_n2237,
         DP_OP_102J5_124_3590_n2236, DP_OP_102J5_124_3590_n2235,
         DP_OP_102J5_124_3590_n2234, DP_OP_102J5_124_3590_n2233,
         DP_OP_102J5_124_3590_n2232, DP_OP_102J5_124_3590_n2231,
         DP_OP_102J5_124_3590_n2230, DP_OP_102J5_124_3590_n2229,
         DP_OP_102J5_124_3590_n2228, DP_OP_102J5_124_3590_n2227,
         DP_OP_102J5_124_3590_n2226, DP_OP_102J5_124_3590_n2225,
         DP_OP_102J5_124_3590_n2224, DP_OP_102J5_124_3590_n2223,
         DP_OP_102J5_124_3590_n2222, DP_OP_102J5_124_3590_n2221,
         DP_OP_102J5_124_3590_n2220, DP_OP_102J5_124_3590_n2219,
         DP_OP_102J5_124_3590_n2218, DP_OP_102J5_124_3590_n2217,
         DP_OP_102J5_124_3590_n2216, DP_OP_102J5_124_3590_n2215,
         DP_OP_102J5_124_3590_n2214, DP_OP_102J5_124_3590_n2213,
         DP_OP_102J5_124_3590_n2212, DP_OP_102J5_124_3590_n2211,
         DP_OP_102J5_124_3590_n2210, DP_OP_102J5_124_3590_n2209,
         DP_OP_102J5_124_3590_n2204, DP_OP_102J5_124_3590_n2203,
         DP_OP_102J5_124_3590_n2202, DP_OP_102J5_124_3590_n2201,
         DP_OP_102J5_124_3590_n2200, DP_OP_102J5_124_3590_n2199,
         DP_OP_102J5_124_3590_n2198, DP_OP_102J5_124_3590_n2197,
         DP_OP_102J5_124_3590_n2196, DP_OP_102J5_124_3590_n2195,
         DP_OP_102J5_124_3590_n2194, DP_OP_102J5_124_3590_n2193,
         DP_OP_102J5_124_3590_n2192, DP_OP_102J5_124_3590_n2191,
         DP_OP_102J5_124_3590_n2190, DP_OP_102J5_124_3590_n2189,
         DP_OP_102J5_124_3590_n2188, DP_OP_102J5_124_3590_n2187,
         DP_OP_102J5_124_3590_n2186, DP_OP_102J5_124_3590_n2185,
         DP_OP_102J5_124_3590_n2184, DP_OP_102J5_124_3590_n2183,
         DP_OP_102J5_124_3590_n2182, DP_OP_102J5_124_3590_n2181,
         DP_OP_102J5_124_3590_n2180, DP_OP_102J5_124_3590_n2179,
         DP_OP_102J5_124_3590_n2178, DP_OP_102J5_124_3590_n2177,
         DP_OP_102J5_124_3590_n2176, DP_OP_102J5_124_3590_n2175,
         DP_OP_102J5_124_3590_n2174, DP_OP_102J5_124_3590_n2173,
         DP_OP_102J5_124_3590_n2172, DP_OP_102J5_124_3590_n2171,
         DP_OP_102J5_124_3590_n2170, DP_OP_102J5_124_3590_n2169,
         DP_OP_102J5_124_3590_n2168, DP_OP_102J5_124_3590_n2167,
         DP_OP_102J5_124_3590_n2166, DP_OP_102J5_124_3590_n2165,
         DP_OP_102J5_124_3590_n2160, DP_OP_102J5_124_3590_n2159,
         DP_OP_102J5_124_3590_n2158, DP_OP_102J5_124_3590_n2157,
         DP_OP_102J5_124_3590_n2156, DP_OP_102J5_124_3590_n2155,
         DP_OP_102J5_124_3590_n2154, DP_OP_102J5_124_3590_n2153,
         DP_OP_102J5_124_3590_n2152, DP_OP_102J5_124_3590_n2151,
         DP_OP_102J5_124_3590_n2150, DP_OP_102J5_124_3590_n2149,
         DP_OP_102J5_124_3590_n2148, DP_OP_102J5_124_3590_n2147,
         DP_OP_102J5_124_3590_n2146, DP_OP_102J5_124_3590_n2145,
         DP_OP_102J5_124_3590_n2144, DP_OP_102J5_124_3590_n2143,
         DP_OP_102J5_124_3590_n2142, DP_OP_102J5_124_3590_n2141,
         DP_OP_102J5_124_3590_n2140, DP_OP_102J5_124_3590_n2139,
         DP_OP_102J5_124_3590_n2138, DP_OP_102J5_124_3590_n2137,
         DP_OP_102J5_124_3590_n2136, DP_OP_102J5_124_3590_n2135,
         DP_OP_102J5_124_3590_n2134, DP_OP_102J5_124_3590_n2133,
         DP_OP_102J5_124_3590_n2132, DP_OP_102J5_124_3590_n2131,
         DP_OP_102J5_124_3590_n2130, DP_OP_102J5_124_3590_n2129,
         DP_OP_102J5_124_3590_n2128, DP_OP_102J5_124_3590_n2127,
         DP_OP_102J5_124_3590_n2126, DP_OP_102J5_124_3590_n2125,
         DP_OP_102J5_124_3590_n2124, DP_OP_102J5_124_3590_n2123,
         DP_OP_102J5_124_3590_n2122, DP_OP_102J5_124_3590_n2121,
         DP_OP_102J5_124_3590_n2116, DP_OP_102J5_124_3590_n2115,
         DP_OP_102J5_124_3590_n2114, DP_OP_102J5_124_3590_n2113,
         DP_OP_102J5_124_3590_n2112, DP_OP_102J5_124_3590_n2111,
         DP_OP_102J5_124_3590_n2110, DP_OP_102J5_124_3590_n2109,
         DP_OP_102J5_124_3590_n2108, DP_OP_102J5_124_3590_n2107,
         DP_OP_102J5_124_3590_n2106, DP_OP_102J5_124_3590_n2105,
         DP_OP_102J5_124_3590_n2104, DP_OP_102J5_124_3590_n2103,
         DP_OP_102J5_124_3590_n2102, DP_OP_102J5_124_3590_n2101,
         DP_OP_102J5_124_3590_n2100, DP_OP_102J5_124_3590_n2099,
         DP_OP_102J5_124_3590_n2098, DP_OP_102J5_124_3590_n2097,
         DP_OP_102J5_124_3590_n2096, DP_OP_102J5_124_3590_n2095,
         DP_OP_102J5_124_3590_n2094, DP_OP_102J5_124_3590_n2093,
         DP_OP_102J5_124_3590_n2092, DP_OP_102J5_124_3590_n2091,
         DP_OP_102J5_124_3590_n2090, DP_OP_102J5_124_3590_n2089,
         DP_OP_102J5_124_3590_n2088, DP_OP_102J5_124_3590_n2087,
         DP_OP_102J5_124_3590_n2086, DP_OP_102J5_124_3590_n2085,
         DP_OP_102J5_124_3590_n2084, DP_OP_102J5_124_3590_n2083,
         DP_OP_102J5_124_3590_n2082, DP_OP_102J5_124_3590_n2081,
         DP_OP_102J5_124_3590_n2080, DP_OP_102J5_124_3590_n2079,
         DP_OP_102J5_124_3590_n2078, DP_OP_102J5_124_3590_n2077,
         DP_OP_102J5_124_3590_n2072, DP_OP_102J5_124_3590_n2071,
         DP_OP_102J5_124_3590_n2070, DP_OP_102J5_124_3590_n2069,
         DP_OP_102J5_124_3590_n2068, DP_OP_102J5_124_3590_n2067,
         DP_OP_102J5_124_3590_n2066, DP_OP_102J5_124_3590_n2065,
         DP_OP_102J5_124_3590_n2064, DP_OP_102J5_124_3590_n2063,
         DP_OP_102J5_124_3590_n2062, DP_OP_102J5_124_3590_n2061,
         DP_OP_102J5_124_3590_n2060, DP_OP_102J5_124_3590_n2059,
         DP_OP_102J5_124_3590_n2058, DP_OP_102J5_124_3590_n2057,
         DP_OP_102J5_124_3590_n2056, DP_OP_102J5_124_3590_n2055,
         DP_OP_102J5_124_3590_n2054, DP_OP_102J5_124_3590_n2053,
         DP_OP_102J5_124_3590_n2052, DP_OP_102J5_124_3590_n2051,
         DP_OP_102J5_124_3590_n2050, DP_OP_102J5_124_3590_n2049,
         DP_OP_102J5_124_3590_n2048, DP_OP_102J5_124_3590_n2047,
         DP_OP_102J5_124_3590_n2046, DP_OP_102J5_124_3590_n2045,
         DP_OP_102J5_124_3590_n2044, DP_OP_102J5_124_3590_n2043,
         DP_OP_102J5_124_3590_n2042, DP_OP_102J5_124_3590_n2041,
         DP_OP_102J5_124_3590_n2040, DP_OP_102J5_124_3590_n2039,
         DP_OP_102J5_124_3590_n2038, DP_OP_102J5_124_3590_n2037,
         DP_OP_102J5_124_3590_n2036, DP_OP_102J5_124_3590_n2035,
         DP_OP_102J5_124_3590_n2034, DP_OP_102J5_124_3590_n2033,
         DP_OP_102J5_124_3590_n2028, DP_OP_102J5_124_3590_n2027,
         DP_OP_102J5_124_3590_n2026, DP_OP_102J5_124_3590_n2025,
         DP_OP_102J5_124_3590_n2024, DP_OP_102J5_124_3590_n2023,
         DP_OP_102J5_124_3590_n2022, DP_OP_102J5_124_3590_n2021,
         DP_OP_102J5_124_3590_n2020, DP_OP_102J5_124_3590_n2019,
         DP_OP_102J5_124_3590_n2018, DP_OP_102J5_124_3590_n2017,
         DP_OP_102J5_124_3590_n2016, DP_OP_102J5_124_3590_n2015,
         DP_OP_102J5_124_3590_n2014, DP_OP_102J5_124_3590_n2013,
         DP_OP_102J5_124_3590_n2012, DP_OP_102J5_124_3590_n2011,
         DP_OP_102J5_124_3590_n2010, DP_OP_102J5_124_3590_n2009,
         DP_OP_102J5_124_3590_n2008, DP_OP_102J5_124_3590_n2007,
         DP_OP_102J5_124_3590_n2006, DP_OP_102J5_124_3590_n2005,
         DP_OP_102J5_124_3590_n2004, DP_OP_102J5_124_3590_n2003,
         DP_OP_102J5_124_3590_n2002, DP_OP_102J5_124_3590_n2001,
         DP_OP_102J5_124_3590_n2000, DP_OP_102J5_124_3590_n1999,
         DP_OP_102J5_124_3590_n1998, DP_OP_102J5_124_3590_n1997,
         DP_OP_102J5_124_3590_n1996, DP_OP_102J5_124_3590_n1995,
         DP_OP_102J5_124_3590_n1994, DP_OP_102J5_124_3590_n1993,
         DP_OP_102J5_124_3590_n1992, DP_OP_102J5_124_3590_n1991,
         DP_OP_102J5_124_3590_n1990, DP_OP_102J5_124_3590_n1989,
         DP_OP_102J5_124_3590_n1984, DP_OP_102J5_124_3590_n1983,
         DP_OP_102J5_124_3590_n1982, DP_OP_102J5_124_3590_n1981,
         DP_OP_102J5_124_3590_n1980, DP_OP_102J5_124_3590_n1979,
         DP_OP_102J5_124_3590_n1978, DP_OP_102J5_124_3590_n1977,
         DP_OP_102J5_124_3590_n1976, DP_OP_102J5_124_3590_n1975,
         DP_OP_102J5_124_3590_n1974, DP_OP_102J5_124_3590_n1973,
         DP_OP_102J5_124_3590_n1972, DP_OP_102J5_124_3590_n1971,
         DP_OP_102J5_124_3590_n1970, DP_OP_102J5_124_3590_n1969,
         DP_OP_102J5_124_3590_n1968, DP_OP_102J5_124_3590_n1967,
         DP_OP_102J5_124_3590_n1966, DP_OP_102J5_124_3590_n1965,
         DP_OP_102J5_124_3590_n1964, DP_OP_102J5_124_3590_n1963,
         DP_OP_102J5_124_3590_n1962, DP_OP_102J5_124_3590_n1961,
         DP_OP_102J5_124_3590_n1960, DP_OP_102J5_124_3590_n1959,
         DP_OP_102J5_124_3590_n1958, DP_OP_102J5_124_3590_n1957,
         DP_OP_102J5_124_3590_n1956, DP_OP_102J5_124_3590_n1955,
         DP_OP_102J5_124_3590_n1954, DP_OP_102J5_124_3590_n1953,
         DP_OP_102J5_124_3590_n1952, DP_OP_102J5_124_3590_n1951,
         DP_OP_102J5_124_3590_n1950, DP_OP_102J5_124_3590_n1949,
         DP_OP_102J5_124_3590_n1948, DP_OP_102J5_124_3590_n1947,
         DP_OP_102J5_124_3590_n1946, DP_OP_102J5_124_3590_n1945,
         DP_OP_102J5_124_3590_n1940, DP_OP_102J5_124_3590_n1939,
         DP_OP_102J5_124_3590_n1938, DP_OP_102J5_124_3590_n1937,
         DP_OP_102J5_124_3590_n1936, DP_OP_102J5_124_3590_n1935,
         DP_OP_102J5_124_3590_n1934, DP_OP_102J5_124_3590_n1933,
         DP_OP_102J5_124_3590_n1932, DP_OP_102J5_124_3590_n1931,
         DP_OP_102J5_124_3590_n1930, DP_OP_102J5_124_3590_n1929,
         DP_OP_102J5_124_3590_n1928, DP_OP_102J5_124_3590_n1927,
         DP_OP_102J5_124_3590_n1926, DP_OP_102J5_124_3590_n1925,
         DP_OP_102J5_124_3590_n1924, DP_OP_102J5_124_3590_n1923,
         DP_OP_102J5_124_3590_n1922, DP_OP_102J5_124_3590_n1921,
         DP_OP_102J5_124_3590_n1920, DP_OP_102J5_124_3590_n1919,
         DP_OP_102J5_124_3590_n1918, DP_OP_102J5_124_3590_n1917,
         DP_OP_102J5_124_3590_n1916, DP_OP_102J5_124_3590_n1915,
         DP_OP_102J5_124_3590_n1914, DP_OP_102J5_124_3590_n1913,
         DP_OP_102J5_124_3590_n1912, DP_OP_102J5_124_3590_n1911,
         DP_OP_102J5_124_3590_n1910, DP_OP_102J5_124_3590_n1909,
         DP_OP_102J5_124_3590_n1908, DP_OP_102J5_124_3590_n1907,
         DP_OP_102J5_124_3590_n1906, DP_OP_102J5_124_3590_n1905,
         DP_OP_102J5_124_3590_n1904, DP_OP_102J5_124_3590_n1903,
         DP_OP_102J5_124_3590_n1902, DP_OP_102J5_124_3590_n1901,
         DP_OP_102J5_124_3590_n1896, DP_OP_102J5_124_3590_n1895,
         DP_OP_102J5_124_3590_n1894, DP_OP_102J5_124_3590_n1893,
         DP_OP_102J5_124_3590_n1892, DP_OP_102J5_124_3590_n1891,
         DP_OP_102J5_124_3590_n1890, DP_OP_102J5_124_3590_n1889,
         DP_OP_102J5_124_3590_n1888, DP_OP_102J5_124_3590_n1887,
         DP_OP_102J5_124_3590_n1886, DP_OP_102J5_124_3590_n1885,
         DP_OP_102J5_124_3590_n1884, DP_OP_102J5_124_3590_n1883,
         DP_OP_102J5_124_3590_n1882, DP_OP_102J5_124_3590_n1881,
         DP_OP_102J5_124_3590_n1880, DP_OP_102J5_124_3590_n1879,
         DP_OP_102J5_124_3590_n1878, DP_OP_102J5_124_3590_n1877,
         DP_OP_102J5_124_3590_n1876, DP_OP_102J5_124_3590_n1875,
         DP_OP_102J5_124_3590_n1874, DP_OP_102J5_124_3590_n1873,
         DP_OP_102J5_124_3590_n1872, DP_OP_102J5_124_3590_n1871,
         DP_OP_102J5_124_3590_n1870, DP_OP_102J5_124_3590_n1869,
         DP_OP_102J5_124_3590_n1868, DP_OP_102J5_124_3590_n1867,
         DP_OP_102J5_124_3590_n1866, DP_OP_102J5_124_3590_n1865,
         DP_OP_102J5_124_3590_n1864, DP_OP_102J5_124_3590_n1863,
         DP_OP_102J5_124_3590_n1862, DP_OP_102J5_124_3590_n1861,
         DP_OP_102J5_124_3590_n1860, DP_OP_102J5_124_3590_n1859,
         DP_OP_102J5_124_3590_n1858, DP_OP_102J5_124_3590_n1857,
         DP_OP_102J5_124_3590_n1852, DP_OP_102J5_124_3590_n1851,
         DP_OP_102J5_124_3590_n1850, DP_OP_102J5_124_3590_n1849,
         DP_OP_102J5_124_3590_n1848, DP_OP_102J5_124_3590_n1847,
         DP_OP_102J5_124_3590_n1846, DP_OP_102J5_124_3590_n1845,
         DP_OP_102J5_124_3590_n1844, DP_OP_102J5_124_3590_n1843,
         DP_OP_102J5_124_3590_n1842, DP_OP_102J5_124_3590_n1841,
         DP_OP_102J5_124_3590_n1840, DP_OP_102J5_124_3590_n1839,
         DP_OP_102J5_124_3590_n1838, DP_OP_102J5_124_3590_n1837,
         DP_OP_102J5_124_3590_n1836, DP_OP_102J5_124_3590_n1835,
         DP_OP_102J5_124_3590_n1834, DP_OP_102J5_124_3590_n1833,
         DP_OP_102J5_124_3590_n1832, DP_OP_102J5_124_3590_n1831,
         DP_OP_102J5_124_3590_n1830, DP_OP_102J5_124_3590_n1829,
         DP_OP_102J5_124_3590_n1828, DP_OP_102J5_124_3590_n1827,
         DP_OP_102J5_124_3590_n1826, DP_OP_102J5_124_3590_n1825,
         DP_OP_102J5_124_3590_n1824, DP_OP_102J5_124_3590_n1823,
         DP_OP_102J5_124_3590_n1822, DP_OP_102J5_124_3590_n1821,
         DP_OP_102J5_124_3590_n1820, DP_OP_102J5_124_3590_n1819,
         DP_OP_102J5_124_3590_n1818, DP_OP_102J5_124_3590_n1817,
         DP_OP_102J5_124_3590_n1816, DP_OP_102J5_124_3590_n1815,
         DP_OP_102J5_124_3590_n1814, DP_OP_102J5_124_3590_n1809,
         DP_OP_102J5_124_3590_n1808, DP_OP_102J5_124_3590_n1807,
         DP_OP_102J5_124_3590_n1806, DP_OP_102J5_124_3590_n1805,
         DP_OP_102J5_124_3590_n1804, DP_OP_102J5_124_3590_n1803,
         DP_OP_102J5_124_3590_n1802, DP_OP_102J5_124_3590_n1801,
         DP_OP_102J5_124_3590_n1800, DP_OP_102J5_124_3590_n1799,
         DP_OP_102J5_124_3590_n1798, DP_OP_102J5_124_3590_n1797,
         DP_OP_102J5_124_3590_n1796, DP_OP_102J5_124_3590_n1795,
         DP_OP_102J5_124_3590_n1794, DP_OP_102J5_124_3590_n1793,
         DP_OP_102J5_124_3590_n1792, DP_OP_102J5_124_3590_n1791,
         DP_OP_102J5_124_3590_n1790, DP_OP_102J5_124_3590_n1789,
         DP_OP_102J5_124_3590_n1788, DP_OP_102J5_124_3590_n1787,
         DP_OP_102J5_124_3590_n1786, DP_OP_102J5_124_3590_n1785,
         DP_OP_102J5_124_3590_n1784, DP_OP_102J5_124_3590_n1783,
         DP_OP_102J5_124_3590_n1782, DP_OP_102J5_124_3590_n1781,
         DP_OP_102J5_124_3590_n1780, DP_OP_102J5_124_3590_n1779,
         DP_OP_102J5_124_3590_n1778, DP_OP_102J5_124_3590_n1777,
         DP_OP_102J5_124_3590_n1776, DP_OP_102J5_124_3590_n1775,
         DP_OP_102J5_124_3590_n1774, DP_OP_102J5_124_3590_n1773,
         DP_OP_102J5_124_3590_n1772, DP_OP_102J5_124_3590_n1771,
         DP_OP_102J5_124_3590_n1770, DP_OP_102J5_124_3590_n1765,
         DP_OP_102J5_124_3590_n1764, DP_OP_102J5_124_3590_n1763,
         DP_OP_102J5_124_3590_n1762, DP_OP_102J5_124_3590_n1761,
         DP_OP_102J5_124_3590_n1760, DP_OP_102J5_124_3590_n1759,
         DP_OP_102J5_124_3590_n1758, DP_OP_102J5_124_3590_n1757,
         DP_OP_102J5_124_3590_n1756, DP_OP_102J5_124_3590_n1755,
         DP_OP_102J5_124_3590_n1754, DP_OP_102J5_124_3590_n1753,
         DP_OP_102J5_124_3590_n1752, DP_OP_102J5_124_3590_n1751,
         DP_OP_102J5_124_3590_n1750, DP_OP_102J5_124_3590_n1749,
         DP_OP_102J5_124_3590_n1748, DP_OP_102J5_124_3590_n1747,
         DP_OP_102J5_124_3590_n1746, DP_OP_102J5_124_3590_n1745,
         DP_OP_102J5_124_3590_n1744, DP_OP_102J5_124_3590_n1743,
         DP_OP_102J5_124_3590_n1742, DP_OP_102J5_124_3590_n1741,
         DP_OP_102J5_124_3590_n1740, DP_OP_102J5_124_3590_n1739,
         DP_OP_102J5_124_3590_n1738, DP_OP_102J5_124_3590_n1737,
         DP_OP_102J5_124_3590_n1736, DP_OP_102J5_124_3590_n1735,
         DP_OP_102J5_124_3590_n1734, DP_OP_102J5_124_3590_n1733,
         DP_OP_102J5_124_3590_n1732, DP_OP_102J5_124_3590_n1731,
         DP_OP_102J5_124_3590_n1730, DP_OP_102J5_124_3590_n1729,
         DP_OP_102J5_124_3590_n1728, DP_OP_102J5_124_3590_n1727,
         DP_OP_102J5_124_3590_n1726, DP_OP_102J5_124_3590_n1721,
         DP_OP_102J5_124_3590_n1720, DP_OP_102J5_124_3590_n1719,
         DP_OP_102J5_124_3590_n1718, DP_OP_102J5_124_3590_n1717,
         DP_OP_102J5_124_3590_n1716, DP_OP_102J5_124_3590_n1715,
         DP_OP_102J5_124_3590_n1714, DP_OP_102J5_124_3590_n1713,
         DP_OP_102J5_124_3590_n1712, DP_OP_102J5_124_3590_n1711,
         DP_OP_102J5_124_3590_n1710, DP_OP_102J5_124_3590_n1709,
         DP_OP_102J5_124_3590_n1708, DP_OP_102J5_124_3590_n1707,
         DP_OP_102J5_124_3590_n1706, DP_OP_102J5_124_3590_n1705,
         DP_OP_102J5_124_3590_n1704, DP_OP_102J5_124_3590_n1703,
         DP_OP_102J5_124_3590_n1702, DP_OP_102J5_124_3590_n1701,
         DP_OP_102J5_124_3590_n1700, DP_OP_102J5_124_3590_n1699,
         DP_OP_102J5_124_3590_n1698, DP_OP_102J5_124_3590_n1697,
         DP_OP_102J5_124_3590_n1696, DP_OP_102J5_124_3590_n1695,
         DP_OP_102J5_124_3590_n1694, DP_OP_102J5_124_3590_n1693,
         DP_OP_102J5_124_3590_n1692, DP_OP_102J5_124_3590_n1691,
         DP_OP_102J5_124_3590_n1690, DP_OP_102J5_124_3590_n1689,
         DP_OP_102J5_124_3590_n1688, DP_OP_102J5_124_3590_n1687,
         DP_OP_102J5_124_3590_n1686, DP_OP_102J5_124_3590_n1685,
         DP_OP_102J5_124_3590_n1684, DP_OP_102J5_124_3590_n1683,
         DP_OP_102J5_124_3590_n1682, DP_OP_102J5_124_3590_n1677,
         DP_OP_102J5_124_3590_n1676, DP_OP_102J5_124_3590_n1675,
         DP_OP_102J5_124_3590_n1674, DP_OP_102J5_124_3590_n1673,
         DP_OP_102J5_124_3590_n1672, DP_OP_102J5_124_3590_n1671,
         DP_OP_102J5_124_3590_n1670, DP_OP_102J5_124_3590_n1669,
         DP_OP_102J5_124_3590_n1668, DP_OP_102J5_124_3590_n1667,
         DP_OP_102J5_124_3590_n1666, DP_OP_102J5_124_3590_n1665,
         DP_OP_102J5_124_3590_n1664, DP_OP_102J5_124_3590_n1663,
         DP_OP_102J5_124_3590_n1662, DP_OP_102J5_124_3590_n1661,
         DP_OP_102J5_124_3590_n1660, DP_OP_102J5_124_3590_n1659,
         DP_OP_102J5_124_3590_n1658, DP_OP_102J5_124_3590_n1657,
         DP_OP_102J5_124_3590_n1656, DP_OP_102J5_124_3590_n1655,
         DP_OP_102J5_124_3590_n1654, DP_OP_102J5_124_3590_n1653,
         DP_OP_102J5_124_3590_n1652, DP_OP_102J5_124_3590_n1651,
         DP_OP_102J5_124_3590_n1650, DP_OP_102J5_124_3590_n1649,
         DP_OP_102J5_124_3590_n1648, DP_OP_102J5_124_3590_n1647,
         DP_OP_102J5_124_3590_n1646, DP_OP_102J5_124_3590_n1645,
         DP_OP_102J5_124_3590_n1644, DP_OP_102J5_124_3590_n1643,
         DP_OP_102J5_124_3590_n1642, DP_OP_102J5_124_3590_n1641,
         DP_OP_102J5_124_3590_n1640, DP_OP_102J5_124_3590_n1639,
         DP_OP_102J5_124_3590_n1638, DP_OP_102J5_124_3590_n1633,
         DP_OP_102J5_124_3590_n1632, DP_OP_102J5_124_3590_n1631,
         DP_OP_102J5_124_3590_n1630, DP_OP_102J5_124_3590_n1629,
         DP_OP_102J5_124_3590_n1628, DP_OP_102J5_124_3590_n1627,
         DP_OP_102J5_124_3590_n1626, DP_OP_102J5_124_3590_n1625,
         DP_OP_102J5_124_3590_n1624, DP_OP_102J5_124_3590_n1623,
         DP_OP_102J5_124_3590_n1622, DP_OP_102J5_124_3590_n1621,
         DP_OP_102J5_124_3590_n1620, DP_OP_102J5_124_3590_n1619,
         DP_OP_102J5_124_3590_n1618, DP_OP_102J5_124_3590_n1617,
         DP_OP_102J5_124_3590_n1616, DP_OP_102J5_124_3590_n1615,
         DP_OP_102J5_124_3590_n1614, DP_OP_102J5_124_3590_n1613,
         DP_OP_102J5_124_3590_n1612, DP_OP_102J5_124_3590_n1611,
         DP_OP_102J5_124_3590_n1610, DP_OP_102J5_124_3590_n1609,
         DP_OP_102J5_124_3590_n1608, DP_OP_102J5_124_3590_n1607,
         DP_OP_102J5_124_3590_n1606, DP_OP_102J5_124_3590_n1605,
         DP_OP_102J5_124_3590_n1604, DP_OP_102J5_124_3590_n1603,
         DP_OP_102J5_124_3590_n1602, DP_OP_102J5_124_3590_n1601,
         DP_OP_102J5_124_3590_n1600, DP_OP_102J5_124_3590_n1599,
         DP_OP_102J5_124_3590_n1598, DP_OP_102J5_124_3590_n1597,
         DP_OP_102J5_124_3590_n1596, DP_OP_102J5_124_3590_n1595,
         DP_OP_102J5_124_3590_n1594, DP_OP_102J5_124_3590_n1589,
         DP_OP_102J5_124_3590_n1588, DP_OP_102J5_124_3590_n1587,
         DP_OP_102J5_124_3590_n1586, DP_OP_102J5_124_3590_n1585,
         DP_OP_102J5_124_3590_n1584, DP_OP_102J5_124_3590_n1583,
         DP_OP_102J5_124_3590_n1582, DP_OP_102J5_124_3590_n1581,
         DP_OP_102J5_124_3590_n1580, DP_OP_102J5_124_3590_n1579,
         DP_OP_102J5_124_3590_n1578, DP_OP_102J5_124_3590_n1577,
         DP_OP_102J5_124_3590_n1576, DP_OP_102J5_124_3590_n1575,
         DP_OP_102J5_124_3590_n1574, DP_OP_102J5_124_3590_n1573,
         DP_OP_102J5_124_3590_n1572, DP_OP_102J5_124_3590_n1571,
         DP_OP_102J5_124_3590_n1570, DP_OP_102J5_124_3590_n1569,
         DP_OP_102J5_124_3590_n1568, DP_OP_102J5_124_3590_n1567,
         DP_OP_102J5_124_3590_n1566, DP_OP_102J5_124_3590_n1565,
         DP_OP_102J5_124_3590_n1564, DP_OP_102J5_124_3590_n1563,
         DP_OP_102J5_124_3590_n1562, DP_OP_102J5_124_3590_n1561,
         DP_OP_102J5_124_3590_n1560, DP_OP_102J5_124_3590_n1559,
         DP_OP_102J5_124_3590_n1558, DP_OP_102J5_124_3590_n1557,
         DP_OP_102J5_124_3590_n1556, DP_OP_102J5_124_3590_n1555,
         DP_OP_102J5_124_3590_n1554, DP_OP_102J5_124_3590_n1553,
         DP_OP_102J5_124_3590_n1552, DP_OP_102J5_124_3590_n1551,
         DP_OP_102J5_124_3590_n1550, DP_OP_102J5_124_3590_n1545,
         DP_OP_102J5_124_3590_n1544, DP_OP_102J5_124_3590_n1543,
         DP_OP_102J5_124_3590_n1542, DP_OP_102J5_124_3590_n1541,
         DP_OP_102J5_124_3590_n1540, DP_OP_102J5_124_3590_n1539,
         DP_OP_102J5_124_3590_n1538, DP_OP_102J5_124_3590_n1537,
         DP_OP_102J5_124_3590_n1536, DP_OP_102J5_124_3590_n1535,
         DP_OP_102J5_124_3590_n1534, DP_OP_102J5_124_3590_n1533,
         DP_OP_102J5_124_3590_n1532, DP_OP_102J5_124_3590_n1531,
         DP_OP_102J5_124_3590_n1530, DP_OP_102J5_124_3590_n1529,
         DP_OP_102J5_124_3590_n1528, DP_OP_102J5_124_3590_n1527,
         DP_OP_102J5_124_3590_n1526, DP_OP_102J5_124_3590_n1525,
         DP_OP_102J5_124_3590_n1524, DP_OP_102J5_124_3590_n1523,
         DP_OP_102J5_124_3590_n1522, DP_OP_102J5_124_3590_n1521,
         DP_OP_102J5_124_3590_n1520, DP_OP_102J5_124_3590_n1519,
         DP_OP_102J5_124_3590_n1518, DP_OP_102J5_124_3590_n1517,
         DP_OP_102J5_124_3590_n1516, DP_OP_102J5_124_3590_n1515,
         DP_OP_102J5_124_3590_n1514, DP_OP_102J5_124_3590_n1513,
         DP_OP_102J5_124_3590_n1512, DP_OP_102J5_124_3590_n1511,
         DP_OP_102J5_124_3590_n1510, DP_OP_102J5_124_3590_n1509,
         DP_OP_102J5_124_3590_n1508, DP_OP_102J5_124_3590_n1507,
         DP_OP_102J5_124_3590_n1506, DP_OP_102J5_124_3590_n1481,
         DP_OP_102J5_124_3590_n1480, DP_OP_102J5_124_3590_n1479,
         DP_OP_102J5_124_3590_n1478, DP_OP_102J5_124_3590_n1477,
         DP_OP_102J5_124_3590_n1476, DP_OP_102J5_124_3590_n1475,
         DP_OP_102J5_124_3590_n1474, DP_OP_102J5_124_3590_n1473,
         DP_OP_102J5_124_3590_n1472, DP_OP_102J5_124_3590_n1471,
         DP_OP_102J5_124_3590_n1470, DP_OP_102J5_124_3590_n1469,
         DP_OP_102J5_124_3590_n1468, DP_OP_102J5_124_3590_n1466,
         DP_OP_102J5_124_3590_n1465, DP_OP_102J5_124_3590_n1464,
         DP_OP_102J5_124_3590_n1463, DP_OP_102J5_124_3590_n1462,
         DP_OP_102J5_124_3590_n1461, DP_OP_102J5_124_3590_n1460,
         DP_OP_102J5_124_3590_n1459, DP_OP_102J5_124_3590_n1458,
         DP_OP_102J5_124_3590_n1457, DP_OP_102J5_124_3590_n1456,
         DP_OP_102J5_124_3590_n1455, DP_OP_102J5_124_3590_n1454,
         DP_OP_102J5_124_3590_n1453, DP_OP_102J5_124_3590_n1452,
         DP_OP_102J5_124_3590_n1451, DP_OP_102J5_124_3590_n1450,
         DP_OP_102J5_124_3590_n1449, DP_OP_102J5_124_3590_n1448,
         DP_OP_102J5_124_3590_n1447, DP_OP_102J5_124_3590_n1446,
         DP_OP_102J5_124_3590_n1445, DP_OP_102J5_124_3590_n1444,
         DP_OP_102J5_124_3590_n1443, DP_OP_102J5_124_3590_n1442,
         DP_OP_102J5_124_3590_n1441, DP_OP_102J5_124_3590_n1440,
         DP_OP_102J5_124_3590_n1439, DP_OP_102J5_124_3590_n1438,
         DP_OP_102J5_124_3590_n1437, DP_OP_102J5_124_3590_n1436,
         DP_OP_102J5_124_3590_n1435, DP_OP_102J5_124_3590_n1434,
         DP_OP_102J5_124_3590_n1433, DP_OP_102J5_124_3590_n1432,
         DP_OP_102J5_124_3590_n1431, DP_OP_102J5_124_3590_n1430,
         DP_OP_102J5_124_3590_n1429, DP_OP_102J5_124_3590_n1428,
         DP_OP_102J5_124_3590_n1427, DP_OP_102J5_124_3590_n1426,
         DP_OP_102J5_124_3590_n1425, DP_OP_102J5_124_3590_n1424,
         DP_OP_102J5_124_3590_n1423, DP_OP_102J5_124_3590_n1422,
         DP_OP_102J5_124_3590_n1421, DP_OP_102J5_124_3590_n1420,
         DP_OP_102J5_124_3590_n1419, DP_OP_102J5_124_3590_n1418,
         DP_OP_102J5_124_3590_n1417, DP_OP_102J5_124_3590_n1416,
         DP_OP_102J5_124_3590_n1415, DP_OP_102J5_124_3590_n1414,
         DP_OP_102J5_124_3590_n1413, DP_OP_102J5_124_3590_n1412,
         DP_OP_102J5_124_3590_n1411, DP_OP_102J5_124_3590_n1410,
         DP_OP_102J5_124_3590_n1409, DP_OP_102J5_124_3590_n1408,
         DP_OP_102J5_124_3590_n1407, DP_OP_102J5_124_3590_n1406,
         DP_OP_102J5_124_3590_n1405, DP_OP_102J5_124_3590_n1404,
         DP_OP_102J5_124_3590_n1403, DP_OP_102J5_124_3590_n1402,
         DP_OP_102J5_124_3590_n1401, DP_OP_102J5_124_3590_n1400,
         DP_OP_102J5_124_3590_n1399, DP_OP_102J5_124_3590_n1398,
         DP_OP_102J5_124_3590_n1397, DP_OP_102J5_124_3590_n1396,
         DP_OP_102J5_124_3590_n1395, DP_OP_102J5_124_3590_n1394,
         DP_OP_102J5_124_3590_n1393, DP_OP_102J5_124_3590_n1392,
         DP_OP_102J5_124_3590_n1391, DP_OP_102J5_124_3590_n1390,
         DP_OP_102J5_124_3590_n1389, DP_OP_102J5_124_3590_n1388,
         DP_OP_102J5_124_3590_n1387, DP_OP_102J5_124_3590_n1386,
         DP_OP_102J5_124_3590_n1385, DP_OP_102J5_124_3590_n1384,
         DP_OP_102J5_124_3590_n1383, DP_OP_102J5_124_3590_n1382,
         DP_OP_102J5_124_3590_n1381, DP_OP_102J5_124_3590_n1380,
         DP_OP_102J5_124_3590_n1379, DP_OP_102J5_124_3590_n1378,
         DP_OP_102J5_124_3590_n1377, DP_OP_102J5_124_3590_n1376,
         DP_OP_102J5_124_3590_n1375, DP_OP_102J5_124_3590_n1374,
         DP_OP_102J5_124_3590_n1373, DP_OP_102J5_124_3590_n1372,
         DP_OP_102J5_124_3590_n1371, DP_OP_102J5_124_3590_n1370,
         DP_OP_102J5_124_3590_n1369, DP_OP_102J5_124_3590_n1368,
         DP_OP_102J5_124_3590_n1367, DP_OP_102J5_124_3590_n1366,
         DP_OP_102J5_124_3590_n1365, DP_OP_102J5_124_3590_n1364,
         DP_OP_102J5_124_3590_n1363, DP_OP_102J5_124_3590_n1362,
         DP_OP_102J5_124_3590_n1361, DP_OP_102J5_124_3590_n1360,
         DP_OP_102J5_124_3590_n1359, DP_OP_102J5_124_3590_n1358,
         DP_OP_102J5_124_3590_n1357, DP_OP_102J5_124_3590_n1356,
         DP_OP_102J5_124_3590_n1355, DP_OP_102J5_124_3590_n1354,
         DP_OP_102J5_124_3590_n1353, DP_OP_102J5_124_3590_n1352,
         DP_OP_102J5_124_3590_n1351, DP_OP_102J5_124_3590_n1350,
         DP_OP_102J5_124_3590_n1349, DP_OP_102J5_124_3590_n1348,
         DP_OP_102J5_124_3590_n1347, DP_OP_102J5_124_3590_n1346,
         DP_OP_102J5_124_3590_n1345, DP_OP_102J5_124_3590_n1344,
         DP_OP_102J5_124_3590_n1343, DP_OP_102J5_124_3590_n1342,
         DP_OP_102J5_124_3590_n1341, DP_OP_102J5_124_3590_n1340,
         DP_OP_102J5_124_3590_n1339, DP_OP_102J5_124_3590_n1338,
         DP_OP_102J5_124_3590_n1337, DP_OP_102J5_124_3590_n1336,
         DP_OP_102J5_124_3590_n1335, DP_OP_102J5_124_3590_n1334,
         DP_OP_102J5_124_3590_n1333, DP_OP_102J5_124_3590_n1332,
         DP_OP_102J5_124_3590_n1331, DP_OP_102J5_124_3590_n1330,
         DP_OP_102J5_124_3590_n1329, DP_OP_102J5_124_3590_n1328,
         DP_OP_102J5_124_3590_n1327, DP_OP_102J5_124_3590_n1326,
         DP_OP_102J5_124_3590_n1325, DP_OP_102J5_124_3590_n1324,
         DP_OP_102J5_124_3590_n1323, DP_OP_102J5_124_3590_n1322,
         DP_OP_102J5_124_3590_n1321, DP_OP_102J5_124_3590_n1320,
         DP_OP_102J5_124_3590_n1319, DP_OP_102J5_124_3590_n1318,
         DP_OP_102J5_124_3590_n1317, DP_OP_102J5_124_3590_n1316,
         DP_OP_102J5_124_3590_n1315, DP_OP_102J5_124_3590_n1314,
         DP_OP_102J5_124_3590_n1313, DP_OP_102J5_124_3590_n1312,
         DP_OP_102J5_124_3590_n1311, DP_OP_102J5_124_3590_n1310,
         DP_OP_102J5_124_3590_n1309, DP_OP_102J5_124_3590_n1308,
         DP_OP_102J5_124_3590_n1307, DP_OP_102J5_124_3590_n1306,
         DP_OP_102J5_124_3590_n1305, DP_OP_102J5_124_3590_n1304,
         DP_OP_102J5_124_3590_n1303, DP_OP_102J5_124_3590_n1302,
         DP_OP_102J5_124_3590_n1301, DP_OP_102J5_124_3590_n1300,
         DP_OP_102J5_124_3590_n1299, DP_OP_102J5_124_3590_n1298,
         DP_OP_102J5_124_3590_n1297, DP_OP_102J5_124_3590_n1296,
         DP_OP_102J5_124_3590_n1295, DP_OP_102J5_124_3590_n1294,
         DP_OP_102J5_124_3590_n1293, DP_OP_102J5_124_3590_n1292,
         DP_OP_102J5_124_3590_n1291, DP_OP_102J5_124_3590_n1290,
         DP_OP_102J5_124_3590_n1289, DP_OP_102J5_124_3590_n1288,
         DP_OP_102J5_124_3590_n1287, DP_OP_102J5_124_3590_n1286,
         DP_OP_102J5_124_3590_n1285, DP_OP_102J5_124_3590_n1284,
         DP_OP_102J5_124_3590_n1283, DP_OP_102J5_124_3590_n1282,
         DP_OP_102J5_124_3590_n1281, DP_OP_102J5_124_3590_n1280,
         DP_OP_102J5_124_3590_n1279, DP_OP_102J5_124_3590_n1278,
         DP_OP_102J5_124_3590_n1277, DP_OP_102J5_124_3590_n1276,
         DP_OP_102J5_124_3590_n1275, DP_OP_102J5_124_3590_n1274,
         DP_OP_102J5_124_3590_n1273, DP_OP_102J5_124_3590_n1272,
         DP_OP_102J5_124_3590_n1271, DP_OP_102J5_124_3590_n1270,
         DP_OP_102J5_124_3590_n1269, DP_OP_102J5_124_3590_n1268,
         DP_OP_102J5_124_3590_n1267, DP_OP_102J5_124_3590_n1266,
         DP_OP_102J5_124_3590_n1265, DP_OP_102J5_124_3590_n1264,
         DP_OP_102J5_124_3590_n1263, DP_OP_102J5_124_3590_n1262,
         DP_OP_102J5_124_3590_n1261, DP_OP_102J5_124_3590_n1260,
         DP_OP_102J5_124_3590_n1259, DP_OP_102J5_124_3590_n1258,
         DP_OP_102J5_124_3590_n1257, DP_OP_102J5_124_3590_n1256,
         DP_OP_102J5_124_3590_n1255, DP_OP_102J5_124_3590_n1254,
         DP_OP_102J5_124_3590_n1253, DP_OP_102J5_124_3590_n1252,
         DP_OP_102J5_124_3590_n1251, DP_OP_102J5_124_3590_n1250,
         DP_OP_102J5_124_3590_n1249, DP_OP_102J5_124_3590_n1248,
         DP_OP_102J5_124_3590_n1247, DP_OP_102J5_124_3590_n1246,
         DP_OP_102J5_124_3590_n1245, DP_OP_102J5_124_3590_n1244,
         DP_OP_102J5_124_3590_n1243, DP_OP_102J5_124_3590_n1242,
         DP_OP_102J5_124_3590_n1241, DP_OP_102J5_124_3590_n1240,
         DP_OP_102J5_124_3590_n1239, DP_OP_102J5_124_3590_n1238,
         DP_OP_102J5_124_3590_n1237, DP_OP_102J5_124_3590_n1236,
         DP_OP_102J5_124_3590_n1235, DP_OP_102J5_124_3590_n1234,
         DP_OP_102J5_124_3590_n1233, DP_OP_102J5_124_3590_n1232,
         DP_OP_102J5_124_3590_n1231, DP_OP_102J5_124_3590_n1230,
         DP_OP_102J5_124_3590_n1229, DP_OP_102J5_124_3590_n1228,
         DP_OP_102J5_124_3590_n1227, DP_OP_102J5_124_3590_n1226,
         DP_OP_102J5_124_3590_n1225, DP_OP_102J5_124_3590_n1224,
         DP_OP_102J5_124_3590_n1223, DP_OP_102J5_124_3590_n1222,
         DP_OP_102J5_124_3590_n1221, DP_OP_102J5_124_3590_n1220,
         DP_OP_102J5_124_3590_n1219, DP_OP_102J5_124_3590_n1218,
         DP_OP_102J5_124_3590_n1217, DP_OP_102J5_124_3590_n1216,
         DP_OP_102J5_124_3590_n1215, DP_OP_102J5_124_3590_n1214,
         DP_OP_102J5_124_3590_n1213, DP_OP_102J5_124_3590_n1212,
         DP_OP_102J5_124_3590_n1211, DP_OP_102J5_124_3590_n1210,
         DP_OP_102J5_124_3590_n1209, DP_OP_102J5_124_3590_n1208,
         DP_OP_102J5_124_3590_n1207, DP_OP_102J5_124_3590_n1206,
         DP_OP_102J5_124_3590_n1205, DP_OP_102J5_124_3590_n1204,
         DP_OP_102J5_124_3590_n1203, DP_OP_102J5_124_3590_n1202,
         DP_OP_102J5_124_3590_n1201, DP_OP_102J5_124_3590_n1200,
         DP_OP_102J5_124_3590_n1199, DP_OP_102J5_124_3590_n1198,
         DP_OP_102J5_124_3590_n1197, DP_OP_102J5_124_3590_n1196,
         DP_OP_102J5_124_3590_n1195, DP_OP_102J5_124_3590_n1194,
         DP_OP_102J5_124_3590_n1193, DP_OP_102J5_124_3590_n1192,
         DP_OP_102J5_124_3590_n1191, DP_OP_102J5_124_3590_n1190,
         DP_OP_102J5_124_3590_n1189, DP_OP_102J5_124_3590_n1188,
         DP_OP_102J5_124_3590_n1187, DP_OP_102J5_124_3590_n1186,
         DP_OP_102J5_124_3590_n1185, DP_OP_102J5_124_3590_n1184,
         DP_OP_102J5_124_3590_n1183, DP_OP_102J5_124_3590_n1182,
         DP_OP_102J5_124_3590_n1181, DP_OP_102J5_124_3590_n1180,
         DP_OP_102J5_124_3590_n1179, DP_OP_102J5_124_3590_n1178,
         DP_OP_102J5_124_3590_n1177, DP_OP_102J5_124_3590_n1176,
         DP_OP_102J5_124_3590_n1175, DP_OP_102J5_124_3590_n1174,
         DP_OP_102J5_124_3590_n1173, DP_OP_102J5_124_3590_n1172,
         DP_OP_102J5_124_3590_n1171, DP_OP_102J5_124_3590_n1170,
         DP_OP_102J5_124_3590_n1169, DP_OP_102J5_124_3590_n1168,
         DP_OP_102J5_124_3590_n1167, DP_OP_102J5_124_3590_n1166,
         DP_OP_102J5_124_3590_n1165, DP_OP_102J5_124_3590_n1164,
         DP_OP_102J5_124_3590_n1163, DP_OP_102J5_124_3590_n1162,
         DP_OP_102J5_124_3590_n1161, DP_OP_102J5_124_3590_n1160,
         DP_OP_102J5_124_3590_n1159, DP_OP_102J5_124_3590_n1158,
         DP_OP_102J5_124_3590_n1157, DP_OP_102J5_124_3590_n1156,
         DP_OP_102J5_124_3590_n1155, DP_OP_102J5_124_3590_n1154,
         DP_OP_102J5_124_3590_n1153, DP_OP_102J5_124_3590_n1152,
         DP_OP_102J5_124_3590_n1151, DP_OP_102J5_124_3590_n1150,
         DP_OP_102J5_124_3590_n1149, DP_OP_102J5_124_3590_n1148,
         DP_OP_102J5_124_3590_n1147, DP_OP_102J5_124_3590_n1146,
         DP_OP_102J5_124_3590_n1145, DP_OP_102J5_124_3590_n1144,
         DP_OP_102J5_124_3590_n1143, DP_OP_102J5_124_3590_n1142,
         DP_OP_102J5_124_3590_n1141, DP_OP_102J5_124_3590_n1140,
         DP_OP_102J5_124_3590_n1139, DP_OP_102J5_124_3590_n1138,
         DP_OP_102J5_124_3590_n1137, DP_OP_102J5_124_3590_n1136,
         DP_OP_102J5_124_3590_n1135, DP_OP_102J5_124_3590_n1134,
         DP_OP_102J5_124_3590_n1133, DP_OP_102J5_124_3590_n1132,
         DP_OP_102J5_124_3590_n1131, DP_OP_102J5_124_3590_n1130,
         DP_OP_102J5_124_3590_n1129, DP_OP_102J5_124_3590_n1128,
         DP_OP_102J5_124_3590_n1127, DP_OP_102J5_124_3590_n1126,
         DP_OP_102J5_124_3590_n1125, DP_OP_102J5_124_3590_n1124,
         DP_OP_102J5_124_3590_n1123, DP_OP_102J5_124_3590_n1122,
         DP_OP_102J5_124_3590_n1121, DP_OP_102J5_124_3590_n1120,
         DP_OP_102J5_124_3590_n1119, DP_OP_102J5_124_3590_n1118,
         DP_OP_102J5_124_3590_n1117, DP_OP_102J5_124_3590_n1116,
         DP_OP_102J5_124_3590_n1115, DP_OP_102J5_124_3590_n1114,
         DP_OP_102J5_124_3590_n1113, DP_OP_102J5_124_3590_n1112,
         DP_OP_102J5_124_3590_n1111, DP_OP_102J5_124_3590_n1110,
         DP_OP_102J5_124_3590_n1109, DP_OP_102J5_124_3590_n1108,
         DP_OP_102J5_124_3590_n1107, DP_OP_102J5_124_3590_n1106,
         DP_OP_102J5_124_3590_n1105, DP_OP_102J5_124_3590_n1104,
         DP_OP_102J5_124_3590_n1103, DP_OP_102J5_124_3590_n1102,
         DP_OP_102J5_124_3590_n1101, DP_OP_102J5_124_3590_n1100,
         DP_OP_102J5_124_3590_n1099, DP_OP_102J5_124_3590_n1098,
         DP_OP_102J5_124_3590_n1097, DP_OP_102J5_124_3590_n1096,
         DP_OP_102J5_124_3590_n1095, DP_OP_102J5_124_3590_n1094,
         DP_OP_102J5_124_3590_n1093, DP_OP_102J5_124_3590_n1092,
         DP_OP_102J5_124_3590_n1091, DP_OP_102J5_124_3590_n1090,
         DP_OP_102J5_124_3590_n1089, DP_OP_102J5_124_3590_n1088,
         DP_OP_102J5_124_3590_n1087, DP_OP_102J5_124_3590_n1086,
         DP_OP_102J5_124_3590_n1085, DP_OP_102J5_124_3590_n1084,
         DP_OP_102J5_124_3590_n1083, DP_OP_102J5_124_3590_n1082,
         DP_OP_102J5_124_3590_n1081, DP_OP_102J5_124_3590_n1080,
         DP_OP_102J5_124_3590_n1079, DP_OP_102J5_124_3590_n1078,
         DP_OP_102J5_124_3590_n1077, DP_OP_102J5_124_3590_n1076,
         DP_OP_102J5_124_3590_n1075, DP_OP_102J5_124_3590_n1074,
         DP_OP_102J5_124_3590_n1073, DP_OP_102J5_124_3590_n1072,
         DP_OP_102J5_124_3590_n1071, DP_OP_102J5_124_3590_n1070,
         DP_OP_102J5_124_3590_n1069, DP_OP_102J5_124_3590_n1068,
         DP_OP_102J5_124_3590_n1067, DP_OP_102J5_124_3590_n1066,
         DP_OP_102J5_124_3590_n1065, DP_OP_102J5_124_3590_n1064,
         DP_OP_102J5_124_3590_n1063, DP_OP_102J5_124_3590_n1062,
         DP_OP_102J5_124_3590_n1061, DP_OP_102J5_124_3590_n1060,
         DP_OP_102J5_124_3590_n1059, DP_OP_102J5_124_3590_n1058,
         DP_OP_102J5_124_3590_n1057, DP_OP_102J5_124_3590_n1056,
         DP_OP_102J5_124_3590_n1055, DP_OP_102J5_124_3590_n1054,
         DP_OP_102J5_124_3590_n1053, DP_OP_102J5_124_3590_n1052,
         DP_OP_102J5_124_3590_n1051, DP_OP_102J5_124_3590_n1050,
         DP_OP_102J5_124_3590_n1049, DP_OP_102J5_124_3590_n1048,
         DP_OP_102J5_124_3590_n1047, DP_OP_102J5_124_3590_n1046,
         DP_OP_102J5_124_3590_n1045, DP_OP_102J5_124_3590_n1044,
         DP_OP_102J5_124_3590_n1043, DP_OP_102J5_124_3590_n1042,
         DP_OP_102J5_124_3590_n1041, DP_OP_102J5_124_3590_n1040,
         DP_OP_102J5_124_3590_n1039, DP_OP_102J5_124_3590_n1038,
         DP_OP_102J5_124_3590_n1037, DP_OP_102J5_124_3590_n1036,
         DP_OP_102J5_124_3590_n1035, DP_OP_102J5_124_3590_n1034,
         DP_OP_102J5_124_3590_n1033, DP_OP_102J5_124_3590_n1032,
         DP_OP_102J5_124_3590_n1031, DP_OP_102J5_124_3590_n1030,
         DP_OP_102J5_124_3590_n1029, DP_OP_102J5_124_3590_n1028,
         DP_OP_102J5_124_3590_n1027, DP_OP_102J5_124_3590_n1026,
         DP_OP_102J5_124_3590_n1025, DP_OP_102J5_124_3590_n1024,
         DP_OP_102J5_124_3590_n1023, DP_OP_102J5_124_3590_n1022,
         DP_OP_102J5_124_3590_n1021, DP_OP_102J5_124_3590_n1020,
         DP_OP_102J5_124_3590_n1019, DP_OP_102J5_124_3590_n1018,
         DP_OP_102J5_124_3590_n1017, DP_OP_102J5_124_3590_n1016,
         DP_OP_102J5_124_3590_n1015, DP_OP_102J5_124_3590_n1014,
         DP_OP_102J5_124_3590_n1013, DP_OP_102J5_124_3590_n1012,
         DP_OP_102J5_124_3590_n1011, DP_OP_102J5_124_3590_n1010,
         DP_OP_102J5_124_3590_n1009, DP_OP_102J5_124_3590_n1008,
         DP_OP_102J5_124_3590_n1007, DP_OP_102J5_124_3590_n1006,
         DP_OP_102J5_124_3590_n1005, DP_OP_102J5_124_3590_n1004,
         DP_OP_102J5_124_3590_n1003, DP_OP_102J5_124_3590_n1002,
         DP_OP_102J5_124_3590_n1001, DP_OP_102J5_124_3590_n1000,
         DP_OP_102J5_124_3590_n999, DP_OP_102J5_124_3590_n998,
         DP_OP_102J5_124_3590_n997, DP_OP_102J5_124_3590_n996,
         DP_OP_102J5_124_3590_n995, DP_OP_102J5_124_3590_n994,
         DP_OP_102J5_124_3590_n993, DP_OP_102J5_124_3590_n992,
         DP_OP_102J5_124_3590_n991, DP_OP_102J5_124_3590_n990,
         DP_OP_102J5_124_3590_n989, DP_OP_102J5_124_3590_n988,
         DP_OP_102J5_124_3590_n987, DP_OP_102J5_124_3590_n986,
         DP_OP_102J5_124_3590_n985, DP_OP_102J5_124_3590_n984,
         DP_OP_102J5_124_3590_n983, DP_OP_102J5_124_3590_n982,
         DP_OP_102J5_124_3590_n981, DP_OP_102J5_124_3590_n980,
         DP_OP_102J5_124_3590_n979, DP_OP_102J5_124_3590_n978,
         DP_OP_102J5_124_3590_n977, DP_OP_102J5_124_3590_n976,
         DP_OP_102J5_124_3590_n975, DP_OP_102J5_124_3590_n974,
         DP_OP_102J5_124_3590_n973, DP_OP_102J5_124_3590_n972,
         DP_OP_102J5_124_3590_n971, DP_OP_102J5_124_3590_n970,
         DP_OP_102J5_124_3590_n969, DP_OP_102J5_124_3590_n968,
         DP_OP_102J5_124_3590_n967, DP_OP_102J5_124_3590_n966,
         DP_OP_102J5_124_3590_n965, DP_OP_102J5_124_3590_n964,
         DP_OP_102J5_124_3590_n963, DP_OP_102J5_124_3590_n962,
         DP_OP_102J5_124_3590_n961, DP_OP_102J5_124_3590_n960,
         DP_OP_102J5_124_3590_n959, DP_OP_102J5_124_3590_n958,
         DP_OP_102J5_124_3590_n957, DP_OP_102J5_124_3590_n956,
         DP_OP_102J5_124_3590_n955, DP_OP_102J5_124_3590_n954,
         DP_OP_102J5_124_3590_n953, DP_OP_102J5_124_3590_n952,
         DP_OP_102J5_124_3590_n951, DP_OP_102J5_124_3590_n950,
         DP_OP_102J5_124_3590_n949, DP_OP_102J5_124_3590_n948,
         DP_OP_102J5_124_3590_n947, DP_OP_102J5_124_3590_n946,
         DP_OP_102J5_124_3590_n945, DP_OP_102J5_124_3590_n944,
         DP_OP_102J5_124_3590_n943, DP_OP_102J5_124_3590_n942,
         DP_OP_102J5_124_3590_n941, DP_OP_102J5_124_3590_n940,
         DP_OP_102J5_124_3590_n939, DP_OP_102J5_124_3590_n938,
         DP_OP_102J5_124_3590_n937, DP_OP_102J5_124_3590_n936,
         DP_OP_102J5_124_3590_n935, DP_OP_102J5_124_3590_n934,
         DP_OP_102J5_124_3590_n933, DP_OP_102J5_124_3590_n932,
         DP_OP_102J5_124_3590_n931, DP_OP_102J5_124_3590_n930,
         DP_OP_102J5_124_3590_n929, DP_OP_102J5_124_3590_n928,
         DP_OP_102J5_124_3590_n927, DP_OP_102J5_124_3590_n926,
         DP_OP_102J5_124_3590_n925, DP_OP_102J5_124_3590_n924,
         DP_OP_102J5_124_3590_n923, DP_OP_102J5_124_3590_n922,
         DP_OP_102J5_124_3590_n921, DP_OP_102J5_124_3590_n920,
         DP_OP_102J5_124_3590_n919, DP_OP_102J5_124_3590_n918,
         DP_OP_102J5_124_3590_n917, DP_OP_102J5_124_3590_n916,
         DP_OP_102J5_124_3590_n915, DP_OP_102J5_124_3590_n914,
         DP_OP_102J5_124_3590_n913, DP_OP_102J5_124_3590_n912,
         DP_OP_102J5_124_3590_n911, DP_OP_102J5_124_3590_n910,
         DP_OP_102J5_124_3590_n909, DP_OP_102J5_124_3590_n908,
         DP_OP_102J5_124_3590_n907, DP_OP_102J5_124_3590_n906,
         DP_OP_102J5_124_3590_n905, DP_OP_102J5_124_3590_n904,
         DP_OP_102J5_124_3590_n903, DP_OP_102J5_124_3590_n902,
         DP_OP_102J5_124_3590_n901, DP_OP_102J5_124_3590_n900,
         DP_OP_102J5_124_3590_n899, DP_OP_102J5_124_3590_n898,
         DP_OP_102J5_124_3590_n897, DP_OP_102J5_124_3590_n896,
         DP_OP_102J5_124_3590_n895, DP_OP_102J5_124_3590_n894,
         DP_OP_102J5_124_3590_n893, DP_OP_102J5_124_3590_n892,
         DP_OP_102J5_124_3590_n891, DP_OP_102J5_124_3590_n890,
         DP_OP_102J5_124_3590_n889, DP_OP_102J5_124_3590_n888,
         DP_OP_102J5_124_3590_n887, DP_OP_102J5_124_3590_n886,
         DP_OP_102J5_124_3590_n885, DP_OP_102J5_124_3590_n884,
         DP_OP_102J5_124_3590_n883, DP_OP_102J5_124_3590_n882,
         DP_OP_102J5_124_3590_n881, DP_OP_102J5_124_3590_n880,
         DP_OP_102J5_124_3590_n879, DP_OP_102J5_124_3590_n878,
         DP_OP_102J5_124_3590_n877, DP_OP_102J5_124_3590_n876,
         DP_OP_102J5_124_3590_n875, DP_OP_102J5_124_3590_n874,
         DP_OP_102J5_124_3590_n873, DP_OP_102J5_124_3590_n872,
         DP_OP_102J5_124_3590_n871, DP_OP_102J5_124_3590_n870,
         DP_OP_102J5_124_3590_n869, DP_OP_102J5_124_3590_n868,
         DP_OP_102J5_124_3590_n867, DP_OP_102J5_124_3590_n866,
         DP_OP_102J5_124_3590_n865, DP_OP_102J5_124_3590_n864,
         DP_OP_102J5_124_3590_n863, DP_OP_102J5_124_3590_n862,
         DP_OP_102J5_124_3590_n861, DP_OP_102J5_124_3590_n860,
         DP_OP_102J5_124_3590_n859, DP_OP_102J5_124_3590_n858,
         DP_OP_102J5_124_3590_n857, DP_OP_102J5_124_3590_n856,
         DP_OP_102J5_124_3590_n855, DP_OP_102J5_124_3590_n854,
         DP_OP_102J5_124_3590_n853, DP_OP_102J5_124_3590_n852,
         DP_OP_102J5_124_3590_n851, DP_OP_102J5_124_3590_n850,
         DP_OP_102J5_124_3590_n849, DP_OP_102J5_124_3590_n848,
         DP_OP_102J5_124_3590_n847, DP_OP_102J5_124_3590_n846,
         DP_OP_102J5_124_3590_n845, DP_OP_102J5_124_3590_n844,
         DP_OP_102J5_124_3590_n843, DP_OP_102J5_124_3590_n842,
         DP_OP_102J5_124_3590_n841, DP_OP_102J5_124_3590_n840,
         DP_OP_102J5_124_3590_n839, DP_OP_102J5_124_3590_n838,
         DP_OP_102J5_124_3590_n837, DP_OP_102J5_124_3590_n836,
         DP_OP_102J5_124_3590_n835, DP_OP_102J5_124_3590_n834,
         DP_OP_102J5_124_3590_n833, DP_OP_102J5_124_3590_n832,
         DP_OP_102J5_124_3590_n831, DP_OP_102J5_124_3590_n830,
         DP_OP_102J5_124_3590_n829, DP_OP_102J5_124_3590_n828,
         DP_OP_102J5_124_3590_n827, DP_OP_102J5_124_3590_n826,
         DP_OP_102J5_124_3590_n825, DP_OP_102J5_124_3590_n824,
         DP_OP_102J5_124_3590_n823, DP_OP_102J5_124_3590_n822,
         DP_OP_102J5_124_3590_n821, DP_OP_102J5_124_3590_n820,
         DP_OP_102J5_124_3590_n819, DP_OP_102J5_124_3590_n818,
         DP_OP_102J5_124_3590_n817, DP_OP_102J5_124_3590_n816,
         DP_OP_102J5_124_3590_n815, DP_OP_102J5_124_3590_n814,
         DP_OP_102J5_124_3590_n813, DP_OP_102J5_124_3590_n812,
         DP_OP_102J5_124_3590_n811, DP_OP_102J5_124_3590_n810,
         DP_OP_102J5_124_3590_n809, DP_OP_102J5_124_3590_n808,
         DP_OP_102J5_124_3590_n807, DP_OP_102J5_124_3590_n806,
         DP_OP_102J5_124_3590_n805, DP_OP_102J5_124_3590_n804,
         DP_OP_102J5_124_3590_n803, DP_OP_102J5_124_3590_n802,
         DP_OP_102J5_124_3590_n801, DP_OP_102J5_124_3590_n800,
         DP_OP_102J5_124_3590_n799, DP_OP_102J5_124_3590_n798,
         DP_OP_102J5_124_3590_n797, DP_OP_102J5_124_3590_n796,
         DP_OP_102J5_124_3590_n795, DP_OP_102J5_124_3590_n794,
         DP_OP_102J5_124_3590_n793, DP_OP_102J5_124_3590_n792,
         DP_OP_102J5_124_3590_n791, DP_OP_102J5_124_3590_n790,
         DP_OP_102J5_124_3590_n789, DP_OP_102J5_124_3590_n788,
         DP_OP_102J5_124_3590_n787, DP_OP_102J5_124_3590_n786,
         DP_OP_102J5_124_3590_n785, DP_OP_102J5_124_3590_n784,
         DP_OP_102J5_124_3590_n783, DP_OP_102J5_124_3590_n782,
         DP_OP_102J5_124_3590_n781, DP_OP_102J5_124_3590_n780,
         DP_OP_102J5_124_3590_n779, DP_OP_102J5_124_3590_n778,
         DP_OP_102J5_124_3590_n777, DP_OP_102J5_124_3590_n776,
         DP_OP_102J5_124_3590_n775, DP_OP_102J5_124_3590_n774,
         DP_OP_102J5_124_3590_n773, DP_OP_102J5_124_3590_n772,
         DP_OP_102J5_124_3590_n771, DP_OP_102J5_124_3590_n770,
         DP_OP_102J5_124_3590_n769, DP_OP_102J5_124_3590_n768,
         DP_OP_102J5_124_3590_n767, DP_OP_102J5_124_3590_n766,
         DP_OP_102J5_124_3590_n765, DP_OP_102J5_124_3590_n764,
         DP_OP_102J5_124_3590_n763, DP_OP_102J5_124_3590_n762,
         DP_OP_102J5_124_3590_n761, DP_OP_102J5_124_3590_n760,
         DP_OP_102J5_124_3590_n759, DP_OP_102J5_124_3590_n758,
         DP_OP_102J5_124_3590_n757, DP_OP_102J5_124_3590_n756,
         DP_OP_102J5_124_3590_n755, DP_OP_102J5_124_3590_n754,
         DP_OP_102J5_124_3590_n753, DP_OP_102J5_124_3590_n752,
         DP_OP_102J5_124_3590_n751, DP_OP_102J5_124_3590_n750,
         DP_OP_102J5_124_3590_n749, DP_OP_102J5_124_3590_n748,
         DP_OP_102J5_124_3590_n747, DP_OP_102J5_124_3590_n746,
         DP_OP_102J5_124_3590_n745, DP_OP_102J5_124_3590_n744,
         DP_OP_102J5_124_3590_n743, DP_OP_102J5_124_3590_n742,
         DP_OP_102J5_124_3590_n741, DP_OP_102J5_124_3590_n740,
         DP_OP_102J5_124_3590_n739, DP_OP_102J5_124_3590_n738,
         DP_OP_102J5_124_3590_n737, DP_OP_102J5_124_3590_n736,
         DP_OP_102J5_124_3590_n735, DP_OP_102J5_124_3590_n734,
         DP_OP_102J5_124_3590_n733, DP_OP_102J5_124_3590_n732,
         DP_OP_102J5_124_3590_n731, DP_OP_102J5_124_3590_n730,
         DP_OP_102J5_124_3590_n729, DP_OP_102J5_124_3590_n728,
         DP_OP_102J5_124_3590_n727, DP_OP_102J5_124_3590_n726,
         DP_OP_102J5_124_3590_n725, DP_OP_102J5_124_3590_n724,
         DP_OP_102J5_124_3590_n723, DP_OP_102J5_124_3590_n722,
         DP_OP_102J5_124_3590_n721, DP_OP_102J5_124_3590_n720,
         DP_OP_102J5_124_3590_n719, DP_OP_102J5_124_3590_n718,
         DP_OP_102J5_124_3590_n717, DP_OP_102J5_124_3590_n716,
         DP_OP_102J5_124_3590_n715, DP_OP_102J5_124_3590_n714,
         DP_OP_102J5_124_3590_n713, DP_OP_102J5_124_3590_n712,
         DP_OP_102J5_124_3590_n711, DP_OP_102J5_124_3590_n710,
         DP_OP_102J5_124_3590_n709, DP_OP_102J5_124_3590_n708,
         DP_OP_102J5_124_3590_n707, DP_OP_102J5_124_3590_n706,
         DP_OP_102J5_124_3590_n705, DP_OP_102J5_124_3590_n704,
         DP_OP_102J5_124_3590_n703, DP_OP_102J5_124_3590_n702,
         DP_OP_102J5_124_3590_n701, DP_OP_102J5_124_3590_n700,
         DP_OP_102J5_124_3590_n699, DP_OP_102J5_124_3590_n698,
         DP_OP_102J5_124_3590_n697, DP_OP_102J5_124_3590_n696,
         DP_OP_102J5_124_3590_n695, DP_OP_102J5_124_3590_n694,
         DP_OP_102J5_124_3590_n693, DP_OP_102J5_124_3590_n692,
         DP_OP_102J5_124_3590_n691, DP_OP_102J5_124_3590_n690,
         DP_OP_102J5_124_3590_n689, DP_OP_102J5_124_3590_n688,
         DP_OP_102J5_124_3590_n687, DP_OP_102J5_124_3590_n686,
         DP_OP_102J5_124_3590_n685, DP_OP_102J5_124_3590_n684,
         DP_OP_102J5_124_3590_n683, DP_OP_102J5_124_3590_n682,
         DP_OP_102J5_124_3590_n681, DP_OP_102J5_124_3590_n680,
         DP_OP_102J5_124_3590_n679, DP_OP_102J5_124_3590_n678,
         DP_OP_102J5_124_3590_n677, DP_OP_102J5_124_3590_n676,
         DP_OP_102J5_124_3590_n675, DP_OP_102J5_124_3590_n674,
         DP_OP_102J5_124_3590_n673, DP_OP_102J5_124_3590_n672,
         DP_OP_102J5_124_3590_n671, DP_OP_102J5_124_3590_n670,
         DP_OP_102J5_124_3590_n669, DP_OP_102J5_124_3590_n668,
         DP_OP_102J5_124_3590_n667, DP_OP_102J5_124_3590_n666,
         DP_OP_102J5_124_3590_n665, DP_OP_102J5_124_3590_n664,
         DP_OP_102J5_124_3590_n663, DP_OP_102J5_124_3590_n662,
         DP_OP_102J5_124_3590_n661, DP_OP_102J5_124_3590_n660,
         DP_OP_102J5_124_3590_n659, DP_OP_102J5_124_3590_n658,
         DP_OP_102J5_124_3590_n657, DP_OP_102J5_124_3590_n656,
         DP_OP_102J5_124_3590_n655, DP_OP_102J5_124_3590_n654,
         DP_OP_102J5_124_3590_n653, DP_OP_102J5_124_3590_n652,
         DP_OP_102J5_124_3590_n651, DP_OP_102J5_124_3590_n650,
         DP_OP_102J5_124_3590_n649, DP_OP_102J5_124_3590_n648,
         DP_OP_102J5_124_3590_n647, DP_OP_102J5_124_3590_n646,
         DP_OP_102J5_124_3590_n645, DP_OP_102J5_124_3590_n644,
         DP_OP_102J5_124_3590_n643, DP_OP_102J5_124_3590_n642,
         DP_OP_102J5_124_3590_n641, DP_OP_102J5_124_3590_n640,
         DP_OP_102J5_124_3590_n639, DP_OP_102J5_124_3590_n638,
         DP_OP_102J5_124_3590_n637, DP_OP_102J5_124_3590_n636,
         DP_OP_102J5_124_3590_n635, DP_OP_102J5_124_3590_n634,
         DP_OP_102J5_124_3590_n633, DP_OP_102J5_124_3590_n632,
         DP_OP_102J5_124_3590_n631, DP_OP_102J5_124_3590_n630,
         DP_OP_102J5_124_3590_n629, DP_OP_102J5_124_3590_n628,
         DP_OP_102J5_124_3590_n627, DP_OP_102J5_124_3590_n626,
         DP_OP_102J5_124_3590_n625, DP_OP_102J5_124_3590_n624,
         DP_OP_102J5_124_3590_n623, DP_OP_102J5_124_3590_n622,
         DP_OP_102J5_124_3590_n621, DP_OP_102J5_124_3590_n620,
         DP_OP_102J5_124_3590_n619, DP_OP_102J5_124_3590_n618,
         DP_OP_102J5_124_3590_n617, DP_OP_102J5_124_3590_n616,
         DP_OP_102J5_124_3590_n615, DP_OP_102J5_124_3590_n614,
         DP_OP_102J5_124_3590_n613, DP_OP_102J5_124_3590_n612,
         DP_OP_102J5_124_3590_n611, DP_OP_102J5_124_3590_n610,
         DP_OP_102J5_124_3590_n609, DP_OP_102J5_124_3590_n608,
         DP_OP_102J5_124_3590_n607, DP_OP_102J5_124_3590_n606,
         DP_OP_102J5_124_3590_n605, DP_OP_102J5_124_3590_n604,
         DP_OP_102J5_124_3590_n603, DP_OP_102J5_124_3590_n602,
         DP_OP_102J5_124_3590_n601, DP_OP_102J5_124_3590_n600,
         DP_OP_102J5_124_3590_n599, DP_OP_102J5_124_3590_n598,
         DP_OP_102J5_124_3590_n597, DP_OP_102J5_124_3590_n596,
         DP_OP_102J5_124_3590_n595, DP_OP_102J5_124_3590_n594,
         DP_OP_102J5_124_3590_n593, DP_OP_102J5_124_3590_n592,
         DP_OP_102J5_124_3590_n591, DP_OP_102J5_124_3590_n590,
         DP_OP_102J5_124_3590_n589, DP_OP_102J5_124_3590_n588,
         DP_OP_102J5_124_3590_n587, DP_OP_102J5_124_3590_n586,
         DP_OP_102J5_124_3590_n585, DP_OP_102J5_124_3590_n584,
         DP_OP_102J5_124_3590_n583, DP_OP_102J5_124_3590_n582,
         DP_OP_102J5_124_3590_n581, DP_OP_102J5_124_3590_n580,
         DP_OP_102J5_124_3590_n579, DP_OP_102J5_124_3590_n578,
         DP_OP_102J5_124_3590_n577, DP_OP_102J5_124_3590_n576,
         DP_OP_102J5_124_3590_n575, DP_OP_102J5_124_3590_n574,
         DP_OP_102J5_124_3590_n573, DP_OP_102J5_124_3590_n572,
         DP_OP_102J5_124_3590_n571, DP_OP_102J5_124_3590_n570,
         DP_OP_102J5_124_3590_n569, DP_OP_102J5_124_3590_n568,
         DP_OP_102J5_124_3590_n567, DP_OP_102J5_124_3590_n566,
         DP_OP_102J5_124_3590_n565, DP_OP_102J5_124_3590_n564,
         DP_OP_102J5_124_3590_n563, DP_OP_102J5_124_3590_n562,
         DP_OP_102J5_124_3590_n561, DP_OP_102J5_124_3590_n560,
         DP_OP_102J5_124_3590_n559, DP_OP_102J5_124_3590_n558,
         DP_OP_102J5_124_3590_n557, DP_OP_102J5_124_3590_n556,
         DP_OP_102J5_124_3590_n555, DP_OP_102J5_124_3590_n554,
         DP_OP_102J5_124_3590_n553, DP_OP_102J5_124_3590_n552,
         DP_OP_102J5_124_3590_n551, DP_OP_102J5_124_3590_n550,
         DP_OP_102J5_124_3590_n549, DP_OP_102J5_124_3590_n548,
         DP_OP_102J5_124_3590_n547, DP_OP_102J5_124_3590_n546,
         DP_OP_102J5_124_3590_n545, DP_OP_102J5_124_3590_n544,
         DP_OP_102J5_124_3590_n543, DP_OP_102J5_124_3590_n542,
         DP_OP_102J5_124_3590_n541, DP_OP_102J5_124_3590_n540,
         DP_OP_102J5_124_3590_n539, DP_OP_102J5_124_3590_n538,
         DP_OP_102J5_124_3590_n537, DP_OP_102J5_124_3590_n536,
         DP_OP_102J5_124_3590_n535, DP_OP_102J5_124_3590_n534,
         DP_OP_102J5_124_3590_n533, DP_OP_102J5_124_3590_n532,
         DP_OP_102J5_124_3590_n531, DP_OP_102J5_124_3590_n530,
         DP_OP_102J5_124_3590_n529, DP_OP_102J5_124_3590_n528,
         DP_OP_102J5_124_3590_n527, DP_OP_102J5_124_3590_n526,
         DP_OP_102J5_124_3590_n525, DP_OP_102J5_124_3590_n524,
         DP_OP_102J5_124_3590_n523, DP_OP_102J5_124_3590_n522,
         DP_OP_102J5_124_3590_n521, DP_OP_102J5_124_3590_n520,
         DP_OP_102J5_124_3590_n519, DP_OP_102J5_124_3590_n518,
         DP_OP_102J5_124_3590_n517, DP_OP_102J5_124_3590_n516,
         DP_OP_102J5_124_3590_n515, DP_OP_102J5_124_3590_n514,
         DP_OP_102J5_124_3590_n513, DP_OP_102J5_124_3590_n512,
         DP_OP_102J5_124_3590_n511, DP_OP_102J5_124_3590_n510,
         DP_OP_102J5_124_3590_n509, DP_OP_102J5_124_3590_n508,
         DP_OP_102J5_124_3590_n507, DP_OP_102J5_124_3590_n506,
         DP_OP_102J5_124_3590_n505, DP_OP_102J5_124_3590_n504,
         DP_OP_102J5_124_3590_n503, DP_OP_102J5_124_3590_n502,
         DP_OP_102J5_124_3590_n501, DP_OP_102J5_124_3590_n500,
         DP_OP_102J5_124_3590_n499, DP_OP_102J5_124_3590_n498,
         DP_OP_102J5_124_3590_n497, DP_OP_102J5_124_3590_n496,
         DP_OP_102J5_124_3590_n495, DP_OP_102J5_124_3590_n494,
         DP_OP_102J5_124_3590_n493, DP_OP_102J5_124_3590_n492,
         DP_OP_102J5_124_3590_n491, DP_OP_102J5_124_3590_n490,
         DP_OP_102J5_124_3590_n489, DP_OP_102J5_124_3590_n488,
         DP_OP_102J5_124_3590_n487, DP_OP_102J5_124_3590_n486,
         DP_OP_102J5_124_3590_n485, DP_OP_102J5_124_3590_n484,
         DP_OP_102J5_124_3590_n483, DP_OP_102J5_124_3590_n482,
         DP_OP_102J5_124_3590_n481, DP_OP_102J5_124_3590_n480,
         DP_OP_102J5_124_3590_n479, DP_OP_102J5_124_3590_n478,
         DP_OP_102J5_124_3590_n477, DP_OP_102J5_124_3590_n476,
         DP_OP_102J5_124_3590_n475, DP_OP_102J5_124_3590_n474,
         DP_OP_102J5_124_3590_n473, DP_OP_102J5_124_3590_n472,
         DP_OP_102J5_124_3590_n471, DP_OP_102J5_124_3590_n470,
         DP_OP_102J5_124_3590_n469, DP_OP_102J5_124_3590_n468,
         DP_OP_102J5_124_3590_n467, DP_OP_102J5_124_3590_n466,
         DP_OP_102J5_124_3590_n465, DP_OP_102J5_124_3590_n464,
         DP_OP_102J5_124_3590_n463, DP_OP_102J5_124_3590_n462,
         DP_OP_102J5_124_3590_n461, DP_OP_102J5_124_3590_n460,
         DP_OP_102J5_124_3590_n459, DP_OP_102J5_124_3590_n458,
         DP_OP_102J5_124_3590_n457, DP_OP_102J5_124_3590_n456,
         DP_OP_102J5_124_3590_n455, DP_OP_102J5_124_3590_n454,
         DP_OP_102J5_124_3590_n453, DP_OP_102J5_124_3590_n452,
         DP_OP_102J5_124_3590_n451, DP_OP_102J5_124_3590_n450,
         DP_OP_102J5_124_3590_n449, DP_OP_102J5_124_3590_n448,
         DP_OP_102J5_124_3590_n447, DP_OP_102J5_124_3590_n446,
         DP_OP_102J5_124_3590_n445, DP_OP_102J5_124_3590_n444,
         DP_OP_102J5_124_3590_n443, DP_OP_102J5_124_3590_n442,
         DP_OP_102J5_124_3590_n441, DP_OP_102J5_124_3590_n440,
         DP_OP_102J5_124_3590_n439, DP_OP_102J5_124_3590_n438,
         DP_OP_102J5_124_3590_n437, DP_OP_102J5_124_3590_n436,
         DP_OP_102J5_124_3590_n435, DP_OP_102J5_124_3590_n434,
         DP_OP_102J5_124_3590_n433, DP_OP_102J5_124_3590_n432,
         DP_OP_102J5_124_3590_n431, DP_OP_102J5_124_3590_n430,
         DP_OP_102J5_124_3590_n429, DP_OP_102J5_124_3590_n428,
         DP_OP_102J5_124_3590_n427, DP_OP_102J5_124_3590_n426,
         DP_OP_102J5_124_3590_n425, DP_OP_102J5_124_3590_n424,
         DP_OP_102J5_124_3590_n423, DP_OP_102J5_124_3590_n422,
         DP_OP_102J5_124_3590_n421, DP_OP_102J5_124_3590_n420,
         DP_OP_102J5_124_3590_n419, DP_OP_102J5_124_3590_n418,
         DP_OP_102J5_124_3590_n417, DP_OP_102J5_124_3590_n416,
         DP_OP_102J5_124_3590_n415, DP_OP_102J5_124_3590_n414,
         DP_OP_102J5_124_3590_n413, DP_OP_102J5_124_3590_n412,
         DP_OP_102J5_124_3590_n411, DP_OP_102J5_124_3590_n410,
         DP_OP_102J5_124_3590_n409, DP_OP_102J5_124_3590_n408,
         DP_OP_102J5_124_3590_n407, DP_OP_102J5_124_3590_n406,
         DP_OP_102J5_124_3590_n405, DP_OP_102J5_124_3590_n404,
         DP_OP_102J5_124_3590_n403, DP_OP_102J5_124_3590_n402,
         DP_OP_102J5_124_3590_n401, DP_OP_102J5_124_3590_n400,
         DP_OP_102J5_124_3590_n399, DP_OP_102J5_124_3590_n398,
         DP_OP_102J5_124_3590_n397, DP_OP_102J5_124_3590_n396,
         DP_OP_102J5_124_3590_n395, DP_OP_102J5_124_3590_n394,
         DP_OP_102J5_124_3590_n393, DP_OP_102J5_124_3590_n392,
         DP_OP_102J5_124_3590_n391, DP_OP_102J5_124_3590_n390,
         DP_OP_102J5_124_3590_n389, DP_OP_102J5_124_3590_n388,
         DP_OP_102J5_124_3590_n387, DP_OP_102J5_124_3590_n386,
         DP_OP_102J5_124_3590_n385, DP_OP_102J5_124_3590_n384,
         DP_OP_102J5_124_3590_n383, DP_OP_102J5_124_3590_n382,
         DP_OP_102J5_124_3590_n381, DP_OP_102J5_124_3590_n380,
         DP_OP_102J5_124_3590_n379, DP_OP_102J5_124_3590_n378,
         DP_OP_102J5_124_3590_n377, DP_OP_102J5_124_3590_n376,
         DP_OP_102J5_124_3590_n375, DP_OP_102J5_124_3590_n374,
         DP_OP_102J5_124_3590_n373, DP_OP_102J5_124_3590_n372,
         DP_OP_102J5_124_3590_n371, DP_OP_102J5_124_3590_n370,
         DP_OP_102J5_124_3590_n369, DP_OP_102J5_124_3590_n368,
         DP_OP_102J5_124_3590_n367, DP_OP_102J5_124_3590_n366,
         DP_OP_102J5_124_3590_n365, DP_OP_102J5_124_3590_n364,
         DP_OP_102J5_124_3590_n363, DP_OP_102J5_124_3590_n362,
         DP_OP_102J5_124_3590_n361, DP_OP_102J5_124_3590_n360,
         DP_OP_102J5_124_3590_n359, DP_OP_102J5_124_3590_n358,
         DP_OP_102J5_124_3590_n357, DP_OP_102J5_124_3590_n356,
         DP_OP_102J5_124_3590_n355, DP_OP_102J5_124_3590_n354,
         DP_OP_102J5_124_3590_n353, DP_OP_102J5_124_3590_n352,
         DP_OP_102J5_124_3590_n351, DP_OP_102J5_124_3590_n350,
         DP_OP_102J5_124_3590_n349, DP_OP_102J5_124_3590_n348,
         DP_OP_102J5_124_3590_n347, DP_OP_102J5_124_3590_n346,
         DP_OP_102J5_124_3590_n345, DP_OP_102J5_124_3590_n344,
         DP_OP_102J5_124_3590_n343, DP_OP_102J5_124_3590_n342,
         DP_OP_102J5_124_3590_n341, DP_OP_102J5_124_3590_n340,
         DP_OP_102J5_124_3590_n339, DP_OP_102J5_124_3590_n338,
         DP_OP_102J5_124_3590_n337, DP_OP_102J5_124_3590_n336,
         DP_OP_102J5_124_3590_n335, DP_OP_102J5_124_3590_n334,
         DP_OP_102J5_124_3590_n333, DP_OP_102J5_124_3590_n332,
         DP_OP_102J5_124_3590_n331, DP_OP_102J5_124_3590_n330,
         DP_OP_102J5_124_3590_n329, DP_OP_102J5_124_3590_n328,
         DP_OP_102J5_124_3590_n327, DP_OP_102J5_124_3590_n326,
         DP_OP_102J5_124_3590_n325, DP_OP_102J5_124_3590_n324,
         DP_OP_102J5_124_3590_n323, DP_OP_102J5_124_3590_n322,
         DP_OP_102J5_124_3590_n321, DP_OP_102J5_124_3590_n320,
         DP_OP_102J5_124_3590_n319, DP_OP_102J5_124_3590_n318,
         DP_OP_102J5_124_3590_n317, DP_OP_102J5_124_3590_n316,
         DP_OP_102J5_124_3590_n315, DP_OP_102J5_124_3590_n314,
         DP_OP_102J5_124_3590_n313, DP_OP_102J5_124_3590_n312,
         DP_OP_102J5_124_3590_n311, DP_OP_102J5_124_3590_n310,
         DP_OP_102J5_124_3590_n309, DP_OP_102J5_124_3590_n308,
         DP_OP_102J5_124_3590_n307, DP_OP_102J5_124_3590_n306,
         DP_OP_102J5_124_3590_n305, DP_OP_102J5_124_3590_n304,
         DP_OP_102J5_124_3590_n303, DP_OP_102J5_124_3590_n302,
         DP_OP_102J5_124_3590_n301, DP_OP_102J5_124_3590_n300,
         DP_OP_102J5_124_3590_n299, DP_OP_102J5_124_3590_n298,
         DP_OP_102J5_124_3590_n297, DP_OP_102J5_124_3590_n296,
         DP_OP_102J5_124_3590_n295, DP_OP_102J5_124_3590_n294,
         DP_OP_102J5_124_3590_n293, DP_OP_102J5_124_3590_n292,
         DP_OP_102J5_124_3590_n291, DP_OP_102J5_124_3590_n290,
         DP_OP_102J5_124_3590_n289, DP_OP_102J5_124_3590_n288,
         DP_OP_102J5_124_3590_n287, DP_OP_102J5_124_3590_n286,
         DP_OP_102J5_124_3590_n285, DP_OP_102J5_124_3590_n284,
         DP_OP_102J5_124_3590_n283, DP_OP_102J5_124_3590_n282,
         DP_OP_102J5_124_3590_n281, DP_OP_102J5_124_3590_n280,
         DP_OP_102J5_124_3590_n279, DP_OP_102J5_124_3590_n278,
         DP_OP_102J5_124_3590_n277, DP_OP_102J5_124_3590_n276,
         DP_OP_102J5_124_3590_n275, DP_OP_102J5_124_3590_n274,
         DP_OP_102J5_124_3590_n273, DP_OP_102J5_124_3590_n272,
         DP_OP_102J5_124_3590_n271, DP_OP_102J5_124_3590_n270,
         DP_OP_102J5_124_3590_n269, DP_OP_102J5_124_3590_n268,
         DP_OP_102J5_124_3590_n267, DP_OP_102J5_124_3590_n266,
         DP_OP_102J5_124_3590_n265, DP_OP_102J5_124_3590_n264,
         DP_OP_102J5_124_3590_n263, DP_OP_102J5_124_3590_n262,
         DP_OP_102J5_124_3590_n261, DP_OP_102J5_124_3590_n260,
         DP_OP_102J5_124_3590_n259, DP_OP_102J5_124_3590_n258,
         DP_OP_102J5_124_3590_n257, DP_OP_102J5_124_3590_n256,
         DP_OP_102J5_124_3590_n255, DP_OP_102J5_124_3590_n254,
         DP_OP_102J5_124_3590_n253, DP_OP_102J5_124_3590_n252,
         DP_OP_102J5_124_3590_n251, DP_OP_102J5_124_3590_n250,
         DP_OP_102J5_124_3590_n249, DP_OP_102J5_124_3590_n248,
         DP_OP_102J5_124_3590_n247, DP_OP_102J5_124_3590_n246,
         DP_OP_102J5_124_3590_n245, DP_OP_102J5_124_3590_n244,
         DP_OP_102J5_124_3590_n243, DP_OP_102J5_124_3590_n242,
         DP_OP_102J5_124_3590_n241, DP_OP_102J5_124_3590_n240,
         DP_OP_102J5_124_3590_n239, DP_OP_102J5_124_3590_n238,
         DP_OP_102J5_124_3590_n237, DP_OP_102J5_124_3590_n236,
         DP_OP_102J5_124_3590_n235, DP_OP_102J5_124_3590_n234,
         DP_OP_102J5_124_3590_n233, DP_OP_102J5_124_3590_n232,
         DP_OP_102J5_124_3590_n231, DP_OP_102J5_124_3590_n230,
         DP_OP_102J5_124_3590_n229, DP_OP_102J5_124_3590_n228,
         DP_OP_102J5_124_3590_n227, DP_OP_102J5_124_3590_n226,
         DP_OP_102J5_124_3590_n225, DP_OP_102J5_124_3590_n224,
         DP_OP_102J5_124_3590_n223, DP_OP_102J5_124_3590_n222,
         DP_OP_102J5_124_3590_n221, DP_OP_102J5_124_3590_n220,
         DP_OP_102J5_124_3590_n219, DP_OP_102J5_124_3590_n218,
         DP_OP_102J5_124_3590_n217, DP_OP_102J5_124_3590_n216,
         DP_OP_102J5_124_3590_n215, DP_OP_102J5_124_3590_n214,
         DP_OP_102J5_124_3590_n213, DP_OP_102J5_124_3590_n212,
         DP_OP_102J5_124_3590_n211, DP_OP_102J5_124_3590_n210,
         DP_OP_102J5_124_3590_n209, DP_OP_102J5_124_3590_n208,
         DP_OP_102J5_124_3590_n207, DP_OP_102J5_124_3590_n206,
         DP_OP_102J5_124_3590_n205, DP_OP_102J5_124_3590_n204,
         DP_OP_102J5_124_3590_n203, DP_OP_102J5_124_3590_n202,
         DP_OP_102J5_124_3590_n201, DP_OP_102J5_124_3590_n200,
         DP_OP_102J5_124_3590_n199, DP_OP_102J5_124_3590_n198,
         DP_OP_102J5_124_3590_n197, DP_OP_102J5_124_3590_n196,
         DP_OP_102J5_124_3590_n195, DP_OP_102J5_124_3590_n194,
         DP_OP_102J5_124_3590_n193, DP_OP_102J5_124_3590_n192,
         DP_OP_102J5_124_3590_n191, DP_OP_102J5_124_3590_n190,
         DP_OP_102J5_124_3590_n189, DP_OP_102J5_124_3590_n188,
         DP_OP_102J5_124_3590_n187, DP_OP_102J5_124_3590_n186,
         DP_OP_102J5_124_3590_n176, DP_OP_102J5_124_3590_n162,
         DP_OP_102J5_124_3590_n161, DP_OP_102J5_124_3590_n160,
         DP_OP_102J5_124_3590_n159, DP_OP_102J5_124_3590_n158,
         DP_OP_102J5_124_3590_n152, DP_OP_102J5_124_3590_n148,
         DP_OP_102J5_124_3590_n147, DP_OP_102J5_124_3590_n146,
         DP_OP_102J5_124_3590_n145, DP_OP_102J5_124_3590_n144,
         DP_OP_102J5_124_3590_n140, DP_OP_102J5_124_3590_n139,
         DP_OP_102J5_124_3590_n138, DP_OP_102J5_124_3590_n137,
         DP_OP_102J5_124_3590_n136, DP_OP_102J5_124_3590_n135,
         DP_OP_102J5_124_3590_n134, DP_OP_102J5_124_3590_n132,
         DP_OP_102J5_124_3590_n131, DP_OP_102J5_124_3590_n128,
         DP_OP_102J5_124_3590_n127, DP_OP_102J5_124_3590_n126,
         DP_OP_102J5_124_3590_n125, DP_OP_102J5_124_3590_n121,
         DP_OP_102J5_124_3590_n120, DP_OP_102J5_124_3590_n119,
         DP_OP_102J5_124_3590_n118, DP_OP_102J5_124_3590_n117,
         DP_OP_102J5_124_3590_n116, DP_OP_102J5_124_3590_n115,
         DP_OP_102J5_124_3590_n113, DP_OP_102J5_124_3590_n112,
         DP_OP_102J5_124_3590_n106, DP_OP_102J5_124_3590_n105,
         DP_OP_102J5_124_3590_n104, DP_OP_102J5_124_3590_n99,
         DP_OP_102J5_124_3590_n98, DP_OP_102J5_124_3590_n97,
         DP_OP_102J5_124_3590_n96, DP_OP_102J5_124_3590_n95,
         DP_OP_102J5_124_3590_n94, DP_OP_102J5_124_3590_n93,
         DP_OP_102J5_124_3590_n91, DP_OP_102J5_124_3590_n89,
         DP_OP_102J5_124_3590_n85, DP_OP_102J5_124_3590_n84,
         DP_OP_102J5_124_3590_n77, DP_OP_102J5_124_3590_n76,
         DP_OP_102J5_124_3590_n75, DP_OP_102J5_124_3590_n71,
         DP_OP_102J5_124_3590_n67, DP_OP_102J5_124_3590_n64,
         DP_OP_102J5_124_3590_n60, DP_OP_102J5_124_3590_n59,
         DP_OP_102J5_124_3590_n57, DP_OP_102J5_124_3590_n56,
         DP_OP_102J5_124_3590_n53, DP_OP_102J5_124_3590_n49,
         DP_OP_102J5_124_3590_n48, DP_OP_102J5_124_3590_n46,
         DP_OP_102J5_124_3590_n44, DP_OP_102J5_124_3590_n43,
         DP_OP_102J5_124_3590_n42, DP_OP_102J5_124_3590_n40,
         DP_OP_102J5_124_3590_n36, DP_OP_102J5_124_3590_n35,
         DP_OP_102J5_124_3590_n31, DP_OP_102J5_124_3590_n30,
         DP_OP_102J5_124_3590_n5, DP_OP_102J5_124_3590_n3, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n140, n141,
         n142, n143, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301;
  wire   [22:0] n_accumulator_sum;

  DFFSSRX1_HVT fc_weight_box_reg_0__3_ ( .D(1'b0), .SETB(n189), .RSTB(
        sram_rdata_weight[79]), .CLK(clk), .QN(n207) );
  DFFSSRX1_HVT fc_weight_box_reg_0__2_ ( .D(1'b0), .SETB(n188), .RSTB(
        sram_rdata_weight[78]), .CLK(clk), .QN(n245) );
  DFFSSRX1_HVT fc_weight_box_reg_0__1_ ( .D(1'b0), .SETB(n187), .RSTB(
        sram_rdata_weight[77]), .CLK(clk), .QN(n246) );
  DFFSSRX1_HVT fc_weight_box_reg_0__0_ ( .D(1'b0), .SETB(n190), .RSTB(
        sram_rdata_weight[76]), .CLK(clk), .QN(n247) );
  DFFSSRX1_HVT fc_weight_box_reg_1__3_ ( .D(1'b0), .SETB(n189), .RSTB(
        sram_rdata_weight[75]), .CLK(clk), .QN(n208) );
  DFFSSRX1_HVT fc_weight_box_reg_1__2_ ( .D(1'b0), .SETB(n188), .RSTB(
        sram_rdata_weight[74]), .CLK(clk), .QN(n248) );
  DFFSSRX1_HVT fc_weight_box_reg_1__1_ ( .D(1'b0), .SETB(n187), .RSTB(
        sram_rdata_weight[73]), .CLK(clk), .QN(n249) );
  DFFSSRX1_HVT fc_weight_box_reg_1__0_ ( .D(1'b0), .SETB(n190), .RSTB(
        sram_rdata_weight[72]), .CLK(clk), .QN(n250) );
  DFFSSRX1_HVT fc_weight_box_reg_2__3_ ( .D(1'b0), .SETB(n189), .RSTB(
        sram_rdata_weight[71]), .CLK(clk), .QN(n206) );
  DFFSSRX1_HVT fc_weight_box_reg_2__2_ ( .D(1'b0), .SETB(n188), .RSTB(
        sram_rdata_weight[70]), .CLK(clk), .QN(n242) );
  DFFSSRX1_HVT fc_weight_box_reg_2__1_ ( .D(1'b0), .SETB(n187), .RSTB(
        sram_rdata_weight[69]), .CLK(clk), .QN(n243) );
  DFFSSRX1_HVT fc_weight_box_reg_2__0_ ( .D(1'b0), .SETB(n190), .RSTB(
        sram_rdata_weight[68]), .CLK(clk), .QN(n244) );
  DFFSSRX1_HVT fc_weight_box_reg_3__3_ ( .D(1'b0), .SETB(n189), .RSTB(
        sram_rdata_weight[67]), .CLK(clk), .QN(n209) );
  DFFSSRX1_HVT fc_weight_box_reg_3__2_ ( .D(1'b0), .SETB(n188), .RSTB(
        sram_rdata_weight[66]), .CLK(clk), .QN(n251) );
  DFFSSRX1_HVT fc_weight_box_reg_3__1_ ( .D(1'b0), .SETB(n187), .RSTB(
        sram_rdata_weight[65]), .CLK(clk), .QN(n252) );
  DFFSSRX1_HVT fc_weight_box_reg_3__0_ ( .D(1'b0), .SETB(n190), .RSTB(
        sram_rdata_weight[64]), .CLK(clk), .QN(n253) );
  DFFSSRX1_HVT fc_weight_box_reg_4__3_ ( .D(1'b0), .SETB(n189), .RSTB(
        sram_rdata_weight[63]), .CLK(clk), .QN(n205) );
  DFFSSRX1_HVT fc_weight_box_reg_4__2_ ( .D(1'b0), .SETB(n188), .RSTB(
        sram_rdata_weight[62]), .CLK(clk), .QN(n239) );
  DFFSSRX1_HVT fc_weight_box_reg_4__1_ ( .D(1'b0), .SETB(n187), .RSTB(
        sram_rdata_weight[61]), .CLK(clk), .QN(n240) );
  DFFSSRX1_HVT fc_weight_box_reg_4__0_ ( .D(1'b0), .SETB(n190), .RSTB(
        sram_rdata_weight[60]), .CLK(clk), .QN(n241) );
  DFFSSRX1_HVT fc_weight_box_reg_5__3_ ( .D(1'b0), .SETB(n189), .RSTB(
        sram_rdata_weight[59]), .CLK(clk), .QN(n210) );
  DFFSSRX1_HVT fc_weight_box_reg_5__2_ ( .D(1'b0), .SETB(n188), .RSTB(
        sram_rdata_weight[58]), .CLK(clk), .QN(n254) );
  DFFSSRX1_HVT fc_weight_box_reg_5__1_ ( .D(1'b0), .SETB(n187), .RSTB(
        sram_rdata_weight[57]), .CLK(clk), .QN(n255) );
  DFFSSRX1_HVT fc_weight_box_reg_5__0_ ( .D(1'b0), .SETB(n190), .RSTB(
        sram_rdata_weight[56]), .CLK(clk), .QN(n256) );
  DFFSSRX1_HVT fc_weight_box_reg_6__3_ ( .D(1'b0), .SETB(n189), .RSTB(
        sram_rdata_weight[55]), .CLK(clk), .QN(n204) );
  DFFSSRX1_HVT fc_weight_box_reg_6__2_ ( .D(1'b0), .SETB(n188), .RSTB(
        sram_rdata_weight[54]), .CLK(clk), .QN(n236) );
  DFFSSRX1_HVT fc_weight_box_reg_6__1_ ( .D(1'b0), .SETB(n187), .RSTB(
        sram_rdata_weight[53]), .CLK(clk), .QN(n237) );
  DFFSSRX1_HVT fc_weight_box_reg_6__0_ ( .D(1'b0), .SETB(n190), .RSTB(
        sram_rdata_weight[52]), .CLK(clk), .QN(n238) );
  DFFSSRX1_HVT fc_weight_box_reg_7__3_ ( .D(1'b0), .SETB(n189), .RSTB(
        sram_rdata_weight[51]), .CLK(clk), .QN(n211) );
  DFFSSRX1_HVT fc_weight_box_reg_7__2_ ( .D(1'b0), .SETB(n188), .RSTB(
        sram_rdata_weight[50]), .CLK(clk), .QN(n257) );
  DFFSSRX1_HVT fc_weight_box_reg_7__1_ ( .D(1'b0), .SETB(n187), .RSTB(
        sram_rdata_weight[49]), .CLK(clk), .QN(n258) );
  DFFSSRX1_HVT fc_weight_box_reg_7__0_ ( .D(1'b0), .SETB(n190), .RSTB(
        sram_rdata_weight[48]), .CLK(clk), .QN(n259) );
  DFFSSRX1_HVT fc_weight_box_reg_8__3_ ( .D(1'b0), .SETB(n189), .RSTB(
        sram_rdata_weight[47]), .CLK(clk), .QN(n203) );
  DFFSSRX1_HVT fc_weight_box_reg_8__2_ ( .D(1'b0), .SETB(n188), .RSTB(
        sram_rdata_weight[46]), .CLK(clk), .QN(n233) );
  DFFSSRX1_HVT fc_weight_box_reg_8__1_ ( .D(1'b0), .SETB(n187), .RSTB(
        sram_rdata_weight[45]), .CLK(clk), .QN(n234) );
  DFFSSRX1_HVT fc_weight_box_reg_8__0_ ( .D(1'b0), .SETB(n190), .RSTB(
        sram_rdata_weight[44]), .CLK(clk), .QN(n235) );
  DFFSSRX1_HVT fc_weight_box_reg_9__3_ ( .D(1'b0), .SETB(n189), .RSTB(
        sram_rdata_weight[43]), .CLK(clk), .QN(n212) );
  DFFSSRX1_HVT fc_weight_box_reg_9__2_ ( .D(1'b0), .SETB(n188), .RSTB(
        sram_rdata_weight[42]), .CLK(clk), .QN(n260) );
  DFFSSRX1_HVT fc_weight_box_reg_9__1_ ( .D(1'b0), .SETB(n187), .RSTB(
        sram_rdata_weight[41]), .CLK(clk), .QN(n261) );
  DFFSSRX1_HVT fc_weight_box_reg_9__0_ ( .D(1'b0), .SETB(n190), .RSTB(
        sram_rdata_weight[40]), .CLK(clk), .QN(n262) );
  DFFSSRX1_HVT fc_weight_box_reg_10__3_ ( .D(1'b0), .SETB(n189), .RSTB(
        sram_rdata_weight[39]), .CLK(clk), .QN(n202) );
  DFFSSRX1_HVT fc_weight_box_reg_10__2_ ( .D(1'b0), .SETB(n188), .RSTB(
        sram_rdata_weight[38]), .CLK(clk), .QN(n230) );
  DFFSSRX1_HVT fc_weight_box_reg_10__1_ ( .D(1'b0), .SETB(n187), .RSTB(
        sram_rdata_weight[37]), .CLK(clk), .QN(n231) );
  DFFSSRX1_HVT fc_weight_box_reg_10__0_ ( .D(1'b0), .SETB(n190), .RSTB(
        sram_rdata_weight[36]), .CLK(clk), .QN(n232) );
  DFFSSRX1_HVT fc_weight_box_reg_11__3_ ( .D(1'b0), .SETB(n189), .RSTB(
        sram_rdata_weight[35]), .CLK(clk), .QN(n213) );
  DFFSSRX1_HVT fc_weight_box_reg_11__2_ ( .D(1'b0), .SETB(n188), .RSTB(
        sram_rdata_weight[34]), .CLK(clk), .QN(n263) );
  DFFSSRX1_HVT fc_weight_box_reg_11__1_ ( .D(1'b0), .SETB(n187), .RSTB(
        sram_rdata_weight[33]), .CLK(clk), .QN(n264) );
  DFFSSRX1_HVT fc_weight_box_reg_11__0_ ( .D(1'b0), .SETB(n190), .RSTB(
        sram_rdata_weight[32]), .CLK(clk), .QN(n265) );
  DFFSSRX1_HVT fc_weight_box_reg_12__3_ ( .D(1'b0), .SETB(n189), .RSTB(
        sram_rdata_weight[31]), .CLK(clk), .QN(n201) );
  DFFSSRX1_HVT fc_weight_box_reg_12__2_ ( .D(1'b0), .SETB(n188), .RSTB(
        sram_rdata_weight[30]), .CLK(clk), .QN(n227) );
  DFFSSRX1_HVT fc_weight_box_reg_12__1_ ( .D(1'b0), .SETB(n187), .RSTB(
        sram_rdata_weight[29]), .CLK(clk), .QN(n228) );
  DFFSSRX1_HVT fc_weight_box_reg_12__0_ ( .D(1'b0), .SETB(n190), .RSTB(
        sram_rdata_weight[28]), .CLK(clk), .QN(n229) );
  DFFSSRX1_HVT fc_weight_box_reg_13__3_ ( .D(1'b0), .SETB(n189), .RSTB(
        sram_rdata_weight[27]), .CLK(clk), .QN(n214) );
  DFFSSRX1_HVT fc_weight_box_reg_13__2_ ( .D(1'b0), .SETB(n188), .RSTB(
        sram_rdata_weight[26]), .CLK(clk), .QN(n266) );
  DFFSSRX1_HVT fc_weight_box_reg_13__1_ ( .D(1'b0), .SETB(n187), .RSTB(
        sram_rdata_weight[25]), .CLK(clk), .QN(n267) );
  DFFSSRX1_HVT fc_weight_box_reg_13__0_ ( .D(1'b0), .SETB(n190), .RSTB(
        sram_rdata_weight[24]), .CLK(clk), .QN(n268) );
  DFFSSRX1_HVT fc_weight_box_reg_14__3_ ( .D(1'b0), .SETB(n189), .RSTB(
        sram_rdata_weight[23]), .CLK(clk), .QN(n200) );
  DFFSSRX1_HVT fc_weight_box_reg_14__2_ ( .D(1'b0), .SETB(n188), .RSTB(
        sram_rdata_weight[22]), .CLK(clk), .QN(n224) );
  DFFSSRX1_HVT fc_weight_box_reg_14__1_ ( .D(1'b0), .SETB(n187), .RSTB(
        sram_rdata_weight[21]), .CLK(clk), .QN(n225) );
  DFFSSRX1_HVT fc_weight_box_reg_14__0_ ( .D(1'b0), .SETB(n190), .RSTB(
        sram_rdata_weight[20]), .CLK(clk), .QN(n226) );
  DFFSSRX1_HVT fc_weight_box_reg_15__3_ ( .D(1'b0), .SETB(n189), .RSTB(
        sram_rdata_weight[19]), .CLK(clk), .QN(n215) );
  DFFSSRX1_HVT fc_weight_box_reg_15__2_ ( .D(1'b0), .SETB(n188), .RSTB(
        sram_rdata_weight[18]), .CLK(clk), .QN(n269) );
  DFFSSRX1_HVT fc_weight_box_reg_15__1_ ( .D(1'b0), .SETB(n187), .RSTB(
        sram_rdata_weight[17]), .CLK(clk), .QN(n270) );
  DFFSSRX1_HVT fc_weight_box_reg_15__0_ ( .D(1'b0), .SETB(n190), .RSTB(
        sram_rdata_weight[16]), .CLK(clk), .QN(n271) );
  DFFSSRX1_HVT fc_weight_box_reg_16__3_ ( .D(1'b0), .SETB(n189), .RSTB(
        sram_rdata_weight[15]), .CLK(clk), .QN(n199) );
  DFFSSRX1_HVT fc_weight_box_reg_16__2_ ( .D(1'b0), .SETB(n188), .RSTB(
        sram_rdata_weight[14]), .CLK(clk), .QN(n221) );
  DFFSSRX1_HVT fc_weight_box_reg_16__1_ ( .D(1'b0), .SETB(n187), .RSTB(
        sram_rdata_weight[13]), .CLK(clk), .QN(n222) );
  DFFSSRX1_HVT fc_weight_box_reg_16__0_ ( .D(1'b0), .SETB(n190), .RSTB(
        sram_rdata_weight[12]), .CLK(clk), .QN(n223) );
  DFFSSRX1_HVT fc_weight_box_reg_17__3_ ( .D(1'b0), .SETB(n189), .RSTB(
        sram_rdata_weight[11]), .CLK(clk), .QN(n216) );
  DFFSSRX1_HVT fc_weight_box_reg_17__2_ ( .D(1'b0), .SETB(n188), .RSTB(
        sram_rdata_weight[10]), .CLK(clk), .QN(n272) );
  DFFSSRX1_HVT fc_weight_box_reg_17__1_ ( .D(1'b0), .SETB(n187), .RSTB(
        sram_rdata_weight[9]), .CLK(clk), .QN(n273) );
  DFFSSRX1_HVT fc_weight_box_reg_17__0_ ( .D(1'b0), .SETB(n190), .RSTB(
        sram_rdata_weight[8]), .CLK(clk), .QN(n274) );
  DFFSSRX1_HVT fc_weight_box_reg_18__3_ ( .D(1'b0), .SETB(n189), .RSTB(
        sram_rdata_weight[7]), .CLK(clk), .QN(n198) );
  DFFSSRX1_HVT fc_weight_box_reg_18__2_ ( .D(1'b0), .SETB(n188), .RSTB(
        sram_rdata_weight[6]), .CLK(clk), .QN(n218) );
  DFFSSRX1_HVT fc_weight_box_reg_18__1_ ( .D(1'b0), .SETB(n187), .RSTB(
        sram_rdata_weight[5]), .CLK(clk), .QN(n219) );
  DFFSSRX1_HVT fc_weight_box_reg_18__0_ ( .D(1'b0), .SETB(n190), .RSTB(
        sram_rdata_weight[4]), .CLK(clk), .QN(n220) );
  DFFSSRX1_HVT fc_weight_box_reg_19__3_ ( .D(1'b0), .SETB(n189), .RSTB(
        sram_rdata_weight[3]), .CLK(clk), .QN(n217) );
  DFFSSRX1_HVT fc_weight_box_reg_19__2_ ( .D(1'b0), .SETB(n188), .RSTB(
        sram_rdata_weight[2]), .CLK(clk), .QN(n275) );
  DFFSSRX1_HVT fc_weight_box_reg_19__1_ ( .D(1'b0), .SETB(n187), .RSTB(
        sram_rdata_weight[1]), .CLK(clk), .QN(n276) );
  DFFSSRX1_HVT fc_weight_box_reg_19__0_ ( .D(1'b0), .SETB(n188), .RSTB(
        sram_rdata_weight[0]), .CLK(clk), .QN(n277) );
  DFFSSRX1_HVT accumulator_sum_reg_22_ ( .D(1'b0), .SETB(n190), .RSTB(
        n_accumulator_sum[22]), .CLK(clk), .Q(data_out[22]), .QN(n301) );
  DFFSSRX1_HVT accumulator_sum_reg_21_ ( .D(1'b0), .SETB(n189), .RSTB(
        n_accumulator_sum[21]), .CLK(clk), .Q(data_out[21]), .QN(n300) );
  DFFSSRX1_HVT accumulator_sum_reg_20_ ( .D(1'b0), .SETB(n188), .RSTB(
        n_accumulator_sum[20]), .CLK(clk), .Q(data_out[20]), .QN(n197) );
  DFFSSRX1_HVT accumulator_sum_reg_19_ ( .D(1'b0), .SETB(n187), .RSTB(
        n_accumulator_sum[19]), .CLK(clk), .Q(data_out[19]), .QN(n299) );
  DFFSSRX1_HVT accumulator_sum_reg_18_ ( .D(1'b0), .SETB(n190), .RSTB(
        n_accumulator_sum[18]), .CLK(clk), .Q(data_out[18]), .QN(n289) );
  DFFSSRX1_HVT accumulator_sum_reg_17_ ( .D(1'b0), .SETB(n189), .RSTB(
        n_accumulator_sum[17]), .CLK(clk), .Q(data_out[17]), .QN(n196) );
  DFFSSRX1_HVT accumulator_sum_reg_16_ ( .D(1'b0), .SETB(n188), .RSTB(
        n_accumulator_sum[16]), .CLK(clk), .Q(data_out[16]), .QN(n288) );
  DFFSSRX1_HVT accumulator_sum_reg_15_ ( .D(1'b0), .SETB(n187), .RSTB(
        n_accumulator_sum[15]), .CLK(clk), .Q(data_out[15]), .QN(n298) );
  DFFSSRX1_HVT accumulator_sum_reg_14_ ( .D(1'b0), .SETB(n190), .RSTB(
        n_accumulator_sum[14]), .CLK(clk), .Q(data_out[14]), .QN(n287) );
  DFFSSRX1_HVT accumulator_sum_reg_13_ ( .D(1'b0), .SETB(n189), .RSTB(
        n_accumulator_sum[13]), .CLK(clk), .Q(data_out[13]), .QN(n297) );
  DFFSSRX1_HVT accumulator_sum_reg_12_ ( .D(1'b0), .SETB(n188), .RSTB(
        n_accumulator_sum[12]), .CLK(clk), .Q(data_out[12]), .QN(n193) );
  DFFSSRX1_HVT accumulator_sum_reg_11_ ( .D(1'b0), .SETB(n187), .RSTB(
        n_accumulator_sum[11]), .CLK(clk), .Q(data_out[11]), .QN(n194) );
  DFFSSRX1_HVT accumulator_sum_reg_10_ ( .D(1'b0), .SETB(n190), .RSTB(
        n_accumulator_sum[10]), .CLK(clk), .Q(data_out[10]), .QN(n292) );
  DFFSSRX1_HVT accumulator_sum_reg_9_ ( .D(1'b0), .SETB(n189), .RSTB(
        n_accumulator_sum[9]), .CLK(clk), .Q(data_out[9]), .QN(n295) );
  DFFSSRX1_HVT accumulator_sum_reg_8_ ( .D(1'b0), .SETB(n188), .RSTB(
        n_accumulator_sum[8]), .CLK(clk), .Q(data_out[8]), .QN(n195) );
  DFFSSRX1_HVT accumulator_sum_reg_7_ ( .D(1'b0), .SETB(n187), .RSTB(
        n_accumulator_sum[7]), .CLK(clk), .Q(data_out[7]), .QN(n296) );
  DFFSSRX1_HVT accumulator_sum_reg_6_ ( .D(1'b0), .SETB(n190), .RSTB(
        n_accumulator_sum[6]), .CLK(clk), .Q(data_out[6]), .QN(n293) );
  DFFSSRX1_HVT accumulator_sum_reg_5_ ( .D(1'b0), .SETB(n189), .RSTB(
        n_accumulator_sum[5]), .CLK(clk), .Q(data_out[5]), .QN(n294) );
  DFFSSRX1_HVT accumulator_sum_reg_4_ ( .D(1'b0), .SETB(n188), .RSTB(
        n_accumulator_sum[4]), .CLK(clk), .Q(data_out[4]), .QN(n278) );
  DFFSSRX1_HVT accumulator_sum_reg_3_ ( .D(1'b0), .SETB(n187), .RSTB(
        n_accumulator_sum[3]), .CLK(clk), .Q(data_out[3]), .QN(n280) );
  DFFSSRX1_HVT accumulator_sum_reg_2_ ( .D(1'b0), .SETB(n190), .RSTB(
        n_accumulator_sum[2]), .CLK(clk), .Q(data_out[2]), .QN(n281) );
  DFFSSRX1_HVT accumulator_sum_reg_1_ ( .D(1'b0), .SETB(n189), .RSTB(
        n_accumulator_sum[1]), .CLK(clk), .Q(data_out[1]), .QN(n282) );
  DFFSSRX1_HVT accumulator_sum_reg_0_ ( .D(1'b0), .SETB(n190), .RSTB(
        n_accumulator_sum[0]), .CLK(clk), .Q(data_out[0]), .QN(n283) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1764 ( .A1(n277), .A2(
        DP_OP_102J5_124_3590_n2379), .Y(DP_OP_102J5_124_3590_n2371) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1763 ( .A1(n277), .A2(
        DP_OP_102J5_124_3590_n2378), .Y(DP_OP_102J5_124_3590_n2370) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1762 ( .A1(n277), .A2(
        DP_OP_102J5_124_3590_n2377), .Y(DP_OP_102J5_124_3590_n2369) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1761 ( .A1(n277), .A2(
        DP_OP_102J5_124_3590_n2376), .Y(DP_OP_102J5_124_3590_n2368) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1760 ( .A1(n277), .A2(
        DP_OP_102J5_124_3590_n2375), .Y(DP_OP_102J5_124_3590_n2367) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1759 ( .A1(n277), .A2(
        DP_OP_102J5_124_3590_n2374), .Y(DP_OP_102J5_124_3590_n2366) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1758 ( .A1(n277), .A2(
        DP_OP_102J5_124_3590_n2373), .Y(DP_OP_102J5_124_3590_n2365) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1757 ( .A1(n277), .A2(
        DP_OP_102J5_124_3590_n2372), .Y(DP_OP_102J5_124_3590_n749) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1756 ( .A1(n276), .A2(
        DP_OP_102J5_124_3590_n2379), .Y(DP_OP_102J5_124_3590_n2364) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1755 ( .A1(n276), .A2(
        DP_OP_102J5_124_3590_n2378), .Y(DP_OP_102J5_124_3590_n2363) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1754 ( .A1(n276), .A2(
        DP_OP_102J5_124_3590_n2377), .Y(DP_OP_102J5_124_3590_n2362) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1753 ( .A1(n276), .A2(
        DP_OP_102J5_124_3590_n2376), .Y(DP_OP_102J5_124_3590_n2361) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1752 ( .A1(n276), .A2(
        DP_OP_102J5_124_3590_n2375), .Y(DP_OP_102J5_124_3590_n2360) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1751 ( .A1(n276), .A2(
        DP_OP_102J5_124_3590_n2374), .Y(DP_OP_102J5_124_3590_n2359) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1750 ( .A1(n276), .A2(
        DP_OP_102J5_124_3590_n2373), .Y(DP_OP_102J5_124_3590_n2358) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1749 ( .A1(n276), .A2(
        DP_OP_102J5_124_3590_n2372), .Y(DP_OP_102J5_124_3590_n2357) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1748 ( .A1(n275), .A2(
        DP_OP_102J5_124_3590_n2379), .Y(DP_OP_102J5_124_3590_n2356) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1747 ( .A1(n275), .A2(
        DP_OP_102J5_124_3590_n2378), .Y(DP_OP_102J5_124_3590_n2355) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1746 ( .A1(n275), .A2(
        DP_OP_102J5_124_3590_n2377), .Y(DP_OP_102J5_124_3590_n2354) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1745 ( .A1(n275), .A2(
        DP_OP_102J5_124_3590_n2376), .Y(DP_OP_102J5_124_3590_n2353) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1744 ( .A1(n275), .A2(
        DP_OP_102J5_124_3590_n2375), .Y(DP_OP_102J5_124_3590_n2352) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1743 ( .A1(n275), .A2(
        DP_OP_102J5_124_3590_n2374), .Y(DP_OP_102J5_124_3590_n2351) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1742 ( .A1(n275), .A2(
        DP_OP_102J5_124_3590_n2373), .Y(DP_OP_102J5_124_3590_n2350) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1741 ( .A1(n275), .A2(
        DP_OP_102J5_124_3590_n2372), .Y(DP_OP_102J5_124_3590_n2349) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1740 ( .A1(n217), .A2(
        DP_OP_102J5_124_3590_n2379), .Y(DP_OP_102J5_124_3590_n2348) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1739 ( .A1(n217), .A2(
        DP_OP_102J5_124_3590_n2378), .Y(DP_OP_102J5_124_3590_n2347) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1738 ( .A1(n217), .A2(
        DP_OP_102J5_124_3590_n2377), .Y(DP_OP_102J5_124_3590_n2346) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1737 ( .A1(n217), .A2(
        DP_OP_102J5_124_3590_n2376), .Y(DP_OP_102J5_124_3590_n2345) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1736 ( .A1(n217), .A2(
        DP_OP_102J5_124_3590_n2375), .Y(DP_OP_102J5_124_3590_n2344) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1735 ( .A1(n217), .A2(
        DP_OP_102J5_124_3590_n2374), .Y(DP_OP_102J5_124_3590_n2343) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1734 ( .A1(n217), .A2(
        DP_OP_102J5_124_3590_n2373), .Y(DP_OP_102J5_124_3590_n2342) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1733 ( .A1(n217), .A2(
        DP_OP_102J5_124_3590_n2372), .Y(DP_OP_102J5_124_3590_n2341) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1720 ( .A1(n274), .A2(
        DP_OP_102J5_124_3590_n2336), .Y(DP_OP_102J5_124_3590_n2328) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1719 ( .A1(n274), .A2(
        DP_OP_102J5_124_3590_n2335), .Y(DP_OP_102J5_124_3590_n2327) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1718 ( .A1(n274), .A2(
        DP_OP_102J5_124_3590_n2334), .Y(DP_OP_102J5_124_3590_n2326) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1717 ( .A1(n274), .A2(
        DP_OP_102J5_124_3590_n2333), .Y(DP_OP_102J5_124_3590_n2325) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1716 ( .A1(n274), .A2(
        DP_OP_102J5_124_3590_n2332), .Y(DP_OP_102J5_124_3590_n2324) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1715 ( .A1(n274), .A2(
        DP_OP_102J5_124_3590_n2331), .Y(DP_OP_102J5_124_3590_n2323) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1714 ( .A1(n274), .A2(
        DP_OP_102J5_124_3590_n2330), .Y(DP_OP_102J5_124_3590_n2322) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1713 ( .A1(n274), .A2(
        DP_OP_102J5_124_3590_n2329), .Y(DP_OP_102J5_124_3590_n2321) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1712 ( .A1(n273), .A2(
        DP_OP_102J5_124_3590_n2336), .Y(DP_OP_102J5_124_3590_n2320) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1711 ( .A1(n273), .A2(
        DP_OP_102J5_124_3590_n2335), .Y(DP_OP_102J5_124_3590_n2319) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1710 ( .A1(n273), .A2(
        DP_OP_102J5_124_3590_n2334), .Y(DP_OP_102J5_124_3590_n2318) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1709 ( .A1(n273), .A2(
        DP_OP_102J5_124_3590_n2333), .Y(DP_OP_102J5_124_3590_n2317) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1708 ( .A1(n273), .A2(
        DP_OP_102J5_124_3590_n2332), .Y(DP_OP_102J5_124_3590_n2316) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1707 ( .A1(n273), .A2(
        DP_OP_102J5_124_3590_n2331), .Y(DP_OP_102J5_124_3590_n2315) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1706 ( .A1(n273), .A2(
        DP_OP_102J5_124_3590_n2330), .Y(DP_OP_102J5_124_3590_n2314) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1705 ( .A1(n273), .A2(
        DP_OP_102J5_124_3590_n2329), .Y(DP_OP_102J5_124_3590_n2313) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1704 ( .A1(n272), .A2(
        DP_OP_102J5_124_3590_n2336), .Y(DP_OP_102J5_124_3590_n2312) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1703 ( .A1(n272), .A2(
        DP_OP_102J5_124_3590_n2335), .Y(DP_OP_102J5_124_3590_n2311) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1702 ( .A1(n272), .A2(
        DP_OP_102J5_124_3590_n2334), .Y(DP_OP_102J5_124_3590_n2310) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1701 ( .A1(n272), .A2(
        DP_OP_102J5_124_3590_n2333), .Y(DP_OP_102J5_124_3590_n2309) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1700 ( .A1(n272), .A2(
        DP_OP_102J5_124_3590_n2332), .Y(DP_OP_102J5_124_3590_n2308) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1699 ( .A1(n272), .A2(
        DP_OP_102J5_124_3590_n2331), .Y(DP_OP_102J5_124_3590_n2307) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1698 ( .A1(n272), .A2(
        DP_OP_102J5_124_3590_n2330), .Y(DP_OP_102J5_124_3590_n2306) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1697 ( .A1(n272), .A2(
        DP_OP_102J5_124_3590_n2329), .Y(DP_OP_102J5_124_3590_n2305) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1696 ( .A1(n216), .A2(
        DP_OP_102J5_124_3590_n2336), .Y(DP_OP_102J5_124_3590_n2304) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1695 ( .A1(n216), .A2(
        DP_OP_102J5_124_3590_n2335), .Y(DP_OP_102J5_124_3590_n2303) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1694 ( .A1(n216), .A2(
        DP_OP_102J5_124_3590_n2334), .Y(DP_OP_102J5_124_3590_n2302) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1693 ( .A1(n216), .A2(
        DP_OP_102J5_124_3590_n2333), .Y(DP_OP_102J5_124_3590_n2301) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1692 ( .A1(n216), .A2(
        DP_OP_102J5_124_3590_n2332), .Y(DP_OP_102J5_124_3590_n2300) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1691 ( .A1(n216), .A2(
        DP_OP_102J5_124_3590_n2331), .Y(DP_OP_102J5_124_3590_n2299) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1690 ( .A1(n216), .A2(
        DP_OP_102J5_124_3590_n2330), .Y(DP_OP_102J5_124_3590_n2298) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1689 ( .A1(n216), .A2(
        DP_OP_102J5_124_3590_n2329), .Y(DP_OP_102J5_124_3590_n2297) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1676 ( .A1(n271), .A2(
        DP_OP_102J5_124_3590_n2292), .Y(DP_OP_102J5_124_3590_n2284) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1675 ( .A1(n271), .A2(
        DP_OP_102J5_124_3590_n2291), .Y(DP_OP_102J5_124_3590_n2283) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1674 ( .A1(n271), .A2(
        DP_OP_102J5_124_3590_n2290), .Y(DP_OP_102J5_124_3590_n2282) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1673 ( .A1(n271), .A2(
        DP_OP_102J5_124_3590_n2289), .Y(DP_OP_102J5_124_3590_n2281) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1672 ( .A1(n271), .A2(
        DP_OP_102J5_124_3590_n2288), .Y(DP_OP_102J5_124_3590_n2280) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1671 ( .A1(n271), .A2(
        DP_OP_102J5_124_3590_n2287), .Y(DP_OP_102J5_124_3590_n2279) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1670 ( .A1(n271), .A2(
        DP_OP_102J5_124_3590_n2286), .Y(DP_OP_102J5_124_3590_n2278) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1669 ( .A1(n271), .A2(
        DP_OP_102J5_124_3590_n2285), .Y(DP_OP_102J5_124_3590_n2277) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1668 ( .A1(n270), .A2(
        DP_OP_102J5_124_3590_n2292), .Y(DP_OP_102J5_124_3590_n2276) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1667 ( .A1(n270), .A2(
        DP_OP_102J5_124_3590_n2291), .Y(DP_OP_102J5_124_3590_n2275) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1666 ( .A1(n270), .A2(
        DP_OP_102J5_124_3590_n2290), .Y(DP_OP_102J5_124_3590_n2274) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1665 ( .A1(n270), .A2(
        DP_OP_102J5_124_3590_n2289), .Y(DP_OP_102J5_124_3590_n2273) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1664 ( .A1(n270), .A2(
        DP_OP_102J5_124_3590_n2288), .Y(DP_OP_102J5_124_3590_n2272) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1663 ( .A1(n270), .A2(
        DP_OP_102J5_124_3590_n2287), .Y(DP_OP_102J5_124_3590_n2271) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1662 ( .A1(n270), .A2(
        DP_OP_102J5_124_3590_n2286), .Y(DP_OP_102J5_124_3590_n2270) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1661 ( .A1(n270), .A2(
        DP_OP_102J5_124_3590_n2285), .Y(DP_OP_102J5_124_3590_n2269) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1660 ( .A1(n269), .A2(
        DP_OP_102J5_124_3590_n2292), .Y(DP_OP_102J5_124_3590_n2268) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1659 ( .A1(n269), .A2(
        DP_OP_102J5_124_3590_n2291), .Y(DP_OP_102J5_124_3590_n2267) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1658 ( .A1(n269), .A2(
        DP_OP_102J5_124_3590_n2290), .Y(DP_OP_102J5_124_3590_n2266) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1657 ( .A1(n269), .A2(
        DP_OP_102J5_124_3590_n2289), .Y(DP_OP_102J5_124_3590_n2265) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1656 ( .A1(n269), .A2(
        DP_OP_102J5_124_3590_n2288), .Y(DP_OP_102J5_124_3590_n2264) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1655 ( .A1(n269), .A2(
        DP_OP_102J5_124_3590_n2287), .Y(DP_OP_102J5_124_3590_n2263) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1654 ( .A1(n269), .A2(
        DP_OP_102J5_124_3590_n2286), .Y(DP_OP_102J5_124_3590_n2262) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1653 ( .A1(n269), .A2(
        DP_OP_102J5_124_3590_n2285), .Y(DP_OP_102J5_124_3590_n2261) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1652 ( .A1(n215), .A2(
        DP_OP_102J5_124_3590_n2292), .Y(DP_OP_102J5_124_3590_n2260) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1651 ( .A1(n215), .A2(
        DP_OP_102J5_124_3590_n2291), .Y(DP_OP_102J5_124_3590_n2259) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1650 ( .A1(n215), .A2(
        DP_OP_102J5_124_3590_n2290), .Y(DP_OP_102J5_124_3590_n2258) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1649 ( .A1(n215), .A2(
        DP_OP_102J5_124_3590_n2289), .Y(DP_OP_102J5_124_3590_n2257) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1648 ( .A1(n215), .A2(
        DP_OP_102J5_124_3590_n2288), .Y(DP_OP_102J5_124_3590_n2256) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1647 ( .A1(n215), .A2(
        DP_OP_102J5_124_3590_n2287), .Y(DP_OP_102J5_124_3590_n2255) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1646 ( .A1(n215), .A2(
        DP_OP_102J5_124_3590_n2286), .Y(DP_OP_102J5_124_3590_n2254) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1645 ( .A1(n215), .A2(
        DP_OP_102J5_124_3590_n2285), .Y(DP_OP_102J5_124_3590_n2253) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1632 ( .A1(n268), .A2(
        DP_OP_102J5_124_3590_n2248), .Y(DP_OP_102J5_124_3590_n2240) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1631 ( .A1(n268), .A2(
        DP_OP_102J5_124_3590_n2247), .Y(DP_OP_102J5_124_3590_n2239) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1630 ( .A1(n268), .A2(
        DP_OP_102J5_124_3590_n2246), .Y(DP_OP_102J5_124_3590_n2238) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1629 ( .A1(n268), .A2(
        DP_OP_102J5_124_3590_n2245), .Y(DP_OP_102J5_124_3590_n2237) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1628 ( .A1(n268), .A2(
        DP_OP_102J5_124_3590_n2244), .Y(DP_OP_102J5_124_3590_n2236) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1627 ( .A1(n268), .A2(
        DP_OP_102J5_124_3590_n2243), .Y(DP_OP_102J5_124_3590_n2235) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1626 ( .A1(n268), .A2(
        DP_OP_102J5_124_3590_n2242), .Y(DP_OP_102J5_124_3590_n2234) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1625 ( .A1(n268), .A2(
        DP_OP_102J5_124_3590_n2241), .Y(DP_OP_102J5_124_3590_n2233) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1624 ( .A1(n267), .A2(
        DP_OP_102J5_124_3590_n2248), .Y(DP_OP_102J5_124_3590_n2232) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1623 ( .A1(n267), .A2(
        DP_OP_102J5_124_3590_n2247), .Y(DP_OP_102J5_124_3590_n2231) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1622 ( .A1(n267), .A2(
        DP_OP_102J5_124_3590_n2246), .Y(DP_OP_102J5_124_3590_n2230) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1621 ( .A1(n267), .A2(
        DP_OP_102J5_124_3590_n2245), .Y(DP_OP_102J5_124_3590_n2229) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1620 ( .A1(n267), .A2(
        DP_OP_102J5_124_3590_n2244), .Y(DP_OP_102J5_124_3590_n2228) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1619 ( .A1(n267), .A2(
        DP_OP_102J5_124_3590_n2243), .Y(DP_OP_102J5_124_3590_n2227) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1618 ( .A1(n267), .A2(
        DP_OP_102J5_124_3590_n2242), .Y(DP_OP_102J5_124_3590_n2226) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1617 ( .A1(n267), .A2(
        DP_OP_102J5_124_3590_n2241), .Y(DP_OP_102J5_124_3590_n2225) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1616 ( .A1(n266), .A2(
        DP_OP_102J5_124_3590_n2248), .Y(DP_OP_102J5_124_3590_n2224) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1615 ( .A1(n266), .A2(
        DP_OP_102J5_124_3590_n2247), .Y(DP_OP_102J5_124_3590_n2223) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1614 ( .A1(n266), .A2(
        DP_OP_102J5_124_3590_n2246), .Y(DP_OP_102J5_124_3590_n2222) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1613 ( .A1(n266), .A2(
        DP_OP_102J5_124_3590_n2245), .Y(DP_OP_102J5_124_3590_n2221) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1612 ( .A1(n266), .A2(
        DP_OP_102J5_124_3590_n2244), .Y(DP_OP_102J5_124_3590_n2220) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1611 ( .A1(n266), .A2(
        DP_OP_102J5_124_3590_n2243), .Y(DP_OP_102J5_124_3590_n2219) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1610 ( .A1(n266), .A2(
        DP_OP_102J5_124_3590_n2242), .Y(DP_OP_102J5_124_3590_n2218) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1609 ( .A1(n266), .A2(
        DP_OP_102J5_124_3590_n2241), .Y(DP_OP_102J5_124_3590_n2217) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1608 ( .A1(n214), .A2(
        DP_OP_102J5_124_3590_n2248), .Y(DP_OP_102J5_124_3590_n2216) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1607 ( .A1(n214), .A2(
        DP_OP_102J5_124_3590_n2247), .Y(DP_OP_102J5_124_3590_n2215) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1606 ( .A1(n214), .A2(
        DP_OP_102J5_124_3590_n2246), .Y(DP_OP_102J5_124_3590_n2214) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1605 ( .A1(n214), .A2(
        DP_OP_102J5_124_3590_n2245), .Y(DP_OP_102J5_124_3590_n2213) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1604 ( .A1(n214), .A2(
        DP_OP_102J5_124_3590_n2244), .Y(DP_OP_102J5_124_3590_n2212) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1603 ( .A1(n214), .A2(
        DP_OP_102J5_124_3590_n2243), .Y(DP_OP_102J5_124_3590_n2211) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1602 ( .A1(n214), .A2(
        DP_OP_102J5_124_3590_n2242), .Y(DP_OP_102J5_124_3590_n2210) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1601 ( .A1(n214), .A2(
        DP_OP_102J5_124_3590_n2241), .Y(DP_OP_102J5_124_3590_n2209) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1588 ( .A1(n265), .A2(
        DP_OP_102J5_124_3590_n2204), .Y(DP_OP_102J5_124_3590_n2196) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1587 ( .A1(n265), .A2(
        DP_OP_102J5_124_3590_n2203), .Y(DP_OP_102J5_124_3590_n2195) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1586 ( .A1(n265), .A2(
        DP_OP_102J5_124_3590_n2202), .Y(DP_OP_102J5_124_3590_n2194) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1585 ( .A1(n265), .A2(
        DP_OP_102J5_124_3590_n2201), .Y(DP_OP_102J5_124_3590_n2193) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1584 ( .A1(n265), .A2(
        DP_OP_102J5_124_3590_n2200), .Y(DP_OP_102J5_124_3590_n2192) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1583 ( .A1(n265), .A2(
        DP_OP_102J5_124_3590_n2199), .Y(DP_OP_102J5_124_3590_n2191) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1582 ( .A1(n265), .A2(
        DP_OP_102J5_124_3590_n2198), .Y(DP_OP_102J5_124_3590_n2190) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1581 ( .A1(n265), .A2(
        DP_OP_102J5_124_3590_n2197), .Y(DP_OP_102J5_124_3590_n2189) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1580 ( .A1(n264), .A2(
        DP_OP_102J5_124_3590_n2204), .Y(DP_OP_102J5_124_3590_n2188) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1579 ( .A1(n264), .A2(
        DP_OP_102J5_124_3590_n2203), .Y(DP_OP_102J5_124_3590_n2187) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1578 ( .A1(n264), .A2(
        DP_OP_102J5_124_3590_n2202), .Y(DP_OP_102J5_124_3590_n2186) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1577 ( .A1(n264), .A2(
        DP_OP_102J5_124_3590_n2201), .Y(DP_OP_102J5_124_3590_n2185) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1576 ( .A1(n264), .A2(
        DP_OP_102J5_124_3590_n2200), .Y(DP_OP_102J5_124_3590_n2184) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1575 ( .A1(n264), .A2(
        DP_OP_102J5_124_3590_n2199), .Y(DP_OP_102J5_124_3590_n2183) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1574 ( .A1(n264), .A2(
        DP_OP_102J5_124_3590_n2198), .Y(DP_OP_102J5_124_3590_n2182) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1573 ( .A1(n264), .A2(
        DP_OP_102J5_124_3590_n2197), .Y(DP_OP_102J5_124_3590_n2181) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1572 ( .A1(n263), .A2(
        DP_OP_102J5_124_3590_n2204), .Y(DP_OP_102J5_124_3590_n2180) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1571 ( .A1(n263), .A2(
        DP_OP_102J5_124_3590_n2203), .Y(DP_OP_102J5_124_3590_n2179) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1570 ( .A1(n263), .A2(
        DP_OP_102J5_124_3590_n2202), .Y(DP_OP_102J5_124_3590_n2178) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1569 ( .A1(n263), .A2(
        DP_OP_102J5_124_3590_n2201), .Y(DP_OP_102J5_124_3590_n2177) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1568 ( .A1(n263), .A2(
        DP_OP_102J5_124_3590_n2200), .Y(DP_OP_102J5_124_3590_n2176) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1567 ( .A1(n263), .A2(
        DP_OP_102J5_124_3590_n2199), .Y(DP_OP_102J5_124_3590_n2175) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1566 ( .A1(n263), .A2(
        DP_OP_102J5_124_3590_n2198), .Y(DP_OP_102J5_124_3590_n2174) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1565 ( .A1(n263), .A2(
        DP_OP_102J5_124_3590_n2197), .Y(DP_OP_102J5_124_3590_n2173) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1564 ( .A1(n213), .A2(
        DP_OP_102J5_124_3590_n2204), .Y(DP_OP_102J5_124_3590_n2172) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1563 ( .A1(n213), .A2(
        DP_OP_102J5_124_3590_n2203), .Y(DP_OP_102J5_124_3590_n2171) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1562 ( .A1(n213), .A2(
        DP_OP_102J5_124_3590_n2202), .Y(DP_OP_102J5_124_3590_n2170) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1561 ( .A1(n213), .A2(
        DP_OP_102J5_124_3590_n2201), .Y(DP_OP_102J5_124_3590_n2169) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1560 ( .A1(n213), .A2(
        DP_OP_102J5_124_3590_n2200), .Y(DP_OP_102J5_124_3590_n2168) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1559 ( .A1(n213), .A2(
        DP_OP_102J5_124_3590_n2199), .Y(DP_OP_102J5_124_3590_n2167) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1558 ( .A1(n213), .A2(
        DP_OP_102J5_124_3590_n2198), .Y(DP_OP_102J5_124_3590_n2166) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1557 ( .A1(n213), .A2(
        DP_OP_102J5_124_3590_n2197), .Y(DP_OP_102J5_124_3590_n2165) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1544 ( .A1(n262), .A2(
        DP_OP_102J5_124_3590_n2160), .Y(DP_OP_102J5_124_3590_n2152) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1543 ( .A1(n262), .A2(
        DP_OP_102J5_124_3590_n2159), .Y(DP_OP_102J5_124_3590_n2151) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1542 ( .A1(n262), .A2(
        DP_OP_102J5_124_3590_n2158), .Y(DP_OP_102J5_124_3590_n2150) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1541 ( .A1(n262), .A2(
        DP_OP_102J5_124_3590_n2157), .Y(DP_OP_102J5_124_3590_n2149) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1540 ( .A1(n262), .A2(
        DP_OP_102J5_124_3590_n2156), .Y(DP_OP_102J5_124_3590_n2148) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1539 ( .A1(n262), .A2(
        DP_OP_102J5_124_3590_n2155), .Y(DP_OP_102J5_124_3590_n2147) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1538 ( .A1(n262), .A2(
        DP_OP_102J5_124_3590_n2154), .Y(DP_OP_102J5_124_3590_n2146) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1537 ( .A1(n262), .A2(
        DP_OP_102J5_124_3590_n2153), .Y(DP_OP_102J5_124_3590_n2145) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1536 ( .A1(n261), .A2(
        DP_OP_102J5_124_3590_n2160), .Y(DP_OP_102J5_124_3590_n2144) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1535 ( .A1(n261), .A2(
        DP_OP_102J5_124_3590_n2159), .Y(DP_OP_102J5_124_3590_n2143) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1534 ( .A1(n261), .A2(
        DP_OP_102J5_124_3590_n2158), .Y(DP_OP_102J5_124_3590_n2142) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1533 ( .A1(n261), .A2(
        DP_OP_102J5_124_3590_n2157), .Y(DP_OP_102J5_124_3590_n2141) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1532 ( .A1(n261), .A2(
        DP_OP_102J5_124_3590_n2156), .Y(DP_OP_102J5_124_3590_n2140) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1531 ( .A1(n261), .A2(
        DP_OP_102J5_124_3590_n2155), .Y(DP_OP_102J5_124_3590_n2139) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1530 ( .A1(n261), .A2(
        DP_OP_102J5_124_3590_n2154), .Y(DP_OP_102J5_124_3590_n2138) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1529 ( .A1(n261), .A2(
        DP_OP_102J5_124_3590_n2153), .Y(DP_OP_102J5_124_3590_n2137) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1528 ( .A1(n260), .A2(
        DP_OP_102J5_124_3590_n2160), .Y(DP_OP_102J5_124_3590_n2136) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1527 ( .A1(n260), .A2(
        DP_OP_102J5_124_3590_n2159), .Y(DP_OP_102J5_124_3590_n2135) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1526 ( .A1(n260), .A2(
        DP_OP_102J5_124_3590_n2158), .Y(DP_OP_102J5_124_3590_n2134) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1525 ( .A1(n260), .A2(
        DP_OP_102J5_124_3590_n2157), .Y(DP_OP_102J5_124_3590_n2133) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1524 ( .A1(n260), .A2(
        DP_OP_102J5_124_3590_n2156), .Y(DP_OP_102J5_124_3590_n2132) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1523 ( .A1(n260), .A2(
        DP_OP_102J5_124_3590_n2155), .Y(DP_OP_102J5_124_3590_n2131) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1522 ( .A1(n260), .A2(
        DP_OP_102J5_124_3590_n2154), .Y(DP_OP_102J5_124_3590_n2130) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1521 ( .A1(n260), .A2(
        DP_OP_102J5_124_3590_n2153), .Y(DP_OP_102J5_124_3590_n2129) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1520 ( .A1(n212), .A2(
        DP_OP_102J5_124_3590_n2160), .Y(DP_OP_102J5_124_3590_n2128) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1519 ( .A1(n212), .A2(
        DP_OP_102J5_124_3590_n2159), .Y(DP_OP_102J5_124_3590_n2127) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1518 ( .A1(n212), .A2(
        DP_OP_102J5_124_3590_n2158), .Y(DP_OP_102J5_124_3590_n2126) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1517 ( .A1(n212), .A2(
        DP_OP_102J5_124_3590_n2157), .Y(DP_OP_102J5_124_3590_n2125) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1516 ( .A1(n212), .A2(
        DP_OP_102J5_124_3590_n2156), .Y(DP_OP_102J5_124_3590_n2124) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1515 ( .A1(n212), .A2(
        DP_OP_102J5_124_3590_n2155), .Y(DP_OP_102J5_124_3590_n2123) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1514 ( .A1(n212), .A2(
        DP_OP_102J5_124_3590_n2154), .Y(DP_OP_102J5_124_3590_n2122) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1513 ( .A1(n212), .A2(
        DP_OP_102J5_124_3590_n2153), .Y(DP_OP_102J5_124_3590_n2121) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1500 ( .A1(n259), .A2(
        DP_OP_102J5_124_3590_n2116), .Y(DP_OP_102J5_124_3590_n2108) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1499 ( .A1(n259), .A2(
        DP_OP_102J5_124_3590_n2115), .Y(DP_OP_102J5_124_3590_n2107) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1498 ( .A1(n259), .A2(
        DP_OP_102J5_124_3590_n2114), .Y(DP_OP_102J5_124_3590_n2106) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1497 ( .A1(n259), .A2(
        DP_OP_102J5_124_3590_n2113), .Y(DP_OP_102J5_124_3590_n2105) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1496 ( .A1(n259), .A2(
        DP_OP_102J5_124_3590_n2112), .Y(DP_OP_102J5_124_3590_n2104) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1495 ( .A1(n259), .A2(
        DP_OP_102J5_124_3590_n2111), .Y(DP_OP_102J5_124_3590_n2103) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1494 ( .A1(n259), .A2(
        DP_OP_102J5_124_3590_n2110), .Y(DP_OP_102J5_124_3590_n2102) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1493 ( .A1(n259), .A2(
        DP_OP_102J5_124_3590_n2109), .Y(DP_OP_102J5_124_3590_n2101) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1492 ( .A1(n258), .A2(
        DP_OP_102J5_124_3590_n2116), .Y(DP_OP_102J5_124_3590_n2100) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1491 ( .A1(n258), .A2(
        DP_OP_102J5_124_3590_n2115), .Y(DP_OP_102J5_124_3590_n2099) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1490 ( .A1(n258), .A2(
        DP_OP_102J5_124_3590_n2114), .Y(DP_OP_102J5_124_3590_n2098) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1489 ( .A1(n258), .A2(
        DP_OP_102J5_124_3590_n2113), .Y(DP_OP_102J5_124_3590_n2097) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1488 ( .A1(n258), .A2(
        DP_OP_102J5_124_3590_n2112), .Y(DP_OP_102J5_124_3590_n2096) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1487 ( .A1(n258), .A2(
        DP_OP_102J5_124_3590_n2111), .Y(DP_OP_102J5_124_3590_n2095) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1486 ( .A1(n258), .A2(
        DP_OP_102J5_124_3590_n2110), .Y(DP_OP_102J5_124_3590_n2094) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1485 ( .A1(n258), .A2(
        DP_OP_102J5_124_3590_n2109), .Y(DP_OP_102J5_124_3590_n2093) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1484 ( .A1(n257), .A2(
        DP_OP_102J5_124_3590_n2116), .Y(DP_OP_102J5_124_3590_n2092) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1483 ( .A1(n257), .A2(
        DP_OP_102J5_124_3590_n2115), .Y(DP_OP_102J5_124_3590_n2091) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1482 ( .A1(n257), .A2(
        DP_OP_102J5_124_3590_n2114), .Y(DP_OP_102J5_124_3590_n2090) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1481 ( .A1(n257), .A2(
        DP_OP_102J5_124_3590_n2113), .Y(DP_OP_102J5_124_3590_n2089) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1480 ( .A1(n257), .A2(
        DP_OP_102J5_124_3590_n2112), .Y(DP_OP_102J5_124_3590_n2088) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1479 ( .A1(n257), .A2(
        DP_OP_102J5_124_3590_n2111), .Y(DP_OP_102J5_124_3590_n2087) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1478 ( .A1(n257), .A2(
        DP_OP_102J5_124_3590_n2110), .Y(DP_OP_102J5_124_3590_n2086) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1477 ( .A1(n257), .A2(
        DP_OP_102J5_124_3590_n2109), .Y(DP_OP_102J5_124_3590_n2085) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1476 ( .A1(n211), .A2(
        DP_OP_102J5_124_3590_n2116), .Y(DP_OP_102J5_124_3590_n2084) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1475 ( .A1(n211), .A2(
        DP_OP_102J5_124_3590_n2115), .Y(DP_OP_102J5_124_3590_n2083) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1474 ( .A1(n211), .A2(
        DP_OP_102J5_124_3590_n2114), .Y(DP_OP_102J5_124_3590_n2082) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1473 ( .A1(n211), .A2(
        DP_OP_102J5_124_3590_n2113), .Y(DP_OP_102J5_124_3590_n2081) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1472 ( .A1(n211), .A2(
        DP_OP_102J5_124_3590_n2112), .Y(DP_OP_102J5_124_3590_n2080) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1471 ( .A1(n211), .A2(
        DP_OP_102J5_124_3590_n2111), .Y(DP_OP_102J5_124_3590_n2079) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1470 ( .A1(n211), .A2(
        DP_OP_102J5_124_3590_n2110), .Y(DP_OP_102J5_124_3590_n2078) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1469 ( .A1(n211), .A2(
        DP_OP_102J5_124_3590_n2109), .Y(DP_OP_102J5_124_3590_n2077) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1456 ( .A1(n256), .A2(
        DP_OP_102J5_124_3590_n2072), .Y(DP_OP_102J5_124_3590_n2064) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1455 ( .A1(n256), .A2(
        DP_OP_102J5_124_3590_n2071), .Y(DP_OP_102J5_124_3590_n2063) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1454 ( .A1(n256), .A2(
        DP_OP_102J5_124_3590_n2070), .Y(DP_OP_102J5_124_3590_n2062) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1453 ( .A1(n256), .A2(
        DP_OP_102J5_124_3590_n2069), .Y(DP_OP_102J5_124_3590_n2061) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1452 ( .A1(n256), .A2(
        DP_OP_102J5_124_3590_n2068), .Y(DP_OP_102J5_124_3590_n2060) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1451 ( .A1(n256), .A2(
        DP_OP_102J5_124_3590_n2067), .Y(DP_OP_102J5_124_3590_n2059) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1450 ( .A1(n256), .A2(
        DP_OP_102J5_124_3590_n2066), .Y(DP_OP_102J5_124_3590_n2058) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1449 ( .A1(n256), .A2(
        DP_OP_102J5_124_3590_n2065), .Y(DP_OP_102J5_124_3590_n2057) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1448 ( .A1(n255), .A2(
        DP_OP_102J5_124_3590_n2072), .Y(DP_OP_102J5_124_3590_n2056) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1447 ( .A1(n255), .A2(
        DP_OP_102J5_124_3590_n2071), .Y(DP_OP_102J5_124_3590_n2055) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1446 ( .A1(n255), .A2(
        DP_OP_102J5_124_3590_n2070), .Y(DP_OP_102J5_124_3590_n2054) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1445 ( .A1(n255), .A2(
        DP_OP_102J5_124_3590_n2069), .Y(DP_OP_102J5_124_3590_n2053) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1444 ( .A1(n255), .A2(
        DP_OP_102J5_124_3590_n2068), .Y(DP_OP_102J5_124_3590_n2052) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1443 ( .A1(n255), .A2(
        DP_OP_102J5_124_3590_n2067), .Y(DP_OP_102J5_124_3590_n2051) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1442 ( .A1(n255), .A2(
        DP_OP_102J5_124_3590_n2066), .Y(DP_OP_102J5_124_3590_n2050) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1441 ( .A1(n255), .A2(
        DP_OP_102J5_124_3590_n2065), .Y(DP_OP_102J5_124_3590_n2049) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1440 ( .A1(n254), .A2(
        DP_OP_102J5_124_3590_n2072), .Y(DP_OP_102J5_124_3590_n2048) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1439 ( .A1(n254), .A2(
        DP_OP_102J5_124_3590_n2071), .Y(DP_OP_102J5_124_3590_n2047) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1438 ( .A1(n254), .A2(
        DP_OP_102J5_124_3590_n2070), .Y(DP_OP_102J5_124_3590_n2046) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1437 ( .A1(n254), .A2(
        DP_OP_102J5_124_3590_n2069), .Y(DP_OP_102J5_124_3590_n2045) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1436 ( .A1(n254), .A2(
        DP_OP_102J5_124_3590_n2068), .Y(DP_OP_102J5_124_3590_n2044) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1435 ( .A1(n254), .A2(
        DP_OP_102J5_124_3590_n2067), .Y(DP_OP_102J5_124_3590_n2043) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1434 ( .A1(n254), .A2(
        DP_OP_102J5_124_3590_n2066), .Y(DP_OP_102J5_124_3590_n2042) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1433 ( .A1(n254), .A2(
        DP_OP_102J5_124_3590_n2065), .Y(DP_OP_102J5_124_3590_n2041) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1432 ( .A1(n210), .A2(
        DP_OP_102J5_124_3590_n2072), .Y(DP_OP_102J5_124_3590_n2040) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1431 ( .A1(n210), .A2(
        DP_OP_102J5_124_3590_n2071), .Y(DP_OP_102J5_124_3590_n2039) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1430 ( .A1(n210), .A2(
        DP_OP_102J5_124_3590_n2070), .Y(DP_OP_102J5_124_3590_n2038) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1429 ( .A1(n210), .A2(
        DP_OP_102J5_124_3590_n2069), .Y(DP_OP_102J5_124_3590_n2037) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1428 ( .A1(n210), .A2(
        DP_OP_102J5_124_3590_n2068), .Y(DP_OP_102J5_124_3590_n2036) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1427 ( .A1(n210), .A2(
        DP_OP_102J5_124_3590_n2067), .Y(DP_OP_102J5_124_3590_n2035) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1426 ( .A1(n210), .A2(
        DP_OP_102J5_124_3590_n2066), .Y(DP_OP_102J5_124_3590_n2034) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1425 ( .A1(n210), .A2(
        DP_OP_102J5_124_3590_n2065), .Y(DP_OP_102J5_124_3590_n2033) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1412 ( .A1(n253), .A2(
        DP_OP_102J5_124_3590_n2028), .Y(DP_OP_102J5_124_3590_n2020) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1411 ( .A1(n253), .A2(
        DP_OP_102J5_124_3590_n2027), .Y(DP_OP_102J5_124_3590_n2019) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1410 ( .A1(n253), .A2(
        DP_OP_102J5_124_3590_n2026), .Y(DP_OP_102J5_124_3590_n2018) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1409 ( .A1(n253), .A2(
        DP_OP_102J5_124_3590_n2025), .Y(DP_OP_102J5_124_3590_n2017) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1408 ( .A1(n253), .A2(
        DP_OP_102J5_124_3590_n2024), .Y(DP_OP_102J5_124_3590_n2016) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1407 ( .A1(n253), .A2(
        DP_OP_102J5_124_3590_n2023), .Y(DP_OP_102J5_124_3590_n2015) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1406 ( .A1(n253), .A2(
        DP_OP_102J5_124_3590_n2022), .Y(DP_OP_102J5_124_3590_n2014) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1405 ( .A1(n253), .A2(
        DP_OP_102J5_124_3590_n2021), .Y(DP_OP_102J5_124_3590_n2013) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1404 ( .A1(n252), .A2(
        DP_OP_102J5_124_3590_n2028), .Y(DP_OP_102J5_124_3590_n2012) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1403 ( .A1(n252), .A2(
        DP_OP_102J5_124_3590_n2027), .Y(DP_OP_102J5_124_3590_n2011) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1402 ( .A1(n252), .A2(
        DP_OP_102J5_124_3590_n2026), .Y(DP_OP_102J5_124_3590_n2010) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1401 ( .A1(n252), .A2(
        DP_OP_102J5_124_3590_n2025), .Y(DP_OP_102J5_124_3590_n2009) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1400 ( .A1(n252), .A2(
        DP_OP_102J5_124_3590_n2024), .Y(DP_OP_102J5_124_3590_n2008) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1399 ( .A1(n252), .A2(
        DP_OP_102J5_124_3590_n2023), .Y(DP_OP_102J5_124_3590_n2007) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1398 ( .A1(n252), .A2(
        DP_OP_102J5_124_3590_n2022), .Y(DP_OP_102J5_124_3590_n2006) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1397 ( .A1(n252), .A2(
        DP_OP_102J5_124_3590_n2021), .Y(DP_OP_102J5_124_3590_n2005) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1396 ( .A1(n251), .A2(
        DP_OP_102J5_124_3590_n2028), .Y(DP_OP_102J5_124_3590_n2004) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1395 ( .A1(n251), .A2(
        DP_OP_102J5_124_3590_n2027), .Y(DP_OP_102J5_124_3590_n2003) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1394 ( .A1(n251), .A2(
        DP_OP_102J5_124_3590_n2026), .Y(DP_OP_102J5_124_3590_n2002) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1393 ( .A1(n251), .A2(
        DP_OP_102J5_124_3590_n2025), .Y(DP_OP_102J5_124_3590_n2001) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1392 ( .A1(n251), .A2(
        DP_OP_102J5_124_3590_n2024), .Y(DP_OP_102J5_124_3590_n2000) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1391 ( .A1(n251), .A2(
        DP_OP_102J5_124_3590_n2023), .Y(DP_OP_102J5_124_3590_n1999) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1390 ( .A1(n251), .A2(
        DP_OP_102J5_124_3590_n2022), .Y(DP_OP_102J5_124_3590_n1998) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1389 ( .A1(n251), .A2(
        DP_OP_102J5_124_3590_n2021), .Y(DP_OP_102J5_124_3590_n1997) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1388 ( .A1(n209), .A2(
        DP_OP_102J5_124_3590_n2028), .Y(DP_OP_102J5_124_3590_n1996) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1387 ( .A1(n209), .A2(
        DP_OP_102J5_124_3590_n2027), .Y(DP_OP_102J5_124_3590_n1995) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1386 ( .A1(n209), .A2(
        DP_OP_102J5_124_3590_n2026), .Y(DP_OP_102J5_124_3590_n1994) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1385 ( .A1(n209), .A2(
        DP_OP_102J5_124_3590_n2025), .Y(DP_OP_102J5_124_3590_n1993) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1384 ( .A1(n209), .A2(
        DP_OP_102J5_124_3590_n2024), .Y(DP_OP_102J5_124_3590_n1992) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1383 ( .A1(n209), .A2(
        DP_OP_102J5_124_3590_n2023), .Y(DP_OP_102J5_124_3590_n1991) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1382 ( .A1(n209), .A2(
        DP_OP_102J5_124_3590_n2022), .Y(DP_OP_102J5_124_3590_n1990) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1381 ( .A1(n209), .A2(
        DP_OP_102J5_124_3590_n2021), .Y(DP_OP_102J5_124_3590_n1989) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1368 ( .A1(n250), .A2(
        DP_OP_102J5_124_3590_n1984), .Y(DP_OP_102J5_124_3590_n1976) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1367 ( .A1(n250), .A2(
        DP_OP_102J5_124_3590_n1983), .Y(DP_OP_102J5_124_3590_n1975) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1366 ( .A1(n250), .A2(
        DP_OP_102J5_124_3590_n1982), .Y(DP_OP_102J5_124_3590_n1974) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1365 ( .A1(n250), .A2(
        DP_OP_102J5_124_3590_n1981), .Y(DP_OP_102J5_124_3590_n1973) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1364 ( .A1(n250), .A2(
        DP_OP_102J5_124_3590_n1980), .Y(DP_OP_102J5_124_3590_n1972) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1363 ( .A1(n250), .A2(
        DP_OP_102J5_124_3590_n1979), .Y(DP_OP_102J5_124_3590_n1971) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1362 ( .A1(n250), .A2(
        DP_OP_102J5_124_3590_n1978), .Y(DP_OP_102J5_124_3590_n1970) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1361 ( .A1(n250), .A2(
        DP_OP_102J5_124_3590_n1977), .Y(DP_OP_102J5_124_3590_n1969) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1360 ( .A1(n249), .A2(
        DP_OP_102J5_124_3590_n1984), .Y(DP_OP_102J5_124_3590_n1968) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1359 ( .A1(n249), .A2(
        DP_OP_102J5_124_3590_n1983), .Y(DP_OP_102J5_124_3590_n1967) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1358 ( .A1(n249), .A2(
        DP_OP_102J5_124_3590_n1982), .Y(DP_OP_102J5_124_3590_n1966) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1357 ( .A1(n249), .A2(
        DP_OP_102J5_124_3590_n1981), .Y(DP_OP_102J5_124_3590_n1965) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1356 ( .A1(n249), .A2(
        DP_OP_102J5_124_3590_n1980), .Y(DP_OP_102J5_124_3590_n1964) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1355 ( .A1(n249), .A2(
        DP_OP_102J5_124_3590_n1979), .Y(DP_OP_102J5_124_3590_n1963) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1354 ( .A1(n249), .A2(
        DP_OP_102J5_124_3590_n1978), .Y(DP_OP_102J5_124_3590_n1962) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1353 ( .A1(n249), .A2(
        DP_OP_102J5_124_3590_n1977), .Y(DP_OP_102J5_124_3590_n1961) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1352 ( .A1(n248), .A2(
        DP_OP_102J5_124_3590_n1984), .Y(DP_OP_102J5_124_3590_n1960) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1351 ( .A1(n248), .A2(
        DP_OP_102J5_124_3590_n1983), .Y(DP_OP_102J5_124_3590_n1959) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1350 ( .A1(n248), .A2(
        DP_OP_102J5_124_3590_n1982), .Y(DP_OP_102J5_124_3590_n1958) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1349 ( .A1(n248), .A2(
        DP_OP_102J5_124_3590_n1981), .Y(DP_OP_102J5_124_3590_n1957) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1348 ( .A1(n248), .A2(
        DP_OP_102J5_124_3590_n1980), .Y(DP_OP_102J5_124_3590_n1956) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1347 ( .A1(n248), .A2(
        DP_OP_102J5_124_3590_n1979), .Y(DP_OP_102J5_124_3590_n1955) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1346 ( .A1(n248), .A2(
        DP_OP_102J5_124_3590_n1978), .Y(DP_OP_102J5_124_3590_n1954) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1345 ( .A1(n248), .A2(
        DP_OP_102J5_124_3590_n1977), .Y(DP_OP_102J5_124_3590_n1953) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1344 ( .A1(n208), .A2(
        DP_OP_102J5_124_3590_n1984), .Y(DP_OP_102J5_124_3590_n1952) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1343 ( .A1(n208), .A2(
        DP_OP_102J5_124_3590_n1983), .Y(DP_OP_102J5_124_3590_n1951) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1342 ( .A1(n208), .A2(
        DP_OP_102J5_124_3590_n1982), .Y(DP_OP_102J5_124_3590_n1950) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1341 ( .A1(n208), .A2(
        DP_OP_102J5_124_3590_n1981), .Y(DP_OP_102J5_124_3590_n1949) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1340 ( .A1(n208), .A2(
        DP_OP_102J5_124_3590_n1980), .Y(DP_OP_102J5_124_3590_n1948) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1339 ( .A1(n208), .A2(
        DP_OP_102J5_124_3590_n1979), .Y(DP_OP_102J5_124_3590_n1947) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1338 ( .A1(n208), .A2(
        DP_OP_102J5_124_3590_n1978), .Y(DP_OP_102J5_124_3590_n1946) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1337 ( .A1(n208), .A2(
        DP_OP_102J5_124_3590_n1977), .Y(DP_OP_102J5_124_3590_n1945) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1324 ( .A1(n247), .A2(
        DP_OP_102J5_124_3590_n1940), .Y(DP_OP_102J5_124_3590_n1932) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1323 ( .A1(n247), .A2(
        DP_OP_102J5_124_3590_n1939), .Y(DP_OP_102J5_124_3590_n1931) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1322 ( .A1(n247), .A2(
        DP_OP_102J5_124_3590_n1938), .Y(DP_OP_102J5_124_3590_n1930) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1321 ( .A1(n247), .A2(
        DP_OP_102J5_124_3590_n1937), .Y(DP_OP_102J5_124_3590_n1929) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1320 ( .A1(n247), .A2(
        DP_OP_102J5_124_3590_n1936), .Y(DP_OP_102J5_124_3590_n1928) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1319 ( .A1(n247), .A2(
        DP_OP_102J5_124_3590_n1935), .Y(DP_OP_102J5_124_3590_n1927) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1318 ( .A1(n247), .A2(
        DP_OP_102J5_124_3590_n1934), .Y(DP_OP_102J5_124_3590_n1926) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1317 ( .A1(n247), .A2(
        DP_OP_102J5_124_3590_n1933), .Y(DP_OP_102J5_124_3590_n1925) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1316 ( .A1(n246), .A2(
        DP_OP_102J5_124_3590_n1940), .Y(DP_OP_102J5_124_3590_n1924) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1315 ( .A1(n246), .A2(
        DP_OP_102J5_124_3590_n1939), .Y(DP_OP_102J5_124_3590_n1923) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1314 ( .A1(n246), .A2(
        DP_OP_102J5_124_3590_n1938), .Y(DP_OP_102J5_124_3590_n1922) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1313 ( .A1(n246), .A2(
        DP_OP_102J5_124_3590_n1937), .Y(DP_OP_102J5_124_3590_n1921) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1312 ( .A1(n246), .A2(
        DP_OP_102J5_124_3590_n1936), .Y(DP_OP_102J5_124_3590_n1920) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1311 ( .A1(n246), .A2(
        DP_OP_102J5_124_3590_n1935), .Y(DP_OP_102J5_124_3590_n1919) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1310 ( .A1(n246), .A2(
        DP_OP_102J5_124_3590_n1934), .Y(DP_OP_102J5_124_3590_n1918) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1309 ( .A1(n246), .A2(
        DP_OP_102J5_124_3590_n1933), .Y(DP_OP_102J5_124_3590_n1917) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1308 ( .A1(n245), .A2(
        DP_OP_102J5_124_3590_n1940), .Y(DP_OP_102J5_124_3590_n1916) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1307 ( .A1(n245), .A2(
        DP_OP_102J5_124_3590_n1939), .Y(DP_OP_102J5_124_3590_n1915) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1306 ( .A1(n245), .A2(
        DP_OP_102J5_124_3590_n1938), .Y(DP_OP_102J5_124_3590_n1914) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1305 ( .A1(n245), .A2(
        DP_OP_102J5_124_3590_n1937), .Y(DP_OP_102J5_124_3590_n1913) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1304 ( .A1(n245), .A2(
        DP_OP_102J5_124_3590_n1936), .Y(DP_OP_102J5_124_3590_n1912) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1303 ( .A1(n245), .A2(
        DP_OP_102J5_124_3590_n1935), .Y(DP_OP_102J5_124_3590_n1911) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1302 ( .A1(n245), .A2(
        DP_OP_102J5_124_3590_n1934), .Y(DP_OP_102J5_124_3590_n1910) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1301 ( .A1(n245), .A2(
        DP_OP_102J5_124_3590_n1933), .Y(DP_OP_102J5_124_3590_n1909) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1300 ( .A1(n207), .A2(
        DP_OP_102J5_124_3590_n1940), .Y(DP_OP_102J5_124_3590_n1908) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1299 ( .A1(n207), .A2(
        DP_OP_102J5_124_3590_n1939), .Y(DP_OP_102J5_124_3590_n1907) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1298 ( .A1(n207), .A2(
        DP_OP_102J5_124_3590_n1938), .Y(DP_OP_102J5_124_3590_n1906) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1297 ( .A1(n207), .A2(
        DP_OP_102J5_124_3590_n1937), .Y(DP_OP_102J5_124_3590_n1905) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1296 ( .A1(n207), .A2(
        DP_OP_102J5_124_3590_n1936), .Y(DP_OP_102J5_124_3590_n1904) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1295 ( .A1(n207), .A2(
        DP_OP_102J5_124_3590_n1935), .Y(DP_OP_102J5_124_3590_n1903) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1294 ( .A1(n207), .A2(
        DP_OP_102J5_124_3590_n1934), .Y(DP_OP_102J5_124_3590_n1902) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1293 ( .A1(n207), .A2(
        DP_OP_102J5_124_3590_n1933), .Y(DP_OP_102J5_124_3590_n1901) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1280 ( .A1(n244), .A2(
        DP_OP_102J5_124_3590_n1896), .Y(DP_OP_102J5_124_3590_n1888) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1279 ( .A1(n244), .A2(
        DP_OP_102J5_124_3590_n1895), .Y(DP_OP_102J5_124_3590_n1887) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1278 ( .A1(n244), .A2(
        DP_OP_102J5_124_3590_n1894), .Y(DP_OP_102J5_124_3590_n1886) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1277 ( .A1(n244), .A2(
        DP_OP_102J5_124_3590_n1893), .Y(DP_OP_102J5_124_3590_n1885) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1276 ( .A1(n244), .A2(
        DP_OP_102J5_124_3590_n1892), .Y(DP_OP_102J5_124_3590_n1884) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1275 ( .A1(n244), .A2(
        DP_OP_102J5_124_3590_n1891), .Y(DP_OP_102J5_124_3590_n1883) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1274 ( .A1(n244), .A2(
        DP_OP_102J5_124_3590_n1890), .Y(DP_OP_102J5_124_3590_n1882) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1273 ( .A1(n244), .A2(
        DP_OP_102J5_124_3590_n1889), .Y(DP_OP_102J5_124_3590_n1881) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1272 ( .A1(n243), .A2(
        DP_OP_102J5_124_3590_n1896), .Y(DP_OP_102J5_124_3590_n1880) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1271 ( .A1(n243), .A2(
        DP_OP_102J5_124_3590_n1895), .Y(DP_OP_102J5_124_3590_n1879) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1270 ( .A1(n243), .A2(
        DP_OP_102J5_124_3590_n1894), .Y(DP_OP_102J5_124_3590_n1878) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1269 ( .A1(n243), .A2(
        DP_OP_102J5_124_3590_n1893), .Y(DP_OP_102J5_124_3590_n1877) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1268 ( .A1(n243), .A2(
        DP_OP_102J5_124_3590_n1892), .Y(DP_OP_102J5_124_3590_n1876) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1267 ( .A1(n243), .A2(
        DP_OP_102J5_124_3590_n1891), .Y(DP_OP_102J5_124_3590_n1875) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1266 ( .A1(n243), .A2(
        DP_OP_102J5_124_3590_n1890), .Y(DP_OP_102J5_124_3590_n1874) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1265 ( .A1(n243), .A2(
        DP_OP_102J5_124_3590_n1889), .Y(DP_OP_102J5_124_3590_n1873) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1264 ( .A1(n242), .A2(
        DP_OP_102J5_124_3590_n1896), .Y(DP_OP_102J5_124_3590_n1872) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1263 ( .A1(n242), .A2(
        DP_OP_102J5_124_3590_n1895), .Y(DP_OP_102J5_124_3590_n1871) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1262 ( .A1(n242), .A2(
        DP_OP_102J5_124_3590_n1894), .Y(DP_OP_102J5_124_3590_n1870) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1261 ( .A1(n242), .A2(
        DP_OP_102J5_124_3590_n1893), .Y(DP_OP_102J5_124_3590_n1869) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1260 ( .A1(n242), .A2(
        DP_OP_102J5_124_3590_n1892), .Y(DP_OP_102J5_124_3590_n1868) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1259 ( .A1(n242), .A2(
        DP_OP_102J5_124_3590_n1891), .Y(DP_OP_102J5_124_3590_n1867) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1258 ( .A1(n242), .A2(
        DP_OP_102J5_124_3590_n1890), .Y(DP_OP_102J5_124_3590_n1866) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1257 ( .A1(n242), .A2(
        DP_OP_102J5_124_3590_n1889), .Y(DP_OP_102J5_124_3590_n1865) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1256 ( .A1(n206), .A2(
        DP_OP_102J5_124_3590_n1896), .Y(DP_OP_102J5_124_3590_n1864) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1255 ( .A1(n206), .A2(
        DP_OP_102J5_124_3590_n1895), .Y(DP_OP_102J5_124_3590_n1863) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1254 ( .A1(n206), .A2(
        DP_OP_102J5_124_3590_n1894), .Y(DP_OP_102J5_124_3590_n1862) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1253 ( .A1(n206), .A2(
        DP_OP_102J5_124_3590_n1893), .Y(DP_OP_102J5_124_3590_n1861) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1252 ( .A1(n206), .A2(
        DP_OP_102J5_124_3590_n1892), .Y(DP_OP_102J5_124_3590_n1860) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1251 ( .A1(n206), .A2(
        DP_OP_102J5_124_3590_n1891), .Y(DP_OP_102J5_124_3590_n1859) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1250 ( .A1(n206), .A2(
        DP_OP_102J5_124_3590_n1890), .Y(DP_OP_102J5_124_3590_n1858) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1249 ( .A1(n206), .A2(
        DP_OP_102J5_124_3590_n1889), .Y(DP_OP_102J5_124_3590_n1857) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1236 ( .A1(n241), .A2(
        DP_OP_102J5_124_3590_n1852), .Y(DP_OP_102J5_124_3590_n1844) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1235 ( .A1(n241), .A2(
        DP_OP_102J5_124_3590_n1851), .Y(DP_OP_102J5_124_3590_n1843) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1234 ( .A1(n241), .A2(
        DP_OP_102J5_124_3590_n1850), .Y(DP_OP_102J5_124_3590_n1842) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1233 ( .A1(n241), .A2(
        DP_OP_102J5_124_3590_n1849), .Y(DP_OP_102J5_124_3590_n1841) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1232 ( .A1(n241), .A2(
        DP_OP_102J5_124_3590_n1848), .Y(DP_OP_102J5_124_3590_n1840) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1231 ( .A1(n241), .A2(
        DP_OP_102J5_124_3590_n1847), .Y(DP_OP_102J5_124_3590_n1839) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1229 ( .A1(n241), .A2(
        DP_OP_102J5_124_3590_n1845), .Y(DP_OP_102J5_124_3590_n1837) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1228 ( .A1(n240), .A2(
        DP_OP_102J5_124_3590_n1852), .Y(DP_OP_102J5_124_3590_n1836) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1227 ( .A1(n240), .A2(
        DP_OP_102J5_124_3590_n1851), .Y(DP_OP_102J5_124_3590_n1835) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1226 ( .A1(n240), .A2(
        DP_OP_102J5_124_3590_n1850), .Y(DP_OP_102J5_124_3590_n1834) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1225 ( .A1(n240), .A2(
        DP_OP_102J5_124_3590_n1849), .Y(DP_OP_102J5_124_3590_n1833) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1224 ( .A1(n240), .A2(
        DP_OP_102J5_124_3590_n1848), .Y(DP_OP_102J5_124_3590_n1832) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1223 ( .A1(n240), .A2(
        DP_OP_102J5_124_3590_n1847), .Y(DP_OP_102J5_124_3590_n1831) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1222 ( .A1(n240), .A2(
        DP_OP_102J5_124_3590_n1846), .Y(DP_OP_102J5_124_3590_n1830) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1221 ( .A1(n240), .A2(
        DP_OP_102J5_124_3590_n1845), .Y(DP_OP_102J5_124_3590_n1829) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1220 ( .A1(n239), .A2(
        DP_OP_102J5_124_3590_n1852), .Y(DP_OP_102J5_124_3590_n1828) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1219 ( .A1(n239), .A2(
        DP_OP_102J5_124_3590_n1851), .Y(DP_OP_102J5_124_3590_n1827) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1218 ( .A1(n239), .A2(
        DP_OP_102J5_124_3590_n1850), .Y(DP_OP_102J5_124_3590_n1826) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1217 ( .A1(n239), .A2(
        DP_OP_102J5_124_3590_n1849), .Y(DP_OP_102J5_124_3590_n1825) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1216 ( .A1(n239), .A2(
        DP_OP_102J5_124_3590_n1848), .Y(DP_OP_102J5_124_3590_n1824) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1215 ( .A1(n239), .A2(
        DP_OP_102J5_124_3590_n1847), .Y(DP_OP_102J5_124_3590_n1823) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1214 ( .A1(n239), .A2(
        DP_OP_102J5_124_3590_n1846), .Y(DP_OP_102J5_124_3590_n1822) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1213 ( .A1(n239), .A2(
        DP_OP_102J5_124_3590_n1845), .Y(DP_OP_102J5_124_3590_n1821) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1212 ( .A1(n205), .A2(
        DP_OP_102J5_124_3590_n1852), .Y(DP_OP_102J5_124_3590_n1820) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1211 ( .A1(n205), .A2(
        DP_OP_102J5_124_3590_n1851), .Y(DP_OP_102J5_124_3590_n1819) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1210 ( .A1(n205), .A2(
        DP_OP_102J5_124_3590_n1850), .Y(DP_OP_102J5_124_3590_n1818) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1209 ( .A1(n205), .A2(
        DP_OP_102J5_124_3590_n1849), .Y(DP_OP_102J5_124_3590_n1817) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1208 ( .A1(n205), .A2(
        DP_OP_102J5_124_3590_n1848), .Y(DP_OP_102J5_124_3590_n1816) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1207 ( .A1(n205), .A2(
        DP_OP_102J5_124_3590_n1847), .Y(DP_OP_102J5_124_3590_n1815) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1206 ( .A1(n205), .A2(
        DP_OP_102J5_124_3590_n1846), .Y(DP_OP_102J5_124_3590_n453) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1205 ( .A1(n205), .A2(
        DP_OP_102J5_124_3590_n1845), .Y(DP_OP_102J5_124_3590_n1814) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1192 ( .A1(n238), .A2(
        DP_OP_102J5_124_3590_n1809), .Y(DP_OP_102J5_124_3590_n1801) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1191 ( .A1(n238), .A2(
        DP_OP_102J5_124_3590_n1808), .Y(DP_OP_102J5_124_3590_n1800) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1190 ( .A1(n238), .A2(
        DP_OP_102J5_124_3590_n1807), .Y(DP_OP_102J5_124_3590_n1799) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1189 ( .A1(n238), .A2(
        DP_OP_102J5_124_3590_n1806), .Y(DP_OP_102J5_124_3590_n1798) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1188 ( .A1(n238), .A2(
        DP_OP_102J5_124_3590_n1805), .Y(DP_OP_102J5_124_3590_n1797) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1187 ( .A1(n238), .A2(
        DP_OP_102J5_124_3590_n1804), .Y(DP_OP_102J5_124_3590_n1796) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1186 ( .A1(n238), .A2(
        DP_OP_102J5_124_3590_n1803), .Y(DP_OP_102J5_124_3590_n1795) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1185 ( .A1(n238), .A2(
        DP_OP_102J5_124_3590_n1802), .Y(DP_OP_102J5_124_3590_n1794) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1184 ( .A1(n237), .A2(
        DP_OP_102J5_124_3590_n1809), .Y(DP_OP_102J5_124_3590_n1793) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1183 ( .A1(n237), .A2(
        DP_OP_102J5_124_3590_n1808), .Y(DP_OP_102J5_124_3590_n1792) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1182 ( .A1(n237), .A2(
        DP_OP_102J5_124_3590_n1807), .Y(DP_OP_102J5_124_3590_n1791) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1181 ( .A1(n237), .A2(
        DP_OP_102J5_124_3590_n1806), .Y(DP_OP_102J5_124_3590_n1790) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1180 ( .A1(n237), .A2(
        DP_OP_102J5_124_3590_n1805), .Y(DP_OP_102J5_124_3590_n1789) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1179 ( .A1(n237), .A2(
        DP_OP_102J5_124_3590_n1804), .Y(DP_OP_102J5_124_3590_n1788) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1178 ( .A1(n237), .A2(
        DP_OP_102J5_124_3590_n1803), .Y(DP_OP_102J5_124_3590_n1787) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1177 ( .A1(n237), .A2(
        DP_OP_102J5_124_3590_n1802), .Y(DP_OP_102J5_124_3590_n1786) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1176 ( .A1(n236), .A2(
        DP_OP_102J5_124_3590_n1809), .Y(DP_OP_102J5_124_3590_n1785) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1175 ( .A1(n236), .A2(
        DP_OP_102J5_124_3590_n1808), .Y(DP_OP_102J5_124_3590_n1784) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1174 ( .A1(n236), .A2(
        DP_OP_102J5_124_3590_n1807), .Y(DP_OP_102J5_124_3590_n1783) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1173 ( .A1(n236), .A2(
        DP_OP_102J5_124_3590_n1806), .Y(DP_OP_102J5_124_3590_n1782) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1172 ( .A1(n236), .A2(
        DP_OP_102J5_124_3590_n1805), .Y(DP_OP_102J5_124_3590_n1781) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1171 ( .A1(n236), .A2(
        DP_OP_102J5_124_3590_n1804), .Y(DP_OP_102J5_124_3590_n1780) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1170 ( .A1(n236), .A2(
        DP_OP_102J5_124_3590_n1803), .Y(DP_OP_102J5_124_3590_n1779) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1169 ( .A1(n236), .A2(
        DP_OP_102J5_124_3590_n1802), .Y(DP_OP_102J5_124_3590_n1778) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1168 ( .A1(n204), .A2(
        DP_OP_102J5_124_3590_n1809), .Y(DP_OP_102J5_124_3590_n1777) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1167 ( .A1(n204), .A2(
        DP_OP_102J5_124_3590_n1808), .Y(DP_OP_102J5_124_3590_n1776) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1166 ( .A1(n204), .A2(
        DP_OP_102J5_124_3590_n1807), .Y(DP_OP_102J5_124_3590_n1775) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1165 ( .A1(n204), .A2(
        DP_OP_102J5_124_3590_n1806), .Y(DP_OP_102J5_124_3590_n1774) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1164 ( .A1(n204), .A2(
        DP_OP_102J5_124_3590_n1805), .Y(DP_OP_102J5_124_3590_n1773) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1163 ( .A1(n204), .A2(
        DP_OP_102J5_124_3590_n1804), .Y(DP_OP_102J5_124_3590_n1772) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1162 ( .A1(n204), .A2(
        DP_OP_102J5_124_3590_n1803), .Y(DP_OP_102J5_124_3590_n1771) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1161 ( .A1(n204), .A2(
        DP_OP_102J5_124_3590_n1802), .Y(DP_OP_102J5_124_3590_n1770) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1148 ( .A1(n235), .A2(
        DP_OP_102J5_124_3590_n1765), .Y(DP_OP_102J5_124_3590_n1757) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1147 ( .A1(n235), .A2(
        DP_OP_102J5_124_3590_n1764), .Y(DP_OP_102J5_124_3590_n1756) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1146 ( .A1(n235), .A2(
        DP_OP_102J5_124_3590_n1763), .Y(DP_OP_102J5_124_3590_n1755) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1145 ( .A1(n235), .A2(
        DP_OP_102J5_124_3590_n1762), .Y(DP_OP_102J5_124_3590_n1754) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1144 ( .A1(n235), .A2(
        DP_OP_102J5_124_3590_n1761), .Y(DP_OP_102J5_124_3590_n1753) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1143 ( .A1(n235), .A2(
        DP_OP_102J5_124_3590_n1760), .Y(DP_OP_102J5_124_3590_n1752) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1142 ( .A1(n235), .A2(
        DP_OP_102J5_124_3590_n1759), .Y(DP_OP_102J5_124_3590_n1751) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1141 ( .A1(n235), .A2(
        DP_OP_102J5_124_3590_n1758), .Y(DP_OP_102J5_124_3590_n1750) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1140 ( .A1(n234), .A2(
        DP_OP_102J5_124_3590_n1765), .Y(DP_OP_102J5_124_3590_n1749) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1139 ( .A1(n234), .A2(
        DP_OP_102J5_124_3590_n1764), .Y(DP_OP_102J5_124_3590_n1748) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1138 ( .A1(n234), .A2(
        DP_OP_102J5_124_3590_n1763), .Y(DP_OP_102J5_124_3590_n1747) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1137 ( .A1(n234), .A2(
        DP_OP_102J5_124_3590_n1762), .Y(DP_OP_102J5_124_3590_n1746) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1136 ( .A1(n234), .A2(
        DP_OP_102J5_124_3590_n1761), .Y(DP_OP_102J5_124_3590_n1745) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1135 ( .A1(n234), .A2(
        DP_OP_102J5_124_3590_n1760), .Y(DP_OP_102J5_124_3590_n1744) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1134 ( .A1(n234), .A2(
        DP_OP_102J5_124_3590_n1759), .Y(DP_OP_102J5_124_3590_n1743) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1133 ( .A1(n234), .A2(
        DP_OP_102J5_124_3590_n1758), .Y(DP_OP_102J5_124_3590_n1742) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1132 ( .A1(n233), .A2(
        DP_OP_102J5_124_3590_n1765), .Y(DP_OP_102J5_124_3590_n1741) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1131 ( .A1(n233), .A2(
        DP_OP_102J5_124_3590_n1764), .Y(DP_OP_102J5_124_3590_n1740) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1130 ( .A1(n233), .A2(
        DP_OP_102J5_124_3590_n1763), .Y(DP_OP_102J5_124_3590_n1739) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1129 ( .A1(n233), .A2(
        DP_OP_102J5_124_3590_n1762), .Y(DP_OP_102J5_124_3590_n1738) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1128 ( .A1(n233), .A2(
        DP_OP_102J5_124_3590_n1761), .Y(DP_OP_102J5_124_3590_n1737) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1127 ( .A1(n233), .A2(
        DP_OP_102J5_124_3590_n1760), .Y(DP_OP_102J5_124_3590_n1736) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1126 ( .A1(n233), .A2(
        DP_OP_102J5_124_3590_n1759), .Y(DP_OP_102J5_124_3590_n1735) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1125 ( .A1(n233), .A2(
        DP_OP_102J5_124_3590_n1758), .Y(DP_OP_102J5_124_3590_n1734) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1124 ( .A1(n203), .A2(
        DP_OP_102J5_124_3590_n1765), .Y(DP_OP_102J5_124_3590_n1733) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1123 ( .A1(n203), .A2(
        DP_OP_102J5_124_3590_n1764), .Y(DP_OP_102J5_124_3590_n1732) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1122 ( .A1(n203), .A2(
        DP_OP_102J5_124_3590_n1763), .Y(DP_OP_102J5_124_3590_n1731) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1121 ( .A1(n203), .A2(
        DP_OP_102J5_124_3590_n1762), .Y(DP_OP_102J5_124_3590_n1730) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1120 ( .A1(n203), .A2(
        DP_OP_102J5_124_3590_n1761), .Y(DP_OP_102J5_124_3590_n1729) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1119 ( .A1(n203), .A2(
        DP_OP_102J5_124_3590_n1760), .Y(DP_OP_102J5_124_3590_n1728) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1118 ( .A1(n203), .A2(
        DP_OP_102J5_124_3590_n1759), .Y(DP_OP_102J5_124_3590_n1727) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1117 ( .A1(n203), .A2(
        DP_OP_102J5_124_3590_n1758), .Y(DP_OP_102J5_124_3590_n1726) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1104 ( .A1(n232), .A2(
        DP_OP_102J5_124_3590_n1721), .Y(DP_OP_102J5_124_3590_n1713) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1103 ( .A1(n232), .A2(
        DP_OP_102J5_124_3590_n1720), .Y(DP_OP_102J5_124_3590_n1712) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1102 ( .A1(n232), .A2(
        DP_OP_102J5_124_3590_n1719), .Y(DP_OP_102J5_124_3590_n1711) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1101 ( .A1(n232), .A2(
        DP_OP_102J5_124_3590_n1718), .Y(DP_OP_102J5_124_3590_n1710) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1100 ( .A1(n232), .A2(
        DP_OP_102J5_124_3590_n1717), .Y(DP_OP_102J5_124_3590_n1709) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1099 ( .A1(n232), .A2(
        DP_OP_102J5_124_3590_n1716), .Y(DP_OP_102J5_124_3590_n1708) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1098 ( .A1(n232), .A2(
        DP_OP_102J5_124_3590_n1715), .Y(DP_OP_102J5_124_3590_n1707) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1097 ( .A1(n232), .A2(
        DP_OP_102J5_124_3590_n1714), .Y(DP_OP_102J5_124_3590_n1706) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1096 ( .A1(n231), .A2(
        DP_OP_102J5_124_3590_n1721), .Y(DP_OP_102J5_124_3590_n1705) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1095 ( .A1(n231), .A2(
        DP_OP_102J5_124_3590_n1720), .Y(DP_OP_102J5_124_3590_n1704) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1094 ( .A1(n231), .A2(
        DP_OP_102J5_124_3590_n1719), .Y(DP_OP_102J5_124_3590_n1703) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1093 ( .A1(n231), .A2(
        DP_OP_102J5_124_3590_n1718), .Y(DP_OP_102J5_124_3590_n1702) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1092 ( .A1(n231), .A2(
        DP_OP_102J5_124_3590_n1717), .Y(DP_OP_102J5_124_3590_n1701) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1091 ( .A1(n231), .A2(
        DP_OP_102J5_124_3590_n1716), .Y(DP_OP_102J5_124_3590_n1700) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1090 ( .A1(n231), .A2(
        DP_OP_102J5_124_3590_n1715), .Y(DP_OP_102J5_124_3590_n1699) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1089 ( .A1(n231), .A2(
        DP_OP_102J5_124_3590_n1714), .Y(DP_OP_102J5_124_3590_n1698) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1088 ( .A1(n230), .A2(
        DP_OP_102J5_124_3590_n1721), .Y(DP_OP_102J5_124_3590_n1697) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1087 ( .A1(n230), .A2(
        DP_OP_102J5_124_3590_n1720), .Y(DP_OP_102J5_124_3590_n1696) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1086 ( .A1(n230), .A2(
        DP_OP_102J5_124_3590_n1719), .Y(DP_OP_102J5_124_3590_n1695) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1085 ( .A1(n230), .A2(
        DP_OP_102J5_124_3590_n1718), .Y(DP_OP_102J5_124_3590_n1694) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1084 ( .A1(n230), .A2(
        DP_OP_102J5_124_3590_n1717), .Y(DP_OP_102J5_124_3590_n1693) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1083 ( .A1(n230), .A2(
        DP_OP_102J5_124_3590_n1716), .Y(DP_OP_102J5_124_3590_n1692) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1082 ( .A1(n230), .A2(
        DP_OP_102J5_124_3590_n1715), .Y(DP_OP_102J5_124_3590_n1691) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1081 ( .A1(n230), .A2(
        DP_OP_102J5_124_3590_n1714), .Y(DP_OP_102J5_124_3590_n1690) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1080 ( .A1(n202), .A2(
        DP_OP_102J5_124_3590_n1721), .Y(DP_OP_102J5_124_3590_n1689) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1079 ( .A1(n202), .A2(
        DP_OP_102J5_124_3590_n1720), .Y(DP_OP_102J5_124_3590_n1688) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1078 ( .A1(n202), .A2(
        DP_OP_102J5_124_3590_n1719), .Y(DP_OP_102J5_124_3590_n1687) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1077 ( .A1(n202), .A2(
        DP_OP_102J5_124_3590_n1718), .Y(DP_OP_102J5_124_3590_n1686) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1076 ( .A1(n202), .A2(
        DP_OP_102J5_124_3590_n1717), .Y(DP_OP_102J5_124_3590_n1685) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1075 ( .A1(n202), .A2(
        DP_OP_102J5_124_3590_n1716), .Y(DP_OP_102J5_124_3590_n1684) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1074 ( .A1(n202), .A2(
        DP_OP_102J5_124_3590_n1715), .Y(DP_OP_102J5_124_3590_n1683) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1073 ( .A1(n202), .A2(
        DP_OP_102J5_124_3590_n1714), .Y(DP_OP_102J5_124_3590_n1682) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1060 ( .A1(n229), .A2(
        DP_OP_102J5_124_3590_n1677), .Y(DP_OP_102J5_124_3590_n1669) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1059 ( .A1(n229), .A2(
        DP_OP_102J5_124_3590_n1676), .Y(DP_OP_102J5_124_3590_n1668) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1058 ( .A1(n229), .A2(
        DP_OP_102J5_124_3590_n1675), .Y(DP_OP_102J5_124_3590_n1667) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1057 ( .A1(n229), .A2(
        DP_OP_102J5_124_3590_n1674), .Y(DP_OP_102J5_124_3590_n1666) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1056 ( .A1(n229), .A2(
        DP_OP_102J5_124_3590_n1673), .Y(DP_OP_102J5_124_3590_n1665) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1055 ( .A1(n229), .A2(
        DP_OP_102J5_124_3590_n1672), .Y(DP_OP_102J5_124_3590_n1664) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1054 ( .A1(n229), .A2(
        DP_OP_102J5_124_3590_n1671), .Y(DP_OP_102J5_124_3590_n1663) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1053 ( .A1(n229), .A2(
        DP_OP_102J5_124_3590_n1670), .Y(DP_OP_102J5_124_3590_n1662) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1052 ( .A1(n228), .A2(
        DP_OP_102J5_124_3590_n1677), .Y(DP_OP_102J5_124_3590_n1661) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1051 ( .A1(n228), .A2(
        DP_OP_102J5_124_3590_n1676), .Y(DP_OP_102J5_124_3590_n1660) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1050 ( .A1(n228), .A2(
        DP_OP_102J5_124_3590_n1675), .Y(DP_OP_102J5_124_3590_n1659) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1049 ( .A1(n228), .A2(
        DP_OP_102J5_124_3590_n1674), .Y(DP_OP_102J5_124_3590_n1658) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1048 ( .A1(n228), .A2(
        DP_OP_102J5_124_3590_n1673), .Y(DP_OP_102J5_124_3590_n1657) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1047 ( .A1(n228), .A2(
        DP_OP_102J5_124_3590_n1672), .Y(DP_OP_102J5_124_3590_n1656) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1046 ( .A1(n228), .A2(
        DP_OP_102J5_124_3590_n1671), .Y(DP_OP_102J5_124_3590_n1655) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1045 ( .A1(n228), .A2(
        DP_OP_102J5_124_3590_n1670), .Y(DP_OP_102J5_124_3590_n1654) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1044 ( .A1(n227), .A2(
        DP_OP_102J5_124_3590_n1677), .Y(DP_OP_102J5_124_3590_n1653) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1043 ( .A1(n227), .A2(
        DP_OP_102J5_124_3590_n1676), .Y(DP_OP_102J5_124_3590_n1652) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1042 ( .A1(n227), .A2(
        DP_OP_102J5_124_3590_n1675), .Y(DP_OP_102J5_124_3590_n1651) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1041 ( .A1(n227), .A2(
        DP_OP_102J5_124_3590_n1674), .Y(DP_OP_102J5_124_3590_n1650) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1040 ( .A1(n227), .A2(
        DP_OP_102J5_124_3590_n1673), .Y(DP_OP_102J5_124_3590_n1649) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1039 ( .A1(n227), .A2(
        DP_OP_102J5_124_3590_n1672), .Y(DP_OP_102J5_124_3590_n1648) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1038 ( .A1(n227), .A2(
        DP_OP_102J5_124_3590_n1671), .Y(DP_OP_102J5_124_3590_n1647) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1037 ( .A1(n227), .A2(
        DP_OP_102J5_124_3590_n1670), .Y(DP_OP_102J5_124_3590_n1646) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1036 ( .A1(n201), .A2(
        DP_OP_102J5_124_3590_n1677), .Y(DP_OP_102J5_124_3590_n1645) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1035 ( .A1(n201), .A2(
        DP_OP_102J5_124_3590_n1676), .Y(DP_OP_102J5_124_3590_n1644) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1034 ( .A1(n201), .A2(
        DP_OP_102J5_124_3590_n1675), .Y(DP_OP_102J5_124_3590_n1643) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1033 ( .A1(n201), .A2(
        DP_OP_102J5_124_3590_n1674), .Y(DP_OP_102J5_124_3590_n1642) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1032 ( .A1(n201), .A2(
        DP_OP_102J5_124_3590_n1673), .Y(DP_OP_102J5_124_3590_n1641) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1031 ( .A1(n201), .A2(
        DP_OP_102J5_124_3590_n1672), .Y(DP_OP_102J5_124_3590_n1640) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1030 ( .A1(n201), .A2(
        DP_OP_102J5_124_3590_n1671), .Y(DP_OP_102J5_124_3590_n1639) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1029 ( .A1(n201), .A2(
        DP_OP_102J5_124_3590_n1670), .Y(DP_OP_102J5_124_3590_n1638) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1016 ( .A1(n226), .A2(
        DP_OP_102J5_124_3590_n1633), .Y(DP_OP_102J5_124_3590_n1625) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1015 ( .A1(n226), .A2(
        DP_OP_102J5_124_3590_n1632), .Y(DP_OP_102J5_124_3590_n1624) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1014 ( .A1(n226), .A2(
        DP_OP_102J5_124_3590_n1631), .Y(DP_OP_102J5_124_3590_n1623) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1013 ( .A1(n226), .A2(
        DP_OP_102J5_124_3590_n1630), .Y(DP_OP_102J5_124_3590_n1622) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1012 ( .A1(n226), .A2(
        DP_OP_102J5_124_3590_n1629), .Y(DP_OP_102J5_124_3590_n1621) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1011 ( .A1(n226), .A2(
        DP_OP_102J5_124_3590_n1628), .Y(DP_OP_102J5_124_3590_n1620) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1010 ( .A1(n226), .A2(
        DP_OP_102J5_124_3590_n1627), .Y(DP_OP_102J5_124_3590_n1619) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1009 ( .A1(n226), .A2(
        DP_OP_102J5_124_3590_n1626), .Y(DP_OP_102J5_124_3590_n1618) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1008 ( .A1(n225), .A2(
        DP_OP_102J5_124_3590_n1633), .Y(DP_OP_102J5_124_3590_n1617) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1007 ( .A1(n225), .A2(
        DP_OP_102J5_124_3590_n1632), .Y(DP_OP_102J5_124_3590_n1616) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1006 ( .A1(n225), .A2(
        DP_OP_102J5_124_3590_n1631), .Y(DP_OP_102J5_124_3590_n1615) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1005 ( .A1(n225), .A2(
        DP_OP_102J5_124_3590_n1630), .Y(DP_OP_102J5_124_3590_n1614) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1004 ( .A1(n225), .A2(
        DP_OP_102J5_124_3590_n1629), .Y(DP_OP_102J5_124_3590_n1613) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1003 ( .A1(n225), .A2(
        DP_OP_102J5_124_3590_n1628), .Y(DP_OP_102J5_124_3590_n1612) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1002 ( .A1(n225), .A2(
        DP_OP_102J5_124_3590_n1627), .Y(DP_OP_102J5_124_3590_n1611) );
  OR2X1_HVT DP_OP_102J5_124_3590_U1001 ( .A1(n225), .A2(
        DP_OP_102J5_124_3590_n1626), .Y(DP_OP_102J5_124_3590_n1610) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U1000 ( .A1(n224), .A2(
        DP_OP_102J5_124_3590_n1633), .Y(DP_OP_102J5_124_3590_n1609) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U999 ( .A1(n224), .A2(
        DP_OP_102J5_124_3590_n1632), .Y(DP_OP_102J5_124_3590_n1608) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U998 ( .A1(n224), .A2(
        DP_OP_102J5_124_3590_n1631), .Y(DP_OP_102J5_124_3590_n1607) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U997 ( .A1(n224), .A2(
        DP_OP_102J5_124_3590_n1630), .Y(DP_OP_102J5_124_3590_n1606) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U996 ( .A1(n224), .A2(
        DP_OP_102J5_124_3590_n1629), .Y(DP_OP_102J5_124_3590_n1605) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U995 ( .A1(n224), .A2(
        DP_OP_102J5_124_3590_n1628), .Y(DP_OP_102J5_124_3590_n1604) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U994 ( .A1(n224), .A2(
        DP_OP_102J5_124_3590_n1627), .Y(DP_OP_102J5_124_3590_n1603) );
  OR2X1_HVT DP_OP_102J5_124_3590_U993 ( .A1(n224), .A2(
        DP_OP_102J5_124_3590_n1626), .Y(DP_OP_102J5_124_3590_n1602) );
  OR2X1_HVT DP_OP_102J5_124_3590_U992 ( .A1(n200), .A2(
        DP_OP_102J5_124_3590_n1633), .Y(DP_OP_102J5_124_3590_n1601) );
  OR2X1_HVT DP_OP_102J5_124_3590_U991 ( .A1(n200), .A2(
        DP_OP_102J5_124_3590_n1632), .Y(DP_OP_102J5_124_3590_n1600) );
  OR2X1_HVT DP_OP_102J5_124_3590_U990 ( .A1(n200), .A2(
        DP_OP_102J5_124_3590_n1631), .Y(DP_OP_102J5_124_3590_n1599) );
  OR2X1_HVT DP_OP_102J5_124_3590_U989 ( .A1(n200), .A2(
        DP_OP_102J5_124_3590_n1630), .Y(DP_OP_102J5_124_3590_n1598) );
  OR2X1_HVT DP_OP_102J5_124_3590_U988 ( .A1(n200), .A2(
        DP_OP_102J5_124_3590_n1629), .Y(DP_OP_102J5_124_3590_n1597) );
  OR2X1_HVT DP_OP_102J5_124_3590_U987 ( .A1(n200), .A2(
        DP_OP_102J5_124_3590_n1628), .Y(DP_OP_102J5_124_3590_n1596) );
  OR2X1_HVT DP_OP_102J5_124_3590_U986 ( .A1(n200), .A2(
        DP_OP_102J5_124_3590_n1627), .Y(DP_OP_102J5_124_3590_n1595) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U985 ( .A1(n200), .A2(
        DP_OP_102J5_124_3590_n1626), .Y(DP_OP_102J5_124_3590_n1594) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U972 ( .A1(n223), .A2(
        DP_OP_102J5_124_3590_n1589), .Y(DP_OP_102J5_124_3590_n1581) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U971 ( .A1(n223), .A2(
        DP_OP_102J5_124_3590_n1588), .Y(DP_OP_102J5_124_3590_n1580) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U970 ( .A1(n223), .A2(
        DP_OP_102J5_124_3590_n1587), .Y(DP_OP_102J5_124_3590_n1579) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U969 ( .A1(n223), .A2(
        DP_OP_102J5_124_3590_n1586), .Y(DP_OP_102J5_124_3590_n1578) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U968 ( .A1(n223), .A2(
        DP_OP_102J5_124_3590_n1585), .Y(DP_OP_102J5_124_3590_n1577) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U967 ( .A1(n223), .A2(
        DP_OP_102J5_124_3590_n1584), .Y(DP_OP_102J5_124_3590_n1576) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U966 ( .A1(n223), .A2(
        DP_OP_102J5_124_3590_n1583), .Y(DP_OP_102J5_124_3590_n1575) );
  OR2X1_HVT DP_OP_102J5_124_3590_U965 ( .A1(n223), .A2(
        DP_OP_102J5_124_3590_n1582), .Y(DP_OP_102J5_124_3590_n1574) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U964 ( .A1(n222), .A2(
        DP_OP_102J5_124_3590_n1589), .Y(DP_OP_102J5_124_3590_n1573) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U963 ( .A1(n222), .A2(
        DP_OP_102J5_124_3590_n1588), .Y(DP_OP_102J5_124_3590_n1572) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U962 ( .A1(n222), .A2(
        DP_OP_102J5_124_3590_n1587), .Y(DP_OP_102J5_124_3590_n1571) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U961 ( .A1(n222), .A2(
        DP_OP_102J5_124_3590_n1586), .Y(DP_OP_102J5_124_3590_n1570) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U960 ( .A1(n222), .A2(
        DP_OP_102J5_124_3590_n1585), .Y(DP_OP_102J5_124_3590_n1569) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U959 ( .A1(n222), .A2(
        DP_OP_102J5_124_3590_n1584), .Y(DP_OP_102J5_124_3590_n1568) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U958 ( .A1(n222), .A2(
        DP_OP_102J5_124_3590_n1583), .Y(DP_OP_102J5_124_3590_n1567) );
  OR2X1_HVT DP_OP_102J5_124_3590_U957 ( .A1(n222), .A2(
        DP_OP_102J5_124_3590_n1582), .Y(DP_OP_102J5_124_3590_n1566) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U956 ( .A1(n221), .A2(
        DP_OP_102J5_124_3590_n1589), .Y(DP_OP_102J5_124_3590_n1565) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U955 ( .A1(n221), .A2(
        DP_OP_102J5_124_3590_n1588), .Y(DP_OP_102J5_124_3590_n1564) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U954 ( .A1(n221), .A2(
        DP_OP_102J5_124_3590_n1587), .Y(DP_OP_102J5_124_3590_n1563) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U953 ( .A1(n221), .A2(
        DP_OP_102J5_124_3590_n1586), .Y(DP_OP_102J5_124_3590_n1562) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U952 ( .A1(n221), .A2(
        DP_OP_102J5_124_3590_n1585), .Y(DP_OP_102J5_124_3590_n1561) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U951 ( .A1(n221), .A2(
        DP_OP_102J5_124_3590_n1584), .Y(DP_OP_102J5_124_3590_n1560) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U950 ( .A1(n221), .A2(
        DP_OP_102J5_124_3590_n1583), .Y(DP_OP_102J5_124_3590_n1559) );
  OR2X1_HVT DP_OP_102J5_124_3590_U949 ( .A1(n221), .A2(
        DP_OP_102J5_124_3590_n1582), .Y(DP_OP_102J5_124_3590_n1558) );
  OR2X1_HVT DP_OP_102J5_124_3590_U948 ( .A1(n199), .A2(
        DP_OP_102J5_124_3590_n1589), .Y(DP_OP_102J5_124_3590_n1557) );
  OR2X1_HVT DP_OP_102J5_124_3590_U947 ( .A1(n199), .A2(
        DP_OP_102J5_124_3590_n1588), .Y(DP_OP_102J5_124_3590_n1556) );
  OR2X1_HVT DP_OP_102J5_124_3590_U946 ( .A1(n199), .A2(
        DP_OP_102J5_124_3590_n1587), .Y(DP_OP_102J5_124_3590_n1555) );
  OR2X1_HVT DP_OP_102J5_124_3590_U945 ( .A1(n199), .A2(
        DP_OP_102J5_124_3590_n1586), .Y(DP_OP_102J5_124_3590_n1554) );
  OR2X1_HVT DP_OP_102J5_124_3590_U944 ( .A1(n199), .A2(
        DP_OP_102J5_124_3590_n1585), .Y(DP_OP_102J5_124_3590_n1553) );
  OR2X1_HVT DP_OP_102J5_124_3590_U943 ( .A1(n199), .A2(
        DP_OP_102J5_124_3590_n1584), .Y(DP_OP_102J5_124_3590_n1552) );
  OR2X1_HVT DP_OP_102J5_124_3590_U942 ( .A1(n199), .A2(
        DP_OP_102J5_124_3590_n1583), .Y(DP_OP_102J5_124_3590_n1551) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U941 ( .A1(n199), .A2(
        DP_OP_102J5_124_3590_n1582), .Y(DP_OP_102J5_124_3590_n1550) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U928 ( .A1(n220), .A2(
        DP_OP_102J5_124_3590_n1545), .Y(DP_OP_102J5_124_3590_n1537) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U927 ( .A1(n220), .A2(
        DP_OP_102J5_124_3590_n1544), .Y(DP_OP_102J5_124_3590_n1536) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U926 ( .A1(n220), .A2(
        DP_OP_102J5_124_3590_n1543), .Y(DP_OP_102J5_124_3590_n1535) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U925 ( .A1(n220), .A2(
        DP_OP_102J5_124_3590_n1542), .Y(DP_OP_102J5_124_3590_n1534) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U924 ( .A1(n220), .A2(
        DP_OP_102J5_124_3590_n1541), .Y(DP_OP_102J5_124_3590_n1533) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U923 ( .A1(n220), .A2(
        DP_OP_102J5_124_3590_n1540), .Y(DP_OP_102J5_124_3590_n1532) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U922 ( .A1(n220), .A2(
        DP_OP_102J5_124_3590_n1539), .Y(DP_OP_102J5_124_3590_n1531) );
  OR2X1_HVT DP_OP_102J5_124_3590_U921 ( .A1(n220), .A2(
        DP_OP_102J5_124_3590_n1538), .Y(DP_OP_102J5_124_3590_n1530) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U920 ( .A1(n219), .A2(
        DP_OP_102J5_124_3590_n1545), .Y(DP_OP_102J5_124_3590_n1529) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U919 ( .A1(n219), .A2(
        DP_OP_102J5_124_3590_n1544), .Y(DP_OP_102J5_124_3590_n1528) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U918 ( .A1(n219), .A2(
        DP_OP_102J5_124_3590_n1543), .Y(DP_OP_102J5_124_3590_n1527) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U917 ( .A1(n219), .A2(
        DP_OP_102J5_124_3590_n1542), .Y(DP_OP_102J5_124_3590_n1526) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U916 ( .A1(n219), .A2(
        DP_OP_102J5_124_3590_n1541), .Y(DP_OP_102J5_124_3590_n1525) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U915 ( .A1(n219), .A2(
        DP_OP_102J5_124_3590_n1540), .Y(DP_OP_102J5_124_3590_n1524) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U914 ( .A1(n219), .A2(
        DP_OP_102J5_124_3590_n1539), .Y(DP_OP_102J5_124_3590_n1523) );
  OR2X1_HVT DP_OP_102J5_124_3590_U913 ( .A1(n219), .A2(
        DP_OP_102J5_124_3590_n1538), .Y(DP_OP_102J5_124_3590_n1522) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U912 ( .A1(n218), .A2(
        DP_OP_102J5_124_3590_n1545), .Y(DP_OP_102J5_124_3590_n1521) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U911 ( .A1(n218), .A2(
        DP_OP_102J5_124_3590_n1544), .Y(DP_OP_102J5_124_3590_n1520) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U910 ( .A1(n218), .A2(
        DP_OP_102J5_124_3590_n1543), .Y(DP_OP_102J5_124_3590_n1519) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U909 ( .A1(n218), .A2(
        DP_OP_102J5_124_3590_n1542), .Y(DP_OP_102J5_124_3590_n1518) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U908 ( .A1(n218), .A2(
        DP_OP_102J5_124_3590_n1541), .Y(DP_OP_102J5_124_3590_n1517) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U907 ( .A1(n218), .A2(
        DP_OP_102J5_124_3590_n1540), .Y(DP_OP_102J5_124_3590_n1516) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U906 ( .A1(n218), .A2(
        DP_OP_102J5_124_3590_n1539), .Y(DP_OP_102J5_124_3590_n1515) );
  OR2X1_HVT DP_OP_102J5_124_3590_U905 ( .A1(n218), .A2(
        DP_OP_102J5_124_3590_n1538), .Y(DP_OP_102J5_124_3590_n1514) );
  OR2X1_HVT DP_OP_102J5_124_3590_U904 ( .A1(n198), .A2(
        DP_OP_102J5_124_3590_n1545), .Y(DP_OP_102J5_124_3590_n1513) );
  OR2X1_HVT DP_OP_102J5_124_3590_U903 ( .A1(n198), .A2(
        DP_OP_102J5_124_3590_n1544), .Y(DP_OP_102J5_124_3590_n1512) );
  OR2X1_HVT DP_OP_102J5_124_3590_U902 ( .A1(n198), .A2(
        DP_OP_102J5_124_3590_n1543), .Y(DP_OP_102J5_124_3590_n1511) );
  OR2X1_HVT DP_OP_102J5_124_3590_U901 ( .A1(n198), .A2(
        DP_OP_102J5_124_3590_n1542), .Y(DP_OP_102J5_124_3590_n1510) );
  OR2X1_HVT DP_OP_102J5_124_3590_U900 ( .A1(n198), .A2(
        DP_OP_102J5_124_3590_n1541), .Y(DP_OP_102J5_124_3590_n1509) );
  OR2X1_HVT DP_OP_102J5_124_3590_U899 ( .A1(n198), .A2(
        DP_OP_102J5_124_3590_n1540), .Y(DP_OP_102J5_124_3590_n1508) );
  OR2X1_HVT DP_OP_102J5_124_3590_U898 ( .A1(n198), .A2(
        DP_OP_102J5_124_3590_n1539), .Y(DP_OP_102J5_124_3590_n1507) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U897 ( .A1(n198), .A2(
        DP_OP_102J5_124_3590_n1538), .Y(DP_OP_102J5_124_3590_n1506) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U858 ( .A1(n287), .A2(n191), .Y(
        DP_OP_102J5_124_3590_n204) );
  FADDX1_HVT DP_OP_102J5_124_3590_U849 ( .A(DP_OP_102J5_124_3590_n1581), .B(
        DP_OP_102J5_124_3590_n1537), .CI(DP_OP_102J5_124_3590_n1625), .CO(
        DP_OP_102J5_124_3590_n1465), .S(DP_OP_102J5_124_3590_n1466) );
  FADDX1_HVT DP_OP_102J5_124_3590_U848 ( .A(DP_OP_102J5_124_3590_n1713), .B(
        DP_OP_102J5_124_3590_n1669), .CI(DP_OP_102J5_124_3590_n1757), .CO(
        DP_OP_102J5_124_3590_n1463), .S(DP_OP_102J5_124_3590_n1464) );
  FADDX1_HVT DP_OP_102J5_124_3590_U847 ( .A(DP_OP_102J5_124_3590_n1844), .B(
        DP_OP_102J5_124_3590_n1801), .CI(DP_OP_102J5_124_3590_n1888), .CO(
        DP_OP_102J5_124_3590_n1461), .S(DP_OP_102J5_124_3590_n1462) );
  FADDX1_HVT DP_OP_102J5_124_3590_U846 ( .A(DP_OP_102J5_124_3590_n1976), .B(
        DP_OP_102J5_124_3590_n1932), .CI(DP_OP_102J5_124_3590_n2020), .CO(
        DP_OP_102J5_124_3590_n1459), .S(DP_OP_102J5_124_3590_n1460) );
  FADDX1_HVT DP_OP_102J5_124_3590_U845 ( .A(DP_OP_102J5_124_3590_n2108), .B(
        DP_OP_102J5_124_3590_n2064), .CI(DP_OP_102J5_124_3590_n2152), .CO(
        DP_OP_102J5_124_3590_n1457), .S(DP_OP_102J5_124_3590_n1458) );
  FADDX1_HVT DP_OP_102J5_124_3590_U844 ( .A(DP_OP_102J5_124_3590_n2371), .B(
        DP_OP_102J5_124_3590_n2196), .CI(DP_OP_102J5_124_3590_n2240), .CO(
        DP_OP_102J5_124_3590_n1455), .S(DP_OP_102J5_124_3590_n1456) );
  FADDX1_HVT DP_OP_102J5_124_3590_U843 ( .A(DP_OP_102J5_124_3590_n2328), .B(
        DP_OP_102J5_124_3590_n2284), .CI(DP_OP_102J5_124_3590_n1460), .CO(
        DP_OP_102J5_124_3590_n1453), .S(DP_OP_102J5_124_3590_n1454) );
  FADDX1_HVT DP_OP_102J5_124_3590_U842 ( .A(DP_OP_102J5_124_3590_n1456), .B(
        DP_OP_102J5_124_3590_n1462), .CI(DP_OP_102J5_124_3590_n1464), .CO(
        DP_OP_102J5_124_3590_n1451), .S(DP_OP_102J5_124_3590_n1452) );
  FADDX1_HVT DP_OP_102J5_124_3590_U841 ( .A(DP_OP_102J5_124_3590_n1458), .B(
        DP_OP_102J5_124_3590_n1466), .CI(DP_OP_102J5_124_3590_n1481), .CO(
        DP_OP_102J5_124_3590_n1449), .S(DP_OP_102J5_124_3590_n1450) );
  FADDX1_HVT DP_OP_102J5_124_3590_U840 ( .A(DP_OP_102J5_124_3590_n1536), .B(
        DP_OP_102J5_124_3590_n1529), .CI(DP_OP_102J5_124_3590_n1573), .CO(
        DP_OP_102J5_124_3590_n1447), .S(DP_OP_102J5_124_3590_n1448) );
  FADDX1_HVT DP_OP_102J5_124_3590_U839 ( .A(DP_OP_102J5_124_3590_n1617), .B(
        DP_OP_102J5_124_3590_n1580), .CI(DP_OP_102J5_124_3590_n1624), .CO(
        DP_OP_102J5_124_3590_n1445), .S(DP_OP_102J5_124_3590_n1446) );
  FADDX1_HVT DP_OP_102J5_124_3590_U838 ( .A(DP_OP_102J5_124_3590_n1668), .B(
        DP_OP_102J5_124_3590_n1661), .CI(DP_OP_102J5_124_3590_n1705), .CO(
        DP_OP_102J5_124_3590_n1443), .S(DP_OP_102J5_124_3590_n1444) );
  FADDX1_HVT DP_OP_102J5_124_3590_U837 ( .A(DP_OP_102J5_124_3590_n1749), .B(
        DP_OP_102J5_124_3590_n1712), .CI(DP_OP_102J5_124_3590_n1756), .CO(
        DP_OP_102J5_124_3590_n1441), .S(DP_OP_102J5_124_3590_n1442) );
  FADDX1_HVT DP_OP_102J5_124_3590_U836 ( .A(DP_OP_102J5_124_3590_n1800), .B(
        DP_OP_102J5_124_3590_n1793), .CI(DP_OP_102J5_124_3590_n1836), .CO(
        DP_OP_102J5_124_3590_n1439), .S(DP_OP_102J5_124_3590_n1440) );
  FADDX1_HVT DP_OP_102J5_124_3590_U835 ( .A(DP_OP_102J5_124_3590_n1880), .B(
        DP_OP_102J5_124_3590_n1843), .CI(DP_OP_102J5_124_3590_n1887), .CO(
        DP_OP_102J5_124_3590_n1437), .S(DP_OP_102J5_124_3590_n1438) );
  FADDX1_HVT DP_OP_102J5_124_3590_U834 ( .A(DP_OP_102J5_124_3590_n1931), .B(
        DP_OP_102J5_124_3590_n1924), .CI(DP_OP_102J5_124_3590_n1968), .CO(
        DP_OP_102J5_124_3590_n1435), .S(DP_OP_102J5_124_3590_n1436) );
  FADDX1_HVT DP_OP_102J5_124_3590_U833 ( .A(DP_OP_102J5_124_3590_n2012), .B(
        DP_OP_102J5_124_3590_n1975), .CI(DP_OP_102J5_124_3590_n2370), .CO(
        DP_OP_102J5_124_3590_n1433), .S(DP_OP_102J5_124_3590_n1434) );
  FADDX1_HVT DP_OP_102J5_124_3590_U832 ( .A(DP_OP_102J5_124_3590_n2364), .B(
        DP_OP_102J5_124_3590_n2019), .CI(DP_OP_102J5_124_3590_n2056), .CO(
        DP_OP_102J5_124_3590_n1431), .S(DP_OP_102J5_124_3590_n1432) );
  FADDX1_HVT DP_OP_102J5_124_3590_U831 ( .A(DP_OP_102J5_124_3590_n2195), .B(
        DP_OP_102J5_124_3590_n2327), .CI(DP_OP_102J5_124_3590_n2320), .CO(
        DP_OP_102J5_124_3590_n1429), .S(DP_OP_102J5_124_3590_n1430) );
  FADDX1_HVT DP_OP_102J5_124_3590_U830 ( .A(DP_OP_102J5_124_3590_n2283), .B(
        DP_OP_102J5_124_3590_n2063), .CI(DP_OP_102J5_124_3590_n2100), .CO(
        DP_OP_102J5_124_3590_n1427), .S(DP_OP_102J5_124_3590_n1428) );
  FADDX1_HVT DP_OP_102J5_124_3590_U829 ( .A(DP_OP_102J5_124_3590_n2276), .B(
        DP_OP_102J5_124_3590_n2107), .CI(DP_OP_102J5_124_3590_n2144), .CO(
        DP_OP_102J5_124_3590_n1425), .S(DP_OP_102J5_124_3590_n1426) );
  FADDX1_HVT DP_OP_102J5_124_3590_U828 ( .A(DP_OP_102J5_124_3590_n2239), .B(
        DP_OP_102J5_124_3590_n2151), .CI(DP_OP_102J5_124_3590_n2188), .CO(
        DP_OP_102J5_124_3590_n1423), .S(DP_OP_102J5_124_3590_n1424) );
  FADDX1_HVT DP_OP_102J5_124_3590_U827 ( .A(DP_OP_102J5_124_3590_n2232), .B(
        DP_OP_102J5_124_3590_n1457), .CI(DP_OP_102J5_124_3590_n1455), .CO(
        DP_OP_102J5_124_3590_n1421), .S(DP_OP_102J5_124_3590_n1422) );
  FADDX1_HVT DP_OP_102J5_124_3590_U826 ( .A(DP_OP_102J5_124_3590_n1463), .B(
        DP_OP_102J5_124_3590_n1459), .CI(DP_OP_102J5_124_3590_n1461), .CO(
        DP_OP_102J5_124_3590_n1419), .S(DP_OP_102J5_124_3590_n1420) );
  FADDX1_HVT DP_OP_102J5_124_3590_U825 ( .A(DP_OP_102J5_124_3590_n1465), .B(
        DP_OP_102J5_124_3590_n1426), .CI(DP_OP_102J5_124_3590_n1428), .CO(
        DP_OP_102J5_124_3590_n1417), .S(DP_OP_102J5_124_3590_n1418) );
  FADDX1_HVT DP_OP_102J5_124_3590_U824 ( .A(DP_OP_102J5_124_3590_n1424), .B(
        DP_OP_102J5_124_3590_n1438), .CI(DP_OP_102J5_124_3590_n1440), .CO(
        DP_OP_102J5_124_3590_n1415), .S(DP_OP_102J5_124_3590_n1416) );
  FADDX1_HVT DP_OP_102J5_124_3590_U823 ( .A(DP_OP_102J5_124_3590_n1430), .B(
        DP_OP_102J5_124_3590_n1444), .CI(DP_OP_102J5_124_3590_n1442), .CO(
        DP_OP_102J5_124_3590_n1413), .S(DP_OP_102J5_124_3590_n1414) );
  FADDX1_HVT DP_OP_102J5_124_3590_U822 ( .A(DP_OP_102J5_124_3590_n1432), .B(
        DP_OP_102J5_124_3590_n1448), .CI(DP_OP_102J5_124_3590_n1446), .CO(
        DP_OP_102J5_124_3590_n1411), .S(DP_OP_102J5_124_3590_n1412) );
  FADDX1_HVT DP_OP_102J5_124_3590_U821 ( .A(DP_OP_102J5_124_3590_n1434), .B(
        DP_OP_102J5_124_3590_n1436), .CI(DP_OP_102J5_124_3590_n1480), .CO(
        DP_OP_102J5_124_3590_n1409), .S(DP_OP_102J5_124_3590_n1410) );
  FADDX1_HVT DP_OP_102J5_124_3590_U820 ( .A(DP_OP_102J5_124_3590_n1453), .B(
        DP_OP_102J5_124_3590_n1422), .CI(DP_OP_102J5_124_3590_n1451), .CO(
        DP_OP_102J5_124_3590_n1407), .S(DP_OP_102J5_124_3590_n1408) );
  FADDX1_HVT DP_OP_102J5_124_3590_U819 ( .A(DP_OP_102J5_124_3590_n1420), .B(
        DP_OP_102J5_124_3590_n1418), .CI(DP_OP_102J5_124_3590_n1412), .CO(
        DP_OP_102J5_124_3590_n1405), .S(DP_OP_102J5_124_3590_n1406) );
  FADDX1_HVT DP_OP_102J5_124_3590_U818 ( .A(DP_OP_102J5_124_3590_n1416), .B(
        DP_OP_102J5_124_3590_n1414), .CI(DP_OP_102J5_124_3590_n1449), .CO(
        DP_OP_102J5_124_3590_n1403), .S(DP_OP_102J5_124_3590_n1404) );
  FADDX1_HVT DP_OP_102J5_124_3590_U817 ( .A(DP_OP_102J5_124_3590_n1410), .B(
        DP_OP_102J5_124_3590_n1408), .CI(DP_OP_102J5_124_3590_n1406), .CO(
        DP_OP_102J5_124_3590_n1401), .S(DP_OP_102J5_124_3590_n1402) );
  HADDX1_HVT DP_OP_102J5_124_3590_U816 ( .A0(DP_OP_102J5_124_3590_n1528), .B0(
        DP_OP_102J5_124_3590_n1535), .C1(DP_OP_102J5_124_3590_n1399), .SO(
        DP_OP_102J5_124_3590_n1400) );
  FADDX1_HVT DP_OP_102J5_124_3590_U815 ( .A(DP_OP_102J5_124_3590_n1565), .B(
        DP_OP_102J5_124_3590_n1521), .CI(DP_OP_102J5_124_3590_n1572), .CO(
        DP_OP_102J5_124_3590_n1397), .S(DP_OP_102J5_124_3590_n1398) );
  FADDX1_HVT DP_OP_102J5_124_3590_U814 ( .A(DP_OP_102J5_124_3590_n1609), .B(
        DP_OP_102J5_124_3590_n1579), .CI(DP_OP_102J5_124_3590_n1616), .CO(
        DP_OP_102J5_124_3590_n1395), .S(DP_OP_102J5_124_3590_n1396) );
  FADDX1_HVT DP_OP_102J5_124_3590_U813 ( .A(DP_OP_102J5_124_3590_n1653), .B(
        DP_OP_102J5_124_3590_n1623), .CI(DP_OP_102J5_124_3590_n1660), .CO(
        DP_OP_102J5_124_3590_n1393), .S(DP_OP_102J5_124_3590_n1394) );
  FADDX1_HVT DP_OP_102J5_124_3590_U812 ( .A(DP_OP_102J5_124_3590_n1697), .B(
        DP_OP_102J5_124_3590_n1667), .CI(DP_OP_102J5_124_3590_n1704), .CO(
        DP_OP_102J5_124_3590_n1391), .S(DP_OP_102J5_124_3590_n1392) );
  FADDX1_HVT DP_OP_102J5_124_3590_U811 ( .A(DP_OP_102J5_124_3590_n1741), .B(
        DP_OP_102J5_124_3590_n1711), .CI(DP_OP_102J5_124_3590_n1748), .CO(
        DP_OP_102J5_124_3590_n1389), .S(DP_OP_102J5_124_3590_n1390) );
  FADDX1_HVT DP_OP_102J5_124_3590_U810 ( .A(DP_OP_102J5_124_3590_n1785), .B(
        DP_OP_102J5_124_3590_n1755), .CI(DP_OP_102J5_124_3590_n1792), .CO(
        DP_OP_102J5_124_3590_n1387), .S(DP_OP_102J5_124_3590_n1388) );
  FADDX1_HVT DP_OP_102J5_124_3590_U809 ( .A(DP_OP_102J5_124_3590_n1828), .B(
        DP_OP_102J5_124_3590_n1799), .CI(DP_OP_102J5_124_3590_n1835), .CO(
        DP_OP_102J5_124_3590_n1385), .S(DP_OP_102J5_124_3590_n1386) );
  FADDX1_HVT DP_OP_102J5_124_3590_U808 ( .A(DP_OP_102J5_124_3590_n1872), .B(
        DP_OP_102J5_124_3590_n1842), .CI(DP_OP_102J5_124_3590_n1879), .CO(
        DP_OP_102J5_124_3590_n1383), .S(DP_OP_102J5_124_3590_n1384) );
  FADDX1_HVT DP_OP_102J5_124_3590_U807 ( .A(DP_OP_102J5_124_3590_n2106), .B(
        DP_OP_102J5_124_3590_n2369), .CI(DP_OP_102J5_124_3590_n2363), .CO(
        DP_OP_102J5_124_3590_n1381), .S(DP_OP_102J5_124_3590_n1382) );
  FADDX1_HVT DP_OP_102J5_124_3590_U806 ( .A(DP_OP_102J5_124_3590_n2092), .B(
        DP_OP_102J5_124_3590_n2356), .CI(DP_OP_102J5_124_3590_n2326), .CO(
        DP_OP_102J5_124_3590_n1379), .S(DP_OP_102J5_124_3590_n1380) );
  FADDX1_HVT DP_OP_102J5_124_3590_U805 ( .A(DP_OP_102J5_124_3590_n2062), .B(
        DP_OP_102J5_124_3590_n1886), .CI(DP_OP_102J5_124_3590_n1916), .CO(
        DP_OP_102J5_124_3590_n1377), .S(DP_OP_102J5_124_3590_n1378) );
  FADDX1_HVT DP_OP_102J5_124_3590_U804 ( .A(DP_OP_102J5_124_3590_n2099), .B(
        DP_OP_102J5_124_3590_n1923), .CI(DP_OP_102J5_124_3590_n1930), .CO(
        DP_OP_102J5_124_3590_n1375), .S(DP_OP_102J5_124_3590_n1376) );
  FADDX1_HVT DP_OP_102J5_124_3590_U803 ( .A(DP_OP_102J5_124_3590_n2136), .B(
        DP_OP_102J5_124_3590_n1960), .CI(DP_OP_102J5_124_3590_n1967), .CO(
        DP_OP_102J5_124_3590_n1373), .S(DP_OP_102J5_124_3590_n1374) );
  FADDX1_HVT DP_OP_102J5_124_3590_U802 ( .A(DP_OP_102J5_124_3590_n2150), .B(
        DP_OP_102J5_124_3590_n1974), .CI(DP_OP_102J5_124_3590_n2319), .CO(
        DP_OP_102J5_124_3590_n1371), .S(DP_OP_102J5_124_3590_n1372) );
  FADDX1_HVT DP_OP_102J5_124_3590_U801 ( .A(DP_OP_102J5_124_3590_n2143), .B(
        DP_OP_102J5_124_3590_n2312), .CI(DP_OP_102J5_124_3590_n2282), .CO(
        DP_OP_102J5_124_3590_n1369), .S(DP_OP_102J5_124_3590_n1370) );
  FADDX1_HVT DP_OP_102J5_124_3590_U800 ( .A(DP_OP_102J5_124_3590_n2275), .B(
        DP_OP_102J5_124_3590_n2004), .CI(DP_OP_102J5_124_3590_n2011), .CO(
        DP_OP_102J5_124_3590_n1367), .S(DP_OP_102J5_124_3590_n1368) );
  FADDX1_HVT DP_OP_102J5_124_3590_U799 ( .A(DP_OP_102J5_124_3590_n2268), .B(
        DP_OP_102J5_124_3590_n2018), .CI(DP_OP_102J5_124_3590_n2048), .CO(
        DP_OP_102J5_124_3590_n1365), .S(DP_OP_102J5_124_3590_n1366) );
  FADDX1_HVT DP_OP_102J5_124_3590_U798 ( .A(DP_OP_102J5_124_3590_n2238), .B(
        DP_OP_102J5_124_3590_n2055), .CI(DP_OP_102J5_124_3590_n2231), .CO(
        DP_OP_102J5_124_3590_n1363), .S(DP_OP_102J5_124_3590_n1364) );
  FADDX1_HVT DP_OP_102J5_124_3590_U797 ( .A(DP_OP_102J5_124_3590_n2224), .B(
        DP_OP_102J5_124_3590_n2180), .CI(DP_OP_102J5_124_3590_n2187), .CO(
        DP_OP_102J5_124_3590_n1361), .S(DP_OP_102J5_124_3590_n1362) );
  FADDX1_HVT DP_OP_102J5_124_3590_U796 ( .A(DP_OP_102J5_124_3590_n2194), .B(
        DP_OP_102J5_124_3590_n1400), .CI(DP_OP_102J5_124_3590_n1425), .CO(
        DP_OP_102J5_124_3590_n1359), .S(DP_OP_102J5_124_3590_n1360) );
  FADDX1_HVT DP_OP_102J5_124_3590_U795 ( .A(DP_OP_102J5_124_3590_n1427), .B(
        DP_OP_102J5_124_3590_n1429), .CI(DP_OP_102J5_124_3590_n1431), .CO(
        DP_OP_102J5_124_3590_n1357), .S(DP_OP_102J5_124_3590_n1358) );
  FADDX1_HVT DP_OP_102J5_124_3590_U794 ( .A(DP_OP_102J5_124_3590_n1441), .B(
        DP_OP_102J5_124_3590_n1433), .CI(DP_OP_102J5_124_3590_n1423), .CO(
        DP_OP_102J5_124_3590_n1355), .S(DP_OP_102J5_124_3590_n1356) );
  FADDX1_HVT DP_OP_102J5_124_3590_U793 ( .A(DP_OP_102J5_124_3590_n1439), .B(
        DP_OP_102J5_124_3590_n1435), .CI(DP_OP_102J5_124_3590_n1437), .CO(
        DP_OP_102J5_124_3590_n1353), .S(DP_OP_102J5_124_3590_n1354) );
  FADDX1_HVT DP_OP_102J5_124_3590_U792 ( .A(DP_OP_102J5_124_3590_n1443), .B(
        DP_OP_102J5_124_3590_n1445), .CI(DP_OP_102J5_124_3590_n1447), .CO(
        DP_OP_102J5_124_3590_n1351), .S(DP_OP_102J5_124_3590_n1352) );
  FADDX1_HVT DP_OP_102J5_124_3590_U791 ( .A(DP_OP_102J5_124_3590_n1376), .B(
        DP_OP_102J5_124_3590_n1388), .CI(DP_OP_102J5_124_3590_n1386), .CO(
        DP_OP_102J5_124_3590_n1349), .S(DP_OP_102J5_124_3590_n1350) );
  FADDX1_HVT DP_OP_102J5_124_3590_U790 ( .A(DP_OP_102J5_124_3590_n1366), .B(
        DP_OP_102J5_124_3590_n1380), .CI(DP_OP_102J5_124_3590_n1378), .CO(
        DP_OP_102J5_124_3590_n1347), .S(DP_OP_102J5_124_3590_n1348) );
  FADDX1_HVT DP_OP_102J5_124_3590_U789 ( .A(DP_OP_102J5_124_3590_n1364), .B(
        DP_OP_102J5_124_3590_n1390), .CI(DP_OP_102J5_124_3590_n1384), .CO(
        DP_OP_102J5_124_3590_n1345), .S(DP_OP_102J5_124_3590_n1346) );
  FADDX1_HVT DP_OP_102J5_124_3590_U788 ( .A(DP_OP_102J5_124_3590_n1370), .B(
        DP_OP_102J5_124_3590_n1392), .CI(DP_OP_102J5_124_3590_n1394), .CO(
        DP_OP_102J5_124_3590_n1343), .S(DP_OP_102J5_124_3590_n1344) );
  FADDX1_HVT DP_OP_102J5_124_3590_U787 ( .A(DP_OP_102J5_124_3590_n1368), .B(
        DP_OP_102J5_124_3590_n1398), .CI(DP_OP_102J5_124_3590_n1396), .CO(
        DP_OP_102J5_124_3590_n1341), .S(DP_OP_102J5_124_3590_n1342) );
  FADDX1_HVT DP_OP_102J5_124_3590_U786 ( .A(DP_OP_102J5_124_3590_n1374), .B(
        DP_OP_102J5_124_3590_n1372), .CI(DP_OP_102J5_124_3590_n1362), .CO(
        DP_OP_102J5_124_3590_n1339), .S(DP_OP_102J5_124_3590_n1340) );
  FADDX1_HVT DP_OP_102J5_124_3590_U785 ( .A(DP_OP_102J5_124_3590_n1382), .B(
        DP_OP_102J5_124_3590_n1421), .CI(DP_OP_102J5_124_3590_n1419), .CO(
        DP_OP_102J5_124_3590_n1337), .S(DP_OP_102J5_124_3590_n1338) );
  FADDX1_HVT DP_OP_102J5_124_3590_U784 ( .A(DP_OP_102J5_124_3590_n1479), .B(
        DP_OP_102J5_124_3590_n1360), .CI(DP_OP_102J5_124_3590_n1417), .CO(
        DP_OP_102J5_124_3590_n1335), .S(DP_OP_102J5_124_3590_n1336) );
  FADDX1_HVT DP_OP_102J5_124_3590_U783 ( .A(DP_OP_102J5_124_3590_n1354), .B(
        DP_OP_102J5_124_3590_n1352), .CI(DP_OP_102J5_124_3590_n1356), .CO(
        DP_OP_102J5_124_3590_n1333), .S(DP_OP_102J5_124_3590_n1334) );
  FADDX1_HVT DP_OP_102J5_124_3590_U782 ( .A(DP_OP_102J5_124_3590_n1415), .B(
        DP_OP_102J5_124_3590_n1358), .CI(DP_OP_102J5_124_3590_n1413), .CO(
        DP_OP_102J5_124_3590_n1331), .S(DP_OP_102J5_124_3590_n1332) );
  FADDX1_HVT DP_OP_102J5_124_3590_U781 ( .A(DP_OP_102J5_124_3590_n1411), .B(
        DP_OP_102J5_124_3590_n1340), .CI(DP_OP_102J5_124_3590_n1342), .CO(
        DP_OP_102J5_124_3590_n1329), .S(DP_OP_102J5_124_3590_n1330) );
  FADDX1_HVT DP_OP_102J5_124_3590_U780 ( .A(DP_OP_102J5_124_3590_n1344), .B(
        DP_OP_102J5_124_3590_n1350), .CI(DP_OP_102J5_124_3590_n1409), .CO(
        DP_OP_102J5_124_3590_n1327), .S(DP_OP_102J5_124_3590_n1328) );
  FADDX1_HVT DP_OP_102J5_124_3590_U779 ( .A(DP_OP_102J5_124_3590_n1348), .B(
        DP_OP_102J5_124_3590_n1346), .CI(DP_OP_102J5_124_3590_n1407), .CO(
        DP_OP_102J5_124_3590_n1325), .S(DP_OP_102J5_124_3590_n1326) );
  FADDX1_HVT DP_OP_102J5_124_3590_U778 ( .A(DP_OP_102J5_124_3590_n1338), .B(
        DP_OP_102J5_124_3590_n1336), .CI(DP_OP_102J5_124_3590_n1405), .CO(
        DP_OP_102J5_124_3590_n1323), .S(DP_OP_102J5_124_3590_n1324) );
  FADDX1_HVT DP_OP_102J5_124_3590_U777 ( .A(DP_OP_102J5_124_3590_n1403), .B(
        DP_OP_102J5_124_3590_n1334), .CI(DP_OP_102J5_124_3590_n1332), .CO(
        DP_OP_102J5_124_3590_n1321), .S(DP_OP_102J5_124_3590_n1322) );
  FADDX1_HVT DP_OP_102J5_124_3590_U776 ( .A(DP_OP_102J5_124_3590_n1330), .B(
        DP_OP_102J5_124_3590_n1328), .CI(DP_OP_102J5_124_3590_n1326), .CO(
        DP_OP_102J5_124_3590_n1319), .S(DP_OP_102J5_124_3590_n1320) );
  FADDX1_HVT DP_OP_102J5_124_3590_U775 ( .A(DP_OP_102J5_124_3590_n1401), .B(
        DP_OP_102J5_124_3590_n1324), .CI(DP_OP_102J5_124_3590_n1322), .CO(
        DP_OP_102J5_124_3590_n1317), .S(DP_OP_102J5_124_3590_n1318) );
  HADDX1_HVT DP_OP_102J5_124_3590_U774 ( .A0(DP_OP_102J5_124_3590_n1689), .B0(
        DP_OP_102J5_124_3590_n1513), .C1(DP_OP_102J5_124_3590_n1315), .SO(
        DP_OP_102J5_124_3590_n1316) );
  FADDX1_HVT DP_OP_102J5_124_3590_U773 ( .A(DP_OP_102J5_124_3590_n2172), .B(
        DP_OP_102J5_124_3590_n1820), .CI(DP_OP_102J5_124_3590_n1952), .CO(
        DP_OP_102J5_124_3590_n1313), .S(DP_OP_102J5_124_3590_n1314) );
  FADDX1_HVT DP_OP_102J5_124_3590_U772 ( .A(DP_OP_102J5_124_3590_n2084), .B(
        DP_OP_102J5_124_3590_n2040), .CI(DP_OP_102J5_124_3590_n2216), .CO(
        DP_OP_102J5_124_3590_n1311), .S(DP_OP_102J5_124_3590_n1312) );
  FADDX1_HVT DP_OP_102J5_124_3590_U771 ( .A(DP_OP_102J5_124_3590_n1864), .B(
        DP_OP_102J5_124_3590_n1996), .CI(DP_OP_102J5_124_3590_n1645), .CO(
        DP_OP_102J5_124_3590_n1309), .S(DP_OP_102J5_124_3590_n1310) );
  FADDX1_HVT DP_OP_102J5_124_3590_U770 ( .A(DP_OP_102J5_124_3590_n1601), .B(
        DP_OP_102J5_124_3590_n1908), .CI(DP_OP_102J5_124_3590_n2304), .CO(
        DP_OP_102J5_124_3590_n1307), .S(DP_OP_102J5_124_3590_n1308) );
  FADDX1_HVT DP_OP_102J5_124_3590_U769 ( .A(DP_OP_102J5_124_3590_n1777), .B(
        DP_OP_102J5_124_3590_n2128), .CI(DP_OP_102J5_124_3590_n2348), .CO(
        DP_OP_102J5_124_3590_n1305), .S(DP_OP_102J5_124_3590_n1306) );
  FADDX1_HVT DP_OP_102J5_124_3590_U768 ( .A(DP_OP_102J5_124_3590_n1557), .B(
        DP_OP_102J5_124_3590_n1733), .CI(DP_OP_102J5_124_3590_n2260), .CO(
        DP_OP_102J5_124_3590_n1303), .S(DP_OP_102J5_124_3590_n1304) );
  FADDX1_HVT DP_OP_102J5_124_3590_U767 ( .A(DP_OP_102J5_124_3590_n1534), .B(
        DP_OP_102J5_124_3590_n1520), .CI(DP_OP_102J5_124_3590_n1527), .CO(
        DP_OP_102J5_124_3590_n1301), .S(DP_OP_102J5_124_3590_n1302) );
  FADDX1_HVT DP_OP_102J5_124_3590_U766 ( .A(DP_OP_102J5_124_3590_n1571), .B(
        DP_OP_102J5_124_3590_n1564), .CI(DP_OP_102J5_124_3590_n1578), .CO(
        DP_OP_102J5_124_3590_n1299), .S(DP_OP_102J5_124_3590_n1300) );
  FADDX1_HVT DP_OP_102J5_124_3590_U765 ( .A(DP_OP_102J5_124_3590_n1615), .B(
        DP_OP_102J5_124_3590_n1608), .CI(DP_OP_102J5_124_3590_n1622), .CO(
        DP_OP_102J5_124_3590_n1297), .S(DP_OP_102J5_124_3590_n1298) );
  FADDX1_HVT DP_OP_102J5_124_3590_U764 ( .A(DP_OP_102J5_124_3590_n2368), .B(
        DP_OP_102J5_124_3590_n1652), .CI(DP_OP_102J5_124_3590_n2362), .CO(
        DP_OP_102J5_124_3590_n1295), .S(DP_OP_102J5_124_3590_n1296) );
  FADDX1_HVT DP_OP_102J5_124_3590_U763 ( .A(DP_OP_102J5_124_3590_n1966), .B(
        DP_OP_102J5_124_3590_n2355), .CI(DP_OP_102J5_124_3590_n1659), .CO(
        DP_OP_102J5_124_3590_n1293), .S(DP_OP_102J5_124_3590_n1294) );
  FADDX1_HVT DP_OP_102J5_124_3590_U762 ( .A(DP_OP_102J5_124_3590_n1959), .B(
        DP_OP_102J5_124_3590_n2325), .CI(DP_OP_102J5_124_3590_n2318), .CO(
        DP_OP_102J5_124_3590_n1291), .S(DP_OP_102J5_124_3590_n1292) );
  FADDX1_HVT DP_OP_102J5_124_3590_U761 ( .A(DP_OP_102J5_124_3590_n1922), .B(
        DP_OP_102J5_124_3590_n1666), .CI(DP_OP_102J5_124_3590_n2311), .CO(
        DP_OP_102J5_124_3590_n1289), .S(DP_OP_102J5_124_3590_n1290) );
  FADDX1_HVT DP_OP_102J5_124_3590_U760 ( .A(DP_OP_102J5_124_3590_n1929), .B(
        DP_OP_102J5_124_3590_n2281), .CI(DP_OP_102J5_124_3590_n1696), .CO(
        DP_OP_102J5_124_3590_n1287), .S(DP_OP_102J5_124_3590_n1288) );
  FADDX1_HVT DP_OP_102J5_124_3590_U759 ( .A(DP_OP_102J5_124_3590_n2274), .B(
        DP_OP_102J5_124_3590_n1703), .CI(DP_OP_102J5_124_3590_n2267), .CO(
        DP_OP_102J5_124_3590_n1285), .S(DP_OP_102J5_124_3590_n1286) );
  FADDX1_HVT DP_OP_102J5_124_3590_U758 ( .A(DP_OP_102J5_124_3590_n1885), .B(
        DP_OP_102J5_124_3590_n2237), .CI(DP_OP_102J5_124_3590_n1710), .CO(
        DP_OP_102J5_124_3590_n1283), .S(DP_OP_102J5_124_3590_n1284) );
  FADDX1_HVT DP_OP_102J5_124_3590_U757 ( .A(DP_OP_102J5_124_3590_n1915), .B(
        DP_OP_102J5_124_3590_n1740), .CI(DP_OP_102J5_124_3590_n2230), .CO(
        DP_OP_102J5_124_3590_n1281), .S(DP_OP_102J5_124_3590_n1282) );
  FADDX1_HVT DP_OP_102J5_124_3590_U756 ( .A(DP_OP_102J5_124_3590_n1878), .B(
        DP_OP_102J5_124_3590_n1747), .CI(DP_OP_102J5_124_3590_n2223), .CO(
        DP_OP_102J5_124_3590_n1279), .S(DP_OP_102J5_124_3590_n1280) );
  FADDX1_HVT DP_OP_102J5_124_3590_U755 ( .A(DP_OP_102J5_124_3590_n1973), .B(
        DP_OP_102J5_124_3590_n1754), .CI(DP_OP_102J5_124_3590_n2193), .CO(
        DP_OP_102J5_124_3590_n1277), .S(DP_OP_102J5_124_3590_n1278) );
  FADDX1_HVT DP_OP_102J5_124_3590_U754 ( .A(DP_OP_102J5_124_3590_n2186), .B(
        DP_OP_102J5_124_3590_n1784), .CI(DP_OP_102J5_124_3590_n1791), .CO(
        DP_OP_102J5_124_3590_n1275), .S(DP_OP_102J5_124_3590_n1276) );
  FADDX1_HVT DP_OP_102J5_124_3590_U753 ( .A(DP_OP_102J5_124_3590_n2010), .B(
        DP_OP_102J5_124_3590_n2179), .CI(DP_OP_102J5_124_3590_n2149), .CO(
        DP_OP_102J5_124_3590_n1273), .S(DP_OP_102J5_124_3590_n1274) );
  FADDX1_HVT DP_OP_102J5_124_3590_U752 ( .A(DP_OP_102J5_124_3590_n1841), .B(
        DP_OP_102J5_124_3590_n2142), .CI(DP_OP_102J5_124_3590_n2135), .CO(
        DP_OP_102J5_124_3590_n1271), .S(DP_OP_102J5_124_3590_n1272) );
  FADDX1_HVT DP_OP_102J5_124_3590_U751 ( .A(DP_OP_102J5_124_3590_n1827), .B(
        DP_OP_102J5_124_3590_n2105), .CI(DP_OP_102J5_124_3590_n2098), .CO(
        DP_OP_102J5_124_3590_n1269), .S(DP_OP_102J5_124_3590_n1270) );
  FADDX1_HVT DP_OP_102J5_124_3590_U750 ( .A(DP_OP_102J5_124_3590_n2017), .B(
        DP_OP_102J5_124_3590_n2091), .CI(DP_OP_102J5_124_3590_n1798), .CO(
        DP_OP_102J5_124_3590_n1267), .S(DP_OP_102J5_124_3590_n1268) );
  FADDX1_HVT DP_OP_102J5_124_3590_U749 ( .A(DP_OP_102J5_124_3590_n1871), .B(
        DP_OP_102J5_124_3590_n2061), .CI(DP_OP_102J5_124_3590_n2054), .CO(
        DP_OP_102J5_124_3590_n1265), .S(DP_OP_102J5_124_3590_n1266) );
  FADDX1_HVT DP_OP_102J5_124_3590_U748 ( .A(DP_OP_102J5_124_3590_n2047), .B(
        DP_OP_102J5_124_3590_n1834), .CI(DP_OP_102J5_124_3590_n2003), .CO(
        DP_OP_102J5_124_3590_n1263), .S(DP_OP_102J5_124_3590_n1264) );
  FADDX1_HVT DP_OP_102J5_124_3590_U747 ( .A(DP_OP_102J5_124_3590_n1399), .B(
        DP_OP_102J5_124_3590_n1316), .CI(DP_OP_102J5_124_3590_n1361), .CO(
        DP_OP_102J5_124_3590_n1261), .S(DP_OP_102J5_124_3590_n1262) );
  FADDX1_HVT DP_OP_102J5_124_3590_U746 ( .A(DP_OP_102J5_124_3590_n1383), .B(
        DP_OP_102J5_124_3590_n1363), .CI(DP_OP_102J5_124_3590_n1367), .CO(
        DP_OP_102J5_124_3590_n1259), .S(DP_OP_102J5_124_3590_n1260) );
  FADDX1_HVT DP_OP_102J5_124_3590_U745 ( .A(DP_OP_102J5_124_3590_n1381), .B(
        DP_OP_102J5_124_3590_n1369), .CI(DP_OP_102J5_124_3590_n1365), .CO(
        DP_OP_102J5_124_3590_n1257), .S(DP_OP_102J5_124_3590_n1258) );
  FADDX1_HVT DP_OP_102J5_124_3590_U744 ( .A(DP_OP_102J5_124_3590_n1385), .B(
        DP_OP_102J5_124_3590_n1371), .CI(DP_OP_102J5_124_3590_n1375), .CO(
        DP_OP_102J5_124_3590_n1255), .S(DP_OP_102J5_124_3590_n1256) );
  FADDX1_HVT DP_OP_102J5_124_3590_U743 ( .A(DP_OP_102J5_124_3590_n1379), .B(
        DP_OP_102J5_124_3590_n1373), .CI(DP_OP_102J5_124_3590_n1377), .CO(
        DP_OP_102J5_124_3590_n1253), .S(DP_OP_102J5_124_3590_n1254) );
  FADDX1_HVT DP_OP_102J5_124_3590_U742 ( .A(DP_OP_102J5_124_3590_n1389), .B(
        DP_OP_102J5_124_3590_n1391), .CI(DP_OP_102J5_124_3590_n1393), .CO(
        DP_OP_102J5_124_3590_n1251), .S(DP_OP_102J5_124_3590_n1252) );
  FADDX1_HVT DP_OP_102J5_124_3590_U741 ( .A(DP_OP_102J5_124_3590_n1395), .B(
        DP_OP_102J5_124_3590_n1397), .CI(DP_OP_102J5_124_3590_n1387), .CO(
        DP_OP_102J5_124_3590_n1249), .S(DP_OP_102J5_124_3590_n1250) );
  FADDX1_HVT DP_OP_102J5_124_3590_U740 ( .A(DP_OP_102J5_124_3590_n1308), .B(
        DP_OP_102J5_124_3590_n1310), .CI(DP_OP_102J5_124_3590_n1314), .CO(
        DP_OP_102J5_124_3590_n1247), .S(DP_OP_102J5_124_3590_n1248) );
  FADDX1_HVT DP_OP_102J5_124_3590_U739 ( .A(DP_OP_102J5_124_3590_n1312), .B(
        DP_OP_102J5_124_3590_n1304), .CI(DP_OP_102J5_124_3590_n1306), .CO(
        DP_OP_102J5_124_3590_n1245), .S(DP_OP_102J5_124_3590_n1246) );
  FADDX1_HVT DP_OP_102J5_124_3590_U738 ( .A(DP_OP_102J5_124_3590_n1268), .B(
        DP_OP_102J5_124_3590_n1296), .CI(DP_OP_102J5_124_3590_n1298), .CO(
        DP_OP_102J5_124_3590_n1243), .S(DP_OP_102J5_124_3590_n1244) );
  FADDX1_HVT DP_OP_102J5_124_3590_U737 ( .A(DP_OP_102J5_124_3590_n1266), .B(
        DP_OP_102J5_124_3590_n1290), .CI(DP_OP_102J5_124_3590_n1292), .CO(
        DP_OP_102J5_124_3590_n1241), .S(DP_OP_102J5_124_3590_n1242) );
  FADDX1_HVT DP_OP_102J5_124_3590_U736 ( .A(DP_OP_102J5_124_3590_n1288), .B(
        DP_OP_102J5_124_3590_n1294), .CI(DP_OP_102J5_124_3590_n1286), .CO(
        DP_OP_102J5_124_3590_n1239), .S(DP_OP_102J5_124_3590_n1240) );
  FADDX1_HVT DP_OP_102J5_124_3590_U735 ( .A(DP_OP_102J5_124_3590_n1264), .B(
        DP_OP_102J5_124_3590_n1302), .CI(DP_OP_102J5_124_3590_n1282), .CO(
        DP_OP_102J5_124_3590_n1237), .S(DP_OP_102J5_124_3590_n1238) );
  FADDX1_HVT DP_OP_102J5_124_3590_U734 ( .A(DP_OP_102J5_124_3590_n1284), .B(
        DP_OP_102J5_124_3590_n1270), .CI(DP_OP_102J5_124_3590_n1276), .CO(
        DP_OP_102J5_124_3590_n1235), .S(DP_OP_102J5_124_3590_n1236) );
  FADDX1_HVT DP_OP_102J5_124_3590_U733 ( .A(DP_OP_102J5_124_3590_n1278), .B(
        DP_OP_102J5_124_3590_n1300), .CI(DP_OP_102J5_124_3590_n1280), .CO(
        DP_OP_102J5_124_3590_n1233), .S(DP_OP_102J5_124_3590_n1234) );
  FADDX1_HVT DP_OP_102J5_124_3590_U732 ( .A(DP_OP_102J5_124_3590_n1272), .B(
        DP_OP_102J5_124_3590_n1274), .CI(DP_OP_102J5_124_3590_n1359), .CO(
        DP_OP_102J5_124_3590_n1231), .S(DP_OP_102J5_124_3590_n1232) );
  FADDX1_HVT DP_OP_102J5_124_3590_U731 ( .A(DP_OP_102J5_124_3590_n1351), .B(
        DP_OP_102J5_124_3590_n1353), .CI(DP_OP_102J5_124_3590_n1478), .CO(
        DP_OP_102J5_124_3590_n1229), .S(DP_OP_102J5_124_3590_n1230) );
  FADDX1_HVT DP_OP_102J5_124_3590_U730 ( .A(DP_OP_102J5_124_3590_n1357), .B(
        DP_OP_102J5_124_3590_n1355), .CI(DP_OP_102J5_124_3590_n1262), .CO(
        DP_OP_102J5_124_3590_n1227), .S(DP_OP_102J5_124_3590_n1228) );
  FADDX1_HVT DP_OP_102J5_124_3590_U729 ( .A(DP_OP_102J5_124_3590_n1252), .B(
        DP_OP_102J5_124_3590_n1250), .CI(DP_OP_102J5_124_3590_n1254), .CO(
        DP_OP_102J5_124_3590_n1225), .S(DP_OP_102J5_124_3590_n1226) );
  FADDX1_HVT DP_OP_102J5_124_3590_U728 ( .A(DP_OP_102J5_124_3590_n1256), .B(
        DP_OP_102J5_124_3590_n1258), .CI(DP_OP_102J5_124_3590_n1260), .CO(
        DP_OP_102J5_124_3590_n1223), .S(DP_OP_102J5_124_3590_n1224) );
  FADDX1_HVT DP_OP_102J5_124_3590_U727 ( .A(DP_OP_102J5_124_3590_n1349), .B(
        DP_OP_102J5_124_3590_n1339), .CI(DP_OP_102J5_124_3590_n1341), .CO(
        DP_OP_102J5_124_3590_n1221), .S(DP_OP_102J5_124_3590_n1222) );
  FADDX1_HVT DP_OP_102J5_124_3590_U726 ( .A(DP_OP_102J5_124_3590_n1343), .B(
        DP_OP_102J5_124_3590_n1347), .CI(DP_OP_102J5_124_3590_n1345), .CO(
        DP_OP_102J5_124_3590_n1219), .S(DP_OP_102J5_124_3590_n1220) );
  FADDX1_HVT DP_OP_102J5_124_3590_U725 ( .A(DP_OP_102J5_124_3590_n1246), .B(
        DP_OP_102J5_124_3590_n1248), .CI(DP_OP_102J5_124_3590_n1236), .CO(
        DP_OP_102J5_124_3590_n1217), .S(DP_OP_102J5_124_3590_n1218) );
  FADDX1_HVT DP_OP_102J5_124_3590_U724 ( .A(DP_OP_102J5_124_3590_n1242), .B(
        DP_OP_102J5_124_3590_n1244), .CI(DP_OP_102J5_124_3590_n1337), .CO(
        DP_OP_102J5_124_3590_n1215), .S(DP_OP_102J5_124_3590_n1216) );
  FADDX1_HVT DP_OP_102J5_124_3590_U723 ( .A(DP_OP_102J5_124_3590_n1240), .B(
        DP_OP_102J5_124_3590_n1238), .CI(DP_OP_102J5_124_3590_n1234), .CO(
        DP_OP_102J5_124_3590_n1213), .S(DP_OP_102J5_124_3590_n1214) );
  FADDX1_HVT DP_OP_102J5_124_3590_U722 ( .A(DP_OP_102J5_124_3590_n1232), .B(
        DP_OP_102J5_124_3590_n1335), .CI(DP_OP_102J5_124_3590_n1331), .CO(
        DP_OP_102J5_124_3590_n1211), .S(DP_OP_102J5_124_3590_n1212) );
  FADDX1_HVT DP_OP_102J5_124_3590_U721 ( .A(DP_OP_102J5_124_3590_n1333), .B(
        DP_OP_102J5_124_3590_n1230), .CI(DP_OP_102J5_124_3590_n1228), .CO(
        DP_OP_102J5_124_3590_n1209), .S(DP_OP_102J5_124_3590_n1210) );
  FADDX1_HVT DP_OP_102J5_124_3590_U720 ( .A(DP_OP_102J5_124_3590_n1329), .B(
        DP_OP_102J5_124_3590_n1327), .CI(DP_OP_102J5_124_3590_n1222), .CO(
        DP_OP_102J5_124_3590_n1207), .S(DP_OP_102J5_124_3590_n1208) );
  FADDX1_HVT DP_OP_102J5_124_3590_U719 ( .A(DP_OP_102J5_124_3590_n1224), .B(
        DP_OP_102J5_124_3590_n1226), .CI(DP_OP_102J5_124_3590_n1220), .CO(
        DP_OP_102J5_124_3590_n1205), .S(DP_OP_102J5_124_3590_n1206) );
  FADDX1_HVT DP_OP_102J5_124_3590_U718 ( .A(DP_OP_102J5_124_3590_n1218), .B(
        DP_OP_102J5_124_3590_n1325), .CI(DP_OP_102J5_124_3590_n1214), .CO(
        DP_OP_102J5_124_3590_n1203), .S(DP_OP_102J5_124_3590_n1204) );
  FADDX1_HVT DP_OP_102J5_124_3590_U717 ( .A(DP_OP_102J5_124_3590_n1216), .B(
        DP_OP_102J5_124_3590_n1323), .CI(DP_OP_102J5_124_3590_n1212), .CO(
        DP_OP_102J5_124_3590_n1201), .S(DP_OP_102J5_124_3590_n1202) );
  FADDX1_HVT DP_OP_102J5_124_3590_U716 ( .A(DP_OP_102J5_124_3590_n1321), .B(
        DP_OP_102J5_124_3590_n1210), .CI(DP_OP_102J5_124_3590_n1208), .CO(
        DP_OP_102J5_124_3590_n1199), .S(DP_OP_102J5_124_3590_n1200) );
  FADDX1_HVT DP_OP_102J5_124_3590_U715 ( .A(DP_OP_102J5_124_3590_n1206), .B(
        DP_OP_102J5_124_3590_n1319), .CI(DP_OP_102J5_124_3590_n1204), .CO(
        DP_OP_102J5_124_3590_n1197), .S(DP_OP_102J5_124_3590_n1198) );
  FADDX1_HVT DP_OP_102J5_124_3590_U714 ( .A(DP_OP_102J5_124_3590_n1202), .B(
        DP_OP_102J5_124_3590_n1317), .CI(DP_OP_102J5_124_3590_n1200), .CO(
        DP_OP_102J5_124_3590_n1195), .S(DP_OP_102J5_124_3590_n1196) );
  FADDX1_HVT DP_OP_102J5_124_3590_U713 ( .A(DP_OP_102J5_124_3590_n1688), .B(
        DP_OP_102J5_124_3590_n2039), .CI(DP_OP_102J5_124_3590_n1512), .CO(
        DP_OP_102J5_124_3590_n1193), .S(DP_OP_102J5_124_3590_n1194) );
  FADDX1_HVT DP_OP_102J5_124_3590_U712 ( .A(DP_OP_102J5_124_3590_n2171), .B(
        DP_OP_102J5_124_3590_n2215), .CI(DP_OP_102J5_124_3590_n1732), .CO(
        DP_OP_102J5_124_3590_n1191), .S(DP_OP_102J5_124_3590_n1192) );
  FADDX1_HVT DP_OP_102J5_124_3590_U711 ( .A(DP_OP_102J5_124_3590_n2303), .B(
        DP_OP_102J5_124_3590_n1819), .CI(DP_OP_102J5_124_3590_n1863), .CO(
        DP_OP_102J5_124_3590_n1189), .S(DP_OP_102J5_124_3590_n1190) );
  FADDX1_HVT DP_OP_102J5_124_3590_U710 ( .A(DP_OP_102J5_124_3590_n2347), .B(
        DP_OP_102J5_124_3590_n1907), .CI(DP_OP_102J5_124_3590_n1776), .CO(
        DP_OP_102J5_124_3590_n1187), .S(DP_OP_102J5_124_3590_n1188) );
  FADDX1_HVT DP_OP_102J5_124_3590_U709 ( .A(DP_OP_102J5_124_3590_n1995), .B(
        DP_OP_102J5_124_3590_n1600), .CI(DP_OP_102J5_124_3590_n2259), .CO(
        DP_OP_102J5_124_3590_n1185), .S(DP_OP_102J5_124_3590_n1186) );
  FADDX1_HVT DP_OP_102J5_124_3590_U708 ( .A(DP_OP_102J5_124_3590_n2127), .B(
        DP_OP_102J5_124_3590_n2083), .CI(DP_OP_102J5_124_3590_n1644), .CO(
        DP_OP_102J5_124_3590_n1183), .S(DP_OP_102J5_124_3590_n1184) );
  FADDX1_HVT DP_OP_102J5_124_3590_U707 ( .A(DP_OP_102J5_124_3590_n1951), .B(
        DP_OP_102J5_124_3590_n1556), .CI(DP_OP_102J5_124_3590_n1965), .CO(
        DP_OP_102J5_124_3590_n1181), .S(DP_OP_102J5_124_3590_n1182) );
  FADDX1_HVT DP_OP_102J5_124_3590_U706 ( .A(DP_OP_102J5_124_3590_n1958), .B(
        DP_OP_102J5_124_3590_n1526), .CI(DP_OP_102J5_124_3590_n1519), .CO(
        DP_OP_102J5_124_3590_n1179), .S(DP_OP_102J5_124_3590_n1180) );
  FADDX1_HVT DP_OP_102J5_124_3590_U705 ( .A(DP_OP_102J5_124_3590_n2367), .B(
        DP_OP_102J5_124_3590_n1533), .CI(DP_OP_102J5_124_3590_n1563), .CO(
        DP_OP_102J5_124_3590_n1177), .S(DP_OP_102J5_124_3590_n1178) );
  FADDX1_HVT DP_OP_102J5_124_3590_U704 ( .A(DP_OP_102J5_124_3590_n1877), .B(
        DP_OP_102J5_124_3590_n1570), .CI(DP_OP_102J5_124_3590_n2361), .CO(
        DP_OP_102J5_124_3590_n1175), .S(DP_OP_102J5_124_3590_n1176) );
  FADDX1_HVT DP_OP_102J5_124_3590_U703 ( .A(DP_OP_102J5_124_3590_n2354), .B(
        DP_OP_102J5_124_3590_n1577), .CI(DP_OP_102J5_124_3590_n1607), .CO(
        DP_OP_102J5_124_3590_n1173), .S(DP_OP_102J5_124_3590_n1174) );
  FADDX1_HVT DP_OP_102J5_124_3590_U702 ( .A(DP_OP_102J5_124_3590_n1870), .B(
        DP_OP_102J5_124_3590_n1614), .CI(DP_OP_102J5_124_3590_n2324), .CO(
        DP_OP_102J5_124_3590_n1171), .S(DP_OP_102J5_124_3590_n1172) );
  FADDX1_HVT DP_OP_102J5_124_3590_U701 ( .A(DP_OP_102J5_124_3590_n1884), .B(
        DP_OP_102J5_124_3590_n2317), .CI(DP_OP_102J5_124_3590_n1621), .CO(
        DP_OP_102J5_124_3590_n1169), .S(DP_OP_102J5_124_3590_n1170) );
  FADDX1_HVT DP_OP_102J5_124_3590_U700 ( .A(DP_OP_102J5_124_3590_n1914), .B(
        DP_OP_102J5_124_3590_n1651), .CI(DP_OP_102J5_124_3590_n2310), .CO(
        DP_OP_102J5_124_3590_n1167), .S(DP_OP_102J5_124_3590_n1168) );
  FADDX1_HVT DP_OP_102J5_124_3590_U699 ( .A(DP_OP_102J5_124_3590_n1840), .B(
        DP_OP_102J5_124_3590_n2280), .CI(DP_OP_102J5_124_3590_n2273), .CO(
        DP_OP_102J5_124_3590_n1165), .S(DP_OP_102J5_124_3590_n1166) );
  FADDX1_HVT DP_OP_102J5_124_3590_U698 ( .A(DP_OP_102J5_124_3590_n1826), .B(
        DP_OP_102J5_124_3590_n2266), .CI(DP_OP_102J5_124_3590_n2236), .CO(
        DP_OP_102J5_124_3590_n1163), .S(DP_OP_102J5_124_3590_n1164) );
  FADDX1_HVT DP_OP_102J5_124_3590_U697 ( .A(DP_OP_102J5_124_3590_n1797), .B(
        DP_OP_102J5_124_3590_n2229), .CI(DP_OP_102J5_124_3590_n2222), .CO(
        DP_OP_102J5_124_3590_n1161), .S(DP_OP_102J5_124_3590_n1162) );
  FADDX1_HVT DP_OP_102J5_124_3590_U696 ( .A(DP_OP_102J5_124_3590_n1783), .B(
        DP_OP_102J5_124_3590_n1658), .CI(DP_OP_102J5_124_3590_n1665), .CO(
        DP_OP_102J5_124_3590_n1159), .S(DP_OP_102J5_124_3590_n1160) );
  FADDX1_HVT DP_OP_102J5_124_3590_U695 ( .A(DP_OP_102J5_124_3590_n2192), .B(
        DP_OP_102J5_124_3590_n1695), .CI(DP_OP_102J5_124_3590_n1702), .CO(
        DP_OP_102J5_124_3590_n1157), .S(DP_OP_102J5_124_3590_n1158) );
  FADDX1_HVT DP_OP_102J5_124_3590_U694 ( .A(DP_OP_102J5_124_3590_n2185), .B(
        DP_OP_102J5_124_3590_n1709), .CI(DP_OP_102J5_124_3590_n1739), .CO(
        DP_OP_102J5_124_3590_n1155), .S(DP_OP_102J5_124_3590_n1156) );
  FADDX1_HVT DP_OP_102J5_124_3590_U693 ( .A(DP_OP_102J5_124_3590_n2178), .B(
        DP_OP_102J5_124_3590_n1746), .CI(DP_OP_102J5_124_3590_n1753), .CO(
        DP_OP_102J5_124_3590_n1153), .S(DP_OP_102J5_124_3590_n1154) );
  FADDX1_HVT DP_OP_102J5_124_3590_U692 ( .A(DP_OP_102J5_124_3590_n2148), .B(
        DP_OP_102J5_124_3590_n1790), .CI(DP_OP_102J5_124_3590_n1833), .CO(
        DP_OP_102J5_124_3590_n1151), .S(DP_OP_102J5_124_3590_n1152) );
  FADDX1_HVT DP_OP_102J5_124_3590_U691 ( .A(DP_OP_102J5_124_3590_n2141), .B(
        DP_OP_102J5_124_3590_n1921), .CI(DP_OP_102J5_124_3590_n1928), .CO(
        DP_OP_102J5_124_3590_n1149), .S(DP_OP_102J5_124_3590_n1150) );
  FADDX1_HVT DP_OP_102J5_124_3590_U690 ( .A(DP_OP_102J5_124_3590_n2134), .B(
        DP_OP_102J5_124_3590_n1972), .CI(DP_OP_102J5_124_3590_n2002), .CO(
        DP_OP_102J5_124_3590_n1147), .S(DP_OP_102J5_124_3590_n1148) );
  FADDX1_HVT DP_OP_102J5_124_3590_U689 ( .A(DP_OP_102J5_124_3590_n2046), .B(
        DP_OP_102J5_124_3590_n2009), .CI(DP_OP_102J5_124_3590_n2104), .CO(
        DP_OP_102J5_124_3590_n1145), .S(DP_OP_102J5_124_3590_n1146) );
  FADDX1_HVT DP_OP_102J5_124_3590_U688 ( .A(DP_OP_102J5_124_3590_n2097), .B(
        DP_OP_102J5_124_3590_n2090), .CI(DP_OP_102J5_124_3590_n2060), .CO(
        DP_OP_102J5_124_3590_n1143), .S(DP_OP_102J5_124_3590_n1144) );
  FADDX1_HVT DP_OP_102J5_124_3590_U687 ( .A(DP_OP_102J5_124_3590_n2053), .B(
        DP_OP_102J5_124_3590_n2016), .CI(DP_OP_102J5_124_3590_n1315), .CO(
        DP_OP_102J5_124_3590_n1141), .S(DP_OP_102J5_124_3590_n1142) );
  FADDX1_HVT DP_OP_102J5_124_3590_U686 ( .A(DP_OP_102J5_124_3590_n1307), .B(
        DP_OP_102J5_124_3590_n1303), .CI(DP_OP_102J5_124_3590_n1309), .CO(
        DP_OP_102J5_124_3590_n1139), .S(DP_OP_102J5_124_3590_n1140) );
  FADDX1_HVT DP_OP_102J5_124_3590_U685 ( .A(DP_OP_102J5_124_3590_n1313), .B(
        DP_OP_102J5_124_3590_n1305), .CI(DP_OP_102J5_124_3590_n1311), .CO(
        DP_OP_102J5_124_3590_n1137), .S(DP_OP_102J5_124_3590_n1138) );
  FADDX1_HVT DP_OP_102J5_124_3590_U684 ( .A(DP_OP_102J5_124_3590_n1263), .B(
        DP_OP_102J5_124_3590_n1265), .CI(DP_OP_102J5_124_3590_n1269), .CO(
        DP_OP_102J5_124_3590_n1135), .S(DP_OP_102J5_124_3590_n1136) );
  FADDX1_HVT DP_OP_102J5_124_3590_U683 ( .A(DP_OP_102J5_124_3590_n1285), .B(
        DP_OP_102J5_124_3590_n1267), .CI(DP_OP_102J5_124_3590_n1271), .CO(
        DP_OP_102J5_124_3590_n1133), .S(DP_OP_102J5_124_3590_n1134) );
  FADDX1_HVT DP_OP_102J5_124_3590_U682 ( .A(DP_OP_102J5_124_3590_n1287), .B(
        DP_OP_102J5_124_3590_n1273), .CI(DP_OP_102J5_124_3590_n1275), .CO(
        DP_OP_102J5_124_3590_n1131), .S(DP_OP_102J5_124_3590_n1132) );
  FADDX1_HVT DP_OP_102J5_124_3590_U681 ( .A(DP_OP_102J5_124_3590_n1289), .B(
        DP_OP_102J5_124_3590_n1277), .CI(DP_OP_102J5_124_3590_n1279), .CO(
        DP_OP_102J5_124_3590_n1129), .S(DP_OP_102J5_124_3590_n1130) );
  FADDX1_HVT DP_OP_102J5_124_3590_U680 ( .A(DP_OP_102J5_124_3590_n1281), .B(
        DP_OP_102J5_124_3590_n1283), .CI(DP_OP_102J5_124_3590_n1293), .CO(
        DP_OP_102J5_124_3590_n1127), .S(DP_OP_102J5_124_3590_n1128) );
  FADDX1_HVT DP_OP_102J5_124_3590_U679 ( .A(DP_OP_102J5_124_3590_n1297), .B(
        DP_OP_102J5_124_3590_n1291), .CI(DP_OP_102J5_124_3590_n1299), .CO(
        DP_OP_102J5_124_3590_n1125), .S(DP_OP_102J5_124_3590_n1126) );
  FADDX1_HVT DP_OP_102J5_124_3590_U678 ( .A(DP_OP_102J5_124_3590_n1301), .B(
        DP_OP_102J5_124_3590_n1295), .CI(DP_OP_102J5_124_3590_n1188), .CO(
        DP_OP_102J5_124_3590_n1123), .S(DP_OP_102J5_124_3590_n1124) );
  FADDX1_HVT DP_OP_102J5_124_3590_U677 ( .A(DP_OP_102J5_124_3590_n1184), .B(
        DP_OP_102J5_124_3590_n1186), .CI(DP_OP_102J5_124_3590_n1182), .CO(
        DP_OP_102J5_124_3590_n1121), .S(DP_OP_102J5_124_3590_n1122) );
  FADDX1_HVT DP_OP_102J5_124_3590_U676 ( .A(DP_OP_102J5_124_3590_n1192), .B(
        DP_OP_102J5_124_3590_n1190), .CI(DP_OP_102J5_124_3590_n1194), .CO(
        DP_OP_102J5_124_3590_n1119), .S(DP_OP_102J5_124_3590_n1120) );
  FADDX1_HVT DP_OP_102J5_124_3590_U675 ( .A(DP_OP_102J5_124_3590_n1174), .B(
        DP_OP_102J5_124_3590_n1180), .CI(DP_OP_102J5_124_3590_n1178), .CO(
        DP_OP_102J5_124_3590_n1117), .S(DP_OP_102J5_124_3590_n1118) );
  FADDX1_HVT DP_OP_102J5_124_3590_U674 ( .A(DP_OP_102J5_124_3590_n1170), .B(
        DP_OP_102J5_124_3590_n1176), .CI(DP_OP_102J5_124_3590_n1164), .CO(
        DP_OP_102J5_124_3590_n1115), .S(DP_OP_102J5_124_3590_n1116) );
  FADDX1_HVT DP_OP_102J5_124_3590_U673 ( .A(DP_OP_102J5_124_3590_n1162), .B(
        DP_OP_102J5_124_3590_n1158), .CI(DP_OP_102J5_124_3590_n1154), .CO(
        DP_OP_102J5_124_3590_n1113), .S(DP_OP_102J5_124_3590_n1114) );
  FADDX1_HVT DP_OP_102J5_124_3590_U672 ( .A(DP_OP_102J5_124_3590_n1166), .B(
        DP_OP_102J5_124_3590_n1148), .CI(DP_OP_102J5_124_3590_n1146), .CO(
        DP_OP_102J5_124_3590_n1111), .S(DP_OP_102J5_124_3590_n1112) );
  FADDX1_HVT DP_OP_102J5_124_3590_U671 ( .A(DP_OP_102J5_124_3590_n1160), .B(
        DP_OP_102J5_124_3590_n1150), .CI(DP_OP_102J5_124_3590_n1152), .CO(
        DP_OP_102J5_124_3590_n1109), .S(DP_OP_102J5_124_3590_n1110) );
  FADDX1_HVT DP_OP_102J5_124_3590_U670 ( .A(DP_OP_102J5_124_3590_n1156), .B(
        DP_OP_102J5_124_3590_n1172), .CI(DP_OP_102J5_124_3590_n1144), .CO(
        DP_OP_102J5_124_3590_n1107), .S(DP_OP_102J5_124_3590_n1108) );
  FADDX1_HVT DP_OP_102J5_124_3590_U669 ( .A(DP_OP_102J5_124_3590_n1168), .B(
        DP_OP_102J5_124_3590_n1142), .CI(DP_OP_102J5_124_3590_n1261), .CO(
        DP_OP_102J5_124_3590_n1105), .S(DP_OP_102J5_124_3590_n1106) );
  FADDX1_HVT DP_OP_102J5_124_3590_U668 ( .A(DP_OP_102J5_124_3590_n1249), .B(
        DP_OP_102J5_124_3590_n1253), .CI(DP_OP_102J5_124_3590_n1477), .CO(
        DP_OP_102J5_124_3590_n1103), .S(DP_OP_102J5_124_3590_n1104) );
  FADDX1_HVT DP_OP_102J5_124_3590_U667 ( .A(DP_OP_102J5_124_3590_n1259), .B(
        DP_OP_102J5_124_3590_n1257), .CI(DP_OP_102J5_124_3590_n1251), .CO(
        DP_OP_102J5_124_3590_n1101), .S(DP_OP_102J5_124_3590_n1102) );
  FADDX1_HVT DP_OP_102J5_124_3590_U666 ( .A(DP_OP_102J5_124_3590_n1255), .B(
        DP_OP_102J5_124_3590_n1245), .CI(DP_OP_102J5_124_3590_n1247), .CO(
        DP_OP_102J5_124_3590_n1099), .S(DP_OP_102J5_124_3590_n1100) );
  FADDX1_HVT DP_OP_102J5_124_3590_U665 ( .A(DP_OP_102J5_124_3590_n1138), .B(
        DP_OP_102J5_124_3590_n1140), .CI(DP_OP_102J5_124_3590_n1243), .CO(
        DP_OP_102J5_124_3590_n1097), .S(DP_OP_102J5_124_3590_n1098) );
  FADDX1_HVT DP_OP_102J5_124_3590_U664 ( .A(DP_OP_102J5_124_3590_n1132), .B(
        DP_OP_102J5_124_3590_n1241), .CI(DP_OP_102J5_124_3590_n1124), .CO(
        DP_OP_102J5_124_3590_n1095), .S(DP_OP_102J5_124_3590_n1096) );
  FADDX1_HVT DP_OP_102J5_124_3590_U663 ( .A(DP_OP_102J5_124_3590_n1239), .B(
        DP_OP_102J5_124_3590_n1126), .CI(DP_OP_102J5_124_3590_n1134), .CO(
        DP_OP_102J5_124_3590_n1093), .S(DP_OP_102J5_124_3590_n1094) );
  FADDX1_HVT DP_OP_102J5_124_3590_U662 ( .A(DP_OP_102J5_124_3590_n1237), .B(
        DP_OP_102J5_124_3590_n1128), .CI(DP_OP_102J5_124_3590_n1130), .CO(
        DP_OP_102J5_124_3590_n1091), .S(DP_OP_102J5_124_3590_n1092) );
  FADDX1_HVT DP_OP_102J5_124_3590_U661 ( .A(DP_OP_102J5_124_3590_n1235), .B(
        DP_OP_102J5_124_3590_n1136), .CI(DP_OP_102J5_124_3590_n1233), .CO(
        DP_OP_102J5_124_3590_n1089), .S(DP_OP_102J5_124_3590_n1090) );
  FADDX1_HVT DP_OP_102J5_124_3590_U660 ( .A(DP_OP_102J5_124_3590_n1231), .B(
        DP_OP_102J5_124_3590_n1122), .CI(DP_OP_102J5_124_3590_n1120), .CO(
        DP_OP_102J5_124_3590_n1087), .S(DP_OP_102J5_124_3590_n1088) );
  FADDX1_HVT DP_OP_102J5_124_3590_U659 ( .A(DP_OP_102J5_124_3590_n1114), .B(
        DP_OP_102J5_124_3590_n1110), .CI(DP_OP_102J5_124_3590_n1112), .CO(
        DP_OP_102J5_124_3590_n1085), .S(DP_OP_102J5_124_3590_n1086) );
  FADDX1_HVT DP_OP_102J5_124_3590_U658 ( .A(DP_OP_102J5_124_3590_n1108), .B(
        DP_OP_102J5_124_3590_n1118), .CI(DP_OP_102J5_124_3590_n1116), .CO(
        DP_OP_102J5_124_3590_n1083), .S(DP_OP_102J5_124_3590_n1084) );
  FADDX1_HVT DP_OP_102J5_124_3590_U657 ( .A(DP_OP_102J5_124_3590_n1229), .B(
        DP_OP_102J5_124_3590_n1106), .CI(DP_OP_102J5_124_3590_n1227), .CO(
        DP_OP_102J5_124_3590_n1081), .S(DP_OP_102J5_124_3590_n1082) );
  FADDX1_HVT DP_OP_102J5_124_3590_U656 ( .A(DP_OP_102J5_124_3590_n1225), .B(
        DP_OP_102J5_124_3590_n1102), .CI(DP_OP_102J5_124_3590_n1104), .CO(
        DP_OP_102J5_124_3590_n1079), .S(DP_OP_102J5_124_3590_n1080) );
  FADDX1_HVT DP_OP_102J5_124_3590_U655 ( .A(DP_OP_102J5_124_3590_n1223), .B(
        DP_OP_102J5_124_3590_n1219), .CI(DP_OP_102J5_124_3590_n1221), .CO(
        DP_OP_102J5_124_3590_n1077), .S(DP_OP_102J5_124_3590_n1078) );
  FADDX1_HVT DP_OP_102J5_124_3590_U654 ( .A(DP_OP_102J5_124_3590_n1100), .B(
        DP_OP_102J5_124_3590_n1217), .CI(DP_OP_102J5_124_3590_n1098), .CO(
        DP_OP_102J5_124_3590_n1075), .S(DP_OP_102J5_124_3590_n1076) );
  FADDX1_HVT DP_OP_102J5_124_3590_U653 ( .A(DP_OP_102J5_124_3590_n1213), .B(
        DP_OP_102J5_124_3590_n1092), .CI(DP_OP_102J5_124_3590_n1090), .CO(
        DP_OP_102J5_124_3590_n1073), .S(DP_OP_102J5_124_3590_n1074) );
  FADDX1_HVT DP_OP_102J5_124_3590_U652 ( .A(DP_OP_102J5_124_3590_n1215), .B(
        DP_OP_102J5_124_3590_n1096), .CI(DP_OP_102J5_124_3590_n1094), .CO(
        DP_OP_102J5_124_3590_n1071), .S(DP_OP_102J5_124_3590_n1072) );
  FADDX1_HVT DP_OP_102J5_124_3590_U651 ( .A(DP_OP_102J5_124_3590_n1088), .B(
        DP_OP_102J5_124_3590_n1086), .CI(DP_OP_102J5_124_3590_n1084), .CO(
        DP_OP_102J5_124_3590_n1069), .S(DP_OP_102J5_124_3590_n1070) );
  FADDX1_HVT DP_OP_102J5_124_3590_U650 ( .A(DP_OP_102J5_124_3590_n1211), .B(
        DP_OP_102J5_124_3590_n1209), .CI(DP_OP_102J5_124_3590_n1082), .CO(
        DP_OP_102J5_124_3590_n1067), .S(DP_OP_102J5_124_3590_n1068) );
  FADDX1_HVT DP_OP_102J5_124_3590_U649 ( .A(DP_OP_102J5_124_3590_n1207), .B(
        DP_OP_102J5_124_3590_n1205), .CI(DP_OP_102J5_124_3590_n1080), .CO(
        DP_OP_102J5_124_3590_n1065), .S(DP_OP_102J5_124_3590_n1066) );
  FADDX1_HVT DP_OP_102J5_124_3590_U648 ( .A(DP_OP_102J5_124_3590_n1078), .B(
        DP_OP_102J5_124_3590_n1076), .CI(DP_OP_102J5_124_3590_n1203), .CO(
        DP_OP_102J5_124_3590_n1063), .S(DP_OP_102J5_124_3590_n1064) );
  FADDX1_HVT DP_OP_102J5_124_3590_U647 ( .A(DP_OP_102J5_124_3590_n1074), .B(
        DP_OP_102J5_124_3590_n1072), .CI(DP_OP_102J5_124_3590_n1201), .CO(
        DP_OP_102J5_124_3590_n1061), .S(DP_OP_102J5_124_3590_n1062) );
  FADDX1_HVT DP_OP_102J5_124_3590_U646 ( .A(DP_OP_102J5_124_3590_n1070), .B(
        DP_OP_102J5_124_3590_n1068), .CI(DP_OP_102J5_124_3590_n1199), .CO(
        DP_OP_102J5_124_3590_n1059), .S(DP_OP_102J5_124_3590_n1060) );
  FADDX1_HVT DP_OP_102J5_124_3590_U645 ( .A(DP_OP_102J5_124_3590_n1066), .B(
        DP_OP_102J5_124_3590_n1197), .CI(DP_OP_102J5_124_3590_n1064), .CO(
        DP_OP_102J5_124_3590_n1057), .S(DP_OP_102J5_124_3590_n1058) );
  FADDX1_HVT DP_OP_102J5_124_3590_U644 ( .A(DP_OP_102J5_124_3590_n1062), .B(
        DP_OP_102J5_124_3590_n1195), .CI(DP_OP_102J5_124_3590_n1060), .CO(
        DP_OP_102J5_124_3590_n1055), .S(DP_OP_102J5_124_3590_n1056) );
  OR2X1_HVT DP_OP_102J5_124_3590_U643 ( .A1(DP_OP_102J5_124_3590_n2082), .A2(
        DP_OP_102J5_124_3590_n1950), .Y(DP_OP_102J5_124_3590_n1053) );
  FADDX1_HVT DP_OP_102J5_124_3590_U641 ( .A(DP_OP_102J5_124_3590_n2170), .B(
        DP_OP_102J5_124_3590_n1994), .CI(DP_OP_102J5_124_3590_n1511), .CO(
        DP_OP_102J5_124_3590_n1051), .S(DP_OP_102J5_124_3590_n1052) );
  FADDX1_HVT DP_OP_102J5_124_3590_U640 ( .A(DP_OP_102J5_124_3590_n1687), .B(
        DP_OP_102J5_124_3590_n1906), .CI(DP_OP_102J5_124_3590_n2038), .CO(
        DP_OP_102J5_124_3590_n1049), .S(DP_OP_102J5_124_3590_n1050) );
  FADDX1_HVT DP_OP_102J5_124_3590_U639 ( .A(DP_OP_102J5_124_3590_n1555), .B(
        DP_OP_102J5_124_3590_n2258), .CI(DP_OP_102J5_124_3590_n1862), .CO(
        DP_OP_102J5_124_3590_n1047), .S(DP_OP_102J5_124_3590_n1048) );
  FADDX1_HVT DP_OP_102J5_124_3590_U638 ( .A(DP_OP_102J5_124_3590_n2214), .B(
        DP_OP_102J5_124_3590_n2302), .CI(DP_OP_102J5_124_3590_n1643), .CO(
        DP_OP_102J5_124_3590_n1045), .S(DP_OP_102J5_124_3590_n1046) );
  FADDX1_HVT DP_OP_102J5_124_3590_U637 ( .A(DP_OP_102J5_124_3590_n1775), .B(
        DP_OP_102J5_124_3590_n1818), .CI(DP_OP_102J5_124_3590_n2346), .CO(
        DP_OP_102J5_124_3590_n1043), .S(DP_OP_102J5_124_3590_n1044) );
  FADDX1_HVT DP_OP_102J5_124_3590_U636 ( .A(DP_OP_102J5_124_3590_n1599), .B(
        DP_OP_102J5_124_3590_n1731), .CI(DP_OP_102J5_124_3590_n2126), .CO(
        DP_OP_102J5_124_3590_n1041), .S(DP_OP_102J5_124_3590_n1042) );
  FADDX1_HVT DP_OP_102J5_124_3590_U635 ( .A(DP_OP_102J5_124_3590_n1869), .B(
        DP_OP_102J5_124_3590_n1518), .CI(DP_OP_102J5_124_3590_n1525), .CO(
        DP_OP_102J5_124_3590_n1039), .S(DP_OP_102J5_124_3590_n1040) );
  FADDX1_HVT DP_OP_102J5_124_3590_U634 ( .A(DP_OP_102J5_124_3590_n1883), .B(
        DP_OP_102J5_124_3590_n2366), .CI(DP_OP_102J5_124_3590_n2360), .CO(
        DP_OP_102J5_124_3590_n1037), .S(DP_OP_102J5_124_3590_n1038) );
  FADDX1_HVT DP_OP_102J5_124_3590_U633 ( .A(DP_OP_102J5_124_3590_n1839), .B(
        DP_OP_102J5_124_3590_n2353), .CI(DP_OP_102J5_124_3590_n2323), .CO(
        DP_OP_102J5_124_3590_n1035), .S(DP_OP_102J5_124_3590_n1036) );
  FADDX1_HVT DP_OP_102J5_124_3590_U632 ( .A(DP_OP_102J5_124_3590_n1832), .B(
        DP_OP_102J5_124_3590_n1532), .CI(DP_OP_102J5_124_3590_n2316), .CO(
        DP_OP_102J5_124_3590_n1033), .S(DP_OP_102J5_124_3590_n1034) );
  FADDX1_HVT DP_OP_102J5_124_3590_U631 ( .A(DP_OP_102J5_124_3590_n1825), .B(
        DP_OP_102J5_124_3590_n2309), .CI(DP_OP_102J5_124_3590_n2279), .CO(
        DP_OP_102J5_124_3590_n1031), .S(DP_OP_102J5_124_3590_n1032) );
  FADDX1_HVT DP_OP_102J5_124_3590_U630 ( .A(DP_OP_102J5_124_3590_n1789), .B(
        DP_OP_102J5_124_3590_n2272), .CI(DP_OP_102J5_124_3590_n1562), .CO(
        DP_OP_102J5_124_3590_n1029), .S(DP_OP_102J5_124_3590_n1030) );
  FADDX1_HVT DP_OP_102J5_124_3590_U629 ( .A(DP_OP_102J5_124_3590_n1796), .B(
        DP_OP_102J5_124_3590_n1569), .CI(DP_OP_102J5_124_3590_n1576), .CO(
        DP_OP_102J5_124_3590_n1027), .S(DP_OP_102J5_124_3590_n1028) );
  FADDX1_HVT DP_OP_102J5_124_3590_U628 ( .A(DP_OP_102J5_124_3590_n1876), .B(
        DP_OP_102J5_124_3590_n1606), .CI(DP_OP_102J5_124_3590_n1613), .CO(
        DP_OP_102J5_124_3590_n1025), .S(DP_OP_102J5_124_3590_n1026) );
  FADDX1_HVT DP_OP_102J5_124_3590_U627 ( .A(DP_OP_102J5_124_3590_n1913), .B(
        DP_OP_102J5_124_3590_n1620), .CI(DP_OP_102J5_124_3590_n2265), .CO(
        DP_OP_102J5_124_3590_n1023), .S(DP_OP_102J5_124_3590_n1024) );
  FADDX1_HVT DP_OP_102J5_124_3590_U626 ( .A(DP_OP_102J5_124_3590_n1708), .B(
        DP_OP_102J5_124_3590_n2235), .CI(DP_OP_102J5_124_3590_n1650), .CO(
        DP_OP_102J5_124_3590_n1021), .S(DP_OP_102J5_124_3590_n1022) );
  FADDX1_HVT DP_OP_102J5_124_3590_U625 ( .A(DP_OP_102J5_124_3590_n2228), .B(
        DP_OP_102J5_124_3590_n1657), .CI(DP_OP_102J5_124_3590_n1664), .CO(
        DP_OP_102J5_124_3590_n1019), .S(DP_OP_102J5_124_3590_n1020) );
  FADDX1_HVT DP_OP_102J5_124_3590_U624 ( .A(DP_OP_102J5_124_3590_n2221), .B(
        DP_OP_102J5_124_3590_n1694), .CI(DP_OP_102J5_124_3590_n1701), .CO(
        DP_OP_102J5_124_3590_n1017), .S(DP_OP_102J5_124_3590_n1018) );
  FADDX1_HVT DP_OP_102J5_124_3590_U623 ( .A(DP_OP_102J5_124_3590_n2191), .B(
        DP_OP_102J5_124_3590_n1738), .CI(DP_OP_102J5_124_3590_n1745), .CO(
        DP_OP_102J5_124_3590_n1015), .S(DP_OP_102J5_124_3590_n1016) );
  FADDX1_HVT DP_OP_102J5_124_3590_U622 ( .A(DP_OP_102J5_124_3590_n2184), .B(
        DP_OP_102J5_124_3590_n1752), .CI(DP_OP_102J5_124_3590_n1782), .CO(
        DP_OP_102J5_124_3590_n1013), .S(DP_OP_102J5_124_3590_n1014) );
  FADDX1_HVT DP_OP_102J5_124_3590_U621 ( .A(DP_OP_102J5_124_3590_n2177), .B(
        DP_OP_102J5_124_3590_n1920), .CI(DP_OP_102J5_124_3590_n1927), .CO(
        DP_OP_102J5_124_3590_n1011), .S(DP_OP_102J5_124_3590_n1012) );
  FADDX1_HVT DP_OP_102J5_124_3590_U620 ( .A(DP_OP_102J5_124_3590_n2147), .B(
        DP_OP_102J5_124_3590_n1957), .CI(DP_OP_102J5_124_3590_n1964), .CO(
        DP_OP_102J5_124_3590_n1009), .S(DP_OP_102J5_124_3590_n1010) );
  FADDX1_HVT DP_OP_102J5_124_3590_U619 ( .A(DP_OP_102J5_124_3590_n2140), .B(
        DP_OP_102J5_124_3590_n1971), .CI(DP_OP_102J5_124_3590_n2001), .CO(
        DP_OP_102J5_124_3590_n1007), .S(DP_OP_102J5_124_3590_n1008) );
  FADDX1_HVT DP_OP_102J5_124_3590_U618 ( .A(DP_OP_102J5_124_3590_n2133), .B(
        DP_OP_102J5_124_3590_n2008), .CI(DP_OP_102J5_124_3590_n2015), .CO(
        DP_OP_102J5_124_3590_n1005), .S(DP_OP_102J5_124_3590_n1006) );
  FADDX1_HVT DP_OP_102J5_124_3590_U617 ( .A(DP_OP_102J5_124_3590_n2045), .B(
        DP_OP_102J5_124_3590_n2103), .CI(DP_OP_102J5_124_3590_n2096), .CO(
        DP_OP_102J5_124_3590_n1003), .S(DP_OP_102J5_124_3590_n1004) );
  FADDX1_HVT DP_OP_102J5_124_3590_U616 ( .A(DP_OP_102J5_124_3590_n2059), .B(
        DP_OP_102J5_124_3590_n2089), .CI(DP_OP_102J5_124_3590_n2052), .CO(
        DP_OP_102J5_124_3590_n1001), .S(DP_OP_102J5_124_3590_n1002) );
  FADDX1_HVT DP_OP_102J5_124_3590_U615 ( .A(DP_OP_102J5_124_3590_n1187), .B(
        DP_OP_102J5_124_3590_n1181), .CI(DP_OP_102J5_124_3590_n1054), .CO(
        DP_OP_102J5_124_3590_n999), .S(DP_OP_102J5_124_3590_n1000) );
  FADDX1_HVT DP_OP_102J5_124_3590_U614 ( .A(DP_OP_102J5_124_3590_n1185), .B(
        DP_OP_102J5_124_3590_n1189), .CI(DP_OP_102J5_124_3590_n1183), .CO(
        DP_OP_102J5_124_3590_n997), .S(DP_OP_102J5_124_3590_n998) );
  FADDX1_HVT DP_OP_102J5_124_3590_U613 ( .A(DP_OP_102J5_124_3590_n1193), .B(
        DP_OP_102J5_124_3590_n1191), .CI(DP_OP_102J5_124_3590_n1163), .CO(
        DP_OP_102J5_124_3590_n995), .S(DP_OP_102J5_124_3590_n996) );
  FADDX1_HVT DP_OP_102J5_124_3590_U612 ( .A(DP_OP_102J5_124_3590_n1161), .B(
        DP_OP_102J5_124_3590_n1145), .CI(DP_OP_102J5_124_3590_n1143), .CO(
        DP_OP_102J5_124_3590_n993), .S(DP_OP_102J5_124_3590_n994) );
  FADDX1_HVT DP_OP_102J5_124_3590_U611 ( .A(DP_OP_102J5_124_3590_n1159), .B(
        DP_OP_102J5_124_3590_n1149), .CI(DP_OP_102J5_124_3590_n1147), .CO(
        DP_OP_102J5_124_3590_n991), .S(DP_OP_102J5_124_3590_n992) );
  FADDX1_HVT DP_OP_102J5_124_3590_U610 ( .A(DP_OP_102J5_124_3590_n1157), .B(
        DP_OP_102J5_124_3590_n1153), .CI(DP_OP_102J5_124_3590_n1151), .CO(
        DP_OP_102J5_124_3590_n989), .S(DP_OP_102J5_124_3590_n990) );
  FADDX1_HVT DP_OP_102J5_124_3590_U609 ( .A(DP_OP_102J5_124_3590_n1155), .B(
        DP_OP_102J5_124_3590_n1167), .CI(DP_OP_102J5_124_3590_n1165), .CO(
        DP_OP_102J5_124_3590_n987), .S(DP_OP_102J5_124_3590_n988) );
  FADDX1_HVT DP_OP_102J5_124_3590_U608 ( .A(DP_OP_102J5_124_3590_n1175), .B(
        DP_OP_102J5_124_3590_n1169), .CI(DP_OP_102J5_124_3590_n1171), .CO(
        DP_OP_102J5_124_3590_n985), .S(DP_OP_102J5_124_3590_n986) );
  FADDX1_HVT DP_OP_102J5_124_3590_U607 ( .A(DP_OP_102J5_124_3590_n1173), .B(
        DP_OP_102J5_124_3590_n1177), .CI(DP_OP_102J5_124_3590_n1179), .CO(
        DP_OP_102J5_124_3590_n983), .S(DP_OP_102J5_124_3590_n984) );
  FADDX1_HVT DP_OP_102J5_124_3590_U606 ( .A(DP_OP_102J5_124_3590_n1141), .B(
        DP_OP_102J5_124_3590_n1042), .CI(DP_OP_102J5_124_3590_n1044), .CO(
        DP_OP_102J5_124_3590_n981), .S(DP_OP_102J5_124_3590_n982) );
  FADDX1_HVT DP_OP_102J5_124_3590_U605 ( .A(DP_OP_102J5_124_3590_n1046), .B(
        DP_OP_102J5_124_3590_n1052), .CI(DP_OP_102J5_124_3590_n1050), .CO(
        DP_OP_102J5_124_3590_n979), .S(DP_OP_102J5_124_3590_n980) );
  FADDX1_HVT DP_OP_102J5_124_3590_U604 ( .A(DP_OP_102J5_124_3590_n1048), .B(
        DP_OP_102J5_124_3590_n1008), .CI(DP_OP_102J5_124_3590_n1006), .CO(
        DP_OP_102J5_124_3590_n977), .S(DP_OP_102J5_124_3590_n978) );
  FADDX1_HVT DP_OP_102J5_124_3590_U603 ( .A(DP_OP_102J5_124_3590_n1002), .B(
        DP_OP_102J5_124_3590_n1040), .CI(DP_OP_102J5_124_3590_n1038), .CO(
        DP_OP_102J5_124_3590_n975), .S(DP_OP_102J5_124_3590_n976) );
  FADDX1_HVT DP_OP_102J5_124_3590_U602 ( .A(DP_OP_102J5_124_3590_n1030), .B(
        DP_OP_102J5_124_3590_n1028), .CI(DP_OP_102J5_124_3590_n1024), .CO(
        DP_OP_102J5_124_3590_n973), .S(DP_OP_102J5_124_3590_n974) );
  FADDX1_HVT DP_OP_102J5_124_3590_U601 ( .A(DP_OP_102J5_124_3590_n1032), .B(
        DP_OP_102J5_124_3590_n1020), .CI(DP_OP_102J5_124_3590_n1018), .CO(
        DP_OP_102J5_124_3590_n971), .S(DP_OP_102J5_124_3590_n972) );
  FADDX1_HVT DP_OP_102J5_124_3590_U600 ( .A(DP_OP_102J5_124_3590_n1022), .B(
        DP_OP_102J5_124_3590_n1004), .CI(DP_OP_102J5_124_3590_n1010), .CO(
        DP_OP_102J5_124_3590_n969), .S(DP_OP_102J5_124_3590_n970) );
  FADDX1_HVT DP_OP_102J5_124_3590_U599 ( .A(DP_OP_102J5_124_3590_n1026), .B(
        DP_OP_102J5_124_3590_n1012), .CI(DP_OP_102J5_124_3590_n1014), .CO(
        DP_OP_102J5_124_3590_n967), .S(DP_OP_102J5_124_3590_n968) );
  FADDX1_HVT DP_OP_102J5_124_3590_U598 ( .A(DP_OP_102J5_124_3590_n1016), .B(
        DP_OP_102J5_124_3590_n1034), .CI(DP_OP_102J5_124_3590_n1036), .CO(
        DP_OP_102J5_124_3590_n965), .S(DP_OP_102J5_124_3590_n966) );
  FADDX1_HVT DP_OP_102J5_124_3590_U597 ( .A(DP_OP_102J5_124_3590_n1137), .B(
        DP_OP_102J5_124_3590_n1139), .CI(DP_OP_102J5_124_3590_n1127), .CO(
        DP_OP_102J5_124_3590_n963), .S(DP_OP_102J5_124_3590_n964) );
  FADDX1_HVT DP_OP_102J5_124_3590_U596 ( .A(DP_OP_102J5_124_3590_n1125), .B(
        DP_OP_102J5_124_3590_n1131), .CI(DP_OP_102J5_124_3590_n1476), .CO(
        DP_OP_102J5_124_3590_n961), .S(DP_OP_102J5_124_3590_n962) );
  FADDX1_HVT DP_OP_102J5_124_3590_U595 ( .A(DP_OP_102J5_124_3590_n1129), .B(
        DP_OP_102J5_124_3590_n1135), .CI(DP_OP_102J5_124_3590_n1123), .CO(
        DP_OP_102J5_124_3590_n959), .S(DP_OP_102J5_124_3590_n960) );
  FADDX1_HVT DP_OP_102J5_124_3590_U594 ( .A(DP_OP_102J5_124_3590_n1133), .B(
        DP_OP_102J5_124_3590_n1121), .CI(DP_OP_102J5_124_3590_n1119), .CO(
        DP_OP_102J5_124_3590_n957), .S(DP_OP_102J5_124_3590_n958) );
  FADDX1_HVT DP_OP_102J5_124_3590_U593 ( .A(DP_OP_102J5_124_3590_n998), .B(
        DP_OP_102J5_124_3590_n1000), .CI(DP_OP_102J5_124_3590_n996), .CO(
        DP_OP_102J5_124_3590_n955), .S(DP_OP_102J5_124_3590_n956) );
  FADDX1_HVT DP_OP_102J5_124_3590_U592 ( .A(DP_OP_102J5_124_3590_n1117), .B(
        DP_OP_102J5_124_3590_n984), .CI(DP_OP_102J5_124_3590_n986), .CO(
        DP_OP_102J5_124_3590_n953), .S(DP_OP_102J5_124_3590_n954) );
  FADDX1_HVT DP_OP_102J5_124_3590_U591 ( .A(DP_OP_102J5_124_3590_n990), .B(
        DP_OP_102J5_124_3590_n994), .CI(DP_OP_102J5_124_3590_n992), .CO(
        DP_OP_102J5_124_3590_n951), .S(DP_OP_102J5_124_3590_n952) );
  FADDX1_HVT DP_OP_102J5_124_3590_U590 ( .A(DP_OP_102J5_124_3590_n1115), .B(
        DP_OP_102J5_124_3590_n988), .CI(DP_OP_102J5_124_3590_n1107), .CO(
        DP_OP_102J5_124_3590_n949), .S(DP_OP_102J5_124_3590_n950) );
  FADDX1_HVT DP_OP_102J5_124_3590_U589 ( .A(DP_OP_102J5_124_3590_n1113), .B(
        DP_OP_102J5_124_3590_n1109), .CI(DP_OP_102J5_124_3590_n1111), .CO(
        DP_OP_102J5_124_3590_n947), .S(DP_OP_102J5_124_3590_n948) );
  FADDX1_HVT DP_OP_102J5_124_3590_U588 ( .A(DP_OP_102J5_124_3590_n982), .B(
        DP_OP_102J5_124_3590_n980), .CI(DP_OP_102J5_124_3590_n978), .CO(
        DP_OP_102J5_124_3590_n945), .S(DP_OP_102J5_124_3590_n946) );
  FADDX1_HVT DP_OP_102J5_124_3590_U587 ( .A(DP_OP_102J5_124_3590_n1105), .B(
        DP_OP_102J5_124_3590_n972), .CI(DP_OP_102J5_124_3590_n974), .CO(
        DP_OP_102J5_124_3590_n943), .S(DP_OP_102J5_124_3590_n944) );
  FADDX1_HVT DP_OP_102J5_124_3590_U586 ( .A(DP_OP_102J5_124_3590_n970), .B(
        DP_OP_102J5_124_3590_n976), .CI(DP_OP_102J5_124_3590_n968), .CO(
        DP_OP_102J5_124_3590_n941), .S(DP_OP_102J5_124_3590_n942) );
  FADDX1_HVT DP_OP_102J5_124_3590_U585 ( .A(DP_OP_102J5_124_3590_n966), .B(
        DP_OP_102J5_124_3590_n1103), .CI(DP_OP_102J5_124_3590_n1101), .CO(
        DP_OP_102J5_124_3590_n939), .S(DP_OP_102J5_124_3590_n940) );
  FADDX1_HVT DP_OP_102J5_124_3590_U584 ( .A(DP_OP_102J5_124_3590_n1099), .B(
        DP_OP_102J5_124_3590_n1097), .CI(DP_OP_102J5_124_3590_n964), .CO(
        DP_OP_102J5_124_3590_n937), .S(DP_OP_102J5_124_3590_n938) );
  FADDX1_HVT DP_OP_102J5_124_3590_U583 ( .A(DP_OP_102J5_124_3590_n1095), .B(
        DP_OP_102J5_124_3590_n962), .CI(DP_OP_102J5_124_3590_n960), .CO(
        DP_OP_102J5_124_3590_n935), .S(DP_OP_102J5_124_3590_n936) );
  FADDX1_HVT DP_OP_102J5_124_3590_U582 ( .A(DP_OP_102J5_124_3590_n1093), .B(
        DP_OP_102J5_124_3590_n1089), .CI(DP_OP_102J5_124_3590_n1091), .CO(
        DP_OP_102J5_124_3590_n933), .S(DP_OP_102J5_124_3590_n934) );
  FADDX1_HVT DP_OP_102J5_124_3590_U581 ( .A(DP_OP_102J5_124_3590_n958), .B(
        DP_OP_102J5_124_3590_n1087), .CI(DP_OP_102J5_124_3590_n956), .CO(
        DP_OP_102J5_124_3590_n931), .S(DP_OP_102J5_124_3590_n932) );
  FADDX1_HVT DP_OP_102J5_124_3590_U580 ( .A(DP_OP_102J5_124_3590_n1085), .B(
        DP_OP_102J5_124_3590_n952), .CI(DP_OP_102J5_124_3590_n954), .CO(
        DP_OP_102J5_124_3590_n929), .S(DP_OP_102J5_124_3590_n930) );
  FADDX1_HVT DP_OP_102J5_124_3590_U579 ( .A(DP_OP_102J5_124_3590_n1083), .B(
        DP_OP_102J5_124_3590_n948), .CI(DP_OP_102J5_124_3590_n950), .CO(
        DP_OP_102J5_124_3590_n927), .S(DP_OP_102J5_124_3590_n928) );
  FADDX1_HVT DP_OP_102J5_124_3590_U578 ( .A(DP_OP_102J5_124_3590_n1081), .B(
        DP_OP_102J5_124_3590_n946), .CI(DP_OP_102J5_124_3590_n944), .CO(
        DP_OP_102J5_124_3590_n925), .S(DP_OP_102J5_124_3590_n926) );
  FADDX1_HVT DP_OP_102J5_124_3590_U577 ( .A(DP_OP_102J5_124_3590_n942), .B(
        DP_OP_102J5_124_3590_n940), .CI(DP_OP_102J5_124_3590_n1079), .CO(
        DP_OP_102J5_124_3590_n923), .S(DP_OP_102J5_124_3590_n924) );
  FADDX1_HVT DP_OP_102J5_124_3590_U576 ( .A(DP_OP_102J5_124_3590_n1077), .B(
        DP_OP_102J5_124_3590_n1075), .CI(DP_OP_102J5_124_3590_n938), .CO(
        DP_OP_102J5_124_3590_n921), .S(DP_OP_102J5_124_3590_n922) );
  FADDX1_HVT DP_OP_102J5_124_3590_U575 ( .A(DP_OP_102J5_124_3590_n1073), .B(
        DP_OP_102J5_124_3590_n934), .CI(DP_OP_102J5_124_3590_n936), .CO(
        DP_OP_102J5_124_3590_n919), .S(DP_OP_102J5_124_3590_n920) );
  FADDX1_HVT DP_OP_102J5_124_3590_U574 ( .A(DP_OP_102J5_124_3590_n1071), .B(
        DP_OP_102J5_124_3590_n932), .CI(DP_OP_102J5_124_3590_n1069), .CO(
        DP_OP_102J5_124_3590_n917), .S(DP_OP_102J5_124_3590_n918) );
  FADDX1_HVT DP_OP_102J5_124_3590_U573 ( .A(DP_OP_102J5_124_3590_n930), .B(
        DP_OP_102J5_124_3590_n928), .CI(DP_OP_102J5_124_3590_n1067), .CO(
        DP_OP_102J5_124_3590_n915), .S(DP_OP_102J5_124_3590_n916) );
  FADDX1_HVT DP_OP_102J5_124_3590_U572 ( .A(DP_OP_102J5_124_3590_n926), .B(
        DP_OP_102J5_124_3590_n924), .CI(DP_OP_102J5_124_3590_n1065), .CO(
        DP_OP_102J5_124_3590_n913), .S(DP_OP_102J5_124_3590_n914) );
  FADDX1_HVT DP_OP_102J5_124_3590_U571 ( .A(DP_OP_102J5_124_3590_n1063), .B(
        DP_OP_102J5_124_3590_n922), .CI(DP_OP_102J5_124_3590_n920), .CO(
        DP_OP_102J5_124_3590_n911), .S(DP_OP_102J5_124_3590_n912) );
  FADDX1_HVT DP_OP_102J5_124_3590_U570 ( .A(DP_OP_102J5_124_3590_n1061), .B(
        DP_OP_102J5_124_3590_n918), .CI(DP_OP_102J5_124_3590_n916), .CO(
        DP_OP_102J5_124_3590_n909), .S(DP_OP_102J5_124_3590_n910) );
  FADDX1_HVT DP_OP_102J5_124_3590_U569 ( .A(DP_OP_102J5_124_3590_n1059), .B(
        DP_OP_102J5_124_3590_n914), .CI(DP_OP_102J5_124_3590_n1057), .CO(
        DP_OP_102J5_124_3590_n907), .S(DP_OP_102J5_124_3590_n908) );
  FADDX1_HVT DP_OP_102J5_124_3590_U568 ( .A(DP_OP_102J5_124_3590_n912), .B(
        DP_OP_102J5_124_3590_n910), .CI(DP_OP_102J5_124_3590_n1055), .CO(
        DP_OP_102J5_124_3590_n905), .S(DP_OP_102J5_124_3590_n906) );
  FADDX1_HVT DP_OP_102J5_124_3590_U567 ( .A(DP_OP_102J5_124_3590_n2081), .B(
        DP_OP_102J5_124_3590_n1905), .CI(DP_OP_102J5_124_3590_n1510), .CO(
        DP_OP_102J5_124_3590_n903), .S(DP_OP_102J5_124_3590_n904) );
  FADDX1_HVT DP_OP_102J5_124_3590_U566 ( .A(DP_OP_102J5_124_3590_n2169), .B(
        DP_OP_102J5_124_3590_n2037), .CI(DP_OP_102J5_124_3590_n1993), .CO(
        DP_OP_102J5_124_3590_n901), .S(DP_OP_102J5_124_3590_n902) );
  FADDX1_HVT DP_OP_102J5_124_3590_U565 ( .A(DP_OP_102J5_124_3590_n1949), .B(
        DP_OP_102J5_124_3590_n1730), .CI(DP_OP_102J5_124_3590_n1817), .CO(
        DP_OP_102J5_124_3590_n899), .S(DP_OP_102J5_124_3590_n900) );
  FADDX1_HVT DP_OP_102J5_124_3590_U564 ( .A(DP_OP_102J5_124_3590_n2213), .B(
        DP_OP_102J5_124_3590_n1598), .CI(DP_OP_102J5_124_3590_n2125), .CO(
        DP_OP_102J5_124_3590_n897), .S(DP_OP_102J5_124_3590_n898) );
  FADDX1_HVT DP_OP_102J5_124_3590_U563 ( .A(DP_OP_102J5_124_3590_n1554), .B(
        DP_OP_102J5_124_3590_n2301), .CI(DP_OP_102J5_124_3590_n1686), .CO(
        DP_OP_102J5_124_3590_n895), .S(DP_OP_102J5_124_3590_n896) );
  FADDX1_HVT DP_OP_102J5_124_3590_U562 ( .A(DP_OP_102J5_124_3590_n2345), .B(
        DP_OP_102J5_124_3590_n1774), .CI(DP_OP_102J5_124_3590_n2257), .CO(
        DP_OP_102J5_124_3590_n893), .S(DP_OP_102J5_124_3590_n894) );
  FADDX1_HVT DP_OP_102J5_124_3590_U561 ( .A(DP_OP_102J5_124_3590_n1642), .B(
        DP_OP_102J5_124_3590_n1861), .CI(DP_OP_102J5_124_3590_n1868), .CO(
        DP_OP_102J5_124_3590_n891), .S(DP_OP_102J5_124_3590_n892) );
  FADDX1_HVT DP_OP_102J5_124_3590_U560 ( .A(DP_OP_102J5_124_3590_n1875), .B(
        DP_OP_102J5_124_3590_n2365), .CI(DP_OP_102J5_124_3590_n2359), .CO(
        DP_OP_102J5_124_3590_n889), .S(DP_OP_102J5_124_3590_n890) );
  FADDX1_HVT DP_OP_102J5_124_3590_U559 ( .A(DP_OP_102J5_124_3590_n1831), .B(
        DP_OP_102J5_124_3590_n2352), .CI(DP_OP_102J5_124_3590_n2322), .CO(
        DP_OP_102J5_124_3590_n887), .S(DP_OP_102J5_124_3590_n888) );
  FADDX1_HVT DP_OP_102J5_124_3590_U558 ( .A(DP_OP_102J5_124_3590_n1824), .B(
        DP_OP_102J5_124_3590_n2315), .CI(DP_OP_102J5_124_3590_n1517), .CO(
        DP_OP_102J5_124_3590_n885), .S(DP_OP_102J5_124_3590_n886) );
  FADDX1_HVT DP_OP_102J5_124_3590_U557 ( .A(DP_OP_102J5_124_3590_n1795), .B(
        DP_OP_102J5_124_3590_n2308), .CI(DP_OP_102J5_124_3590_n2278), .CO(
        DP_OP_102J5_124_3590_n883), .S(DP_OP_102J5_124_3590_n884) );
  FADDX1_HVT DP_OP_102J5_124_3590_U556 ( .A(DP_OP_102J5_124_3590_n1788), .B(
        DP_OP_102J5_124_3590_n2271), .CI(DP_OP_102J5_124_3590_n2264), .CO(
        DP_OP_102J5_124_3590_n881), .S(DP_OP_102J5_124_3590_n882) );
  FADDX1_HVT DP_OP_102J5_124_3590_U555 ( .A(DP_OP_102J5_124_3590_n1751), .B(
        DP_OP_102J5_124_3590_n2234), .CI(DP_OP_102J5_124_3590_n2227), .CO(
        DP_OP_102J5_124_3590_n879), .S(DP_OP_102J5_124_3590_n880) );
  FADDX1_HVT DP_OP_102J5_124_3590_U554 ( .A(DP_OP_102J5_124_3590_n1744), .B(
        DP_OP_102J5_124_3590_n2220), .CI(DP_OP_102J5_124_3590_n2190), .CO(
        DP_OP_102J5_124_3590_n877), .S(DP_OP_102J5_124_3590_n878) );
  FADDX1_HVT DP_OP_102J5_124_3590_U553 ( .A(DP_OP_102J5_124_3590_n2183), .B(
        DP_OP_102J5_124_3590_n1524), .CI(DP_OP_102J5_124_3590_n1531), .CO(
        DP_OP_102J5_124_3590_n875), .S(DP_OP_102J5_124_3590_n876) );
  FADDX1_HVT DP_OP_102J5_124_3590_U552 ( .A(DP_OP_102J5_124_3590_n1956), .B(
        DP_OP_102J5_124_3590_n2176), .CI(DP_OP_102J5_124_3590_n2146), .CO(
        DP_OP_102J5_124_3590_n873), .S(DP_OP_102J5_124_3590_n874) );
  FADDX1_HVT DP_OP_102J5_124_3590_U551 ( .A(DP_OP_102J5_124_3590_n2139), .B(
        DP_OP_102J5_124_3590_n1561), .CI(DP_OP_102J5_124_3590_n1568), .CO(
        DP_OP_102J5_124_3590_n871), .S(DP_OP_102J5_124_3590_n872) );
  FADDX1_HVT DP_OP_102J5_124_3590_U550 ( .A(DP_OP_102J5_124_3590_n2132), .B(
        DP_OP_102J5_124_3590_n1575), .CI(DP_OP_102J5_124_3590_n1605), .CO(
        DP_OP_102J5_124_3590_n869), .S(DP_OP_102J5_124_3590_n870) );
  FADDX1_HVT DP_OP_102J5_124_3590_U549 ( .A(DP_OP_102J5_124_3590_n2102), .B(
        DP_OP_102J5_124_3590_n1612), .CI(DP_OP_102J5_124_3590_n1619), .CO(
        DP_OP_102J5_124_3590_n867), .S(DP_OP_102J5_124_3590_n868) );
  FADDX1_HVT DP_OP_102J5_124_3590_U548 ( .A(DP_OP_102J5_124_3590_n2095), .B(
        DP_OP_102J5_124_3590_n1649), .CI(DP_OP_102J5_124_3590_n1656), .CO(
        DP_OP_102J5_124_3590_n865), .S(DP_OP_102J5_124_3590_n866) );
  FADDX1_HVT DP_OP_102J5_124_3590_U547 ( .A(DP_OP_102J5_124_3590_n2088), .B(
        DP_OP_102J5_124_3590_n1663), .CI(DP_OP_102J5_124_3590_n1693), .CO(
        DP_OP_102J5_124_3590_n863), .S(DP_OP_102J5_124_3590_n864) );
  FADDX1_HVT DP_OP_102J5_124_3590_U546 ( .A(DP_OP_102J5_124_3590_n2058), .B(
        DP_OP_102J5_124_3590_n1700), .CI(DP_OP_102J5_124_3590_n1707), .CO(
        DP_OP_102J5_124_3590_n861), .S(DP_OP_102J5_124_3590_n862) );
  FADDX1_HVT DP_OP_102J5_124_3590_U545 ( .A(DP_OP_102J5_124_3590_n2051), .B(
        DP_OP_102J5_124_3590_n1737), .CI(DP_OP_102J5_124_3590_n1781), .CO(
        DP_OP_102J5_124_3590_n859), .S(DP_OP_102J5_124_3590_n860) );
  FADDX1_HVT DP_OP_102J5_124_3590_U544 ( .A(DP_OP_102J5_124_3590_n2044), .B(
        DP_OP_102J5_124_3590_n1838), .CI(DP_OP_102J5_124_3590_n1882), .CO(
        DP_OP_102J5_124_3590_n857), .S(DP_OP_102J5_124_3590_n858) );
  FADDX1_HVT DP_OP_102J5_124_3590_U543 ( .A(DP_OP_102J5_124_3590_n2014), .B(
        DP_OP_102J5_124_3590_n1912), .CI(DP_OP_102J5_124_3590_n1919), .CO(
        DP_OP_102J5_124_3590_n855), .S(DP_OP_102J5_124_3590_n856) );
  FADDX1_HVT DP_OP_102J5_124_3590_U542 ( .A(DP_OP_102J5_124_3590_n2007), .B(
        DP_OP_102J5_124_3590_n1926), .CI(DP_OP_102J5_124_3590_n1963), .CO(
        DP_OP_102J5_124_3590_n853), .S(DP_OP_102J5_124_3590_n854) );
  FADDX1_HVT DP_OP_102J5_124_3590_U541 ( .A(DP_OP_102J5_124_3590_n2000), .B(
        DP_OP_102J5_124_3590_n1970), .CI(DP_OP_102J5_124_3590_n1053), .CO(
        DP_OP_102J5_124_3590_n851), .S(DP_OP_102J5_124_3590_n852) );
  FADDX1_HVT DP_OP_102J5_124_3590_U540 ( .A(DP_OP_102J5_124_3590_n1045), .B(
        DP_OP_102J5_124_3590_n1041), .CI(DP_OP_102J5_124_3590_n1047), .CO(
        DP_OP_102J5_124_3590_n849), .S(DP_OP_102J5_124_3590_n850) );
  FADDX1_HVT DP_OP_102J5_124_3590_U539 ( .A(DP_OP_102J5_124_3590_n1051), .B(
        DP_OP_102J5_124_3590_n1043), .CI(DP_OP_102J5_124_3590_n1049), .CO(
        DP_OP_102J5_124_3590_n847), .S(DP_OP_102J5_124_3590_n848) );
  FADDX1_HVT DP_OP_102J5_124_3590_U538 ( .A(DP_OP_102J5_124_3590_n1021), .B(
        DP_OP_102J5_124_3590_n1001), .CI(DP_OP_102J5_124_3590_n1005), .CO(
        DP_OP_102J5_124_3590_n845), .S(DP_OP_102J5_124_3590_n846) );
  FADDX1_HVT DP_OP_102J5_124_3590_U537 ( .A(DP_OP_102J5_124_3590_n1023), .B(
        DP_OP_102J5_124_3590_n1003), .CI(DP_OP_102J5_124_3590_n1007), .CO(
        DP_OP_102J5_124_3590_n843), .S(DP_OP_102J5_124_3590_n844) );
  FADDX1_HVT DP_OP_102J5_124_3590_U536 ( .A(DP_OP_102J5_124_3590_n1019), .B(
        DP_OP_102J5_124_3590_n1009), .CI(DP_OP_102J5_124_3590_n1011), .CO(
        DP_OP_102J5_124_3590_n841), .S(DP_OP_102J5_124_3590_n842) );
  FADDX1_HVT DP_OP_102J5_124_3590_U535 ( .A(DP_OP_102J5_124_3590_n1017), .B(
        DP_OP_102J5_124_3590_n1013), .CI(DP_OP_102J5_124_3590_n1025), .CO(
        DP_OP_102J5_124_3590_n839), .S(DP_OP_102J5_124_3590_n840) );
  FADDX1_HVT DP_OP_102J5_124_3590_U534 ( .A(DP_OP_102J5_124_3590_n1033), .B(
        DP_OP_102J5_124_3590_n1015), .CI(DP_OP_102J5_124_3590_n1029), .CO(
        DP_OP_102J5_124_3590_n837), .S(DP_OP_102J5_124_3590_n838) );
  FADDX1_HVT DP_OP_102J5_124_3590_U533 ( .A(DP_OP_102J5_124_3590_n1035), .B(
        DP_OP_102J5_124_3590_n1027), .CI(DP_OP_102J5_124_3590_n1037), .CO(
        DP_OP_102J5_124_3590_n835), .S(DP_OP_102J5_124_3590_n836) );
  FADDX1_HVT DP_OP_102J5_124_3590_U532 ( .A(DP_OP_102J5_124_3590_n1039), .B(
        DP_OP_102J5_124_3590_n1031), .CI(DP_OP_102J5_124_3590_n896), .CO(
        DP_OP_102J5_124_3590_n833), .S(DP_OP_102J5_124_3590_n834) );
  FADDX1_HVT DP_OP_102J5_124_3590_U531 ( .A(DP_OP_102J5_124_3590_n898), .B(
        DP_OP_102J5_124_3590_n904), .CI(DP_OP_102J5_124_3590_n892), .CO(
        DP_OP_102J5_124_3590_n831), .S(DP_OP_102J5_124_3590_n832) );
  FADDX1_HVT DP_OP_102J5_124_3590_U530 ( .A(DP_OP_102J5_124_3590_n894), .B(
        DP_OP_102J5_124_3590_n902), .CI(DP_OP_102J5_124_3590_n900), .CO(
        DP_OP_102J5_124_3590_n829), .S(DP_OP_102J5_124_3590_n830) );
  FADDX1_HVT DP_OP_102J5_124_3590_U529 ( .A(DP_OP_102J5_124_3590_n858), .B(
        DP_OP_102J5_124_3590_n884), .CI(DP_OP_102J5_124_3590_n890), .CO(
        DP_OP_102J5_124_3590_n827), .S(DP_OP_102J5_124_3590_n828) );
  FADDX1_HVT DP_OP_102J5_124_3590_U528 ( .A(DP_OP_102J5_124_3590_n880), .B(
        DP_OP_102J5_124_3590_n874), .CI(DP_OP_102J5_124_3590_n872), .CO(
        DP_OP_102J5_124_3590_n825), .S(DP_OP_102J5_124_3590_n826) );
  FADDX1_HVT DP_OP_102J5_124_3590_U527 ( .A(DP_OP_102J5_124_3590_n882), .B(
        DP_OP_102J5_124_3590_n870), .CI(DP_OP_102J5_124_3590_n868), .CO(
        DP_OP_102J5_124_3590_n823), .S(DP_OP_102J5_124_3590_n824) );
  FADDX1_HVT DP_OP_102J5_124_3590_U526 ( .A(DP_OP_102J5_124_3590_n876), .B(
        DP_OP_102J5_124_3590_n866), .CI(DP_OP_102J5_124_3590_n854), .CO(
        DP_OP_102J5_124_3590_n821), .S(DP_OP_102J5_124_3590_n822) );
  FADDX1_HVT DP_OP_102J5_124_3590_U525 ( .A(DP_OP_102J5_124_3590_n878), .B(
        DP_OP_102J5_124_3590_n860), .CI(DP_OP_102J5_124_3590_n856), .CO(
        DP_OP_102J5_124_3590_n819), .S(DP_OP_102J5_124_3590_n820) );
  FADDX1_HVT DP_OP_102J5_124_3590_U524 ( .A(DP_OP_102J5_124_3590_n864), .B(
        DP_OP_102J5_124_3590_n888), .CI(DP_OP_102J5_124_3590_n886), .CO(
        DP_OP_102J5_124_3590_n817), .S(DP_OP_102J5_124_3590_n818) );
  FADDX1_HVT DP_OP_102J5_124_3590_U523 ( .A(DP_OP_102J5_124_3590_n862), .B(
        DP_OP_102J5_124_3590_n852), .CI(DP_OP_102J5_124_3590_n997), .CO(
        DP_OP_102J5_124_3590_n815), .S(DP_OP_102J5_124_3590_n816) );
  FADDX1_HVT DP_OP_102J5_124_3590_U522 ( .A(DP_OP_102J5_124_3590_n995), .B(
        DP_OP_102J5_124_3590_n999), .CI(DP_OP_102J5_124_3590_n985), .CO(
        DP_OP_102J5_124_3590_n813), .S(DP_OP_102J5_124_3590_n814) );
  FADDX1_HVT DP_OP_102J5_124_3590_U521 ( .A(DP_OP_102J5_124_3590_n983), .B(
        DP_OP_102J5_124_3590_n989), .CI(DP_OP_102J5_124_3590_n1475), .CO(
        DP_OP_102J5_124_3590_n811), .S(DP_OP_102J5_124_3590_n812) );
  FADDX1_HVT DP_OP_102J5_124_3590_U520 ( .A(DP_OP_102J5_124_3590_n987), .B(
        DP_OP_102J5_124_3590_n991), .CI(DP_OP_102J5_124_3590_n993), .CO(
        DP_OP_102J5_124_3590_n809), .S(DP_OP_102J5_124_3590_n810) );
  FADDX1_HVT DP_OP_102J5_124_3590_U519 ( .A(DP_OP_102J5_124_3590_n981), .B(
        DP_OP_102J5_124_3590_n979), .CI(DP_OP_102J5_124_3590_n977), .CO(
        DP_OP_102J5_124_3590_n807), .S(DP_OP_102J5_124_3590_n808) );
  FADDX1_HVT DP_OP_102J5_124_3590_U518 ( .A(DP_OP_102J5_124_3590_n848), .B(
        DP_OP_102J5_124_3590_n850), .CI(DP_OP_102J5_124_3590_n844), .CO(
        DP_OP_102J5_124_3590_n805), .S(DP_OP_102J5_124_3590_n806) );
  FADDX1_HVT DP_OP_102J5_124_3590_U517 ( .A(DP_OP_102J5_124_3590_n840), .B(
        DP_OP_102J5_124_3590_n846), .CI(DP_OP_102J5_124_3590_n834), .CO(
        DP_OP_102J5_124_3590_n803), .S(DP_OP_102J5_124_3590_n804) );
  FADDX1_HVT DP_OP_102J5_124_3590_U516 ( .A(DP_OP_102J5_124_3590_n975), .B(
        DP_OP_102J5_124_3590_n842), .CI(DP_OP_102J5_124_3590_n838), .CO(
        DP_OP_102J5_124_3590_n801), .S(DP_OP_102J5_124_3590_n802) );
  FADDX1_HVT DP_OP_102J5_124_3590_U515 ( .A(DP_OP_102J5_124_3590_n973), .B(
        DP_OP_102J5_124_3590_n836), .CI(DP_OP_102J5_124_3590_n965), .CO(
        DP_OP_102J5_124_3590_n799), .S(DP_OP_102J5_124_3590_n800) );
  FADDX1_HVT DP_OP_102J5_124_3590_U514 ( .A(DP_OP_102J5_124_3590_n971), .B(
        DP_OP_102J5_124_3590_n967), .CI(DP_OP_102J5_124_3590_n969), .CO(
        DP_OP_102J5_124_3590_n797), .S(DP_OP_102J5_124_3590_n798) );
  FADDX1_HVT DP_OP_102J5_124_3590_U513 ( .A(DP_OP_102J5_124_3590_n830), .B(
        DP_OP_102J5_124_3590_n832), .CI(DP_OP_102J5_124_3590_n826), .CO(
        DP_OP_102J5_124_3590_n795), .S(DP_OP_102J5_124_3590_n796) );
  FADDX1_HVT DP_OP_102J5_124_3590_U512 ( .A(DP_OP_102J5_124_3590_n824), .B(
        DP_OP_102J5_124_3590_n820), .CI(DP_OP_102J5_124_3590_n963), .CO(
        DP_OP_102J5_124_3590_n793), .S(DP_OP_102J5_124_3590_n794) );
  FADDX1_HVT DP_OP_102J5_124_3590_U511 ( .A(DP_OP_102J5_124_3590_n822), .B(
        DP_OP_102J5_124_3590_n828), .CI(DP_OP_102J5_124_3590_n818), .CO(
        DP_OP_102J5_124_3590_n791), .S(DP_OP_102J5_124_3590_n792) );
  FADDX1_HVT DP_OP_102J5_124_3590_U510 ( .A(DP_OP_102J5_124_3590_n961), .B(
        DP_OP_102J5_124_3590_n959), .CI(DP_OP_102J5_124_3590_n816), .CO(
        DP_OP_102J5_124_3590_n789), .S(DP_OP_102J5_124_3590_n790) );
  FADDX1_HVT DP_OP_102J5_124_3590_U509 ( .A(DP_OP_102J5_124_3590_n957), .B(
        DP_OP_102J5_124_3590_n955), .CI(DP_OP_102J5_124_3590_n814), .CO(
        DP_OP_102J5_124_3590_n787), .S(DP_OP_102J5_124_3590_n788) );
  FADDX1_HVT DP_OP_102J5_124_3590_U508 ( .A(DP_OP_102J5_124_3590_n953), .B(
        DP_OP_102J5_124_3590_n812), .CI(DP_OP_102J5_124_3590_n810), .CO(
        DP_OP_102J5_124_3590_n785), .S(DP_OP_102J5_124_3590_n786) );
  FADDX1_HVT DP_OP_102J5_124_3590_U507 ( .A(DP_OP_102J5_124_3590_n951), .B(
        DP_OP_102J5_124_3590_n947), .CI(DP_OP_102J5_124_3590_n949), .CO(
        DP_OP_102J5_124_3590_n783), .S(DP_OP_102J5_124_3590_n784) );
  FADDX1_HVT DP_OP_102J5_124_3590_U506 ( .A(DP_OP_102J5_124_3590_n945), .B(
        DP_OP_102J5_124_3590_n806), .CI(DP_OP_102J5_124_3590_n943), .CO(
        DP_OP_102J5_124_3590_n781), .S(DP_OP_102J5_124_3590_n782) );
  FADDX1_HVT DP_OP_102J5_124_3590_U505 ( .A(DP_OP_102J5_124_3590_n808), .B(
        DP_OP_102J5_124_3590_n941), .CI(DP_OP_102J5_124_3590_n802), .CO(
        DP_OP_102J5_124_3590_n779), .S(DP_OP_102J5_124_3590_n780) );
  FADDX1_HVT DP_OP_102J5_124_3590_U504 ( .A(DP_OP_102J5_124_3590_n798), .B(
        DP_OP_102J5_124_3590_n804), .CI(DP_OP_102J5_124_3590_n939), .CO(
        DP_OP_102J5_124_3590_n777), .S(DP_OP_102J5_124_3590_n778) );
  FADDX1_HVT DP_OP_102J5_124_3590_U503 ( .A(DP_OP_102J5_124_3590_n800), .B(
        DP_OP_102J5_124_3590_n796), .CI(DP_OP_102J5_124_3590_n937), .CO(
        DP_OP_102J5_124_3590_n775), .S(DP_OP_102J5_124_3590_n776) );
  FADDX1_HVT DP_OP_102J5_124_3590_U502 ( .A(DP_OP_102J5_124_3590_n792), .B(
        DP_OP_102J5_124_3590_n794), .CI(DP_OP_102J5_124_3590_n935), .CO(
        DP_OP_102J5_124_3590_n773), .S(DP_OP_102J5_124_3590_n774) );
  FADDX1_HVT DP_OP_102J5_124_3590_U501 ( .A(DP_OP_102J5_124_3590_n933), .B(
        DP_OP_102J5_124_3590_n790), .CI(DP_OP_102J5_124_3590_n931), .CO(
        DP_OP_102J5_124_3590_n771), .S(DP_OP_102J5_124_3590_n772) );
  FADDX1_HVT DP_OP_102J5_124_3590_U500 ( .A(DP_OP_102J5_124_3590_n788), .B(
        DP_OP_102J5_124_3590_n929), .CI(DP_OP_102J5_124_3590_n927), .CO(
        DP_OP_102J5_124_3590_n769), .S(DP_OP_102J5_124_3590_n770) );
  FADDX1_HVT DP_OP_102J5_124_3590_U499 ( .A(DP_OP_102J5_124_3590_n786), .B(
        DP_OP_102J5_124_3590_n784), .CI(DP_OP_102J5_124_3590_n925), .CO(
        DP_OP_102J5_124_3590_n767), .S(DP_OP_102J5_124_3590_n768) );
  FADDX1_HVT DP_OP_102J5_124_3590_U498 ( .A(DP_OP_102J5_124_3590_n782), .B(
        DP_OP_102J5_124_3590_n780), .CI(DP_OP_102J5_124_3590_n778), .CO(
        DP_OP_102J5_124_3590_n765), .S(DP_OP_102J5_124_3590_n766) );
  FADDX1_HVT DP_OP_102J5_124_3590_U497 ( .A(DP_OP_102J5_124_3590_n923), .B(
        DP_OP_102J5_124_3590_n776), .CI(DP_OP_102J5_124_3590_n921), .CO(
        DP_OP_102J5_124_3590_n763), .S(DP_OP_102J5_124_3590_n764) );
  FADDX1_HVT DP_OP_102J5_124_3590_U496 ( .A(DP_OP_102J5_124_3590_n774), .B(
        DP_OP_102J5_124_3590_n919), .CI(DP_OP_102J5_124_3590_n772), .CO(
        DP_OP_102J5_124_3590_n761), .S(DP_OP_102J5_124_3590_n762) );
  FADDX1_HVT DP_OP_102J5_124_3590_U495 ( .A(DP_OP_102J5_124_3590_n917), .B(
        DP_OP_102J5_124_3590_n770), .CI(DP_OP_102J5_124_3590_n915), .CO(
        DP_OP_102J5_124_3590_n759), .S(DP_OP_102J5_124_3590_n760) );
  FADDX1_HVT DP_OP_102J5_124_3590_U494 ( .A(DP_OP_102J5_124_3590_n768), .B(
        DP_OP_102J5_124_3590_n766), .CI(DP_OP_102J5_124_3590_n913), .CO(
        DP_OP_102J5_124_3590_n757), .S(DP_OP_102J5_124_3590_n758) );
  FADDX1_HVT DP_OP_102J5_124_3590_U493 ( .A(DP_OP_102J5_124_3590_n764), .B(
        DP_OP_102J5_124_3590_n911), .CI(DP_OP_102J5_124_3590_n762), .CO(
        DP_OP_102J5_124_3590_n755), .S(DP_OP_102J5_124_3590_n756) );
  FADDX1_HVT DP_OP_102J5_124_3590_U492 ( .A(DP_OP_102J5_124_3590_n909), .B(
        DP_OP_102J5_124_3590_n760), .CI(DP_OP_102J5_124_3590_n758), .CO(
        DP_OP_102J5_124_3590_n753), .S(DP_OP_102J5_124_3590_n754) );
  FADDX1_HVT DP_OP_102J5_124_3590_U491 ( .A(DP_OP_102J5_124_3590_n907), .B(
        DP_OP_102J5_124_3590_n756), .CI(DP_OP_102J5_124_3590_n905), .CO(
        DP_OP_102J5_124_3590_n751), .S(DP_OP_102J5_124_3590_n752) );
  FADDX1_HVT DP_OP_102J5_124_3590_U489 ( .A(DP_OP_102J5_124_3590_n1881), .B(
        DP_OP_102J5_124_3590_n1530), .CI(DP_OP_102J5_124_3590_n1509), .CO(
        DP_OP_102J5_124_3590_n747), .S(DP_OP_102J5_124_3590_n748) );
  FADDX1_HVT DP_OP_102J5_124_3590_U488 ( .A(DP_OP_102J5_124_3590_n2277), .B(
        DP_OP_102J5_124_3590_n1729), .CI(DP_OP_102J5_124_3590_n1860), .CO(
        DP_OP_102J5_124_3590_n745), .S(DP_OP_102J5_124_3590_n746) );
  FADDX1_HVT DP_OP_102J5_124_3590_U487 ( .A(DP_OP_102J5_124_3590_n1553), .B(
        DP_OP_102J5_124_3590_n1618), .CI(DP_OP_102J5_124_3590_n1750), .CO(
        DP_OP_102J5_124_3590_n743), .S(DP_OP_102J5_124_3590_n744) );
  FADDX1_HVT DP_OP_102J5_124_3590_U486 ( .A(DP_OP_102J5_124_3590_n1992), .B(
        DP_OP_102J5_124_3590_n1948), .CI(DP_OP_102J5_124_3590_n1816), .CO(
        DP_OP_102J5_124_3590_n741), .S(DP_OP_102J5_124_3590_n742) );
  FADDX1_HVT DP_OP_102J5_124_3590_U485 ( .A(DP_OP_102J5_124_3590_n2168), .B(
        DP_OP_102J5_124_3590_n2013), .CI(DP_OP_102J5_124_3590_n2057), .CO(
        DP_OP_102J5_124_3590_n739), .S(DP_OP_102J5_124_3590_n740) );
  FADDX1_HVT DP_OP_102J5_124_3590_U484 ( .A(DP_OP_102J5_124_3590_n1904), .B(
        DP_OP_102J5_124_3590_n1837), .CI(DP_OP_102J5_124_3590_n1597), .CO(
        DP_OP_102J5_124_3590_n737), .S(DP_OP_102J5_124_3590_n738) );
  FADDX1_HVT DP_OP_102J5_124_3590_U483 ( .A(DP_OP_102J5_124_3590_n1662), .B(
        DP_OP_102J5_124_3590_n2080), .CI(DP_OP_102J5_124_3590_n1925), .CO(
        DP_OP_102J5_124_3590_n735), .S(DP_OP_102J5_124_3590_n736) );
  FADDX1_HVT DP_OP_102J5_124_3590_U482 ( .A(DP_OP_102J5_124_3590_n2300), .B(
        DP_OP_102J5_124_3590_n1641), .CI(DP_OP_102J5_124_3590_n2036), .CO(
        DP_OP_102J5_124_3590_n733), .S(DP_OP_102J5_124_3590_n734) );
  FADDX1_HVT DP_OP_102J5_124_3590_U481 ( .A(DP_OP_102J5_124_3590_n2101), .B(
        DP_OP_102J5_124_3590_n1706), .CI(DP_OP_102J5_124_3590_n1685), .CO(
        DP_OP_102J5_124_3590_n731), .S(DP_OP_102J5_124_3590_n732) );
  FADDX1_HVT DP_OP_102J5_124_3590_U480 ( .A(DP_OP_102J5_124_3590_n2212), .B(
        DP_OP_102J5_124_3590_n2189), .CI(DP_OP_102J5_124_3590_n1969), .CO(
        DP_OP_102J5_124_3590_n729), .S(DP_OP_102J5_124_3590_n730) );
  FADDX1_HVT DP_OP_102J5_124_3590_U479 ( .A(DP_OP_102J5_124_3590_n1773), .B(
        DP_OP_102J5_124_3590_n2233), .CI(DP_OP_102J5_124_3590_n2256), .CO(
        DP_OP_102J5_124_3590_n727), .S(DP_OP_102J5_124_3590_n728) );
  FADDX1_HVT DP_OP_102J5_124_3590_U478 ( .A(DP_OP_102J5_124_3590_n2145), .B(
        DP_OP_102J5_124_3590_n2124), .CI(DP_OP_102J5_124_3590_n2321), .CO(
        DP_OP_102J5_124_3590_n725), .S(DP_OP_102J5_124_3590_n726) );
  FADDX1_HVT DP_OP_102J5_124_3590_U477 ( .A(DP_OP_102J5_124_3590_n1794), .B(
        DP_OP_102J5_124_3590_n2344), .CI(DP_OP_102J5_124_3590_n1574), .CO(
        DP_OP_102J5_124_3590_n723), .S(DP_OP_102J5_124_3590_n724) );
  FADDX1_HVT DP_OP_102J5_124_3590_U476 ( .A(DP_OP_102J5_124_3590_n1823), .B(
        DP_OP_102J5_124_3590_n1516), .CI(DP_OP_102J5_124_3590_n750), .CO(
        DP_OP_102J5_124_3590_n721), .S(DP_OP_102J5_124_3590_n722) );
  FADDX1_HVT DP_OP_102J5_124_3590_U475 ( .A(DP_OP_102J5_124_3590_n2358), .B(
        DP_OP_102J5_124_3590_n1523), .CI(DP_OP_102J5_124_3590_n2351), .CO(
        DP_OP_102J5_124_3590_n719), .S(DP_OP_102J5_124_3590_n720) );
  FADDX1_HVT DP_OP_102J5_124_3590_U474 ( .A(DP_OP_102J5_124_3590_n1999), .B(
        DP_OP_102J5_124_3590_n1560), .CI(DP_OP_102J5_124_3590_n2314), .CO(
        DP_OP_102J5_124_3590_n717), .S(DP_OP_102J5_124_3590_n718) );
  FADDX1_HVT DP_OP_102J5_124_3590_U473 ( .A(DP_OP_102J5_124_3590_n2307), .B(
        DP_OP_102J5_124_3590_n1567), .CI(DP_OP_102J5_124_3590_n1604), .CO(
        DP_OP_102J5_124_3590_n715), .S(DP_OP_102J5_124_3590_n716) );
  FADDX1_HVT DP_OP_102J5_124_3590_U472 ( .A(DP_OP_102J5_124_3590_n2270), .B(
        DP_OP_102J5_124_3590_n1611), .CI(DP_OP_102J5_124_3590_n1648), .CO(
        DP_OP_102J5_124_3590_n713), .S(DP_OP_102J5_124_3590_n714) );
  FADDX1_HVT DP_OP_102J5_124_3590_U471 ( .A(DP_OP_102J5_124_3590_n2263), .B(
        DP_OP_102J5_124_3590_n1655), .CI(DP_OP_102J5_124_3590_n1692), .CO(
        DP_OP_102J5_124_3590_n711), .S(DP_OP_102J5_124_3590_n712) );
  FADDX1_HVT DP_OP_102J5_124_3590_U470 ( .A(DP_OP_102J5_124_3590_n2226), .B(
        DP_OP_102J5_124_3590_n1699), .CI(DP_OP_102J5_124_3590_n1736), .CO(
        DP_OP_102J5_124_3590_n709), .S(DP_OP_102J5_124_3590_n710) );
  FADDX1_HVT DP_OP_102J5_124_3590_U469 ( .A(DP_OP_102J5_124_3590_n2219), .B(
        DP_OP_102J5_124_3590_n1743), .CI(DP_OP_102J5_124_3590_n1780), .CO(
        DP_OP_102J5_124_3590_n707), .S(DP_OP_102J5_124_3590_n708) );
  FADDX1_HVT DP_OP_102J5_124_3590_U468 ( .A(DP_OP_102J5_124_3590_n2182), .B(
        DP_OP_102J5_124_3590_n1787), .CI(DP_OP_102J5_124_3590_n1830), .CO(
        DP_OP_102J5_124_3590_n705), .S(DP_OP_102J5_124_3590_n706) );
  FADDX1_HVT DP_OP_102J5_124_3590_U467 ( .A(DP_OP_102J5_124_3590_n2175), .B(
        DP_OP_102J5_124_3590_n1867), .CI(DP_OP_102J5_124_3590_n1874), .CO(
        DP_OP_102J5_124_3590_n703), .S(DP_OP_102J5_124_3590_n704) );
  FADDX1_HVT DP_OP_102J5_124_3590_U466 ( .A(DP_OP_102J5_124_3590_n2138), .B(
        DP_OP_102J5_124_3590_n1911), .CI(DP_OP_102J5_124_3590_n1918), .CO(
        DP_OP_102J5_124_3590_n701), .S(DP_OP_102J5_124_3590_n702) );
  FADDX1_HVT DP_OP_102J5_124_3590_U465 ( .A(DP_OP_102J5_124_3590_n2131), .B(
        DP_OP_102J5_124_3590_n1955), .CI(DP_OP_102J5_124_3590_n1962), .CO(
        DP_OP_102J5_124_3590_n699), .S(DP_OP_102J5_124_3590_n700) );
  FADDX1_HVT DP_OP_102J5_124_3590_U464 ( .A(DP_OP_102J5_124_3590_n2094), .B(
        DP_OP_102J5_124_3590_n2006), .CI(DP_OP_102J5_124_3590_n2043), .CO(
        DP_OP_102J5_124_3590_n697), .S(DP_OP_102J5_124_3590_n698) );
  FADDX1_HVT DP_OP_102J5_124_3590_U463 ( .A(DP_OP_102J5_124_3590_n2087), .B(
        DP_OP_102J5_124_3590_n2050), .CI(DP_OP_102J5_124_3590_n897), .CO(
        DP_OP_102J5_124_3590_n695), .S(DP_OP_102J5_124_3590_n696) );
  FADDX1_HVT DP_OP_102J5_124_3590_U462 ( .A(DP_OP_102J5_124_3590_n895), .B(
        DP_OP_102J5_124_3590_n891), .CI(DP_OP_102J5_124_3590_n899), .CO(
        DP_OP_102J5_124_3590_n693), .S(DP_OP_102J5_124_3590_n694) );
  FADDX1_HVT DP_OP_102J5_124_3590_U461 ( .A(DP_OP_102J5_124_3590_n903), .B(
        DP_OP_102J5_124_3590_n893), .CI(DP_OP_102J5_124_3590_n901), .CO(
        DP_OP_102J5_124_3590_n691), .S(DP_OP_102J5_124_3590_n692) );
  FADDX1_HVT DP_OP_102J5_124_3590_U460 ( .A(DP_OP_102J5_124_3590_n873), .B(
        DP_OP_102J5_124_3590_n855), .CI(DP_OP_102J5_124_3590_n851), .CO(
        DP_OP_102J5_124_3590_n689), .S(DP_OP_102J5_124_3590_n690) );
  FADDX1_HVT DP_OP_102J5_124_3590_U459 ( .A(DP_OP_102J5_124_3590_n871), .B(
        DP_OP_102J5_124_3590_n853), .CI(DP_OP_102J5_124_3590_n857), .CO(
        DP_OP_102J5_124_3590_n687), .S(DP_OP_102J5_124_3590_n688) );
  FADDX1_HVT DP_OP_102J5_124_3590_U458 ( .A(DP_OP_102J5_124_3590_n867), .B(
        DP_OP_102J5_124_3590_n861), .CI(DP_OP_102J5_124_3590_n859), .CO(
        DP_OP_102J5_124_3590_n685), .S(DP_OP_102J5_124_3590_n686) );
  FADDX1_HVT DP_OP_102J5_124_3590_U457 ( .A(DP_OP_102J5_124_3590_n869), .B(
        DP_OP_102J5_124_3590_n863), .CI(DP_OP_102J5_124_3590_n875), .CO(
        DP_OP_102J5_124_3590_n683), .S(DP_OP_102J5_124_3590_n684) );
  FADDX1_HVT DP_OP_102J5_124_3590_U456 ( .A(DP_OP_102J5_124_3590_n865), .B(
        DP_OP_102J5_124_3590_n877), .CI(DP_OP_102J5_124_3590_n881), .CO(
        DP_OP_102J5_124_3590_n681), .S(DP_OP_102J5_124_3590_n682) );
  FADDX1_HVT DP_OP_102J5_124_3590_U455 ( .A(DP_OP_102J5_124_3590_n885), .B(
        DP_OP_102J5_124_3590_n879), .CI(DP_OP_102J5_124_3590_n887), .CO(
        DP_OP_102J5_124_3590_n679), .S(DP_OP_102J5_124_3590_n680) );
  FADDX1_HVT DP_OP_102J5_124_3590_U454 ( .A(DP_OP_102J5_124_3590_n889), .B(
        DP_OP_102J5_124_3590_n883), .CI(DP_OP_102J5_124_3590_n742), .CO(
        DP_OP_102J5_124_3590_n677), .S(DP_OP_102J5_124_3590_n678) );
  FADDX1_HVT DP_OP_102J5_124_3590_U453 ( .A(DP_OP_102J5_124_3590_n738), .B(
        DP_OP_102J5_124_3590_n726), .CI(DP_OP_102J5_124_3590_n724), .CO(
        DP_OP_102J5_124_3590_n675), .S(DP_OP_102J5_124_3590_n676) );
  FADDX1_HVT DP_OP_102J5_124_3590_U452 ( .A(DP_OP_102J5_124_3590_n740), .B(
        DP_OP_102J5_124_3590_n736), .CI(DP_OP_102J5_124_3590_n732), .CO(
        DP_OP_102J5_124_3590_n673), .S(DP_OP_102J5_124_3590_n674) );
  FADDX1_HVT DP_OP_102J5_124_3590_U451 ( .A(DP_OP_102J5_124_3590_n744), .B(
        DP_OP_102J5_124_3590_n728), .CI(DP_OP_102J5_124_3590_n730), .CO(
        DP_OP_102J5_124_3590_n671), .S(DP_OP_102J5_124_3590_n672) );
  FADDX1_HVT DP_OP_102J5_124_3590_U450 ( .A(DP_OP_102J5_124_3590_n746), .B(
        DP_OP_102J5_124_3590_n748), .CI(DP_OP_102J5_124_3590_n734), .CO(
        DP_OP_102J5_124_3590_n669), .S(DP_OP_102J5_124_3590_n670) );
  FADDX1_HVT DP_OP_102J5_124_3590_U449 ( .A(DP_OP_102J5_124_3590_n716), .B(
        DP_OP_102J5_124_3590_n714), .CI(DP_OP_102J5_124_3590_n710), .CO(
        DP_OP_102J5_124_3590_n667), .S(DP_OP_102J5_124_3590_n668) );
  FADDX1_HVT DP_OP_102J5_124_3590_U448 ( .A(DP_OP_102J5_124_3590_n718), .B(
        DP_OP_102J5_124_3590_n700), .CI(DP_OP_102J5_124_3590_n698), .CO(
        DP_OP_102J5_124_3590_n665), .S(DP_OP_102J5_124_3590_n666) );
  FADDX1_HVT DP_OP_102J5_124_3590_U447 ( .A(DP_OP_102J5_124_3590_n708), .B(
        DP_OP_102J5_124_3590_n706), .CI(DP_OP_102J5_124_3590_n702), .CO(
        DP_OP_102J5_124_3590_n663), .S(DP_OP_102J5_124_3590_n664) );
  FADDX1_HVT DP_OP_102J5_124_3590_U446 ( .A(DP_OP_102J5_124_3590_n712), .B(
        DP_OP_102J5_124_3590_n722), .CI(DP_OP_102J5_124_3590_n720), .CO(
        DP_OP_102J5_124_3590_n661), .S(DP_OP_102J5_124_3590_n662) );
  FADDX1_HVT DP_OP_102J5_124_3590_U445 ( .A(DP_OP_102J5_124_3590_n704), .B(
        DP_OP_102J5_124_3590_n847), .CI(DP_OP_102J5_124_3590_n849), .CO(
        DP_OP_102J5_124_3590_n659), .S(DP_OP_102J5_124_3590_n660) );
  FADDX1_HVT DP_OP_102J5_124_3590_U444 ( .A(DP_OP_102J5_124_3590_n837), .B(
        DP_OP_102J5_124_3590_n839), .CI(DP_OP_102J5_124_3590_n696), .CO(
        DP_OP_102J5_124_3590_n657), .S(DP_OP_102J5_124_3590_n658) );
  FADDX1_HVT DP_OP_102J5_124_3590_U443 ( .A(DP_OP_102J5_124_3590_n843), .B(
        DP_OP_102J5_124_3590_n835), .CI(DP_OP_102J5_124_3590_n1474), .CO(
        DP_OP_102J5_124_3590_n655), .S(DP_OP_102J5_124_3590_n656) );
  FADDX1_HVT DP_OP_102J5_124_3590_U442 ( .A(DP_OP_102J5_124_3590_n845), .B(
        DP_OP_102J5_124_3590_n841), .CI(DP_OP_102J5_124_3590_n833), .CO(
        DP_OP_102J5_124_3590_n653), .S(DP_OP_102J5_124_3590_n654) );
  FADDX1_HVT DP_OP_102J5_124_3590_U441 ( .A(DP_OP_102J5_124_3590_n831), .B(
        DP_OP_102J5_124_3590_n829), .CI(DP_OP_102J5_124_3590_n694), .CO(
        DP_OP_102J5_124_3590_n651), .S(DP_OP_102J5_124_3590_n652) );
  FADDX1_HVT DP_OP_102J5_124_3590_U440 ( .A(DP_OP_102J5_124_3590_n692), .B(
        DP_OP_102J5_124_3590_n688), .CI(DP_OP_102J5_124_3590_n684), .CO(
        DP_OP_102J5_124_3590_n649), .S(DP_OP_102J5_124_3590_n650) );
  FADDX1_HVT DP_OP_102J5_124_3590_U439 ( .A(DP_OP_102J5_124_3590_n686), .B(
        DP_OP_102J5_124_3590_n690), .CI(DP_OP_102J5_124_3590_n678), .CO(
        DP_OP_102J5_124_3590_n647), .S(DP_OP_102J5_124_3590_n648) );
  FADDX1_HVT DP_OP_102J5_124_3590_U438 ( .A(DP_OP_102J5_124_3590_n827), .B(
        DP_OP_102J5_124_3590_n682), .CI(DP_OP_102J5_124_3590_n680), .CO(
        DP_OP_102J5_124_3590_n645), .S(DP_OP_102J5_124_3590_n646) );
  FADDX1_HVT DP_OP_102J5_124_3590_U437 ( .A(DP_OP_102J5_124_3590_n817), .B(
        DP_OP_102J5_124_3590_n825), .CI(DP_OP_102J5_124_3590_n819), .CO(
        DP_OP_102J5_124_3590_n643), .S(DP_OP_102J5_124_3590_n644) );
  FADDX1_HVT DP_OP_102J5_124_3590_U436 ( .A(DP_OP_102J5_124_3590_n823), .B(
        DP_OP_102J5_124_3590_n821), .CI(DP_OP_102J5_124_3590_n672), .CO(
        DP_OP_102J5_124_3590_n641), .S(DP_OP_102J5_124_3590_n642) );
  FADDX1_HVT DP_OP_102J5_124_3590_U435 ( .A(DP_OP_102J5_124_3590_n674), .B(
        DP_OP_102J5_124_3590_n676), .CI(DP_OP_102J5_124_3590_n815), .CO(
        DP_OP_102J5_124_3590_n639), .S(DP_OP_102J5_124_3590_n640) );
  FADDX1_HVT DP_OP_102J5_124_3590_U434 ( .A(DP_OP_102J5_124_3590_n670), .B(
        DP_OP_102J5_124_3590_n664), .CI(DP_OP_102J5_124_3590_n666), .CO(
        DP_OP_102J5_124_3590_n637), .S(DP_OP_102J5_124_3590_n638) );
  FADDX1_HVT DP_OP_102J5_124_3590_U433 ( .A(DP_OP_102J5_124_3590_n662), .B(
        DP_OP_102J5_124_3590_n668), .CI(DP_OP_102J5_124_3590_n813), .CO(
        DP_OP_102J5_124_3590_n635), .S(DP_OP_102J5_124_3590_n636) );
  FADDX1_HVT DP_OP_102J5_124_3590_U432 ( .A(DP_OP_102J5_124_3590_n811), .B(
        DP_OP_102J5_124_3590_n809), .CI(DP_OP_102J5_124_3590_n660), .CO(
        DP_OP_102J5_124_3590_n633), .S(DP_OP_102J5_124_3590_n634) );
  FADDX1_HVT DP_OP_102J5_124_3590_U431 ( .A(DP_OP_102J5_124_3590_n807), .B(
        DP_OP_102J5_124_3590_n805), .CI(DP_OP_102J5_124_3590_n803), .CO(
        DP_OP_102J5_124_3590_n631), .S(DP_OP_102J5_124_3590_n632) );
  FADDX1_HVT DP_OP_102J5_124_3590_U430 ( .A(DP_OP_102J5_124_3590_n801), .B(
        DP_OP_102J5_124_3590_n654), .CI(DP_OP_102J5_124_3590_n658), .CO(
        DP_OP_102J5_124_3590_n629), .S(DP_OP_102J5_124_3590_n630) );
  FADDX1_HVT DP_OP_102J5_124_3590_U429 ( .A(DP_OP_102J5_124_3590_n799), .B(
        DP_OP_102J5_124_3590_n656), .CI(DP_OP_102J5_124_3590_n797), .CO(
        DP_OP_102J5_124_3590_n627), .S(DP_OP_102J5_124_3590_n628) );
  FADDX1_HVT DP_OP_102J5_124_3590_U428 ( .A(DP_OP_102J5_124_3590_n795), .B(
        DP_OP_102J5_124_3590_n652), .CI(DP_OP_102J5_124_3590_n650), .CO(
        DP_OP_102J5_124_3590_n625), .S(DP_OP_102J5_124_3590_n626) );
  FADDX1_HVT DP_OP_102J5_124_3590_U427 ( .A(DP_OP_102J5_124_3590_n793), .B(
        DP_OP_102J5_124_3590_n646), .CI(DP_OP_102J5_124_3590_n642), .CO(
        DP_OP_102J5_124_3590_n623), .S(DP_OP_102J5_124_3590_n624) );
  FADDX1_HVT DP_OP_102J5_124_3590_U426 ( .A(DP_OP_102J5_124_3590_n791), .B(
        DP_OP_102J5_124_3590_n644), .CI(DP_OP_102J5_124_3590_n648), .CO(
        DP_OP_102J5_124_3590_n621), .S(DP_OP_102J5_124_3590_n622) );
  FADDX1_HVT DP_OP_102J5_124_3590_U425 ( .A(DP_OP_102J5_124_3590_n789), .B(
        DP_OP_102J5_124_3590_n640), .CI(DP_OP_102J5_124_3590_n638), .CO(
        DP_OP_102J5_124_3590_n619), .S(DP_OP_102J5_124_3590_n620) );
  FADDX1_HVT DP_OP_102J5_124_3590_U424 ( .A(DP_OP_102J5_124_3590_n787), .B(
        DP_OP_102J5_124_3590_n636), .CI(DP_OP_102J5_124_3590_n785), .CO(
        DP_OP_102J5_124_3590_n617), .S(DP_OP_102J5_124_3590_n618) );
  FADDX1_HVT DP_OP_102J5_124_3590_U423 ( .A(DP_OP_102J5_124_3590_n783), .B(
        DP_OP_102J5_124_3590_n634), .CI(DP_OP_102J5_124_3590_n781), .CO(
        DP_OP_102J5_124_3590_n615), .S(DP_OP_102J5_124_3590_n616) );
  FADDX1_HVT DP_OP_102J5_124_3590_U422 ( .A(DP_OP_102J5_124_3590_n632), .B(
        DP_OP_102J5_124_3590_n779), .CI(DP_OP_102J5_124_3590_n777), .CO(
        DP_OP_102J5_124_3590_n613), .S(DP_OP_102J5_124_3590_n614) );
  FADDX1_HVT DP_OP_102J5_124_3590_U421 ( .A(DP_OP_102J5_124_3590_n630), .B(
        DP_OP_102J5_124_3590_n628), .CI(DP_OP_102J5_124_3590_n775), .CO(
        DP_OP_102J5_124_3590_n611), .S(DP_OP_102J5_124_3590_n612) );
  FADDX1_HVT DP_OP_102J5_124_3590_U420 ( .A(DP_OP_102J5_124_3590_n626), .B(
        DP_OP_102J5_124_3590_n622), .CI(DP_OP_102J5_124_3590_n624), .CO(
        DP_OP_102J5_124_3590_n609), .S(DP_OP_102J5_124_3590_n610) );
  FADDX1_HVT DP_OP_102J5_124_3590_U419 ( .A(DP_OP_102J5_124_3590_n773), .B(
        DP_OP_102J5_124_3590_n771), .CI(DP_OP_102J5_124_3590_n620), .CO(
        DP_OP_102J5_124_3590_n607), .S(DP_OP_102J5_124_3590_n608) );
  FADDX1_HVT DP_OP_102J5_124_3590_U418 ( .A(DP_OP_102J5_124_3590_n618), .B(
        DP_OP_102J5_124_3590_n769), .CI(DP_OP_102J5_124_3590_n767), .CO(
        DP_OP_102J5_124_3590_n605), .S(DP_OP_102J5_124_3590_n606) );
  FADDX1_HVT DP_OP_102J5_124_3590_U417 ( .A(DP_OP_102J5_124_3590_n616), .B(
        DP_OP_102J5_124_3590_n765), .CI(DP_OP_102J5_124_3590_n614), .CO(
        DP_OP_102J5_124_3590_n603), .S(DP_OP_102J5_124_3590_n604) );
  FADDX1_HVT DP_OP_102J5_124_3590_U416 ( .A(DP_OP_102J5_124_3590_n612), .B(
        DP_OP_102J5_124_3590_n763), .CI(DP_OP_102J5_124_3590_n610), .CO(
        DP_OP_102J5_124_3590_n601), .S(DP_OP_102J5_124_3590_n602) );
  FADDX1_HVT DP_OP_102J5_124_3590_U415 ( .A(DP_OP_102J5_124_3590_n761), .B(
        DP_OP_102J5_124_3590_n608), .CI(DP_OP_102J5_124_3590_n759), .CO(
        DP_OP_102J5_124_3590_n599), .S(DP_OP_102J5_124_3590_n600) );
  FADDX1_HVT DP_OP_102J5_124_3590_U414 ( .A(DP_OP_102J5_124_3590_n606), .B(
        DP_OP_102J5_124_3590_n604), .CI(DP_OP_102J5_124_3590_n757), .CO(
        DP_OP_102J5_124_3590_n597), .S(DP_OP_102J5_124_3590_n598) );
  FADDX1_HVT DP_OP_102J5_124_3590_U413 ( .A(DP_OP_102J5_124_3590_n602), .B(
        DP_OP_102J5_124_3590_n755), .CI(DP_OP_102J5_124_3590_n600), .CO(
        DP_OP_102J5_124_3590_n595), .S(DP_OP_102J5_124_3590_n596) );
  FADDX1_HVT DP_OP_102J5_124_3590_U412 ( .A(DP_OP_102J5_124_3590_n753), .B(
        DP_OP_102J5_124_3590_n598), .CI(DP_OP_102J5_124_3590_n596), .CO(
        DP_OP_102J5_124_3590_n593), .S(DP_OP_102J5_124_3590_n594) );
  FADDX1_HVT DP_OP_102J5_124_3590_U411 ( .A(DP_OP_102J5_124_3590_n1917), .B(
        DP_OP_102J5_124_3590_n2357), .CI(DP_OP_102J5_124_3590_n1508), .CO(
        DP_OP_102J5_124_3590_n591), .S(DP_OP_102J5_124_3590_n592) );
  FADDX1_HVT DP_OP_102J5_124_3590_U410 ( .A(DP_OP_102J5_124_3590_n749), .B(
        DP_OP_102J5_124_3590_n1596), .CI(DP_OP_102J5_124_3590_n1522), .CO(
        DP_OP_102J5_124_3590_n589), .S(DP_OP_102J5_124_3590_n590) );
  FADDX1_HVT DP_OP_102J5_124_3590_U409 ( .A(DP_OP_102J5_124_3590_n1772), .B(
        DP_OP_102J5_124_3590_n1552), .CI(DP_OP_102J5_124_3590_n1610), .CO(
        DP_OP_102J5_124_3590_n587), .S(DP_OP_102J5_124_3590_n588) );
  FADDX1_HVT DP_OP_102J5_124_3590_U408 ( .A(DP_OP_102J5_124_3590_n2137), .B(
        DP_OP_102J5_124_3590_n1829), .CI(DP_OP_102J5_124_3590_n1684), .CO(
        DP_OP_102J5_124_3590_n585), .S(DP_OP_102J5_124_3590_n586) );
  FADDX1_HVT DP_OP_102J5_124_3590_U407 ( .A(DP_OP_102J5_124_3590_n1873), .B(
        DP_OP_102J5_124_3590_n1786), .CI(DP_OP_102J5_124_3590_n1859), .CO(
        DP_OP_102J5_124_3590_n583), .S(DP_OP_102J5_124_3590_n584) );
  FADDX1_HVT DP_OP_102J5_124_3590_U406 ( .A(DP_OP_102J5_124_3590_n1903), .B(
        DP_OP_102J5_124_3590_n1815), .CI(DP_OP_102J5_124_3590_n1961), .CO(
        DP_OP_102J5_124_3590_n581), .S(DP_OP_102J5_124_3590_n582) );
  FADDX1_HVT DP_OP_102J5_124_3590_U405 ( .A(DP_OP_102J5_124_3590_n1566), .B(
        DP_OP_102J5_124_3590_n1640), .CI(DP_OP_102J5_124_3590_n1742), .CO(
        DP_OP_102J5_124_3590_n579), .S(DP_OP_102J5_124_3590_n580) );
  FADDX1_HVT DP_OP_102J5_124_3590_U404 ( .A(DP_OP_102J5_124_3590_n1947), .B(
        DP_OP_102J5_124_3590_n2035), .CI(DP_OP_102J5_124_3590_n2005), .CO(
        DP_OP_102J5_124_3590_n577), .S(DP_OP_102J5_124_3590_n578) );
  FADDX1_HVT DP_OP_102J5_124_3590_U403 ( .A(DP_OP_102J5_124_3590_n2181), .B(
        DP_OP_102J5_124_3590_n2079), .CI(DP_OP_102J5_124_3590_n1698), .CO(
        DP_OP_102J5_124_3590_n575), .S(DP_OP_102J5_124_3590_n576) );
  FADDX1_HVT DP_OP_102J5_124_3590_U402 ( .A(DP_OP_102J5_124_3590_n2123), .B(
        DP_OP_102J5_124_3590_n2167), .CI(DP_OP_102J5_124_3590_n2049), .CO(
        DP_OP_102J5_124_3590_n573), .S(DP_OP_102J5_124_3590_n574) );
  FADDX1_HVT DP_OP_102J5_124_3590_U401 ( .A(DP_OP_102J5_124_3590_n2093), .B(
        DP_OP_102J5_124_3590_n1728), .CI(DP_OP_102J5_124_3590_n2225), .CO(
        DP_OP_102J5_124_3590_n571), .S(DP_OP_102J5_124_3590_n572) );
  FADDX1_HVT DP_OP_102J5_124_3590_U400 ( .A(DP_OP_102J5_124_3590_n2269), .B(
        DP_OP_102J5_124_3590_n1991), .CI(DP_OP_102J5_124_3590_n1654), .CO(
        DP_OP_102J5_124_3590_n569), .S(DP_OP_102J5_124_3590_n570) );
  FADDX1_HVT DP_OP_102J5_124_3590_U399 ( .A(DP_OP_102J5_124_3590_n2313), .B(
        DP_OP_102J5_124_3590_n2299), .CI(DP_OP_102J5_124_3590_n2211), .CO(
        DP_OP_102J5_124_3590_n567), .S(DP_OP_102J5_124_3590_n568) );
  FADDX1_HVT DP_OP_102J5_124_3590_U398 ( .A(DP_OP_102J5_124_3590_n2255), .B(
        DP_OP_102J5_124_3590_n2343), .CI(DP_OP_102J5_124_3590_n1779), .CO(
        DP_OP_102J5_124_3590_n565), .S(DP_OP_102J5_124_3590_n566) );
  FADDX1_HVT DP_OP_102J5_124_3590_U397 ( .A(DP_OP_102J5_124_3590_n1691), .B(
        DP_OP_102J5_124_3590_n1515), .CI(DP_OP_102J5_124_3590_n1559), .CO(
        DP_OP_102J5_124_3590_n563), .S(DP_OP_102J5_124_3590_n564) );
  FADDX1_HVT DP_OP_102J5_124_3590_U396 ( .A(DP_OP_102J5_124_3590_n2350), .B(
        DP_OP_102J5_124_3590_n1603), .CI(DP_OP_102J5_124_3590_n1647), .CO(
        DP_OP_102J5_124_3590_n561), .S(DP_OP_102J5_124_3590_n562) );
  FADDX1_HVT DP_OP_102J5_124_3590_U395 ( .A(DP_OP_102J5_124_3590_n2306), .B(
        DP_OP_102J5_124_3590_n1735), .CI(DP_OP_102J5_124_3590_n1822), .CO(
        DP_OP_102J5_124_3590_n559), .S(DP_OP_102J5_124_3590_n560) );
  FADDX1_HVT DP_OP_102J5_124_3590_U394 ( .A(DP_OP_102J5_124_3590_n2262), .B(
        DP_OP_102J5_124_3590_n1866), .CI(DP_OP_102J5_124_3590_n1910), .CO(
        DP_OP_102J5_124_3590_n557), .S(DP_OP_102J5_124_3590_n558) );
  FADDX1_HVT DP_OP_102J5_124_3590_U393 ( .A(DP_OP_102J5_124_3590_n2218), .B(
        DP_OP_102J5_124_3590_n1954), .CI(DP_OP_102J5_124_3590_n1998), .CO(
        DP_OP_102J5_124_3590_n555), .S(DP_OP_102J5_124_3590_n556) );
  FADDX1_HVT DP_OP_102J5_124_3590_U392 ( .A(DP_OP_102J5_124_3590_n2174), .B(
        DP_OP_102J5_124_3590_n2042), .CI(DP_OP_102J5_124_3590_n2086), .CO(
        DP_OP_102J5_124_3590_n553), .S(DP_OP_102J5_124_3590_n554) );
  FADDX1_HVT DP_OP_102J5_124_3590_U391 ( .A(DP_OP_102J5_124_3590_n2130), .B(
        DP_OP_102J5_124_3590_n731), .CI(DP_OP_102J5_124_3590_n733), .CO(
        DP_OP_102J5_124_3590_n551), .S(DP_OP_102J5_124_3590_n552) );
  FADDX1_HVT DP_OP_102J5_124_3590_U390 ( .A(DP_OP_102J5_124_3590_n723), .B(
        DP_OP_102J5_124_3590_n727), .CI(DP_OP_102J5_124_3590_n725), .CO(
        DP_OP_102J5_124_3590_n549), .S(DP_OP_102J5_124_3590_n550) );
  FADDX1_HVT DP_OP_102J5_124_3590_U389 ( .A(DP_OP_102J5_124_3590_n741), .B(
        DP_OP_102J5_124_3590_n729), .CI(DP_OP_102J5_124_3590_n735), .CO(
        DP_OP_102J5_124_3590_n547), .S(DP_OP_102J5_124_3590_n548) );
  FADDX1_HVT DP_OP_102J5_124_3590_U388 ( .A(DP_OP_102J5_124_3590_n743), .B(
        DP_OP_102J5_124_3590_n737), .CI(DP_OP_102J5_124_3590_n745), .CO(
        DP_OP_102J5_124_3590_n545), .S(DP_OP_102J5_124_3590_n546) );
  FADDX1_HVT DP_OP_102J5_124_3590_U387 ( .A(DP_OP_102J5_124_3590_n747), .B(
        DP_OP_102J5_124_3590_n739), .CI(DP_OP_102J5_124_3590_n709), .CO(
        DP_OP_102J5_124_3590_n543), .S(DP_OP_102J5_124_3590_n544) );
  FADDX1_HVT DP_OP_102J5_124_3590_U386 ( .A(DP_OP_102J5_124_3590_n705), .B(
        DP_OP_102J5_124_3590_n699), .CI(DP_OP_102J5_124_3590_n697), .CO(
        DP_OP_102J5_124_3590_n541), .S(DP_OP_102J5_124_3590_n542) );
  FADDX1_HVT DP_OP_102J5_124_3590_U385 ( .A(DP_OP_102J5_124_3590_n707), .B(
        DP_OP_102J5_124_3590_n701), .CI(DP_OP_102J5_124_3590_n711), .CO(
        DP_OP_102J5_124_3590_n539), .S(DP_OP_102J5_124_3590_n540) );
  FADDX1_HVT DP_OP_102J5_124_3590_U384 ( .A(DP_OP_102J5_124_3590_n717), .B(
        DP_OP_102J5_124_3590_n703), .CI(DP_OP_102J5_124_3590_n715), .CO(
        DP_OP_102J5_124_3590_n537), .S(DP_OP_102J5_124_3590_n538) );
  FADDX1_HVT DP_OP_102J5_124_3590_U383 ( .A(DP_OP_102J5_124_3590_n719), .B(
        DP_OP_102J5_124_3590_n721), .CI(DP_OP_102J5_124_3590_n713), .CO(
        DP_OP_102J5_124_3590_n535), .S(DP_OP_102J5_124_3590_n536) );
  FADDX1_HVT DP_OP_102J5_124_3590_U382 ( .A(DP_OP_102J5_124_3590_n586), .B(
        DP_OP_102J5_124_3590_n582), .CI(DP_OP_102J5_124_3590_n566), .CO(
        DP_OP_102J5_124_3590_n533), .S(DP_OP_102J5_124_3590_n534) );
  FADDX1_HVT DP_OP_102J5_124_3590_U381 ( .A(DP_OP_102J5_124_3590_n588), .B(
        DP_OP_102J5_124_3590_n580), .CI(DP_OP_102J5_124_3590_n572), .CO(
        DP_OP_102J5_124_3590_n531), .S(DP_OP_102J5_124_3590_n532) );
  FADDX1_HVT DP_OP_102J5_124_3590_U380 ( .A(DP_OP_102J5_124_3590_n584), .B(
        DP_OP_102J5_124_3590_n568), .CI(DP_OP_102J5_124_3590_n576), .CO(
        DP_OP_102J5_124_3590_n529), .S(DP_OP_102J5_124_3590_n530) );
  FADDX1_HVT DP_OP_102J5_124_3590_U379 ( .A(DP_OP_102J5_124_3590_n574), .B(
        DP_OP_102J5_124_3590_n570), .CI(DP_OP_102J5_124_3590_n578), .CO(
        DP_OP_102J5_124_3590_n527), .S(DP_OP_102J5_124_3590_n528) );
  FADDX1_HVT DP_OP_102J5_124_3590_U378 ( .A(DP_OP_102J5_124_3590_n590), .B(
        DP_OP_102J5_124_3590_n592), .CI(DP_OP_102J5_124_3590_n562), .CO(
        DP_OP_102J5_124_3590_n525), .S(DP_OP_102J5_124_3590_n526) );
  FADDX1_HVT DP_OP_102J5_124_3590_U377 ( .A(DP_OP_102J5_124_3590_n556), .B(
        DP_OP_102J5_124_3590_n564), .CI(DP_OP_102J5_124_3590_n560), .CO(
        DP_OP_102J5_124_3590_n523), .S(DP_OP_102J5_124_3590_n524) );
  FADDX1_HVT DP_OP_102J5_124_3590_U376 ( .A(DP_OP_102J5_124_3590_n554), .B(
        DP_OP_102J5_124_3590_n558), .CI(DP_OP_102J5_124_3590_n695), .CO(
        DP_OP_102J5_124_3590_n521), .S(DP_OP_102J5_124_3590_n522) );
  FADDX1_HVT DP_OP_102J5_124_3590_U375 ( .A(DP_OP_102J5_124_3590_n691), .B(
        DP_OP_102J5_124_3590_n693), .CI(DP_OP_102J5_124_3590_n679), .CO(
        DP_OP_102J5_124_3590_n519), .S(DP_OP_102J5_124_3590_n520) );
  FADDX1_HVT DP_OP_102J5_124_3590_U374 ( .A(DP_OP_102J5_124_3590_n685), .B(
        DP_OP_102J5_124_3590_n681), .CI(DP_OP_102J5_124_3590_n1473), .CO(
        DP_OP_102J5_124_3590_n517), .S(DP_OP_102J5_124_3590_n518) );
  FADDX1_HVT DP_OP_102J5_124_3590_U373 ( .A(DP_OP_102J5_124_3590_n687), .B(
        DP_OP_102J5_124_3590_n689), .CI(DP_OP_102J5_124_3590_n677), .CO(
        DP_OP_102J5_124_3590_n515), .S(DP_OP_102J5_124_3590_n516) );
  FADDX1_HVT DP_OP_102J5_124_3590_U372 ( .A(DP_OP_102J5_124_3590_n683), .B(
        DP_OP_102J5_124_3590_n552), .CI(DP_OP_102J5_124_3590_n675), .CO(
        DP_OP_102J5_124_3590_n513), .S(DP_OP_102J5_124_3590_n514) );
  FADDX1_HVT DP_OP_102J5_124_3590_U371 ( .A(DP_OP_102J5_124_3590_n548), .B(
        DP_OP_102J5_124_3590_n673), .CI(DP_OP_102J5_124_3590_n544), .CO(
        DP_OP_102J5_124_3590_n511), .S(DP_OP_102J5_124_3590_n512) );
  FADDX1_HVT DP_OP_102J5_124_3590_U370 ( .A(DP_OP_102J5_124_3590_n546), .B(
        DP_OP_102J5_124_3590_n671), .CI(DP_OP_102J5_124_3590_n669), .CO(
        DP_OP_102J5_124_3590_n509), .S(DP_OP_102J5_124_3590_n510) );
  FADDX1_HVT DP_OP_102J5_124_3590_U369 ( .A(DP_OP_102J5_124_3590_n550), .B(
        DP_OP_102J5_124_3590_n540), .CI(DP_OP_102J5_124_3590_n667), .CO(
        DP_OP_102J5_124_3590_n507), .S(DP_OP_102J5_124_3590_n508) );
  FADDX1_HVT DP_OP_102J5_124_3590_U368 ( .A(DP_OP_102J5_124_3590_n665), .B(
        DP_OP_102J5_124_3590_n538), .CI(DP_OP_102J5_124_3590_n536), .CO(
        DP_OP_102J5_124_3590_n505), .S(DP_OP_102J5_124_3590_n506) );
  FADDX1_HVT DP_OP_102J5_124_3590_U367 ( .A(DP_OP_102J5_124_3590_n663), .B(
        DP_OP_102J5_124_3590_n542), .CI(DP_OP_102J5_124_3590_n661), .CO(
        DP_OP_102J5_124_3590_n503), .S(DP_OP_102J5_124_3590_n504) );
  FADDX1_HVT DP_OP_102J5_124_3590_U366 ( .A(DP_OP_102J5_124_3590_n530), .B(
        DP_OP_102J5_124_3590_n526), .CI(DP_OP_102J5_124_3590_n659), .CO(
        DP_OP_102J5_124_3590_n501), .S(DP_OP_102J5_124_3590_n502) );
  FADDX1_HVT DP_OP_102J5_124_3590_U365 ( .A(DP_OP_102J5_124_3590_n528), .B(
        DP_OP_102J5_124_3590_n534), .CI(DP_OP_102J5_124_3590_n532), .CO(
        DP_OP_102J5_124_3590_n499), .S(DP_OP_102J5_124_3590_n500) );
  FADDX1_HVT DP_OP_102J5_124_3590_U364 ( .A(DP_OP_102J5_124_3590_n524), .B(
        DP_OP_102J5_124_3590_n522), .CI(DP_OP_102J5_124_3590_n657), .CO(
        DP_OP_102J5_124_3590_n497), .S(DP_OP_102J5_124_3590_n498) );
  FADDX1_HVT DP_OP_102J5_124_3590_U363 ( .A(DP_OP_102J5_124_3590_n655), .B(
        DP_OP_102J5_124_3590_n653), .CI(DP_OP_102J5_124_3590_n651), .CO(
        DP_OP_102J5_124_3590_n495), .S(DP_OP_102J5_124_3590_n496) );
  FADDX1_HVT DP_OP_102J5_124_3590_U362 ( .A(DP_OP_102J5_124_3590_n520), .B(
        DP_OP_102J5_124_3590_n649), .CI(DP_OP_102J5_124_3590_n647), .CO(
        DP_OP_102J5_124_3590_n493), .S(DP_OP_102J5_124_3590_n494) );
  FADDX1_HVT DP_OP_102J5_124_3590_U361 ( .A(DP_OP_102J5_124_3590_n645), .B(
        DP_OP_102J5_124_3590_n516), .CI(DP_OP_102J5_124_3590_n514), .CO(
        DP_OP_102J5_124_3590_n491), .S(DP_OP_102J5_124_3590_n492) );
  FADDX1_HVT DP_OP_102J5_124_3590_U360 ( .A(DP_OP_102J5_124_3590_n643), .B(
        DP_OP_102J5_124_3590_n518), .CI(DP_OP_102J5_124_3590_n641), .CO(
        DP_OP_102J5_124_3590_n489), .S(DP_OP_102J5_124_3590_n490) );
  FADDX1_HVT DP_OP_102J5_124_3590_U359 ( .A(DP_OP_102J5_124_3590_n639), .B(
        DP_OP_102J5_124_3590_n512), .CI(DP_OP_102J5_124_3590_n508), .CO(
        DP_OP_102J5_124_3590_n487), .S(DP_OP_102J5_124_3590_n488) );
  FADDX1_HVT DP_OP_102J5_124_3590_U358 ( .A(DP_OP_102J5_124_3590_n510), .B(
        DP_OP_102J5_124_3590_n637), .CI(DP_OP_102J5_124_3590_n635), .CO(
        DP_OP_102J5_124_3590_n485), .S(DP_OP_102J5_124_3590_n486) );
  FADDX1_HVT DP_OP_102J5_124_3590_U357 ( .A(DP_OP_102J5_124_3590_n506), .B(
        DP_OP_102J5_124_3590_n504), .CI(DP_OP_102J5_124_3590_n633), .CO(
        DP_OP_102J5_124_3590_n483), .S(DP_OP_102J5_124_3590_n484) );
  FADDX1_HVT DP_OP_102J5_124_3590_U356 ( .A(DP_OP_102J5_124_3590_n500), .B(
        DP_OP_102J5_124_3590_n502), .CI(DP_OP_102J5_124_3590_n631), .CO(
        DP_OP_102J5_124_3590_n481), .S(DP_OP_102J5_124_3590_n482) );
  FADDX1_HVT DP_OP_102J5_124_3590_U355 ( .A(DP_OP_102J5_124_3590_n498), .B(
        DP_OP_102J5_124_3590_n629), .CI(DP_OP_102J5_124_3590_n627), .CO(
        DP_OP_102J5_124_3590_n479), .S(DP_OP_102J5_124_3590_n480) );
  FADDX1_HVT DP_OP_102J5_124_3590_U354 ( .A(DP_OP_102J5_124_3590_n496), .B(
        DP_OP_102J5_124_3590_n625), .CI(DP_OP_102J5_124_3590_n494), .CO(
        DP_OP_102J5_124_3590_n477), .S(DP_OP_102J5_124_3590_n478) );
  FADDX1_HVT DP_OP_102J5_124_3590_U353 ( .A(DP_OP_102J5_124_3590_n623), .B(
        DP_OP_102J5_124_3590_n492), .CI(DP_OP_102J5_124_3590_n490), .CO(
        DP_OP_102J5_124_3590_n475), .S(DP_OP_102J5_124_3590_n476) );
  FADDX1_HVT DP_OP_102J5_124_3590_U352 ( .A(DP_OP_102J5_124_3590_n621), .B(
        DP_OP_102J5_124_3590_n619), .CI(DP_OP_102J5_124_3590_n488), .CO(
        DP_OP_102J5_124_3590_n473), .S(DP_OP_102J5_124_3590_n474) );
  FADDX1_HVT DP_OP_102J5_124_3590_U351 ( .A(DP_OP_102J5_124_3590_n486), .B(
        DP_OP_102J5_124_3590_n617), .CI(DP_OP_102J5_124_3590_n484), .CO(
        DP_OP_102J5_124_3590_n471), .S(DP_OP_102J5_124_3590_n472) );
  FADDX1_HVT DP_OP_102J5_124_3590_U350 ( .A(DP_OP_102J5_124_3590_n615), .B(
        DP_OP_102J5_124_3590_n482), .CI(DP_OP_102J5_124_3590_n613), .CO(
        DP_OP_102J5_124_3590_n469), .S(DP_OP_102J5_124_3590_n470) );
  FADDX1_HVT DP_OP_102J5_124_3590_U349 ( .A(DP_OP_102J5_124_3590_n480), .B(
        DP_OP_102J5_124_3590_n611), .CI(DP_OP_102J5_124_3590_n478), .CO(
        DP_OP_102J5_124_3590_n467), .S(DP_OP_102J5_124_3590_n468) );
  FADDX1_HVT DP_OP_102J5_124_3590_U348 ( .A(DP_OP_102J5_124_3590_n609), .B(
        DP_OP_102J5_124_3590_n476), .CI(DP_OP_102J5_124_3590_n607), .CO(
        DP_OP_102J5_124_3590_n465), .S(DP_OP_102J5_124_3590_n466) );
  FADDX1_HVT DP_OP_102J5_124_3590_U347 ( .A(DP_OP_102J5_124_3590_n474), .B(
        DP_OP_102J5_124_3590_n472), .CI(DP_OP_102J5_124_3590_n605), .CO(
        DP_OP_102J5_124_3590_n463), .S(DP_OP_102J5_124_3590_n464) );
  FADDX1_HVT DP_OP_102J5_124_3590_U346 ( .A(DP_OP_102J5_124_3590_n470), .B(
        DP_OP_102J5_124_3590_n603), .CI(DP_OP_102J5_124_3590_n468), .CO(
        DP_OP_102J5_124_3590_n461), .S(DP_OP_102J5_124_3590_n462) );
  FADDX1_HVT DP_OP_102J5_124_3590_U345 ( .A(DP_OP_102J5_124_3590_n601), .B(
        DP_OP_102J5_124_3590_n466), .CI(DP_OP_102J5_124_3590_n599), .CO(
        DP_OP_102J5_124_3590_n459), .S(DP_OP_102J5_124_3590_n460) );
  FADDX1_HVT DP_OP_102J5_124_3590_U344 ( .A(DP_OP_102J5_124_3590_n464), .B(
        DP_OP_102J5_124_3590_n597), .CI(DP_OP_102J5_124_3590_n462), .CO(
        DP_OP_102J5_124_3590_n457), .S(DP_OP_102J5_124_3590_n458) );
  FADDX1_HVT DP_OP_102J5_124_3590_U343 ( .A(DP_OP_102J5_124_3590_n595), .B(
        DP_OP_102J5_124_3590_n460), .CI(DP_OP_102J5_124_3590_n458), .CO(
        DP_OP_102J5_124_3590_n455), .S(DP_OP_102J5_124_3590_n456) );
  FADDX1_HVT DP_OP_102J5_124_3590_U341 ( .A(DP_OP_102J5_124_3590_n1778), .B(
        DP_OP_102J5_124_3590_n2349), .CI(DP_OP_102J5_124_3590_n1507), .CO(
        DP_OP_102J5_124_3590_n451), .S(DP_OP_102J5_124_3590_n452) );
  FADDX1_HVT DP_OP_102J5_124_3590_U340 ( .A(DP_OP_102J5_124_3590_n1771), .B(
        DP_OP_102J5_124_3590_n1514), .CI(DP_OP_102J5_124_3590_n2342), .CO(
        DP_OP_102J5_124_3590_n449), .S(DP_OP_102J5_124_3590_n450) );
  FADDX1_HVT DP_OP_102J5_124_3590_U339 ( .A(DP_OP_102J5_124_3590_n1821), .B(
        DP_OP_102J5_124_3590_n1551), .CI(DP_OP_102J5_124_3590_n1558), .CO(
        DP_OP_102J5_124_3590_n447), .S(DP_OP_102J5_124_3590_n448) );
  FADDX1_HVT DP_OP_102J5_124_3590_U338 ( .A(DP_OP_102J5_124_3590_n1683), .B(
        DP_OP_102J5_124_3590_n2305), .CI(DP_OP_102J5_124_3590_n2298), .CO(
        DP_OP_102J5_124_3590_n445), .S(DP_OP_102J5_124_3590_n446) );
  FADDX1_HVT DP_OP_102J5_124_3590_U337 ( .A(DP_OP_102J5_124_3590_n1639), .B(
        DP_OP_102J5_124_3590_n1595), .CI(DP_OP_102J5_124_3590_n1602), .CO(
        DP_OP_102J5_124_3590_n443), .S(DP_OP_102J5_124_3590_n444) );
  FADDX1_HVT DP_OP_102J5_124_3590_U336 ( .A(DP_OP_102J5_124_3590_n2261), .B(
        DP_OP_102J5_124_3590_n2254), .CI(DP_OP_102J5_124_3590_n2217), .CO(
        DP_OP_102J5_124_3590_n441), .S(DP_OP_102J5_124_3590_n442) );
  FADDX1_HVT DP_OP_102J5_124_3590_U335 ( .A(DP_OP_102J5_124_3590_n1990), .B(
        DP_OP_102J5_124_3590_n2210), .CI(DP_OP_102J5_124_3590_n2173), .CO(
        DP_OP_102J5_124_3590_n439), .S(DP_OP_102J5_124_3590_n440) );
  FADDX1_HVT DP_OP_102J5_124_3590_U334 ( .A(DP_OP_102J5_124_3590_n1902), .B(
        DP_OP_102J5_124_3590_n1646), .CI(DP_OP_102J5_124_3590_n2166), .CO(
        DP_OP_102J5_124_3590_n437), .S(DP_OP_102J5_124_3590_n438) );
  FADDX1_HVT DP_OP_102J5_124_3590_U333 ( .A(DP_OP_102J5_124_3590_n1865), .B(
        DP_OP_102J5_124_3590_n1690), .CI(DP_OP_102J5_124_3590_n1727), .CO(
        DP_OP_102J5_124_3590_n435), .S(DP_OP_102J5_124_3590_n436) );
  FADDX1_HVT DP_OP_102J5_124_3590_U332 ( .A(DP_OP_102J5_124_3590_n2129), .B(
        DP_OP_102J5_124_3590_n2122), .CI(DP_OP_102J5_124_3590_n1734), .CO(
        DP_OP_102J5_124_3590_n433), .S(DP_OP_102J5_124_3590_n434) );
  FADDX1_HVT DP_OP_102J5_124_3590_U331 ( .A(DP_OP_102J5_124_3590_n1953), .B(
        DP_OP_102J5_124_3590_n2085), .CI(DP_OP_102J5_124_3590_n2078), .CO(
        DP_OP_102J5_124_3590_n431), .S(DP_OP_102J5_124_3590_n432) );
  FADDX1_HVT DP_OP_102J5_124_3590_U330 ( .A(DP_OP_102J5_124_3590_n2041), .B(
        DP_OP_102J5_124_3590_n1858), .CI(DP_OP_102J5_124_3590_n1909), .CO(
        DP_OP_102J5_124_3590_n429), .S(DP_OP_102J5_124_3590_n430) );
  FADDX1_HVT DP_OP_102J5_124_3590_U329 ( .A(DP_OP_102J5_124_3590_n2034), .B(
        DP_OP_102J5_124_3590_n1946), .CI(DP_OP_102J5_124_3590_n1997), .CO(
        DP_OP_102J5_124_3590_n427), .S(DP_OP_102J5_124_3590_n428) );
  FADDX1_HVT DP_OP_102J5_124_3590_U328 ( .A(DP_OP_102J5_124_3590_n454), .B(
        DP_OP_102J5_124_3590_n565), .CI(DP_OP_102J5_124_3590_n581), .CO(
        DP_OP_102J5_124_3590_n425), .S(DP_OP_102J5_124_3590_n426) );
  FADDX1_HVT DP_OP_102J5_124_3590_U327 ( .A(DP_OP_102J5_124_3590_n575), .B(
        DP_OP_102J5_124_3590_n569), .CI(DP_OP_102J5_124_3590_n571), .CO(
        DP_OP_102J5_124_3590_n423), .S(DP_OP_102J5_124_3590_n424) );
  FADDX1_HVT DP_OP_102J5_124_3590_U326 ( .A(DP_OP_102J5_124_3590_n577), .B(
        DP_OP_102J5_124_3590_n567), .CI(DP_OP_102J5_124_3590_n579), .CO(
        DP_OP_102J5_124_3590_n421), .S(DP_OP_102J5_124_3590_n422) );
  FADDX1_HVT DP_OP_102J5_124_3590_U325 ( .A(DP_OP_102J5_124_3590_n587), .B(
        DP_OP_102J5_124_3590_n573), .CI(DP_OP_102J5_124_3590_n585), .CO(
        DP_OP_102J5_124_3590_n419), .S(DP_OP_102J5_124_3590_n420) );
  FADDX1_HVT DP_OP_102J5_124_3590_U324 ( .A(DP_OP_102J5_124_3590_n589), .B(
        DP_OP_102J5_124_3590_n591), .CI(DP_OP_102J5_124_3590_n583), .CO(
        DP_OP_102J5_124_3590_n417), .S(DP_OP_102J5_124_3590_n418) );
  FADDX1_HVT DP_OP_102J5_124_3590_U323 ( .A(DP_OP_102J5_124_3590_n553), .B(
        DP_OP_102J5_124_3590_n555), .CI(DP_OP_102J5_124_3590_n559), .CO(
        DP_OP_102J5_124_3590_n415), .S(DP_OP_102J5_124_3590_n416) );
  FADDX1_HVT DP_OP_102J5_124_3590_U322 ( .A(DP_OP_102J5_124_3590_n561), .B(
        DP_OP_102J5_124_3590_n557), .CI(DP_OP_102J5_124_3590_n563), .CO(
        DP_OP_102J5_124_3590_n413), .S(DP_OP_102J5_124_3590_n414) );
  FADDX1_HVT DP_OP_102J5_124_3590_U321 ( .A(DP_OP_102J5_124_3590_n428), .B(
        DP_OP_102J5_124_3590_n452), .CI(DP_OP_102J5_124_3590_n450), .CO(
        DP_OP_102J5_124_3590_n411), .S(DP_OP_102J5_124_3590_n412) );
  FADDX1_HVT DP_OP_102J5_124_3590_U320 ( .A(DP_OP_102J5_124_3590_n430), .B(
        DP_OP_102J5_124_3590_n446), .CI(DP_OP_102J5_124_3590_n438), .CO(
        DP_OP_102J5_124_3590_n409), .S(DP_OP_102J5_124_3590_n410) );
  FADDX1_HVT DP_OP_102J5_124_3590_U319 ( .A(DP_OP_102J5_124_3590_n440), .B(
        DP_OP_102J5_124_3590_n436), .CI(DP_OP_102J5_124_3590_n432), .CO(
        DP_OP_102J5_124_3590_n407), .S(DP_OP_102J5_124_3590_n408) );
  FADDX1_HVT DP_OP_102J5_124_3590_U318 ( .A(DP_OP_102J5_124_3590_n434), .B(
        DP_OP_102J5_124_3590_n448), .CI(DP_OP_102J5_124_3590_n444), .CO(
        DP_OP_102J5_124_3590_n405), .S(DP_OP_102J5_124_3590_n406) );
  FADDX1_HVT DP_OP_102J5_124_3590_U317 ( .A(DP_OP_102J5_124_3590_n442), .B(
        DP_OP_102J5_124_3590_n551), .CI(DP_OP_102J5_124_3590_n547), .CO(
        DP_OP_102J5_124_3590_n403), .S(DP_OP_102J5_124_3590_n404) );
  FADDX1_HVT DP_OP_102J5_124_3590_U316 ( .A(DP_OP_102J5_124_3590_n545), .B(
        DP_OP_102J5_124_3590_n549), .CI(DP_OP_102J5_124_3590_n543), .CO(
        DP_OP_102J5_124_3590_n401), .S(DP_OP_102J5_124_3590_n402) );
  FADDX1_HVT DP_OP_102J5_124_3590_U315 ( .A(DP_OP_102J5_124_3590_n539), .B(
        DP_OP_102J5_124_3590_n535), .CI(DP_OP_102J5_124_3590_n1472), .CO(
        DP_OP_102J5_124_3590_n399), .S(DP_OP_102J5_124_3590_n400) );
  FADDX1_HVT DP_OP_102J5_124_3590_U314 ( .A(DP_OP_102J5_124_3590_n541), .B(
        DP_OP_102J5_124_3590_n537), .CI(DP_OP_102J5_124_3590_n426), .CO(
        DP_OP_102J5_124_3590_n397), .S(DP_OP_102J5_124_3590_n398) );
  FADDX1_HVT DP_OP_102J5_124_3590_U313 ( .A(DP_OP_102J5_124_3590_n420), .B(
        DP_OP_102J5_124_3590_n424), .CI(DP_OP_102J5_124_3590_n418), .CO(
        DP_OP_102J5_124_3590_n395), .S(DP_OP_102J5_124_3590_n396) );
  FADDX1_HVT DP_OP_102J5_124_3590_U312 ( .A(DP_OP_102J5_124_3590_n533), .B(
        DP_OP_102J5_124_3590_n422), .CI(DP_OP_102J5_124_3590_n525), .CO(
        DP_OP_102J5_124_3590_n393), .S(DP_OP_102J5_124_3590_n394) );
  FADDX1_HVT DP_OP_102J5_124_3590_U311 ( .A(DP_OP_102J5_124_3590_n531), .B(
        DP_OP_102J5_124_3590_n527), .CI(DP_OP_102J5_124_3590_n529), .CO(
        DP_OP_102J5_124_3590_n391), .S(DP_OP_102J5_124_3590_n392) );
  FADDX1_HVT DP_OP_102J5_124_3590_U310 ( .A(DP_OP_102J5_124_3590_n416), .B(
        DP_OP_102J5_124_3590_n414), .CI(DP_OP_102J5_124_3590_n521), .CO(
        DP_OP_102J5_124_3590_n389), .S(DP_OP_102J5_124_3590_n390) );
  FADDX1_HVT DP_OP_102J5_124_3590_U309 ( .A(DP_OP_102J5_124_3590_n523), .B(
        DP_OP_102J5_124_3590_n408), .CI(DP_OP_102J5_124_3590_n410), .CO(
        DP_OP_102J5_124_3590_n387), .S(DP_OP_102J5_124_3590_n388) );
  FADDX1_HVT DP_OP_102J5_124_3590_U308 ( .A(DP_OP_102J5_124_3590_n406), .B(
        DP_OP_102J5_124_3590_n412), .CI(DP_OP_102J5_124_3590_n519), .CO(
        DP_OP_102J5_124_3590_n385), .S(DP_OP_102J5_124_3590_n386) );
  FADDX1_HVT DP_OP_102J5_124_3590_U307 ( .A(DP_OP_102J5_124_3590_n517), .B(
        DP_OP_102J5_124_3590_n515), .CI(DP_OP_102J5_124_3590_n404), .CO(
        DP_OP_102J5_124_3590_n383), .S(DP_OP_102J5_124_3590_n384) );
  FADDX1_HVT DP_OP_102J5_124_3590_U306 ( .A(DP_OP_102J5_124_3590_n513), .B(
        DP_OP_102J5_124_3590_n511), .CI(DP_OP_102J5_124_3590_n402), .CO(
        DP_OP_102J5_124_3590_n381), .S(DP_OP_102J5_124_3590_n382) );
  FADDX1_HVT DP_OP_102J5_124_3590_U305 ( .A(DP_OP_102J5_124_3590_n509), .B(
        DP_OP_102J5_124_3590_n507), .CI(DP_OP_102J5_124_3590_n505), .CO(
        DP_OP_102J5_124_3590_n379), .S(DP_OP_102J5_124_3590_n380) );
  FADDX1_HVT DP_OP_102J5_124_3590_U304 ( .A(DP_OP_102J5_124_3590_n400), .B(
        DP_OP_102J5_124_3590_n503), .CI(DP_OP_102J5_124_3590_n398), .CO(
        DP_OP_102J5_124_3590_n377), .S(DP_OP_102J5_124_3590_n378) );
  FADDX1_HVT DP_OP_102J5_124_3590_U303 ( .A(DP_OP_102J5_124_3590_n501), .B(
        DP_OP_102J5_124_3590_n394), .CI(DP_OP_102J5_124_3590_n396), .CO(
        DP_OP_102J5_124_3590_n375), .S(DP_OP_102J5_124_3590_n376) );
  FADDX1_HVT DP_OP_102J5_124_3590_U302 ( .A(DP_OP_102J5_124_3590_n499), .B(
        DP_OP_102J5_124_3590_n392), .CI(DP_OP_102J5_124_3590_n390), .CO(
        DP_OP_102J5_124_3590_n373), .S(DP_OP_102J5_124_3590_n374) );
  FADDX1_HVT DP_OP_102J5_124_3590_U301 ( .A(DP_OP_102J5_124_3590_n497), .B(
        DP_OP_102J5_124_3590_n388), .CI(DP_OP_102J5_124_3590_n495), .CO(
        DP_OP_102J5_124_3590_n371), .S(DP_OP_102J5_124_3590_n372) );
  FADDX1_HVT DP_OP_102J5_124_3590_U300 ( .A(DP_OP_102J5_124_3590_n386), .B(
        DP_OP_102J5_124_3590_n493), .CI(DP_OP_102J5_124_3590_n491), .CO(
        DP_OP_102J5_124_3590_n369), .S(DP_OP_102J5_124_3590_n370) );
  FADDX1_HVT DP_OP_102J5_124_3590_U299 ( .A(DP_OP_102J5_124_3590_n489), .B(
        DP_OP_102J5_124_3590_n384), .CI(DP_OP_102J5_124_3590_n382), .CO(
        DP_OP_102J5_124_3590_n367), .S(DP_OP_102J5_124_3590_n368) );
  FADDX1_HVT DP_OP_102J5_124_3590_U298 ( .A(DP_OP_102J5_124_3590_n487), .B(
        DP_OP_102J5_124_3590_n485), .CI(DP_OP_102J5_124_3590_n380), .CO(
        DP_OP_102J5_124_3590_n365), .S(DP_OP_102J5_124_3590_n366) );
  FADDX1_HVT DP_OP_102J5_124_3590_U297 ( .A(DP_OP_102J5_124_3590_n378), .B(
        DP_OP_102J5_124_3590_n483), .CI(DP_OP_102J5_124_3590_n481), .CO(
        DP_OP_102J5_124_3590_n363), .S(DP_OP_102J5_124_3590_n364) );
  FADDX1_HVT DP_OP_102J5_124_3590_U296 ( .A(DP_OP_102J5_124_3590_n376), .B(
        DP_OP_102J5_124_3590_n374), .CI(DP_OP_102J5_124_3590_n479), .CO(
        DP_OP_102J5_124_3590_n361), .S(DP_OP_102J5_124_3590_n362) );
  FADDX1_HVT DP_OP_102J5_124_3590_U295 ( .A(DP_OP_102J5_124_3590_n372), .B(
        DP_OP_102J5_124_3590_n477), .CI(DP_OP_102J5_124_3590_n370), .CO(
        DP_OP_102J5_124_3590_n359), .S(DP_OP_102J5_124_3590_n360) );
  FADDX1_HVT DP_OP_102J5_124_3590_U294 ( .A(DP_OP_102J5_124_3590_n475), .B(
        DP_OP_102J5_124_3590_n368), .CI(DP_OP_102J5_124_3590_n473), .CO(
        DP_OP_102J5_124_3590_n357), .S(DP_OP_102J5_124_3590_n358) );
  FADDX1_HVT DP_OP_102J5_124_3590_U293 ( .A(DP_OP_102J5_124_3590_n366), .B(
        DP_OP_102J5_124_3590_n471), .CI(DP_OP_102J5_124_3590_n364), .CO(
        DP_OP_102J5_124_3590_n355), .S(DP_OP_102J5_124_3590_n356) );
  FADDX1_HVT DP_OP_102J5_124_3590_U292 ( .A(DP_OP_102J5_124_3590_n469), .B(
        DP_OP_102J5_124_3590_n362), .CI(DP_OP_102J5_124_3590_n467), .CO(
        DP_OP_102J5_124_3590_n353), .S(DP_OP_102J5_124_3590_n354) );
  FADDX1_HVT DP_OP_102J5_124_3590_U291 ( .A(DP_OP_102J5_124_3590_n360), .B(
        DP_OP_102J5_124_3590_n465), .CI(DP_OP_102J5_124_3590_n358), .CO(
        DP_OP_102J5_124_3590_n351), .S(DP_OP_102J5_124_3590_n352) );
  FADDX1_HVT DP_OP_102J5_124_3590_U290 ( .A(DP_OP_102J5_124_3590_n463), .B(
        DP_OP_102J5_124_3590_n356), .CI(DP_OP_102J5_124_3590_n461), .CO(
        DP_OP_102J5_124_3590_n349), .S(DP_OP_102J5_124_3590_n350) );
  FADDX1_HVT DP_OP_102J5_124_3590_U289 ( .A(DP_OP_102J5_124_3590_n354), .B(
        DP_OP_102J5_124_3590_n352), .CI(DP_OP_102J5_124_3590_n459), .CO(
        DP_OP_102J5_124_3590_n347), .S(DP_OP_102J5_124_3590_n348) );
  FADDX1_HVT DP_OP_102J5_124_3590_U288 ( .A(DP_OP_102J5_124_3590_n457), .B(
        DP_OP_102J5_124_3590_n350), .CI(DP_OP_102J5_124_3590_n348), .CO(
        DP_OP_102J5_124_3590_n345), .S(DP_OP_102J5_124_3590_n346) );
  FADDX1_HVT DP_OP_102J5_124_3590_U287 ( .A(DP_OP_102J5_124_3590_n453), .B(
        DP_OP_102J5_124_3590_n2341), .CI(DP_OP_102J5_124_3590_n2297), .CO(
        DP_OP_102J5_124_3590_n270), .S(DP_OP_102J5_124_3590_n344) );
  FADDX1_HVT DP_OP_102J5_124_3590_U286 ( .A(DP_OP_102J5_124_3590_n1945), .B(
        DP_OP_102J5_124_3590_n2253), .CI(DP_OP_102J5_124_3590_n1506), .CO(
        DP_OP_102J5_124_3590_n342), .S(DP_OP_102J5_124_3590_n343) );
  FADDX1_HVT DP_OP_102J5_124_3590_U285 ( .A(DP_OP_102J5_124_3590_n1857), .B(
        DP_OP_102J5_124_3590_n2209), .CI(DP_OP_102J5_124_3590_n1550), .CO(
        DP_OP_102J5_124_3590_n340), .S(DP_OP_102J5_124_3590_n341) );
  FADDX1_HVT DP_OP_102J5_124_3590_U284 ( .A(DP_OP_102J5_124_3590_n1770), .B(
        DP_OP_102J5_124_3590_n2165), .CI(DP_OP_102J5_124_3590_n2121), .CO(
        DP_OP_102J5_124_3590_n338), .S(DP_OP_102J5_124_3590_n339) );
  FADDX1_HVT DP_OP_102J5_124_3590_U283 ( .A(DP_OP_102J5_124_3590_n2077), .B(
        DP_OP_102J5_124_3590_n2033), .CI(DP_OP_102J5_124_3590_n1989), .CO(
        DP_OP_102J5_124_3590_n336), .S(DP_OP_102J5_124_3590_n337) );
  FADDX1_HVT DP_OP_102J5_124_3590_U282 ( .A(DP_OP_102J5_124_3590_n1682), .B(
        DP_OP_102J5_124_3590_n1594), .CI(DP_OP_102J5_124_3590_n1638), .CO(
        DP_OP_102J5_124_3590_n334), .S(DP_OP_102J5_124_3590_n335) );
  FADDX1_HVT DP_OP_102J5_124_3590_U281 ( .A(DP_OP_102J5_124_3590_n1814), .B(
        DP_OP_102J5_124_3590_n1901), .CI(DP_OP_102J5_124_3590_n1726), .CO(
        DP_OP_102J5_124_3590_n332), .S(DP_OP_102J5_124_3590_n333) );
  FADDX1_HVT DP_OP_102J5_124_3590_U280 ( .A(DP_OP_102J5_124_3590_n439), .B(
        DP_OP_102J5_124_3590_n429), .CI(DP_OP_102J5_124_3590_n427), .CO(
        DP_OP_102J5_124_3590_n330), .S(DP_OP_102J5_124_3590_n331) );
  FADDX1_HVT DP_OP_102J5_124_3590_U279 ( .A(DP_OP_102J5_124_3590_n443), .B(
        DP_OP_102J5_124_3590_n431), .CI(DP_OP_102J5_124_3590_n435), .CO(
        DP_OP_102J5_124_3590_n328), .S(DP_OP_102J5_124_3590_n329) );
  FADDX1_HVT DP_OP_102J5_124_3590_U278 ( .A(DP_OP_102J5_124_3590_n445), .B(
        DP_OP_102J5_124_3590_n433), .CI(DP_OP_102J5_124_3590_n437), .CO(
        DP_OP_102J5_124_3590_n326), .S(DP_OP_102J5_124_3590_n327) );
  FADDX1_HVT DP_OP_102J5_124_3590_U277 ( .A(DP_OP_102J5_124_3590_n441), .B(
        DP_OP_102J5_124_3590_n447), .CI(DP_OP_102J5_124_3590_n449), .CO(
        DP_OP_102J5_124_3590_n324), .S(DP_OP_102J5_124_3590_n325) );
  FADDX1_HVT DP_OP_102J5_124_3590_U276 ( .A(DP_OP_102J5_124_3590_n451), .B(
        DP_OP_102J5_124_3590_n344), .CI(DP_OP_102J5_124_3590_n339), .CO(
        DP_OP_102J5_124_3590_n322), .S(DP_OP_102J5_124_3590_n323) );
  FADDX1_HVT DP_OP_102J5_124_3590_U275 ( .A(DP_OP_102J5_124_3590_n341), .B(
        DP_OP_102J5_124_3590_n333), .CI(DP_OP_102J5_124_3590_n335), .CO(
        DP_OP_102J5_124_3590_n320), .S(DP_OP_102J5_124_3590_n321) );
  FADDX1_HVT DP_OP_102J5_124_3590_U274 ( .A(DP_OP_102J5_124_3590_n337), .B(
        DP_OP_102J5_124_3590_n343), .CI(DP_OP_102J5_124_3590_n425), .CO(
        DP_OP_102J5_124_3590_n318), .S(DP_OP_102J5_124_3590_n319) );
  FADDX1_HVT DP_OP_102J5_124_3590_U273 ( .A(DP_OP_102J5_124_3590_n417), .B(
        DP_OP_102J5_124_3590_n419), .CI(DP_OP_102J5_124_3590_n421), .CO(
        DP_OP_102J5_124_3590_n316), .S(DP_OP_102J5_124_3590_n317) );
  FADDX1_HVT DP_OP_102J5_124_3590_U272 ( .A(DP_OP_102J5_124_3590_n423), .B(
        DP_OP_102J5_124_3590_n415), .CI(DP_OP_102J5_124_3590_n413), .CO(
        DP_OP_102J5_124_3590_n314), .S(DP_OP_102J5_124_3590_n315) );
  FADDX1_HVT DP_OP_102J5_124_3590_U271 ( .A(DP_OP_102J5_124_3590_n1471), .B(
        DP_OP_102J5_124_3590_n411), .CI(DP_OP_102J5_124_3590_n409), .CO(
        DP_OP_102J5_124_3590_n312), .S(DP_OP_102J5_124_3590_n313) );
  FADDX1_HVT DP_OP_102J5_124_3590_U270 ( .A(DP_OP_102J5_124_3590_n407), .B(
        DP_OP_102J5_124_3590_n327), .CI(DP_OP_102J5_124_3590_n325), .CO(
        DP_OP_102J5_124_3590_n310), .S(DP_OP_102J5_124_3590_n311) );
  FADDX1_HVT DP_OP_102J5_124_3590_U269 ( .A(DP_OP_102J5_124_3590_n405), .B(
        DP_OP_102J5_124_3590_n329), .CI(DP_OP_102J5_124_3590_n331), .CO(
        DP_OP_102J5_124_3590_n308), .S(DP_OP_102J5_124_3590_n309) );
  FADDX1_HVT DP_OP_102J5_124_3590_U268 ( .A(DP_OP_102J5_124_3590_n403), .B(
        DP_OP_102J5_124_3590_n323), .CI(DP_OP_102J5_124_3590_n321), .CO(
        DP_OP_102J5_124_3590_n306), .S(DP_OP_102J5_124_3590_n307) );
  FADDX1_HVT DP_OP_102J5_124_3590_U267 ( .A(DP_OP_102J5_124_3590_n401), .B(
        DP_OP_102J5_124_3590_n399), .CI(DP_OP_102J5_124_3590_n397), .CO(
        DP_OP_102J5_124_3590_n304), .S(DP_OP_102J5_124_3590_n305) );
  FADDX1_HVT DP_OP_102J5_124_3590_U266 ( .A(DP_OP_102J5_124_3590_n319), .B(
        DP_OP_102J5_124_3590_n395), .CI(DP_OP_102J5_124_3590_n393), .CO(
        DP_OP_102J5_124_3590_n302), .S(DP_OP_102J5_124_3590_n303) );
  FADDX1_HVT DP_OP_102J5_124_3590_U265 ( .A(DP_OP_102J5_124_3590_n391), .B(
        DP_OP_102J5_124_3590_n317), .CI(DP_OP_102J5_124_3590_n315), .CO(
        DP_OP_102J5_124_3590_n300), .S(DP_OP_102J5_124_3590_n301) );
  FADDX1_HVT DP_OP_102J5_124_3590_U264 ( .A(DP_OP_102J5_124_3590_n389), .B(
        DP_OP_102J5_124_3590_n387), .CI(DP_OP_102J5_124_3590_n313), .CO(
        DP_OP_102J5_124_3590_n298), .S(DP_OP_102J5_124_3590_n299) );
  FADDX1_HVT DP_OP_102J5_124_3590_U263 ( .A(DP_OP_102J5_124_3590_n311), .B(
        DP_OP_102J5_124_3590_n309), .CI(DP_OP_102J5_124_3590_n385), .CO(
        DP_OP_102J5_124_3590_n296), .S(DP_OP_102J5_124_3590_n297) );
  FADDX1_HVT DP_OP_102J5_124_3590_U262 ( .A(DP_OP_102J5_124_3590_n383), .B(
        DP_OP_102J5_124_3590_n307), .CI(DP_OP_102J5_124_3590_n381), .CO(
        DP_OP_102J5_124_3590_n294), .S(DP_OP_102J5_124_3590_n295) );
  FADDX1_HVT DP_OP_102J5_124_3590_U261 ( .A(DP_OP_102J5_124_3590_n379), .B(
        DP_OP_102J5_124_3590_n305), .CI(DP_OP_102J5_124_3590_n377), .CO(
        DP_OP_102J5_124_3590_n292), .S(DP_OP_102J5_124_3590_n293) );
  FADDX1_HVT DP_OP_102J5_124_3590_U260 ( .A(DP_OP_102J5_124_3590_n303), .B(
        DP_OP_102J5_124_3590_n373), .CI(DP_OP_102J5_124_3590_n301), .CO(
        DP_OP_102J5_124_3590_n290), .S(DP_OP_102J5_124_3590_n291) );
  FADDX1_HVT DP_OP_102J5_124_3590_U259 ( .A(DP_OP_102J5_124_3590_n375), .B(
        DP_OP_102J5_124_3590_n371), .CI(DP_OP_102J5_124_3590_n299), .CO(
        DP_OP_102J5_124_3590_n288), .S(DP_OP_102J5_124_3590_n289) );
  FADDX1_HVT DP_OP_102J5_124_3590_U258 ( .A(DP_OP_102J5_124_3590_n297), .B(
        DP_OP_102J5_124_3590_n369), .CI(DP_OP_102J5_124_3590_n367), .CO(
        DP_OP_102J5_124_3590_n286), .S(DP_OP_102J5_124_3590_n287) );
  FADDX1_HVT DP_OP_102J5_124_3590_U257 ( .A(DP_OP_102J5_124_3590_n295), .B(
        DP_OP_102J5_124_3590_n365), .CI(DP_OP_102J5_124_3590_n293), .CO(
        DP_OP_102J5_124_3590_n284), .S(DP_OP_102J5_124_3590_n285) );
  FADDX1_HVT DP_OP_102J5_124_3590_U256 ( .A(DP_OP_102J5_124_3590_n363), .B(
        DP_OP_102J5_124_3590_n291), .CI(DP_OP_102J5_124_3590_n361), .CO(
        DP_OP_102J5_124_3590_n282), .S(DP_OP_102J5_124_3590_n283) );
  FADDX1_HVT DP_OP_102J5_124_3590_U255 ( .A(DP_OP_102J5_124_3590_n289), .B(
        DP_OP_102J5_124_3590_n359), .CI(DP_OP_102J5_124_3590_n287), .CO(
        DP_OP_102J5_124_3590_n280), .S(DP_OP_102J5_124_3590_n281) );
  FADDX1_HVT DP_OP_102J5_124_3590_U254 ( .A(DP_OP_102J5_124_3590_n357), .B(
        DP_OP_102J5_124_3590_n285), .CI(DP_OP_102J5_124_3590_n355), .CO(
        DP_OP_102J5_124_3590_n278), .S(DP_OP_102J5_124_3590_n279) );
  FADDX1_HVT DP_OP_102J5_124_3590_U253 ( .A(DP_OP_102J5_124_3590_n283), .B(
        DP_OP_102J5_124_3590_n353), .CI(DP_OP_102J5_124_3590_n281), .CO(
        DP_OP_102J5_124_3590_n276), .S(DP_OP_102J5_124_3590_n277) );
  FADDX1_HVT DP_OP_102J5_124_3590_U252 ( .A(DP_OP_102J5_124_3590_n351), .B(
        DP_OP_102J5_124_3590_n279), .CI(DP_OP_102J5_124_3590_n349), .CO(
        DP_OP_102J5_124_3590_n274), .S(DP_OP_102J5_124_3590_n275) );
  FADDX1_HVT DP_OP_102J5_124_3590_U251 ( .A(DP_OP_102J5_124_3590_n277), .B(
        DP_OP_102J5_124_3590_n347), .CI(DP_OP_102J5_124_3590_n275), .CO(
        DP_OP_102J5_124_3590_n272), .S(DP_OP_102J5_124_3590_n273) );
  FADDX1_HVT DP_OP_102J5_124_3590_U249 ( .A(DP_OP_102J5_124_3590_n336), .B(
        DP_OP_102J5_124_3590_n332), .CI(DP_OP_102J5_124_3590_n271), .CO(
        DP_OP_102J5_124_3590_n268), .S(DP_OP_102J5_124_3590_n269) );
  FADDX1_HVT DP_OP_102J5_124_3590_U248 ( .A(DP_OP_102J5_124_3590_n338), .B(
        DP_OP_102J5_124_3590_n340), .CI(DP_OP_102J5_124_3590_n334), .CO(
        DP_OP_102J5_124_3590_n266), .S(DP_OP_102J5_124_3590_n267) );
  FADDX1_HVT DP_OP_102J5_124_3590_U247 ( .A(DP_OP_102J5_124_3590_n342), .B(
        DP_OP_102J5_124_3590_n326), .CI(DP_OP_102J5_124_3590_n324), .CO(
        DP_OP_102J5_124_3590_n264), .S(DP_OP_102J5_124_3590_n265) );
  FADDX1_HVT DP_OP_102J5_124_3590_U246 ( .A(DP_OP_102J5_124_3590_n330), .B(
        DP_OP_102J5_124_3590_n328), .CI(DP_OP_102J5_124_3590_n1470), .CO(
        DP_OP_102J5_124_3590_n262), .S(DP_OP_102J5_124_3590_n263) );
  FADDX1_HVT DP_OP_102J5_124_3590_U245 ( .A(DP_OP_102J5_124_3590_n322), .B(
        DP_OP_102J5_124_3590_n320), .CI(DP_OP_102J5_124_3590_n267), .CO(
        DP_OP_102J5_124_3590_n260), .S(DP_OP_102J5_124_3590_n261) );
  FADDX1_HVT DP_OP_102J5_124_3590_U244 ( .A(DP_OP_102J5_124_3590_n269), .B(
        DP_OP_102J5_124_3590_n318), .CI(DP_OP_102J5_124_3590_n316), .CO(
        DP_OP_102J5_124_3590_n258), .S(DP_OP_102J5_124_3590_n259) );
  FADDX1_HVT DP_OP_102J5_124_3590_U243 ( .A(DP_OP_102J5_124_3590_n314), .B(
        DP_OP_102J5_124_3590_n312), .CI(DP_OP_102J5_124_3590_n265), .CO(
        DP_OP_102J5_124_3590_n256), .S(DP_OP_102J5_124_3590_n257) );
  FADDX1_HVT DP_OP_102J5_124_3590_U242 ( .A(DP_OP_102J5_124_3590_n310), .B(
        DP_OP_102J5_124_3590_n308), .CI(DP_OP_102J5_124_3590_n263), .CO(
        DP_OP_102J5_124_3590_n254), .S(DP_OP_102J5_124_3590_n255) );
  FADDX1_HVT DP_OP_102J5_124_3590_U241 ( .A(DP_OP_102J5_124_3590_n306), .B(
        DP_OP_102J5_124_3590_n261), .CI(DP_OP_102J5_124_3590_n304), .CO(
        DP_OP_102J5_124_3590_n252), .S(DP_OP_102J5_124_3590_n253) );
  FADDX1_HVT DP_OP_102J5_124_3590_U240 ( .A(DP_OP_102J5_124_3590_n259), .B(
        DP_OP_102J5_124_3590_n302), .CI(DP_OP_102J5_124_3590_n300), .CO(
        DP_OP_102J5_124_3590_n250), .S(DP_OP_102J5_124_3590_n251) );
  FADDX1_HVT DP_OP_102J5_124_3590_U239 ( .A(DP_OP_102J5_124_3590_n298), .B(
        DP_OP_102J5_124_3590_n257), .CI(DP_OP_102J5_124_3590_n296), .CO(
        DP_OP_102J5_124_3590_n248), .S(DP_OP_102J5_124_3590_n249) );
  FADDX1_HVT DP_OP_102J5_124_3590_U238 ( .A(DP_OP_102J5_124_3590_n255), .B(
        DP_OP_102J5_124_3590_n294), .CI(DP_OP_102J5_124_3590_n253), .CO(
        DP_OP_102J5_124_3590_n246), .S(DP_OP_102J5_124_3590_n247) );
  FADDX1_HVT DP_OP_102J5_124_3590_U237 ( .A(DP_OP_102J5_124_3590_n292), .B(
        DP_OP_102J5_124_3590_n251), .CI(DP_OP_102J5_124_3590_n290), .CO(
        DP_OP_102J5_124_3590_n244), .S(DP_OP_102J5_124_3590_n245) );
  FADDX1_HVT DP_OP_102J5_124_3590_U236 ( .A(DP_OP_102J5_124_3590_n288), .B(
        DP_OP_102J5_124_3590_n249), .CI(DP_OP_102J5_124_3590_n286), .CO(
        DP_OP_102J5_124_3590_n242), .S(DP_OP_102J5_124_3590_n243) );
  FADDX1_HVT DP_OP_102J5_124_3590_U235 ( .A(DP_OP_102J5_124_3590_n247), .B(
        DP_OP_102J5_124_3590_n284), .CI(DP_OP_102J5_124_3590_n245), .CO(
        DP_OP_102J5_124_3590_n240), .S(DP_OP_102J5_124_3590_n241) );
  FADDX1_HVT DP_OP_102J5_124_3590_U234 ( .A(DP_OP_102J5_124_3590_n282), .B(
        DP_OP_102J5_124_3590_n280), .CI(DP_OP_102J5_124_3590_n243), .CO(
        DP_OP_102J5_124_3590_n238), .S(DP_OP_102J5_124_3590_n239) );
  FADDX1_HVT DP_OP_102J5_124_3590_U233 ( .A(DP_OP_102J5_124_3590_n278), .B(
        DP_OP_102J5_124_3590_n241), .CI(DP_OP_102J5_124_3590_n276), .CO(
        DP_OP_102J5_124_3590_n236), .S(DP_OP_102J5_124_3590_n237) );
  FADDX1_HVT DP_OP_102J5_124_3590_U232 ( .A(DP_OP_102J5_124_3590_n239), .B(
        DP_OP_102J5_124_3590_n274), .CI(DP_OP_102J5_124_3590_n237), .CO(
        DP_OP_102J5_124_3590_n234), .S(DP_OP_102J5_124_3590_n235) );
  FADDX1_HVT DP_OP_102J5_124_3590_U231 ( .A(DP_OP_102J5_124_3590_n270), .B(
        DP_OP_102J5_124_3590_n268), .CI(DP_OP_102J5_124_3590_n266), .CO(
        DP_OP_102J5_124_3590_n232), .S(DP_OP_102J5_124_3590_n233) );
  FADDX1_HVT DP_OP_102J5_124_3590_U230 ( .A(DP_OP_102J5_124_3590_n1469), .B(
        DP_OP_102J5_124_3590_n264), .CI(DP_OP_102J5_124_3590_n262), .CO(
        DP_OP_102J5_124_3590_n230), .S(DP_OP_102J5_124_3590_n231) );
  FADDX1_HVT DP_OP_102J5_124_3590_U229 ( .A(DP_OP_102J5_124_3590_n260), .B(
        DP_OP_102J5_124_3590_n233), .CI(DP_OP_102J5_124_3590_n258), .CO(
        DP_OP_102J5_124_3590_n228), .S(DP_OP_102J5_124_3590_n229) );
  FADDX1_HVT DP_OP_102J5_124_3590_U228 ( .A(DP_OP_102J5_124_3590_n256), .B(
        DP_OP_102J5_124_3590_n231), .CI(DP_OP_102J5_124_3590_n254), .CO(
        DP_OP_102J5_124_3590_n226), .S(DP_OP_102J5_124_3590_n227) );
  FADDX1_HVT DP_OP_102J5_124_3590_U227 ( .A(DP_OP_102J5_124_3590_n252), .B(
        DP_OP_102J5_124_3590_n229), .CI(DP_OP_102J5_124_3590_n250), .CO(
        DP_OP_102J5_124_3590_n224), .S(DP_OP_102J5_124_3590_n225) );
  FADDX1_HVT DP_OP_102J5_124_3590_U226 ( .A(DP_OP_102J5_124_3590_n248), .B(
        DP_OP_102J5_124_3590_n227), .CI(DP_OP_102J5_124_3590_n246), .CO(
        DP_OP_102J5_124_3590_n222), .S(DP_OP_102J5_124_3590_n223) );
  FADDX1_HVT DP_OP_102J5_124_3590_U225 ( .A(DP_OP_102J5_124_3590_n225), .B(
        DP_OP_102J5_124_3590_n244), .CI(DP_OP_102J5_124_3590_n242), .CO(
        DP_OP_102J5_124_3590_n220), .S(DP_OP_102J5_124_3590_n221) );
  FADDX1_HVT DP_OP_102J5_124_3590_U224 ( .A(DP_OP_102J5_124_3590_n223), .B(
        DP_OP_102J5_124_3590_n240), .CI(DP_OP_102J5_124_3590_n221), .CO(
        DP_OP_102J5_124_3590_n218), .S(DP_OP_102J5_124_3590_n219) );
  FADDX1_HVT DP_OP_102J5_124_3590_U223 ( .A(DP_OP_102J5_124_3590_n238), .B(
        DP_OP_102J5_124_3590_n236), .CI(DP_OP_102J5_124_3590_n219), .CO(
        DP_OP_102J5_124_3590_n216), .S(DP_OP_102J5_124_3590_n217) );
  FADDX1_HVT DP_OP_102J5_124_3590_U221 ( .A(DP_OP_102J5_124_3590_n215), .B(
        DP_OP_102J5_124_3590_n232), .CI(DP_OP_102J5_124_3590_n230), .CO(
        DP_OP_102J5_124_3590_n212), .S(DP_OP_102J5_124_3590_n213) );
  FADDX1_HVT DP_OP_102J5_124_3590_U220 ( .A(DP_OP_102J5_124_3590_n228), .B(
        DP_OP_102J5_124_3590_n213), .CI(DP_OP_102J5_124_3590_n226), .CO(
        DP_OP_102J5_124_3590_n210), .S(DP_OP_102J5_124_3590_n211) );
  FADDX1_HVT DP_OP_102J5_124_3590_U219 ( .A(DP_OP_102J5_124_3590_n224), .B(
        DP_OP_102J5_124_3590_n211), .CI(DP_OP_102J5_124_3590_n222), .CO(
        DP_OP_102J5_124_3590_n208), .S(DP_OP_102J5_124_3590_n209) );
  FADDX1_HVT DP_OP_102J5_124_3590_U218 ( .A(DP_OP_102J5_124_3590_n220), .B(
        DP_OP_102J5_124_3590_n209), .CI(DP_OP_102J5_124_3590_n218), .CO(
        DP_OP_102J5_124_3590_n206), .S(DP_OP_102J5_124_3590_n207) );
  FADDX1_HVT DP_OP_102J5_124_3590_U216 ( .A(DP_OP_102J5_124_3590_n214), .B(
        DP_OP_102J5_124_3590_n205), .CI(DP_OP_102J5_124_3590_n212), .CO(
        DP_OP_102J5_124_3590_n202), .S(DP_OP_102J5_124_3590_n203) );
  FADDX1_HVT DP_OP_102J5_124_3590_U215 ( .A(DP_OP_102J5_124_3590_n203), .B(
        DP_OP_102J5_124_3590_n210), .CI(DP_OP_102J5_124_3590_n208), .CO(
        DP_OP_102J5_124_3590_n200), .S(DP_OP_102J5_124_3590_n201) );
  FADDX1_HVT DP_OP_102J5_124_3590_U214 ( .A(DP_OP_102J5_124_3590_n1468), .B(
        DP_OP_102J5_124_3590_n204), .CI(DP_OP_102J5_124_3590_n202), .CO(
        DP_OP_102J5_124_3590_n198), .S(DP_OP_102J5_124_3590_n199) );
  FADDX1_HVT DP_OP_102J5_124_3590_U206 ( .A(DP_OP_102J5_124_3590_n1454), .B(
        DP_OP_102J5_124_3590_n1452), .CI(DP_OP_102J5_124_3590_n1450), .CO(
        DP_OP_102J5_124_3590_n162), .S(n_accumulator_sum[0]) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U205 ( .A1(DP_OP_102J5_124_3590_n1402), 
        .A2(DP_OP_102J5_124_3590_n1404), .Y(DP_OP_102J5_124_3590_n161) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U204 ( .A1(DP_OP_102J5_124_3590_n1404), .A2(
        DP_OP_102J5_124_3590_n1402), .Y(DP_OP_102J5_124_3590_n160) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U198 ( .A1(DP_OP_102J5_124_3590_n1318), 
        .A2(DP_OP_102J5_124_3590_n1320), .Y(DP_OP_102J5_124_3590_n158) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U189 ( .A1(DP_OP_102J5_124_3590_n1196), 
        .A2(DP_OP_102J5_124_3590_n1198), .Y(DP_OP_102J5_124_3590_n152) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U181 ( .A1(DP_OP_102J5_124_3590_n1056), 
        .A2(DP_OP_102J5_124_3590_n1058), .Y(DP_OP_102J5_124_3590_n147) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U180 ( .A1(DP_OP_102J5_124_3590_n1058), .A2(
        DP_OP_102J5_124_3590_n1056), .Y(DP_OP_102J5_124_3590_n146) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U175 ( .A1(DP_OP_102J5_124_3590_n906), .A2(
        DP_OP_102J5_124_3590_n908), .Y(DP_OP_102J5_124_3590_n144) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U167 ( .A1(DP_OP_102J5_124_3590_n752), .A2(
        DP_OP_102J5_124_3590_n754), .Y(DP_OP_102J5_124_3590_n139) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U154 ( .A1(DP_OP_102J5_124_3590_n456), .A2(
        DP_OP_102J5_124_3590_n593), .Y(DP_OP_102J5_124_3590_n132) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U145 ( .A1(DP_OP_102J5_124_3590_n346), .A2(
        DP_OP_102J5_124_3590_n455), .Y(DP_OP_102J5_124_3590_n126) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U144 ( .A1(DP_OP_102J5_124_3590_n455), .A2(
        DP_OP_102J5_124_3590_n346), .Y(DP_OP_102J5_124_3590_n125) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U137 ( .A1(DP_OP_102J5_124_3590_n273), .A2(
        DP_OP_102J5_124_3590_n345), .Y(DP_OP_102J5_124_3590_n121) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U136 ( .A1(DP_OP_102J5_124_3590_n345), .A2(
        DP_OP_102J5_124_3590_n273), .Y(DP_OP_102J5_124_3590_n120) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U132 ( .A1(DP_OP_102J5_124_3590_n125), .A2(
        DP_OP_102J5_124_3590_n120), .Y(DP_OP_102J5_124_3590_n118) );
  AOI21X1_HVT DP_OP_102J5_124_3590_U131 ( .A1(DP_OP_102J5_124_3590_n127), .A2(
        DP_OP_102J5_124_3590_n118), .A3(DP_OP_102J5_124_3590_n119), .Y(
        DP_OP_102J5_124_3590_n117) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U129 ( .A1(DP_OP_102J5_124_3590_n235), .A2(
        DP_OP_102J5_124_3590_n272), .Y(DP_OP_102J5_124_3590_n116) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U128 ( .A1(DP_OP_102J5_124_3590_n272), .A2(
        DP_OP_102J5_124_3590_n235), .Y(DP_OP_102J5_124_3590_n115) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U123 ( .A1(DP_OP_102J5_124_3590_n217), .A2(
        DP_OP_102J5_124_3590_n234), .Y(DP_OP_102J5_124_3590_n113) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U122 ( .A1(DP_OP_102J5_124_3590_n234), .A2(
        DP_OP_102J5_124_3590_n217), .Y(DP_OP_102J5_124_3590_n112) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U112 ( .A1(DP_OP_102J5_124_3590_n216), .A2(
        DP_OP_102J5_124_3590_n207), .Y(DP_OP_102J5_124_3590_n105) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U111 ( .A1(DP_OP_102J5_124_3590_n207), .A2(
        DP_OP_102J5_124_3590_n216), .Y(DP_OP_102J5_124_3590_n104) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U106 ( .A1(DP_OP_102J5_124_3590_n206), .A2(
        DP_OP_102J5_124_3590_n201), .Y(DP_OP_102J5_124_3590_n98) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U105 ( .A1(DP_OP_102J5_124_3590_n201), .A2(
        DP_OP_102J5_124_3590_n206), .Y(DP_OP_102J5_124_3590_n97) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U97 ( .A1(DP_OP_102J5_124_3590_n97), .A2(
        DP_OP_102J5_124_3590_n104), .Y(DP_OP_102J5_124_3590_n95) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U92 ( .A1(DP_OP_102J5_124_3590_n200), .A2(
        DP_OP_102J5_124_3590_n199), .Y(DP_OP_102J5_124_3590_n91) );
  AOI21X1_HVT DP_OP_102J5_124_3590_U84 ( .A1(DP_OP_102J5_124_3590_n96), .A2(
        n279), .A3(DP_OP_102J5_124_3590_n89), .Y(DP_OP_102J5_124_3590_n85) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U83 ( .A1(DP_OP_102J5_124_3590_n95), .A2(
        n279), .Y(DP_OP_102J5_124_3590_n84) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U78 ( .A1(DP_OP_102J5_124_3590_n198), .A2(
        DP_OP_102J5_124_3590_n197), .Y(DP_OP_102J5_124_3590_n76) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U77 ( .A1(DP_OP_102J5_124_3590_n197), .A2(
        DP_OP_102J5_124_3590_n198), .Y(DP_OP_102J5_124_3590_n75) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U66 ( .A1(DP_OP_102J5_124_3590_n195), .A2(
        DP_OP_102J5_124_3590_n196), .Y(DP_OP_102J5_124_3590_n71) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U59 ( .A1(DP_OP_102J5_124_3590_n77), .A2(
        n291), .Y(DP_OP_102J5_124_3590_n64) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U52 ( .A1(DP_OP_102J5_124_3590_n193), .A2(
        DP_OP_102J5_124_3590_n194), .Y(DP_OP_102J5_124_3590_n60) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U51 ( .A1(DP_OP_102J5_124_3590_n194), .A2(
        DP_OP_102J5_124_3590_n193), .Y(DP_OP_102J5_124_3590_n59) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U45 ( .A1(n279), .A2(
        DP_OP_102J5_124_3590_n57), .Y(DP_OP_102J5_124_3590_n53) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U38 ( .A1(DP_OP_102J5_124_3590_n191), .A2(
        DP_OP_102J5_124_3590_n192), .Y(DP_OP_102J5_124_3590_n49) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U37 ( .A1(DP_OP_102J5_124_3590_n192), .A2(
        DP_OP_102J5_124_3590_n191), .Y(DP_OP_102J5_124_3590_n48) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U31 ( .A1(DP_OP_102J5_124_3590_n99), .A2(
        DP_OP_102J5_124_3590_n46), .Y(DP_OP_102J5_124_3590_n44) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U29 ( .A1(DP_OP_102J5_124_3590_n44), .A2(
        DP_OP_102J5_124_3590_n104), .Y(DP_OP_102J5_124_3590_n42) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U26 ( .A1(DP_OP_102J5_124_3590_n189), .A2(
        DP_OP_102J5_124_3590_n190), .Y(DP_OP_102J5_124_3590_n40) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U19 ( .A1(DP_OP_102J5_124_3590_n42), .A2(
        n290), .Y(DP_OP_102J5_124_3590_n35) );
  NAND2X0_HVT DP_OP_102J5_124_3590_U14 ( .A1(DP_OP_102J5_124_3590_n187), .A2(
        DP_OP_102J5_124_3590_n188), .Y(DP_OP_102J5_124_3590_n31) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U13 ( .A1(DP_OP_102J5_124_3590_n188), .A2(
        DP_OP_102J5_124_3590_n187), .Y(DP_OP_102J5_124_3590_n30) );
  XNOR2X1_HVT DP_OP_102J5_124_3590_U642 ( .A1(DP_OP_102J5_124_3590_n1950), 
        .A2(DP_OP_102J5_124_3590_n2082), .Y(DP_OP_102J5_124_3590_n1054) );
  OAI21X1_HVT DP_OP_102J5_124_3590_U200 ( .A1(DP_OP_102J5_124_3590_n5), .A2(
        DP_OP_102J5_124_3590_n160), .A3(DP_OP_102J5_124_3590_n161), .Y(
        DP_OP_102J5_124_3590_n159) );
  OAI21X1_HVT DP_OP_102J5_124_3590_U177 ( .A1(DP_OP_102J5_124_3590_n148), .A2(
        DP_OP_102J5_124_3590_n146), .A3(DP_OP_102J5_124_3590_n147), .Y(
        DP_OP_102J5_124_3590_n145) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U867 ( .A1(n294), .A2(accumulate_reset), .Y(
        DP_OP_102J5_124_3590_n1476) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U856 ( .A1(n288), .A2(n191), .Y(
        DP_OP_102J5_124_3590_n196) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U855 ( .A1(n196), .A2(n191), .Y(
        DP_OP_102J5_124_3590_n194) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U854 ( .A1(n289), .A2(n191), .Y(
        DP_OP_102J5_124_3590_n192) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U868 ( .A1(n278), .A2(accumulate_reset), .Y(
        DP_OP_102J5_124_3590_n1477) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U853 ( .A1(n299), .A2(n191), .Y(
        DP_OP_102J5_124_3590_n190) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U852 ( .A1(n197), .A2(n191), .Y(
        DP_OP_102J5_124_3590_n188) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U851 ( .A1(n300), .A2(n191), .Y(
        DP_OP_102J5_124_3590_n186) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U872 ( .A1(n283), .A2(accumulate_reset), .Y(
        DP_OP_102J5_124_3590_n1481) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U871 ( .A1(n282), .A2(accumulate_reset), .Y(
        DP_OP_102J5_124_3590_n1480) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U869 ( .A1(n280), .A2(accumulate_reset), .Y(
        DP_OP_102J5_124_3590_n1478) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U870 ( .A1(n281), .A2(accumulate_reset), .Y(
        DP_OP_102J5_124_3590_n1479) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U862 ( .A1(n292), .A2(accumulate_reset), .Y(
        DP_OP_102J5_124_3590_n1471) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U860 ( .A1(n193), .A2(n191), .Y(
        DP_OP_102J5_124_3590_n1469) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U863 ( .A1(n295), .A2(accumulate_reset), .Y(
        DP_OP_102J5_124_3590_n1472) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U864 ( .A1(n195), .A2(accumulate_reset), .Y(
        DP_OP_102J5_124_3590_n1473) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U857 ( .A1(n298), .A2(n191), .Y(
        DP_OP_102J5_124_3590_n1468) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U865 ( .A1(n296), .A2(accumulate_reset), .Y(
        DP_OP_102J5_124_3590_n1474) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U861 ( .A1(n194), .A2(n191), .Y(
        DP_OP_102J5_124_3590_n1470) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U866 ( .A1(n293), .A2(accumulate_reset), .Y(
        DP_OP_102J5_124_3590_n1475) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U47 ( .A1(DP_OP_102J5_124_3590_n59), .A2(
        DP_OP_102J5_124_3590_n64), .Y(DP_OP_102J5_124_3590_n57) );
  OAI21X1_HVT DP_OP_102J5_124_3590_U133 ( .A1(DP_OP_102J5_124_3590_n126), .A2(
        DP_OP_102J5_124_3590_n120), .A3(DP_OP_102J5_124_3590_n121), .Y(
        DP_OP_102J5_124_3590_n119) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U33 ( .A1(DP_OP_102J5_124_3590_n48), .A2(
        DP_OP_102J5_124_3590_n53), .Y(DP_OP_102J5_124_3590_n46) );
  OAI21X1_HVT DP_OP_102J5_124_3590_U98 ( .A1(DP_OP_102J5_124_3590_n97), .A2(
        DP_OP_102J5_124_3590_n105), .A3(DP_OP_102J5_124_3590_n98), .Y(
        DP_OP_102J5_124_3590_n96) );
  NOR2X1_HVT DP_OP_102J5_124_3590_U1230 ( .A1(n241), .A2(
        DP_OP_102J5_124_3590_n1846), .Y(DP_OP_102J5_124_3590_n1838) );
  NOR2X0_HVT DP_OP_102J5_124_3590_U859 ( .A1(n297), .A2(n191), .Y(
        DP_OP_102J5_124_3590_n214) );
  OA221X1_HVT U106 ( .A1(1'b0), .A2(DP_OP_102J5_124_3590_n31), .A3(
        DP_OP_102J5_124_3590_n30), .A4(DP_OP_102J5_124_3590_n36), .A5(n183), 
        .Y(n185) );
  OA221X1_HVT U107 ( .A1(1'b0), .A2(DP_OP_102J5_124_3590_n56), .A3(
        DP_OP_102J5_124_3590_n53), .A4(DP_OP_102J5_124_3590_n94), .A5(n153), 
        .Y(n155) );
  OA221X1_HVT U108 ( .A1(1'b0), .A2(DP_OP_102J5_124_3590_n67), .A3(
        DP_OP_102J5_124_3590_n64), .A4(DP_OP_102J5_124_3590_n85), .A5(n146), 
        .Y(n147) );
  OA221X1_HVT U109 ( .A1(1'b0), .A2(DP_OP_102J5_124_3590_n76), .A3(
        DP_OP_102J5_124_3590_n75), .A4(DP_OP_102J5_124_3590_n85), .A5(n138), 
        .Y(n140) );
  OA221X1_HVT U110 ( .A1(1'b0), .A2(DP_OP_102J5_124_3590_n60), .A3(
        DP_OP_102J5_124_3590_n67), .A4(DP_OP_102J5_124_3590_n59), .A5(n123), 
        .Y(DP_OP_102J5_124_3590_n56) );
  OA221X1_HVT U111 ( .A1(DP_OP_102J5_124_3590_n56), .A2(
        DP_OP_102J5_124_3590_n48), .A3(DP_OP_102J5_124_3590_n98), .A4(n113), 
        .A5(DP_OP_102J5_124_3590_n49), .Y(n114) );
  INVX2_HVT U112 ( .A(n110), .Y(DP_OP_102J5_124_3590_n138) );
  INVX2_HVT U113 ( .A(n107), .Y(DP_OP_102J5_124_3590_n134) );
  INVX2_HVT U114 ( .A(n108), .Y(DP_OP_102J5_124_3590_n131) );
  AND3X1_HVT U115 ( .A1(n106), .A2(DP_OP_102J5_124_3590_n132), .A3(n104), .Y(
        DP_OP_102J5_124_3590_n128) );
  NAND2X0_HVT U116 ( .A1(n105), .A2(n108), .Y(n104) );
  INVX2_HVT U117 ( .A(DP_OP_102J5_124_3590_n135), .Y(n105) );
  NAND2X0_HVT U118 ( .A1(DP_OP_102J5_124_3590_n594), .A2(
        DP_OP_102J5_124_3590_n751), .Y(DP_OP_102J5_124_3590_n135) );
  NAND3X0_HVT U119 ( .A1(DP_OP_102J5_124_3590_n137), .A2(n108), .A3(n107), .Y(
        n106) );
  OR2X1_HVT U120 ( .A1(DP_OP_102J5_124_3590_n751), .A2(
        DP_OP_102J5_124_3590_n594), .Y(n107) );
  OR2X1_HVT U121 ( .A1(DP_OP_102J5_124_3590_n593), .A2(
        DP_OP_102J5_124_3590_n456), .Y(n108) );
  AO21X1_HVT U122 ( .A1(n111), .A2(n110), .A3(n109), .Y(
        DP_OP_102J5_124_3590_n137) );
  INVX2_HVT U123 ( .A(DP_OP_102J5_124_3590_n139), .Y(n109) );
  OR2X1_HVT U124 ( .A1(DP_OP_102J5_124_3590_n754), .A2(
        DP_OP_102J5_124_3590_n752), .Y(n110) );
  INVX2_HVT U125 ( .A(DP_OP_102J5_124_3590_n140), .Y(n111) );
  AND2X1_HVT U126 ( .A1(n112), .A2(DP_OP_102J5_124_3590_n144), .Y(
        DP_OP_102J5_124_3590_n140) );
  NAND2X0_HVT U127 ( .A1(DP_OP_102J5_124_3590_n145), .A2(n286), .Y(n112) );
  INVX0_HVT U128 ( .A(DP_OP_102J5_124_3590_n46), .Y(n113) );
  OAI21X1_HVT U129 ( .A1(DP_OP_102J5_124_3590_n105), .A2(
        DP_OP_102J5_124_3590_n44), .A3(n114), .Y(DP_OP_102J5_124_3590_n43) );
  NOR2X0_HVT U130 ( .A1(DP_OP_102J5_124_3590_n112), .A2(
        DP_OP_102J5_124_3590_n115), .Y(n115) );
  INVX0_HVT U131 ( .A(DP_OP_102J5_124_3590_n128), .Y(n116) );
  NAND3X0_HVT U132 ( .A1(DP_OP_102J5_124_3590_n118), .A2(n115), .A3(n116), .Y(
        n117) );
  NAND2X0_HVT U133 ( .A1(n115), .A2(DP_OP_102J5_124_3590_n119), .Y(n118) );
  OR2X1_HVT U134 ( .A1(DP_OP_102J5_124_3590_n112), .A2(
        DP_OP_102J5_124_3590_n116), .Y(n119) );
  NAND4X0_HVT U135 ( .A1(DP_OP_102J5_124_3590_n113), .A2(n117), .A3(n118), 
        .A4(n119), .Y(DP_OP_102J5_124_3590_n3) );
  INVX0_HVT U136 ( .A(DP_OP_102J5_124_3590_n104), .Y(n120) );
  NAND2X0_HVT U137 ( .A1(n120), .A2(DP_OP_102J5_124_3590_n105), .Y(n121) );
  HADDX1_HVT U138 ( .A0(DP_OP_102J5_124_3590_n106), .B0(n121), .SO(
        n_accumulator_sum[13]) );
  NAND2X0_HVT U140 ( .A1(DP_OP_102J5_124_3590_n57), .A2(
        DP_OP_102J5_124_3590_n89), .Y(n123) );
  AND2X1_HVT U141 ( .A1(DP_OP_102J5_124_3590_n176), .A2(
        DP_OP_102J5_124_3590_n126), .Y(n124) );
  HADDX1_HVT U142 ( .A0(n124), .B0(DP_OP_102J5_124_3590_n127), .SO(
        n_accumulator_sum[9]) );
  OA21X1_HVT U143 ( .A1(DP_OP_102J5_124_3590_n106), .A2(
        DP_OP_102J5_124_3590_n104), .A3(DP_OP_102J5_124_3590_n105), .Y(n125)
         );
  NAND2X0_HVT U144 ( .A1(DP_OP_102J5_124_3590_n99), .A2(
        DP_OP_102J5_124_3590_n98), .Y(n126) );
  HADDX1_HVT U145 ( .A0(n125), .B0(n126), .SO(n_accumulator_sum[14]) );
  INVX0_HVT U146 ( .A(DP_OP_102J5_124_3590_n120), .Y(n127) );
  NAND2X0_HVT U147 ( .A1(DP_OP_102J5_124_3590_n127), .A2(
        DP_OP_102J5_124_3590_n176), .Y(n128) );
  AO22X1_HVT U148 ( .A1(n127), .A2(DP_OP_102J5_124_3590_n121), .A3(
        DP_OP_102J5_124_3590_n126), .A4(n128), .Y(n129) );
  NAND4X0_HVT U149 ( .A1(n127), .A2(DP_OP_102J5_124_3590_n121), .A3(
        DP_OP_102J5_124_3590_n126), .A4(n128), .Y(n130) );
  NAND2X0_HVT U150 ( .A1(n129), .A2(n130), .Y(n_accumulator_sum[10]) );
  OA21X1_HVT U151 ( .A1(DP_OP_102J5_124_3590_n106), .A2(
        DP_OP_102J5_124_3590_n93), .A3(DP_OP_102J5_124_3590_n94), .Y(n131) );
  NAND2X0_HVT U152 ( .A1(n279), .A2(DP_OP_102J5_124_3590_n91), .Y(n132) );
  HADDX1_HVT U153 ( .A0(n131), .B0(n132), .SO(n_accumulator_sum[15]) );
  INVX0_HVT U154 ( .A(DP_OP_102J5_124_3590_n3), .Y(n133) );
  OA21X1_HVT U155 ( .A1(DP_OP_102J5_124_3590_n84), .A2(n133), .A3(
        DP_OP_102J5_124_3590_n85), .Y(n134) );
  NAND2X0_HVT U156 ( .A1(DP_OP_102J5_124_3590_n77), .A2(
        DP_OP_102J5_124_3590_n76), .Y(n135) );
  HADDX1_HVT U157 ( .A0(n134), .B0(n135), .SO(n_accumulator_sum[16]) );
  NAND2X0_HVT U158 ( .A1(DP_OP_102J5_124_3590_n159), .A2(n285), .Y(n136) );
  NAND2X0_HVT U159 ( .A1(DP_OP_102J5_124_3590_n158), .A2(n136), .Y(n192) );
  OR3X1_HVT U160 ( .A1(n137), .A2(DP_OP_102J5_124_3590_n75), .A3(
        DP_OP_102J5_124_3590_n84), .Y(n138) );
  NAND2X0_HVT U162 ( .A1(n291), .A2(DP_OP_102J5_124_3590_n71), .Y(n141) );
  HADDX1_HVT U163 ( .A0(n140), .B0(n141), .SO(n_accumulator_sum[17]) );
  INVX0_HVT U164 ( .A(DP_OP_102J5_124_3590_n3), .Y(n137) );
  NAND2X0_HVT U165 ( .A1(n284), .A2(n192), .Y(n142) );
  AND2X1_HVT U166 ( .A1(n142), .A2(DP_OP_102J5_124_3590_n152), .Y(
        DP_OP_102J5_124_3590_n148) );
  NAND2X0_HVT U167 ( .A1(DP_OP_102J5_124_3590_n43), .A2(n290), .Y(n143) );
  AND2X1_HVT U168 ( .A1(n143), .A2(DP_OP_102J5_124_3590_n40), .Y(
        DP_OP_102J5_124_3590_n36) );
  INVX0_HVT U170 ( .A(DP_OP_102J5_124_3590_n3), .Y(n145) );
  OR3X1_HVT U171 ( .A1(n145), .A2(DP_OP_102J5_124_3590_n64), .A3(
        DP_OP_102J5_124_3590_n84), .Y(n146) );
  INVX0_HVT U172 ( .A(DP_OP_102J5_124_3590_n59), .Y(n148) );
  NAND2X0_HVT U173 ( .A1(n148), .A2(DP_OP_102J5_124_3590_n60), .Y(n149) );
  HADDX1_HVT U174 ( .A0(n147), .B0(n149), .SO(n_accumulator_sum[18]) );
  INVX0_HVT U175 ( .A(DP_OP_102J5_124_3590_n146), .Y(n150) );
  NAND2X0_HVT U176 ( .A1(n150), .A2(DP_OP_102J5_124_3590_n147), .Y(n151) );
  HADDX1_HVT U177 ( .A0(DP_OP_102J5_124_3590_n148), .B0(n151), .SO(
        n_accumulator_sum[4]) );
  OR3X1_HVT U178 ( .A1(n152), .A2(DP_OP_102J5_124_3590_n53), .A3(
        DP_OP_102J5_124_3590_n93), .Y(n153) );
  INVX0_HVT U180 ( .A(DP_OP_102J5_124_3590_n48), .Y(n156) );
  NAND2X0_HVT U181 ( .A1(n156), .A2(DP_OP_102J5_124_3590_n49), .Y(n157) );
  HADDX1_HVT U182 ( .A0(n155), .B0(n157), .SO(n_accumulator_sum[19]) );
  INVX0_HVT U183 ( .A(DP_OP_102J5_124_3590_n3), .Y(n152) );
  INVX0_HVT U184 ( .A(DP_OP_102J5_124_3590_n138), .Y(n158) );
  NAND2X0_HVT U185 ( .A1(n158), .A2(DP_OP_102J5_124_3590_n139), .Y(n159) );
  HADDX1_HVT U186 ( .A0(DP_OP_102J5_124_3590_n140), .B0(n159), .SO(
        n_accumulator_sum[6]) );
  AOI21X1_HVT U187 ( .A1(DP_OP_102J5_124_3590_n3), .A2(
        DP_OP_102J5_124_3590_n42), .A3(DP_OP_102J5_124_3590_n43), .Y(n160) );
  NAND2X0_HVT U188 ( .A1(DP_OP_102J5_124_3590_n40), .A2(n290), .Y(n161) );
  HADDX1_HVT U189 ( .A0(n160), .B0(n161), .SO(n_accumulator_sum[20]) );
  AND2X1_HVT U190 ( .A1(DP_OP_102J5_124_3590_n158), .A2(n285), .Y(n162) );
  HADDX1_HVT U191 ( .A0(n162), .B0(DP_OP_102J5_124_3590_n159), .SO(
        n_accumulator_sum[2]) );
  INVX0_HVT U192 ( .A(DP_OP_102J5_124_3590_n134), .Y(n163) );
  NAND2X0_HVT U193 ( .A1(n163), .A2(DP_OP_102J5_124_3590_n135), .Y(n164) );
  HADDX1_HVT U194 ( .A0(DP_OP_102J5_124_3590_n136), .B0(n164), .SO(
        n_accumulator_sum[7]) );
  INVX0_HVT U195 ( .A(DP_OP_102J5_124_3590_n115), .Y(n165) );
  NAND2X0_HVT U196 ( .A1(n165), .A2(DP_OP_102J5_124_3590_n116), .Y(n166) );
  HADDX1_HVT U197 ( .A0(DP_OP_102J5_124_3590_n117), .B0(n166), .SO(
        n_accumulator_sum[11]) );
  INVX0_HVT U198 ( .A(DP_OP_102J5_124_3590_n3), .Y(n167) );
  OA21X1_HVT U199 ( .A1(DP_OP_102J5_124_3590_n35), .A2(n167), .A3(
        DP_OP_102J5_124_3590_n36), .Y(n168) );
  INVX0_HVT U200 ( .A(DP_OP_102J5_124_3590_n30), .Y(n169) );
  NAND2X0_HVT U201 ( .A1(n169), .A2(DP_OP_102J5_124_3590_n31), .Y(n170) );
  HADDX1_HVT U202 ( .A0(n168), .B0(n170), .SO(n_accumulator_sum[21]) );
  INVX0_HVT U203 ( .A(n291), .Y(n171) );
  OA21X1_HVT U204 ( .A1(DP_OP_102J5_124_3590_n76), .A2(n171), .A3(
        DP_OP_102J5_124_3590_n71), .Y(DP_OP_102J5_124_3590_n67) );
  INVX0_HVT U205 ( .A(DP_OP_102J5_124_3590_n160), .Y(n172) );
  AND2X1_HVT U206 ( .A1(n172), .A2(DP_OP_102J5_124_3590_n161), .Y(n173) );
  HADDX1_HVT U207 ( .A0(n173), .B0(DP_OP_102J5_124_3590_n162), .SO(
        n_accumulator_sum[1]) );
  AND2X1_HVT U208 ( .A1(DP_OP_102J5_124_3590_n152), .A2(n284), .Y(n174) );
  HADDX1_HVT U209 ( .A0(n174), .B0(n192), .SO(n_accumulator_sum[3]) );
  AND2X1_HVT U210 ( .A1(DP_OP_102J5_124_3590_n144), .A2(n286), .Y(n175) );
  HADDX1_HVT U211 ( .A0(n175), .B0(DP_OP_102J5_124_3590_n145), .SO(
        n_accumulator_sum[5]) );
  OA21X1_HVT U212 ( .A1(DP_OP_102J5_124_3590_n134), .A2(
        DP_OP_102J5_124_3590_n136), .A3(DP_OP_102J5_124_3590_n135), .Y(n176)
         );
  INVX0_HVT U213 ( .A(DP_OP_102J5_124_3590_n131), .Y(n177) );
  NAND2X0_HVT U214 ( .A1(n177), .A2(DP_OP_102J5_124_3590_n132), .Y(n178) );
  HADDX1_HVT U215 ( .A0(n176), .B0(n178), .SO(n_accumulator_sum[8]) );
  OA21X1_HVT U216 ( .A1(DP_OP_102J5_124_3590_n115), .A2(
        DP_OP_102J5_124_3590_n117), .A3(DP_OP_102J5_124_3590_n116), .Y(n179)
         );
  INVX0_HVT U217 ( .A(DP_OP_102J5_124_3590_n112), .Y(n180) );
  NAND2X0_HVT U218 ( .A1(n180), .A2(DP_OP_102J5_124_3590_n113), .Y(n181) );
  HADDX1_HVT U219 ( .A0(n179), .B0(n181), .SO(n_accumulator_sum[12]) );
  OR3X1_HVT U220 ( .A1(n182), .A2(DP_OP_102J5_124_3590_n30), .A3(
        DP_OP_102J5_124_3590_n35), .Y(n183) );
  NOR2X0_HVT U222 ( .A1(n191), .A2(n301), .Y(n186) );
  FADDX1_HVT U223 ( .A(n186), .B(n185), .CI(DP_OP_102J5_124_3590_n186), .S(
        n_accumulator_sum[22]) );
  INVX0_HVT U224 ( .A(DP_OP_102J5_124_3590_n3), .Y(n182) );
  INVX0_HVT U225 ( .A(DP_OP_102J5_124_3590_n91), .Y(DP_OP_102J5_124_3590_n89)
         );
  INVX0_HVT U226 ( .A(DP_OP_102J5_124_3590_n162), .Y(DP_OP_102J5_124_3590_n5)
         );
  INVX1_HVT U227 ( .A(DP_OP_102J5_124_3590_n2411), .Y(n191) );
  INVX2_HVT U228 ( .A(srstn), .Y(n187) );
  INVX2_HVT U229 ( .A(srstn), .Y(n188) );
  INVX2_HVT U230 ( .A(srstn), .Y(n189) );
  INVX2_HVT U231 ( .A(srstn), .Y(n190) );
  OR2X1_HVT U232 ( .A1(DP_OP_102J5_124_3590_n199), .A2(
        DP_OP_102J5_124_3590_n200), .Y(n279) );
  INVX1_HVT U233 ( .A(DP_OP_102J5_124_3590_n137), .Y(DP_OP_102J5_124_3590_n136) );
  INVX1_HVT U234 ( .A(DP_OP_102J5_124_3590_n3), .Y(DP_OP_102J5_124_3590_n106)
         );
  INVX1_HVT U235 ( .A(accumulate_reset), .Y(DP_OP_102J5_124_3590_n2411) );
  OR2X1_HVT U236 ( .A1(DP_OP_102J5_124_3590_n1198), .A2(
        DP_OP_102J5_124_3590_n1196), .Y(n284) );
  OR2X1_HVT U237 ( .A1(DP_OP_102J5_124_3590_n1320), .A2(
        DP_OP_102J5_124_3590_n1318), .Y(n285) );
  OR2X1_HVT U238 ( .A1(DP_OP_102J5_124_3590_n908), .A2(
        DP_OP_102J5_124_3590_n906), .Y(n286) );
  OR2X1_HVT U239 ( .A1(DP_OP_102J5_124_3590_n190), .A2(
        DP_OP_102J5_124_3590_n189), .Y(n290) );
  OR2X1_HVT U240 ( .A1(DP_OP_102J5_124_3590_n196), .A2(
        DP_OP_102J5_124_3590_n195), .Y(n291) );
  INVX1_HVT U241 ( .A(DP_OP_102J5_124_3590_n125), .Y(DP_OP_102J5_124_3590_n176) );
  INVX1_HVT U242 ( .A(DP_OP_102J5_124_3590_n128), .Y(DP_OP_102J5_124_3590_n127) );
  INVX1_HVT U243 ( .A(src_window[15]), .Y(DP_OP_102J5_124_3590_n1538) );
  INVX1_HVT U244 ( .A(src_window[14]), .Y(DP_OP_102J5_124_3590_n1539) );
  INVX1_HVT U245 ( .A(src_window[13]), .Y(DP_OP_102J5_124_3590_n1540) );
  INVX1_HVT U246 ( .A(src_window[12]), .Y(DP_OP_102J5_124_3590_n1541) );
  INVX1_HVT U247 ( .A(src_window[11]), .Y(DP_OP_102J5_124_3590_n1542) );
  INVX1_HVT U248 ( .A(src_window[10]), .Y(DP_OP_102J5_124_3590_n1543) );
  INVX1_HVT U249 ( .A(src_window[9]), .Y(DP_OP_102J5_124_3590_n1544) );
  INVX1_HVT U250 ( .A(src_window[8]), .Y(DP_OP_102J5_124_3590_n1545) );
  INVX1_HVT U251 ( .A(src_window[31]), .Y(DP_OP_102J5_124_3590_n1582) );
  INVX1_HVT U252 ( .A(src_window[30]), .Y(DP_OP_102J5_124_3590_n1583) );
  INVX1_HVT U253 ( .A(src_window[29]), .Y(DP_OP_102J5_124_3590_n1584) );
  INVX1_HVT U254 ( .A(src_window[28]), .Y(DP_OP_102J5_124_3590_n1585) );
  INVX1_HVT U255 ( .A(src_window[27]), .Y(DP_OP_102J5_124_3590_n1586) );
  INVX1_HVT U256 ( .A(src_window[26]), .Y(DP_OP_102J5_124_3590_n1587) );
  INVX1_HVT U257 ( .A(src_window[25]), .Y(DP_OP_102J5_124_3590_n1588) );
  INVX1_HVT U258 ( .A(src_window[24]), .Y(DP_OP_102J5_124_3590_n1589) );
  INVX1_HVT U259 ( .A(src_window[47]), .Y(DP_OP_102J5_124_3590_n1626) );
  INVX1_HVT U260 ( .A(src_window[46]), .Y(DP_OP_102J5_124_3590_n1627) );
  INVX1_HVT U261 ( .A(src_window[45]), .Y(DP_OP_102J5_124_3590_n1628) );
  INVX1_HVT U262 ( .A(src_window[44]), .Y(DP_OP_102J5_124_3590_n1629) );
  INVX1_HVT U263 ( .A(src_window[43]), .Y(DP_OP_102J5_124_3590_n1630) );
  INVX1_HVT U264 ( .A(src_window[42]), .Y(DP_OP_102J5_124_3590_n1631) );
  INVX1_HVT U265 ( .A(src_window[41]), .Y(DP_OP_102J5_124_3590_n1632) );
  INVX1_HVT U266 ( .A(src_window[40]), .Y(DP_OP_102J5_124_3590_n1633) );
  INVX1_HVT U267 ( .A(src_window[63]), .Y(DP_OP_102J5_124_3590_n1670) );
  INVX1_HVT U268 ( .A(src_window[62]), .Y(DP_OP_102J5_124_3590_n1671) );
  INVX1_HVT U269 ( .A(src_window[61]), .Y(DP_OP_102J5_124_3590_n1672) );
  INVX1_HVT U270 ( .A(src_window[60]), .Y(DP_OP_102J5_124_3590_n1673) );
  INVX1_HVT U271 ( .A(src_window[59]), .Y(DP_OP_102J5_124_3590_n1674) );
  INVX1_HVT U272 ( .A(src_window[58]), .Y(DP_OP_102J5_124_3590_n1675) );
  INVX1_HVT U273 ( .A(src_window[57]), .Y(DP_OP_102J5_124_3590_n1676) );
  INVX1_HVT U274 ( .A(src_window[56]), .Y(DP_OP_102J5_124_3590_n1677) );
  INVX1_HVT U275 ( .A(DP_OP_102J5_124_3590_n75), .Y(DP_OP_102J5_124_3590_n77)
         );
  INVX1_HVT U276 ( .A(DP_OP_102J5_124_3590_n97), .Y(DP_OP_102J5_124_3590_n99)
         );
  INVX1_HVT U277 ( .A(src_window[79]), .Y(DP_OP_102J5_124_3590_n1714) );
  INVX1_HVT U278 ( .A(src_window[78]), .Y(DP_OP_102J5_124_3590_n1715) );
  INVX1_HVT U279 ( .A(src_window[77]), .Y(DP_OP_102J5_124_3590_n1716) );
  INVX1_HVT U280 ( .A(src_window[76]), .Y(DP_OP_102J5_124_3590_n1717) );
  INVX1_HVT U281 ( .A(src_window[75]), .Y(DP_OP_102J5_124_3590_n1718) );
  INVX1_HVT U282 ( .A(src_window[74]), .Y(DP_OP_102J5_124_3590_n1719) );
  INVX1_HVT U283 ( .A(src_window[73]), .Y(DP_OP_102J5_124_3590_n1720) );
  INVX1_HVT U284 ( .A(src_window[72]), .Y(DP_OP_102J5_124_3590_n1721) );
  INVX1_HVT U285 ( .A(src_window[95]), .Y(DP_OP_102J5_124_3590_n1758) );
  INVX1_HVT U286 ( .A(src_window[94]), .Y(DP_OP_102J5_124_3590_n1759) );
  INVX1_HVT U287 ( .A(src_window[93]), .Y(DP_OP_102J5_124_3590_n1760) );
  INVX1_HVT U288 ( .A(src_window[92]), .Y(DP_OP_102J5_124_3590_n1761) );
  INVX1_HVT U289 ( .A(src_window[91]), .Y(DP_OP_102J5_124_3590_n1762) );
  INVX1_HVT U290 ( .A(src_window[90]), .Y(DP_OP_102J5_124_3590_n1763) );
  INVX1_HVT U291 ( .A(src_window[89]), .Y(DP_OP_102J5_124_3590_n1764) );
  INVX1_HVT U292 ( .A(src_window[88]), .Y(DP_OP_102J5_124_3590_n1765) );
  INVX1_HVT U293 ( .A(src_window[111]), .Y(DP_OP_102J5_124_3590_n1802) );
  INVX1_HVT U294 ( .A(src_window[110]), .Y(DP_OP_102J5_124_3590_n1803) );
  INVX1_HVT U295 ( .A(src_window[109]), .Y(DP_OP_102J5_124_3590_n1804) );
  INVX1_HVT U296 ( .A(src_window[108]), .Y(DP_OP_102J5_124_3590_n1805) );
  INVX1_HVT U297 ( .A(src_window[107]), .Y(DP_OP_102J5_124_3590_n1806) );
  INVX1_HVT U298 ( .A(src_window[106]), .Y(DP_OP_102J5_124_3590_n1807) );
  INVX1_HVT U299 ( .A(src_window[105]), .Y(DP_OP_102J5_124_3590_n1808) );
  INVX1_HVT U300 ( .A(src_window[104]), .Y(DP_OP_102J5_124_3590_n1809) );
  INVX1_HVT U301 ( .A(src_window[127]), .Y(DP_OP_102J5_124_3590_n1845) );
  INVX1_HVT U302 ( .A(src_window[126]), .Y(DP_OP_102J5_124_3590_n1846) );
  INVX1_HVT U303 ( .A(src_window[125]), .Y(DP_OP_102J5_124_3590_n1847) );
  INVX1_HVT U304 ( .A(src_window[124]), .Y(DP_OP_102J5_124_3590_n1848) );
  INVX1_HVT U305 ( .A(src_window[123]), .Y(DP_OP_102J5_124_3590_n1849) );
  INVX1_HVT U306 ( .A(src_window[122]), .Y(DP_OP_102J5_124_3590_n1850) );
  INVX1_HVT U307 ( .A(src_window[121]), .Y(DP_OP_102J5_124_3590_n1851) );
  INVX1_HVT U308 ( .A(src_window[120]), .Y(DP_OP_102J5_124_3590_n1852) );
  INVX1_HVT U309 ( .A(DP_OP_102J5_124_3590_n186), .Y(DP_OP_102J5_124_3590_n187) );
  INVX1_HVT U310 ( .A(src_window[143]), .Y(DP_OP_102J5_124_3590_n1889) );
  INVX1_HVT U311 ( .A(DP_OP_102J5_124_3590_n188), .Y(DP_OP_102J5_124_3590_n189) );
  INVX1_HVT U312 ( .A(src_window[142]), .Y(DP_OP_102J5_124_3590_n1890) );
  INVX1_HVT U313 ( .A(src_window[141]), .Y(DP_OP_102J5_124_3590_n1891) );
  INVX1_HVT U314 ( .A(src_window[140]), .Y(DP_OP_102J5_124_3590_n1892) );
  INVX1_HVT U315 ( .A(src_window[139]), .Y(DP_OP_102J5_124_3590_n1893) );
  INVX1_HVT U316 ( .A(src_window[138]), .Y(DP_OP_102J5_124_3590_n1894) );
  INVX1_HVT U317 ( .A(src_window[137]), .Y(DP_OP_102J5_124_3590_n1895) );
  INVX1_HVT U318 ( .A(src_window[136]), .Y(DP_OP_102J5_124_3590_n1896) );
  INVX1_HVT U319 ( .A(DP_OP_102J5_124_3590_n190), .Y(DP_OP_102J5_124_3590_n191) );
  INVX1_HVT U320 ( .A(DP_OP_102J5_124_3590_n192), .Y(DP_OP_102J5_124_3590_n193) );
  INVX1_HVT U321 ( .A(src_window[159]), .Y(DP_OP_102J5_124_3590_n1933) );
  INVX1_HVT U322 ( .A(src_window[158]), .Y(DP_OP_102J5_124_3590_n1934) );
  INVX1_HVT U323 ( .A(src_window[157]), .Y(DP_OP_102J5_124_3590_n1935) );
  INVX1_HVT U324 ( .A(src_window[156]), .Y(DP_OP_102J5_124_3590_n1936) );
  INVX1_HVT U325 ( .A(src_window[155]), .Y(DP_OP_102J5_124_3590_n1937) );
  INVX1_HVT U326 ( .A(src_window[154]), .Y(DP_OP_102J5_124_3590_n1938) );
  INVX1_HVT U327 ( .A(src_window[153]), .Y(DP_OP_102J5_124_3590_n1939) );
  INVX1_HVT U328 ( .A(src_window[152]), .Y(DP_OP_102J5_124_3590_n1940) );
  INVX1_HVT U329 ( .A(DP_OP_102J5_124_3590_n194), .Y(DP_OP_102J5_124_3590_n195) );
  INVX1_HVT U330 ( .A(DP_OP_102J5_124_3590_n196), .Y(DP_OP_102J5_124_3590_n197) );
  INVX1_HVT U331 ( .A(src_window[151]), .Y(DP_OP_102J5_124_3590_n1977) );
  INVX1_HVT U332 ( .A(src_window[150]), .Y(DP_OP_102J5_124_3590_n1978) );
  INVX1_HVT U333 ( .A(src_window[149]), .Y(DP_OP_102J5_124_3590_n1979) );
  INVX1_HVT U334 ( .A(src_window[148]), .Y(DP_OP_102J5_124_3590_n1980) );
  INVX1_HVT U335 ( .A(src_window[147]), .Y(DP_OP_102J5_124_3590_n1981) );
  INVX1_HVT U336 ( .A(src_window[146]), .Y(DP_OP_102J5_124_3590_n1982) );
  INVX1_HVT U337 ( .A(src_window[145]), .Y(DP_OP_102J5_124_3590_n1983) );
  INVX1_HVT U338 ( .A(src_window[144]), .Y(DP_OP_102J5_124_3590_n1984) );
  INVX1_HVT U339 ( .A(src_window[135]), .Y(DP_OP_102J5_124_3590_n2021) );
  INVX1_HVT U340 ( .A(src_window[134]), .Y(DP_OP_102J5_124_3590_n2022) );
  INVX1_HVT U341 ( .A(src_window[133]), .Y(DP_OP_102J5_124_3590_n2023) );
  INVX1_HVT U342 ( .A(src_window[132]), .Y(DP_OP_102J5_124_3590_n2024) );
  INVX1_HVT U343 ( .A(src_window[131]), .Y(DP_OP_102J5_124_3590_n2025) );
  INVX1_HVT U344 ( .A(src_window[130]), .Y(DP_OP_102J5_124_3590_n2026) );
  INVX1_HVT U345 ( .A(src_window[129]), .Y(DP_OP_102J5_124_3590_n2027) );
  INVX1_HVT U346 ( .A(src_window[128]), .Y(DP_OP_102J5_124_3590_n2028) );
  INVX1_HVT U347 ( .A(DP_OP_102J5_124_3590_n204), .Y(DP_OP_102J5_124_3590_n205) );
  INVX1_HVT U348 ( .A(src_window[119]), .Y(DP_OP_102J5_124_3590_n2065) );
  INVX1_HVT U349 ( .A(src_window[118]), .Y(DP_OP_102J5_124_3590_n2066) );
  INVX1_HVT U350 ( .A(src_window[117]), .Y(DP_OP_102J5_124_3590_n2067) );
  INVX1_HVT U351 ( .A(src_window[116]), .Y(DP_OP_102J5_124_3590_n2068) );
  INVX1_HVT U352 ( .A(src_window[115]), .Y(DP_OP_102J5_124_3590_n2069) );
  INVX1_HVT U353 ( .A(src_window[114]), .Y(DP_OP_102J5_124_3590_n2070) );
  INVX1_HVT U354 ( .A(src_window[113]), .Y(DP_OP_102J5_124_3590_n2071) );
  INVX1_HVT U355 ( .A(src_window[112]), .Y(DP_OP_102J5_124_3590_n2072) );
  INVX1_HVT U356 ( .A(src_window[103]), .Y(DP_OP_102J5_124_3590_n2109) );
  INVX1_HVT U357 ( .A(src_window[102]), .Y(DP_OP_102J5_124_3590_n2110) );
  INVX1_HVT U358 ( .A(src_window[101]), .Y(DP_OP_102J5_124_3590_n2111) );
  INVX1_HVT U359 ( .A(src_window[100]), .Y(DP_OP_102J5_124_3590_n2112) );
  INVX1_HVT U360 ( .A(src_window[99]), .Y(DP_OP_102J5_124_3590_n2113) );
  INVX1_HVT U361 ( .A(src_window[98]), .Y(DP_OP_102J5_124_3590_n2114) );
  INVX1_HVT U362 ( .A(src_window[97]), .Y(DP_OP_102J5_124_3590_n2115) );
  INVX1_HVT U363 ( .A(src_window[96]), .Y(DP_OP_102J5_124_3590_n2116) );
  INVX1_HVT U364 ( .A(DP_OP_102J5_124_3590_n214), .Y(DP_OP_102J5_124_3590_n215) );
  INVX1_HVT U365 ( .A(src_window[87]), .Y(DP_OP_102J5_124_3590_n2153) );
  INVX1_HVT U366 ( .A(src_window[86]), .Y(DP_OP_102J5_124_3590_n2154) );
  INVX1_HVT U367 ( .A(src_window[85]), .Y(DP_OP_102J5_124_3590_n2155) );
  INVX1_HVT U368 ( .A(src_window[84]), .Y(DP_OP_102J5_124_3590_n2156) );
  INVX1_HVT U369 ( .A(src_window[83]), .Y(DP_OP_102J5_124_3590_n2157) );
  INVX1_HVT U370 ( .A(src_window[82]), .Y(DP_OP_102J5_124_3590_n2158) );
  INVX1_HVT U371 ( .A(src_window[81]), .Y(DP_OP_102J5_124_3590_n2159) );
  INVX1_HVT U372 ( .A(src_window[80]), .Y(DP_OP_102J5_124_3590_n2160) );
  INVX1_HVT U373 ( .A(src_window[71]), .Y(DP_OP_102J5_124_3590_n2197) );
  INVX1_HVT U374 ( .A(src_window[70]), .Y(DP_OP_102J5_124_3590_n2198) );
  INVX1_HVT U375 ( .A(src_window[69]), .Y(DP_OP_102J5_124_3590_n2199) );
  INVX1_HVT U376 ( .A(src_window[68]), .Y(DP_OP_102J5_124_3590_n2200) );
  INVX1_HVT U377 ( .A(src_window[67]), .Y(DP_OP_102J5_124_3590_n2201) );
  INVX1_HVT U378 ( .A(src_window[66]), .Y(DP_OP_102J5_124_3590_n2202) );
  INVX1_HVT U379 ( .A(src_window[65]), .Y(DP_OP_102J5_124_3590_n2203) );
  INVX1_HVT U380 ( .A(src_window[64]), .Y(DP_OP_102J5_124_3590_n2204) );
  INVX1_HVT U381 ( .A(src_window[55]), .Y(DP_OP_102J5_124_3590_n2241) );
  INVX1_HVT U382 ( .A(src_window[54]), .Y(DP_OP_102J5_124_3590_n2242) );
  INVX1_HVT U383 ( .A(src_window[53]), .Y(DP_OP_102J5_124_3590_n2243) );
  INVX1_HVT U384 ( .A(src_window[52]), .Y(DP_OP_102J5_124_3590_n2244) );
  INVX1_HVT U385 ( .A(src_window[51]), .Y(DP_OP_102J5_124_3590_n2245) );
  INVX1_HVT U386 ( .A(src_window[50]), .Y(DP_OP_102J5_124_3590_n2246) );
  INVX1_HVT U387 ( .A(src_window[49]), .Y(DP_OP_102J5_124_3590_n2247) );
  INVX1_HVT U388 ( .A(src_window[48]), .Y(DP_OP_102J5_124_3590_n2248) );
  INVX1_HVT U389 ( .A(src_window[39]), .Y(DP_OP_102J5_124_3590_n2285) );
  INVX1_HVT U390 ( .A(src_window[38]), .Y(DP_OP_102J5_124_3590_n2286) );
  INVX1_HVT U391 ( .A(src_window[37]), .Y(DP_OP_102J5_124_3590_n2287) );
  INVX1_HVT U392 ( .A(src_window[36]), .Y(DP_OP_102J5_124_3590_n2288) );
  INVX1_HVT U393 ( .A(src_window[35]), .Y(DP_OP_102J5_124_3590_n2289) );
  INVX1_HVT U394 ( .A(src_window[34]), .Y(DP_OP_102J5_124_3590_n2290) );
  INVX1_HVT U395 ( .A(src_window[33]), .Y(DP_OP_102J5_124_3590_n2291) );
  INVX1_HVT U396 ( .A(src_window[32]), .Y(DP_OP_102J5_124_3590_n2292) );
  INVX1_HVT U397 ( .A(src_window[23]), .Y(DP_OP_102J5_124_3590_n2329) );
  INVX1_HVT U398 ( .A(src_window[22]), .Y(DP_OP_102J5_124_3590_n2330) );
  INVX1_HVT U399 ( .A(src_window[21]), .Y(DP_OP_102J5_124_3590_n2331) );
  INVX1_HVT U400 ( .A(src_window[20]), .Y(DP_OP_102J5_124_3590_n2332) );
  INVX1_HVT U401 ( .A(src_window[19]), .Y(DP_OP_102J5_124_3590_n2333) );
  INVX1_HVT U402 ( .A(src_window[18]), .Y(DP_OP_102J5_124_3590_n2334) );
  INVX1_HVT U403 ( .A(src_window[17]), .Y(DP_OP_102J5_124_3590_n2335) );
  INVX1_HVT U404 ( .A(src_window[16]), .Y(DP_OP_102J5_124_3590_n2336) );
  INVX1_HVT U405 ( .A(src_window[7]), .Y(DP_OP_102J5_124_3590_n2372) );
  INVX1_HVT U406 ( .A(src_window[6]), .Y(DP_OP_102J5_124_3590_n2373) );
  INVX1_HVT U407 ( .A(src_window[5]), .Y(DP_OP_102J5_124_3590_n2374) );
  INVX1_HVT U408 ( .A(src_window[4]), .Y(DP_OP_102J5_124_3590_n2375) );
  INVX1_HVT U409 ( .A(src_window[3]), .Y(DP_OP_102J5_124_3590_n2376) );
  INVX1_HVT U410 ( .A(src_window[2]), .Y(DP_OP_102J5_124_3590_n2377) );
  INVX1_HVT U411 ( .A(src_window[1]), .Y(DP_OP_102J5_124_3590_n2378) );
  INVX1_HVT U412 ( .A(src_window[0]), .Y(DP_OP_102J5_124_3590_n2379) );
  INVX1_HVT U413 ( .A(DP_OP_102J5_124_3590_n270), .Y(DP_OP_102J5_124_3590_n271) );
  INVX1_HVT U414 ( .A(DP_OP_102J5_124_3590_n453), .Y(DP_OP_102J5_124_3590_n454) );
  INVX1_HVT U415 ( .A(DP_OP_102J5_124_3590_n749), .Y(DP_OP_102J5_124_3590_n750) );
  INVX1_HVT U416 ( .A(DP_OP_102J5_124_3590_n95), .Y(DP_OP_102J5_124_3590_n93)
         );
  INVX1_HVT U417 ( .A(DP_OP_102J5_124_3590_n96), .Y(DP_OP_102J5_124_3590_n94)
         );
endmodule


module fc_quantize ( clk, srstn, fc_state, quantized_data, 
        unquautized_data_22_, unquautized_data_21_, unquautized_data_20_, 
        unquautized_data_19_, unquautized_data_18_, unquautized_data_17_, 
        unquautized_data_16_, unquautized_data_15_, unquautized_data_14_, 
        unquautized_data_13_, unquautized_data_12_, unquautized_data_11_, 
        unquautized_data_10_, unquautized_data_9_, unquautized_data_8_, 
        unquautized_data_7_, unquautized_data_6_, unquautized_data_5_, 
        unquautized_data_4_ );
  output [7:0] quantized_data;
  input clk, srstn, fc_state, unquautized_data_22_, unquautized_data_21_,
         unquautized_data_20_, unquautized_data_19_, unquautized_data_18_,
         unquautized_data_17_, unquautized_data_16_, unquautized_data_15_,
         unquautized_data_14_, unquautized_data_13_, unquautized_data_12_,
         unquautized_data_11_, unquautized_data_10_, unquautized_data_9_,
         unquautized_data_8_, unquautized_data_7_, unquautized_data_6_,
         unquautized_data_5_, unquautized_data_4_;
  wire   n13, n1, n2, n4, n5, n6, n7, n10, n11, n12, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82;
  wire   [7:0] n_quantized_data;

  DFFSSRX1_HVT quantized_data_reg_7_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[7]), .CLK(clk), .Q(quantized_data[7]) );
  DFFSSRX1_HVT quantized_data_reg_6_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[6]), .CLK(clk), .Q(quantized_data[6]) );
  DFFSSRX1_HVT quantized_data_reg_5_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[5]), .CLK(clk), .Q(quantized_data[5]) );
  DFFSSRX1_HVT quantized_data_reg_4_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[4]), .CLK(clk), .Q(quantized_data[4]) );
  DFFSSRX1_HVT quantized_data_reg_3_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[3]), .CLK(clk), .Q(quantized_data[3]) );
  DFFSSRX1_HVT quantized_data_reg_2_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[2]), .CLK(clk), .Q(quantized_data[2]) );
  DFFSSRX1_HVT quantized_data_reg_1_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[1]), .CLK(clk), .Q(quantized_data[1]) );
  DFFSSRX1_HVT quantized_data_reg_0_ ( .D(1'b0), .SETB(n13), .RSTB(
        n_quantized_data[0]), .CLK(clk), .Q(quantized_data[0]) );
  AO221X1_HVT U3 ( .A1(1'b1), .A2(n67), .A3(n59), .A4(n6), .A5(n7), .Y(n10) );
  AO221X1_HVT U4 ( .A1(1'b1), .A2(n58), .A3(n49), .A4(n1), .A5(n2), .Y(n4) );
  NAND3X0_HVT U5 ( .A1(unquautized_data_6_), .A2(unquautized_data_5_), .A3(
        unquautized_data_4_), .Y(n1) );
  INVX0_HVT U6 ( .A(n66), .Y(n2) );
  AO21X1_HVT U8 ( .A1(n55), .A2(n50), .A3(n53), .Y(n5) );
  NAND3X0_HVT U9 ( .A1(n81), .A2(n4), .A3(n5), .Y(n_quantized_data[2]) );
  NAND2X0_HVT U10 ( .A1(unquautized_data_8_), .A2(n58), .Y(n6) );
  INVX0_HVT U11 ( .A(n66), .Y(n7) );
  AO21X1_HVT U13 ( .A1(n65), .A2(n60), .A3(n63), .Y(n11) );
  NAND3X0_HVT U14 ( .A1(n81), .A2(n10), .A3(n11), .Y(n_quantized_data[4]) );
  INVX1_HVT U15 ( .A(n33), .Y(n78) );
  INVX0_HVT U16 ( .A(n21), .Y(n73) );
  INVX0_HVT U17 ( .A(unquautized_data_9_), .Y(n59) );
  INVX0_HVT U18 ( .A(unquautized_data_15_), .Y(n25) );
  INVX0_HVT U19 ( .A(unquautized_data_19_), .Y(n27) );
  INVX0_HVT U20 ( .A(unquautized_data_20_), .Y(n23) );
  INVX0_HVT U21 ( .A(unquautized_data_21_), .Y(n24) );
  INVX0_HVT U22 ( .A(unquautized_data_13_), .Y(n22) );
  INVX0_HVT U23 ( .A(unquautized_data_7_), .Y(n49) );
  INVX0_HVT U24 ( .A(unquautized_data_6_), .Y(n45) );
  INVX0_HVT U25 ( .A(unquautized_data_5_), .Y(n39) );
  INVX1_HVT U26 ( .A(srstn), .Y(n13) );
  INVX1_HVT U27 ( .A(n70), .Y(n66) );
  INVX1_HVT U28 ( .A(n41), .Y(n81) );
  OR2X1_HVT U29 ( .A1(n72), .A2(n71), .Y(n21) );
  INVX1_HVT U30 ( .A(unquautized_data_22_), .Y(n36) );
  INVX1_HVT U31 ( .A(unquautized_data_10_), .Y(n65) );
  INVX1_HVT U32 ( .A(unquautized_data_8_), .Y(n55) );
  INVX1_HVT U33 ( .A(n75), .Y(n61) );
  INVX1_HVT U34 ( .A(fc_state), .Y(n20) );
  INVX1_HVT U35 ( .A(unquautized_data_17_), .Y(n34) );
  INVX1_HVT U36 ( .A(n60), .Y(n74) );
  INVX1_HVT U37 ( .A(n50), .Y(n51) );
  INVX1_HVT U38 ( .A(unquautized_data_12_), .Y(n77) );
  INVX1_HVT U39 ( .A(unquautized_data_11_), .Y(n71) );
  NAND2X0_HVT U40 ( .A1(n77), .A2(n76), .Y(n12) );
  NAND3X0_HVT U41 ( .A1(n61), .A2(n33), .A3(n12), .Y(n79) );
  NAND2X0_HVT U42 ( .A1(n72), .A2(n71), .Y(n14) );
  NAND3X0_HVT U43 ( .A1(n66), .A2(n21), .A3(n14), .Y(n80) );
  AND4X1_HVT U44 ( .A1(unquautized_data_20_), .A2(unquautized_data_19_), .A3(
        unquautized_data_18_), .A4(unquautized_data_17_), .Y(n15) );
  AND4X1_HVT U45 ( .A1(unquautized_data_16_), .A2(unquautized_data_14_), .A3(
        unquautized_data_21_), .A4(n15), .Y(n16) );
  NAND3X0_HVT U46 ( .A1(unquautized_data_13_), .A2(unquautized_data_15_), .A3(
        n16), .Y(n19) );
  AND4X1_HVT U47 ( .A1(unquautized_data_6_), .A2(unquautized_data_5_), .A3(
        unquautized_data_4_), .A4(unquautized_data_7_), .Y(n58) );
  AND3X1_HVT U48 ( .A1(n58), .A2(unquautized_data_8_), .A3(unquautized_data_9_), .Y(n67) );
  NAND2X0_HVT U49 ( .A1(n67), .A2(unquautized_data_10_), .Y(n72) );
  OR3X1_HVT U50 ( .A1(n19), .A2(n21), .A3(n77), .Y(n17) );
  HADDX1_HVT U51 ( .A0(n36), .B0(n17), .SO(n82) );
  HADDX1_HVT U52 ( .A0(unquautized_data_12_), .B0(n21), .SO(n18) );
  AO221X1_HVT U53 ( .A1(n82), .A2(n19), .A3(n82), .A4(n18), .A5(n20), .Y(n70)
         );
  NAND2X0_HVT U54 ( .A1(n36), .A2(n20), .Y(n75) );
  OAI22X1_HVT U55 ( .A1(unquautized_data_4_), .A2(n70), .A3(
        unquautized_data_6_), .A4(n75), .Y(n40) );
  AO22X1_HVT U56 ( .A1(unquautized_data_6_), .A2(n61), .A3(unquautized_data_4_), .A4(n66), .Y(n38) );
  OA221X1_HVT U57 ( .A1(unquautized_data_12_), .A2(n73), .A3(n77), .A4(n21), 
        .A5(n36), .Y(n37) );
  NAND3X0_HVT U58 ( .A1(unquautized_data_6_), .A2(unquautized_data_5_), .A3(
        unquautized_data_7_), .Y(n50) );
  NAND3X0_HVT U59 ( .A1(unquautized_data_8_), .A2(unquautized_data_9_), .A3(
        n51), .Y(n60) );
  NAND4X0_HVT U60 ( .A1(unquautized_data_10_), .A2(unquautized_data_12_), .A3(
        unquautized_data_11_), .A4(n74), .Y(n33) );
  OA222X1_HVT U61 ( .A1(n22), .A2(n78), .A3(n22), .A4(unquautized_data_15_), 
        .A5(n33), .A6(unquautized_data_13_), .Y(n31) );
  OA222X1_HVT U62 ( .A1(unquautized_data_20_), .A2(n24), .A3(n23), .A4(n78), 
        .A5(unquautized_data_21_), .A6(n33), .Y(n30) );
  OA22X1_HVT U63 ( .A1(unquautized_data_16_), .A2(n34), .A3(
        unquautized_data_14_), .A4(n25), .Y(n26) );
  OA221X1_HVT U64 ( .A1(unquautized_data_19_), .A2(n33), .A3(n27), .A4(
        unquautized_data_18_), .A5(n26), .Y(n29) );
  OAI21X1_HVT U65 ( .A1(unquautized_data_18_), .A2(unquautized_data_16_), .A3(
        n33), .Y(n28) );
  NAND4X0_HVT U66 ( .A1(n31), .A2(n30), .A3(n29), .A4(n28), .Y(n32) );
  AO221X1_HVT U67 ( .A1(n78), .A2(n34), .A3(n33), .A4(unquautized_data_14_), 
        .A5(n32), .Y(n35) );
  AO22X1_HVT U68 ( .A1(n37), .A2(fc_state), .A3(n36), .A4(n35), .Y(n41) );
  AO221X1_HVT U69 ( .A1(unquautized_data_5_), .A2(n40), .A3(n39), .A4(n38), 
        .A5(n41), .Y(n_quantized_data[0]) );
  NAND3X0_HVT U70 ( .A1(unquautized_data_5_), .A2(n61), .A3(n49), .Y(n44) );
  NAND2X0_HVT U71 ( .A1(unquautized_data_5_), .A2(unquautized_data_4_), .Y(n42) );
  HADDX1_HVT U72 ( .A0(unquautized_data_6_), .B0(n42), .SO(n43) );
  OA22X1_HVT U73 ( .A1(n45), .A2(n44), .A3(n70), .A4(n43), .Y(n48) );
  NAND2X0_HVT U74 ( .A1(unquautized_data_6_), .A2(unquautized_data_5_), .Y(n46) );
  NAND3X0_HVT U75 ( .A1(unquautized_data_7_), .A2(n61), .A3(n46), .Y(n47) );
  NAND3X0_HVT U76 ( .A1(n81), .A2(n48), .A3(n47), .Y(n_quantized_data[1]) );
  AO21X1_HVT U77 ( .A1(unquautized_data_8_), .A2(n51), .A3(n75), .Y(n53) );
  NAND2X0_HVT U78 ( .A1(n51), .A2(n61), .Y(n52) );
  OA22X1_HVT U79 ( .A1(unquautized_data_9_), .A2(n52), .A3(n58), .A4(n70), .Y(
        n54) );
  OA22X1_HVT U80 ( .A1(n54), .A2(n55), .A3(n59), .A4(n53), .Y(n57) );
  NAND3X0_HVT U81 ( .A1(n58), .A2(n66), .A3(n55), .Y(n56) );
  NAND3X0_HVT U82 ( .A1(n81), .A2(n57), .A3(n56), .Y(n_quantized_data[3]) );
  AO21X1_HVT U83 ( .A1(unquautized_data_10_), .A2(n74), .A3(n75), .Y(n63) );
  NAND2X0_HVT U84 ( .A1(n74), .A2(n61), .Y(n62) );
  OA22X1_HVT U85 ( .A1(unquautized_data_11_), .A2(n62), .A3(n67), .A4(n70), 
        .Y(n64) );
  OA22X1_HVT U86 ( .A1(n64), .A2(n65), .A3(n71), .A4(n63), .Y(n69) );
  NAND3X0_HVT U87 ( .A1(n67), .A2(n66), .A3(n65), .Y(n68) );
  NAND3X0_HVT U88 ( .A1(n81), .A2(n69), .A3(n68), .Y(n_quantized_data[5]) );
  NAND3X0_HVT U89 ( .A1(unquautized_data_10_), .A2(unquautized_data_11_), .A3(
        n74), .Y(n76) );
  NAND3X0_HVT U90 ( .A1(n81), .A2(n80), .A3(n79), .Y(n_quantized_data[6]) );
  AND2X1_HVT U91 ( .A1(n82), .A2(fc_state), .Y(n_quantized_data[7]) );
endmodule


module fc_top ( clk, srstn, conv_done, mem_sel, sram_rdata_c0, sram_rdata_c1, 
        sram_rdata_c2, sram_rdata_c3, sram_rdata_c4, sram_raddr_c0, 
        sram_raddr_c1, sram_raddr_c2, sram_raddr_c3, sram_raddr_c4, 
        sram_rdata_d0, sram_rdata_d1, sram_rdata_d2, sram_rdata_d3, 
        sram_rdata_d4, sram_raddr_d0, sram_raddr_d1, sram_raddr_d2, 
        sram_raddr_d3, sram_raddr_d4, sram_rdata_e0, sram_rdata_e1, 
        sram_rdata_e2, sram_rdata_e3, sram_rdata_e4, sram_raddr_e0, 
        sram_raddr_e1, sram_raddr_e2, sram_raddr_e3, sram_raddr_e4, 
        sram_write_enable_e0, sram_write_enable_e1, sram_write_enable_e2, 
        sram_write_enable_e3, sram_write_enable_e4, sram_bytemask_e, 
        sram_waddr_e, sram_wdata_e, sram_write_enable_f, sram_bytemask_f, 
        sram_waddr_f, sram_wdata_f, sram_rdata_weight, sram_raddr_weight, 
        fc1_done, fc2_done );
  input [31:0] sram_rdata_c0;
  input [31:0] sram_rdata_c1;
  input [31:0] sram_rdata_c2;
  input [31:0] sram_rdata_c3;
  input [31:0] sram_rdata_c4;
  output [5:0] sram_raddr_c0;
  output [5:0] sram_raddr_c1;
  output [5:0] sram_raddr_c2;
  output [5:0] sram_raddr_c3;
  output [5:0] sram_raddr_c4;
  input [31:0] sram_rdata_d0;
  input [31:0] sram_rdata_d1;
  input [31:0] sram_rdata_d2;
  input [31:0] sram_rdata_d3;
  input [31:0] sram_rdata_d4;
  output [5:0] sram_raddr_d0;
  output [5:0] sram_raddr_d1;
  output [5:0] sram_raddr_d2;
  output [5:0] sram_raddr_d3;
  output [5:0] sram_raddr_d4;
  input [31:0] sram_rdata_e0;
  input [31:0] sram_rdata_e1;
  input [31:0] sram_rdata_e2;
  input [31:0] sram_rdata_e3;
  input [31:0] sram_rdata_e4;
  output [4:0] sram_raddr_e0;
  output [4:0] sram_raddr_e1;
  output [4:0] sram_raddr_e2;
  output [4:0] sram_raddr_e3;
  output [4:0] sram_raddr_e4;
  output [3:0] sram_bytemask_e;
  output [4:0] sram_waddr_e;
  output [7:0] sram_wdata_e;
  output [3:0] sram_bytemask_f;
  output [1:0] sram_waddr_f;
  output [7:0] sram_wdata_f;
  input [79:0] sram_rdata_weight;
  output [14:0] sram_raddr_weight;
  input clk, srstn, conv_done, mem_sel;
  output sram_write_enable_e0, sram_write_enable_e1, sram_write_enable_e2,
         sram_write_enable_e3, sram_write_enable_e4, sram_write_enable_f,
         fc1_done, fc2_done;
  wire   accumulate_reset, fc_state, data_out_22_, data_out_21_, data_out_20_,
         data_out_19_, data_out_18_, data_out_17_, data_out_16_, data_out_15_,
         data_out_14_, data_out_13_, data_out_12_, data_out_11_, data_out_10_,
         data_out_9_, data_out_8_, data_out_7_, data_out_6_, data_out_5_,
         data_out_4_, data_out_3_, data_out_2_, data_out_1_, data_out_0_,
         SYNOPSYS_UNCONNECTED_1;
  wire   [1:0] sram_sel;
  wire   [159:0] src_window;

  fc_controller fc_controller ( .clk(clk), .srstn(srstn), .conv_done(conv_done), .mem_sel(mem_sel), .accumulate_reset(accumulate_reset), .fc_state(fc_state), 
        .sram_sel(sram_sel), .sram_raddr_c0(sram_raddr_c0), .sram_raddr_c1(
        sram_raddr_c1), .sram_raddr_c2(sram_raddr_c2), .sram_raddr_c3(
        sram_raddr_c3), .sram_raddr_c4(sram_raddr_c4), .sram_raddr_d0(
        sram_raddr_d0), .sram_raddr_d1(sram_raddr_d1), .sram_raddr_d2(
        sram_raddr_d2), .sram_raddr_d3(sram_raddr_d3), .sram_raddr_d4(
        sram_raddr_d4), .sram_raddr_e0(sram_raddr_e0), .sram_raddr_e1(
        sram_raddr_e1), .sram_raddr_e2(sram_raddr_e2), .sram_raddr_e3(
        sram_raddr_e3), .sram_raddr_e4(sram_raddr_e4), .sram_write_enable_e0(
        sram_write_enable_e0), .sram_write_enable_e1(sram_write_enable_e1), 
        .sram_write_enable_e2(sram_write_enable_e2), .sram_write_enable_e3(
        sram_write_enable_e3), .sram_write_enable_e4(sram_write_enable_e4), 
        .sram_write_enable_f(sram_write_enable_f), .sram_waddr({
        SYNOPSYS_UNCONNECTED_1, sram_waddr_e}), .sram_bytemask(sram_bytemask_e), .sram_raddr_weight(sram_raddr_weight), .fc1_done(fc1_done), .fc2_done(
        fc2_done) );
  fc_data_reg fc_data_reg ( .clk(clk), .srstn(srstn), .sram_rdata_c0(
        sram_rdata_c0), .sram_rdata_c1(sram_rdata_c1), .sram_rdata_c2(
        sram_rdata_c2), .sram_rdata_c3(sram_rdata_c3), .sram_rdata_c4(
        sram_rdata_c4), .sram_rdata_d0(sram_rdata_d0), .sram_rdata_d1(
        sram_rdata_d1), .sram_rdata_d2(sram_rdata_d2), .sram_rdata_d3(
        sram_rdata_d3), .sram_rdata_d4(sram_rdata_d4), .sram_rdata_e0(
        sram_rdata_e0), .sram_rdata_e1(sram_rdata_e1), .sram_rdata_e2(
        sram_rdata_e2), .sram_rdata_e3(sram_rdata_e3), .sram_rdata_e4(
        sram_rdata_e4), .sram_sel(sram_sel), .src_window(src_window) );
  fc_multiplier_accumulator fc_multiplier_accumulator ( .clk(clk), .srstn(
        srstn), .src_window(src_window), .sram_rdata_weight(sram_rdata_weight), 
        .accumulate_reset(accumulate_reset), .data_out({data_out_22_, 
        data_out_21_, data_out_20_, data_out_19_, data_out_18_, data_out_17_, 
        data_out_16_, data_out_15_, data_out_14_, data_out_13_, data_out_12_, 
        data_out_11_, data_out_10_, data_out_9_, data_out_8_, data_out_7_, 
        data_out_6_, data_out_5_, data_out_4_, data_out_3_, data_out_2_, 
        data_out_1_, data_out_0_}) );
  fc_quantize fc_quantize ( .clk(clk), .srstn(srstn), .fc_state(fc_state), 
        .quantized_data(sram_wdata_e), .unquautized_data_22_(data_out_22_), 
        .unquautized_data_21_(data_out_21_), .unquautized_data_20_(
        data_out_20_), .unquautized_data_19_(data_out_19_), 
        .unquautized_data_18_(data_out_18_), .unquautized_data_17_(
        data_out_17_), .unquautized_data_16_(data_out_16_), 
        .unquautized_data_15_(data_out_15_), .unquautized_data_14_(
        data_out_14_), .unquautized_data_13_(data_out_13_), 
        .unquautized_data_12_(data_out_12_), .unquautized_data_11_(
        data_out_11_), .unquautized_data_10_(data_out_10_), 
        .unquautized_data_9_(data_out_9_), .unquautized_data_8_(data_out_8_), 
        .unquautized_data_7_(data_out_7_), .unquautized_data_6_(data_out_6_), 
        .unquautized_data_5_(data_out_5_), .unquautized_data_4_(data_out_4_)
         );
  NBUFFX2_HVT U1 ( .A(sram_wdata_e[7]), .Y(sram_wdata_f[7]) );
  NBUFFX2_HVT U2 ( .A(sram_wdata_e[6]), .Y(sram_wdata_f[6]) );
  NBUFFX2_HVT U3 ( .A(sram_wdata_e[1]), .Y(sram_wdata_f[1]) );
  NBUFFX2_HVT U4 ( .A(sram_wdata_e[3]), .Y(sram_wdata_f[3]) );
  NBUFFX2_HVT U5 ( .A(sram_wdata_e[4]), .Y(sram_wdata_f[4]) );
  NBUFFX2_HVT U6 ( .A(sram_wdata_e[0]), .Y(sram_wdata_f[0]) );
  NBUFFX2_HVT U7 ( .A(sram_wdata_e[5]), .Y(sram_wdata_f[5]) );
  NBUFFX2_HVT U8 ( .A(sram_wdata_e[2]), .Y(sram_wdata_f[2]) );
  NBUFFX2_HVT U9 ( .A(sram_bytemask_e[3]), .Y(sram_bytemask_f[3]) );
  NBUFFX2_HVT U10 ( .A(sram_waddr_e[1]), .Y(sram_waddr_f[1]) );
  NBUFFX2_HVT U11 ( .A(sram_waddr_e[0]), .Y(sram_waddr_f[0]) );
  NBUFFX2_HVT U12 ( .A(sram_bytemask_e[1]), .Y(sram_bytemask_f[1]) );
  NBUFFX2_HVT U13 ( .A(sram_bytemask_e[0]), .Y(sram_bytemask_f[0]) );
  NBUFFX2_HVT U14 ( .A(sram_bytemask_e[2]), .Y(sram_bytemask_f[2]) );
endmodule


module lenet ( clk, srstn, conv_start, sram_rdata_a0, sram_rdata_a1, 
        sram_rdata_a2, sram_rdata_a3, sram_rdata_a4, sram_rdata_a5, 
        sram_rdata_a6, sram_rdata_a7, sram_rdata_a8, sram_rdata_b0, 
        sram_rdata_b1, sram_rdata_b2, sram_rdata_b3, sram_rdata_b4, 
        sram_rdata_b5, sram_rdata_b6, sram_rdata_b7, sram_rdata_b8, 
        conv_sram_rdata_weight, conv_sram_raddr_weight, sram_raddr_a0, 
        sram_raddr_a1, sram_raddr_a2, sram_raddr_a3, sram_raddr_a4, 
        sram_raddr_a5, sram_raddr_a6, sram_raddr_a7, sram_raddr_a8, 
        sram_write_enable_b0, sram_write_enable_b1, sram_write_enable_b2, 
        sram_write_enable_b3, sram_write_enable_b4, sram_write_enable_b5, 
        sram_write_enable_b6, sram_write_enable_b7, sram_write_enable_b8, 
        sram_bytemask_b, sram_waddr_b, sram_wdata_b, sram_raddr_b0, 
        sram_raddr_b1, sram_raddr_b2, sram_raddr_b3, sram_raddr_b4, 
        sram_raddr_b5, sram_raddr_b6, sram_raddr_b7, sram_raddr_b8, 
        sram_write_enable_c0, sram_write_enable_c1, sram_write_enable_c2, 
        sram_write_enable_c3, sram_write_enable_c4, sram_bytemask_c, 
        sram_waddr_c, sram_wdata_c, sram_write_enable_d0, sram_write_enable_d1, 
        sram_write_enable_d2, sram_write_enable_d3, sram_write_enable_d4, 
        sram_bytemask_d, sram_waddr_d, sram_wdata_d, conv_done, mem_sel, 
        sram_rdata_c0, sram_rdata_c1, sram_rdata_c2, sram_rdata_c3, 
        sram_rdata_c4, sram_raddr_c0, sram_raddr_c1, sram_raddr_c2, 
        sram_raddr_c3, sram_raddr_c4, sram_rdata_d0, sram_rdata_d1, 
        sram_rdata_d2, sram_rdata_d3, sram_rdata_d4, sram_raddr_d0, 
        sram_raddr_d1, sram_raddr_d2, sram_raddr_d3, sram_raddr_d4, 
        sram_rdata_e0, sram_rdata_e1, sram_rdata_e2, sram_rdata_e3, 
        sram_rdata_e4, sram_raddr_e0, sram_raddr_e1, sram_raddr_e2, 
        sram_raddr_e3, sram_raddr_e4, sram_write_enable_e0, 
        sram_write_enable_e1, sram_write_enable_e2, sram_write_enable_e3, 
        sram_write_enable_e4, sram_bytemask_e, sram_waddr_e, sram_wdata_e, 
        sram_write_enable_f, sram_bytemask_f, sram_waddr_f, sram_wdata_f, 
        fc_sram_rdata_weight, fc_sram_raddr_weight, fc1_done, fc2_done );
  input [31:0] sram_rdata_a0;
  input [31:0] sram_rdata_a1;
  input [31:0] sram_rdata_a2;
  input [31:0] sram_rdata_a3;
  input [31:0] sram_rdata_a4;
  input [31:0] sram_rdata_a5;
  input [31:0] sram_rdata_a6;
  input [31:0] sram_rdata_a7;
  input [31:0] sram_rdata_a8;
  input [31:0] sram_rdata_b0;
  input [31:0] sram_rdata_b1;
  input [31:0] sram_rdata_b2;
  input [31:0] sram_rdata_b3;
  input [31:0] sram_rdata_b4;
  input [31:0] sram_rdata_b5;
  input [31:0] sram_rdata_b6;
  input [31:0] sram_rdata_b7;
  input [31:0] sram_rdata_b8;
  input [99:0] conv_sram_rdata_weight;
  output [16:0] conv_sram_raddr_weight;
  output [9:0] sram_raddr_a0;
  output [9:0] sram_raddr_a1;
  output [9:0] sram_raddr_a2;
  output [9:0] sram_raddr_a3;
  output [9:0] sram_raddr_a4;
  output [9:0] sram_raddr_a5;
  output [9:0] sram_raddr_a6;
  output [9:0] sram_raddr_a7;
  output [9:0] sram_raddr_a8;
  output [3:0] sram_bytemask_b;
  output [9:0] sram_waddr_b;
  output [7:0] sram_wdata_b;
  output [9:0] sram_raddr_b0;
  output [9:0] sram_raddr_b1;
  output [9:0] sram_raddr_b2;
  output [9:0] sram_raddr_b3;
  output [9:0] sram_raddr_b4;
  output [9:0] sram_raddr_b5;
  output [9:0] sram_raddr_b6;
  output [9:0] sram_raddr_b7;
  output [9:0] sram_raddr_b8;
  output [3:0] sram_bytemask_c;
  output [9:0] sram_waddr_c;
  output [7:0] sram_wdata_c;
  output [3:0] sram_bytemask_d;
  output [9:0] sram_waddr_d;
  output [7:0] sram_wdata_d;
  input [31:0] sram_rdata_c0;
  input [31:0] sram_rdata_c1;
  input [31:0] sram_rdata_c2;
  input [31:0] sram_rdata_c3;
  input [31:0] sram_rdata_c4;
  output [5:0] sram_raddr_c0;
  output [5:0] sram_raddr_c1;
  output [5:0] sram_raddr_c2;
  output [5:0] sram_raddr_c3;
  output [5:0] sram_raddr_c4;
  input [31:0] sram_rdata_d0;
  input [31:0] sram_rdata_d1;
  input [31:0] sram_rdata_d2;
  input [31:0] sram_rdata_d3;
  input [31:0] sram_rdata_d4;
  output [5:0] sram_raddr_d0;
  output [5:0] sram_raddr_d1;
  output [5:0] sram_raddr_d2;
  output [5:0] sram_raddr_d3;
  output [5:0] sram_raddr_d4;
  input [31:0] sram_rdata_e0;
  input [31:0] sram_rdata_e1;
  input [31:0] sram_rdata_e2;
  input [31:0] sram_rdata_e3;
  input [31:0] sram_rdata_e4;
  output [4:0] sram_raddr_e0;
  output [4:0] sram_raddr_e1;
  output [4:0] sram_raddr_e2;
  output [4:0] sram_raddr_e3;
  output [4:0] sram_raddr_e4;
  output [3:0] sram_bytemask_e;
  output [4:0] sram_waddr_e;
  output [7:0] sram_wdata_e;
  output [3:0] sram_bytemask_f;
  output [1:0] sram_waddr_f;
  output [7:0] sram_wdata_f;
  input [79:0] fc_sram_rdata_weight;
  output [14:0] fc_sram_raddr_weight;
  input clk, srstn, conv_start;
  output sram_write_enable_b0, sram_write_enable_b1, sram_write_enable_b2,
         sram_write_enable_b3, sram_write_enable_b4, sram_write_enable_b5,
         sram_write_enable_b6, sram_write_enable_b7, sram_write_enable_b8,
         sram_write_enable_c0, sram_write_enable_c1, sram_write_enable_c2,
         sram_write_enable_c3, sram_write_enable_c4, sram_write_enable_d0,
         sram_write_enable_d1, sram_write_enable_d2, sram_write_enable_d3,
         sram_write_enable_d4, conv_done, mem_sel, sram_write_enable_e0,
         sram_write_enable_e1, sram_write_enable_e2, sram_write_enable_e3,
         sram_write_enable_e4, sram_write_enable_f, fc1_done, fc2_done;


  conv_top conv_top ( .clk(clk), .srstn(srstn), .conv_start(conv_start), 
        .fc_done(fc2_done), .sram_rdata_a0(sram_rdata_a0), .sram_rdata_a1(
        sram_rdata_a1), .sram_rdata_a2(sram_rdata_a2), .sram_rdata_a3(
        sram_rdata_a3), .sram_rdata_a4(sram_rdata_a4), .sram_rdata_a5(
        sram_rdata_a5), .sram_rdata_a6(sram_rdata_a6), .sram_rdata_a7(
        sram_rdata_a7), .sram_rdata_a8(sram_rdata_a8), .sram_rdata_b0(
        sram_rdata_b0), .sram_rdata_b1(sram_rdata_b1), .sram_rdata_b2(
        sram_rdata_b2), .sram_rdata_b3(sram_rdata_b3), .sram_rdata_b4(
        sram_rdata_b4), .sram_rdata_b5(sram_rdata_b5), .sram_rdata_b6(
        sram_rdata_b6), .sram_rdata_b7(sram_rdata_b7), .sram_rdata_b8(
        sram_rdata_b8), .sram_rdata_weight(conv_sram_rdata_weight), 
        .sram_raddr_weight(conv_sram_raddr_weight), .sram_raddr_a0(
        sram_raddr_a0), .sram_raddr_a1(sram_raddr_a1), .sram_raddr_a2(
        sram_raddr_a2), .sram_raddr_a3(sram_raddr_a3), .sram_raddr_a4(
        sram_raddr_a4), .sram_raddr_a5(sram_raddr_a5), .sram_raddr_a6(
        sram_raddr_a6), .sram_raddr_a7(sram_raddr_a7), .sram_raddr_a8(
        sram_raddr_a8), .sram_write_enable_b0(sram_write_enable_b0), 
        .sram_write_enable_b1(sram_write_enable_b1), .sram_write_enable_b2(
        sram_write_enable_b2), .sram_write_enable_b3(sram_write_enable_b3), 
        .sram_write_enable_b4(sram_write_enable_b4), .sram_write_enable_b5(
        sram_write_enable_b5), .sram_write_enable_b6(sram_write_enable_b6), 
        .sram_write_enable_b7(sram_write_enable_b7), .sram_write_enable_b8(
        sram_write_enable_b8), .sram_bytemask_b(sram_bytemask_b), 
        .sram_waddr_b(sram_waddr_b), .sram_wdata_b(sram_wdata_b), 
        .sram_raddr_b0(sram_raddr_b0), .sram_raddr_b1(sram_raddr_b1), 
        .sram_raddr_b2(sram_raddr_b2), .sram_raddr_b3(sram_raddr_b3), 
        .sram_raddr_b4(sram_raddr_b4), .sram_raddr_b5(sram_raddr_b5), 
        .sram_raddr_b6(sram_raddr_b6), .sram_raddr_b7(sram_raddr_b7), 
        .sram_raddr_b8(sram_raddr_b8), .sram_write_enable_c0(
        sram_write_enable_c0), .sram_write_enable_c1(sram_write_enable_c1), 
        .sram_write_enable_c2(sram_write_enable_c2), .sram_write_enable_c3(
        sram_write_enable_c3), .sram_write_enable_c4(sram_write_enable_c4), 
        .sram_bytemask_c(sram_bytemask_c), .sram_waddr_c(sram_waddr_c), 
        .sram_wdata_c(sram_wdata_c), .sram_write_enable_d0(
        sram_write_enable_d0), .sram_write_enable_d1(sram_write_enable_d1), 
        .sram_write_enable_d2(sram_write_enable_d2), .sram_write_enable_d3(
        sram_write_enable_d3), .sram_write_enable_d4(sram_write_enable_d4), 
        .sram_bytemask_d(sram_bytemask_d), .sram_waddr_d(sram_waddr_d), 
        .sram_wdata_d(sram_wdata_d), .conv_done(conv_done), .mem_sel(mem_sel)
         );
  fc_top fc_top ( .clk(clk), .srstn(srstn), .conv_done(conv_done), .mem_sel(
        mem_sel), .sram_rdata_c0(sram_rdata_c0), .sram_rdata_c1(sram_rdata_c1), 
        .sram_rdata_c2(sram_rdata_c2), .sram_rdata_c3(sram_rdata_c3), 
        .sram_rdata_c4(sram_rdata_c4), .sram_raddr_c0(sram_raddr_c0), 
        .sram_raddr_c1(sram_raddr_c1), .sram_raddr_c2(sram_raddr_c2), 
        .sram_raddr_c3(sram_raddr_c3), .sram_raddr_c4(sram_raddr_c4), 
        .sram_rdata_d0(sram_rdata_d0), .sram_rdata_d1(sram_rdata_d1), 
        .sram_rdata_d2(sram_rdata_d2), .sram_rdata_d3(sram_rdata_d3), 
        .sram_rdata_d4(sram_rdata_d4), .sram_raddr_d0(sram_raddr_d0), 
        .sram_raddr_d1(sram_raddr_d1), .sram_raddr_d2(sram_raddr_d2), 
        .sram_raddr_d3(sram_raddr_d3), .sram_raddr_d4(sram_raddr_d4), 
        .sram_rdata_e0(sram_rdata_e0), .sram_rdata_e1(sram_rdata_e1), 
        .sram_rdata_e2(sram_rdata_e2), .sram_rdata_e3(sram_rdata_e3), 
        .sram_rdata_e4(sram_rdata_e4), .sram_raddr_e0(sram_raddr_e0), 
        .sram_raddr_e1(sram_raddr_e1), .sram_raddr_e2(sram_raddr_e2), 
        .sram_raddr_e3(sram_raddr_e3), .sram_raddr_e4(sram_raddr_e4), 
        .sram_write_enable_e0(sram_write_enable_e0), .sram_write_enable_e1(
        sram_write_enable_e1), .sram_write_enable_e2(sram_write_enable_e2), 
        .sram_write_enable_e3(sram_write_enable_e3), .sram_write_enable_e4(
        sram_write_enable_e4), .sram_bytemask_e(sram_bytemask_e), 
        .sram_waddr_e(sram_waddr_e), .sram_wdata_e(sram_wdata_e), 
        .sram_write_enable_f(sram_write_enable_f), .sram_bytemask_f(
        sram_bytemask_f), .sram_waddr_f(sram_waddr_f), .sram_wdata_f(
        sram_wdata_f), .sram_rdata_weight(fc_sram_rdata_weight), 
        .sram_raddr_weight(fc_sram_raddr_weight), .fc1_done(fc1_done), 
        .fc2_done(fc2_done) );
endmodule

